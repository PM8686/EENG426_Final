magic
tech sky130l
timestamp 1731220607
<< m1 >>
rect 392 3511 396 3535
rect 536 3511 540 3535
rect 680 3511 684 3535
rect 944 3511 948 3535
rect 1168 3511 1172 3535
rect 1304 3511 1308 3535
rect 1416 3511 1420 3535
rect 1536 3511 1540 3535
rect 1968 3523 1972 3547
rect 2056 3523 2060 3547
rect 2144 3523 2148 3547
rect 2232 3523 2236 3547
rect 2320 3523 2324 3547
rect 2408 3523 2412 3547
rect 2496 3523 2500 3547
rect 2672 3523 2676 3547
rect 2760 3523 2764 3547
rect 2848 3523 2852 3547
rect 2936 3523 2940 3547
rect 3024 3523 3028 3547
rect 3112 3523 3116 3547
rect 3200 3523 3204 3547
rect 3288 3523 3292 3547
rect 256 3471 260 3495
rect 608 3471 612 3495
rect 1040 3475 1044 3495
rect 1296 3475 1300 3495
rect 1416 3475 1420 3495
rect 1520 3475 1524 3495
rect 1984 3475 1988 3499
rect 3032 3475 3036 3499
rect 408 3375 412 3399
rect 576 3375 580 3399
rect 752 3375 756 3399
rect 1472 3375 1476 3399
rect 2064 3371 2068 3395
rect 2624 3371 2628 3395
rect 3016 3371 3020 3395
rect 328 3331 332 3351
rect 472 3331 476 3351
rect 632 3331 636 3351
rect 960 3331 964 3351
rect 1064 3331 1068 3351
rect 1352 3327 1356 3351
rect 1504 3327 1508 3351
rect 2336 3331 2340 3351
rect 2472 3331 2476 3351
rect 368 3227 372 3251
rect 504 3227 508 3251
rect 656 3227 660 3251
rect 816 3227 820 3251
rect 1512 3227 1516 3251
rect 2056 3227 2060 3251
rect 2976 3227 2980 3251
rect 3472 3227 3476 3251
rect 512 3187 516 3207
rect 632 3187 636 3207
rect 752 3187 756 3207
rect 1024 3187 1028 3207
rect 1192 3187 1196 3207
rect 1480 3183 1484 3207
rect 2424 3191 2428 3211
rect 3280 3191 3284 3223
rect 3296 3187 3300 3211
rect 544 3083 548 3107
rect 632 3083 636 3107
rect 728 3083 732 3107
rect 840 3083 844 3107
rect 960 3083 964 3107
rect 1512 3083 1516 3107
rect 2072 3087 2076 3111
rect 3032 3087 3036 3111
rect 3184 3087 3188 3111
rect 3336 3087 3340 3111
rect 312 3039 316 3059
rect 392 3039 396 3059
rect 480 3039 484 3059
rect 568 3039 572 3059
rect 656 3039 660 3059
rect 744 3039 748 3059
rect 832 3039 836 3059
rect 920 3039 924 3059
rect 1008 3039 1012 3059
rect 1184 3039 1188 3059
rect 1272 3039 1276 3059
rect 1360 3039 1364 3059
rect 1368 3035 1372 3079
rect 1712 3039 1716 3059
rect 1808 3039 1812 3083
rect 2376 3039 2380 3059
rect 2664 3039 2668 3083
rect 2672 3035 2676 3059
rect 3024 3039 3028 3059
rect 1704 2931 1708 2955
rect 2856 2935 2860 2959
rect 1544 2895 1548 2915
rect 2760 2883 2764 2903
rect 2960 2883 2964 2903
rect 3120 2883 3124 2903
rect 3280 2883 3284 2903
rect 208 2779 212 2807
rect 296 2791 300 2815
rect 960 2791 964 2815
rect 1208 2791 1212 2815
rect 280 2755 284 2775
rect 376 2755 380 2775
rect 640 2755 644 2775
rect 776 2755 780 2775
rect 888 2755 892 2787
rect 1976 2779 1980 2803
rect 2064 2779 2068 2803
rect 2152 2779 2156 2803
rect 2240 2779 2244 2803
rect 2328 2779 2332 2803
rect 1032 2755 1036 2775
rect 1280 2755 1284 2775
rect 1392 2755 1396 2775
rect 1504 2755 1508 2775
rect 1608 2755 1612 2775
rect 1712 2755 1716 2775
rect 2416 2771 2420 2803
rect 2680 2779 2684 2803
rect 2784 2779 2788 2803
rect 2896 2779 2900 2803
rect 3024 2779 3028 2803
rect 2112 2731 2116 2751
rect 2240 2731 2244 2751
rect 2248 2727 2252 2767
rect 2904 2727 2908 2751
rect 3336 2731 3340 2775
rect 2400 2631 2404 2655
rect 2624 2631 2628 2655
rect 2728 2631 2732 2655
rect 2840 2631 2844 2655
rect 2952 2631 2956 2655
rect 3064 2631 3068 2655
rect 336 2595 340 2615
rect 440 2595 444 2615
rect 1328 2595 1332 2615
rect 1528 2595 1532 2615
rect 2000 2591 2004 2611
rect 2184 2591 2188 2611
rect 2584 2591 2588 2611
rect 3152 2587 3156 2611
rect 3272 2535 3276 2611
rect 848 2495 852 2519
rect 1312 2495 1316 2519
rect 2568 2491 2572 2515
rect 2896 2491 2900 2515
rect 3048 2491 3052 2515
rect 408 2455 412 2475
rect 568 2391 572 2475
rect 696 2455 700 2475
rect 832 2455 836 2475
rect 840 2451 844 2491
rect 1312 2455 1316 2475
rect 1416 2455 1420 2475
rect 1520 2455 1524 2475
rect 1616 2455 1620 2475
rect 1712 2455 1716 2475
rect 1808 2455 1812 2475
rect 1960 2455 1964 2475
rect 2080 2455 2084 2475
rect 2216 2455 2220 2475
rect 3368 2455 3372 2487
rect 1040 2347 1044 2371
rect 1296 2347 1300 2371
rect 1424 2347 1428 2371
rect 2800 2347 2804 2371
rect 2960 2347 2964 2371
rect 3128 2347 3132 2371
rect 232 2307 236 2327
rect 496 2307 500 2327
rect 632 2307 636 2327
rect 752 2307 756 2343
rect 784 2251 788 2327
rect 888 2307 892 2327
rect 1000 2307 1004 2327
rect 2840 2307 2844 2327
rect 128 2191 132 2231
rect 1048 2207 1052 2231
rect 2440 2207 2444 2231
rect 208 2167 212 2187
rect 472 2167 476 2187
rect 608 2167 612 2187
rect 864 2167 868 2187
rect 1120 2163 1124 2187
rect 1256 2103 1260 2187
rect 2944 2171 2948 2191
rect 3200 2171 3204 2191
rect 208 2035 212 2075
rect 824 2059 828 2083
rect 936 2059 940 2083
rect 1048 2059 1052 2083
rect 1168 2059 1172 2083
rect 2232 2063 2236 2087
rect 2408 2063 2412 2087
rect 2496 2063 2500 2087
rect 2744 2063 2748 2087
rect 2912 2063 2916 2087
rect 3200 2055 3204 2103
rect 3296 2063 3300 2087
rect 528 2011 532 2031
rect 1296 2007 1300 2031
rect 2080 2023 2084 2043
rect 2464 2023 2468 2043
rect 288 1911 292 1935
rect 432 1891 436 1935
rect 1232 1911 1236 1935
rect 2392 1915 2396 1939
rect 320 1863 324 1887
rect 1040 1867 1044 1887
rect 1232 1867 1236 1887
rect 1392 1867 1396 1887
rect 1552 1867 1556 1887
rect 2048 1879 2052 1899
rect 2056 1875 2060 1907
rect 2608 1903 2612 1939
rect 2808 1915 2812 1939
rect 2992 1915 2996 1939
rect 3160 1915 3164 1939
rect 3328 1915 3332 1939
rect 2248 1879 2252 1899
rect 2392 1879 2396 1899
rect 2696 1879 2700 1899
rect 3016 1879 3020 1899
rect 3160 1879 3164 1899
rect 408 1767 412 1791
rect 416 1727 420 1747
rect 864 1727 868 1747
rect 1208 1727 1212 1747
rect 1320 1727 1324 1747
rect 1624 1727 1628 1747
rect 2008 1735 2012 1771
rect 2432 1759 2436 1799
rect 2632 1775 2636 1799
rect 3336 1775 3340 1859
rect 2224 1675 2228 1755
rect 2528 1735 2532 1755
rect 2912 1735 2916 1755
rect 880 1623 884 1647
rect 1416 1603 1420 1639
rect 2024 1631 2028 1655
rect 2144 1631 2148 1655
rect 2392 1631 2396 1655
rect 328 1579 332 1599
rect 440 1579 444 1599
rect 712 1579 716 1599
rect 1000 1579 1004 1599
rect 1480 1579 1484 1599
rect 2112 1523 2116 1607
rect 2360 1583 2364 1607
rect 2680 1587 2684 1607
rect 2864 1587 2868 1607
rect 3024 1587 3028 1607
rect 208 1475 212 1499
rect 1336 1475 1340 1499
rect 2016 1479 2020 1503
rect 2336 1479 2340 1503
rect 2496 1479 2500 1503
rect 2976 1479 2980 1503
rect 3144 1479 3148 1503
rect 208 1431 212 1451
rect 352 1431 356 1451
rect 616 1431 620 1451
rect 728 1431 732 1471
rect 872 1431 876 1451
rect 984 1431 988 1451
rect 1464 1431 1468 1451
rect 1592 1375 1596 1451
rect 1704 1431 1708 1451
rect 1808 1431 1812 1475
rect 2288 1435 2292 1455
rect 2824 1435 2828 1455
rect 2944 1435 2948 1455
rect 3112 1435 3116 1455
rect 3280 1435 3284 1455
rect 208 1331 212 1355
rect 1496 1331 1500 1355
rect 2256 1327 2260 1351
rect 2608 1327 2612 1351
rect 2928 1327 2932 1351
rect 3072 1327 3076 1351
rect 3216 1327 3220 1351
rect 208 1287 212 1307
rect 640 1287 644 1307
rect 832 1287 836 1307
rect 984 1287 988 1327
rect 1328 1287 1332 1307
rect 1480 1287 1484 1307
rect 1632 1287 1636 1307
rect 1752 1287 1756 1327
rect 3352 1315 3356 1351
rect 2432 1291 2436 1311
rect 2816 1291 2820 1311
rect 3288 1287 3292 1311
rect 288 1183 292 1207
rect 472 1183 476 1207
rect 1104 1183 1108 1207
rect 1240 1183 1244 1207
rect 1376 1183 1380 1207
rect 1520 1183 1524 1207
rect 2624 1187 2628 1211
rect 3056 1187 3060 1211
rect 3200 1187 3204 1211
rect 704 1143 708 1163
rect 824 1143 828 1179
rect 1008 1143 1012 1163
rect 1168 1143 1172 1163
rect 1336 1143 1340 1163
rect 1528 1143 1532 1163
rect 2176 1147 2180 1167
rect 2512 1147 2516 1183
rect 2720 1147 2724 1167
rect 2896 1147 2900 1167
rect 3056 1147 3060 1167
rect 320 1039 324 1063
rect 432 1039 436 1063
rect 544 1039 548 1063
rect 552 1019 556 1063
rect 936 1039 940 1063
rect 1032 1039 1036 1063
rect 1240 1039 1244 1063
rect 1400 1039 1404 1063
rect 2400 1035 2404 1059
rect 2856 1035 2860 1059
rect 1624 995 1628 1015
rect 2152 995 2156 1015
rect 2272 995 2276 1015
rect 2392 995 2396 1015
rect 2664 995 2668 1015
rect 2824 995 2828 1015
rect 2968 995 2972 1015
rect 3264 995 3268 1031
rect 3288 991 3292 1015
rect 456 891 460 915
rect 696 891 700 915
rect 840 891 844 915
rect 1520 891 1524 915
rect 2016 891 2020 915
rect 2624 891 2628 915
rect 3016 891 3020 915
rect 992 851 996 887
rect 2264 855 2268 875
rect 2760 851 2764 875
rect 3160 855 3164 875
rect 528 751 532 775
rect 816 751 820 775
rect 1120 751 1124 775
rect 448 711 452 731
rect 1000 711 1004 747
rect 1432 735 1436 775
rect 1592 751 1596 775
rect 2128 755 2132 779
rect 2792 755 2796 779
rect 2960 755 2964 771
rect 3312 755 3316 779
rect 1232 711 1236 731
rect 1520 711 1524 731
rect 2176 715 2180 735
rect 2368 715 2372 735
rect 3104 715 3108 735
rect 200 595 204 627
rect 768 611 772 635
rect 1024 611 1028 635
rect 1336 611 1340 635
rect 208 571 212 591
rect 416 571 420 591
rect 1000 567 1004 607
rect 1664 571 1668 591
rect 2264 571 2268 591
rect 2352 571 2356 591
rect 2440 571 2444 591
rect 2536 571 2540 607
rect 2640 571 2644 591
rect 3256 571 3260 591
rect 200 451 204 483
rect 1344 467 1348 491
rect 3088 467 3092 491
rect 3344 467 3348 491
rect 208 427 212 447
rect 376 427 380 447
rect 664 371 668 447
rect 760 427 764 447
rect 1664 427 1668 447
rect 2304 431 2308 451
rect 2400 431 2404 451
rect 2512 431 2516 451
rect 2632 431 2636 451
rect 2944 431 2948 451
rect 3408 375 3412 451
rect 208 327 212 351
rect 1576 327 1580 351
rect 2280 331 2284 355
rect 2392 331 2396 355
rect 2520 331 2524 355
rect 2744 331 2748 355
rect 3288 331 3292 355
rect 3456 331 3460 355
rect 560 311 568 314
rect 304 291 308 311
rect 560 310 572 311
rect 560 291 564 310
rect 736 291 740 311
rect 1024 287 1028 311
rect 1312 291 1316 311
rect 1424 291 1428 311
rect 1696 291 1700 311
rect 1808 291 1812 307
rect 2160 291 2164 327
rect 2632 287 2636 307
rect 3216 283 3220 307
rect 480 183 484 207
rect 1024 183 1028 207
rect 1288 183 1292 207
rect 1992 187 1996 211
rect 2136 187 2140 211
rect 240 123 244 143
rect 328 123 332 143
rect 416 123 420 143
rect 504 123 508 143
rect 592 123 596 143
rect 680 123 684 143
rect 768 123 772 143
rect 1040 119 1044 143
rect 1384 123 1388 143
rect 1472 123 1476 143
rect 1480 119 1484 151
rect 2688 147 2692 203
rect 1968 123 1972 143
rect 2048 123 2052 143
rect 2136 123 2140 143
rect 2224 123 2228 143
rect 2312 123 2316 143
rect 2408 123 2412 143
rect 2712 123 2716 143
rect 2824 123 2828 143
rect 2904 123 2908 143
rect 3000 123 3004 143
rect 3096 123 3100 143
rect 3192 123 3196 143
rect 3288 123 3292 143
<< m2c >>
rect 268 3639 272 3643
rect 356 3639 360 3643
rect 444 3639 448 3643
rect 532 3639 536 3643
rect 620 3639 624 3643
rect 280 3583 284 3587
rect 1968 3547 1972 3551
rect 392 3535 396 3539
rect 536 3535 540 3539
rect 680 3535 684 3539
rect 944 3535 948 3539
rect 1168 3535 1172 3539
rect 1304 3535 1308 3539
rect 1416 3535 1420 3539
rect 1536 3535 1540 3539
rect 2056 3547 2060 3551
rect 2144 3547 2148 3551
rect 2232 3547 2236 3551
rect 2320 3547 2324 3551
rect 2408 3547 2412 3551
rect 2496 3547 2500 3551
rect 2672 3547 2676 3551
rect 2760 3547 2764 3551
rect 2848 3547 2852 3551
rect 2936 3547 2940 3551
rect 3024 3547 3028 3551
rect 3112 3547 3116 3551
rect 3200 3547 3204 3551
rect 3288 3547 3292 3551
rect 1924 3519 1928 3523
rect 1968 3519 1972 3523
rect 2012 3519 2016 3523
rect 2056 3519 2060 3523
rect 2100 3519 2104 3523
rect 2144 3519 2148 3523
rect 2188 3519 2192 3523
rect 2232 3519 2236 3523
rect 2276 3519 2280 3523
rect 2320 3519 2324 3523
rect 2364 3519 2368 3523
rect 2408 3519 2412 3523
rect 2452 3519 2456 3523
rect 2496 3519 2500 3523
rect 2540 3519 2544 3523
rect 2628 3519 2632 3523
rect 2672 3519 2676 3523
rect 2716 3519 2720 3523
rect 2760 3519 2764 3523
rect 2804 3519 2808 3523
rect 2848 3519 2852 3523
rect 2892 3519 2896 3523
rect 2936 3519 2940 3523
rect 2980 3519 2984 3523
rect 3024 3519 3028 3523
rect 3068 3519 3072 3523
rect 3112 3519 3116 3523
rect 3156 3519 3160 3523
rect 3200 3519 3204 3523
rect 3244 3519 3248 3523
rect 3288 3519 3292 3523
rect 3332 3519 3336 3523
rect 284 3507 288 3511
rect 392 3507 396 3511
rect 436 3507 440 3511
rect 536 3507 540 3511
rect 580 3507 584 3511
rect 680 3507 684 3511
rect 724 3507 728 3511
rect 860 3507 864 3511
rect 944 3507 948 3511
rect 988 3507 992 3511
rect 1116 3507 1120 3511
rect 1168 3507 1172 3511
rect 1236 3507 1240 3511
rect 1304 3507 1308 3511
rect 1348 3507 1352 3511
rect 1416 3507 1420 3511
rect 1460 3507 1464 3511
rect 1536 3507 1540 3511
rect 1580 3507 1584 3511
rect 1940 3499 1944 3503
rect 1984 3499 1988 3503
rect 2044 3499 2048 3503
rect 2164 3499 2168 3503
rect 2292 3499 2296 3503
rect 2420 3499 2424 3503
rect 2556 3499 2560 3503
rect 2692 3499 2696 3503
rect 2828 3499 2832 3503
rect 2972 3499 2976 3503
rect 3032 3499 3036 3503
rect 3116 3499 3120 3503
rect 212 3495 216 3499
rect 256 3495 260 3499
rect 380 3495 384 3499
rect 548 3495 552 3499
rect 608 3495 612 3499
rect 708 3495 712 3499
rect 860 3495 864 3499
rect 996 3495 1000 3499
rect 1040 3495 1044 3499
rect 1124 3495 1128 3499
rect 1244 3495 1248 3499
rect 1296 3495 1300 3499
rect 1364 3495 1368 3499
rect 1416 3495 1420 3499
rect 1484 3495 1488 3499
rect 1520 3495 1524 3499
rect 1604 3495 1608 3499
rect 256 3467 260 3471
rect 1040 3471 1044 3475
rect 1296 3471 1300 3475
rect 1416 3471 1420 3475
rect 1520 3471 1524 3475
rect 1984 3471 1988 3475
rect 3032 3471 3036 3475
rect 608 3467 612 3471
rect 408 3399 412 3403
rect 576 3399 580 3403
rect 752 3399 756 3403
rect 1472 3399 1476 3403
rect 2064 3395 2068 3399
rect 172 3371 176 3375
rect 292 3371 296 3375
rect 408 3371 412 3375
rect 452 3371 456 3375
rect 576 3371 580 3375
rect 620 3371 624 3375
rect 752 3371 756 3375
rect 796 3371 800 3375
rect 972 3371 976 3375
rect 1148 3371 1152 3375
rect 1332 3371 1336 3375
rect 1472 3371 1476 3375
rect 1516 3371 1520 3375
rect 2624 3395 2628 3399
rect 3016 3395 3020 3399
rect 1948 3367 1952 3371
rect 2064 3367 2068 3371
rect 2108 3367 2112 3371
rect 2260 3367 2264 3371
rect 2404 3367 2408 3371
rect 2540 3367 2544 3371
rect 2624 3367 2628 3371
rect 2668 3367 2672 3371
rect 2796 3367 2800 3371
rect 2924 3367 2928 3371
rect 3016 3367 3020 3371
rect 3060 3367 3064 3371
rect 236 3353 240 3357
rect 328 3351 332 3355
rect 396 3351 400 3355
rect 472 3351 476 3355
rect 564 3351 568 3355
rect 632 3351 636 3355
rect 724 3351 728 3355
rect 884 3351 888 3355
rect 960 3351 964 3355
rect 1028 3351 1032 3355
rect 1064 3351 1068 3355
rect 1172 3351 1176 3355
rect 1308 3351 1312 3355
rect 1352 3351 1356 3355
rect 1444 3351 1448 3355
rect 1504 3351 1508 3355
rect 1588 3351 1592 3355
rect 1924 3351 1928 3355
rect 2076 3351 2080 3355
rect 2236 3351 2240 3355
rect 2336 3351 2340 3355
rect 2396 3351 2400 3355
rect 2472 3351 2476 3355
rect 2564 3351 2568 3355
rect 2732 3351 2736 3355
rect 2908 3351 2912 3355
rect 3084 3351 3088 3355
rect 328 3327 332 3331
rect 472 3327 476 3331
rect 632 3327 636 3331
rect 960 3327 964 3331
rect 1064 3327 1068 3331
rect 1352 3323 1356 3327
rect 2336 3327 2340 3331
rect 2472 3327 2476 3331
rect 1504 3323 1508 3327
rect 368 3251 372 3255
rect 504 3251 508 3255
rect 656 3251 660 3255
rect 816 3251 820 3255
rect 1512 3251 1516 3255
rect 2056 3251 2060 3255
rect 2976 3251 2980 3255
rect 3472 3251 3476 3255
rect 292 3223 296 3227
rect 368 3223 372 3227
rect 412 3223 416 3227
rect 504 3223 508 3227
rect 548 3223 552 3227
rect 656 3223 660 3227
rect 700 3223 704 3227
rect 816 3223 820 3227
rect 860 3223 864 3227
rect 1028 3223 1032 3227
rect 1204 3223 1208 3227
rect 1380 3223 1384 3227
rect 1512 3223 1516 3227
rect 1556 3223 1560 3227
rect 1924 3223 1928 3227
rect 2056 3223 2060 3227
rect 2100 3223 2104 3227
rect 2300 3223 2304 3227
rect 2492 3223 2496 3227
rect 2676 3223 2680 3227
rect 2852 3223 2856 3227
rect 2976 3223 2980 3227
rect 3020 3223 3024 3227
rect 3188 3223 3192 3227
rect 3280 3223 3284 3227
rect 3356 3223 3360 3227
rect 3472 3223 3476 3227
rect 3516 3223 3520 3227
rect 1924 3211 1928 3215
rect 2116 3211 2120 3215
rect 2332 3211 2336 3215
rect 2424 3211 2428 3215
rect 2540 3211 2544 3215
rect 2732 3211 2736 3215
rect 2908 3211 2912 3215
rect 3068 3211 3072 3215
rect 3228 3211 3232 3215
rect 460 3207 464 3211
rect 512 3207 516 3211
rect 580 3207 584 3211
rect 632 3207 636 3211
rect 700 3207 704 3211
rect 752 3207 756 3211
rect 828 3207 832 3211
rect 964 3207 968 3211
rect 1024 3207 1028 3211
rect 1108 3207 1112 3211
rect 1192 3207 1196 3211
rect 1260 3207 1264 3211
rect 1412 3207 1416 3211
rect 1480 3207 1484 3211
rect 1564 3207 1568 3211
rect 512 3183 516 3187
rect 632 3183 636 3187
rect 752 3183 756 3187
rect 1024 3183 1028 3187
rect 1192 3183 1196 3187
rect 2424 3187 2428 3191
rect 3280 3187 3284 3191
rect 3296 3211 3300 3215
rect 3380 3211 3384 3215
rect 3516 3211 3520 3215
rect 3296 3183 3300 3187
rect 1480 3179 1484 3183
rect 2552 3155 2556 3159
rect 2920 3155 2924 3159
rect 3528 3155 3532 3159
rect 1424 3151 1428 3155
rect 2072 3111 2076 3115
rect 544 3107 548 3111
rect 632 3107 636 3111
rect 728 3107 732 3111
rect 840 3107 844 3111
rect 960 3107 964 3111
rect 1512 3107 1516 3111
rect 3032 3111 3036 3115
rect 3184 3111 3188 3115
rect 3336 3111 3340 3115
rect 1808 3083 1812 3087
rect 1924 3083 1928 3087
rect 2072 3083 2076 3087
rect 2116 3083 2120 3087
rect 2332 3083 2336 3087
rect 2540 3083 2544 3087
rect 2664 3083 2668 3087
rect 2732 3083 2736 3087
rect 2908 3083 2912 3087
rect 3032 3083 3036 3087
rect 3076 3083 3080 3087
rect 3184 3083 3188 3087
rect 3228 3083 3232 3087
rect 3336 3083 3340 3087
rect 3380 3083 3384 3087
rect 3516 3083 3520 3087
rect 500 3079 504 3083
rect 544 3079 548 3083
rect 588 3079 592 3083
rect 632 3079 636 3083
rect 676 3079 680 3083
rect 728 3079 732 3083
rect 772 3079 776 3083
rect 840 3079 844 3083
rect 884 3079 888 3083
rect 960 3079 964 3083
rect 1004 3079 1008 3083
rect 1132 3079 1136 3083
rect 1268 3079 1272 3083
rect 1368 3079 1372 3083
rect 1412 3079 1416 3083
rect 1512 3079 1516 3083
rect 1556 3079 1560 3083
rect 180 3059 184 3063
rect 268 3059 272 3063
rect 312 3059 316 3063
rect 356 3059 360 3063
rect 392 3059 396 3063
rect 444 3059 448 3063
rect 480 3059 484 3063
rect 532 3059 536 3063
rect 568 3059 572 3063
rect 620 3059 624 3063
rect 656 3059 660 3063
rect 708 3059 712 3063
rect 744 3059 748 3063
rect 796 3059 800 3063
rect 832 3059 836 3063
rect 884 3059 888 3063
rect 920 3059 924 3063
rect 972 3059 976 3063
rect 1008 3059 1012 3063
rect 1060 3059 1064 3063
rect 1148 3059 1152 3063
rect 1184 3059 1188 3063
rect 1236 3059 1240 3063
rect 1272 3059 1276 3063
rect 1324 3059 1328 3063
rect 1360 3059 1364 3063
rect 312 3035 316 3039
rect 392 3035 396 3039
rect 480 3035 484 3039
rect 568 3035 572 3039
rect 656 3035 660 3039
rect 744 3035 748 3039
rect 832 3035 836 3039
rect 920 3035 924 3039
rect 1008 3035 1012 3039
rect 1184 3035 1188 3039
rect 1272 3035 1276 3039
rect 1360 3035 1364 3039
rect 1412 3059 1416 3063
rect 1500 3059 1504 3063
rect 1588 3059 1592 3063
rect 1676 3059 1680 3063
rect 1712 3059 1716 3063
rect 1764 3059 1768 3063
rect 1712 3035 1716 3039
rect 2284 3059 2288 3063
rect 2376 3059 2380 3063
rect 2452 3059 2456 3063
rect 2620 3059 2624 3063
rect 1808 3035 1812 3039
rect 2376 3035 2380 3039
rect 2664 3035 2668 3039
rect 2672 3059 2676 3063
rect 2780 3059 2784 3063
rect 2948 3059 2952 3063
rect 3024 3059 3028 3063
rect 3116 3059 3120 3063
rect 3024 3035 3028 3039
rect 1368 3031 1372 3035
rect 2672 3031 2676 3035
rect 2856 2959 2860 2963
rect 1704 2955 1708 2959
rect 2276 2931 2280 2935
rect 2500 2931 2504 2935
rect 2708 2931 2712 2935
rect 2856 2931 2860 2935
rect 2900 2931 2904 2935
rect 3068 2931 3072 2935
rect 3228 2931 3232 2935
rect 3380 2931 3384 2935
rect 3516 2931 3520 2935
rect 1444 2927 1448 2931
rect 1556 2927 1560 2931
rect 1668 2927 1672 2931
rect 1704 2927 1708 2931
rect 1764 2927 1768 2931
rect 1388 2917 1392 2921
rect 1500 2915 1504 2919
rect 1544 2915 1548 2919
rect 1612 2915 1616 2919
rect 1732 2915 1736 2919
rect 2268 2903 2272 2907
rect 2492 2903 2496 2907
rect 2700 2903 2704 2907
rect 2760 2903 2764 2907
rect 2884 2903 2888 2907
rect 2960 2903 2964 2907
rect 3052 2903 3056 2907
rect 3120 2903 3124 2907
rect 3212 2903 3216 2907
rect 3280 2903 3284 2907
rect 3364 2903 3368 2907
rect 3516 2903 3520 2907
rect 1544 2891 1548 2895
rect 2760 2879 2764 2883
rect 2960 2879 2964 2883
rect 3120 2879 3124 2883
rect 3280 2879 3284 2883
rect 1400 2859 1404 2863
rect 3528 2847 3532 2851
rect 296 2815 300 2819
rect 208 2807 212 2811
rect 172 2787 176 2791
rect 960 2815 964 2819
rect 260 2787 264 2791
rect 296 2787 300 2791
rect 348 2787 352 2791
rect 436 2787 440 2791
rect 524 2787 528 2791
rect 636 2787 640 2791
rect 764 2789 768 2793
rect 1208 2815 1212 2819
rect 1976 2803 1980 2807
rect 888 2787 892 2791
rect 900 2787 904 2791
rect 960 2787 964 2791
rect 1036 2787 1040 2791
rect 1172 2787 1176 2791
rect 1208 2787 1212 2791
rect 1300 2787 1304 2791
rect 1420 2787 1424 2791
rect 1540 2789 1544 2793
rect 1660 2787 1664 2791
rect 1764 2787 1768 2791
rect 208 2775 212 2779
rect 220 2775 224 2779
rect 280 2775 284 2779
rect 324 2775 328 2779
rect 376 2775 380 2779
rect 444 2775 448 2779
rect 580 2775 584 2779
rect 640 2775 644 2779
rect 716 2775 720 2779
rect 776 2775 780 2779
rect 852 2775 856 2779
rect 280 2751 284 2755
rect 376 2751 380 2755
rect 640 2751 644 2755
rect 776 2751 780 2755
rect 2064 2803 2068 2807
rect 2152 2803 2156 2807
rect 2240 2803 2244 2807
rect 2328 2803 2332 2807
rect 2416 2803 2420 2807
rect 988 2775 992 2779
rect 1032 2775 1036 2779
rect 1116 2775 1120 2779
rect 1236 2775 1240 2779
rect 1280 2775 1284 2779
rect 1348 2775 1352 2779
rect 1392 2775 1396 2779
rect 1460 2775 1464 2779
rect 1504 2775 1508 2779
rect 1564 2775 1568 2779
rect 1608 2775 1612 2779
rect 1676 2775 1680 2779
rect 1712 2775 1716 2779
rect 1764 2775 1768 2779
rect 1932 2775 1936 2779
rect 1976 2775 1980 2779
rect 2020 2775 2024 2779
rect 2064 2775 2068 2779
rect 2108 2775 2112 2779
rect 2152 2775 2156 2779
rect 2196 2775 2200 2779
rect 2240 2775 2244 2779
rect 2284 2775 2288 2779
rect 2328 2775 2332 2779
rect 2372 2775 2376 2779
rect 888 2751 892 2755
rect 1032 2751 1036 2755
rect 1280 2751 1284 2755
rect 1392 2751 1396 2755
rect 1504 2751 1508 2755
rect 1608 2751 1612 2755
rect 2680 2803 2684 2807
rect 2784 2803 2788 2807
rect 2896 2803 2900 2807
rect 3024 2803 3028 2807
rect 2460 2775 2464 2779
rect 2548 2775 2552 2779
rect 2636 2775 2640 2779
rect 2680 2775 2684 2779
rect 2724 2775 2728 2779
rect 2784 2775 2788 2779
rect 2828 2775 2832 2779
rect 2896 2775 2900 2779
rect 2940 2775 2944 2779
rect 3024 2775 3028 2779
rect 3068 2775 3072 2779
rect 3212 2775 3216 2779
rect 3336 2775 3340 2779
rect 3364 2775 3368 2779
rect 3516 2775 3520 2779
rect 2248 2767 2252 2771
rect 2416 2767 2420 2771
rect 1712 2751 1716 2755
rect 2076 2751 2080 2755
rect 2112 2751 2116 2755
rect 2196 2751 2200 2755
rect 2240 2751 2244 2755
rect 2112 2727 2116 2731
rect 2240 2727 2244 2731
rect 2324 2751 2328 2755
rect 2476 2751 2480 2755
rect 2652 2751 2656 2755
rect 2852 2751 2856 2755
rect 2904 2751 2908 2755
rect 3068 2751 3072 2755
rect 3300 2751 3304 2755
rect 2248 2723 2252 2727
rect 3516 2751 3520 2755
rect 3336 2727 3340 2731
rect 2904 2723 2908 2727
rect 3528 2695 3532 2699
rect 2400 2655 2404 2659
rect 204 2643 208 2647
rect 316 2643 320 2647
rect 428 2643 432 2647
rect 540 2643 544 2647
rect 652 2643 656 2647
rect 2624 2655 2628 2659
rect 2728 2655 2732 2659
rect 2840 2655 2844 2659
rect 2952 2655 2956 2659
rect 3064 2655 3068 2659
rect 1980 2627 1984 2631
rect 2092 2627 2096 2631
rect 2204 2627 2208 2631
rect 2324 2627 2328 2631
rect 2400 2627 2404 2631
rect 2444 2627 2448 2631
rect 2556 2627 2560 2631
rect 2624 2627 2628 2631
rect 2668 2627 2672 2631
rect 2728 2627 2732 2631
rect 2772 2627 2776 2631
rect 2840 2627 2844 2631
rect 2884 2627 2888 2631
rect 2952 2627 2956 2631
rect 2996 2627 3000 2631
rect 3064 2627 3068 2631
rect 3108 2627 3112 2631
rect 252 2615 256 2619
rect 336 2615 340 2619
rect 380 2615 384 2619
rect 440 2615 444 2619
rect 524 2615 528 2619
rect 692 2615 696 2619
rect 868 2615 872 2619
rect 1052 2615 1056 2619
rect 1244 2615 1248 2619
rect 1328 2615 1332 2619
rect 1436 2615 1440 2619
rect 1528 2615 1532 2619
rect 1636 2615 1640 2619
rect 336 2591 340 2595
rect 440 2591 444 2595
rect 1328 2591 1332 2595
rect 1924 2611 1928 2615
rect 2000 2611 2004 2615
rect 2100 2611 2104 2615
rect 2184 2611 2188 2615
rect 2292 2611 2296 2615
rect 2492 2611 2496 2615
rect 2584 2611 2588 2615
rect 2692 2611 2696 2615
rect 2900 2611 2904 2615
rect 3108 2611 3112 2615
rect 3152 2611 3156 2615
rect 1528 2591 1532 2595
rect 2000 2587 2004 2591
rect 2184 2587 2188 2591
rect 2584 2587 2588 2591
rect 3152 2583 3156 2587
rect 3272 2611 3276 2615
rect 3324 2611 3328 2615
rect 3516 2611 3520 2615
rect 3528 2555 3532 2559
rect 3272 2531 3276 2535
rect 848 2519 852 2523
rect 1312 2519 1316 2523
rect 2568 2515 2572 2519
rect 308 2491 312 2495
rect 508 2491 512 2495
rect 708 2491 712 2495
rect 840 2491 844 2495
rect 848 2491 852 2495
rect 892 2491 896 2495
rect 1060 2491 1064 2495
rect 1212 2491 1216 2495
rect 1312 2491 1316 2495
rect 1356 2491 1360 2495
rect 1492 2491 1496 2495
rect 1628 2491 1632 2495
rect 1764 2491 1768 2495
rect 2896 2515 2900 2519
rect 3048 2515 3052 2519
rect 212 2475 216 2479
rect 348 2475 352 2479
rect 408 2475 412 2479
rect 492 2475 496 2479
rect 568 2475 572 2479
rect 636 2475 640 2479
rect 696 2475 700 2479
rect 772 2475 776 2479
rect 832 2475 836 2479
rect 408 2451 412 2455
rect 696 2451 700 2455
rect 832 2451 836 2455
rect 1924 2487 1928 2491
rect 2076 2487 2080 2491
rect 2252 2487 2256 2491
rect 2436 2487 2440 2491
rect 2568 2487 2572 2491
rect 2612 2487 2616 2491
rect 2780 2487 2784 2491
rect 2896 2487 2900 2491
rect 2940 2487 2944 2491
rect 3048 2487 3052 2491
rect 3092 2487 3096 2491
rect 3236 2487 3240 2491
rect 3368 2487 3372 2491
rect 3380 2487 3384 2491
rect 3516 2487 3520 2491
rect 908 2475 912 2479
rect 1036 2475 1040 2479
rect 1156 2475 1160 2479
rect 1268 2477 1272 2481
rect 1312 2475 1316 2479
rect 1372 2475 1376 2479
rect 1416 2475 1420 2479
rect 1476 2475 1480 2479
rect 1520 2475 1524 2479
rect 1580 2475 1584 2479
rect 1616 2475 1620 2479
rect 1676 2475 1680 2479
rect 1712 2475 1716 2479
rect 1764 2475 1768 2479
rect 1808 2475 1812 2479
rect 1924 2475 1928 2479
rect 1960 2475 1964 2479
rect 2020 2475 2024 2479
rect 2080 2475 2084 2479
rect 2156 2475 2160 2479
rect 2216 2475 2220 2479
rect 2308 2475 2312 2479
rect 2468 2475 2472 2479
rect 2628 2475 2632 2479
rect 2796 2475 2800 2479
rect 2972 2475 2976 2479
rect 3148 2475 3152 2479
rect 3324 2475 3328 2479
rect 1312 2451 1316 2455
rect 1416 2451 1420 2455
rect 1520 2451 1524 2455
rect 1616 2451 1620 2455
rect 1712 2451 1716 2455
rect 1808 2451 1812 2455
rect 1960 2451 1964 2455
rect 2080 2451 2084 2455
rect 2216 2451 2220 2455
rect 3500 2475 3504 2479
rect 3368 2451 3372 2455
rect 840 2447 844 2451
rect 3512 2419 3516 2423
rect 568 2387 572 2391
rect 1040 2371 1044 2375
rect 1296 2371 1300 2375
rect 1424 2371 1428 2375
rect 2800 2371 2804 2375
rect 2960 2371 2964 2375
rect 3128 2371 3132 2375
rect 188 2343 192 2347
rect 356 2343 360 2347
rect 516 2343 520 2347
rect 676 2343 680 2347
rect 752 2343 756 2347
rect 820 2343 824 2347
rect 956 2343 960 2347
rect 1040 2343 1044 2347
rect 1084 2343 1088 2347
rect 1212 2343 1216 2347
rect 1296 2343 1300 2347
rect 1340 2343 1344 2347
rect 1424 2343 1428 2347
rect 1468 2343 1472 2347
rect 2388 2343 2392 2347
rect 2540 2343 2544 2347
rect 2692 2343 2696 2347
rect 2800 2343 2804 2347
rect 2844 2343 2848 2347
rect 2960 2343 2964 2347
rect 3004 2343 3008 2347
rect 3128 2343 3132 2347
rect 3172 2343 3176 2347
rect 3340 2343 3344 2347
rect 3508 2343 3512 2347
rect 172 2327 176 2331
rect 232 2327 236 2331
rect 292 2327 296 2331
rect 436 2327 440 2331
rect 496 2327 500 2331
rect 572 2327 576 2331
rect 632 2327 636 2331
rect 708 2327 712 2331
rect 232 2303 236 2307
rect 496 2303 500 2307
rect 632 2303 636 2307
rect 752 2303 756 2307
rect 784 2327 788 2331
rect 836 2327 840 2331
rect 888 2327 892 2331
rect 956 2327 960 2331
rect 1000 2327 1004 2331
rect 1068 2327 1072 2331
rect 1188 2327 1192 2331
rect 1308 2327 1312 2331
rect 2380 2327 2384 2331
rect 2476 2327 2480 2331
rect 2588 2327 2592 2331
rect 2732 2329 2736 2333
rect 2840 2327 2844 2331
rect 2908 2327 2912 2331
rect 3108 2327 3112 2331
rect 3316 2327 3320 2331
rect 3516 2327 3520 2331
rect 888 2303 892 2307
rect 1000 2303 1004 2307
rect 2840 2303 2844 2307
rect 2392 2271 2396 2275
rect 3528 2271 3532 2275
rect 784 2247 788 2251
rect 128 2231 132 2235
rect 1048 2231 1052 2235
rect 172 2203 176 2207
rect 268 2203 272 2207
rect 388 2203 392 2207
rect 508 2203 512 2207
rect 628 2203 632 2207
rect 748 2203 752 2207
rect 860 2205 864 2209
rect 2440 2231 2444 2235
rect 972 2203 976 2207
rect 1048 2203 1052 2207
rect 1092 2203 1096 2207
rect 1212 2203 1216 2207
rect 2372 2203 2376 2207
rect 2440 2203 2444 2207
rect 2484 2203 2488 2207
rect 2620 2203 2624 2207
rect 2772 2205 2776 2209
rect 2948 2203 2952 2207
rect 3140 2203 3144 2207
rect 3340 2203 3344 2207
rect 3516 2203 3520 2207
rect 128 2187 132 2191
rect 172 2187 176 2191
rect 208 2187 212 2191
rect 276 2187 280 2191
rect 412 2187 416 2191
rect 472 2187 476 2191
rect 548 2187 552 2191
rect 608 2187 612 2191
rect 684 2187 688 2191
rect 812 2189 816 2193
rect 2284 2191 2288 2195
rect 2372 2191 2376 2195
rect 2468 2191 2472 2195
rect 2580 2191 2584 2195
rect 2724 2191 2728 2195
rect 2900 2191 2904 2195
rect 2944 2191 2948 2195
rect 3100 2191 3104 2195
rect 3200 2191 3204 2195
rect 3316 2191 3320 2195
rect 3516 2191 3520 2195
rect 864 2187 868 2191
rect 940 2187 944 2191
rect 1060 2187 1064 2191
rect 1120 2187 1124 2191
rect 1188 2187 1192 2191
rect 1256 2187 1260 2191
rect 1316 2187 1320 2191
rect 208 2163 212 2167
rect 472 2163 476 2167
rect 608 2163 612 2167
rect 864 2163 868 2167
rect 1120 2159 1124 2163
rect 288 2131 292 2135
rect 2944 2167 2948 2171
rect 3200 2167 3204 2171
rect 3528 2135 3532 2139
rect 1256 2099 1260 2103
rect 3200 2103 3204 2107
rect 2232 2087 2236 2091
rect 824 2083 828 2087
rect 208 2075 212 2079
rect 172 2055 176 2059
rect 936 2083 940 2087
rect 1048 2083 1052 2087
rect 1168 2083 1172 2087
rect 2408 2087 2412 2091
rect 2496 2087 2500 2091
rect 2744 2087 2748 2091
rect 2912 2087 2916 2091
rect 2188 2059 2192 2063
rect 2232 2059 2236 2063
rect 2276 2059 2280 2063
rect 2364 2059 2368 2063
rect 2408 2059 2412 2063
rect 2452 2059 2456 2063
rect 2496 2059 2500 2063
rect 2540 2059 2544 2063
rect 2652 2059 2656 2063
rect 2744 2059 2748 2063
rect 2788 2059 2792 2063
rect 2912 2059 2916 2063
rect 2956 2059 2960 2063
rect 3140 2059 3144 2063
rect 268 2055 272 2059
rect 396 2055 400 2059
rect 516 2055 520 2059
rect 636 2055 640 2059
rect 756 2055 760 2059
rect 824 2055 828 2059
rect 868 2055 872 2059
rect 936 2055 940 2059
rect 980 2055 984 2059
rect 1048 2055 1052 2059
rect 1092 2055 1096 2059
rect 1168 2055 1172 2059
rect 1212 2055 1216 2059
rect 3296 2087 3300 2091
rect 3296 2059 3300 2063
rect 3340 2059 3344 2063
rect 3516 2059 3520 2063
rect 3200 2051 3204 2055
rect 2028 2043 2032 2047
rect 2080 2043 2084 2047
rect 2156 2043 2160 2047
rect 2284 2043 2288 2047
rect 2428 2043 2432 2047
rect 2464 2043 2468 2047
rect 2580 2043 2584 2047
rect 2740 2045 2744 2049
rect 2908 2043 2912 2047
rect 3092 2043 3096 2047
rect 3276 2043 3280 2047
rect 3468 2043 3472 2047
rect 196 2031 200 2035
rect 208 2031 212 2035
rect 340 2031 344 2035
rect 476 2031 480 2035
rect 528 2031 532 2035
rect 604 2031 608 2035
rect 724 2031 728 2035
rect 836 2031 840 2035
rect 940 2031 944 2035
rect 1044 2031 1048 2035
rect 1148 2031 1152 2035
rect 1252 2031 1256 2035
rect 1296 2031 1300 2035
rect 1356 2031 1360 2035
rect 528 2007 532 2011
rect 2080 2019 2084 2023
rect 2464 2019 2468 2023
rect 1296 2003 1300 2007
rect 208 1975 212 1979
rect 2392 1939 2396 1943
rect 288 1935 292 1939
rect 432 1935 436 1939
rect 196 1907 200 1911
rect 288 1907 292 1911
rect 332 1907 336 1911
rect 1232 1935 1236 1939
rect 476 1907 480 1911
rect 620 1909 624 1913
rect 2608 1939 2612 1943
rect 1940 1911 1944 1915
rect 2196 1911 2200 1915
rect 2392 1911 2396 1915
rect 2436 1911 2440 1915
rect 756 1907 760 1911
rect 892 1907 896 1911
rect 1028 1907 1032 1911
rect 1156 1907 1160 1911
rect 1232 1907 1236 1911
rect 1276 1907 1280 1911
rect 1396 1907 1400 1911
rect 1516 1907 1520 1911
rect 1636 1907 1640 1911
rect 2056 1907 2060 1911
rect 1924 1901 1928 1905
rect 2012 1899 2016 1903
rect 2048 1899 2052 1903
rect 252 1887 256 1891
rect 320 1887 324 1891
rect 432 1887 436 1891
rect 508 1887 512 1891
rect 748 1887 752 1891
rect 964 1887 968 1891
rect 1040 1887 1044 1891
rect 1156 1887 1160 1891
rect 1232 1887 1236 1891
rect 1324 1887 1328 1891
rect 1392 1887 1396 1891
rect 1484 1887 1488 1891
rect 1552 1887 1556 1891
rect 1636 1887 1640 1891
rect 1764 1887 1768 1891
rect 1040 1863 1044 1867
rect 1232 1863 1236 1867
rect 1392 1863 1396 1867
rect 2048 1875 2052 1879
rect 2808 1939 2812 1943
rect 2992 1939 2996 1943
rect 3160 1939 3164 1943
rect 3328 1939 3332 1943
rect 2652 1911 2656 1915
rect 2808 1911 2812 1915
rect 2852 1911 2856 1915
rect 2992 1911 2996 1915
rect 3036 1911 3040 1915
rect 3160 1911 3164 1915
rect 3204 1911 3208 1915
rect 3328 1911 3332 1915
rect 3372 1911 3376 1915
rect 3516 1911 3520 1915
rect 2100 1899 2104 1903
rect 2196 1899 2200 1903
rect 2248 1899 2252 1903
rect 2324 1899 2328 1903
rect 2392 1899 2396 1903
rect 2476 1899 2480 1903
rect 2608 1899 2612 1903
rect 2636 1899 2640 1903
rect 2696 1899 2700 1903
rect 2796 1899 2800 1903
rect 2948 1899 2952 1903
rect 3016 1899 3020 1903
rect 3100 1899 3104 1903
rect 3160 1899 3164 1903
rect 3244 1899 3248 1903
rect 3388 1899 3392 1903
rect 3516 1899 3520 1903
rect 2248 1875 2252 1879
rect 2392 1875 2396 1879
rect 2696 1875 2700 1879
rect 3016 1875 3020 1879
rect 3160 1875 3164 1879
rect 2056 1871 2060 1875
rect 1552 1863 1556 1867
rect 320 1859 324 1863
rect 3336 1859 3340 1863
rect 264 1831 268 1835
rect 1776 1831 1780 1835
rect 2432 1799 2436 1803
rect 408 1791 412 1795
rect 2008 1771 2012 1775
rect 2036 1771 2040 1775
rect 2260 1771 2264 1775
rect 284 1763 288 1767
rect 408 1763 412 1767
rect 452 1763 456 1767
rect 628 1763 632 1767
rect 796 1763 800 1767
rect 964 1763 968 1767
rect 1116 1763 1120 1767
rect 1260 1763 1264 1767
rect 1396 1763 1400 1767
rect 1524 1763 1528 1767
rect 1652 1763 1656 1767
rect 1764 1763 1768 1767
rect 1972 1755 1976 1759
rect 356 1749 360 1753
rect 416 1747 420 1751
rect 500 1747 504 1751
rect 644 1747 648 1751
rect 796 1747 800 1751
rect 864 1747 868 1751
rect 948 1747 952 1751
rect 1100 1747 1104 1751
rect 1208 1747 1212 1751
rect 1252 1747 1256 1751
rect 1320 1747 1324 1751
rect 1404 1747 1408 1751
rect 1556 1749 1560 1753
rect 1624 1747 1628 1751
rect 1716 1747 1720 1751
rect 416 1723 420 1727
rect 864 1723 868 1727
rect 1208 1723 1212 1727
rect 1320 1723 1324 1727
rect 2632 1799 2636 1803
rect 2476 1771 2480 1775
rect 2632 1771 2636 1775
rect 2676 1771 2680 1775
rect 2868 1771 2872 1775
rect 3052 1771 3056 1775
rect 3236 1771 3240 1775
rect 3336 1771 3340 1775
rect 3428 1771 3432 1775
rect 2116 1755 2120 1759
rect 2224 1755 2228 1759
rect 2276 1755 2280 1759
rect 2432 1755 2436 1759
rect 2444 1755 2448 1759
rect 2528 1755 2532 1759
rect 2628 1755 2632 1759
rect 2820 1755 2824 1759
rect 2912 1755 2916 1759
rect 3020 1755 3024 1759
rect 3228 1755 3232 1759
rect 3444 1755 3448 1759
rect 2008 1731 2012 1735
rect 1624 1723 1628 1727
rect 2528 1731 2532 1735
rect 2912 1731 2916 1735
rect 3456 1699 3460 1703
rect 2224 1671 2228 1675
rect 2024 1655 2028 1659
rect 880 1647 884 1651
rect 1416 1639 1420 1643
rect 348 1619 352 1623
rect 484 1619 488 1623
rect 628 1619 632 1623
rect 772 1619 776 1623
rect 880 1619 884 1623
rect 924 1619 928 1623
rect 1076 1619 1080 1623
rect 1228 1619 1232 1623
rect 1380 1619 1384 1623
rect 2144 1655 2148 1659
rect 2392 1655 2396 1659
rect 1948 1627 1952 1631
rect 2024 1627 2028 1631
rect 2068 1627 2072 1631
rect 2144 1627 2148 1631
rect 2188 1627 2192 1631
rect 2308 1627 2312 1631
rect 2392 1627 2396 1631
rect 2436 1627 2440 1631
rect 2580 1627 2584 1631
rect 2732 1627 2736 1631
rect 2900 1627 2904 1631
rect 3084 1627 3088 1631
rect 3276 1627 3280 1631
rect 3468 1627 3472 1631
rect 1532 1619 1536 1623
rect 1684 1619 1688 1623
rect 1924 1607 1928 1611
rect 2044 1607 2048 1611
rect 2112 1607 2116 1611
rect 2180 1607 2184 1611
rect 2316 1607 2320 1611
rect 2360 1607 2364 1611
rect 2460 1607 2464 1611
rect 2612 1609 2616 1613
rect 2680 1607 2684 1611
rect 2772 1607 2776 1611
rect 2864 1607 2868 1611
rect 2940 1607 2944 1611
rect 3024 1607 3028 1611
rect 3124 1607 3128 1611
rect 3308 1607 3312 1611
rect 3500 1607 3504 1611
rect 252 1599 256 1603
rect 328 1599 332 1603
rect 380 1599 384 1603
rect 440 1599 444 1603
rect 516 1599 520 1603
rect 652 1599 656 1603
rect 712 1599 716 1603
rect 788 1599 792 1603
rect 932 1599 936 1603
rect 1000 1599 1004 1603
rect 1084 1599 1088 1603
rect 1244 1599 1248 1603
rect 1404 1599 1408 1603
rect 1416 1599 1420 1603
rect 1480 1599 1484 1603
rect 1572 1599 1576 1603
rect 328 1575 332 1579
rect 440 1575 444 1579
rect 712 1575 716 1579
rect 1000 1575 1004 1579
rect 1480 1575 1484 1579
rect 2680 1583 2684 1587
rect 2864 1583 2868 1587
rect 3024 1583 3028 1587
rect 2360 1579 2364 1583
rect 3512 1551 3516 1555
rect 2112 1519 2116 1523
rect 2016 1503 2020 1507
rect 208 1499 212 1503
rect 1336 1499 1340 1503
rect 2336 1503 2340 1507
rect 2496 1503 2500 1507
rect 2976 1503 2980 1507
rect 3144 1503 3148 1507
rect 1808 1475 1812 1479
rect 1924 1475 1928 1479
rect 2016 1475 2020 1479
rect 2060 1475 2064 1479
rect 2220 1475 2224 1479
rect 2336 1475 2340 1479
rect 2380 1475 2384 1479
rect 2496 1475 2500 1479
rect 2540 1475 2544 1479
rect 2700 1475 2704 1479
rect 2860 1475 2864 1479
rect 2976 1475 2980 1479
rect 3020 1475 3024 1479
rect 3144 1475 3148 1479
rect 3188 1475 3192 1479
rect 3356 1475 3360 1479
rect 3516 1475 3520 1479
rect 172 1471 176 1475
rect 208 1471 212 1475
rect 308 1471 312 1475
rect 460 1471 464 1475
rect 620 1471 624 1475
rect 728 1471 732 1475
rect 772 1471 776 1475
rect 924 1471 928 1475
rect 1076 1471 1080 1475
rect 1228 1471 1232 1475
rect 1336 1471 1340 1475
rect 1380 1471 1384 1475
rect 1532 1471 1536 1475
rect 172 1451 176 1455
rect 208 1451 212 1455
rect 292 1451 296 1455
rect 352 1451 356 1455
rect 428 1451 432 1455
rect 564 1451 568 1455
rect 616 1451 620 1455
rect 692 1451 696 1455
rect 208 1427 212 1431
rect 352 1427 356 1431
rect 616 1427 620 1431
rect 820 1453 824 1457
rect 728 1427 732 1431
rect 872 1451 876 1455
rect 940 1451 944 1455
rect 984 1451 988 1455
rect 1052 1451 1056 1455
rect 1172 1451 1176 1455
rect 1292 1451 1296 1455
rect 1412 1451 1416 1455
rect 1464 1451 1468 1455
rect 1532 1451 1536 1455
rect 1592 1451 1596 1455
rect 1660 1451 1664 1455
rect 1704 1451 1708 1455
rect 1764 1451 1768 1455
rect 872 1427 876 1431
rect 984 1427 988 1431
rect 1464 1427 1468 1431
rect 1704 1427 1708 1431
rect 2212 1455 2216 1459
rect 2288 1455 2292 1459
rect 2388 1455 2392 1459
rect 2556 1455 2560 1459
rect 2716 1455 2720 1459
rect 2824 1455 2828 1459
rect 2876 1455 2880 1459
rect 2944 1455 2948 1459
rect 3036 1455 3040 1459
rect 3112 1455 3116 1459
rect 3204 1455 3208 1459
rect 3280 1455 3284 1459
rect 3372 1455 3376 1459
rect 3516 1455 3520 1459
rect 2288 1431 2292 1435
rect 2824 1431 2828 1435
rect 2944 1431 2948 1435
rect 3112 1431 3116 1435
rect 3280 1431 3284 1435
rect 1808 1427 1812 1431
rect 3528 1399 3532 1403
rect 1592 1371 1596 1375
rect 208 1355 212 1359
rect 1496 1355 1500 1359
rect 2256 1351 2260 1355
rect 172 1327 176 1331
rect 208 1327 212 1331
rect 364 1327 368 1331
rect 588 1327 592 1331
rect 820 1327 824 1331
rect 984 1327 988 1331
rect 1060 1327 1064 1331
rect 1300 1327 1304 1331
rect 1496 1327 1500 1331
rect 1540 1327 1544 1331
rect 1752 1327 1756 1331
rect 1764 1327 1768 1331
rect 2608 1351 2612 1355
rect 2928 1351 2932 1355
rect 3072 1351 3076 1355
rect 3216 1351 3220 1355
rect 3352 1351 3356 1355
rect 172 1307 176 1311
rect 208 1307 212 1311
rect 356 1307 360 1311
rect 556 1307 560 1311
rect 640 1307 644 1311
rect 748 1307 752 1311
rect 832 1307 836 1311
rect 932 1307 936 1311
rect 208 1283 212 1287
rect 640 1283 644 1287
rect 832 1283 836 1287
rect 1100 1309 1104 1313
rect 1260 1307 1264 1311
rect 1328 1307 1332 1311
rect 1412 1307 1416 1311
rect 1480 1307 1484 1311
rect 1564 1307 1568 1311
rect 1632 1307 1636 1311
rect 1716 1307 1720 1311
rect 984 1283 988 1287
rect 1328 1283 1332 1287
rect 1480 1283 1484 1287
rect 1632 1283 1636 1287
rect 2116 1323 2120 1327
rect 2256 1323 2260 1327
rect 2300 1323 2304 1327
rect 2476 1323 2480 1327
rect 2608 1323 2612 1327
rect 2652 1323 2656 1327
rect 2820 1323 2824 1327
rect 2928 1323 2932 1327
rect 2972 1323 2976 1327
rect 3072 1323 3076 1327
rect 3116 1323 3120 1327
rect 3216 1323 3220 1327
rect 3260 1323 3264 1327
rect 3396 1323 3400 1327
rect 3516 1323 3520 1327
rect 2116 1311 2120 1315
rect 2340 1311 2344 1315
rect 2432 1311 2436 1315
rect 2548 1311 2552 1315
rect 2740 1311 2744 1315
rect 2816 1311 2820 1315
rect 2916 1311 2920 1315
rect 3076 1311 3080 1315
rect 3228 1311 3232 1315
rect 3288 1311 3292 1315
rect 3352 1311 3356 1315
rect 3380 1311 3384 1315
rect 3516 1311 3520 1315
rect 2432 1287 2436 1291
rect 2816 1287 2820 1291
rect 1752 1283 1756 1287
rect 3288 1283 3292 1287
rect 2128 1255 2132 1259
rect 2928 1255 2932 1259
rect 3528 1255 3532 1259
rect 2624 1211 2628 1215
rect 288 1207 292 1211
rect 472 1207 476 1211
rect 1104 1207 1108 1211
rect 1240 1207 1244 1211
rect 1376 1207 1380 1211
rect 1520 1207 1524 1211
rect 1940 1183 1944 1187
rect 2028 1185 2032 1189
rect 2132 1183 2136 1187
rect 2252 1183 2256 1187
rect 2388 1185 2392 1189
rect 3056 1211 3060 1215
rect 3200 1211 3204 1215
rect 2512 1183 2516 1187
rect 2524 1183 2528 1187
rect 2624 1183 2628 1187
rect 2668 1183 2672 1187
rect 2812 1183 2816 1187
rect 2956 1183 2960 1187
rect 3056 1183 3060 1187
rect 3100 1183 3104 1187
rect 3200 1183 3204 1187
rect 3244 1183 3248 1187
rect 3388 1183 3392 1187
rect 3516 1183 3520 1187
rect 172 1179 176 1183
rect 288 1179 292 1183
rect 332 1179 336 1183
rect 472 1179 476 1183
rect 516 1179 520 1183
rect 692 1179 696 1183
rect 824 1179 828 1183
rect 852 1179 856 1183
rect 1004 1179 1008 1183
rect 1104 1179 1108 1183
rect 1148 1179 1152 1183
rect 1240 1179 1244 1183
rect 1284 1179 1288 1183
rect 1376 1179 1380 1183
rect 1420 1179 1424 1183
rect 1520 1179 1524 1183
rect 1564 1179 1568 1183
rect 196 1163 200 1167
rect 348 1163 352 1167
rect 500 1163 504 1167
rect 644 1163 648 1167
rect 704 1163 708 1167
rect 788 1163 792 1167
rect 704 1139 708 1143
rect 1924 1167 1928 1171
rect 2092 1167 2096 1171
rect 2176 1167 2180 1171
rect 2284 1167 2288 1171
rect 2468 1167 2472 1171
rect 940 1163 944 1167
rect 1008 1163 1012 1167
rect 1092 1163 1096 1167
rect 1168 1163 1172 1167
rect 1260 1163 1264 1167
rect 1336 1163 1340 1167
rect 1428 1163 1432 1167
rect 1528 1163 1532 1167
rect 1604 1163 1608 1167
rect 1764 1163 1768 1167
rect 824 1139 828 1143
rect 1008 1139 1012 1143
rect 1168 1139 1172 1143
rect 1336 1139 1340 1143
rect 2176 1143 2180 1147
rect 2644 1167 2648 1171
rect 2720 1167 2724 1171
rect 2820 1167 2824 1171
rect 2896 1167 2900 1171
rect 2996 1167 3000 1171
rect 3056 1167 3060 1171
rect 3172 1167 3176 1171
rect 3356 1167 3360 1171
rect 3516 1167 3520 1171
rect 2512 1143 2516 1147
rect 2720 1143 2724 1147
rect 2896 1143 2900 1147
rect 3056 1143 3060 1147
rect 1528 1139 1532 1143
rect 3528 1111 3532 1115
rect 1776 1107 1780 1111
rect 320 1063 324 1067
rect 432 1063 436 1067
rect 544 1063 548 1067
rect 252 1035 256 1039
rect 320 1035 324 1039
rect 364 1035 368 1039
rect 432 1035 436 1039
rect 476 1035 480 1039
rect 544 1035 548 1039
rect 552 1063 556 1067
rect 936 1063 940 1067
rect 1032 1063 1036 1067
rect 1240 1063 1244 1067
rect 1400 1063 1404 1067
rect 2400 1059 2404 1063
rect 596 1035 600 1039
rect 716 1035 720 1039
rect 844 1035 848 1039
rect 936 1035 940 1039
rect 980 1035 984 1039
rect 1032 1035 1036 1039
rect 1124 1035 1128 1039
rect 1240 1035 1244 1039
rect 1284 1035 1288 1039
rect 1400 1035 1404 1039
rect 1444 1035 1448 1039
rect 1612 1035 1616 1039
rect 1764 1035 1768 1039
rect 2856 1059 2860 1063
rect 1972 1031 1976 1035
rect 2132 1031 2136 1035
rect 2284 1031 2288 1035
rect 2400 1031 2404 1035
rect 2444 1031 2448 1035
rect 2604 1031 2608 1035
rect 2772 1031 2776 1035
rect 2856 1031 2860 1035
rect 2948 1031 2952 1035
rect 3132 1031 3136 1035
rect 3264 1031 3268 1035
rect 3324 1031 3328 1035
rect 3516 1031 3520 1035
rect 372 1015 376 1019
rect 460 1015 464 1019
rect 552 1015 556 1019
rect 564 1015 568 1019
rect 684 1015 688 1019
rect 820 1015 824 1019
rect 980 1015 984 1019
rect 1164 1015 1168 1019
rect 1356 1015 1360 1019
rect 1564 1015 1568 1019
rect 1624 1015 1628 1019
rect 1764 1015 1768 1019
rect 1972 1015 1976 1019
rect 2100 1015 2104 1019
rect 2152 1015 2156 1019
rect 2220 1015 2224 1019
rect 2272 1015 2276 1019
rect 2340 1015 2344 1019
rect 2392 1015 2396 1019
rect 2468 1015 2472 1019
rect 2604 1015 2608 1019
rect 2664 1015 2668 1019
rect 2748 1015 2752 1019
rect 2824 1015 2828 1019
rect 2900 1015 2904 1019
rect 2968 1015 2972 1019
rect 3060 1015 3064 1019
rect 3220 1015 3224 1019
rect 1624 991 1628 995
rect 2152 991 2156 995
rect 2272 991 2276 995
rect 2392 991 2396 995
rect 2664 991 2668 995
rect 2824 991 2828 995
rect 2968 991 2972 995
rect 3264 991 3268 995
rect 3288 1015 3292 1019
rect 3380 1015 3384 1019
rect 3516 1015 3520 1019
rect 3288 987 3292 991
rect 384 959 388 963
rect 456 915 460 919
rect 696 915 700 919
rect 840 915 844 919
rect 1520 915 1524 919
rect 2016 915 2020 919
rect 2624 915 2628 919
rect 3016 915 3020 919
rect 404 887 408 891
rect 456 887 460 891
rect 500 887 504 891
rect 612 887 616 891
rect 696 887 700 891
rect 740 887 744 891
rect 840 887 844 891
rect 884 887 888 891
rect 992 887 996 891
rect 1044 887 1048 891
rect 1212 887 1216 891
rect 1388 887 1392 891
rect 1520 887 1524 891
rect 1564 887 1568 891
rect 1748 887 1752 891
rect 1924 887 1928 891
rect 2016 887 2020 891
rect 2084 887 2088 891
rect 2236 887 2240 891
rect 2388 887 2392 891
rect 2532 887 2536 891
rect 2624 887 2628 891
rect 2668 887 2672 891
rect 2796 887 2800 891
rect 2924 887 2928 891
rect 3016 887 3020 891
rect 3060 887 3064 891
rect 372 871 376 875
rect 460 871 464 875
rect 564 871 568 875
rect 676 871 680 875
rect 812 871 816 875
rect 956 871 960 875
rect 1924 875 1928 879
rect 2044 875 2048 879
rect 2196 875 2200 879
rect 2264 875 2268 879
rect 2348 875 2352 879
rect 2516 875 2520 879
rect 2692 875 2696 879
rect 2760 875 2764 879
rect 2876 875 2880 879
rect 3068 875 3072 879
rect 3160 875 3164 879
rect 3268 875 3272 879
rect 3468 875 3472 879
rect 1116 871 1120 875
rect 1292 871 1296 875
rect 1476 871 1480 875
rect 1660 871 1664 875
rect 2264 851 2268 855
rect 3160 851 3164 855
rect 992 847 996 851
rect 2760 847 2764 851
rect 1936 819 1940 823
rect 1488 815 1492 819
rect 2128 779 2132 783
rect 528 775 532 779
rect 324 749 328 753
rect 816 775 820 779
rect 1120 775 1124 779
rect 1432 775 1436 779
rect 444 747 448 751
rect 528 747 532 751
rect 572 747 576 751
rect 716 747 720 751
rect 816 747 820 751
rect 860 747 864 751
rect 1000 747 1004 751
rect 1012 747 1016 751
rect 1120 747 1124 751
rect 1164 747 1168 751
rect 1316 747 1320 751
rect 244 731 248 735
rect 388 731 392 735
rect 448 731 452 735
rect 532 731 536 735
rect 676 731 680 735
rect 820 731 824 735
rect 964 733 968 737
rect 448 707 452 711
rect 1592 775 1596 779
rect 2792 779 2796 783
rect 3312 779 3316 783
rect 2960 771 2964 775
rect 1924 751 1928 755
rect 2028 751 2032 755
rect 2128 751 2132 755
rect 2172 751 2176 755
rect 2324 751 2328 755
rect 2492 751 2496 755
rect 2660 751 2664 755
rect 2792 751 2796 755
rect 2836 751 2840 755
rect 2960 751 2964 755
rect 3004 751 3008 755
rect 3180 751 3184 755
rect 3312 751 3316 755
rect 3356 751 3360 755
rect 3516 751 3520 755
rect 1476 747 1480 751
rect 1592 747 1596 751
rect 1636 747 1640 751
rect 1924 735 1928 739
rect 2092 735 2096 739
rect 2176 735 2180 739
rect 2284 735 2288 739
rect 2368 735 2372 739
rect 2476 735 2480 739
rect 2668 735 2672 739
rect 2852 735 2856 739
rect 3028 735 3032 739
rect 3104 735 3108 739
rect 3196 735 3200 739
rect 3364 735 3368 739
rect 3516 735 3520 739
rect 1116 731 1120 735
rect 1232 731 1236 735
rect 1276 731 1280 735
rect 1432 731 1436 735
rect 1444 731 1448 735
rect 1520 731 1524 735
rect 1612 731 1616 735
rect 1764 731 1768 735
rect 1000 707 1004 711
rect 1232 707 1236 711
rect 2176 711 2180 715
rect 2368 711 2372 715
rect 3104 711 3108 715
rect 1520 707 1524 711
rect 3528 679 3532 683
rect 1776 675 1780 679
rect 768 635 772 639
rect 200 627 204 631
rect 172 607 176 611
rect 1024 635 1028 639
rect 1336 635 1340 639
rect 332 607 336 611
rect 500 607 504 611
rect 660 607 664 611
rect 768 607 772 611
rect 812 607 816 611
rect 964 607 968 611
rect 1000 607 1004 611
rect 1024 607 1028 611
rect 1108 607 1112 611
rect 1244 609 1248 613
rect 1336 607 1340 611
rect 1380 607 1384 611
rect 1516 607 1520 611
rect 1652 607 1656 611
rect 1764 607 1768 611
rect 2252 607 2256 611
rect 2396 607 2400 611
rect 2536 607 2540 611
rect 2548 607 2552 611
rect 2708 607 2712 611
rect 2868 607 2872 611
rect 3028 607 3032 611
rect 3196 607 3200 611
rect 3364 607 3368 611
rect 3516 607 3520 611
rect 172 591 176 595
rect 200 591 204 595
rect 208 591 212 595
rect 332 591 336 595
rect 416 591 420 595
rect 516 591 520 595
rect 700 591 704 595
rect 876 591 880 595
rect 208 567 212 571
rect 416 567 420 571
rect 1052 591 1056 595
rect 1228 591 1232 595
rect 1404 591 1408 595
rect 1588 591 1592 595
rect 1664 591 1668 595
rect 1764 591 1768 595
rect 2228 591 2232 595
rect 2264 591 2268 595
rect 2316 591 2320 595
rect 2352 591 2356 595
rect 2404 591 2408 595
rect 2440 591 2444 595
rect 2492 591 2496 595
rect 1664 567 1668 571
rect 2264 567 2268 571
rect 2352 567 2356 571
rect 2440 567 2444 571
rect 2596 593 2600 597
rect 2536 567 2540 571
rect 2640 591 2644 595
rect 2708 591 2712 595
rect 2844 591 2848 595
rect 3004 591 3008 595
rect 3172 591 3176 595
rect 3256 591 3260 595
rect 3356 591 3360 595
rect 3516 591 3520 595
rect 2640 567 2644 571
rect 3256 567 3260 571
rect 1000 563 1004 567
rect 528 535 532 539
rect 1240 535 1244 539
rect 3528 535 3532 539
rect 1344 491 1348 495
rect 200 483 204 487
rect 172 463 176 467
rect 3088 491 3092 495
rect 3344 491 3348 495
rect 340 463 344 467
rect 532 463 536 467
rect 716 463 720 467
rect 900 463 904 467
rect 1068 463 1072 467
rect 1228 463 1232 467
rect 1344 463 1348 467
rect 1388 463 1392 467
rect 1540 463 1544 467
rect 1700 463 1704 467
rect 2340 463 2344 467
rect 2436 463 2440 467
rect 2540 463 2544 467
rect 2644 463 2648 467
rect 2756 463 2760 467
rect 2876 463 2880 467
rect 3004 463 3008 467
rect 3088 463 3092 467
rect 3132 463 3136 467
rect 3260 463 3264 467
rect 3344 463 3348 467
rect 3388 463 3392 467
rect 3516 463 3520 467
rect 2268 451 2272 455
rect 2304 451 2308 455
rect 2356 451 2360 455
rect 2400 451 2404 455
rect 2460 451 2464 455
rect 2512 451 2516 455
rect 2588 451 2592 455
rect 2632 451 2636 455
rect 2724 451 2728 455
rect 2876 451 2880 455
rect 2944 451 2948 455
rect 3028 451 3032 455
rect 3188 451 3192 455
rect 3356 451 3360 455
rect 3408 451 3412 455
rect 3516 451 3520 455
rect 172 447 176 451
rect 200 447 204 451
rect 208 447 212 451
rect 332 447 336 451
rect 376 447 380 451
rect 524 447 528 451
rect 664 447 668 451
rect 716 447 720 451
rect 760 447 764 451
rect 908 447 912 451
rect 1084 447 1088 451
rect 1252 447 1256 451
rect 1420 447 1424 451
rect 1588 447 1592 451
rect 1664 447 1668 451
rect 1756 447 1760 451
rect 208 423 212 427
rect 376 423 380 427
rect 760 423 764 427
rect 2304 427 2308 431
rect 2400 427 2404 431
rect 2512 427 2516 431
rect 2632 427 2636 431
rect 2944 427 2948 431
rect 1664 423 1668 427
rect 1768 391 1772 395
rect 3528 395 3532 399
rect 3408 371 3412 375
rect 664 367 668 371
rect 2280 355 2284 359
rect 208 351 212 355
rect 1576 351 1580 355
rect 172 323 176 327
rect 208 323 212 327
rect 300 323 304 327
rect 460 323 464 327
rect 628 323 632 327
rect 804 323 808 327
rect 972 323 976 327
rect 1140 323 1144 327
rect 1300 323 1304 327
rect 1460 325 1464 329
rect 2392 355 2396 359
rect 2520 355 2524 359
rect 2744 355 2748 359
rect 3288 355 3292 359
rect 3456 355 3460 359
rect 2160 327 2164 331
rect 2220 327 2224 331
rect 2280 327 2284 331
rect 2324 327 2328 331
rect 2392 327 2396 331
rect 2436 327 2440 331
rect 2520 327 2524 331
rect 2564 327 2568 331
rect 2708 327 2712 331
rect 2744 327 2748 331
rect 2852 327 2856 331
rect 3004 327 3008 331
rect 3164 327 3168 331
rect 3288 327 3292 331
rect 3332 327 3336 331
rect 3456 327 3460 331
rect 3500 327 3504 331
rect 1576 323 1580 327
rect 1620 323 1624 327
rect 1764 323 1768 327
rect 244 311 248 315
rect 304 311 308 315
rect 380 311 384 315
rect 524 311 528 315
rect 568 311 572 315
rect 668 311 672 315
rect 736 311 740 315
rect 820 311 824 315
rect 964 311 968 315
rect 1024 311 1028 315
rect 1108 311 1112 315
rect 1252 311 1256 315
rect 1312 311 1316 315
rect 1388 311 1392 315
rect 1424 311 1428 315
rect 1516 311 1520 315
rect 1652 311 1656 315
rect 1696 311 1700 315
rect 1764 311 1768 315
rect 304 287 308 291
rect 560 287 564 291
rect 736 287 740 291
rect 1312 287 1316 291
rect 1424 287 1428 291
rect 1696 287 1700 291
rect 1808 307 1812 311
rect 1924 307 1928 311
rect 2116 307 2120 311
rect 1808 287 1812 291
rect 2332 307 2336 311
rect 2540 307 2544 311
rect 2632 307 2636 311
rect 2740 307 2744 311
rect 2932 307 2936 311
rect 3124 307 3128 311
rect 3216 307 3220 311
rect 3324 307 3328 311
rect 3516 307 3520 311
rect 2160 287 2164 291
rect 1024 283 1028 287
rect 2632 283 2636 287
rect 3216 279 3220 283
rect 392 255 396 259
rect 1936 251 1940 255
rect 3528 251 3532 255
rect 1992 211 1996 215
rect 480 207 484 211
rect 268 181 272 185
rect 1024 207 1028 211
rect 1288 207 1292 211
rect 2136 211 2140 215
rect 2688 203 2692 207
rect 1924 183 1928 187
rect 1992 183 1996 187
rect 2036 183 2040 187
rect 2136 183 2140 187
rect 2180 183 2184 187
rect 2332 183 2336 187
rect 2492 183 2496 187
rect 2652 183 2656 187
rect 396 179 400 183
rect 480 179 484 183
rect 524 179 528 183
rect 660 179 664 183
rect 796 179 800 183
rect 932 179 936 183
rect 1024 179 1028 183
rect 1068 179 1072 183
rect 1196 179 1200 183
rect 1288 179 1292 183
rect 1332 179 1336 183
rect 1468 179 1472 183
rect 1480 151 1484 155
rect 204 143 208 147
rect 240 143 244 147
rect 292 143 296 147
rect 328 143 332 147
rect 380 143 384 147
rect 416 143 420 147
rect 468 143 472 147
rect 504 143 508 147
rect 556 143 560 147
rect 592 143 596 147
rect 644 143 648 147
rect 680 143 684 147
rect 732 143 736 147
rect 768 143 772 147
rect 820 143 824 147
rect 908 143 912 147
rect 996 143 1000 147
rect 1040 143 1044 147
rect 1084 143 1088 147
rect 1172 143 1176 147
rect 1260 145 1264 149
rect 1348 143 1352 147
rect 1384 143 1388 147
rect 1436 143 1440 147
rect 1472 143 1476 147
rect 240 119 244 123
rect 328 119 332 123
rect 416 119 420 123
rect 504 119 508 123
rect 592 119 596 123
rect 680 119 684 123
rect 768 119 772 123
rect 1384 119 1388 123
rect 1472 119 1476 123
rect 1532 143 1536 147
rect 1924 145 1928 149
rect 2820 183 2824 187
rect 2988 183 2992 187
rect 3164 183 3168 187
rect 3348 183 3352 187
rect 3516 183 3520 187
rect 1968 143 1972 147
rect 2012 143 2016 147
rect 2048 143 2052 147
rect 2100 143 2104 147
rect 2136 143 2140 147
rect 2188 143 2192 147
rect 2224 143 2228 147
rect 2276 143 2280 147
rect 2312 143 2316 147
rect 2364 143 2368 147
rect 2408 143 2412 147
rect 2468 143 2472 147
rect 2572 143 2576 147
rect 2676 143 2680 147
rect 2688 143 2692 147
rect 2712 143 2716 147
rect 2772 143 2776 147
rect 2824 143 2828 147
rect 2868 143 2872 147
rect 2904 143 2908 147
rect 2964 143 2968 147
rect 3000 143 3004 147
rect 3060 143 3064 147
rect 3096 143 3100 147
rect 3156 143 3160 147
rect 3192 143 3196 147
rect 3252 143 3256 147
rect 3288 143 3292 147
rect 3340 143 3344 147
rect 3428 143 3432 147
rect 3516 143 3520 147
rect 1968 119 1972 123
rect 2048 119 2052 123
rect 2136 119 2140 123
rect 2224 119 2228 123
rect 2312 119 2316 123
rect 2408 119 2412 123
rect 2712 119 2716 123
rect 2824 119 2828 123
rect 2904 119 2908 123
rect 3000 119 3004 123
rect 3096 119 3100 123
rect 3192 119 3196 123
rect 3288 119 3292 123
rect 1040 115 1044 119
rect 1480 115 1484 119
<< m2 >>
rect 267 3643 273 3644
rect 267 3639 268 3643
rect 272 3642 273 3643
rect 306 3643 312 3644
rect 306 3642 307 3643
rect 272 3640 307 3642
rect 272 3639 273 3640
rect 267 3638 273 3639
rect 306 3639 307 3640
rect 311 3639 312 3643
rect 306 3638 312 3639
rect 355 3643 361 3644
rect 355 3639 356 3643
rect 360 3642 361 3643
rect 394 3643 400 3644
rect 394 3642 395 3643
rect 360 3640 395 3642
rect 360 3639 361 3640
rect 355 3638 361 3639
rect 394 3639 395 3640
rect 399 3639 400 3643
rect 394 3638 400 3639
rect 443 3643 449 3644
rect 443 3639 444 3643
rect 448 3642 449 3643
rect 482 3643 488 3644
rect 482 3642 483 3643
rect 448 3640 483 3642
rect 448 3639 449 3640
rect 443 3638 449 3639
rect 482 3639 483 3640
rect 487 3639 488 3643
rect 482 3638 488 3639
rect 531 3643 537 3644
rect 531 3639 532 3643
rect 536 3642 537 3643
rect 570 3643 576 3644
rect 570 3642 571 3643
rect 536 3640 571 3642
rect 536 3639 537 3640
rect 531 3638 537 3639
rect 570 3639 571 3640
rect 575 3639 576 3643
rect 570 3638 576 3639
rect 619 3643 625 3644
rect 619 3639 620 3643
rect 624 3642 625 3643
rect 658 3643 664 3644
rect 658 3642 659 3643
rect 624 3640 659 3642
rect 624 3639 625 3640
rect 619 3638 625 3639
rect 658 3639 659 3640
rect 663 3639 664 3643
rect 658 3638 664 3639
rect 238 3633 244 3634
rect 238 3629 239 3633
rect 243 3629 244 3633
rect 238 3628 244 3629
rect 326 3633 332 3634
rect 326 3629 327 3633
rect 331 3629 332 3633
rect 326 3628 332 3629
rect 414 3633 420 3634
rect 414 3629 415 3633
rect 419 3629 420 3633
rect 414 3628 420 3629
rect 502 3633 508 3634
rect 502 3629 503 3633
rect 507 3629 508 3633
rect 502 3628 508 3629
rect 590 3633 596 3634
rect 590 3629 591 3633
rect 595 3629 596 3633
rect 590 3628 596 3629
rect 678 3633 684 3634
rect 678 3629 679 3633
rect 683 3629 684 3633
rect 678 3628 684 3629
rect 110 3620 116 3621
rect 110 3616 111 3620
rect 115 3616 116 3620
rect 1822 3620 1828 3621
rect 1822 3616 1823 3620
rect 1827 3616 1828 3620
rect 110 3615 116 3616
rect 306 3615 312 3616
rect 306 3611 307 3615
rect 311 3614 312 3615
rect 394 3615 400 3616
rect 311 3612 345 3614
rect 311 3611 312 3612
rect 306 3610 312 3611
rect 394 3611 395 3615
rect 399 3614 400 3615
rect 482 3615 488 3616
rect 399 3612 433 3614
rect 399 3611 400 3612
rect 394 3610 400 3611
rect 482 3611 483 3615
rect 487 3614 488 3615
rect 570 3615 576 3616
rect 487 3612 521 3614
rect 487 3611 488 3612
rect 482 3610 488 3611
rect 570 3611 571 3615
rect 575 3614 576 3615
rect 658 3615 664 3616
rect 1822 3615 1828 3616
rect 575 3612 609 3614
rect 575 3611 576 3612
rect 570 3610 576 3611
rect 658 3611 659 3615
rect 663 3614 664 3615
rect 663 3612 697 3614
rect 663 3611 664 3612
rect 658 3610 664 3611
rect 110 3603 116 3604
rect 110 3599 111 3603
rect 115 3599 116 3603
rect 110 3598 116 3599
rect 1822 3603 1828 3604
rect 1822 3599 1823 3603
rect 1827 3599 1828 3603
rect 1822 3598 1828 3599
rect 230 3593 236 3594
rect 230 3589 231 3593
rect 235 3589 236 3593
rect 230 3588 236 3589
rect 318 3593 324 3594
rect 318 3589 319 3593
rect 323 3589 324 3593
rect 318 3588 324 3589
rect 406 3593 412 3594
rect 406 3589 407 3593
rect 411 3589 412 3593
rect 406 3588 412 3589
rect 494 3593 500 3594
rect 494 3589 495 3593
rect 499 3589 500 3593
rect 494 3588 500 3589
rect 582 3593 588 3594
rect 582 3589 583 3593
rect 587 3589 588 3593
rect 582 3588 588 3589
rect 670 3593 676 3594
rect 670 3589 671 3593
rect 675 3589 676 3593
rect 670 3588 676 3589
rect 279 3587 288 3588
rect 279 3583 280 3587
rect 287 3583 288 3587
rect 279 3582 288 3583
rect 1886 3575 1892 3576
rect 1886 3571 1887 3575
rect 1891 3571 1892 3575
rect 1886 3570 1892 3571
rect 1974 3575 1980 3576
rect 1974 3571 1975 3575
rect 1979 3571 1980 3575
rect 1974 3570 1980 3571
rect 2062 3575 2068 3576
rect 2062 3571 2063 3575
rect 2067 3571 2068 3575
rect 2062 3570 2068 3571
rect 2150 3575 2156 3576
rect 2150 3571 2151 3575
rect 2155 3571 2156 3575
rect 2150 3570 2156 3571
rect 2238 3575 2244 3576
rect 2238 3571 2239 3575
rect 2243 3571 2244 3575
rect 2238 3570 2244 3571
rect 2326 3575 2332 3576
rect 2326 3571 2327 3575
rect 2331 3571 2332 3575
rect 2326 3570 2332 3571
rect 2414 3575 2420 3576
rect 2414 3571 2415 3575
rect 2419 3571 2420 3575
rect 2414 3570 2420 3571
rect 2502 3575 2508 3576
rect 2502 3571 2503 3575
rect 2507 3571 2508 3575
rect 2502 3570 2508 3571
rect 2590 3575 2596 3576
rect 2590 3571 2591 3575
rect 2595 3571 2596 3575
rect 2590 3570 2596 3571
rect 2678 3575 2684 3576
rect 2678 3571 2679 3575
rect 2683 3571 2684 3575
rect 2678 3570 2684 3571
rect 2766 3575 2772 3576
rect 2766 3571 2767 3575
rect 2771 3571 2772 3575
rect 2766 3570 2772 3571
rect 2854 3575 2860 3576
rect 2854 3571 2855 3575
rect 2859 3571 2860 3575
rect 2854 3570 2860 3571
rect 2942 3575 2948 3576
rect 2942 3571 2943 3575
rect 2947 3571 2948 3575
rect 2942 3570 2948 3571
rect 3030 3575 3036 3576
rect 3030 3571 3031 3575
rect 3035 3571 3036 3575
rect 3030 3570 3036 3571
rect 3118 3575 3124 3576
rect 3118 3571 3119 3575
rect 3123 3571 3124 3575
rect 3118 3570 3124 3571
rect 3206 3575 3212 3576
rect 3206 3571 3207 3575
rect 3211 3571 3212 3575
rect 3206 3570 3212 3571
rect 3294 3575 3300 3576
rect 3294 3571 3295 3575
rect 3299 3571 3300 3575
rect 3294 3570 3300 3571
rect 3274 3567 3280 3568
rect 1862 3565 1868 3566
rect 246 3563 252 3564
rect 246 3559 247 3563
rect 251 3559 252 3563
rect 246 3558 252 3559
rect 398 3563 404 3564
rect 398 3559 399 3563
rect 403 3559 404 3563
rect 398 3558 404 3559
rect 542 3563 548 3564
rect 542 3559 543 3563
rect 547 3559 548 3563
rect 542 3558 548 3559
rect 686 3563 692 3564
rect 686 3559 687 3563
rect 691 3559 692 3563
rect 686 3558 692 3559
rect 822 3563 828 3564
rect 822 3559 823 3563
rect 827 3559 828 3563
rect 822 3558 828 3559
rect 950 3563 956 3564
rect 950 3559 951 3563
rect 955 3559 956 3563
rect 950 3558 956 3559
rect 1078 3563 1084 3564
rect 1078 3559 1079 3563
rect 1083 3559 1084 3563
rect 1078 3558 1084 3559
rect 1198 3563 1204 3564
rect 1198 3559 1199 3563
rect 1203 3559 1204 3563
rect 1198 3558 1204 3559
rect 1310 3563 1316 3564
rect 1310 3559 1311 3563
rect 1315 3559 1316 3563
rect 1310 3558 1316 3559
rect 1422 3563 1428 3564
rect 1422 3559 1423 3563
rect 1427 3559 1428 3563
rect 1422 3558 1428 3559
rect 1542 3563 1548 3564
rect 1542 3559 1543 3563
rect 1547 3559 1548 3563
rect 1862 3561 1863 3565
rect 1867 3561 1868 3565
rect 3274 3563 3275 3567
rect 3279 3566 3280 3567
rect 3279 3564 3313 3566
rect 3574 3565 3580 3566
rect 3279 3563 3280 3564
rect 3274 3562 3280 3563
rect 1862 3560 1868 3561
rect 3574 3561 3575 3565
rect 3579 3561 3580 3565
rect 3574 3560 3580 3561
rect 1542 3558 1548 3559
rect 1490 3555 1496 3556
rect 110 3553 116 3554
rect 110 3549 111 3553
rect 115 3549 116 3553
rect 1490 3551 1491 3555
rect 1495 3554 1496 3555
rect 1495 3552 1561 3554
rect 1822 3553 1828 3554
rect 1495 3551 1496 3552
rect 1490 3550 1496 3551
rect 110 3548 116 3549
rect 1822 3549 1823 3553
rect 1827 3549 1828 3553
rect 1967 3551 1973 3552
rect 1967 3550 1968 3551
rect 1822 3548 1828 3549
rect 1862 3548 1868 3549
rect 1949 3548 1968 3550
rect 1862 3544 1863 3548
rect 1867 3544 1868 3548
rect 1967 3547 1968 3548
rect 1972 3547 1973 3551
rect 2055 3551 2061 3552
rect 2055 3550 2056 3551
rect 2037 3548 2056 3550
rect 1967 3546 1973 3547
rect 2055 3547 2056 3548
rect 2060 3547 2061 3551
rect 2143 3551 2149 3552
rect 2143 3550 2144 3551
rect 2125 3548 2144 3550
rect 2055 3546 2061 3547
rect 2143 3547 2144 3548
rect 2148 3547 2149 3551
rect 2231 3551 2237 3552
rect 2231 3550 2232 3551
rect 2213 3548 2232 3550
rect 2143 3546 2149 3547
rect 2231 3547 2232 3548
rect 2236 3547 2237 3551
rect 2319 3551 2325 3552
rect 2319 3550 2320 3551
rect 2301 3548 2320 3550
rect 2231 3546 2237 3547
rect 2319 3547 2320 3548
rect 2324 3547 2325 3551
rect 2407 3551 2413 3552
rect 2407 3550 2408 3551
rect 2389 3548 2408 3550
rect 2319 3546 2325 3547
rect 2407 3547 2408 3548
rect 2412 3547 2413 3551
rect 2495 3551 2501 3552
rect 2495 3550 2496 3551
rect 2477 3548 2496 3550
rect 2407 3546 2413 3547
rect 2495 3547 2496 3548
rect 2500 3547 2501 3551
rect 2570 3551 2576 3552
rect 2570 3550 2571 3551
rect 2565 3548 2571 3550
rect 2495 3546 2501 3547
rect 2570 3547 2571 3548
rect 2575 3547 2576 3551
rect 2671 3551 2677 3552
rect 2671 3550 2672 3551
rect 2653 3548 2672 3550
rect 2570 3546 2576 3547
rect 2671 3547 2672 3548
rect 2676 3547 2677 3551
rect 2759 3551 2765 3552
rect 2759 3550 2760 3551
rect 2741 3548 2760 3550
rect 2671 3546 2677 3547
rect 2759 3547 2760 3548
rect 2764 3547 2765 3551
rect 2847 3551 2853 3552
rect 2847 3550 2848 3551
rect 2829 3548 2848 3550
rect 2759 3546 2765 3547
rect 2847 3547 2848 3548
rect 2852 3547 2853 3551
rect 2935 3551 2941 3552
rect 2935 3550 2936 3551
rect 2917 3548 2936 3550
rect 2847 3546 2853 3547
rect 2935 3547 2936 3548
rect 2940 3547 2941 3551
rect 3023 3551 3029 3552
rect 3023 3550 3024 3551
rect 3005 3548 3024 3550
rect 2935 3546 2941 3547
rect 3023 3547 3024 3548
rect 3028 3547 3029 3551
rect 3111 3551 3117 3552
rect 3111 3550 3112 3551
rect 3093 3548 3112 3550
rect 3023 3546 3029 3547
rect 3111 3547 3112 3548
rect 3116 3547 3117 3551
rect 3199 3551 3205 3552
rect 3199 3550 3200 3551
rect 3181 3548 3200 3550
rect 3111 3546 3117 3547
rect 3199 3547 3200 3548
rect 3204 3547 3205 3551
rect 3287 3551 3293 3552
rect 3287 3550 3288 3551
rect 3269 3548 3288 3550
rect 3199 3546 3205 3547
rect 3287 3547 3288 3548
rect 3292 3547 3293 3551
rect 3287 3546 3293 3547
rect 3574 3548 3580 3549
rect 1862 3543 1868 3544
rect 3574 3544 3575 3548
rect 3579 3544 3580 3548
rect 3574 3543 3580 3544
rect 391 3539 397 3540
rect 391 3538 392 3539
rect 110 3536 116 3537
rect 309 3536 392 3538
rect 110 3532 111 3536
rect 115 3532 116 3536
rect 391 3535 392 3536
rect 396 3535 397 3539
rect 535 3539 541 3540
rect 535 3538 536 3539
rect 461 3536 536 3538
rect 391 3534 397 3535
rect 535 3535 536 3536
rect 540 3535 541 3539
rect 679 3539 685 3540
rect 679 3538 680 3539
rect 605 3536 680 3538
rect 535 3534 541 3535
rect 679 3535 680 3536
rect 684 3535 685 3539
rect 754 3539 760 3540
rect 754 3538 755 3539
rect 749 3536 755 3538
rect 679 3534 685 3535
rect 754 3535 755 3536
rect 759 3535 760 3539
rect 943 3539 949 3540
rect 943 3538 944 3539
rect 885 3536 944 3538
rect 754 3534 760 3535
rect 943 3535 944 3536
rect 948 3535 949 3539
rect 1034 3539 1040 3540
rect 1034 3538 1035 3539
rect 1013 3536 1035 3538
rect 943 3534 949 3535
rect 1034 3535 1035 3536
rect 1039 3535 1040 3539
rect 1167 3539 1173 3540
rect 1167 3538 1168 3539
rect 1141 3536 1168 3538
rect 1034 3534 1040 3535
rect 1167 3535 1168 3536
rect 1172 3535 1173 3539
rect 1303 3539 1309 3540
rect 1303 3538 1304 3539
rect 1261 3536 1304 3538
rect 1167 3534 1173 3535
rect 1303 3535 1304 3536
rect 1308 3535 1309 3539
rect 1415 3539 1421 3540
rect 1415 3538 1416 3539
rect 1373 3536 1416 3538
rect 1303 3534 1309 3535
rect 1415 3535 1416 3536
rect 1420 3535 1421 3539
rect 1535 3539 1541 3540
rect 1535 3538 1536 3539
rect 1485 3536 1536 3538
rect 1415 3534 1421 3535
rect 1535 3535 1536 3536
rect 1540 3535 1541 3539
rect 1535 3534 1541 3535
rect 1822 3536 1828 3537
rect 110 3531 116 3532
rect 1822 3532 1823 3536
rect 1827 3532 1828 3536
rect 1822 3531 1828 3532
rect 1894 3535 1900 3536
rect 1894 3531 1895 3535
rect 1899 3531 1900 3535
rect 1894 3530 1900 3531
rect 1982 3535 1988 3536
rect 1982 3531 1983 3535
rect 1987 3531 1988 3535
rect 1982 3530 1988 3531
rect 2070 3535 2076 3536
rect 2070 3531 2071 3535
rect 2075 3531 2076 3535
rect 2070 3530 2076 3531
rect 2158 3535 2164 3536
rect 2158 3531 2159 3535
rect 2163 3531 2164 3535
rect 2158 3530 2164 3531
rect 2246 3535 2252 3536
rect 2246 3531 2247 3535
rect 2251 3531 2252 3535
rect 2246 3530 2252 3531
rect 2334 3535 2340 3536
rect 2334 3531 2335 3535
rect 2339 3531 2340 3535
rect 2334 3530 2340 3531
rect 2422 3535 2428 3536
rect 2422 3531 2423 3535
rect 2427 3531 2428 3535
rect 2422 3530 2428 3531
rect 2510 3535 2516 3536
rect 2510 3531 2511 3535
rect 2515 3531 2516 3535
rect 2510 3530 2516 3531
rect 2598 3535 2604 3536
rect 2598 3531 2599 3535
rect 2603 3531 2604 3535
rect 2598 3530 2604 3531
rect 2686 3535 2692 3536
rect 2686 3531 2687 3535
rect 2691 3531 2692 3535
rect 2686 3530 2692 3531
rect 2774 3535 2780 3536
rect 2774 3531 2775 3535
rect 2779 3531 2780 3535
rect 2774 3530 2780 3531
rect 2862 3535 2868 3536
rect 2862 3531 2863 3535
rect 2867 3531 2868 3535
rect 2862 3530 2868 3531
rect 2950 3535 2956 3536
rect 2950 3531 2951 3535
rect 2955 3531 2956 3535
rect 2950 3530 2956 3531
rect 3038 3535 3044 3536
rect 3038 3531 3039 3535
rect 3043 3531 3044 3535
rect 3038 3530 3044 3531
rect 3126 3535 3132 3536
rect 3126 3531 3127 3535
rect 3131 3531 3132 3535
rect 3126 3530 3132 3531
rect 3214 3535 3220 3536
rect 3214 3531 3215 3535
rect 3219 3531 3220 3535
rect 3214 3530 3220 3531
rect 3302 3535 3308 3536
rect 3302 3531 3303 3535
rect 3307 3531 3308 3535
rect 3302 3530 3308 3531
rect 254 3523 260 3524
rect 254 3519 255 3523
rect 259 3519 260 3523
rect 254 3518 260 3519
rect 406 3523 412 3524
rect 406 3519 407 3523
rect 411 3519 412 3523
rect 406 3518 412 3519
rect 550 3523 556 3524
rect 550 3519 551 3523
rect 555 3519 556 3523
rect 550 3518 556 3519
rect 694 3523 700 3524
rect 694 3519 695 3523
rect 699 3519 700 3523
rect 694 3518 700 3519
rect 830 3523 836 3524
rect 830 3519 831 3523
rect 835 3519 836 3523
rect 830 3518 836 3519
rect 958 3523 964 3524
rect 958 3519 959 3523
rect 963 3519 964 3523
rect 958 3518 964 3519
rect 1086 3523 1092 3524
rect 1086 3519 1087 3523
rect 1091 3519 1092 3523
rect 1086 3518 1092 3519
rect 1206 3523 1212 3524
rect 1206 3519 1207 3523
rect 1211 3519 1212 3523
rect 1206 3518 1212 3519
rect 1318 3523 1324 3524
rect 1318 3519 1319 3523
rect 1323 3519 1324 3523
rect 1318 3518 1324 3519
rect 1430 3523 1436 3524
rect 1430 3519 1431 3523
rect 1435 3519 1436 3523
rect 1430 3518 1436 3519
rect 1550 3523 1556 3524
rect 1550 3519 1551 3523
rect 1555 3519 1556 3523
rect 1550 3518 1556 3519
rect 1902 3523 1908 3524
rect 1902 3519 1903 3523
rect 1907 3522 1908 3523
rect 1923 3523 1929 3524
rect 1923 3522 1924 3523
rect 1907 3520 1924 3522
rect 1907 3519 1908 3520
rect 1902 3518 1908 3519
rect 1923 3519 1924 3520
rect 1928 3519 1929 3523
rect 1923 3518 1929 3519
rect 1967 3523 1973 3524
rect 1967 3519 1968 3523
rect 1972 3522 1973 3523
rect 2011 3523 2017 3524
rect 2011 3522 2012 3523
rect 1972 3520 2012 3522
rect 1972 3519 1973 3520
rect 1967 3518 1973 3519
rect 2011 3519 2012 3520
rect 2016 3519 2017 3523
rect 2011 3518 2017 3519
rect 2055 3523 2061 3524
rect 2055 3519 2056 3523
rect 2060 3522 2061 3523
rect 2099 3523 2105 3524
rect 2099 3522 2100 3523
rect 2060 3520 2100 3522
rect 2060 3519 2061 3520
rect 2055 3518 2061 3519
rect 2099 3519 2100 3520
rect 2104 3519 2105 3523
rect 2099 3518 2105 3519
rect 2143 3523 2149 3524
rect 2143 3519 2144 3523
rect 2148 3522 2149 3523
rect 2187 3523 2193 3524
rect 2187 3522 2188 3523
rect 2148 3520 2188 3522
rect 2148 3519 2149 3520
rect 2143 3518 2149 3519
rect 2187 3519 2188 3520
rect 2192 3519 2193 3523
rect 2187 3518 2193 3519
rect 2231 3523 2237 3524
rect 2231 3519 2232 3523
rect 2236 3522 2237 3523
rect 2275 3523 2281 3524
rect 2275 3522 2276 3523
rect 2236 3520 2276 3522
rect 2236 3519 2237 3520
rect 2231 3518 2237 3519
rect 2275 3519 2276 3520
rect 2280 3519 2281 3523
rect 2275 3518 2281 3519
rect 2319 3523 2325 3524
rect 2319 3519 2320 3523
rect 2324 3522 2325 3523
rect 2363 3523 2369 3524
rect 2363 3522 2364 3523
rect 2324 3520 2364 3522
rect 2324 3519 2325 3520
rect 2319 3518 2325 3519
rect 2363 3519 2364 3520
rect 2368 3519 2369 3523
rect 2363 3518 2369 3519
rect 2407 3523 2413 3524
rect 2407 3519 2408 3523
rect 2412 3522 2413 3523
rect 2451 3523 2457 3524
rect 2451 3522 2452 3523
rect 2412 3520 2452 3522
rect 2412 3519 2413 3520
rect 2407 3518 2413 3519
rect 2451 3519 2452 3520
rect 2456 3519 2457 3523
rect 2451 3518 2457 3519
rect 2495 3523 2501 3524
rect 2495 3519 2496 3523
rect 2500 3522 2501 3523
rect 2539 3523 2545 3524
rect 2539 3522 2540 3523
rect 2500 3520 2540 3522
rect 2500 3519 2501 3520
rect 2495 3518 2501 3519
rect 2539 3519 2540 3520
rect 2544 3519 2545 3523
rect 2539 3518 2545 3519
rect 2627 3523 2636 3524
rect 2627 3519 2628 3523
rect 2635 3519 2636 3523
rect 2627 3518 2636 3519
rect 2671 3523 2677 3524
rect 2671 3519 2672 3523
rect 2676 3522 2677 3523
rect 2715 3523 2721 3524
rect 2715 3522 2716 3523
rect 2676 3520 2716 3522
rect 2676 3519 2677 3520
rect 2671 3518 2677 3519
rect 2715 3519 2716 3520
rect 2720 3519 2721 3523
rect 2715 3518 2721 3519
rect 2759 3523 2765 3524
rect 2759 3519 2760 3523
rect 2764 3522 2765 3523
rect 2803 3523 2809 3524
rect 2803 3522 2804 3523
rect 2764 3520 2804 3522
rect 2764 3519 2765 3520
rect 2759 3518 2765 3519
rect 2803 3519 2804 3520
rect 2808 3519 2809 3523
rect 2803 3518 2809 3519
rect 2847 3523 2853 3524
rect 2847 3519 2848 3523
rect 2852 3522 2853 3523
rect 2891 3523 2897 3524
rect 2891 3522 2892 3523
rect 2852 3520 2892 3522
rect 2852 3519 2853 3520
rect 2847 3518 2853 3519
rect 2891 3519 2892 3520
rect 2896 3519 2897 3523
rect 2891 3518 2897 3519
rect 2935 3523 2941 3524
rect 2935 3519 2936 3523
rect 2940 3522 2941 3523
rect 2979 3523 2985 3524
rect 2979 3522 2980 3523
rect 2940 3520 2980 3522
rect 2940 3519 2941 3520
rect 2935 3518 2941 3519
rect 2979 3519 2980 3520
rect 2984 3519 2985 3523
rect 2979 3518 2985 3519
rect 3023 3523 3029 3524
rect 3023 3519 3024 3523
rect 3028 3522 3029 3523
rect 3067 3523 3073 3524
rect 3067 3522 3068 3523
rect 3028 3520 3068 3522
rect 3028 3519 3029 3520
rect 3023 3518 3029 3519
rect 3067 3519 3068 3520
rect 3072 3519 3073 3523
rect 3067 3518 3073 3519
rect 3111 3523 3117 3524
rect 3111 3519 3112 3523
rect 3116 3522 3117 3523
rect 3155 3523 3161 3524
rect 3155 3522 3156 3523
rect 3116 3520 3156 3522
rect 3116 3519 3117 3520
rect 3111 3518 3117 3519
rect 3155 3519 3156 3520
rect 3160 3519 3161 3523
rect 3155 3518 3161 3519
rect 3199 3523 3205 3524
rect 3199 3519 3200 3523
rect 3204 3522 3205 3523
rect 3243 3523 3249 3524
rect 3243 3522 3244 3523
rect 3204 3520 3244 3522
rect 3204 3519 3205 3520
rect 3199 3518 3205 3519
rect 3243 3519 3244 3520
rect 3248 3519 3249 3523
rect 3243 3518 3249 3519
rect 3287 3523 3293 3524
rect 3287 3519 3288 3523
rect 3292 3522 3293 3523
rect 3331 3523 3337 3524
rect 3331 3522 3332 3523
rect 3292 3520 3332 3522
rect 3292 3519 3293 3520
rect 3287 3518 3293 3519
rect 3331 3519 3332 3520
rect 3336 3519 3337 3523
rect 3331 3518 3337 3519
rect 282 3511 289 3512
rect 282 3507 283 3511
rect 288 3507 289 3511
rect 282 3506 289 3507
rect 391 3511 397 3512
rect 391 3507 392 3511
rect 396 3510 397 3511
rect 435 3511 441 3512
rect 435 3510 436 3511
rect 396 3508 436 3510
rect 396 3507 397 3508
rect 391 3506 397 3507
rect 435 3507 436 3508
rect 440 3507 441 3511
rect 435 3506 441 3507
rect 535 3511 541 3512
rect 535 3507 536 3511
rect 540 3510 541 3511
rect 579 3511 585 3512
rect 579 3510 580 3511
rect 540 3508 580 3510
rect 540 3507 541 3508
rect 535 3506 541 3507
rect 579 3507 580 3508
rect 584 3507 585 3511
rect 579 3506 585 3507
rect 679 3511 685 3512
rect 679 3507 680 3511
rect 684 3510 685 3511
rect 723 3511 729 3512
rect 723 3510 724 3511
rect 684 3508 724 3510
rect 684 3507 685 3508
rect 679 3506 685 3507
rect 723 3507 724 3508
rect 728 3507 729 3511
rect 723 3506 729 3507
rect 859 3511 865 3512
rect 859 3507 860 3511
rect 864 3510 865 3511
rect 890 3511 896 3512
rect 890 3510 891 3511
rect 864 3508 891 3510
rect 864 3507 865 3508
rect 859 3506 865 3507
rect 890 3507 891 3508
rect 895 3507 896 3511
rect 890 3506 896 3507
rect 943 3511 949 3512
rect 943 3507 944 3511
rect 948 3510 949 3511
rect 987 3511 993 3512
rect 987 3510 988 3511
rect 948 3508 988 3510
rect 948 3507 949 3508
rect 943 3506 949 3507
rect 987 3507 988 3508
rect 992 3507 993 3511
rect 987 3506 993 3507
rect 1034 3511 1040 3512
rect 1034 3507 1035 3511
rect 1039 3510 1040 3511
rect 1115 3511 1121 3512
rect 1115 3510 1116 3511
rect 1039 3508 1116 3510
rect 1039 3507 1040 3508
rect 1034 3506 1040 3507
rect 1115 3507 1116 3508
rect 1120 3507 1121 3511
rect 1115 3506 1121 3507
rect 1167 3511 1173 3512
rect 1167 3507 1168 3511
rect 1172 3510 1173 3511
rect 1235 3511 1241 3512
rect 1235 3510 1236 3511
rect 1172 3508 1236 3510
rect 1172 3507 1173 3508
rect 1167 3506 1173 3507
rect 1235 3507 1236 3508
rect 1240 3507 1241 3511
rect 1235 3506 1241 3507
rect 1303 3511 1309 3512
rect 1303 3507 1304 3511
rect 1308 3510 1309 3511
rect 1347 3511 1353 3512
rect 1347 3510 1348 3511
rect 1308 3508 1348 3510
rect 1308 3507 1309 3508
rect 1303 3506 1309 3507
rect 1347 3507 1348 3508
rect 1352 3507 1353 3511
rect 1347 3506 1353 3507
rect 1415 3511 1421 3512
rect 1415 3507 1416 3511
rect 1420 3510 1421 3511
rect 1459 3511 1465 3512
rect 1459 3510 1460 3511
rect 1420 3508 1460 3510
rect 1420 3507 1421 3508
rect 1415 3506 1421 3507
rect 1459 3507 1460 3508
rect 1464 3507 1465 3511
rect 1459 3506 1465 3507
rect 1535 3511 1541 3512
rect 1535 3507 1536 3511
rect 1540 3510 1541 3511
rect 1579 3511 1585 3512
rect 1579 3510 1580 3511
rect 1540 3508 1580 3510
rect 1540 3507 1541 3508
rect 1535 3506 1541 3507
rect 1579 3507 1580 3508
rect 1584 3507 1585 3511
rect 1579 3506 1585 3507
rect 1939 3503 1945 3504
rect 211 3499 217 3500
rect 211 3495 212 3499
rect 216 3498 217 3499
rect 255 3499 261 3500
rect 255 3498 256 3499
rect 216 3496 256 3498
rect 216 3495 217 3496
rect 211 3494 217 3495
rect 255 3495 256 3496
rect 260 3495 261 3499
rect 255 3494 261 3495
rect 379 3499 385 3500
rect 379 3495 380 3499
rect 384 3498 385 3499
rect 454 3499 460 3500
rect 454 3498 455 3499
rect 384 3496 455 3498
rect 384 3495 385 3496
rect 379 3494 385 3495
rect 454 3495 455 3496
rect 459 3495 460 3499
rect 454 3494 460 3495
rect 547 3499 553 3500
rect 547 3495 548 3499
rect 552 3498 553 3499
rect 607 3499 613 3500
rect 607 3498 608 3499
rect 552 3496 608 3498
rect 552 3495 553 3496
rect 547 3494 553 3495
rect 607 3495 608 3496
rect 612 3495 613 3499
rect 607 3494 613 3495
rect 707 3499 713 3500
rect 707 3495 708 3499
rect 712 3498 713 3499
rect 754 3499 760 3500
rect 754 3498 755 3499
rect 712 3496 755 3498
rect 712 3495 713 3496
rect 707 3494 713 3495
rect 754 3495 755 3496
rect 759 3495 760 3499
rect 754 3494 760 3495
rect 859 3499 865 3500
rect 859 3495 860 3499
rect 864 3498 865 3499
rect 978 3499 984 3500
rect 978 3498 979 3499
rect 864 3496 979 3498
rect 864 3495 865 3496
rect 859 3494 865 3495
rect 978 3495 979 3496
rect 983 3495 984 3499
rect 978 3494 984 3495
rect 995 3499 1001 3500
rect 995 3495 996 3499
rect 1000 3498 1001 3499
rect 1006 3499 1012 3500
rect 1006 3498 1007 3499
rect 1000 3496 1007 3498
rect 1000 3495 1001 3496
rect 995 3494 1001 3495
rect 1006 3495 1007 3496
rect 1011 3495 1012 3499
rect 1006 3494 1012 3495
rect 1039 3499 1045 3500
rect 1039 3495 1040 3499
rect 1044 3498 1045 3499
rect 1123 3499 1129 3500
rect 1123 3498 1124 3499
rect 1044 3496 1124 3498
rect 1044 3495 1045 3496
rect 1039 3494 1045 3495
rect 1123 3495 1124 3496
rect 1128 3495 1129 3499
rect 1123 3494 1129 3495
rect 1243 3499 1252 3500
rect 1243 3495 1244 3499
rect 1251 3495 1252 3499
rect 1243 3494 1252 3495
rect 1295 3499 1301 3500
rect 1295 3495 1296 3499
rect 1300 3498 1301 3499
rect 1363 3499 1369 3500
rect 1363 3498 1364 3499
rect 1300 3496 1364 3498
rect 1300 3495 1301 3496
rect 1295 3494 1301 3495
rect 1363 3495 1364 3496
rect 1368 3495 1369 3499
rect 1363 3494 1369 3495
rect 1415 3499 1421 3500
rect 1415 3495 1416 3499
rect 1420 3498 1421 3499
rect 1483 3499 1489 3500
rect 1483 3498 1484 3499
rect 1420 3496 1484 3498
rect 1420 3495 1421 3496
rect 1415 3494 1421 3495
rect 1483 3495 1484 3496
rect 1488 3495 1489 3499
rect 1483 3494 1489 3495
rect 1519 3499 1525 3500
rect 1519 3495 1520 3499
rect 1524 3498 1525 3499
rect 1603 3499 1609 3500
rect 1603 3498 1604 3499
rect 1524 3496 1604 3498
rect 1524 3495 1525 3496
rect 1519 3494 1525 3495
rect 1603 3495 1604 3496
rect 1608 3495 1609 3499
rect 1939 3499 1940 3503
rect 1944 3502 1945 3503
rect 1983 3503 1989 3504
rect 1983 3502 1984 3503
rect 1944 3500 1984 3502
rect 1944 3499 1945 3500
rect 1939 3498 1945 3499
rect 1983 3499 1984 3500
rect 1988 3499 1989 3503
rect 1983 3498 1989 3499
rect 2043 3503 2049 3504
rect 2043 3499 2044 3503
rect 2048 3502 2049 3503
rect 2082 3503 2088 3504
rect 2082 3502 2083 3503
rect 2048 3500 2083 3502
rect 2048 3499 2049 3500
rect 2043 3498 2049 3499
rect 2082 3499 2083 3500
rect 2087 3499 2088 3503
rect 2082 3498 2088 3499
rect 2142 3503 2148 3504
rect 2142 3499 2143 3503
rect 2147 3502 2148 3503
rect 2163 3503 2169 3504
rect 2163 3502 2164 3503
rect 2147 3500 2164 3502
rect 2147 3499 2148 3500
rect 2142 3498 2148 3499
rect 2163 3499 2164 3500
rect 2168 3499 2169 3503
rect 2163 3498 2169 3499
rect 2291 3503 2297 3504
rect 2291 3499 2292 3503
rect 2296 3502 2297 3503
rect 2350 3503 2356 3504
rect 2350 3502 2351 3503
rect 2296 3500 2351 3502
rect 2296 3499 2297 3500
rect 2291 3498 2297 3499
rect 2350 3499 2351 3500
rect 2355 3499 2356 3503
rect 2350 3498 2356 3499
rect 2419 3503 2425 3504
rect 2419 3499 2420 3503
rect 2424 3502 2425 3503
rect 2458 3503 2464 3504
rect 2458 3502 2459 3503
rect 2424 3500 2459 3502
rect 2424 3499 2425 3500
rect 2419 3498 2425 3499
rect 2458 3499 2459 3500
rect 2463 3499 2464 3503
rect 2458 3498 2464 3499
rect 2555 3503 2561 3504
rect 2555 3499 2556 3503
rect 2560 3502 2561 3503
rect 2570 3503 2576 3504
rect 2570 3502 2571 3503
rect 2560 3500 2571 3502
rect 2560 3499 2561 3500
rect 2555 3498 2561 3499
rect 2570 3499 2571 3500
rect 2575 3499 2576 3503
rect 2570 3498 2576 3499
rect 2691 3503 2697 3504
rect 2691 3499 2692 3503
rect 2696 3502 2697 3503
rect 2702 3503 2708 3504
rect 2702 3502 2703 3503
rect 2696 3500 2703 3502
rect 2696 3499 2697 3500
rect 2691 3498 2697 3499
rect 2702 3499 2703 3500
rect 2707 3499 2708 3503
rect 2702 3498 2708 3499
rect 2827 3503 2833 3504
rect 2827 3499 2828 3503
rect 2832 3502 2833 3503
rect 2890 3503 2896 3504
rect 2890 3502 2891 3503
rect 2832 3500 2891 3502
rect 2832 3499 2833 3500
rect 2827 3498 2833 3499
rect 2890 3499 2891 3500
rect 2895 3499 2896 3503
rect 2890 3498 2896 3499
rect 2971 3503 2977 3504
rect 2971 3499 2972 3503
rect 2976 3502 2977 3503
rect 3031 3503 3037 3504
rect 3031 3502 3032 3503
rect 2976 3500 3032 3502
rect 2976 3499 2977 3500
rect 2971 3498 2977 3499
rect 3031 3499 3032 3500
rect 3036 3499 3037 3503
rect 3031 3498 3037 3499
rect 3115 3503 3121 3504
rect 3115 3499 3116 3503
rect 3120 3502 3121 3503
rect 3274 3503 3280 3504
rect 3274 3502 3275 3503
rect 3120 3500 3275 3502
rect 3120 3499 3121 3500
rect 3115 3498 3121 3499
rect 3274 3499 3275 3500
rect 3279 3499 3280 3503
rect 3274 3498 3280 3499
rect 1603 3494 1609 3495
rect 1910 3493 1916 3494
rect 182 3489 188 3490
rect 182 3485 183 3489
rect 187 3485 188 3489
rect 182 3484 188 3485
rect 350 3489 356 3490
rect 350 3485 351 3489
rect 355 3485 356 3489
rect 350 3484 356 3485
rect 518 3489 524 3490
rect 518 3485 519 3489
rect 523 3485 524 3489
rect 518 3484 524 3485
rect 678 3489 684 3490
rect 678 3485 679 3489
rect 683 3485 684 3489
rect 678 3484 684 3485
rect 830 3489 836 3490
rect 830 3485 831 3489
rect 835 3485 836 3489
rect 830 3484 836 3485
rect 966 3489 972 3490
rect 966 3485 967 3489
rect 971 3485 972 3489
rect 966 3484 972 3485
rect 1094 3489 1100 3490
rect 1094 3485 1095 3489
rect 1099 3485 1100 3489
rect 1094 3484 1100 3485
rect 1214 3489 1220 3490
rect 1214 3485 1215 3489
rect 1219 3485 1220 3489
rect 1214 3484 1220 3485
rect 1334 3489 1340 3490
rect 1334 3485 1335 3489
rect 1339 3485 1340 3489
rect 1334 3484 1340 3485
rect 1454 3489 1460 3490
rect 1454 3485 1455 3489
rect 1459 3485 1460 3489
rect 1454 3484 1460 3485
rect 1574 3489 1580 3490
rect 1574 3485 1575 3489
rect 1579 3485 1580 3489
rect 1910 3489 1911 3493
rect 1915 3489 1916 3493
rect 1910 3488 1916 3489
rect 2014 3493 2020 3494
rect 2014 3489 2015 3493
rect 2019 3489 2020 3493
rect 2014 3488 2020 3489
rect 2134 3493 2140 3494
rect 2134 3489 2135 3493
rect 2139 3489 2140 3493
rect 2134 3488 2140 3489
rect 2262 3493 2268 3494
rect 2262 3489 2263 3493
rect 2267 3489 2268 3493
rect 2262 3488 2268 3489
rect 2390 3493 2396 3494
rect 2390 3489 2391 3493
rect 2395 3489 2396 3493
rect 2390 3488 2396 3489
rect 2526 3493 2532 3494
rect 2526 3489 2527 3493
rect 2531 3489 2532 3493
rect 2526 3488 2532 3489
rect 2662 3493 2668 3494
rect 2662 3489 2663 3493
rect 2667 3489 2668 3493
rect 2662 3488 2668 3489
rect 2798 3493 2804 3494
rect 2798 3489 2799 3493
rect 2803 3489 2804 3493
rect 2798 3488 2804 3489
rect 2942 3493 2948 3494
rect 2942 3489 2943 3493
rect 2947 3489 2948 3493
rect 2942 3488 2948 3489
rect 3086 3493 3092 3494
rect 3086 3489 3087 3493
rect 3091 3489 3092 3493
rect 3086 3488 3092 3489
rect 1574 3484 1580 3485
rect 1862 3480 1868 3481
rect 110 3476 116 3477
rect 1822 3476 1828 3477
rect 110 3472 111 3476
rect 115 3472 116 3476
rect 890 3475 896 3476
rect 890 3474 891 3475
rect 885 3472 891 3474
rect 110 3471 116 3472
rect 255 3471 261 3472
rect 255 3467 256 3471
rect 260 3470 261 3471
rect 454 3471 460 3472
rect 260 3468 369 3470
rect 260 3467 261 3468
rect 255 3466 261 3467
rect 454 3467 455 3471
rect 459 3470 460 3471
rect 607 3471 613 3472
rect 459 3468 537 3470
rect 459 3467 460 3468
rect 454 3466 460 3467
rect 607 3467 608 3471
rect 612 3470 613 3471
rect 890 3471 891 3472
rect 895 3471 896 3475
rect 1039 3475 1045 3476
rect 1039 3474 1040 3475
rect 1021 3472 1040 3474
rect 890 3470 896 3471
rect 1039 3471 1040 3472
rect 1044 3471 1045 3475
rect 1295 3475 1301 3476
rect 1295 3474 1296 3475
rect 1269 3472 1296 3474
rect 1039 3470 1045 3471
rect 1295 3471 1296 3472
rect 1300 3471 1301 3475
rect 1415 3475 1421 3476
rect 1415 3474 1416 3475
rect 1389 3472 1416 3474
rect 1295 3470 1301 3471
rect 1415 3471 1416 3472
rect 1420 3471 1421 3475
rect 1519 3475 1525 3476
rect 1519 3474 1520 3475
rect 1509 3472 1520 3474
rect 1415 3470 1421 3471
rect 1519 3471 1520 3472
rect 1524 3471 1525 3475
rect 1822 3472 1823 3476
rect 1827 3472 1828 3476
rect 1862 3476 1863 3480
rect 1867 3476 1868 3480
rect 3574 3480 3580 3481
rect 3574 3476 3575 3480
rect 3579 3476 3580 3480
rect 1862 3475 1868 3476
rect 1902 3475 1908 3476
rect 1822 3471 1828 3472
rect 1902 3471 1903 3475
rect 1907 3474 1908 3475
rect 1983 3475 1989 3476
rect 1907 3472 1929 3474
rect 1907 3471 1908 3472
rect 1519 3470 1525 3471
rect 1902 3470 1908 3471
rect 1983 3471 1984 3475
rect 1988 3474 1989 3475
rect 2082 3475 2088 3476
rect 1988 3472 2033 3474
rect 1988 3471 1989 3472
rect 1983 3470 1989 3471
rect 2082 3471 2083 3475
rect 2087 3474 2088 3475
rect 2350 3475 2356 3476
rect 2087 3472 2153 3474
rect 2087 3471 2088 3472
rect 2082 3470 2088 3471
rect 2350 3471 2351 3475
rect 2355 3474 2356 3475
rect 2458 3475 2464 3476
rect 2355 3472 2409 3474
rect 2355 3471 2356 3472
rect 2350 3470 2356 3471
rect 2458 3471 2459 3475
rect 2463 3474 2464 3475
rect 2630 3475 2636 3476
rect 2463 3472 2545 3474
rect 2463 3471 2464 3472
rect 2458 3470 2464 3471
rect 2630 3471 2631 3475
rect 2635 3474 2636 3475
rect 2890 3475 2896 3476
rect 2635 3472 2681 3474
rect 2635 3471 2636 3472
rect 2630 3470 2636 3471
rect 2890 3471 2891 3475
rect 2895 3474 2896 3475
rect 3031 3475 3037 3476
rect 3574 3475 3580 3476
rect 2895 3472 2961 3474
rect 2895 3471 2896 3472
rect 2890 3470 2896 3471
rect 3031 3471 3032 3475
rect 3036 3474 3037 3475
rect 3036 3472 3105 3474
rect 3036 3471 3037 3472
rect 3031 3470 3037 3471
rect 612 3468 697 3470
rect 612 3467 613 3468
rect 607 3466 613 3467
rect 1862 3463 1868 3464
rect 110 3459 116 3460
rect 110 3455 111 3459
rect 115 3455 116 3459
rect 270 3459 276 3460
rect 270 3458 271 3459
rect 233 3456 271 3458
rect 110 3454 116 3455
rect 270 3455 271 3456
rect 275 3455 276 3459
rect 1822 3459 1828 3460
rect 270 3454 276 3455
rect 1028 3456 1105 3458
rect 1516 3456 1585 3458
rect 174 3449 180 3450
rect 174 3445 175 3449
rect 179 3445 180 3449
rect 174 3444 180 3445
rect 342 3449 348 3450
rect 342 3445 343 3449
rect 347 3445 348 3449
rect 342 3444 348 3445
rect 510 3449 516 3450
rect 510 3445 511 3449
rect 515 3445 516 3449
rect 510 3444 516 3445
rect 670 3449 676 3450
rect 670 3445 671 3449
rect 675 3445 676 3449
rect 670 3444 676 3445
rect 822 3449 828 3450
rect 822 3445 823 3449
rect 827 3445 828 3449
rect 822 3444 828 3445
rect 958 3449 964 3450
rect 958 3445 959 3449
rect 963 3445 964 3449
rect 958 3444 964 3445
rect 978 3443 984 3444
rect 978 3439 979 3443
rect 983 3442 984 3443
rect 1028 3442 1030 3456
rect 1086 3449 1092 3450
rect 1086 3445 1087 3449
rect 1091 3445 1092 3449
rect 1086 3444 1092 3445
rect 1206 3449 1212 3450
rect 1206 3445 1207 3449
rect 1211 3445 1212 3449
rect 1206 3444 1212 3445
rect 1326 3449 1332 3450
rect 1326 3445 1327 3449
rect 1331 3445 1332 3449
rect 1326 3444 1332 3445
rect 1446 3449 1452 3450
rect 1446 3445 1447 3449
rect 1451 3445 1452 3449
rect 1446 3444 1452 3445
rect 983 3440 1030 3442
rect 1334 3443 1340 3444
rect 983 3439 984 3440
rect 978 3438 984 3439
rect 1334 3439 1335 3443
rect 1339 3442 1340 3443
rect 1516 3442 1518 3456
rect 1822 3455 1823 3459
rect 1827 3455 1828 3459
rect 1862 3459 1863 3463
rect 1867 3459 1868 3463
rect 2390 3463 2396 3464
rect 2390 3462 2391 3463
rect 2313 3460 2391 3462
rect 1862 3458 1868 3459
rect 2390 3459 2391 3460
rect 2395 3459 2396 3463
rect 2390 3458 2396 3459
rect 2798 3463 2804 3464
rect 2798 3459 2799 3463
rect 2803 3462 2804 3463
rect 3574 3463 3580 3464
rect 2803 3460 2809 3462
rect 2803 3459 2804 3460
rect 2798 3458 2804 3459
rect 3574 3459 3575 3463
rect 3579 3459 3580 3463
rect 3574 3458 3580 3459
rect 1822 3454 1828 3455
rect 1902 3453 1908 3454
rect 1566 3449 1572 3450
rect 1566 3445 1567 3449
rect 1571 3445 1572 3449
rect 1902 3449 1903 3453
rect 1907 3449 1908 3453
rect 1902 3448 1908 3449
rect 2006 3453 2012 3454
rect 2006 3449 2007 3453
rect 2011 3449 2012 3453
rect 2006 3448 2012 3449
rect 2126 3453 2132 3454
rect 2126 3449 2127 3453
rect 2131 3449 2132 3453
rect 2126 3448 2132 3449
rect 2254 3453 2260 3454
rect 2254 3449 2255 3453
rect 2259 3449 2260 3453
rect 2254 3448 2260 3449
rect 2382 3453 2388 3454
rect 2382 3449 2383 3453
rect 2387 3449 2388 3453
rect 2382 3448 2388 3449
rect 2518 3453 2524 3454
rect 2518 3449 2519 3453
rect 2523 3449 2524 3453
rect 2518 3448 2524 3449
rect 2654 3453 2660 3454
rect 2654 3449 2655 3453
rect 2659 3449 2660 3453
rect 2654 3448 2660 3449
rect 2790 3453 2796 3454
rect 2790 3449 2791 3453
rect 2795 3449 2796 3453
rect 2790 3448 2796 3449
rect 2934 3453 2940 3454
rect 2934 3449 2935 3453
rect 2939 3449 2940 3453
rect 2934 3448 2940 3449
rect 3078 3453 3084 3454
rect 3078 3449 3079 3453
rect 3083 3449 3084 3453
rect 3078 3448 3084 3449
rect 1566 3444 1572 3445
rect 1339 3440 1518 3442
rect 1339 3439 1340 3440
rect 1334 3438 1340 3439
rect 134 3427 140 3428
rect 134 3423 135 3427
rect 139 3423 140 3427
rect 134 3422 140 3423
rect 254 3427 260 3428
rect 254 3423 255 3427
rect 259 3423 260 3427
rect 254 3422 260 3423
rect 414 3427 420 3428
rect 414 3423 415 3427
rect 419 3423 420 3427
rect 414 3422 420 3423
rect 582 3427 588 3428
rect 582 3423 583 3427
rect 587 3423 588 3427
rect 582 3422 588 3423
rect 758 3427 764 3428
rect 758 3423 759 3427
rect 763 3423 764 3427
rect 758 3422 764 3423
rect 934 3427 940 3428
rect 934 3423 935 3427
rect 939 3423 940 3427
rect 934 3422 940 3423
rect 1110 3427 1116 3428
rect 1110 3423 1111 3427
rect 1115 3423 1116 3427
rect 1110 3422 1116 3423
rect 1294 3427 1300 3428
rect 1294 3423 1295 3427
rect 1299 3423 1300 3427
rect 1294 3422 1300 3423
rect 1478 3427 1484 3428
rect 1478 3423 1479 3427
rect 1483 3423 1484 3427
rect 1478 3422 1484 3423
rect 1910 3423 1916 3424
rect 678 3419 684 3420
rect 110 3417 116 3418
rect 110 3413 111 3417
rect 115 3413 116 3417
rect 678 3415 679 3419
rect 683 3418 684 3419
rect 1006 3419 1012 3420
rect 1006 3418 1007 3419
rect 683 3416 777 3418
rect 993 3416 1007 3418
rect 683 3415 684 3416
rect 678 3414 684 3415
rect 1006 3415 1007 3416
rect 1011 3415 1012 3419
rect 1910 3419 1911 3423
rect 1915 3419 1916 3423
rect 1910 3418 1916 3419
rect 2070 3423 2076 3424
rect 2070 3419 2071 3423
rect 2075 3419 2076 3423
rect 2070 3418 2076 3419
rect 2222 3423 2228 3424
rect 2222 3419 2223 3423
rect 2227 3419 2228 3423
rect 2222 3418 2228 3419
rect 2366 3423 2372 3424
rect 2366 3419 2367 3423
rect 2371 3419 2372 3423
rect 2366 3418 2372 3419
rect 2502 3423 2508 3424
rect 2502 3419 2503 3423
rect 2507 3419 2508 3423
rect 2502 3418 2508 3419
rect 2630 3423 2636 3424
rect 2630 3419 2631 3423
rect 2635 3419 2636 3423
rect 2630 3418 2636 3419
rect 2758 3423 2764 3424
rect 2758 3419 2759 3423
rect 2763 3419 2764 3423
rect 2758 3418 2764 3419
rect 2886 3423 2892 3424
rect 2886 3419 2887 3423
rect 2891 3419 2892 3423
rect 2886 3418 2892 3419
rect 3022 3423 3028 3424
rect 3022 3419 3023 3423
rect 3027 3419 3028 3423
rect 3022 3418 3028 3419
rect 1006 3414 1012 3415
rect 1822 3417 1828 3418
rect 110 3412 116 3413
rect 1822 3413 1823 3417
rect 1827 3413 1828 3417
rect 2142 3415 2148 3416
rect 2142 3414 2143 3415
rect 1822 3412 1828 3413
rect 1862 3413 1868 3414
rect 1862 3409 1863 3413
rect 1867 3409 1868 3413
rect 2129 3412 2143 3414
rect 2142 3411 2143 3412
rect 2147 3411 2148 3415
rect 2702 3415 2708 3416
rect 2702 3414 2703 3415
rect 2689 3412 2703 3414
rect 2142 3410 2148 3411
rect 2702 3411 2703 3412
rect 2707 3411 2708 3415
rect 2702 3410 2708 3411
rect 3574 3413 3580 3414
rect 1862 3408 1868 3409
rect 3574 3409 3575 3413
rect 3579 3409 3580 3413
rect 3574 3408 3580 3409
rect 218 3403 224 3404
rect 218 3402 219 3403
rect 110 3400 116 3401
rect 197 3400 219 3402
rect 110 3396 111 3400
rect 115 3396 116 3400
rect 218 3399 219 3400
rect 223 3399 224 3403
rect 407 3403 413 3404
rect 407 3402 408 3403
rect 317 3400 408 3402
rect 218 3398 224 3399
rect 407 3399 408 3400
rect 412 3399 413 3403
rect 575 3403 581 3404
rect 575 3402 576 3403
rect 477 3400 576 3402
rect 407 3398 413 3399
rect 575 3399 576 3400
rect 580 3399 581 3403
rect 751 3403 757 3404
rect 751 3402 752 3403
rect 645 3400 752 3402
rect 575 3398 581 3399
rect 751 3399 752 3400
rect 756 3399 757 3403
rect 751 3398 757 3399
rect 1002 3403 1008 3404
rect 1002 3399 1003 3403
rect 1007 3402 1008 3403
rect 1471 3403 1477 3404
rect 1471 3402 1472 3403
rect 1007 3400 1137 3402
rect 1357 3400 1472 3402
rect 1007 3399 1008 3400
rect 1002 3398 1008 3399
rect 1471 3399 1472 3400
rect 1476 3399 1477 3403
rect 1586 3403 1592 3404
rect 1586 3402 1587 3403
rect 1541 3400 1587 3402
rect 1471 3398 1477 3399
rect 1586 3399 1587 3400
rect 1591 3399 1592 3403
rect 1586 3398 1592 3399
rect 1822 3400 1828 3401
rect 110 3395 116 3396
rect 1822 3396 1823 3400
rect 1827 3396 1828 3400
rect 2063 3399 2069 3400
rect 2063 3398 2064 3399
rect 1822 3395 1828 3396
rect 1862 3396 1868 3397
rect 1973 3396 2064 3398
rect 1862 3392 1863 3396
rect 1867 3392 1868 3396
rect 2063 3395 2064 3396
rect 2068 3395 2069 3399
rect 2063 3394 2069 3395
rect 2214 3399 2220 3400
rect 2214 3395 2215 3399
rect 2219 3398 2220 3399
rect 2290 3399 2296 3400
rect 2219 3396 2249 3398
rect 2219 3395 2220 3396
rect 2214 3394 2220 3395
rect 2290 3395 2291 3399
rect 2295 3398 2296 3399
rect 2623 3399 2629 3400
rect 2623 3398 2624 3399
rect 2295 3396 2393 3398
rect 2565 3396 2624 3398
rect 2295 3395 2296 3396
rect 2290 3394 2296 3395
rect 2623 3395 2624 3396
rect 2628 3395 2629 3399
rect 2842 3399 2848 3400
rect 2842 3398 2843 3399
rect 2821 3396 2843 3398
rect 2623 3394 2629 3395
rect 2842 3395 2843 3396
rect 2847 3395 2848 3399
rect 3015 3399 3021 3400
rect 3015 3398 3016 3399
rect 2949 3396 3016 3398
rect 2842 3394 2848 3395
rect 3015 3395 3016 3396
rect 3020 3395 3021 3399
rect 3090 3399 3096 3400
rect 3090 3398 3091 3399
rect 3085 3396 3091 3398
rect 3015 3394 3021 3395
rect 3090 3395 3091 3396
rect 3095 3395 3096 3399
rect 3090 3394 3096 3395
rect 3574 3396 3580 3397
rect 1862 3391 1868 3392
rect 3574 3392 3575 3396
rect 3579 3392 3580 3396
rect 3574 3391 3580 3392
rect 142 3387 148 3388
rect 142 3383 143 3387
rect 147 3383 148 3387
rect 142 3382 148 3383
rect 262 3387 268 3388
rect 262 3383 263 3387
rect 267 3383 268 3387
rect 262 3382 268 3383
rect 422 3387 428 3388
rect 422 3383 423 3387
rect 427 3383 428 3387
rect 422 3382 428 3383
rect 590 3387 596 3388
rect 590 3383 591 3387
rect 595 3383 596 3387
rect 590 3382 596 3383
rect 766 3387 772 3388
rect 766 3383 767 3387
rect 771 3383 772 3387
rect 766 3382 772 3383
rect 942 3387 948 3388
rect 942 3383 943 3387
rect 947 3383 948 3387
rect 942 3382 948 3383
rect 1118 3387 1124 3388
rect 1118 3383 1119 3387
rect 1123 3383 1124 3387
rect 1118 3382 1124 3383
rect 1302 3387 1308 3388
rect 1302 3383 1303 3387
rect 1307 3383 1308 3387
rect 1302 3382 1308 3383
rect 1486 3387 1492 3388
rect 1486 3383 1487 3387
rect 1491 3383 1492 3387
rect 1486 3382 1492 3383
rect 1918 3383 1924 3384
rect 1918 3379 1919 3383
rect 1923 3379 1924 3383
rect 1918 3378 1924 3379
rect 2078 3383 2084 3384
rect 2078 3379 2079 3383
rect 2083 3379 2084 3383
rect 2078 3378 2084 3379
rect 2230 3383 2236 3384
rect 2230 3379 2231 3383
rect 2235 3379 2236 3383
rect 2230 3378 2236 3379
rect 2374 3383 2380 3384
rect 2374 3379 2375 3383
rect 2379 3379 2380 3383
rect 2374 3378 2380 3379
rect 2510 3383 2516 3384
rect 2510 3379 2511 3383
rect 2515 3379 2516 3383
rect 2510 3378 2516 3379
rect 2638 3383 2644 3384
rect 2638 3379 2639 3383
rect 2643 3379 2644 3383
rect 2638 3378 2644 3379
rect 2766 3383 2772 3384
rect 2766 3379 2767 3383
rect 2771 3379 2772 3383
rect 2766 3378 2772 3379
rect 2894 3383 2900 3384
rect 2894 3379 2895 3383
rect 2899 3379 2900 3383
rect 2894 3378 2900 3379
rect 3030 3383 3036 3384
rect 3030 3379 3031 3383
rect 3035 3379 3036 3383
rect 3030 3378 3036 3379
rect 171 3375 177 3376
rect 171 3371 172 3375
rect 176 3374 177 3375
rect 270 3375 276 3376
rect 270 3374 271 3375
rect 176 3372 271 3374
rect 176 3371 177 3372
rect 171 3370 177 3371
rect 270 3371 271 3372
rect 275 3371 276 3375
rect 291 3375 297 3376
rect 291 3374 292 3375
rect 270 3370 276 3371
rect 280 3372 292 3374
rect 218 3367 224 3368
rect 218 3363 219 3367
rect 223 3366 224 3367
rect 280 3366 282 3372
rect 291 3371 292 3372
rect 296 3371 297 3375
rect 291 3370 297 3371
rect 407 3375 413 3376
rect 407 3371 408 3375
rect 412 3374 413 3375
rect 451 3375 457 3376
rect 451 3374 452 3375
rect 412 3372 452 3374
rect 412 3371 413 3372
rect 407 3370 413 3371
rect 451 3371 452 3372
rect 456 3371 457 3375
rect 451 3370 457 3371
rect 575 3375 581 3376
rect 575 3371 576 3375
rect 580 3374 581 3375
rect 619 3375 625 3376
rect 619 3374 620 3375
rect 580 3372 620 3374
rect 580 3371 581 3372
rect 575 3370 581 3371
rect 619 3371 620 3372
rect 624 3371 625 3375
rect 619 3370 625 3371
rect 751 3375 757 3376
rect 751 3371 752 3375
rect 756 3374 757 3375
rect 795 3375 801 3376
rect 795 3374 796 3375
rect 756 3372 796 3374
rect 756 3371 757 3372
rect 751 3370 757 3371
rect 795 3371 796 3372
rect 800 3371 801 3375
rect 795 3370 801 3371
rect 971 3375 977 3376
rect 971 3371 972 3375
rect 976 3374 977 3375
rect 1002 3375 1008 3376
rect 1002 3374 1003 3375
rect 976 3372 1003 3374
rect 976 3371 977 3372
rect 971 3370 977 3371
rect 1002 3371 1003 3372
rect 1007 3371 1008 3375
rect 1002 3370 1008 3371
rect 1134 3375 1140 3376
rect 1134 3371 1135 3375
rect 1139 3374 1140 3375
rect 1147 3375 1153 3376
rect 1147 3374 1148 3375
rect 1139 3372 1148 3374
rect 1139 3371 1140 3372
rect 1134 3370 1140 3371
rect 1147 3371 1148 3372
rect 1152 3371 1153 3375
rect 1147 3370 1153 3371
rect 1331 3375 1340 3376
rect 1331 3371 1332 3375
rect 1339 3371 1340 3375
rect 1331 3370 1340 3371
rect 1471 3375 1477 3376
rect 1471 3371 1472 3375
rect 1476 3374 1477 3375
rect 1515 3375 1521 3376
rect 1515 3374 1516 3375
rect 1476 3372 1516 3374
rect 1476 3371 1477 3372
rect 1471 3370 1477 3371
rect 1515 3371 1516 3372
rect 1520 3371 1521 3375
rect 1515 3370 1521 3371
rect 1947 3371 1956 3372
rect 1947 3367 1948 3371
rect 1955 3367 1956 3371
rect 1947 3366 1956 3367
rect 2063 3371 2069 3372
rect 2063 3367 2064 3371
rect 2068 3370 2069 3371
rect 2107 3371 2113 3372
rect 2107 3370 2108 3371
rect 2068 3368 2108 3370
rect 2068 3367 2069 3368
rect 2063 3366 2069 3367
rect 2107 3367 2108 3368
rect 2112 3367 2113 3371
rect 2107 3366 2113 3367
rect 2259 3371 2265 3372
rect 2259 3367 2260 3371
rect 2264 3370 2265 3371
rect 2290 3371 2296 3372
rect 2290 3370 2291 3371
rect 2264 3368 2291 3370
rect 2264 3367 2265 3368
rect 2259 3366 2265 3367
rect 2290 3367 2291 3368
rect 2295 3367 2296 3371
rect 2290 3366 2296 3367
rect 2390 3371 2396 3372
rect 2390 3367 2391 3371
rect 2395 3370 2396 3371
rect 2403 3371 2409 3372
rect 2403 3370 2404 3371
rect 2395 3368 2404 3370
rect 2395 3367 2396 3368
rect 2390 3366 2396 3367
rect 2403 3367 2404 3368
rect 2408 3367 2409 3371
rect 2403 3366 2409 3367
rect 2539 3371 2545 3372
rect 2539 3367 2540 3371
rect 2544 3370 2545 3371
rect 2602 3371 2608 3372
rect 2602 3370 2603 3371
rect 2544 3368 2603 3370
rect 2544 3367 2545 3368
rect 2539 3366 2545 3367
rect 2602 3367 2603 3368
rect 2607 3367 2608 3371
rect 2602 3366 2608 3367
rect 2623 3371 2629 3372
rect 2623 3367 2624 3371
rect 2628 3370 2629 3371
rect 2667 3371 2673 3372
rect 2667 3370 2668 3371
rect 2628 3368 2668 3370
rect 2628 3367 2629 3368
rect 2623 3366 2629 3367
rect 2667 3367 2668 3368
rect 2672 3367 2673 3371
rect 2667 3366 2673 3367
rect 2795 3371 2804 3372
rect 2795 3367 2796 3371
rect 2803 3367 2804 3371
rect 2795 3366 2804 3367
rect 2842 3371 2848 3372
rect 2842 3367 2843 3371
rect 2847 3370 2848 3371
rect 2923 3371 2929 3372
rect 2923 3370 2924 3371
rect 2847 3368 2924 3370
rect 2847 3367 2848 3368
rect 2842 3366 2848 3367
rect 2923 3367 2924 3368
rect 2928 3367 2929 3371
rect 2923 3366 2929 3367
rect 3015 3371 3021 3372
rect 3015 3367 3016 3371
rect 3020 3370 3021 3371
rect 3059 3371 3065 3372
rect 3059 3370 3060 3371
rect 3020 3368 3060 3370
rect 3020 3367 3021 3368
rect 3015 3366 3021 3367
rect 3059 3367 3060 3368
rect 3064 3367 3065 3371
rect 3059 3366 3065 3367
rect 223 3364 282 3366
rect 223 3363 224 3364
rect 218 3362 224 3363
rect 678 3363 684 3364
rect 678 3362 679 3363
rect 236 3360 679 3362
rect 236 3358 238 3360
rect 678 3359 679 3360
rect 683 3359 684 3363
rect 678 3358 684 3359
rect 235 3357 241 3358
rect 235 3353 236 3357
rect 240 3353 241 3357
rect 235 3352 241 3353
rect 327 3355 333 3356
rect 327 3351 328 3355
rect 332 3354 333 3355
rect 395 3355 401 3356
rect 395 3354 396 3355
rect 332 3352 396 3354
rect 332 3351 333 3352
rect 327 3350 333 3351
rect 395 3351 396 3352
rect 400 3351 401 3355
rect 395 3350 401 3351
rect 471 3355 477 3356
rect 471 3351 472 3355
rect 476 3354 477 3355
rect 563 3355 569 3356
rect 563 3354 564 3355
rect 476 3352 564 3354
rect 476 3351 477 3352
rect 471 3350 477 3351
rect 563 3351 564 3352
rect 568 3351 569 3355
rect 563 3350 569 3351
rect 631 3355 637 3356
rect 631 3351 632 3355
rect 636 3354 637 3355
rect 723 3355 729 3356
rect 723 3354 724 3355
rect 636 3352 724 3354
rect 636 3351 637 3352
rect 631 3350 637 3351
rect 723 3351 724 3352
rect 728 3351 729 3355
rect 723 3350 729 3351
rect 883 3355 889 3356
rect 883 3351 884 3355
rect 888 3354 889 3355
rect 950 3355 956 3356
rect 950 3354 951 3355
rect 888 3352 951 3354
rect 888 3351 889 3352
rect 883 3350 889 3351
rect 950 3351 951 3352
rect 955 3351 956 3355
rect 950 3350 956 3351
rect 959 3355 965 3356
rect 959 3351 960 3355
rect 964 3354 965 3355
rect 1027 3355 1033 3356
rect 1027 3354 1028 3355
rect 964 3352 1028 3354
rect 964 3351 965 3352
rect 959 3350 965 3351
rect 1027 3351 1028 3352
rect 1032 3351 1033 3355
rect 1027 3350 1033 3351
rect 1063 3355 1069 3356
rect 1063 3351 1064 3355
rect 1068 3354 1069 3355
rect 1171 3355 1177 3356
rect 1171 3354 1172 3355
rect 1068 3352 1172 3354
rect 1068 3351 1069 3352
rect 1063 3350 1069 3351
rect 1171 3351 1172 3352
rect 1176 3351 1177 3355
rect 1171 3350 1177 3351
rect 1307 3355 1313 3356
rect 1307 3351 1308 3355
rect 1312 3354 1313 3355
rect 1351 3355 1357 3356
rect 1351 3354 1352 3355
rect 1312 3352 1352 3354
rect 1312 3351 1313 3352
rect 1307 3350 1313 3351
rect 1351 3351 1352 3352
rect 1356 3351 1357 3355
rect 1351 3350 1357 3351
rect 1443 3355 1449 3356
rect 1443 3351 1444 3355
rect 1448 3354 1449 3355
rect 1503 3355 1509 3356
rect 1503 3354 1504 3355
rect 1448 3352 1504 3354
rect 1448 3351 1449 3352
rect 1443 3350 1449 3351
rect 1503 3351 1504 3352
rect 1508 3351 1509 3355
rect 1503 3350 1509 3351
rect 1586 3355 1593 3356
rect 1586 3351 1587 3355
rect 1592 3351 1593 3355
rect 1586 3350 1593 3351
rect 1923 3355 1929 3356
rect 1923 3351 1924 3355
rect 1928 3354 1929 3355
rect 1990 3355 1996 3356
rect 1990 3354 1991 3355
rect 1928 3352 1991 3354
rect 1928 3351 1929 3352
rect 1923 3350 1929 3351
rect 1990 3351 1991 3352
rect 1995 3351 1996 3355
rect 1990 3350 1996 3351
rect 2070 3355 2081 3356
rect 2070 3351 2071 3355
rect 2075 3351 2076 3355
rect 2080 3351 2081 3355
rect 2070 3350 2081 3351
rect 2214 3355 2220 3356
rect 2214 3351 2215 3355
rect 2219 3354 2220 3355
rect 2235 3355 2241 3356
rect 2235 3354 2236 3355
rect 2219 3352 2236 3354
rect 2219 3351 2220 3352
rect 2214 3350 2220 3351
rect 2235 3351 2236 3352
rect 2240 3351 2241 3355
rect 2235 3350 2241 3351
rect 2335 3355 2341 3356
rect 2335 3351 2336 3355
rect 2340 3354 2341 3355
rect 2395 3355 2401 3356
rect 2395 3354 2396 3355
rect 2340 3352 2396 3354
rect 2340 3351 2341 3352
rect 2335 3350 2341 3351
rect 2395 3351 2396 3352
rect 2400 3351 2401 3355
rect 2395 3350 2401 3351
rect 2471 3355 2477 3356
rect 2471 3351 2472 3355
rect 2476 3354 2477 3355
rect 2563 3355 2569 3356
rect 2563 3354 2564 3355
rect 2476 3352 2564 3354
rect 2476 3351 2477 3352
rect 2471 3350 2477 3351
rect 2563 3351 2564 3352
rect 2568 3351 2569 3355
rect 2563 3350 2569 3351
rect 2710 3355 2716 3356
rect 2710 3351 2711 3355
rect 2715 3354 2716 3355
rect 2731 3355 2737 3356
rect 2731 3354 2732 3355
rect 2715 3352 2732 3354
rect 2715 3351 2716 3352
rect 2710 3350 2716 3351
rect 2731 3351 2732 3352
rect 2736 3351 2737 3355
rect 2731 3350 2737 3351
rect 2907 3355 2913 3356
rect 2907 3351 2908 3355
rect 2912 3354 2913 3355
rect 2986 3355 2992 3356
rect 2986 3354 2987 3355
rect 2912 3352 2987 3354
rect 2912 3351 2913 3352
rect 2907 3350 2913 3351
rect 2986 3351 2987 3352
rect 2991 3351 2992 3355
rect 2986 3350 2992 3351
rect 3083 3355 3092 3356
rect 3083 3351 3084 3355
rect 3091 3351 3092 3355
rect 3083 3350 3092 3351
rect 206 3345 212 3346
rect 206 3341 207 3345
rect 211 3341 212 3345
rect 206 3340 212 3341
rect 366 3345 372 3346
rect 366 3341 367 3345
rect 371 3341 372 3345
rect 366 3340 372 3341
rect 534 3345 540 3346
rect 534 3341 535 3345
rect 539 3341 540 3345
rect 534 3340 540 3341
rect 694 3345 700 3346
rect 694 3341 695 3345
rect 699 3341 700 3345
rect 694 3340 700 3341
rect 854 3345 860 3346
rect 854 3341 855 3345
rect 859 3341 860 3345
rect 854 3340 860 3341
rect 998 3345 1004 3346
rect 998 3341 999 3345
rect 1003 3341 1004 3345
rect 998 3340 1004 3341
rect 1142 3345 1148 3346
rect 1142 3341 1143 3345
rect 1147 3341 1148 3345
rect 1142 3340 1148 3341
rect 1278 3345 1284 3346
rect 1278 3341 1279 3345
rect 1283 3341 1284 3345
rect 1278 3340 1284 3341
rect 1414 3345 1420 3346
rect 1414 3341 1415 3345
rect 1419 3341 1420 3345
rect 1414 3340 1420 3341
rect 1558 3345 1564 3346
rect 1558 3341 1559 3345
rect 1563 3341 1564 3345
rect 1558 3340 1564 3341
rect 1894 3345 1900 3346
rect 1894 3341 1895 3345
rect 1899 3341 1900 3345
rect 1894 3340 1900 3341
rect 2046 3345 2052 3346
rect 2046 3341 2047 3345
rect 2051 3341 2052 3345
rect 2046 3340 2052 3341
rect 2206 3345 2212 3346
rect 2206 3341 2207 3345
rect 2211 3341 2212 3345
rect 2206 3340 2212 3341
rect 2366 3345 2372 3346
rect 2366 3341 2367 3345
rect 2371 3341 2372 3345
rect 2366 3340 2372 3341
rect 2534 3345 2540 3346
rect 2534 3341 2535 3345
rect 2539 3341 2540 3345
rect 2534 3340 2540 3341
rect 2702 3345 2708 3346
rect 2702 3341 2703 3345
rect 2707 3341 2708 3345
rect 2702 3340 2708 3341
rect 2878 3345 2884 3346
rect 2878 3341 2879 3345
rect 2883 3341 2884 3345
rect 2878 3340 2884 3341
rect 3054 3345 3060 3346
rect 3054 3341 3055 3345
rect 3059 3341 3060 3345
rect 3054 3340 3060 3341
rect 1950 3339 1956 3340
rect 1950 3338 1951 3339
rect 1948 3335 1951 3338
rect 1955 3335 1956 3339
rect 1948 3334 1956 3335
rect 110 3332 116 3333
rect 1822 3332 1828 3333
rect 110 3328 111 3332
rect 115 3328 116 3332
rect 327 3331 333 3332
rect 327 3330 328 3331
rect 261 3328 328 3330
rect 110 3327 116 3328
rect 327 3327 328 3328
rect 332 3327 333 3331
rect 471 3331 477 3332
rect 471 3330 472 3331
rect 421 3328 472 3330
rect 327 3326 333 3327
rect 471 3327 472 3328
rect 476 3327 477 3331
rect 631 3331 637 3332
rect 631 3330 632 3331
rect 589 3328 632 3330
rect 471 3326 477 3327
rect 631 3327 632 3328
rect 636 3327 637 3331
rect 959 3331 965 3332
rect 959 3330 960 3331
rect 909 3328 960 3330
rect 631 3326 637 3327
rect 959 3327 960 3328
rect 964 3327 965 3331
rect 1063 3331 1069 3332
rect 1063 3330 1064 3331
rect 1053 3328 1064 3330
rect 959 3326 965 3327
rect 1063 3327 1064 3328
rect 1068 3327 1069 3331
rect 1822 3328 1823 3332
rect 1827 3328 1828 3332
rect 1063 3326 1069 3327
rect 1134 3327 1140 3328
rect 1134 3323 1135 3327
rect 1139 3326 1140 3327
rect 1351 3327 1357 3328
rect 1139 3324 1161 3326
rect 1139 3323 1140 3324
rect 1134 3322 1140 3323
rect 1351 3323 1352 3327
rect 1356 3326 1357 3327
rect 1503 3327 1509 3328
rect 1822 3327 1828 3328
rect 1862 3332 1868 3333
rect 1862 3328 1863 3332
rect 1867 3328 1868 3332
rect 1948 3329 1950 3334
rect 3574 3332 3580 3333
rect 2335 3331 2341 3332
rect 2335 3330 2336 3331
rect 2261 3328 2336 3330
rect 1862 3327 1868 3328
rect 1990 3327 1996 3328
rect 1356 3324 1433 3326
rect 1356 3323 1357 3324
rect 1351 3322 1357 3323
rect 1503 3323 1504 3327
rect 1508 3326 1509 3327
rect 1508 3324 1577 3326
rect 1508 3323 1509 3324
rect 1503 3322 1509 3323
rect 1990 3323 1991 3327
rect 1995 3326 1996 3327
rect 2335 3327 2336 3328
rect 2340 3327 2341 3331
rect 2471 3331 2477 3332
rect 2471 3330 2472 3331
rect 2421 3328 2472 3330
rect 2335 3326 2341 3327
rect 2471 3327 2472 3328
rect 2476 3327 2477 3331
rect 3574 3328 3575 3332
rect 3579 3328 3580 3332
rect 2471 3326 2477 3327
rect 2602 3327 2608 3328
rect 1995 3324 2065 3326
rect 1995 3323 1996 3324
rect 1990 3322 1996 3323
rect 2602 3323 2603 3327
rect 2607 3326 2608 3327
rect 2986 3327 2992 3328
rect 3574 3327 3580 3328
rect 2607 3324 2721 3326
rect 2607 3323 2608 3324
rect 2602 3322 2608 3323
rect 2986 3323 2987 3327
rect 2991 3326 2992 3327
rect 2991 3324 3073 3326
rect 2991 3323 2992 3324
rect 2986 3322 2992 3323
rect 110 3315 116 3316
rect 110 3311 111 3315
rect 115 3311 116 3315
rect 110 3310 116 3311
rect 618 3315 624 3316
rect 618 3311 619 3315
rect 623 3314 624 3315
rect 1378 3315 1384 3316
rect 1378 3314 1379 3315
rect 623 3312 705 3314
rect 1329 3312 1379 3314
rect 623 3311 624 3312
rect 618 3310 624 3311
rect 1378 3311 1379 3312
rect 1383 3311 1384 3315
rect 1378 3310 1384 3311
rect 1822 3315 1828 3316
rect 1822 3311 1823 3315
rect 1827 3311 1828 3315
rect 1822 3310 1828 3311
rect 1862 3315 1868 3316
rect 1862 3311 1863 3315
rect 1867 3311 1868 3315
rect 1862 3310 1868 3311
rect 2494 3315 2500 3316
rect 2494 3311 2495 3315
rect 2499 3314 2500 3315
rect 2854 3315 2860 3316
rect 2499 3312 2545 3314
rect 2499 3311 2500 3312
rect 2494 3310 2500 3311
rect 2854 3311 2855 3315
rect 2859 3314 2860 3315
rect 3574 3315 3580 3316
rect 2859 3312 2889 3314
rect 2859 3311 2860 3312
rect 2854 3310 2860 3311
rect 3574 3311 3575 3315
rect 3579 3311 3580 3315
rect 3574 3310 3580 3311
rect 198 3305 204 3306
rect 198 3301 199 3305
rect 203 3301 204 3305
rect 198 3300 204 3301
rect 358 3305 364 3306
rect 358 3301 359 3305
rect 363 3301 364 3305
rect 358 3300 364 3301
rect 526 3305 532 3306
rect 526 3301 527 3305
rect 531 3301 532 3305
rect 526 3300 532 3301
rect 686 3305 692 3306
rect 686 3301 687 3305
rect 691 3301 692 3305
rect 686 3300 692 3301
rect 846 3305 852 3306
rect 846 3301 847 3305
rect 851 3301 852 3305
rect 846 3300 852 3301
rect 990 3305 996 3306
rect 990 3301 991 3305
rect 995 3301 996 3305
rect 990 3300 996 3301
rect 1134 3305 1140 3306
rect 1134 3301 1135 3305
rect 1139 3301 1140 3305
rect 1134 3300 1140 3301
rect 1270 3305 1276 3306
rect 1270 3301 1271 3305
rect 1275 3301 1276 3305
rect 1270 3300 1276 3301
rect 1406 3305 1412 3306
rect 1406 3301 1407 3305
rect 1411 3301 1412 3305
rect 1406 3300 1412 3301
rect 1550 3305 1556 3306
rect 1550 3301 1551 3305
rect 1555 3301 1556 3305
rect 1550 3300 1556 3301
rect 1886 3305 1892 3306
rect 1886 3301 1887 3305
rect 1891 3301 1892 3305
rect 1886 3300 1892 3301
rect 2038 3305 2044 3306
rect 2038 3301 2039 3305
rect 2043 3301 2044 3305
rect 2038 3300 2044 3301
rect 2198 3305 2204 3306
rect 2198 3301 2199 3305
rect 2203 3301 2204 3305
rect 2198 3300 2204 3301
rect 2358 3305 2364 3306
rect 2358 3301 2359 3305
rect 2363 3301 2364 3305
rect 2358 3300 2364 3301
rect 2526 3305 2532 3306
rect 2526 3301 2527 3305
rect 2531 3301 2532 3305
rect 2526 3300 2532 3301
rect 2694 3305 2700 3306
rect 2694 3301 2695 3305
rect 2699 3301 2700 3305
rect 2694 3300 2700 3301
rect 2870 3305 2876 3306
rect 2870 3301 2871 3305
rect 2875 3301 2876 3305
rect 2870 3300 2876 3301
rect 3046 3305 3052 3306
rect 3046 3301 3047 3305
rect 3051 3301 3052 3305
rect 3046 3300 3052 3301
rect 254 3279 260 3280
rect 254 3275 255 3279
rect 259 3275 260 3279
rect 254 3274 260 3275
rect 374 3279 380 3280
rect 374 3275 375 3279
rect 379 3275 380 3279
rect 374 3274 380 3275
rect 510 3279 516 3280
rect 510 3275 511 3279
rect 515 3275 516 3279
rect 510 3274 516 3275
rect 662 3279 668 3280
rect 662 3275 663 3279
rect 667 3275 668 3279
rect 662 3274 668 3275
rect 822 3279 828 3280
rect 822 3275 823 3279
rect 827 3275 828 3279
rect 822 3274 828 3275
rect 990 3279 996 3280
rect 990 3275 991 3279
rect 995 3275 996 3279
rect 990 3274 996 3275
rect 1166 3279 1172 3280
rect 1166 3275 1167 3279
rect 1171 3275 1172 3279
rect 1166 3274 1172 3275
rect 1342 3279 1348 3280
rect 1342 3275 1343 3279
rect 1347 3275 1348 3279
rect 1342 3274 1348 3275
rect 1518 3279 1524 3280
rect 1518 3275 1519 3279
rect 1523 3275 1524 3279
rect 1518 3274 1524 3275
rect 1886 3279 1892 3280
rect 1886 3275 1887 3279
rect 1891 3275 1892 3279
rect 1886 3274 1892 3275
rect 2062 3279 2068 3280
rect 2062 3275 2063 3279
rect 2067 3275 2068 3279
rect 2062 3274 2068 3275
rect 2262 3279 2268 3280
rect 2262 3275 2263 3279
rect 2267 3275 2268 3279
rect 2262 3274 2268 3275
rect 2454 3279 2460 3280
rect 2454 3275 2455 3279
rect 2459 3275 2460 3279
rect 2454 3274 2460 3275
rect 2638 3279 2644 3280
rect 2638 3275 2639 3279
rect 2643 3275 2644 3279
rect 2638 3274 2644 3275
rect 2814 3279 2820 3280
rect 2814 3275 2815 3279
rect 2819 3275 2820 3279
rect 2814 3274 2820 3275
rect 2982 3279 2988 3280
rect 2982 3275 2983 3279
rect 2987 3275 2988 3279
rect 2982 3274 2988 3275
rect 3150 3279 3156 3280
rect 3150 3275 3151 3279
rect 3155 3275 3156 3279
rect 3150 3274 3156 3275
rect 3318 3279 3324 3280
rect 3318 3275 3319 3279
rect 3323 3275 3324 3279
rect 3318 3274 3324 3275
rect 3478 3279 3484 3280
rect 3478 3275 3479 3279
rect 3483 3275 3484 3279
rect 3478 3274 3484 3275
rect 738 3271 744 3272
rect 110 3269 116 3270
rect 110 3265 111 3269
rect 115 3265 116 3269
rect 738 3267 739 3271
rect 743 3270 744 3271
rect 950 3271 956 3272
rect 743 3268 841 3270
rect 743 3267 744 3268
rect 738 3266 744 3267
rect 950 3267 951 3271
rect 955 3270 956 3271
rect 2710 3271 2716 3272
rect 2710 3270 2711 3271
rect 955 3268 1009 3270
rect 1822 3269 1828 3270
rect 955 3267 956 3268
rect 950 3266 956 3267
rect 110 3264 116 3265
rect 1822 3265 1823 3269
rect 1827 3265 1828 3269
rect 1822 3264 1828 3265
rect 1862 3269 1868 3270
rect 1862 3265 1863 3269
rect 1867 3265 1868 3269
rect 2072 3268 2081 3270
rect 2697 3268 2711 3270
rect 1862 3264 1868 3265
rect 2070 3267 2076 3268
rect 2070 3263 2071 3267
rect 2075 3263 2076 3267
rect 2710 3267 2711 3268
rect 2715 3267 2716 3271
rect 2710 3266 2716 3267
rect 3574 3269 3580 3270
rect 3574 3265 3575 3269
rect 3579 3265 3580 3269
rect 3574 3264 3580 3265
rect 2070 3262 2076 3263
rect 367 3255 373 3256
rect 367 3254 368 3255
rect 110 3252 116 3253
rect 317 3252 368 3254
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 367 3251 368 3252
rect 372 3251 373 3255
rect 503 3255 509 3256
rect 503 3254 504 3255
rect 437 3252 504 3254
rect 367 3250 373 3251
rect 503 3251 504 3252
rect 508 3251 509 3255
rect 655 3255 661 3256
rect 655 3254 656 3255
rect 573 3252 656 3254
rect 503 3250 509 3251
rect 655 3251 656 3252
rect 660 3251 661 3255
rect 815 3255 821 3256
rect 815 3254 816 3255
rect 725 3252 816 3254
rect 655 3250 661 3251
rect 815 3251 816 3252
rect 820 3251 821 3255
rect 815 3250 821 3251
rect 1058 3255 1064 3256
rect 1058 3251 1059 3255
rect 1063 3254 1064 3255
rect 1511 3255 1517 3256
rect 1511 3254 1512 3255
rect 1063 3252 1193 3254
rect 1405 3252 1512 3254
rect 1063 3251 1064 3252
rect 1058 3250 1064 3251
rect 1511 3251 1512 3252
rect 1516 3251 1517 3255
rect 1586 3255 1592 3256
rect 1586 3254 1587 3255
rect 1581 3252 1587 3254
rect 1511 3250 1517 3251
rect 1586 3251 1587 3252
rect 1591 3251 1592 3255
rect 2055 3255 2061 3256
rect 2055 3254 2056 3255
rect 1586 3250 1592 3251
rect 1822 3252 1828 3253
rect 110 3247 116 3248
rect 1822 3248 1823 3252
rect 1827 3248 1828 3252
rect 1822 3247 1828 3248
rect 1862 3252 1868 3253
rect 1949 3252 2056 3254
rect 1862 3248 1863 3252
rect 1867 3248 1868 3252
rect 2055 3251 2056 3252
rect 2060 3251 2061 3255
rect 2330 3255 2336 3256
rect 2330 3254 2331 3255
rect 2325 3252 2331 3254
rect 2055 3250 2061 3251
rect 2330 3251 2331 3252
rect 2335 3251 2336 3255
rect 2330 3250 2336 3251
rect 2338 3255 2344 3256
rect 2338 3251 2339 3255
rect 2343 3254 2344 3255
rect 2975 3255 2981 3256
rect 2975 3254 2976 3255
rect 2343 3252 2481 3254
rect 2877 3252 2976 3254
rect 2343 3251 2344 3252
rect 2338 3250 2344 3251
rect 2975 3251 2976 3252
rect 2980 3251 2981 3255
rect 3062 3255 3068 3256
rect 3062 3254 3063 3255
rect 3045 3252 3063 3254
rect 2975 3250 2981 3251
rect 3062 3251 3063 3252
rect 3067 3251 3068 3255
rect 3062 3250 3068 3251
rect 3070 3255 3076 3256
rect 3070 3251 3071 3255
rect 3075 3254 3076 3255
rect 3471 3255 3477 3256
rect 3471 3254 3472 3255
rect 3075 3252 3177 3254
rect 3381 3252 3472 3254
rect 3075 3251 3076 3252
rect 3070 3250 3076 3251
rect 3471 3251 3472 3252
rect 3476 3251 3477 3255
rect 3546 3255 3552 3256
rect 3546 3254 3547 3255
rect 3541 3252 3547 3254
rect 3471 3250 3477 3251
rect 3546 3251 3547 3252
rect 3551 3251 3552 3255
rect 3546 3250 3552 3251
rect 3574 3252 3580 3253
rect 1862 3247 1868 3248
rect 3574 3248 3575 3252
rect 3579 3248 3580 3252
rect 3574 3247 3580 3248
rect 262 3239 268 3240
rect 262 3235 263 3239
rect 267 3235 268 3239
rect 262 3234 268 3235
rect 382 3239 388 3240
rect 382 3235 383 3239
rect 387 3235 388 3239
rect 382 3234 388 3235
rect 518 3239 524 3240
rect 518 3235 519 3239
rect 523 3235 524 3239
rect 518 3234 524 3235
rect 670 3239 676 3240
rect 670 3235 671 3239
rect 675 3235 676 3239
rect 670 3234 676 3235
rect 830 3239 836 3240
rect 830 3235 831 3239
rect 835 3235 836 3239
rect 830 3234 836 3235
rect 998 3239 1004 3240
rect 998 3235 999 3239
rect 1003 3235 1004 3239
rect 998 3234 1004 3235
rect 1174 3239 1180 3240
rect 1174 3235 1175 3239
rect 1179 3235 1180 3239
rect 1174 3234 1180 3235
rect 1350 3239 1356 3240
rect 1350 3235 1351 3239
rect 1355 3235 1356 3239
rect 1350 3234 1356 3235
rect 1526 3239 1532 3240
rect 1526 3235 1527 3239
rect 1531 3235 1532 3239
rect 1526 3234 1532 3235
rect 1894 3239 1900 3240
rect 1894 3235 1895 3239
rect 1899 3235 1900 3239
rect 1894 3234 1900 3235
rect 2070 3239 2076 3240
rect 2070 3235 2071 3239
rect 2075 3235 2076 3239
rect 2070 3234 2076 3235
rect 2270 3239 2276 3240
rect 2270 3235 2271 3239
rect 2275 3235 2276 3239
rect 2270 3234 2276 3235
rect 2462 3239 2468 3240
rect 2462 3235 2463 3239
rect 2467 3235 2468 3239
rect 2462 3234 2468 3235
rect 2646 3239 2652 3240
rect 2646 3235 2647 3239
rect 2651 3235 2652 3239
rect 2646 3234 2652 3235
rect 2822 3239 2828 3240
rect 2822 3235 2823 3239
rect 2827 3235 2828 3239
rect 2822 3234 2828 3235
rect 2990 3239 2996 3240
rect 2990 3235 2991 3239
rect 2995 3235 2996 3239
rect 2990 3234 2996 3235
rect 3158 3239 3164 3240
rect 3158 3235 3159 3239
rect 3163 3235 3164 3239
rect 3158 3234 3164 3235
rect 3326 3239 3332 3240
rect 3326 3235 3327 3239
rect 3331 3235 3332 3239
rect 3326 3234 3332 3235
rect 3486 3239 3492 3240
rect 3486 3235 3487 3239
rect 3491 3235 3492 3239
rect 3486 3234 3492 3235
rect 291 3227 300 3228
rect 291 3223 292 3227
rect 299 3223 300 3227
rect 291 3222 300 3223
rect 367 3227 373 3228
rect 367 3223 368 3227
rect 372 3226 373 3227
rect 411 3227 417 3228
rect 411 3226 412 3227
rect 372 3224 412 3226
rect 372 3223 373 3224
rect 367 3222 373 3223
rect 411 3223 412 3224
rect 416 3223 417 3227
rect 411 3222 417 3223
rect 503 3227 509 3228
rect 503 3223 504 3227
rect 508 3226 509 3227
rect 547 3227 553 3228
rect 547 3226 548 3227
rect 508 3224 548 3226
rect 508 3223 509 3224
rect 503 3222 509 3223
rect 547 3223 548 3224
rect 552 3223 553 3227
rect 547 3222 553 3223
rect 655 3227 661 3228
rect 655 3223 656 3227
rect 660 3226 661 3227
rect 699 3227 705 3228
rect 699 3226 700 3227
rect 660 3224 700 3226
rect 660 3223 661 3224
rect 655 3222 661 3223
rect 699 3223 700 3224
rect 704 3223 705 3227
rect 699 3222 705 3223
rect 815 3227 821 3228
rect 815 3223 816 3227
rect 820 3226 821 3227
rect 859 3227 865 3228
rect 859 3226 860 3227
rect 820 3224 860 3226
rect 820 3223 821 3224
rect 815 3222 821 3223
rect 859 3223 860 3224
rect 864 3223 865 3227
rect 859 3222 865 3223
rect 1027 3227 1033 3228
rect 1027 3223 1028 3227
rect 1032 3226 1033 3227
rect 1058 3227 1064 3228
rect 1058 3226 1059 3227
rect 1032 3224 1059 3226
rect 1032 3223 1033 3224
rect 1027 3222 1033 3223
rect 1058 3223 1059 3224
rect 1063 3223 1064 3227
rect 1058 3222 1064 3223
rect 1203 3227 1212 3228
rect 1203 3223 1204 3227
rect 1211 3223 1212 3227
rect 1203 3222 1212 3223
rect 1378 3227 1385 3228
rect 1378 3223 1379 3227
rect 1384 3223 1385 3227
rect 1378 3222 1385 3223
rect 1511 3227 1517 3228
rect 1511 3223 1512 3227
rect 1516 3226 1517 3227
rect 1555 3227 1561 3228
rect 1555 3226 1556 3227
rect 1516 3224 1556 3226
rect 1516 3223 1517 3224
rect 1511 3222 1517 3223
rect 1555 3223 1556 3224
rect 1560 3223 1561 3227
rect 1555 3222 1561 3223
rect 1923 3227 1929 3228
rect 1923 3223 1924 3227
rect 1928 3226 1929 3227
rect 1954 3227 1960 3228
rect 1954 3226 1955 3227
rect 1928 3224 1955 3226
rect 1928 3223 1929 3224
rect 1923 3222 1929 3223
rect 1954 3223 1955 3224
rect 1959 3223 1960 3227
rect 1954 3222 1960 3223
rect 2055 3227 2061 3228
rect 2055 3223 2056 3227
rect 2060 3226 2061 3227
rect 2099 3227 2105 3228
rect 2099 3226 2100 3227
rect 2060 3224 2100 3226
rect 2060 3223 2061 3224
rect 2055 3222 2061 3223
rect 2099 3223 2100 3224
rect 2104 3223 2105 3227
rect 2099 3222 2105 3223
rect 2299 3227 2305 3228
rect 2299 3223 2300 3227
rect 2304 3226 2305 3227
rect 2338 3227 2344 3228
rect 2338 3226 2339 3227
rect 2304 3224 2339 3226
rect 2304 3223 2305 3224
rect 2299 3222 2305 3223
rect 2338 3223 2339 3224
rect 2343 3223 2344 3227
rect 2338 3222 2344 3223
rect 2491 3227 2500 3228
rect 2491 3223 2492 3227
rect 2499 3223 2500 3227
rect 2491 3222 2500 3223
rect 2675 3227 2684 3228
rect 2675 3223 2676 3227
rect 2683 3223 2684 3227
rect 2675 3222 2684 3223
rect 2851 3227 2860 3228
rect 2851 3223 2852 3227
rect 2859 3223 2860 3227
rect 2851 3222 2860 3223
rect 2975 3227 2981 3228
rect 2975 3223 2976 3227
rect 2980 3226 2981 3227
rect 3019 3227 3025 3228
rect 3019 3226 3020 3227
rect 2980 3224 3020 3226
rect 2980 3223 2981 3224
rect 2975 3222 2981 3223
rect 3019 3223 3020 3224
rect 3024 3223 3025 3227
rect 3019 3222 3025 3223
rect 3062 3227 3068 3228
rect 3062 3223 3063 3227
rect 3067 3226 3068 3227
rect 3187 3227 3193 3228
rect 3187 3226 3188 3227
rect 3067 3224 3188 3226
rect 3067 3223 3068 3224
rect 3062 3222 3068 3223
rect 3187 3223 3188 3224
rect 3192 3223 3193 3227
rect 3187 3222 3193 3223
rect 3279 3227 3285 3228
rect 3279 3223 3280 3227
rect 3284 3226 3285 3227
rect 3355 3227 3361 3228
rect 3355 3226 3356 3227
rect 3284 3224 3356 3226
rect 3284 3223 3285 3224
rect 3279 3222 3285 3223
rect 3355 3223 3356 3224
rect 3360 3223 3361 3227
rect 3355 3222 3361 3223
rect 3471 3227 3477 3228
rect 3471 3223 3472 3227
rect 3476 3226 3477 3227
rect 3515 3227 3521 3228
rect 3515 3226 3516 3227
rect 3476 3224 3516 3226
rect 3476 3223 3477 3224
rect 3471 3222 3477 3223
rect 3515 3223 3516 3224
rect 3520 3223 3521 3227
rect 3515 3222 3521 3223
rect 1923 3215 1929 3216
rect 459 3211 468 3212
rect 459 3207 460 3211
rect 467 3207 468 3211
rect 459 3206 468 3207
rect 511 3211 517 3212
rect 511 3207 512 3211
rect 516 3210 517 3211
rect 579 3211 585 3212
rect 579 3210 580 3211
rect 516 3208 580 3210
rect 516 3207 517 3208
rect 511 3206 517 3207
rect 579 3207 580 3208
rect 584 3207 585 3211
rect 579 3206 585 3207
rect 631 3211 637 3212
rect 631 3207 632 3211
rect 636 3210 637 3211
rect 699 3211 705 3212
rect 699 3210 700 3211
rect 636 3208 700 3210
rect 636 3207 637 3208
rect 631 3206 637 3207
rect 699 3207 700 3208
rect 704 3207 705 3211
rect 699 3206 705 3207
rect 751 3211 757 3212
rect 751 3207 752 3211
rect 756 3210 757 3211
rect 827 3211 833 3212
rect 827 3210 828 3211
rect 756 3208 828 3210
rect 756 3207 757 3208
rect 751 3206 757 3207
rect 827 3207 828 3208
rect 832 3207 833 3211
rect 827 3206 833 3207
rect 963 3211 969 3212
rect 963 3207 964 3211
rect 968 3210 969 3211
rect 1023 3211 1029 3212
rect 968 3208 1018 3210
rect 968 3207 969 3208
rect 963 3206 969 3207
rect 1016 3202 1018 3208
rect 1023 3207 1024 3211
rect 1028 3210 1029 3211
rect 1107 3211 1113 3212
rect 1107 3210 1108 3211
rect 1028 3208 1108 3210
rect 1028 3207 1029 3208
rect 1023 3206 1029 3207
rect 1107 3207 1108 3208
rect 1112 3207 1113 3211
rect 1107 3206 1113 3207
rect 1191 3211 1197 3212
rect 1191 3207 1192 3211
rect 1196 3210 1197 3211
rect 1259 3211 1265 3212
rect 1259 3210 1260 3211
rect 1196 3208 1260 3210
rect 1196 3207 1197 3208
rect 1191 3206 1197 3207
rect 1259 3207 1260 3208
rect 1264 3207 1265 3211
rect 1259 3206 1265 3207
rect 1411 3211 1417 3212
rect 1411 3207 1412 3211
rect 1416 3210 1417 3211
rect 1479 3211 1485 3212
rect 1479 3210 1480 3211
rect 1416 3208 1480 3210
rect 1416 3207 1417 3208
rect 1411 3206 1417 3207
rect 1479 3207 1480 3208
rect 1484 3207 1485 3211
rect 1479 3206 1485 3207
rect 1563 3211 1569 3212
rect 1563 3207 1564 3211
rect 1568 3210 1569 3211
rect 1586 3211 1592 3212
rect 1586 3210 1587 3211
rect 1568 3208 1587 3210
rect 1568 3207 1569 3208
rect 1563 3206 1569 3207
rect 1586 3207 1587 3208
rect 1591 3207 1592 3211
rect 1923 3211 1924 3215
rect 1928 3214 1929 3215
rect 1962 3215 1968 3216
rect 1962 3214 1963 3215
rect 1928 3212 1963 3214
rect 1928 3211 1929 3212
rect 1923 3210 1929 3211
rect 1962 3211 1963 3212
rect 1967 3211 1968 3215
rect 1962 3210 1968 3211
rect 2115 3215 2121 3216
rect 2115 3211 2116 3215
rect 2120 3214 2121 3215
rect 2146 3215 2152 3216
rect 2146 3214 2147 3215
rect 2120 3212 2147 3214
rect 2120 3211 2121 3212
rect 2115 3210 2121 3211
rect 2146 3211 2147 3212
rect 2151 3211 2152 3215
rect 2146 3210 2152 3211
rect 2330 3215 2337 3216
rect 2330 3211 2331 3215
rect 2336 3211 2337 3215
rect 2330 3210 2337 3211
rect 2423 3215 2429 3216
rect 2423 3211 2424 3215
rect 2428 3214 2429 3215
rect 2539 3215 2545 3216
rect 2539 3214 2540 3215
rect 2428 3212 2540 3214
rect 2428 3211 2429 3212
rect 2423 3210 2429 3211
rect 2539 3211 2540 3212
rect 2544 3211 2545 3215
rect 2539 3210 2545 3211
rect 2731 3215 2737 3216
rect 2731 3211 2732 3215
rect 2736 3214 2737 3215
rect 2762 3215 2768 3216
rect 2762 3214 2763 3215
rect 2736 3212 2763 3214
rect 2736 3211 2737 3212
rect 2731 3210 2737 3211
rect 2762 3211 2763 3212
rect 2767 3211 2768 3215
rect 2762 3210 2768 3211
rect 2907 3215 2913 3216
rect 2907 3211 2908 3215
rect 2912 3214 2913 3215
rect 2978 3215 2984 3216
rect 2978 3214 2979 3215
rect 2912 3212 2979 3214
rect 2912 3211 2913 3212
rect 2907 3210 2913 3211
rect 2978 3211 2979 3212
rect 2983 3211 2984 3215
rect 2978 3210 2984 3211
rect 3067 3215 3076 3216
rect 3067 3211 3068 3215
rect 3075 3211 3076 3215
rect 3067 3210 3076 3211
rect 3227 3215 3233 3216
rect 3227 3211 3228 3215
rect 3232 3214 3233 3215
rect 3295 3215 3301 3216
rect 3295 3214 3296 3215
rect 3232 3212 3296 3214
rect 3232 3211 3233 3212
rect 3227 3210 3233 3211
rect 3295 3211 3296 3212
rect 3300 3211 3301 3215
rect 3295 3210 3301 3211
rect 3379 3215 3385 3216
rect 3379 3211 3380 3215
rect 3384 3214 3385 3215
rect 3410 3215 3416 3216
rect 3410 3214 3411 3215
rect 3384 3212 3411 3214
rect 3384 3211 3385 3212
rect 3379 3210 3385 3211
rect 3410 3211 3411 3212
rect 3415 3211 3416 3215
rect 3410 3210 3416 3211
rect 3515 3215 3521 3216
rect 3515 3211 3516 3215
rect 3520 3214 3521 3215
rect 3546 3215 3552 3216
rect 3546 3214 3547 3215
rect 3520 3212 3547 3214
rect 3520 3211 3521 3212
rect 3515 3210 3521 3211
rect 3546 3211 3547 3212
rect 3551 3211 3552 3215
rect 3546 3210 3552 3211
rect 1586 3206 1592 3207
rect 1894 3205 1900 3206
rect 1034 3203 1040 3204
rect 1034 3202 1035 3203
rect 430 3201 436 3202
rect 430 3197 431 3201
rect 435 3197 436 3201
rect 430 3196 436 3197
rect 550 3201 556 3202
rect 550 3197 551 3201
rect 555 3197 556 3201
rect 550 3196 556 3197
rect 670 3201 676 3202
rect 670 3197 671 3201
rect 675 3197 676 3201
rect 670 3196 676 3197
rect 798 3201 804 3202
rect 798 3197 799 3201
rect 803 3197 804 3201
rect 798 3196 804 3197
rect 934 3201 940 3202
rect 934 3197 935 3201
rect 939 3197 940 3201
rect 1016 3200 1035 3202
rect 1034 3199 1035 3200
rect 1039 3199 1040 3203
rect 1034 3198 1040 3199
rect 1078 3201 1084 3202
rect 934 3196 940 3197
rect 1078 3197 1079 3201
rect 1083 3197 1084 3201
rect 1078 3196 1084 3197
rect 1230 3201 1236 3202
rect 1230 3197 1231 3201
rect 1235 3197 1236 3201
rect 1230 3196 1236 3197
rect 1382 3201 1388 3202
rect 1382 3197 1383 3201
rect 1387 3197 1388 3201
rect 1382 3196 1388 3197
rect 1534 3201 1540 3202
rect 1534 3197 1535 3201
rect 1539 3197 1540 3201
rect 1894 3201 1895 3205
rect 1899 3201 1900 3205
rect 1894 3200 1900 3201
rect 2086 3205 2092 3206
rect 2086 3201 2087 3205
rect 2091 3201 2092 3205
rect 2086 3200 2092 3201
rect 2302 3205 2308 3206
rect 2302 3201 2303 3205
rect 2307 3201 2308 3205
rect 2302 3200 2308 3201
rect 2510 3205 2516 3206
rect 2510 3201 2511 3205
rect 2515 3201 2516 3205
rect 2510 3200 2516 3201
rect 2702 3205 2708 3206
rect 2702 3201 2703 3205
rect 2707 3201 2708 3205
rect 2702 3200 2708 3201
rect 2878 3205 2884 3206
rect 2878 3201 2879 3205
rect 2883 3201 2884 3205
rect 2878 3200 2884 3201
rect 3038 3205 3044 3206
rect 3038 3201 3039 3205
rect 3043 3201 3044 3205
rect 3038 3200 3044 3201
rect 3198 3205 3204 3206
rect 3198 3201 3199 3205
rect 3203 3201 3204 3205
rect 3198 3200 3204 3201
rect 3350 3205 3356 3206
rect 3350 3201 3351 3205
rect 3355 3201 3356 3205
rect 3350 3200 3356 3201
rect 3486 3205 3492 3206
rect 3486 3201 3487 3205
rect 3491 3201 3492 3205
rect 3486 3200 3492 3201
rect 1534 3196 1540 3197
rect 1862 3192 1868 3193
rect 3574 3192 3580 3193
rect 110 3188 116 3189
rect 1822 3188 1828 3189
rect 110 3184 111 3188
rect 115 3184 116 3188
rect 511 3187 517 3188
rect 511 3186 512 3187
rect 485 3184 512 3186
rect 110 3183 116 3184
rect 511 3183 512 3184
rect 516 3183 517 3187
rect 631 3187 637 3188
rect 631 3186 632 3187
rect 605 3184 632 3186
rect 511 3182 517 3183
rect 631 3183 632 3184
rect 636 3183 637 3187
rect 751 3187 757 3188
rect 751 3186 752 3187
rect 725 3184 752 3186
rect 631 3182 637 3183
rect 751 3183 752 3184
rect 756 3183 757 3187
rect 1023 3187 1029 3188
rect 1023 3186 1024 3187
rect 989 3184 1024 3186
rect 751 3182 757 3183
rect 1023 3183 1024 3184
rect 1028 3183 1029 3187
rect 1191 3187 1197 3188
rect 1191 3186 1192 3187
rect 1133 3184 1192 3186
rect 1023 3182 1029 3183
rect 1191 3183 1192 3184
rect 1196 3183 1197 3187
rect 1822 3184 1823 3188
rect 1827 3184 1828 3188
rect 1862 3188 1863 3192
rect 1867 3188 1868 3192
rect 1954 3191 1960 3192
rect 1954 3190 1955 3191
rect 1949 3188 1955 3190
rect 1862 3187 1868 3188
rect 1954 3187 1955 3188
rect 1959 3187 1960 3191
rect 2423 3191 2429 3192
rect 2423 3190 2424 3191
rect 2357 3188 2424 3190
rect 1954 3186 1960 3187
rect 1962 3187 1968 3188
rect 1191 3182 1197 3183
rect 1206 3183 1212 3184
rect 1206 3179 1207 3183
rect 1211 3182 1212 3183
rect 1479 3183 1485 3184
rect 1822 3183 1828 3184
rect 1962 3183 1963 3187
rect 1967 3186 1968 3187
rect 2423 3187 2424 3188
rect 2428 3187 2429 3191
rect 3279 3191 3285 3192
rect 3279 3190 3280 3191
rect 3253 3188 3280 3190
rect 2423 3186 2429 3187
rect 2678 3187 2684 3188
rect 1967 3184 2105 3186
rect 1967 3183 1968 3184
rect 1211 3180 1249 3182
rect 1211 3179 1212 3180
rect 1206 3178 1212 3179
rect 1479 3179 1480 3183
rect 1484 3182 1485 3183
rect 1962 3182 1968 3183
rect 2678 3183 2679 3187
rect 2683 3186 2684 3187
rect 2978 3187 2984 3188
rect 2683 3184 2721 3186
rect 2683 3183 2684 3184
rect 2678 3182 2684 3183
rect 2978 3183 2979 3187
rect 2983 3186 2984 3187
rect 3279 3187 3280 3188
rect 3284 3187 3285 3191
rect 3574 3188 3575 3192
rect 3579 3188 3580 3192
rect 3279 3186 3285 3187
rect 3295 3187 3301 3188
rect 3574 3187 3580 3188
rect 2983 3184 3057 3186
rect 2983 3183 2984 3184
rect 2978 3182 2984 3183
rect 3295 3183 3296 3187
rect 3300 3186 3301 3187
rect 3300 3184 3369 3186
rect 3300 3183 3301 3184
rect 3295 3182 3301 3183
rect 1484 3180 1553 3182
rect 1484 3179 1485 3180
rect 1479 3178 1485 3179
rect 1862 3175 1868 3176
rect 110 3171 116 3172
rect 110 3167 111 3171
rect 115 3167 116 3171
rect 1822 3171 1828 3172
rect 110 3166 116 3167
rect 732 3168 809 3170
rect 422 3161 428 3162
rect 422 3157 423 3161
rect 427 3157 428 3161
rect 422 3156 428 3157
rect 542 3161 548 3162
rect 542 3157 543 3161
rect 547 3157 548 3161
rect 542 3156 548 3157
rect 662 3161 668 3162
rect 662 3157 663 3161
rect 667 3157 668 3161
rect 662 3156 668 3157
rect 502 3155 508 3156
rect 502 3151 503 3155
rect 507 3154 508 3155
rect 732 3154 734 3168
rect 1822 3167 1823 3171
rect 1827 3167 1828 3171
rect 1862 3171 1863 3175
rect 1867 3171 1868 3175
rect 1862 3170 1868 3171
rect 3574 3175 3580 3176
rect 3574 3171 3575 3175
rect 3579 3171 3580 3175
rect 3574 3170 3580 3171
rect 1822 3166 1828 3167
rect 1886 3165 1892 3166
rect 790 3161 796 3162
rect 790 3157 791 3161
rect 795 3157 796 3161
rect 790 3156 796 3157
rect 926 3161 932 3162
rect 926 3157 927 3161
rect 931 3157 932 3161
rect 926 3156 932 3157
rect 1070 3161 1076 3162
rect 1070 3157 1071 3161
rect 1075 3157 1076 3161
rect 1070 3156 1076 3157
rect 1222 3161 1228 3162
rect 1222 3157 1223 3161
rect 1227 3157 1228 3161
rect 1222 3156 1228 3157
rect 1374 3161 1380 3162
rect 1374 3157 1375 3161
rect 1379 3157 1380 3161
rect 1374 3156 1380 3157
rect 1526 3161 1532 3162
rect 1526 3157 1527 3161
rect 1531 3157 1532 3161
rect 1886 3161 1887 3165
rect 1891 3161 1892 3165
rect 1886 3160 1892 3161
rect 2078 3165 2084 3166
rect 2078 3161 2079 3165
rect 2083 3161 2084 3165
rect 2078 3160 2084 3161
rect 2294 3165 2300 3166
rect 2294 3161 2295 3165
rect 2299 3161 2300 3165
rect 2294 3160 2300 3161
rect 2502 3165 2508 3166
rect 2502 3161 2503 3165
rect 2507 3161 2508 3165
rect 2502 3160 2508 3161
rect 2694 3165 2700 3166
rect 2694 3161 2695 3165
rect 2699 3161 2700 3165
rect 2694 3160 2700 3161
rect 2870 3165 2876 3166
rect 2870 3161 2871 3165
rect 2875 3161 2876 3165
rect 2870 3160 2876 3161
rect 3030 3165 3036 3166
rect 3030 3161 3031 3165
rect 3035 3161 3036 3165
rect 3030 3160 3036 3161
rect 3190 3165 3196 3166
rect 3190 3161 3191 3165
rect 3195 3161 3196 3165
rect 3190 3160 3196 3161
rect 3342 3165 3348 3166
rect 3342 3161 3343 3165
rect 3347 3161 3348 3165
rect 3342 3160 3348 3161
rect 3478 3165 3484 3166
rect 3478 3161 3479 3165
rect 3483 3161 3484 3165
rect 3478 3160 3484 3161
rect 1526 3156 1532 3157
rect 2542 3159 2548 3160
rect 507 3152 734 3154
rect 1414 3155 1420 3156
rect 507 3151 508 3152
rect 502 3150 508 3151
rect 1414 3151 1415 3155
rect 1419 3154 1420 3155
rect 1423 3155 1429 3156
rect 1423 3154 1424 3155
rect 1419 3152 1424 3154
rect 1419 3151 1420 3152
rect 1414 3150 1420 3151
rect 1423 3151 1424 3152
rect 1428 3151 1429 3155
rect 2542 3155 2543 3159
rect 2547 3158 2548 3159
rect 2551 3159 2557 3160
rect 2551 3158 2552 3159
rect 2547 3156 2552 3158
rect 2547 3155 2548 3156
rect 2542 3154 2548 3155
rect 2551 3155 2552 3156
rect 2556 3155 2557 3159
rect 2551 3154 2557 3155
rect 2910 3159 2916 3160
rect 2910 3155 2911 3159
rect 2915 3158 2916 3159
rect 2919 3159 2925 3160
rect 2919 3158 2920 3159
rect 2915 3156 2920 3158
rect 2915 3155 2916 3156
rect 2910 3154 2916 3155
rect 2919 3155 2920 3156
rect 2924 3155 2925 3159
rect 2919 3154 2925 3155
rect 3518 3159 3524 3160
rect 3518 3155 3519 3159
rect 3523 3158 3524 3159
rect 3527 3159 3533 3160
rect 3527 3158 3528 3159
rect 3523 3156 3528 3158
rect 3523 3155 3524 3156
rect 3518 3154 3524 3155
rect 3527 3155 3528 3156
rect 3532 3155 3533 3159
rect 3527 3154 3533 3155
rect 1423 3150 1429 3151
rect 1886 3139 1892 3140
rect 462 3135 468 3136
rect 462 3131 463 3135
rect 467 3131 468 3135
rect 462 3130 468 3131
rect 550 3135 556 3136
rect 550 3131 551 3135
rect 555 3131 556 3135
rect 550 3130 556 3131
rect 638 3135 644 3136
rect 638 3131 639 3135
rect 643 3131 644 3135
rect 638 3130 644 3131
rect 734 3135 740 3136
rect 734 3131 735 3135
rect 739 3131 740 3135
rect 734 3130 740 3131
rect 846 3135 852 3136
rect 846 3131 847 3135
rect 851 3131 852 3135
rect 846 3130 852 3131
rect 966 3135 972 3136
rect 966 3131 967 3135
rect 971 3131 972 3135
rect 966 3130 972 3131
rect 1094 3135 1100 3136
rect 1094 3131 1095 3135
rect 1099 3131 1100 3135
rect 1094 3130 1100 3131
rect 1230 3135 1236 3136
rect 1230 3131 1231 3135
rect 1235 3131 1236 3135
rect 1230 3130 1236 3131
rect 1374 3135 1380 3136
rect 1374 3131 1375 3135
rect 1379 3131 1380 3135
rect 1374 3130 1380 3131
rect 1518 3135 1524 3136
rect 1518 3131 1519 3135
rect 1523 3131 1524 3135
rect 1886 3135 1887 3139
rect 1891 3135 1892 3139
rect 1886 3134 1892 3135
rect 2078 3139 2084 3140
rect 2078 3135 2079 3139
rect 2083 3135 2084 3139
rect 2078 3134 2084 3135
rect 2294 3139 2300 3140
rect 2294 3135 2295 3139
rect 2299 3135 2300 3139
rect 2294 3134 2300 3135
rect 2502 3139 2508 3140
rect 2502 3135 2503 3139
rect 2507 3135 2508 3139
rect 2502 3134 2508 3135
rect 2694 3139 2700 3140
rect 2694 3135 2695 3139
rect 2699 3135 2700 3139
rect 2694 3134 2700 3135
rect 2870 3139 2876 3140
rect 2870 3135 2871 3139
rect 2875 3135 2876 3139
rect 2870 3134 2876 3135
rect 3038 3139 3044 3140
rect 3038 3135 3039 3139
rect 3043 3135 3044 3139
rect 3038 3134 3044 3135
rect 3190 3139 3196 3140
rect 3190 3135 3191 3139
rect 3195 3135 3196 3139
rect 3190 3134 3196 3135
rect 3342 3139 3348 3140
rect 3342 3135 3343 3139
rect 3347 3135 3348 3139
rect 3342 3134 3348 3135
rect 3478 3139 3484 3140
rect 3478 3135 3479 3139
rect 3483 3135 3484 3139
rect 3478 3134 3484 3135
rect 1518 3130 1524 3131
rect 2146 3131 2152 3132
rect 2146 3130 2147 3131
rect 1862 3129 1868 3130
rect 914 3127 920 3128
rect 110 3125 116 3126
rect 110 3121 111 3125
rect 115 3121 116 3125
rect 914 3123 915 3127
rect 919 3126 920 3127
rect 1034 3127 1040 3128
rect 919 3124 985 3126
rect 919 3123 920 3124
rect 914 3122 920 3123
rect 1034 3123 1035 3127
rect 1039 3126 1040 3127
rect 1039 3124 1113 3126
rect 1822 3125 1828 3126
rect 1039 3123 1040 3124
rect 1034 3122 1040 3123
rect 110 3120 116 3121
rect 1822 3121 1823 3125
rect 1827 3121 1828 3125
rect 1862 3125 1863 3129
rect 1867 3125 1868 3129
rect 2137 3128 2147 3130
rect 2146 3127 2147 3128
rect 2151 3127 2152 3131
rect 2762 3131 2768 3132
rect 2762 3130 2763 3131
rect 2753 3128 2763 3130
rect 2146 3126 2152 3127
rect 2762 3127 2763 3128
rect 2767 3127 2768 3131
rect 3410 3131 3416 3132
rect 3410 3130 3411 3131
rect 3401 3128 3411 3130
rect 2762 3126 2768 3127
rect 3410 3127 3411 3128
rect 3415 3127 3416 3131
rect 3410 3126 3416 3127
rect 3574 3129 3580 3130
rect 1862 3124 1868 3125
rect 3574 3125 3575 3129
rect 3579 3125 3580 3129
rect 3574 3124 3580 3125
rect 1822 3120 1828 3121
rect 2071 3115 2077 3116
rect 2071 3114 2072 3115
rect 1862 3112 1868 3113
rect 1949 3112 2072 3114
rect 543 3111 549 3112
rect 543 3110 544 3111
rect 110 3108 116 3109
rect 525 3108 544 3110
rect 110 3104 111 3108
rect 115 3104 116 3108
rect 543 3107 544 3108
rect 548 3107 549 3111
rect 631 3111 637 3112
rect 631 3110 632 3111
rect 613 3108 632 3110
rect 543 3106 549 3107
rect 631 3107 632 3108
rect 636 3107 637 3111
rect 727 3111 733 3112
rect 727 3110 728 3111
rect 701 3108 728 3110
rect 631 3106 637 3107
rect 727 3107 728 3108
rect 732 3107 733 3111
rect 839 3111 845 3112
rect 839 3110 840 3111
rect 797 3108 840 3110
rect 727 3106 733 3107
rect 839 3107 840 3108
rect 844 3107 845 3111
rect 959 3111 965 3112
rect 959 3110 960 3111
rect 909 3108 960 3110
rect 839 3106 845 3107
rect 959 3107 960 3108
rect 964 3107 965 3111
rect 959 3106 965 3107
rect 1162 3111 1168 3112
rect 1162 3107 1163 3111
rect 1167 3110 1168 3111
rect 1511 3111 1517 3112
rect 1511 3110 1512 3111
rect 1167 3108 1257 3110
rect 1437 3108 1512 3110
rect 1167 3107 1168 3108
rect 1162 3106 1168 3107
rect 1511 3107 1512 3108
rect 1516 3107 1517 3111
rect 1586 3111 1592 3112
rect 1586 3110 1587 3111
rect 1581 3108 1587 3110
rect 1511 3106 1517 3107
rect 1586 3107 1587 3108
rect 1591 3107 1592 3111
rect 1586 3106 1592 3107
rect 1822 3108 1828 3109
rect 110 3103 116 3104
rect 1822 3104 1823 3108
rect 1827 3104 1828 3108
rect 1862 3108 1863 3112
rect 1867 3108 1868 3112
rect 2071 3111 2072 3112
rect 2076 3111 2077 3115
rect 2071 3110 2077 3111
rect 2286 3115 2292 3116
rect 2286 3111 2287 3115
rect 2291 3114 2292 3115
rect 2362 3115 2368 3116
rect 2291 3112 2321 3114
rect 2291 3111 2292 3112
rect 2286 3110 2292 3111
rect 2362 3111 2363 3115
rect 2367 3114 2368 3115
rect 3031 3115 3037 3116
rect 3031 3114 3032 3115
rect 2367 3112 2529 3114
rect 2933 3112 3032 3114
rect 2367 3111 2368 3112
rect 2362 3110 2368 3111
rect 3031 3111 3032 3112
rect 3036 3111 3037 3115
rect 3183 3115 3189 3116
rect 3183 3114 3184 3115
rect 3101 3112 3184 3114
rect 3031 3110 3037 3111
rect 3183 3111 3184 3112
rect 3188 3111 3189 3115
rect 3335 3115 3341 3116
rect 3335 3114 3336 3115
rect 3253 3112 3336 3114
rect 3183 3110 3189 3111
rect 3335 3111 3336 3112
rect 3340 3111 3341 3115
rect 3554 3115 3560 3116
rect 3554 3114 3555 3115
rect 3541 3112 3555 3114
rect 3335 3110 3341 3111
rect 3554 3111 3555 3112
rect 3559 3111 3560 3115
rect 3554 3110 3560 3111
rect 3574 3112 3580 3113
rect 1862 3107 1868 3108
rect 3574 3108 3575 3112
rect 3579 3108 3580 3112
rect 3574 3107 3580 3108
rect 1822 3103 1828 3104
rect 1894 3099 1900 3100
rect 470 3095 476 3096
rect 470 3091 471 3095
rect 475 3091 476 3095
rect 470 3090 476 3091
rect 558 3095 564 3096
rect 558 3091 559 3095
rect 563 3091 564 3095
rect 558 3090 564 3091
rect 646 3095 652 3096
rect 646 3091 647 3095
rect 651 3091 652 3095
rect 646 3090 652 3091
rect 742 3095 748 3096
rect 742 3091 743 3095
rect 747 3091 748 3095
rect 742 3090 748 3091
rect 854 3095 860 3096
rect 854 3091 855 3095
rect 859 3091 860 3095
rect 854 3090 860 3091
rect 974 3095 980 3096
rect 974 3091 975 3095
rect 979 3091 980 3095
rect 974 3090 980 3091
rect 1102 3095 1108 3096
rect 1102 3091 1103 3095
rect 1107 3091 1108 3095
rect 1102 3090 1108 3091
rect 1238 3095 1244 3096
rect 1238 3091 1239 3095
rect 1243 3091 1244 3095
rect 1238 3090 1244 3091
rect 1382 3095 1388 3096
rect 1382 3091 1383 3095
rect 1387 3091 1388 3095
rect 1382 3090 1388 3091
rect 1526 3095 1532 3096
rect 1526 3091 1527 3095
rect 1531 3091 1532 3095
rect 1894 3095 1895 3099
rect 1899 3095 1900 3099
rect 1894 3094 1900 3095
rect 2086 3099 2092 3100
rect 2086 3095 2087 3099
rect 2091 3095 2092 3099
rect 2086 3094 2092 3095
rect 2302 3099 2308 3100
rect 2302 3095 2303 3099
rect 2307 3095 2308 3099
rect 2302 3094 2308 3095
rect 2510 3099 2516 3100
rect 2510 3095 2511 3099
rect 2515 3095 2516 3099
rect 2510 3094 2516 3095
rect 2702 3099 2708 3100
rect 2702 3095 2703 3099
rect 2707 3095 2708 3099
rect 2702 3094 2708 3095
rect 2878 3099 2884 3100
rect 2878 3095 2879 3099
rect 2883 3095 2884 3099
rect 2878 3094 2884 3095
rect 3046 3099 3052 3100
rect 3046 3095 3047 3099
rect 3051 3095 3052 3099
rect 3046 3094 3052 3095
rect 3198 3099 3204 3100
rect 3198 3095 3199 3099
rect 3203 3095 3204 3099
rect 3198 3094 3204 3095
rect 3350 3099 3356 3100
rect 3350 3095 3351 3099
rect 3355 3095 3356 3099
rect 3350 3094 3356 3095
rect 3486 3099 3492 3100
rect 3486 3095 3487 3099
rect 3491 3095 3492 3099
rect 3486 3094 3492 3095
rect 1526 3090 1532 3091
rect 1807 3087 1813 3088
rect 499 3083 508 3084
rect 499 3079 500 3083
rect 507 3079 508 3083
rect 499 3078 508 3079
rect 543 3083 549 3084
rect 543 3079 544 3083
rect 548 3082 549 3083
rect 587 3083 593 3084
rect 587 3082 588 3083
rect 548 3080 588 3082
rect 548 3079 549 3080
rect 543 3078 549 3079
rect 587 3079 588 3080
rect 592 3079 593 3083
rect 587 3078 593 3079
rect 631 3083 637 3084
rect 631 3079 632 3083
rect 636 3082 637 3083
rect 675 3083 681 3084
rect 675 3082 676 3083
rect 636 3080 676 3082
rect 636 3079 637 3080
rect 631 3078 637 3079
rect 675 3079 676 3080
rect 680 3079 681 3083
rect 675 3078 681 3079
rect 727 3083 733 3084
rect 727 3079 728 3083
rect 732 3082 733 3083
rect 771 3083 777 3084
rect 771 3082 772 3083
rect 732 3080 772 3082
rect 732 3079 733 3080
rect 727 3078 733 3079
rect 771 3079 772 3080
rect 776 3079 777 3083
rect 771 3078 777 3079
rect 839 3083 845 3084
rect 839 3079 840 3083
rect 844 3082 845 3083
rect 883 3083 889 3084
rect 883 3082 884 3083
rect 844 3080 884 3082
rect 844 3079 845 3080
rect 839 3078 845 3079
rect 883 3079 884 3080
rect 888 3079 889 3083
rect 883 3078 889 3079
rect 959 3083 965 3084
rect 959 3079 960 3083
rect 964 3082 965 3083
rect 1003 3083 1009 3084
rect 1003 3082 1004 3083
rect 964 3080 1004 3082
rect 964 3079 965 3080
rect 959 3078 965 3079
rect 1003 3079 1004 3080
rect 1008 3079 1009 3083
rect 1003 3078 1009 3079
rect 1131 3083 1137 3084
rect 1131 3079 1132 3083
rect 1136 3082 1137 3083
rect 1162 3083 1168 3084
rect 1162 3082 1163 3083
rect 1136 3080 1163 3082
rect 1136 3079 1137 3080
rect 1131 3078 1137 3079
rect 1162 3079 1163 3080
rect 1167 3079 1168 3083
rect 1162 3078 1168 3079
rect 1267 3083 1273 3084
rect 1267 3079 1268 3083
rect 1272 3082 1273 3083
rect 1367 3083 1373 3084
rect 1367 3082 1368 3083
rect 1272 3080 1368 3082
rect 1272 3079 1273 3080
rect 1267 3078 1273 3079
rect 1367 3079 1368 3080
rect 1372 3079 1373 3083
rect 1367 3078 1373 3079
rect 1411 3083 1420 3084
rect 1411 3079 1412 3083
rect 1419 3079 1420 3083
rect 1411 3078 1420 3079
rect 1511 3083 1517 3084
rect 1511 3079 1512 3083
rect 1516 3082 1517 3083
rect 1555 3083 1561 3084
rect 1555 3082 1556 3083
rect 1516 3080 1556 3082
rect 1516 3079 1517 3080
rect 1511 3078 1517 3079
rect 1555 3079 1556 3080
rect 1560 3079 1561 3083
rect 1807 3083 1808 3087
rect 1812 3086 1813 3087
rect 1923 3087 1929 3088
rect 1923 3086 1924 3087
rect 1812 3084 1924 3086
rect 1812 3083 1813 3084
rect 1807 3082 1813 3083
rect 1923 3083 1924 3084
rect 1928 3083 1929 3087
rect 1923 3082 1929 3083
rect 2071 3087 2077 3088
rect 2071 3083 2072 3087
rect 2076 3086 2077 3087
rect 2115 3087 2121 3088
rect 2115 3086 2116 3087
rect 2076 3084 2116 3086
rect 2076 3083 2077 3084
rect 2071 3082 2077 3083
rect 2115 3083 2116 3084
rect 2120 3083 2121 3087
rect 2115 3082 2121 3083
rect 2331 3087 2337 3088
rect 2331 3083 2332 3087
rect 2336 3086 2337 3087
rect 2362 3087 2368 3088
rect 2362 3086 2363 3087
rect 2336 3084 2363 3086
rect 2336 3083 2337 3084
rect 2331 3082 2337 3083
rect 2362 3083 2363 3084
rect 2367 3083 2368 3087
rect 2362 3082 2368 3083
rect 2539 3087 2548 3088
rect 2539 3083 2540 3087
rect 2547 3083 2548 3087
rect 2539 3082 2548 3083
rect 2663 3087 2669 3088
rect 2663 3083 2664 3087
rect 2668 3086 2669 3087
rect 2731 3087 2737 3088
rect 2731 3086 2732 3087
rect 2668 3084 2732 3086
rect 2668 3083 2669 3084
rect 2663 3082 2669 3083
rect 2731 3083 2732 3084
rect 2736 3083 2737 3087
rect 2731 3082 2737 3083
rect 2907 3087 2916 3088
rect 2907 3083 2908 3087
rect 2915 3083 2916 3087
rect 2907 3082 2916 3083
rect 3031 3087 3037 3088
rect 3031 3083 3032 3087
rect 3036 3086 3037 3087
rect 3075 3087 3081 3088
rect 3075 3086 3076 3087
rect 3036 3084 3076 3086
rect 3036 3083 3037 3084
rect 3031 3082 3037 3083
rect 3075 3083 3076 3084
rect 3080 3083 3081 3087
rect 3075 3082 3081 3083
rect 3183 3087 3189 3088
rect 3183 3083 3184 3087
rect 3188 3086 3189 3087
rect 3227 3087 3233 3088
rect 3227 3086 3228 3087
rect 3188 3084 3228 3086
rect 3188 3083 3189 3084
rect 3183 3082 3189 3083
rect 3227 3083 3228 3084
rect 3232 3083 3233 3087
rect 3227 3082 3233 3083
rect 3335 3087 3341 3088
rect 3335 3083 3336 3087
rect 3340 3086 3341 3087
rect 3379 3087 3385 3088
rect 3379 3086 3380 3087
rect 3340 3084 3380 3086
rect 3340 3083 3341 3084
rect 3335 3082 3341 3083
rect 3379 3083 3380 3084
rect 3384 3083 3385 3087
rect 3379 3082 3385 3083
rect 3515 3087 3524 3088
rect 3515 3083 3516 3087
rect 3523 3083 3524 3087
rect 3515 3082 3524 3083
rect 1555 3078 1561 3079
rect 179 3063 185 3064
rect 179 3059 180 3063
rect 184 3062 185 3063
rect 222 3063 228 3064
rect 222 3062 223 3063
rect 184 3060 223 3062
rect 184 3059 185 3060
rect 179 3058 185 3059
rect 222 3059 223 3060
rect 227 3059 228 3063
rect 222 3058 228 3059
rect 230 3063 236 3064
rect 230 3059 231 3063
rect 235 3062 236 3063
rect 267 3063 273 3064
rect 267 3062 268 3063
rect 235 3060 268 3062
rect 235 3059 236 3060
rect 230 3058 236 3059
rect 267 3059 268 3060
rect 272 3059 273 3063
rect 267 3058 273 3059
rect 311 3063 317 3064
rect 311 3059 312 3063
rect 316 3062 317 3063
rect 355 3063 361 3064
rect 355 3062 356 3063
rect 316 3060 356 3062
rect 316 3059 317 3060
rect 311 3058 317 3059
rect 355 3059 356 3060
rect 360 3059 361 3063
rect 355 3058 361 3059
rect 391 3063 397 3064
rect 391 3059 392 3063
rect 396 3062 397 3063
rect 443 3063 449 3064
rect 443 3062 444 3063
rect 396 3060 444 3062
rect 396 3059 397 3060
rect 391 3058 397 3059
rect 443 3059 444 3060
rect 448 3059 449 3063
rect 443 3058 449 3059
rect 479 3063 485 3064
rect 479 3059 480 3063
rect 484 3062 485 3063
rect 531 3063 537 3064
rect 531 3062 532 3063
rect 484 3060 532 3062
rect 484 3059 485 3060
rect 479 3058 485 3059
rect 531 3059 532 3060
rect 536 3059 537 3063
rect 531 3058 537 3059
rect 567 3063 573 3064
rect 567 3059 568 3063
rect 572 3062 573 3063
rect 619 3063 625 3064
rect 619 3062 620 3063
rect 572 3060 620 3062
rect 572 3059 573 3060
rect 567 3058 573 3059
rect 619 3059 620 3060
rect 624 3059 625 3063
rect 619 3058 625 3059
rect 655 3063 661 3064
rect 655 3059 656 3063
rect 660 3062 661 3063
rect 707 3063 713 3064
rect 707 3062 708 3063
rect 660 3060 708 3062
rect 660 3059 661 3060
rect 655 3058 661 3059
rect 707 3059 708 3060
rect 712 3059 713 3063
rect 707 3058 713 3059
rect 743 3063 749 3064
rect 743 3059 744 3063
rect 748 3062 749 3063
rect 795 3063 801 3064
rect 795 3062 796 3063
rect 748 3060 796 3062
rect 748 3059 749 3060
rect 743 3058 749 3059
rect 795 3059 796 3060
rect 800 3059 801 3063
rect 795 3058 801 3059
rect 831 3063 837 3064
rect 831 3059 832 3063
rect 836 3062 837 3063
rect 883 3063 889 3064
rect 883 3062 884 3063
rect 836 3060 884 3062
rect 836 3059 837 3060
rect 831 3058 837 3059
rect 883 3059 884 3060
rect 888 3059 889 3063
rect 883 3058 889 3059
rect 919 3063 925 3064
rect 919 3059 920 3063
rect 924 3062 925 3063
rect 971 3063 977 3064
rect 971 3062 972 3063
rect 924 3060 972 3062
rect 924 3059 925 3060
rect 919 3058 925 3059
rect 971 3059 972 3060
rect 976 3059 977 3063
rect 971 3058 977 3059
rect 1007 3063 1013 3064
rect 1007 3059 1008 3063
rect 1012 3062 1013 3063
rect 1059 3063 1065 3064
rect 1059 3062 1060 3063
rect 1012 3060 1060 3062
rect 1012 3059 1013 3060
rect 1007 3058 1013 3059
rect 1059 3059 1060 3060
rect 1064 3059 1065 3063
rect 1059 3058 1065 3059
rect 1090 3063 1096 3064
rect 1090 3059 1091 3063
rect 1095 3062 1096 3063
rect 1147 3063 1153 3064
rect 1147 3062 1148 3063
rect 1095 3060 1148 3062
rect 1095 3059 1096 3060
rect 1090 3058 1096 3059
rect 1147 3059 1148 3060
rect 1152 3059 1153 3063
rect 1147 3058 1153 3059
rect 1183 3063 1189 3064
rect 1183 3059 1184 3063
rect 1188 3062 1189 3063
rect 1235 3063 1241 3064
rect 1235 3062 1236 3063
rect 1188 3060 1236 3062
rect 1188 3059 1189 3060
rect 1183 3058 1189 3059
rect 1235 3059 1236 3060
rect 1240 3059 1241 3063
rect 1235 3058 1241 3059
rect 1271 3063 1277 3064
rect 1271 3059 1272 3063
rect 1276 3062 1277 3063
rect 1323 3063 1329 3064
rect 1323 3062 1324 3063
rect 1276 3060 1324 3062
rect 1276 3059 1277 3060
rect 1271 3058 1277 3059
rect 1323 3059 1324 3060
rect 1328 3059 1329 3063
rect 1323 3058 1329 3059
rect 1359 3063 1365 3064
rect 1359 3059 1360 3063
rect 1364 3062 1365 3063
rect 1411 3063 1417 3064
rect 1411 3062 1412 3063
rect 1364 3060 1412 3062
rect 1364 3059 1365 3060
rect 1359 3058 1365 3059
rect 1411 3059 1412 3060
rect 1416 3059 1417 3063
rect 1411 3058 1417 3059
rect 1499 3063 1505 3064
rect 1499 3059 1500 3063
rect 1504 3062 1505 3063
rect 1538 3063 1544 3064
rect 1538 3062 1539 3063
rect 1504 3060 1539 3062
rect 1504 3059 1505 3060
rect 1499 3058 1505 3059
rect 1538 3059 1539 3060
rect 1543 3059 1544 3063
rect 1538 3058 1544 3059
rect 1586 3063 1593 3064
rect 1586 3059 1587 3063
rect 1592 3059 1593 3063
rect 1586 3058 1593 3059
rect 1675 3063 1681 3064
rect 1675 3059 1676 3063
rect 1680 3062 1681 3063
rect 1698 3063 1704 3064
rect 1698 3062 1699 3063
rect 1680 3060 1699 3062
rect 1680 3059 1681 3060
rect 1675 3058 1681 3059
rect 1698 3059 1699 3060
rect 1703 3059 1704 3063
rect 1698 3058 1704 3059
rect 1711 3063 1717 3064
rect 1711 3059 1712 3063
rect 1716 3062 1717 3063
rect 1763 3063 1769 3064
rect 1763 3062 1764 3063
rect 1716 3060 1764 3062
rect 1716 3059 1717 3060
rect 1711 3058 1717 3059
rect 1763 3059 1764 3060
rect 1768 3059 1769 3063
rect 1763 3058 1769 3059
rect 2283 3063 2292 3064
rect 2283 3059 2284 3063
rect 2291 3059 2292 3063
rect 2283 3058 2292 3059
rect 2375 3063 2381 3064
rect 2375 3059 2376 3063
rect 2380 3062 2381 3063
rect 2451 3063 2457 3064
rect 2451 3062 2452 3063
rect 2380 3060 2452 3062
rect 2380 3059 2381 3060
rect 2375 3058 2381 3059
rect 2451 3059 2452 3060
rect 2456 3059 2457 3063
rect 2451 3058 2457 3059
rect 2619 3063 2625 3064
rect 2619 3059 2620 3063
rect 2624 3062 2625 3063
rect 2671 3063 2677 3064
rect 2671 3062 2672 3063
rect 2624 3060 2672 3062
rect 2624 3059 2625 3060
rect 2619 3058 2625 3059
rect 2671 3059 2672 3060
rect 2676 3059 2677 3063
rect 2671 3058 2677 3059
rect 2779 3063 2788 3064
rect 2779 3059 2780 3063
rect 2787 3059 2788 3063
rect 2779 3058 2788 3059
rect 2930 3063 2936 3064
rect 2930 3059 2931 3063
rect 2935 3062 2936 3063
rect 2947 3063 2953 3064
rect 2947 3062 2948 3063
rect 2935 3060 2948 3062
rect 2935 3059 2936 3060
rect 2930 3058 2936 3059
rect 2947 3059 2948 3060
rect 2952 3059 2953 3063
rect 2947 3058 2953 3059
rect 3023 3063 3029 3064
rect 3023 3059 3024 3063
rect 3028 3062 3029 3063
rect 3115 3063 3121 3064
rect 3115 3062 3116 3063
rect 3028 3060 3116 3062
rect 3028 3059 3029 3060
rect 3023 3058 3029 3059
rect 3115 3059 3116 3060
rect 3120 3059 3121 3063
rect 3115 3058 3121 3059
rect 150 3053 156 3054
rect 150 3049 151 3053
rect 155 3049 156 3053
rect 150 3048 156 3049
rect 238 3053 244 3054
rect 238 3049 239 3053
rect 243 3049 244 3053
rect 238 3048 244 3049
rect 326 3053 332 3054
rect 326 3049 327 3053
rect 331 3049 332 3053
rect 326 3048 332 3049
rect 414 3053 420 3054
rect 414 3049 415 3053
rect 419 3049 420 3053
rect 414 3048 420 3049
rect 502 3053 508 3054
rect 502 3049 503 3053
rect 507 3049 508 3053
rect 502 3048 508 3049
rect 590 3053 596 3054
rect 590 3049 591 3053
rect 595 3049 596 3053
rect 590 3048 596 3049
rect 678 3053 684 3054
rect 678 3049 679 3053
rect 683 3049 684 3053
rect 678 3048 684 3049
rect 766 3053 772 3054
rect 766 3049 767 3053
rect 771 3049 772 3053
rect 766 3048 772 3049
rect 854 3053 860 3054
rect 854 3049 855 3053
rect 859 3049 860 3053
rect 854 3048 860 3049
rect 942 3053 948 3054
rect 942 3049 943 3053
rect 947 3049 948 3053
rect 942 3048 948 3049
rect 1030 3053 1036 3054
rect 1030 3049 1031 3053
rect 1035 3049 1036 3053
rect 1030 3048 1036 3049
rect 1118 3053 1124 3054
rect 1118 3049 1119 3053
rect 1123 3049 1124 3053
rect 1118 3048 1124 3049
rect 1206 3053 1212 3054
rect 1206 3049 1207 3053
rect 1211 3049 1212 3053
rect 1206 3048 1212 3049
rect 1294 3053 1300 3054
rect 1294 3049 1295 3053
rect 1299 3049 1300 3053
rect 1294 3048 1300 3049
rect 1382 3053 1388 3054
rect 1382 3049 1383 3053
rect 1387 3049 1388 3053
rect 1382 3048 1388 3049
rect 1470 3053 1476 3054
rect 1470 3049 1471 3053
rect 1475 3049 1476 3053
rect 1470 3048 1476 3049
rect 1558 3053 1564 3054
rect 1558 3049 1559 3053
rect 1563 3049 1564 3053
rect 1558 3048 1564 3049
rect 1646 3053 1652 3054
rect 1646 3049 1647 3053
rect 1651 3049 1652 3053
rect 1646 3048 1652 3049
rect 1734 3053 1740 3054
rect 1734 3049 1735 3053
rect 1739 3049 1740 3053
rect 1734 3048 1740 3049
rect 2254 3053 2260 3054
rect 2254 3049 2255 3053
rect 2259 3049 2260 3053
rect 2254 3048 2260 3049
rect 2422 3053 2428 3054
rect 2422 3049 2423 3053
rect 2427 3049 2428 3053
rect 2422 3048 2428 3049
rect 2590 3053 2596 3054
rect 2590 3049 2591 3053
rect 2595 3049 2596 3053
rect 2590 3048 2596 3049
rect 2750 3053 2756 3054
rect 2750 3049 2751 3053
rect 2755 3049 2756 3053
rect 2750 3048 2756 3049
rect 2918 3053 2924 3054
rect 2918 3049 2919 3053
rect 2923 3049 2924 3053
rect 2918 3048 2924 3049
rect 3086 3053 3092 3054
rect 3086 3049 3087 3053
rect 3091 3049 3092 3053
rect 3086 3048 3092 3049
rect 110 3040 116 3041
rect 1822 3040 1828 3041
rect 110 3036 111 3040
rect 115 3036 116 3040
rect 311 3039 317 3040
rect 311 3038 312 3039
rect 293 3036 312 3038
rect 110 3035 116 3036
rect 230 3035 236 3036
rect 230 3034 231 3035
rect 205 3032 231 3034
rect 230 3031 231 3032
rect 235 3031 236 3035
rect 311 3035 312 3036
rect 316 3035 317 3039
rect 391 3039 397 3040
rect 391 3038 392 3039
rect 381 3036 392 3038
rect 311 3034 317 3035
rect 391 3035 392 3036
rect 396 3035 397 3039
rect 479 3039 485 3040
rect 479 3038 480 3039
rect 469 3036 480 3038
rect 391 3034 397 3035
rect 479 3035 480 3036
rect 484 3035 485 3039
rect 567 3039 573 3040
rect 567 3038 568 3039
rect 557 3036 568 3038
rect 479 3034 485 3035
rect 567 3035 568 3036
rect 572 3035 573 3039
rect 655 3039 661 3040
rect 655 3038 656 3039
rect 645 3036 656 3038
rect 567 3034 573 3035
rect 655 3035 656 3036
rect 660 3035 661 3039
rect 743 3039 749 3040
rect 743 3038 744 3039
rect 733 3036 744 3038
rect 655 3034 661 3035
rect 743 3035 744 3036
rect 748 3035 749 3039
rect 831 3039 837 3040
rect 831 3038 832 3039
rect 821 3036 832 3038
rect 743 3034 749 3035
rect 831 3035 832 3036
rect 836 3035 837 3039
rect 919 3039 925 3040
rect 919 3038 920 3039
rect 909 3036 920 3038
rect 831 3034 837 3035
rect 919 3035 920 3036
rect 924 3035 925 3039
rect 1007 3039 1013 3040
rect 1007 3038 1008 3039
rect 997 3036 1008 3038
rect 919 3034 925 3035
rect 1007 3035 1008 3036
rect 1012 3035 1013 3039
rect 1090 3039 1096 3040
rect 1090 3038 1091 3039
rect 1085 3036 1091 3038
rect 1007 3034 1013 3035
rect 1090 3035 1091 3036
rect 1095 3035 1096 3039
rect 1183 3039 1189 3040
rect 1183 3038 1184 3039
rect 1173 3036 1184 3038
rect 1090 3034 1096 3035
rect 1183 3035 1184 3036
rect 1188 3035 1189 3039
rect 1271 3039 1277 3040
rect 1271 3038 1272 3039
rect 1261 3036 1272 3038
rect 1183 3034 1189 3035
rect 1271 3035 1272 3036
rect 1276 3035 1277 3039
rect 1359 3039 1365 3040
rect 1359 3038 1360 3039
rect 1349 3036 1360 3038
rect 1271 3034 1277 3035
rect 1359 3035 1360 3036
rect 1364 3035 1365 3039
rect 1711 3039 1717 3040
rect 1711 3038 1712 3039
rect 1701 3036 1712 3038
rect 1359 3034 1365 3035
rect 1367 3035 1373 3036
rect 230 3030 236 3031
rect 1367 3031 1368 3035
rect 1372 3034 1373 3035
rect 1538 3035 1544 3036
rect 1372 3032 1401 3034
rect 1372 3031 1373 3032
rect 1367 3030 1373 3031
rect 1538 3031 1539 3035
rect 1543 3034 1544 3035
rect 1711 3035 1712 3036
rect 1716 3035 1717 3039
rect 1807 3039 1813 3040
rect 1807 3038 1808 3039
rect 1789 3036 1808 3038
rect 1711 3034 1717 3035
rect 1807 3035 1808 3036
rect 1812 3035 1813 3039
rect 1822 3036 1823 3040
rect 1827 3036 1828 3040
rect 1822 3035 1828 3036
rect 1862 3040 1868 3041
rect 3574 3040 3580 3041
rect 1862 3036 1863 3040
rect 1867 3036 1868 3040
rect 2375 3039 2381 3040
rect 2375 3038 2376 3039
rect 2309 3036 2376 3038
rect 1862 3035 1868 3036
rect 2375 3035 2376 3036
rect 2380 3035 2381 3039
rect 2663 3039 2669 3040
rect 2663 3038 2664 3039
rect 2645 3036 2664 3038
rect 1807 3034 1813 3035
rect 2375 3034 2381 3035
rect 2663 3035 2664 3036
rect 2668 3035 2669 3039
rect 3023 3039 3029 3040
rect 3023 3038 3024 3039
rect 2973 3036 3024 3038
rect 2663 3034 2669 3035
rect 2671 3035 2677 3036
rect 1543 3032 1577 3034
rect 1543 3031 1544 3032
rect 1538 3030 1544 3031
rect 2671 3031 2672 3035
rect 2676 3034 2677 3035
rect 3023 3035 3024 3036
rect 3028 3035 3029 3039
rect 3574 3036 3575 3040
rect 3579 3036 3580 3040
rect 3023 3034 3029 3035
rect 3034 3035 3040 3036
rect 3574 3035 3580 3036
rect 2676 3032 2769 3034
rect 2676 3031 2677 3032
rect 2671 3030 2677 3031
rect 3034 3031 3035 3035
rect 3039 3034 3040 3035
rect 3039 3032 3105 3034
rect 3039 3031 3040 3032
rect 3034 3030 3040 3031
rect 110 3023 116 3024
rect 110 3019 111 3023
rect 115 3019 116 3023
rect 1542 3023 1548 3024
rect 1542 3022 1543 3023
rect 1521 3020 1543 3022
rect 110 3018 116 3019
rect 1542 3019 1543 3020
rect 1547 3019 1548 3023
rect 1542 3018 1548 3019
rect 1822 3023 1828 3024
rect 1822 3019 1823 3023
rect 1827 3019 1828 3023
rect 1822 3018 1828 3019
rect 1862 3023 1868 3024
rect 1862 3019 1863 3023
rect 1867 3019 1868 3023
rect 2498 3023 2504 3024
rect 2498 3022 2499 3023
rect 2473 3020 2499 3022
rect 1862 3018 1868 3019
rect 2498 3019 2499 3020
rect 2503 3019 2504 3023
rect 2498 3018 2504 3019
rect 3574 3023 3580 3024
rect 3574 3019 3575 3023
rect 3579 3019 3580 3023
rect 3574 3018 3580 3019
rect 142 3013 148 3014
rect 142 3009 143 3013
rect 147 3009 148 3013
rect 142 3008 148 3009
rect 230 3013 236 3014
rect 230 3009 231 3013
rect 235 3009 236 3013
rect 230 3008 236 3009
rect 318 3013 324 3014
rect 318 3009 319 3013
rect 323 3009 324 3013
rect 318 3008 324 3009
rect 406 3013 412 3014
rect 406 3009 407 3013
rect 411 3009 412 3013
rect 406 3008 412 3009
rect 494 3013 500 3014
rect 494 3009 495 3013
rect 499 3009 500 3013
rect 494 3008 500 3009
rect 582 3013 588 3014
rect 582 3009 583 3013
rect 587 3009 588 3013
rect 582 3008 588 3009
rect 670 3013 676 3014
rect 670 3009 671 3013
rect 675 3009 676 3013
rect 670 3008 676 3009
rect 758 3013 764 3014
rect 758 3009 759 3013
rect 763 3009 764 3013
rect 758 3008 764 3009
rect 846 3013 852 3014
rect 846 3009 847 3013
rect 851 3009 852 3013
rect 846 3008 852 3009
rect 934 3013 940 3014
rect 934 3009 935 3013
rect 939 3009 940 3013
rect 934 3008 940 3009
rect 1022 3013 1028 3014
rect 1022 3009 1023 3013
rect 1027 3009 1028 3013
rect 1022 3008 1028 3009
rect 1110 3013 1116 3014
rect 1110 3009 1111 3013
rect 1115 3009 1116 3013
rect 1110 3008 1116 3009
rect 1198 3013 1204 3014
rect 1198 3009 1199 3013
rect 1203 3009 1204 3013
rect 1198 3008 1204 3009
rect 1286 3013 1292 3014
rect 1286 3009 1287 3013
rect 1291 3009 1292 3013
rect 1286 3008 1292 3009
rect 1374 3013 1380 3014
rect 1374 3009 1375 3013
rect 1379 3009 1380 3013
rect 1374 3008 1380 3009
rect 1462 3013 1468 3014
rect 1462 3009 1463 3013
rect 1467 3009 1468 3013
rect 1462 3008 1468 3009
rect 1550 3013 1556 3014
rect 1550 3009 1551 3013
rect 1555 3009 1556 3013
rect 1550 3008 1556 3009
rect 1638 3013 1644 3014
rect 1638 3009 1639 3013
rect 1643 3009 1644 3013
rect 1638 3008 1644 3009
rect 1726 3013 1732 3014
rect 1726 3009 1727 3013
rect 1731 3009 1732 3013
rect 1726 3008 1732 3009
rect 2246 3013 2252 3014
rect 2246 3009 2247 3013
rect 2251 3009 2252 3013
rect 2246 3008 2252 3009
rect 2414 3013 2420 3014
rect 2414 3009 2415 3013
rect 2419 3009 2420 3013
rect 2414 3008 2420 3009
rect 2582 3013 2588 3014
rect 2582 3009 2583 3013
rect 2587 3009 2588 3013
rect 2582 3008 2588 3009
rect 2742 3013 2748 3014
rect 2742 3009 2743 3013
rect 2747 3009 2748 3013
rect 2742 3008 2748 3009
rect 2910 3013 2916 3014
rect 2910 3009 2911 3013
rect 2915 3009 2916 3013
rect 2910 3008 2916 3009
rect 3078 3013 3084 3014
rect 3078 3009 3079 3013
rect 3083 3009 3084 3013
rect 3078 3008 3084 3009
rect 2238 2987 2244 2988
rect 1406 2983 1412 2984
rect 1406 2979 1407 2983
rect 1411 2979 1412 2983
rect 1406 2978 1412 2979
rect 1518 2983 1524 2984
rect 1518 2979 1519 2983
rect 1523 2979 1524 2983
rect 1518 2978 1524 2979
rect 1630 2983 1636 2984
rect 1630 2979 1631 2983
rect 1635 2979 1636 2983
rect 1630 2978 1636 2979
rect 1726 2983 1732 2984
rect 1726 2979 1727 2983
rect 1731 2979 1732 2983
rect 2238 2983 2239 2987
rect 2243 2983 2244 2987
rect 2238 2982 2244 2983
rect 2462 2987 2468 2988
rect 2462 2983 2463 2987
rect 2467 2983 2468 2987
rect 2462 2982 2468 2983
rect 2670 2987 2676 2988
rect 2670 2983 2671 2987
rect 2675 2983 2676 2987
rect 2670 2982 2676 2983
rect 2862 2987 2868 2988
rect 2862 2983 2863 2987
rect 2867 2983 2868 2987
rect 2862 2982 2868 2983
rect 3030 2987 3036 2988
rect 3030 2983 3031 2987
rect 3035 2983 3036 2987
rect 3030 2982 3036 2983
rect 3190 2987 3196 2988
rect 3190 2983 3191 2987
rect 3195 2983 3196 2987
rect 3190 2982 3196 2983
rect 3342 2987 3348 2988
rect 3342 2983 3343 2987
rect 3347 2983 3348 2987
rect 3342 2982 3348 2983
rect 3478 2987 3484 2988
rect 3478 2983 3479 2987
rect 3483 2983 3484 2987
rect 3478 2982 3484 2983
rect 1726 2978 1732 2979
rect 2930 2979 2936 2980
rect 2930 2978 2931 2979
rect 1862 2977 1868 2978
rect 1698 2975 1704 2976
rect 1698 2974 1699 2975
rect 110 2973 116 2974
rect 110 2969 111 2973
rect 115 2969 116 2973
rect 1689 2972 1699 2974
rect 1698 2971 1699 2972
rect 1703 2971 1704 2975
rect 1698 2970 1704 2971
rect 1822 2973 1828 2974
rect 110 2968 116 2969
rect 1822 2969 1823 2973
rect 1827 2969 1828 2973
rect 1862 2973 1863 2977
rect 1867 2973 1868 2977
rect 2921 2976 2931 2978
rect 2930 2975 2931 2976
rect 2935 2975 2936 2979
rect 2930 2974 2936 2975
rect 3574 2977 3580 2978
rect 1862 2972 1868 2973
rect 3574 2973 3575 2977
rect 3579 2973 3580 2977
rect 3574 2972 3580 2973
rect 1822 2968 1828 2969
rect 2306 2963 2312 2964
rect 2306 2962 2307 2963
rect 1862 2960 1868 2961
rect 2301 2960 2307 2962
rect 1478 2959 1484 2960
rect 110 2956 116 2957
rect 110 2952 111 2956
rect 115 2952 116 2956
rect 110 2951 116 2952
rect 1468 2950 1470 2957
rect 1478 2955 1479 2959
rect 1483 2958 1484 2959
rect 1703 2959 1709 2960
rect 1483 2956 1545 2958
rect 1483 2955 1484 2956
rect 1478 2954 1484 2955
rect 1703 2955 1704 2959
rect 1708 2958 1709 2959
rect 1708 2956 1753 2958
rect 1822 2956 1828 2957
rect 1708 2955 1709 2956
rect 1703 2954 1709 2955
rect 1822 2952 1823 2956
rect 1827 2952 1828 2956
rect 1862 2956 1863 2960
rect 1867 2956 1868 2960
rect 2306 2959 2307 2960
rect 2311 2959 2312 2963
rect 2306 2958 2312 2959
rect 2350 2963 2356 2964
rect 2350 2959 2351 2963
rect 2355 2962 2356 2963
rect 2855 2963 2861 2964
rect 2855 2962 2856 2963
rect 2355 2960 2489 2962
rect 2733 2960 2856 2962
rect 2355 2959 2356 2960
rect 2350 2958 2356 2959
rect 2855 2959 2856 2960
rect 2860 2959 2861 2963
rect 2855 2958 2861 2959
rect 2958 2963 2964 2964
rect 2958 2959 2959 2963
rect 2963 2962 2964 2963
rect 3098 2963 3104 2964
rect 2963 2960 3057 2962
rect 2963 2959 2964 2960
rect 2958 2958 2964 2959
rect 3098 2959 3099 2963
rect 3103 2962 3104 2963
rect 3258 2963 3264 2964
rect 3103 2960 3217 2962
rect 3103 2959 3104 2960
rect 3098 2958 3104 2959
rect 3258 2959 3259 2963
rect 3263 2962 3264 2963
rect 3546 2963 3552 2964
rect 3546 2962 3547 2963
rect 3263 2960 3369 2962
rect 3541 2960 3547 2962
rect 3263 2959 3264 2960
rect 3258 2958 3264 2959
rect 3546 2959 3547 2960
rect 3551 2959 3552 2963
rect 3546 2958 3552 2959
rect 3574 2960 3580 2961
rect 1862 2955 1868 2956
rect 3574 2956 3575 2960
rect 3579 2956 3580 2960
rect 3574 2955 3580 2956
rect 1498 2951 1504 2952
rect 1822 2951 1828 2952
rect 1498 2950 1499 2951
rect 1468 2948 1499 2950
rect 1498 2947 1499 2948
rect 1503 2947 1504 2951
rect 1498 2946 1504 2947
rect 2246 2947 2252 2948
rect 1414 2943 1420 2944
rect 1414 2939 1415 2943
rect 1419 2939 1420 2943
rect 1414 2938 1420 2939
rect 1526 2943 1532 2944
rect 1526 2939 1527 2943
rect 1531 2939 1532 2943
rect 1526 2938 1532 2939
rect 1638 2943 1644 2944
rect 1638 2939 1639 2943
rect 1643 2939 1644 2943
rect 1638 2938 1644 2939
rect 1734 2943 1740 2944
rect 1734 2939 1735 2943
rect 1739 2939 1740 2943
rect 2246 2943 2247 2947
rect 2251 2943 2252 2947
rect 2246 2942 2252 2943
rect 2470 2947 2476 2948
rect 2470 2943 2471 2947
rect 2475 2943 2476 2947
rect 2470 2942 2476 2943
rect 2678 2947 2684 2948
rect 2678 2943 2679 2947
rect 2683 2943 2684 2947
rect 2678 2942 2684 2943
rect 2870 2947 2876 2948
rect 2870 2943 2871 2947
rect 2875 2943 2876 2947
rect 2870 2942 2876 2943
rect 3038 2947 3044 2948
rect 3038 2943 3039 2947
rect 3043 2943 3044 2947
rect 3038 2942 3044 2943
rect 3198 2947 3204 2948
rect 3198 2943 3199 2947
rect 3203 2943 3204 2947
rect 3198 2942 3204 2943
rect 3350 2947 3356 2948
rect 3350 2943 3351 2947
rect 3355 2943 3356 2947
rect 3350 2942 3356 2943
rect 3486 2947 3492 2948
rect 3486 2943 3487 2947
rect 3491 2943 3492 2947
rect 3486 2942 3492 2943
rect 1734 2938 1740 2939
rect 2275 2935 2281 2936
rect 1443 2931 1449 2932
rect 1443 2927 1444 2931
rect 1448 2930 1449 2931
rect 1478 2931 1484 2932
rect 1478 2930 1479 2931
rect 1448 2928 1479 2930
rect 1448 2927 1449 2928
rect 1443 2926 1449 2927
rect 1478 2927 1479 2928
rect 1483 2927 1484 2931
rect 1542 2931 1548 2932
rect 1478 2926 1484 2927
rect 1534 2927 1540 2928
rect 1534 2926 1535 2927
rect 1488 2924 1535 2926
rect 1488 2922 1490 2924
rect 1534 2923 1535 2924
rect 1539 2923 1540 2927
rect 1542 2927 1543 2931
rect 1547 2930 1548 2931
rect 1555 2931 1561 2932
rect 1555 2930 1556 2931
rect 1547 2928 1556 2930
rect 1547 2927 1548 2928
rect 1542 2926 1548 2927
rect 1555 2927 1556 2928
rect 1560 2927 1561 2931
rect 1555 2926 1561 2927
rect 1667 2931 1673 2932
rect 1667 2927 1668 2931
rect 1672 2930 1673 2931
rect 1703 2931 1709 2932
rect 1703 2930 1704 2931
rect 1672 2928 1704 2930
rect 1672 2927 1673 2928
rect 1667 2926 1673 2927
rect 1703 2927 1704 2928
rect 1708 2927 1709 2931
rect 1703 2926 1709 2927
rect 1762 2931 1769 2932
rect 1762 2927 1763 2931
rect 1768 2927 1769 2931
rect 2275 2931 2276 2935
rect 2280 2934 2281 2935
rect 2350 2935 2356 2936
rect 2350 2934 2351 2935
rect 2280 2932 2351 2934
rect 2280 2931 2281 2932
rect 2275 2930 2281 2931
rect 2350 2931 2351 2932
rect 2355 2931 2356 2935
rect 2350 2930 2356 2931
rect 2498 2935 2505 2936
rect 2498 2931 2499 2935
rect 2504 2931 2505 2935
rect 2498 2930 2505 2931
rect 2707 2935 2716 2936
rect 2707 2931 2708 2935
rect 2715 2931 2716 2935
rect 2707 2930 2716 2931
rect 2855 2935 2861 2936
rect 2855 2931 2856 2935
rect 2860 2934 2861 2935
rect 2899 2935 2905 2936
rect 2899 2934 2900 2935
rect 2860 2932 2900 2934
rect 2860 2931 2861 2932
rect 2855 2930 2861 2931
rect 2899 2931 2900 2932
rect 2904 2931 2905 2935
rect 2899 2930 2905 2931
rect 3067 2935 3073 2936
rect 3067 2931 3068 2935
rect 3072 2934 3073 2935
rect 3098 2935 3104 2936
rect 3098 2934 3099 2935
rect 3072 2932 3099 2934
rect 3072 2931 3073 2932
rect 3067 2930 3073 2931
rect 3098 2931 3099 2932
rect 3103 2931 3104 2935
rect 3098 2930 3104 2931
rect 3227 2935 3233 2936
rect 3227 2931 3228 2935
rect 3232 2934 3233 2935
rect 3258 2935 3264 2936
rect 3258 2934 3259 2935
rect 3232 2932 3259 2934
rect 3232 2931 3233 2932
rect 3227 2930 3233 2931
rect 3258 2931 3259 2932
rect 3263 2931 3264 2935
rect 3258 2930 3264 2931
rect 3379 2935 3385 2936
rect 3379 2931 3380 2935
rect 3384 2934 3385 2935
rect 3394 2935 3400 2936
rect 3394 2934 3395 2935
rect 3384 2932 3395 2934
rect 3384 2931 3385 2932
rect 3379 2930 3385 2931
rect 3394 2931 3395 2932
rect 3399 2931 3400 2935
rect 3394 2930 3400 2931
rect 3515 2935 3521 2936
rect 3515 2931 3516 2935
rect 3520 2934 3521 2935
rect 3554 2935 3560 2936
rect 3554 2934 3555 2935
rect 3520 2932 3555 2934
rect 3520 2931 3521 2932
rect 3515 2930 3521 2931
rect 3554 2931 3555 2932
rect 3559 2931 3560 2935
rect 3554 2930 3560 2931
rect 1762 2926 1769 2927
rect 1534 2922 1540 2923
rect 1387 2921 1490 2922
rect 1387 2917 1388 2921
rect 1392 2920 1490 2921
rect 1392 2917 1393 2920
rect 1387 2916 1393 2917
rect 1498 2919 1505 2920
rect 1498 2915 1499 2919
rect 1504 2915 1505 2919
rect 1498 2914 1505 2915
rect 1543 2919 1549 2920
rect 1543 2915 1544 2919
rect 1548 2918 1549 2919
rect 1611 2919 1617 2920
rect 1611 2918 1612 2919
rect 1548 2916 1612 2918
rect 1548 2915 1549 2916
rect 1543 2914 1549 2915
rect 1611 2915 1612 2916
rect 1616 2915 1617 2919
rect 1611 2914 1617 2915
rect 1710 2919 1716 2920
rect 1710 2915 1711 2919
rect 1715 2918 1716 2919
rect 1731 2919 1737 2920
rect 1731 2918 1732 2919
rect 1715 2916 1732 2918
rect 1715 2915 1716 2916
rect 1710 2914 1716 2915
rect 1731 2915 1732 2916
rect 1736 2915 1737 2919
rect 1731 2914 1737 2915
rect 1358 2909 1364 2910
rect 1358 2905 1359 2909
rect 1363 2905 1364 2909
rect 1358 2904 1364 2905
rect 1470 2909 1476 2910
rect 1470 2905 1471 2909
rect 1475 2905 1476 2909
rect 1470 2904 1476 2905
rect 1582 2909 1588 2910
rect 1582 2905 1583 2909
rect 1587 2905 1588 2909
rect 1582 2904 1588 2905
rect 1702 2909 1708 2910
rect 1702 2905 1703 2909
rect 1707 2905 1708 2909
rect 1702 2904 1708 2905
rect 2267 2907 2273 2908
rect 2267 2903 2268 2907
rect 2272 2906 2273 2907
rect 2306 2907 2312 2908
rect 2306 2906 2307 2907
rect 2272 2904 2307 2906
rect 2272 2903 2273 2904
rect 2267 2902 2273 2903
rect 2306 2903 2307 2904
rect 2311 2903 2312 2907
rect 2306 2902 2312 2903
rect 2394 2907 2400 2908
rect 2394 2903 2395 2907
rect 2399 2906 2400 2907
rect 2491 2907 2497 2908
rect 2491 2906 2492 2907
rect 2399 2904 2492 2906
rect 2399 2903 2400 2904
rect 2394 2902 2400 2903
rect 2491 2903 2492 2904
rect 2496 2903 2497 2907
rect 2491 2902 2497 2903
rect 2699 2907 2705 2908
rect 2699 2903 2700 2907
rect 2704 2906 2705 2907
rect 2750 2907 2756 2908
rect 2750 2906 2751 2907
rect 2704 2904 2751 2906
rect 2704 2903 2705 2904
rect 2699 2902 2705 2903
rect 2750 2903 2751 2904
rect 2755 2903 2756 2907
rect 2750 2902 2756 2903
rect 2759 2907 2765 2908
rect 2759 2903 2760 2907
rect 2764 2906 2765 2907
rect 2883 2907 2889 2908
rect 2883 2906 2884 2907
rect 2764 2904 2884 2906
rect 2764 2903 2765 2904
rect 2759 2902 2765 2903
rect 2883 2903 2884 2904
rect 2888 2903 2889 2907
rect 2883 2902 2889 2903
rect 2959 2907 2965 2908
rect 2959 2903 2960 2907
rect 2964 2906 2965 2907
rect 3051 2907 3057 2908
rect 3051 2906 3052 2907
rect 2964 2904 3052 2906
rect 2964 2903 2965 2904
rect 2959 2902 2965 2903
rect 3051 2903 3052 2904
rect 3056 2903 3057 2907
rect 3051 2902 3057 2903
rect 3119 2907 3125 2908
rect 3119 2903 3120 2907
rect 3124 2906 3125 2907
rect 3211 2907 3217 2908
rect 3211 2906 3212 2907
rect 3124 2904 3212 2906
rect 3124 2903 3125 2904
rect 3119 2902 3125 2903
rect 3211 2903 3212 2904
rect 3216 2903 3217 2907
rect 3211 2902 3217 2903
rect 3279 2907 3285 2908
rect 3279 2903 3280 2907
rect 3284 2906 3285 2907
rect 3363 2907 3369 2908
rect 3363 2906 3364 2907
rect 3284 2904 3364 2906
rect 3284 2903 3285 2904
rect 3279 2902 3285 2903
rect 3363 2903 3364 2904
rect 3368 2903 3369 2907
rect 3363 2902 3369 2903
rect 3515 2907 3521 2908
rect 3515 2903 3516 2907
rect 3520 2906 3521 2907
rect 3546 2907 3552 2908
rect 3546 2906 3547 2907
rect 3520 2904 3547 2906
rect 3520 2903 3521 2904
rect 3515 2902 3521 2903
rect 3546 2903 3547 2904
rect 3551 2903 3552 2907
rect 3546 2902 3552 2903
rect 2238 2897 2244 2898
rect 110 2896 116 2897
rect 1822 2896 1828 2897
rect 110 2892 111 2896
rect 115 2892 116 2896
rect 1543 2895 1549 2896
rect 1543 2894 1544 2895
rect 1525 2892 1544 2894
rect 110 2891 116 2892
rect 1543 2891 1544 2892
rect 1548 2891 1549 2895
rect 1762 2895 1768 2896
rect 1762 2894 1763 2895
rect 1757 2892 1763 2894
rect 1543 2890 1549 2891
rect 1762 2891 1763 2892
rect 1767 2891 1768 2895
rect 1822 2892 1823 2896
rect 1827 2892 1828 2896
rect 2238 2893 2239 2897
rect 2243 2893 2244 2897
rect 2238 2892 2244 2893
rect 2462 2897 2468 2898
rect 2462 2893 2463 2897
rect 2467 2893 2468 2897
rect 2462 2892 2468 2893
rect 2670 2897 2676 2898
rect 2670 2893 2671 2897
rect 2675 2893 2676 2897
rect 2670 2892 2676 2893
rect 2854 2897 2860 2898
rect 2854 2893 2855 2897
rect 2859 2893 2860 2897
rect 2854 2892 2860 2893
rect 3022 2897 3028 2898
rect 3022 2893 3023 2897
rect 3027 2893 3028 2897
rect 3022 2892 3028 2893
rect 3182 2897 3188 2898
rect 3182 2893 3183 2897
rect 3187 2893 3188 2897
rect 3182 2892 3188 2893
rect 3334 2897 3340 2898
rect 3334 2893 3335 2897
rect 3339 2893 3340 2897
rect 3334 2892 3340 2893
rect 3486 2897 3492 2898
rect 3486 2893 3487 2897
rect 3491 2893 3492 2897
rect 3486 2892 3492 2893
rect 1822 2891 1828 2892
rect 1762 2890 1768 2891
rect 1862 2884 1868 2885
rect 3574 2884 3580 2885
rect 1862 2880 1863 2884
rect 1867 2880 1868 2884
rect 2394 2883 2400 2884
rect 2394 2882 2395 2883
rect 2293 2880 2395 2882
rect 110 2879 116 2880
rect 110 2875 111 2879
rect 115 2875 116 2879
rect 110 2874 116 2875
rect 1538 2879 1544 2880
rect 1538 2875 1539 2879
rect 1543 2878 1544 2879
rect 1822 2879 1828 2880
rect 1862 2879 1868 2880
rect 2394 2879 2395 2880
rect 2399 2879 2400 2883
rect 2759 2883 2765 2884
rect 2759 2882 2760 2883
rect 2725 2880 2760 2882
rect 1543 2876 1593 2878
rect 1543 2875 1544 2876
rect 1538 2874 1544 2875
rect 1822 2875 1823 2879
rect 1827 2875 1828 2879
rect 2394 2878 2400 2879
rect 2759 2879 2760 2880
rect 2764 2879 2765 2883
rect 2959 2883 2965 2884
rect 2959 2882 2960 2883
rect 2909 2880 2960 2882
rect 2759 2878 2765 2879
rect 2959 2879 2960 2880
rect 2964 2879 2965 2883
rect 3119 2883 3125 2884
rect 3119 2882 3120 2883
rect 3077 2880 3120 2882
rect 2959 2878 2965 2879
rect 3119 2879 3120 2880
rect 3124 2879 3125 2883
rect 3279 2883 3285 2884
rect 3279 2882 3280 2883
rect 3237 2880 3280 2882
rect 3119 2878 3125 2879
rect 3279 2879 3280 2880
rect 3284 2879 3285 2883
rect 3394 2883 3400 2884
rect 3394 2882 3395 2883
rect 3389 2880 3395 2882
rect 3279 2878 3285 2879
rect 3394 2879 3395 2880
rect 3399 2879 3400 2883
rect 3574 2880 3575 2884
rect 3579 2880 3580 2884
rect 3574 2879 3580 2880
rect 3394 2878 3400 2879
rect 1822 2874 1828 2875
rect 1350 2869 1356 2870
rect 1350 2865 1351 2869
rect 1355 2865 1356 2869
rect 1350 2864 1356 2865
rect 1462 2869 1468 2870
rect 1462 2865 1463 2869
rect 1467 2865 1468 2869
rect 1462 2864 1468 2865
rect 1574 2869 1580 2870
rect 1574 2865 1575 2869
rect 1579 2865 1580 2869
rect 1574 2864 1580 2865
rect 1694 2869 1700 2870
rect 1694 2865 1695 2869
rect 1699 2865 1700 2869
rect 1694 2864 1700 2865
rect 1862 2867 1868 2868
rect 1399 2863 1405 2864
rect 1399 2859 1400 2863
rect 1404 2862 1405 2863
rect 1418 2863 1424 2864
rect 1418 2862 1419 2863
rect 1404 2860 1419 2862
rect 1404 2859 1405 2860
rect 1399 2858 1405 2859
rect 1418 2859 1419 2860
rect 1423 2859 1424 2863
rect 1862 2863 1863 2867
rect 1867 2863 1868 2867
rect 2546 2867 2552 2868
rect 2546 2866 2547 2867
rect 2513 2864 2547 2866
rect 1862 2862 1868 2863
rect 2546 2863 2547 2864
rect 2551 2863 2552 2867
rect 2546 2862 2552 2863
rect 3574 2867 3580 2868
rect 3574 2863 3575 2867
rect 3579 2863 3580 2867
rect 3574 2862 3580 2863
rect 1418 2858 1424 2859
rect 2230 2857 2236 2858
rect 2230 2853 2231 2857
rect 2235 2853 2236 2857
rect 2230 2852 2236 2853
rect 2454 2857 2460 2858
rect 2454 2853 2455 2857
rect 2459 2853 2460 2857
rect 2454 2852 2460 2853
rect 2662 2857 2668 2858
rect 2662 2853 2663 2857
rect 2667 2853 2668 2857
rect 2662 2852 2668 2853
rect 2846 2857 2852 2858
rect 2846 2853 2847 2857
rect 2851 2853 2852 2857
rect 2846 2852 2852 2853
rect 3014 2857 3020 2858
rect 3014 2853 3015 2857
rect 3019 2853 3020 2857
rect 3014 2852 3020 2853
rect 3174 2857 3180 2858
rect 3174 2853 3175 2857
rect 3179 2853 3180 2857
rect 3174 2852 3180 2853
rect 3326 2857 3332 2858
rect 3326 2853 3327 2857
rect 3331 2853 3332 2857
rect 3326 2852 3332 2853
rect 3478 2857 3484 2858
rect 3478 2853 3479 2857
rect 3483 2853 3484 2857
rect 3478 2852 3484 2853
rect 3518 2851 3524 2852
rect 3518 2847 3519 2851
rect 3523 2850 3524 2851
rect 3527 2851 3533 2852
rect 3527 2850 3528 2851
rect 3523 2848 3528 2850
rect 3523 2847 3524 2848
rect 3518 2846 3524 2847
rect 3527 2847 3528 2848
rect 3532 2847 3533 2851
rect 3527 2846 3533 2847
rect 134 2843 140 2844
rect 134 2839 135 2843
rect 139 2839 140 2843
rect 134 2838 140 2839
rect 222 2843 228 2844
rect 222 2839 223 2843
rect 227 2839 228 2843
rect 222 2838 228 2839
rect 310 2843 316 2844
rect 310 2839 311 2843
rect 315 2839 316 2843
rect 310 2838 316 2839
rect 398 2843 404 2844
rect 398 2839 399 2843
rect 403 2839 404 2843
rect 398 2838 404 2839
rect 486 2843 492 2844
rect 486 2839 487 2843
rect 491 2839 492 2843
rect 486 2838 492 2839
rect 598 2843 604 2844
rect 598 2839 599 2843
rect 603 2839 604 2843
rect 598 2838 604 2839
rect 726 2843 732 2844
rect 726 2839 727 2843
rect 731 2839 732 2843
rect 726 2838 732 2839
rect 862 2843 868 2844
rect 862 2839 863 2843
rect 867 2839 868 2843
rect 862 2838 868 2839
rect 998 2843 1004 2844
rect 998 2839 999 2843
rect 1003 2839 1004 2843
rect 998 2838 1004 2839
rect 1134 2843 1140 2844
rect 1134 2839 1135 2843
rect 1139 2839 1140 2843
rect 1134 2838 1140 2839
rect 1262 2843 1268 2844
rect 1262 2839 1263 2843
rect 1267 2839 1268 2843
rect 1262 2838 1268 2839
rect 1382 2843 1388 2844
rect 1382 2839 1383 2843
rect 1387 2839 1388 2843
rect 1382 2838 1388 2839
rect 1502 2843 1508 2844
rect 1502 2839 1503 2843
rect 1507 2839 1508 2843
rect 1502 2838 1508 2839
rect 1622 2843 1628 2844
rect 1622 2839 1623 2843
rect 1627 2839 1628 2843
rect 1622 2838 1628 2839
rect 1726 2843 1732 2844
rect 1726 2839 1727 2843
rect 1731 2839 1732 2843
rect 1726 2838 1732 2839
rect 930 2835 936 2836
rect 110 2833 116 2834
rect 110 2829 111 2833
rect 115 2829 116 2833
rect 930 2831 931 2835
rect 935 2834 936 2835
rect 1710 2835 1716 2836
rect 1710 2834 1711 2835
rect 935 2832 1017 2834
rect 1681 2832 1711 2834
rect 935 2831 936 2832
rect 930 2830 936 2831
rect 1710 2831 1711 2832
rect 1715 2831 1716 2835
rect 1710 2830 1716 2831
rect 1822 2833 1828 2834
rect 110 2828 116 2829
rect 1822 2829 1823 2833
rect 1827 2829 1828 2833
rect 1822 2828 1828 2829
rect 1894 2831 1900 2832
rect 1894 2827 1895 2831
rect 1899 2827 1900 2831
rect 1894 2826 1900 2827
rect 1982 2831 1988 2832
rect 1982 2827 1983 2831
rect 1987 2827 1988 2831
rect 1982 2826 1988 2827
rect 2070 2831 2076 2832
rect 2070 2827 2071 2831
rect 2075 2827 2076 2831
rect 2070 2826 2076 2827
rect 2158 2831 2164 2832
rect 2158 2827 2159 2831
rect 2163 2827 2164 2831
rect 2158 2826 2164 2827
rect 2246 2831 2252 2832
rect 2246 2827 2247 2831
rect 2251 2827 2252 2831
rect 2246 2826 2252 2827
rect 2334 2831 2340 2832
rect 2334 2827 2335 2831
rect 2339 2827 2340 2831
rect 2334 2826 2340 2827
rect 2422 2831 2428 2832
rect 2422 2827 2423 2831
rect 2427 2827 2428 2831
rect 2422 2826 2428 2827
rect 2510 2831 2516 2832
rect 2510 2827 2511 2831
rect 2515 2827 2516 2831
rect 2510 2826 2516 2827
rect 2598 2831 2604 2832
rect 2598 2827 2599 2831
rect 2603 2827 2604 2831
rect 2598 2826 2604 2827
rect 2686 2831 2692 2832
rect 2686 2827 2687 2831
rect 2691 2827 2692 2831
rect 2686 2826 2692 2827
rect 2790 2831 2796 2832
rect 2790 2827 2791 2831
rect 2795 2827 2796 2831
rect 2790 2826 2796 2827
rect 2902 2831 2908 2832
rect 2902 2827 2903 2831
rect 2907 2827 2908 2831
rect 2902 2826 2908 2827
rect 3030 2831 3036 2832
rect 3030 2827 3031 2831
rect 3035 2827 3036 2831
rect 3030 2826 3036 2827
rect 3174 2831 3180 2832
rect 3174 2827 3175 2831
rect 3179 2827 3180 2831
rect 3174 2826 3180 2827
rect 3326 2831 3332 2832
rect 3326 2827 3327 2831
rect 3331 2827 3332 2831
rect 3326 2826 3332 2827
rect 3478 2831 3484 2832
rect 3478 2827 3479 2831
rect 3483 2827 3484 2831
rect 3478 2826 3484 2827
rect 2498 2823 2504 2824
rect 2498 2822 2499 2823
rect 1862 2821 1868 2822
rect 202 2819 208 2820
rect 110 2816 116 2817
rect 110 2812 111 2816
rect 115 2812 116 2816
rect 110 2811 116 2812
rect 196 2810 198 2817
rect 202 2815 203 2819
rect 207 2818 208 2819
rect 295 2819 301 2820
rect 207 2816 249 2818
rect 207 2815 208 2816
rect 202 2814 208 2815
rect 295 2815 296 2819
rect 300 2818 301 2819
rect 378 2819 384 2820
rect 300 2816 337 2818
rect 300 2815 301 2816
rect 295 2814 301 2815
rect 378 2815 379 2819
rect 383 2818 384 2819
rect 466 2819 472 2820
rect 383 2816 425 2818
rect 383 2815 384 2816
rect 378 2814 384 2815
rect 466 2815 467 2819
rect 471 2818 472 2819
rect 558 2819 564 2820
rect 471 2816 513 2818
rect 471 2815 472 2816
rect 466 2814 472 2815
rect 558 2815 559 2819
rect 563 2818 564 2819
rect 666 2819 672 2820
rect 563 2816 625 2818
rect 563 2815 564 2816
rect 558 2814 564 2815
rect 666 2815 667 2819
rect 671 2818 672 2819
rect 959 2819 965 2820
rect 959 2818 960 2819
rect 671 2816 753 2818
rect 925 2816 960 2818
rect 671 2815 672 2816
rect 666 2814 672 2815
rect 959 2815 960 2816
rect 964 2815 965 2819
rect 959 2814 965 2815
rect 1066 2819 1072 2820
rect 1066 2815 1067 2819
rect 1071 2818 1072 2819
rect 1207 2819 1213 2820
rect 1071 2816 1161 2818
rect 1071 2815 1072 2816
rect 1066 2814 1072 2815
rect 1207 2815 1208 2819
rect 1212 2818 1213 2819
rect 1330 2819 1336 2820
rect 1212 2816 1289 2818
rect 1212 2815 1213 2816
rect 1207 2814 1213 2815
rect 1330 2815 1331 2819
rect 1335 2818 1336 2819
rect 1578 2819 1584 2820
rect 1578 2818 1579 2819
rect 1335 2816 1409 2818
rect 1565 2816 1579 2818
rect 1335 2815 1336 2816
rect 1330 2814 1336 2815
rect 1578 2815 1579 2816
rect 1583 2815 1584 2819
rect 1578 2814 1584 2815
rect 1690 2819 1696 2820
rect 1690 2815 1691 2819
rect 1695 2818 1696 2819
rect 1695 2816 1753 2818
rect 1862 2817 1863 2821
rect 1867 2817 1868 2821
rect 2481 2820 2499 2822
rect 2498 2819 2499 2820
rect 2503 2819 2504 2823
rect 2498 2818 2504 2819
rect 3098 2823 3104 2824
rect 3098 2819 3099 2823
rect 3103 2822 3104 2823
rect 3103 2820 3193 2822
rect 3574 2821 3580 2822
rect 3103 2819 3104 2820
rect 3098 2818 3104 2819
rect 1822 2816 1828 2817
rect 1862 2816 1868 2817
rect 3574 2817 3575 2821
rect 3579 2817 3580 2821
rect 3574 2816 3580 2817
rect 1695 2815 1696 2816
rect 1690 2814 1696 2815
rect 1822 2812 1823 2816
rect 1827 2812 1828 2816
rect 207 2811 213 2812
rect 1822 2811 1828 2812
rect 207 2810 208 2811
rect 196 2808 208 2810
rect 207 2807 208 2808
rect 212 2807 213 2811
rect 207 2806 213 2807
rect 1975 2807 1981 2808
rect 1975 2806 1976 2807
rect 1862 2804 1868 2805
rect 1957 2804 1976 2806
rect 142 2803 148 2804
rect 142 2799 143 2803
rect 147 2799 148 2803
rect 142 2798 148 2799
rect 230 2803 236 2804
rect 230 2799 231 2803
rect 235 2799 236 2803
rect 230 2798 236 2799
rect 318 2803 324 2804
rect 318 2799 319 2803
rect 323 2799 324 2803
rect 318 2798 324 2799
rect 406 2803 412 2804
rect 406 2799 407 2803
rect 411 2799 412 2803
rect 406 2798 412 2799
rect 494 2803 500 2804
rect 494 2799 495 2803
rect 499 2799 500 2803
rect 494 2798 500 2799
rect 606 2803 612 2804
rect 606 2799 607 2803
rect 611 2799 612 2803
rect 606 2798 612 2799
rect 734 2803 740 2804
rect 734 2799 735 2803
rect 739 2799 740 2803
rect 734 2798 740 2799
rect 870 2803 876 2804
rect 870 2799 871 2803
rect 875 2799 876 2803
rect 1006 2803 1012 2804
rect 870 2798 876 2799
rect 930 2799 936 2800
rect 930 2798 931 2799
rect 880 2796 931 2798
rect 880 2794 882 2796
rect 930 2795 931 2796
rect 935 2795 936 2799
rect 1006 2799 1007 2803
rect 1011 2799 1012 2803
rect 1006 2798 1012 2799
rect 1142 2803 1148 2804
rect 1142 2799 1143 2803
rect 1147 2799 1148 2803
rect 1142 2798 1148 2799
rect 1270 2803 1276 2804
rect 1270 2799 1271 2803
rect 1275 2799 1276 2803
rect 1270 2798 1276 2799
rect 1390 2803 1396 2804
rect 1390 2799 1391 2803
rect 1395 2799 1396 2803
rect 1390 2798 1396 2799
rect 1510 2803 1516 2804
rect 1510 2799 1511 2803
rect 1515 2799 1516 2803
rect 1510 2798 1516 2799
rect 1630 2803 1636 2804
rect 1630 2799 1631 2803
rect 1635 2799 1636 2803
rect 1734 2803 1740 2804
rect 1630 2798 1636 2799
rect 1690 2799 1696 2800
rect 1690 2798 1691 2799
rect 930 2794 936 2795
rect 1540 2796 1590 2798
rect 1540 2794 1542 2796
rect 1588 2794 1590 2796
rect 1640 2796 1691 2798
rect 1640 2794 1642 2796
rect 1690 2795 1691 2796
rect 1695 2795 1696 2799
rect 1734 2799 1735 2803
rect 1739 2799 1740 2803
rect 1862 2800 1863 2804
rect 1867 2800 1868 2804
rect 1975 2803 1976 2804
rect 1980 2803 1981 2807
rect 2063 2807 2069 2808
rect 2063 2806 2064 2807
rect 2045 2804 2064 2806
rect 1975 2802 1981 2803
rect 2063 2803 2064 2804
rect 2068 2803 2069 2807
rect 2151 2807 2157 2808
rect 2151 2806 2152 2807
rect 2133 2804 2152 2806
rect 2063 2802 2069 2803
rect 2151 2803 2152 2804
rect 2156 2803 2157 2807
rect 2239 2807 2245 2808
rect 2239 2806 2240 2807
rect 2221 2804 2240 2806
rect 2151 2802 2157 2803
rect 2239 2803 2240 2804
rect 2244 2803 2245 2807
rect 2327 2807 2333 2808
rect 2327 2806 2328 2807
rect 2309 2804 2328 2806
rect 2239 2802 2245 2803
rect 2327 2803 2328 2804
rect 2332 2803 2333 2807
rect 2415 2807 2421 2808
rect 2415 2806 2416 2807
rect 2397 2804 2416 2806
rect 2327 2802 2333 2803
rect 2415 2803 2416 2804
rect 2420 2803 2421 2807
rect 2415 2802 2421 2803
rect 2490 2807 2496 2808
rect 2490 2803 2491 2807
rect 2495 2806 2496 2807
rect 2679 2807 2685 2808
rect 2679 2806 2680 2807
rect 2495 2804 2537 2806
rect 2661 2804 2680 2806
rect 2495 2803 2496 2804
rect 2490 2802 2496 2803
rect 2679 2803 2680 2804
rect 2684 2803 2685 2807
rect 2783 2807 2789 2808
rect 2783 2806 2784 2807
rect 2749 2804 2784 2806
rect 2679 2802 2685 2803
rect 2783 2803 2784 2804
rect 2788 2803 2789 2807
rect 2895 2807 2901 2808
rect 2895 2806 2896 2807
rect 2853 2804 2896 2806
rect 2783 2802 2789 2803
rect 2895 2803 2896 2804
rect 2900 2803 2901 2807
rect 3023 2807 3029 2808
rect 3023 2806 3024 2807
rect 2965 2804 3024 2806
rect 2895 2802 2901 2803
rect 3023 2803 3024 2804
rect 3028 2803 3029 2807
rect 3098 2807 3104 2808
rect 3098 2806 3099 2807
rect 3093 2804 3099 2806
rect 3023 2802 3029 2803
rect 3098 2803 3099 2804
rect 3103 2803 3104 2807
rect 3098 2802 3104 2803
rect 3242 2807 3248 2808
rect 3242 2803 3243 2807
rect 3247 2806 3248 2807
rect 3546 2807 3552 2808
rect 3546 2806 3547 2807
rect 3247 2804 3353 2806
rect 3541 2804 3547 2806
rect 3247 2803 3248 2804
rect 3242 2802 3248 2803
rect 3546 2803 3547 2804
rect 3551 2803 3552 2807
rect 3546 2802 3552 2803
rect 3574 2804 3580 2805
rect 1862 2799 1868 2800
rect 3574 2800 3575 2804
rect 3579 2800 3580 2804
rect 3574 2799 3580 2800
rect 1734 2798 1740 2799
rect 1690 2794 1696 2795
rect 763 2793 882 2794
rect 171 2791 177 2792
rect 171 2787 172 2791
rect 176 2790 177 2791
rect 202 2791 208 2792
rect 202 2790 203 2791
rect 176 2788 203 2790
rect 176 2787 177 2788
rect 171 2786 177 2787
rect 202 2787 203 2788
rect 207 2787 208 2791
rect 202 2786 208 2787
rect 259 2791 265 2792
rect 259 2787 260 2791
rect 264 2790 265 2791
rect 295 2791 301 2792
rect 295 2790 296 2791
rect 264 2788 296 2790
rect 264 2787 265 2788
rect 259 2786 265 2787
rect 295 2787 296 2788
rect 300 2787 301 2791
rect 295 2786 301 2787
rect 347 2791 353 2792
rect 347 2787 348 2791
rect 352 2790 353 2791
rect 378 2791 384 2792
rect 378 2790 379 2791
rect 352 2788 379 2790
rect 352 2787 353 2788
rect 347 2786 353 2787
rect 378 2787 379 2788
rect 383 2787 384 2791
rect 378 2786 384 2787
rect 435 2791 441 2792
rect 435 2787 436 2791
rect 440 2790 441 2791
rect 466 2791 472 2792
rect 466 2790 467 2791
rect 440 2788 467 2790
rect 440 2787 441 2788
rect 435 2786 441 2787
rect 466 2787 467 2788
rect 471 2787 472 2791
rect 466 2786 472 2787
rect 523 2791 529 2792
rect 523 2787 524 2791
rect 528 2790 529 2791
rect 558 2791 564 2792
rect 558 2790 559 2791
rect 528 2788 559 2790
rect 528 2787 529 2788
rect 523 2786 529 2787
rect 558 2787 559 2788
rect 563 2787 564 2791
rect 558 2786 564 2787
rect 635 2791 641 2792
rect 635 2787 636 2791
rect 640 2790 641 2791
rect 666 2791 672 2792
rect 666 2790 667 2791
rect 640 2788 667 2790
rect 640 2787 641 2788
rect 635 2786 641 2787
rect 666 2787 667 2788
rect 671 2787 672 2791
rect 763 2789 764 2793
rect 768 2792 882 2793
rect 1539 2793 1545 2794
rect 768 2789 769 2792
rect 763 2788 769 2789
rect 887 2791 893 2792
rect 666 2786 672 2787
rect 887 2787 888 2791
rect 892 2790 893 2791
rect 899 2791 905 2792
rect 899 2790 900 2791
rect 892 2788 900 2790
rect 892 2787 893 2788
rect 887 2786 893 2787
rect 899 2787 900 2788
rect 904 2787 905 2791
rect 899 2786 905 2787
rect 959 2791 965 2792
rect 959 2787 960 2791
rect 964 2790 965 2791
rect 1035 2791 1041 2792
rect 1035 2790 1036 2791
rect 964 2788 1036 2790
rect 964 2787 965 2788
rect 959 2786 965 2787
rect 1035 2787 1036 2788
rect 1040 2787 1041 2791
rect 1035 2786 1041 2787
rect 1171 2791 1177 2792
rect 1171 2787 1172 2791
rect 1176 2790 1177 2791
rect 1207 2791 1213 2792
rect 1207 2790 1208 2791
rect 1176 2788 1208 2790
rect 1176 2787 1177 2788
rect 1171 2786 1177 2787
rect 1207 2787 1208 2788
rect 1212 2787 1213 2791
rect 1207 2786 1213 2787
rect 1299 2791 1305 2792
rect 1299 2787 1300 2791
rect 1304 2790 1305 2791
rect 1330 2791 1336 2792
rect 1330 2790 1331 2791
rect 1304 2788 1331 2790
rect 1304 2787 1305 2788
rect 1299 2786 1305 2787
rect 1330 2787 1331 2788
rect 1335 2787 1336 2791
rect 1330 2786 1336 2787
rect 1418 2791 1425 2792
rect 1418 2787 1419 2791
rect 1424 2787 1425 2791
rect 1539 2789 1540 2793
rect 1544 2789 1545 2793
rect 1588 2792 1642 2794
rect 1539 2788 1545 2789
rect 1578 2791 1584 2792
rect 1418 2786 1425 2787
rect 1578 2787 1579 2791
rect 1583 2790 1584 2791
rect 1659 2791 1665 2792
rect 1659 2790 1660 2791
rect 1583 2788 1660 2790
rect 1583 2787 1584 2788
rect 1578 2786 1584 2787
rect 1659 2787 1660 2788
rect 1664 2787 1665 2791
rect 1659 2786 1665 2787
rect 1763 2791 1769 2792
rect 1763 2787 1764 2791
rect 1768 2790 1769 2791
rect 1794 2791 1800 2792
rect 1794 2790 1795 2791
rect 1768 2788 1795 2790
rect 1768 2787 1769 2788
rect 1763 2786 1769 2787
rect 1794 2787 1795 2788
rect 1799 2787 1800 2791
rect 1794 2786 1800 2787
rect 1902 2791 1908 2792
rect 1902 2787 1903 2791
rect 1907 2787 1908 2791
rect 1902 2786 1908 2787
rect 1990 2791 1996 2792
rect 1990 2787 1991 2791
rect 1995 2787 1996 2791
rect 1990 2786 1996 2787
rect 2078 2791 2084 2792
rect 2078 2787 2079 2791
rect 2083 2787 2084 2791
rect 2078 2786 2084 2787
rect 2166 2791 2172 2792
rect 2166 2787 2167 2791
rect 2171 2787 2172 2791
rect 2166 2786 2172 2787
rect 2254 2791 2260 2792
rect 2254 2787 2255 2791
rect 2259 2787 2260 2791
rect 2254 2786 2260 2787
rect 2342 2791 2348 2792
rect 2342 2787 2343 2791
rect 2347 2787 2348 2791
rect 2342 2786 2348 2787
rect 2430 2791 2436 2792
rect 2430 2787 2431 2791
rect 2435 2787 2436 2791
rect 2430 2786 2436 2787
rect 2518 2791 2524 2792
rect 2518 2787 2519 2791
rect 2523 2787 2524 2791
rect 2518 2786 2524 2787
rect 2606 2791 2612 2792
rect 2606 2787 2607 2791
rect 2611 2787 2612 2791
rect 2606 2786 2612 2787
rect 2694 2791 2700 2792
rect 2694 2787 2695 2791
rect 2699 2787 2700 2791
rect 2694 2786 2700 2787
rect 2798 2791 2804 2792
rect 2798 2787 2799 2791
rect 2803 2787 2804 2791
rect 2798 2786 2804 2787
rect 2910 2791 2916 2792
rect 2910 2787 2911 2791
rect 2915 2787 2916 2791
rect 2910 2786 2916 2787
rect 3038 2791 3044 2792
rect 3038 2787 3039 2791
rect 3043 2787 3044 2791
rect 3038 2786 3044 2787
rect 3182 2791 3188 2792
rect 3182 2787 3183 2791
rect 3187 2787 3188 2791
rect 3182 2786 3188 2787
rect 3334 2791 3340 2792
rect 3334 2787 3335 2791
rect 3339 2787 3340 2791
rect 3334 2786 3340 2787
rect 3486 2791 3492 2792
rect 3486 2787 3487 2791
rect 3491 2787 3492 2791
rect 3486 2786 3492 2787
rect 207 2779 213 2780
rect 207 2775 208 2779
rect 212 2778 213 2779
rect 219 2779 225 2780
rect 219 2778 220 2779
rect 212 2776 220 2778
rect 212 2775 213 2776
rect 207 2774 213 2775
rect 219 2775 220 2776
rect 224 2775 225 2779
rect 219 2774 225 2775
rect 279 2779 285 2780
rect 279 2775 280 2779
rect 284 2778 285 2779
rect 323 2779 329 2780
rect 323 2778 324 2779
rect 284 2776 324 2778
rect 284 2775 285 2776
rect 279 2774 285 2775
rect 323 2775 324 2776
rect 328 2775 329 2779
rect 323 2774 329 2775
rect 375 2779 381 2780
rect 375 2775 376 2779
rect 380 2778 381 2779
rect 443 2779 449 2780
rect 443 2778 444 2779
rect 380 2776 444 2778
rect 380 2775 381 2776
rect 375 2774 381 2775
rect 443 2775 444 2776
rect 448 2775 449 2779
rect 443 2774 449 2775
rect 570 2779 576 2780
rect 570 2775 571 2779
rect 575 2778 576 2779
rect 579 2779 585 2780
rect 579 2778 580 2779
rect 575 2776 580 2778
rect 575 2775 576 2776
rect 570 2774 576 2775
rect 579 2775 580 2776
rect 584 2775 585 2779
rect 579 2774 585 2775
rect 639 2779 645 2780
rect 639 2775 640 2779
rect 644 2778 645 2779
rect 715 2779 721 2780
rect 715 2778 716 2779
rect 644 2776 716 2778
rect 644 2775 645 2776
rect 639 2774 645 2775
rect 715 2775 716 2776
rect 720 2775 721 2779
rect 715 2774 721 2775
rect 775 2779 781 2780
rect 775 2775 776 2779
rect 780 2778 781 2779
rect 851 2779 857 2780
rect 851 2778 852 2779
rect 780 2776 852 2778
rect 780 2775 781 2776
rect 775 2774 781 2775
rect 851 2775 852 2776
rect 856 2775 857 2779
rect 851 2774 857 2775
rect 987 2779 993 2780
rect 987 2775 988 2779
rect 992 2778 993 2779
rect 1031 2779 1037 2780
rect 992 2776 1026 2778
rect 992 2775 993 2776
rect 987 2774 993 2775
rect 1024 2770 1026 2776
rect 1031 2775 1032 2779
rect 1036 2778 1037 2779
rect 1115 2779 1121 2780
rect 1115 2778 1116 2779
rect 1036 2776 1116 2778
rect 1036 2775 1037 2776
rect 1031 2774 1037 2775
rect 1115 2775 1116 2776
rect 1120 2775 1121 2779
rect 1115 2774 1121 2775
rect 1190 2779 1196 2780
rect 1190 2775 1191 2779
rect 1195 2778 1196 2779
rect 1235 2779 1241 2780
rect 1235 2778 1236 2779
rect 1195 2776 1236 2778
rect 1195 2775 1196 2776
rect 1190 2774 1196 2775
rect 1235 2775 1236 2776
rect 1240 2775 1241 2779
rect 1235 2774 1241 2775
rect 1279 2779 1285 2780
rect 1279 2775 1280 2779
rect 1284 2778 1285 2779
rect 1347 2779 1353 2780
rect 1347 2778 1348 2779
rect 1284 2776 1348 2778
rect 1284 2775 1285 2776
rect 1279 2774 1285 2775
rect 1347 2775 1348 2776
rect 1352 2775 1353 2779
rect 1347 2774 1353 2775
rect 1391 2779 1397 2780
rect 1391 2775 1392 2779
rect 1396 2778 1397 2779
rect 1459 2779 1465 2780
rect 1459 2778 1460 2779
rect 1396 2776 1460 2778
rect 1396 2775 1397 2776
rect 1391 2774 1397 2775
rect 1459 2775 1460 2776
rect 1464 2775 1465 2779
rect 1459 2774 1465 2775
rect 1503 2779 1509 2780
rect 1503 2775 1504 2779
rect 1508 2778 1509 2779
rect 1563 2779 1569 2780
rect 1563 2778 1564 2779
rect 1508 2776 1564 2778
rect 1508 2775 1509 2776
rect 1503 2774 1509 2775
rect 1563 2775 1564 2776
rect 1568 2775 1569 2779
rect 1563 2774 1569 2775
rect 1607 2779 1613 2780
rect 1607 2775 1608 2779
rect 1612 2778 1613 2779
rect 1675 2779 1681 2780
rect 1675 2778 1676 2779
rect 1612 2776 1676 2778
rect 1612 2775 1613 2776
rect 1607 2774 1613 2775
rect 1675 2775 1676 2776
rect 1680 2775 1681 2779
rect 1675 2774 1681 2775
rect 1711 2779 1717 2780
rect 1711 2775 1712 2779
rect 1716 2778 1717 2779
rect 1763 2779 1769 2780
rect 1763 2778 1764 2779
rect 1716 2776 1764 2778
rect 1716 2775 1717 2776
rect 1711 2774 1717 2775
rect 1763 2775 1764 2776
rect 1768 2775 1769 2779
rect 1763 2774 1769 2775
rect 1931 2779 1937 2780
rect 1931 2775 1932 2779
rect 1936 2778 1937 2779
rect 1975 2779 1981 2780
rect 1936 2776 1970 2778
rect 1936 2775 1937 2776
rect 1931 2774 1937 2775
rect 1066 2771 1072 2772
rect 1066 2770 1067 2771
rect 190 2769 196 2770
rect 190 2765 191 2769
rect 195 2765 196 2769
rect 190 2764 196 2765
rect 294 2769 300 2770
rect 294 2765 295 2769
rect 299 2765 300 2769
rect 294 2764 300 2765
rect 414 2769 420 2770
rect 414 2765 415 2769
rect 419 2765 420 2769
rect 414 2764 420 2765
rect 550 2769 556 2770
rect 550 2765 551 2769
rect 555 2765 556 2769
rect 550 2764 556 2765
rect 686 2769 692 2770
rect 686 2765 687 2769
rect 691 2765 692 2769
rect 686 2764 692 2765
rect 822 2769 828 2770
rect 822 2765 823 2769
rect 827 2765 828 2769
rect 822 2764 828 2765
rect 958 2769 964 2770
rect 958 2765 959 2769
rect 963 2765 964 2769
rect 1024 2768 1067 2770
rect 1066 2767 1067 2768
rect 1071 2767 1072 2771
rect 1968 2770 1970 2776
rect 1975 2775 1976 2779
rect 1980 2778 1981 2779
rect 2019 2779 2025 2780
rect 2019 2778 2020 2779
rect 1980 2776 2020 2778
rect 1980 2775 1981 2776
rect 1975 2774 1981 2775
rect 2019 2775 2020 2776
rect 2024 2775 2025 2779
rect 2019 2774 2025 2775
rect 2063 2779 2069 2780
rect 2063 2775 2064 2779
rect 2068 2778 2069 2779
rect 2107 2779 2113 2780
rect 2107 2778 2108 2779
rect 2068 2776 2108 2778
rect 2068 2775 2069 2776
rect 2063 2774 2069 2775
rect 2107 2775 2108 2776
rect 2112 2775 2113 2779
rect 2107 2774 2113 2775
rect 2151 2779 2157 2780
rect 2151 2775 2152 2779
rect 2156 2778 2157 2779
rect 2195 2779 2201 2780
rect 2195 2778 2196 2779
rect 2156 2776 2196 2778
rect 2156 2775 2157 2776
rect 2151 2774 2157 2775
rect 2195 2775 2196 2776
rect 2200 2775 2201 2779
rect 2195 2774 2201 2775
rect 2239 2779 2245 2780
rect 2239 2775 2240 2779
rect 2244 2778 2245 2779
rect 2283 2779 2289 2780
rect 2283 2778 2284 2779
rect 2244 2776 2284 2778
rect 2244 2775 2245 2776
rect 2239 2774 2245 2775
rect 2283 2775 2284 2776
rect 2288 2775 2289 2779
rect 2283 2774 2289 2775
rect 2327 2779 2333 2780
rect 2327 2775 2328 2779
rect 2332 2778 2333 2779
rect 2371 2779 2377 2780
rect 2371 2778 2372 2779
rect 2332 2776 2372 2778
rect 2332 2775 2333 2776
rect 2327 2774 2333 2775
rect 2371 2775 2372 2776
rect 2376 2775 2377 2779
rect 2371 2774 2377 2775
rect 2459 2779 2465 2780
rect 2459 2775 2460 2779
rect 2464 2778 2465 2779
rect 2490 2779 2496 2780
rect 2490 2778 2491 2779
rect 2464 2776 2491 2778
rect 2464 2775 2465 2776
rect 2459 2774 2465 2775
rect 2490 2775 2491 2776
rect 2495 2775 2496 2779
rect 2490 2774 2496 2775
rect 2546 2779 2553 2780
rect 2546 2775 2547 2779
rect 2552 2775 2553 2779
rect 2635 2779 2641 2780
rect 2635 2778 2636 2779
rect 2546 2774 2553 2775
rect 2556 2776 2636 2778
rect 2247 2771 2253 2772
rect 2247 2770 2248 2771
rect 1066 2766 1072 2767
rect 1086 2769 1092 2770
rect 958 2764 964 2765
rect 1086 2765 1087 2769
rect 1091 2765 1092 2769
rect 1086 2764 1092 2765
rect 1206 2769 1212 2770
rect 1206 2765 1207 2769
rect 1211 2765 1212 2769
rect 1206 2764 1212 2765
rect 1318 2769 1324 2770
rect 1318 2765 1319 2769
rect 1323 2765 1324 2769
rect 1318 2764 1324 2765
rect 1430 2769 1436 2770
rect 1430 2765 1431 2769
rect 1435 2765 1436 2769
rect 1430 2764 1436 2765
rect 1534 2769 1540 2770
rect 1534 2765 1535 2769
rect 1539 2765 1540 2769
rect 1534 2764 1540 2765
rect 1646 2769 1652 2770
rect 1646 2765 1647 2769
rect 1651 2765 1652 2769
rect 1646 2764 1652 2765
rect 1734 2769 1740 2770
rect 1734 2765 1735 2769
rect 1739 2765 1740 2769
rect 1968 2768 2248 2770
rect 2247 2767 2248 2768
rect 2252 2767 2253 2771
rect 2247 2766 2253 2767
rect 2415 2771 2421 2772
rect 2415 2767 2416 2771
rect 2420 2770 2421 2771
rect 2556 2770 2558 2776
rect 2635 2775 2636 2776
rect 2640 2775 2641 2779
rect 2635 2774 2641 2775
rect 2679 2779 2685 2780
rect 2679 2775 2680 2779
rect 2684 2778 2685 2779
rect 2723 2779 2729 2780
rect 2723 2778 2724 2779
rect 2684 2776 2724 2778
rect 2684 2775 2685 2776
rect 2679 2774 2685 2775
rect 2723 2775 2724 2776
rect 2728 2775 2729 2779
rect 2723 2774 2729 2775
rect 2783 2779 2789 2780
rect 2783 2775 2784 2779
rect 2788 2778 2789 2779
rect 2827 2779 2833 2780
rect 2827 2778 2828 2779
rect 2788 2776 2828 2778
rect 2788 2775 2789 2776
rect 2783 2774 2789 2775
rect 2827 2775 2828 2776
rect 2832 2775 2833 2779
rect 2827 2774 2833 2775
rect 2895 2779 2901 2780
rect 2895 2775 2896 2779
rect 2900 2778 2901 2779
rect 2939 2779 2945 2780
rect 2939 2778 2940 2779
rect 2900 2776 2940 2778
rect 2900 2775 2901 2776
rect 2895 2774 2901 2775
rect 2939 2775 2940 2776
rect 2944 2775 2945 2779
rect 2939 2774 2945 2775
rect 3023 2779 3029 2780
rect 3023 2775 3024 2779
rect 3028 2778 3029 2779
rect 3067 2779 3073 2780
rect 3067 2778 3068 2779
rect 3028 2776 3068 2778
rect 3028 2775 3029 2776
rect 3023 2774 3029 2775
rect 3067 2775 3068 2776
rect 3072 2775 3073 2779
rect 3067 2774 3073 2775
rect 3211 2779 3217 2780
rect 3211 2775 3212 2779
rect 3216 2778 3217 2779
rect 3242 2779 3248 2780
rect 3242 2778 3243 2779
rect 3216 2776 3243 2778
rect 3216 2775 3217 2776
rect 3211 2774 3217 2775
rect 3242 2775 3243 2776
rect 3247 2775 3248 2779
rect 3242 2774 3248 2775
rect 3335 2779 3341 2780
rect 3335 2775 3336 2779
rect 3340 2778 3341 2779
rect 3363 2779 3369 2780
rect 3363 2778 3364 2779
rect 3340 2776 3364 2778
rect 3340 2775 3341 2776
rect 3335 2774 3341 2775
rect 3363 2775 3364 2776
rect 3368 2775 3369 2779
rect 3363 2774 3369 2775
rect 3515 2779 3524 2780
rect 3515 2775 3516 2779
rect 3523 2775 3524 2779
rect 3515 2774 3524 2775
rect 2420 2768 2558 2770
rect 2420 2767 2421 2768
rect 2415 2766 2421 2767
rect 1734 2764 1740 2765
rect 110 2756 116 2757
rect 1822 2756 1828 2757
rect 110 2752 111 2756
rect 115 2752 116 2756
rect 279 2755 285 2756
rect 279 2754 280 2755
rect 245 2752 280 2754
rect 110 2751 116 2752
rect 279 2751 280 2752
rect 284 2751 285 2755
rect 375 2755 381 2756
rect 375 2754 376 2755
rect 349 2752 376 2754
rect 279 2750 285 2751
rect 375 2751 376 2752
rect 380 2751 381 2755
rect 639 2755 645 2756
rect 639 2754 640 2755
rect 605 2752 640 2754
rect 375 2750 381 2751
rect 639 2751 640 2752
rect 644 2751 645 2755
rect 775 2755 781 2756
rect 775 2754 776 2755
rect 741 2752 776 2754
rect 639 2750 645 2751
rect 775 2751 776 2752
rect 780 2751 781 2755
rect 887 2755 893 2756
rect 887 2754 888 2755
rect 877 2752 888 2754
rect 775 2750 781 2751
rect 887 2751 888 2752
rect 892 2751 893 2755
rect 1031 2755 1037 2756
rect 1031 2754 1032 2755
rect 1013 2752 1032 2754
rect 887 2750 893 2751
rect 1031 2751 1032 2752
rect 1036 2751 1037 2755
rect 1190 2755 1196 2756
rect 1190 2754 1191 2755
rect 1141 2752 1191 2754
rect 1031 2750 1037 2751
rect 1190 2751 1191 2752
rect 1195 2751 1196 2755
rect 1279 2755 1285 2756
rect 1279 2754 1280 2755
rect 1261 2752 1280 2754
rect 1190 2750 1196 2751
rect 1279 2751 1280 2752
rect 1284 2751 1285 2755
rect 1391 2755 1397 2756
rect 1391 2754 1392 2755
rect 1373 2752 1392 2754
rect 1279 2750 1285 2751
rect 1391 2751 1392 2752
rect 1396 2751 1397 2755
rect 1503 2755 1509 2756
rect 1503 2754 1504 2755
rect 1485 2752 1504 2754
rect 1391 2750 1397 2751
rect 1503 2751 1504 2752
rect 1508 2751 1509 2755
rect 1607 2755 1613 2756
rect 1607 2754 1608 2755
rect 1589 2752 1608 2754
rect 1503 2750 1509 2751
rect 1607 2751 1608 2752
rect 1612 2751 1613 2755
rect 1711 2755 1717 2756
rect 1711 2754 1712 2755
rect 1701 2752 1712 2754
rect 1607 2750 1613 2751
rect 1711 2751 1712 2752
rect 1716 2751 1717 2755
rect 1794 2755 1800 2756
rect 1794 2754 1795 2755
rect 1789 2752 1795 2754
rect 1711 2750 1717 2751
rect 1794 2751 1795 2752
rect 1799 2751 1800 2755
rect 1822 2752 1823 2756
rect 1827 2752 1828 2756
rect 1822 2751 1828 2752
rect 2022 2755 2028 2756
rect 2022 2751 2023 2755
rect 2027 2754 2028 2755
rect 2075 2755 2081 2756
rect 2075 2754 2076 2755
rect 2027 2752 2076 2754
rect 2027 2751 2028 2752
rect 1794 2750 1800 2751
rect 2022 2750 2028 2751
rect 2075 2751 2076 2752
rect 2080 2751 2081 2755
rect 2075 2750 2081 2751
rect 2111 2755 2117 2756
rect 2111 2751 2112 2755
rect 2116 2754 2117 2755
rect 2195 2755 2201 2756
rect 2195 2754 2196 2755
rect 2116 2752 2196 2754
rect 2116 2751 2117 2752
rect 2111 2750 2117 2751
rect 2195 2751 2196 2752
rect 2200 2751 2201 2755
rect 2195 2750 2201 2751
rect 2239 2755 2245 2756
rect 2239 2751 2240 2755
rect 2244 2754 2245 2755
rect 2323 2755 2329 2756
rect 2323 2754 2324 2755
rect 2244 2752 2324 2754
rect 2244 2751 2245 2752
rect 2239 2750 2245 2751
rect 2323 2751 2324 2752
rect 2328 2751 2329 2755
rect 2323 2750 2329 2751
rect 2475 2755 2481 2756
rect 2475 2751 2476 2755
rect 2480 2754 2481 2755
rect 2498 2755 2504 2756
rect 2498 2754 2499 2755
rect 2480 2752 2499 2754
rect 2480 2751 2481 2752
rect 2475 2750 2481 2751
rect 2498 2751 2499 2752
rect 2503 2751 2504 2755
rect 2498 2750 2504 2751
rect 2651 2755 2657 2756
rect 2651 2751 2652 2755
rect 2656 2754 2657 2755
rect 2706 2755 2712 2756
rect 2706 2754 2707 2755
rect 2656 2752 2707 2754
rect 2656 2751 2657 2752
rect 2651 2750 2657 2751
rect 2706 2751 2707 2752
rect 2711 2751 2712 2755
rect 2706 2750 2712 2751
rect 2851 2755 2857 2756
rect 2851 2751 2852 2755
rect 2856 2754 2857 2755
rect 2903 2755 2909 2756
rect 2903 2754 2904 2755
rect 2856 2752 2904 2754
rect 2856 2751 2857 2752
rect 2851 2750 2857 2751
rect 2903 2751 2904 2752
rect 2908 2751 2909 2755
rect 2903 2750 2909 2751
rect 3067 2755 3073 2756
rect 3067 2751 3068 2755
rect 3072 2754 3073 2755
rect 3098 2755 3104 2756
rect 3098 2754 3099 2755
rect 3072 2752 3099 2754
rect 3072 2751 3073 2752
rect 3067 2750 3073 2751
rect 3098 2751 3099 2752
rect 3103 2751 3104 2755
rect 3098 2750 3104 2751
rect 3198 2755 3204 2756
rect 3198 2751 3199 2755
rect 3203 2754 3204 2755
rect 3299 2755 3305 2756
rect 3299 2754 3300 2755
rect 3203 2752 3300 2754
rect 3203 2751 3204 2752
rect 3198 2750 3204 2751
rect 3299 2751 3300 2752
rect 3304 2751 3305 2755
rect 3299 2750 3305 2751
rect 3515 2755 3521 2756
rect 3515 2751 3516 2755
rect 3520 2754 3521 2755
rect 3546 2755 3552 2756
rect 3546 2754 3547 2755
rect 3520 2752 3547 2754
rect 3520 2751 3521 2752
rect 3515 2750 3521 2751
rect 3546 2751 3547 2752
rect 3551 2751 3552 2755
rect 3546 2750 3552 2751
rect 2046 2745 2052 2746
rect 2046 2741 2047 2745
rect 2051 2741 2052 2745
rect 2046 2740 2052 2741
rect 2166 2745 2172 2746
rect 2166 2741 2167 2745
rect 2171 2741 2172 2745
rect 2166 2740 2172 2741
rect 2294 2745 2300 2746
rect 2294 2741 2295 2745
rect 2299 2741 2300 2745
rect 2294 2740 2300 2741
rect 2446 2745 2452 2746
rect 2446 2741 2447 2745
rect 2451 2741 2452 2745
rect 2446 2740 2452 2741
rect 2622 2745 2628 2746
rect 2622 2741 2623 2745
rect 2627 2741 2628 2745
rect 2622 2740 2628 2741
rect 2822 2745 2828 2746
rect 2822 2741 2823 2745
rect 2827 2741 2828 2745
rect 2822 2740 2828 2741
rect 3038 2745 3044 2746
rect 3038 2741 3039 2745
rect 3043 2741 3044 2745
rect 3038 2740 3044 2741
rect 3270 2745 3276 2746
rect 3270 2741 3271 2745
rect 3275 2741 3276 2745
rect 3270 2740 3276 2741
rect 3486 2745 3492 2746
rect 3486 2741 3487 2745
rect 3491 2741 3492 2745
rect 3486 2740 3492 2741
rect 110 2739 116 2740
rect 110 2735 111 2739
rect 115 2735 116 2739
rect 110 2734 116 2735
rect 414 2739 420 2740
rect 414 2735 415 2739
rect 419 2738 420 2739
rect 1822 2739 1828 2740
rect 419 2736 425 2738
rect 419 2735 420 2736
rect 414 2734 420 2735
rect 1822 2735 1823 2739
rect 1827 2735 1828 2739
rect 1822 2734 1828 2735
rect 1862 2732 1868 2733
rect 3574 2732 3580 2733
rect 182 2729 188 2730
rect 182 2725 183 2729
rect 187 2725 188 2729
rect 182 2724 188 2725
rect 286 2729 292 2730
rect 286 2725 287 2729
rect 291 2725 292 2729
rect 286 2724 292 2725
rect 406 2729 412 2730
rect 406 2725 407 2729
rect 411 2725 412 2729
rect 406 2724 412 2725
rect 542 2729 548 2730
rect 542 2725 543 2729
rect 547 2725 548 2729
rect 542 2724 548 2725
rect 678 2729 684 2730
rect 678 2725 679 2729
rect 683 2725 684 2729
rect 678 2724 684 2725
rect 814 2729 820 2730
rect 814 2725 815 2729
rect 819 2725 820 2729
rect 814 2724 820 2725
rect 950 2729 956 2730
rect 950 2725 951 2729
rect 955 2725 956 2729
rect 950 2724 956 2725
rect 1078 2729 1084 2730
rect 1078 2725 1079 2729
rect 1083 2725 1084 2729
rect 1078 2724 1084 2725
rect 1198 2729 1204 2730
rect 1198 2725 1199 2729
rect 1203 2725 1204 2729
rect 1198 2724 1204 2725
rect 1310 2729 1316 2730
rect 1310 2725 1311 2729
rect 1315 2725 1316 2729
rect 1310 2724 1316 2725
rect 1422 2729 1428 2730
rect 1422 2725 1423 2729
rect 1427 2725 1428 2729
rect 1422 2724 1428 2725
rect 1526 2729 1532 2730
rect 1526 2725 1527 2729
rect 1531 2725 1532 2729
rect 1526 2724 1532 2725
rect 1638 2729 1644 2730
rect 1638 2725 1639 2729
rect 1643 2725 1644 2729
rect 1638 2724 1644 2725
rect 1726 2729 1732 2730
rect 1726 2725 1727 2729
rect 1731 2725 1732 2729
rect 1862 2728 1863 2732
rect 1867 2728 1868 2732
rect 2111 2731 2117 2732
rect 2111 2730 2112 2731
rect 2101 2728 2112 2730
rect 1862 2727 1868 2728
rect 2111 2727 2112 2728
rect 2116 2727 2117 2731
rect 2239 2731 2245 2732
rect 2239 2730 2240 2731
rect 2221 2728 2240 2730
rect 2111 2726 2117 2727
rect 2239 2727 2240 2728
rect 2244 2727 2245 2731
rect 3335 2731 3341 2732
rect 3335 2730 3336 2731
rect 3325 2728 3336 2730
rect 2239 2726 2245 2727
rect 2247 2727 2253 2728
rect 1726 2724 1732 2725
rect 2247 2723 2248 2727
rect 2252 2726 2253 2727
rect 2706 2727 2712 2728
rect 2252 2724 2313 2726
rect 2252 2723 2253 2724
rect 2247 2722 2253 2723
rect 2706 2723 2707 2727
rect 2711 2726 2712 2727
rect 2903 2727 2909 2728
rect 2711 2724 2841 2726
rect 2711 2723 2712 2724
rect 2706 2722 2712 2723
rect 2903 2723 2904 2727
rect 2908 2726 2909 2727
rect 3335 2727 3336 2728
rect 3340 2727 3341 2731
rect 3574 2728 3575 2732
rect 3579 2728 3580 2732
rect 3574 2727 3580 2728
rect 3335 2726 3341 2727
rect 2908 2724 3057 2726
rect 2908 2723 2909 2724
rect 2903 2722 2909 2723
rect 1862 2715 1868 2716
rect 1862 2711 1863 2715
rect 1867 2711 1868 2715
rect 1862 2710 1868 2711
rect 2370 2715 2376 2716
rect 2370 2711 2371 2715
rect 2375 2714 2376 2715
rect 2558 2715 2564 2716
rect 2375 2712 2457 2714
rect 2375 2711 2376 2712
rect 2370 2710 2376 2711
rect 2558 2711 2559 2715
rect 2563 2714 2564 2715
rect 3574 2715 3580 2716
rect 2563 2712 2633 2714
rect 2563 2711 2564 2712
rect 2558 2710 2564 2711
rect 3574 2711 3575 2715
rect 3579 2711 3580 2715
rect 3574 2710 3580 2711
rect 2038 2705 2044 2706
rect 2038 2701 2039 2705
rect 2043 2701 2044 2705
rect 2038 2700 2044 2701
rect 2158 2705 2164 2706
rect 2158 2701 2159 2705
rect 2163 2701 2164 2705
rect 2158 2700 2164 2701
rect 2286 2705 2292 2706
rect 2286 2701 2287 2705
rect 2291 2701 2292 2705
rect 2286 2700 2292 2701
rect 2438 2705 2444 2706
rect 2438 2701 2439 2705
rect 2443 2701 2444 2705
rect 2438 2700 2444 2701
rect 2614 2705 2620 2706
rect 2614 2701 2615 2705
rect 2619 2701 2620 2705
rect 2614 2700 2620 2701
rect 2814 2705 2820 2706
rect 2814 2701 2815 2705
rect 2819 2701 2820 2705
rect 2814 2700 2820 2701
rect 3030 2705 3036 2706
rect 3030 2701 3031 2705
rect 3035 2701 3036 2705
rect 3030 2700 3036 2701
rect 3262 2705 3268 2706
rect 3262 2701 3263 2705
rect 3267 2701 3268 2705
rect 3262 2700 3268 2701
rect 3478 2705 3484 2706
rect 3478 2701 3479 2705
rect 3483 2701 3484 2705
rect 3478 2700 3484 2701
rect 166 2699 172 2700
rect 166 2695 167 2699
rect 171 2695 172 2699
rect 166 2694 172 2695
rect 278 2699 284 2700
rect 278 2695 279 2699
rect 283 2695 284 2699
rect 278 2694 284 2695
rect 390 2699 396 2700
rect 390 2695 391 2699
rect 395 2695 396 2699
rect 390 2694 396 2695
rect 502 2699 508 2700
rect 502 2695 503 2699
rect 507 2695 508 2699
rect 502 2694 508 2695
rect 614 2699 620 2700
rect 614 2695 615 2699
rect 619 2695 620 2699
rect 614 2694 620 2695
rect 3518 2699 3524 2700
rect 3518 2695 3519 2699
rect 3523 2698 3524 2699
rect 3527 2699 3533 2700
rect 3527 2698 3528 2699
rect 3523 2696 3528 2698
rect 3523 2695 3524 2696
rect 3518 2694 3524 2695
rect 3527 2695 3528 2696
rect 3532 2695 3533 2699
rect 3527 2694 3533 2695
rect 570 2691 576 2692
rect 570 2690 571 2691
rect 110 2689 116 2690
rect 110 2685 111 2689
rect 115 2685 116 2689
rect 561 2688 571 2690
rect 570 2687 571 2688
rect 575 2687 576 2691
rect 570 2686 576 2687
rect 1822 2689 1828 2690
rect 110 2684 116 2685
rect 1822 2685 1823 2689
rect 1827 2685 1828 2689
rect 1822 2684 1828 2685
rect 1942 2683 1948 2684
rect 1942 2679 1943 2683
rect 1947 2679 1948 2683
rect 1942 2678 1948 2679
rect 2054 2683 2060 2684
rect 2054 2679 2055 2683
rect 2059 2679 2060 2683
rect 2054 2678 2060 2679
rect 2166 2683 2172 2684
rect 2166 2679 2167 2683
rect 2171 2679 2172 2683
rect 2166 2678 2172 2679
rect 2286 2683 2292 2684
rect 2286 2679 2287 2683
rect 2291 2679 2292 2683
rect 2286 2678 2292 2679
rect 2406 2683 2412 2684
rect 2406 2679 2407 2683
rect 2411 2679 2412 2683
rect 2406 2678 2412 2679
rect 2518 2683 2524 2684
rect 2518 2679 2519 2683
rect 2523 2679 2524 2683
rect 2518 2678 2524 2679
rect 2630 2683 2636 2684
rect 2630 2679 2631 2683
rect 2635 2679 2636 2683
rect 2630 2678 2636 2679
rect 2734 2683 2740 2684
rect 2734 2679 2735 2683
rect 2739 2679 2740 2683
rect 2734 2678 2740 2679
rect 2846 2683 2852 2684
rect 2846 2679 2847 2683
rect 2851 2679 2852 2683
rect 2846 2678 2852 2679
rect 2958 2683 2964 2684
rect 2958 2679 2959 2683
rect 2963 2679 2964 2683
rect 2958 2678 2964 2679
rect 3070 2683 3076 2684
rect 3070 2679 3071 2683
rect 3075 2679 3076 2683
rect 3070 2678 3076 2679
rect 234 2675 240 2676
rect 110 2672 116 2673
rect 110 2668 111 2672
rect 115 2668 116 2672
rect 110 2667 116 2668
rect 228 2666 230 2673
rect 234 2671 235 2675
rect 239 2674 240 2675
rect 346 2675 352 2676
rect 239 2672 305 2674
rect 239 2671 240 2672
rect 234 2670 240 2671
rect 346 2671 347 2675
rect 351 2674 352 2675
rect 570 2675 576 2676
rect 351 2672 417 2674
rect 351 2671 352 2672
rect 346 2670 352 2671
rect 570 2671 571 2675
rect 575 2674 576 2675
rect 2022 2675 2028 2676
rect 2022 2674 2023 2675
rect 575 2672 641 2674
rect 1862 2673 1868 2674
rect 1822 2672 1828 2673
rect 575 2671 576 2672
rect 570 2670 576 2671
rect 1822 2668 1823 2672
rect 1827 2668 1828 2672
rect 1862 2669 1863 2673
rect 1867 2669 1868 2673
rect 2001 2672 2023 2674
rect 2022 2671 2023 2672
rect 2027 2671 2028 2675
rect 3198 2675 3204 2676
rect 3198 2674 3199 2675
rect 3129 2672 3199 2674
rect 2022 2670 2028 2671
rect 3198 2671 3199 2672
rect 3203 2671 3204 2675
rect 3198 2670 3204 2671
rect 3574 2673 3580 2674
rect 1862 2668 1868 2669
rect 3574 2669 3575 2673
rect 3579 2669 3580 2673
rect 3574 2668 3580 2669
rect 250 2667 256 2668
rect 1822 2667 1828 2668
rect 250 2666 251 2667
rect 228 2664 251 2666
rect 250 2663 251 2664
rect 255 2663 256 2667
rect 250 2662 256 2663
rect 174 2659 180 2660
rect 174 2655 175 2659
rect 179 2655 180 2659
rect 174 2654 180 2655
rect 286 2659 292 2660
rect 286 2655 287 2659
rect 291 2655 292 2659
rect 286 2654 292 2655
rect 398 2659 404 2660
rect 398 2655 399 2659
rect 403 2655 404 2659
rect 398 2654 404 2655
rect 510 2659 516 2660
rect 510 2655 511 2659
rect 515 2655 516 2659
rect 510 2654 516 2655
rect 622 2659 628 2660
rect 622 2655 623 2659
rect 627 2655 628 2659
rect 2010 2659 2016 2660
rect 622 2654 628 2655
rect 1862 2656 1868 2657
rect 1862 2652 1863 2656
rect 1867 2652 1868 2656
rect 2010 2655 2011 2659
rect 2015 2658 2016 2659
rect 2122 2659 2128 2660
rect 2015 2656 2081 2658
rect 2015 2655 2016 2656
rect 2010 2654 2016 2655
rect 2122 2655 2123 2659
rect 2127 2658 2128 2659
rect 2399 2659 2405 2660
rect 2399 2658 2400 2659
rect 2127 2656 2193 2658
rect 2349 2656 2400 2658
rect 2127 2655 2128 2656
rect 2122 2654 2128 2655
rect 2399 2655 2400 2656
rect 2404 2655 2405 2659
rect 2490 2659 2496 2660
rect 2490 2658 2491 2659
rect 2469 2656 2491 2658
rect 2399 2654 2405 2655
rect 2490 2655 2491 2656
rect 2495 2655 2496 2659
rect 2623 2659 2629 2660
rect 2623 2658 2624 2659
rect 2581 2656 2624 2658
rect 2490 2654 2496 2655
rect 2623 2655 2624 2656
rect 2628 2655 2629 2659
rect 2727 2659 2733 2660
rect 2727 2658 2728 2659
rect 2693 2656 2728 2658
rect 2623 2654 2629 2655
rect 2727 2655 2728 2656
rect 2732 2655 2733 2659
rect 2839 2659 2845 2660
rect 2839 2658 2840 2659
rect 2797 2656 2840 2658
rect 2727 2654 2733 2655
rect 2839 2655 2840 2656
rect 2844 2655 2845 2659
rect 2951 2659 2957 2660
rect 2951 2658 2952 2659
rect 2909 2656 2952 2658
rect 2839 2654 2845 2655
rect 2951 2655 2952 2656
rect 2956 2655 2957 2659
rect 3063 2659 3069 2660
rect 3063 2658 3064 2659
rect 3021 2656 3064 2658
rect 2951 2654 2957 2655
rect 3063 2655 3064 2656
rect 3068 2655 3069 2659
rect 3063 2654 3069 2655
rect 3574 2656 3580 2657
rect 1862 2651 1868 2652
rect 3574 2652 3575 2656
rect 3579 2652 3580 2656
rect 3574 2651 3580 2652
rect 203 2647 209 2648
rect 203 2643 204 2647
rect 208 2646 209 2647
rect 234 2647 240 2648
rect 234 2646 235 2647
rect 208 2644 235 2646
rect 208 2643 209 2644
rect 203 2642 209 2643
rect 234 2643 235 2644
rect 239 2643 240 2647
rect 234 2642 240 2643
rect 315 2647 321 2648
rect 315 2643 316 2647
rect 320 2646 321 2647
rect 346 2647 352 2648
rect 346 2646 347 2647
rect 320 2644 347 2646
rect 320 2643 321 2644
rect 315 2642 321 2643
rect 346 2643 347 2644
rect 351 2643 352 2647
rect 346 2642 352 2643
rect 414 2647 420 2648
rect 414 2643 415 2647
rect 419 2646 420 2647
rect 427 2647 433 2648
rect 427 2646 428 2647
rect 419 2644 428 2646
rect 419 2643 420 2644
rect 414 2642 420 2643
rect 427 2643 428 2644
rect 432 2643 433 2647
rect 427 2642 433 2643
rect 539 2647 545 2648
rect 539 2643 540 2647
rect 544 2646 545 2647
rect 570 2647 576 2648
rect 570 2646 571 2647
rect 544 2644 571 2646
rect 544 2643 545 2644
rect 539 2642 545 2643
rect 570 2643 571 2644
rect 575 2643 576 2647
rect 570 2642 576 2643
rect 651 2647 660 2648
rect 651 2643 652 2647
rect 659 2643 660 2647
rect 651 2642 660 2643
rect 1950 2643 1956 2644
rect 1950 2639 1951 2643
rect 1955 2639 1956 2643
rect 1950 2638 1956 2639
rect 2062 2643 2068 2644
rect 2062 2639 2063 2643
rect 2067 2639 2068 2643
rect 2062 2638 2068 2639
rect 2174 2643 2180 2644
rect 2174 2639 2175 2643
rect 2179 2639 2180 2643
rect 2174 2638 2180 2639
rect 2294 2643 2300 2644
rect 2294 2639 2295 2643
rect 2299 2639 2300 2643
rect 2294 2638 2300 2639
rect 2414 2643 2420 2644
rect 2414 2639 2415 2643
rect 2419 2639 2420 2643
rect 2414 2638 2420 2639
rect 2526 2643 2532 2644
rect 2526 2639 2527 2643
rect 2531 2639 2532 2643
rect 2526 2638 2532 2639
rect 2638 2643 2644 2644
rect 2638 2639 2639 2643
rect 2643 2639 2644 2643
rect 2638 2638 2644 2639
rect 2742 2643 2748 2644
rect 2742 2639 2743 2643
rect 2747 2639 2748 2643
rect 2742 2638 2748 2639
rect 2854 2643 2860 2644
rect 2854 2639 2855 2643
rect 2859 2639 2860 2643
rect 2854 2638 2860 2639
rect 2966 2643 2972 2644
rect 2966 2639 2967 2643
rect 2971 2639 2972 2643
rect 2966 2638 2972 2639
rect 3078 2643 3084 2644
rect 3078 2639 3079 2643
rect 3083 2639 3084 2643
rect 3078 2638 3084 2639
rect 1979 2631 1985 2632
rect 1979 2627 1980 2631
rect 1984 2630 1985 2631
rect 2010 2631 2016 2632
rect 2010 2630 2011 2631
rect 1984 2628 2011 2630
rect 1984 2627 1985 2628
rect 1979 2626 1985 2627
rect 2010 2627 2011 2628
rect 2015 2627 2016 2631
rect 2010 2626 2016 2627
rect 2091 2631 2097 2632
rect 2091 2627 2092 2631
rect 2096 2630 2097 2631
rect 2122 2631 2128 2632
rect 2122 2630 2123 2631
rect 2096 2628 2123 2630
rect 2096 2627 2097 2628
rect 2091 2626 2097 2627
rect 2122 2627 2123 2628
rect 2127 2627 2128 2631
rect 2122 2626 2128 2627
rect 2203 2631 2209 2632
rect 2203 2627 2204 2631
rect 2208 2630 2209 2631
rect 2238 2631 2244 2632
rect 2238 2630 2239 2631
rect 2208 2628 2239 2630
rect 2208 2627 2209 2628
rect 2203 2626 2209 2627
rect 2238 2627 2239 2628
rect 2243 2627 2244 2631
rect 2238 2626 2244 2627
rect 2323 2631 2329 2632
rect 2323 2627 2324 2631
rect 2328 2630 2329 2631
rect 2370 2631 2376 2632
rect 2370 2630 2371 2631
rect 2328 2628 2371 2630
rect 2328 2627 2329 2628
rect 2323 2626 2329 2627
rect 2370 2627 2371 2628
rect 2375 2627 2376 2631
rect 2370 2626 2376 2627
rect 2399 2631 2405 2632
rect 2399 2627 2400 2631
rect 2404 2630 2405 2631
rect 2443 2631 2449 2632
rect 2443 2630 2444 2631
rect 2404 2628 2444 2630
rect 2404 2627 2405 2628
rect 2399 2626 2405 2627
rect 2443 2627 2444 2628
rect 2448 2627 2449 2631
rect 2443 2626 2449 2627
rect 2555 2631 2564 2632
rect 2555 2627 2556 2631
rect 2563 2627 2564 2631
rect 2555 2626 2564 2627
rect 2623 2631 2629 2632
rect 2623 2627 2624 2631
rect 2628 2630 2629 2631
rect 2667 2631 2673 2632
rect 2667 2630 2668 2631
rect 2628 2628 2668 2630
rect 2628 2627 2629 2628
rect 2623 2626 2629 2627
rect 2667 2627 2668 2628
rect 2672 2627 2673 2631
rect 2667 2626 2673 2627
rect 2727 2631 2733 2632
rect 2727 2627 2728 2631
rect 2732 2630 2733 2631
rect 2771 2631 2777 2632
rect 2771 2630 2772 2631
rect 2732 2628 2772 2630
rect 2732 2627 2733 2628
rect 2727 2626 2733 2627
rect 2771 2627 2772 2628
rect 2776 2627 2777 2631
rect 2771 2626 2777 2627
rect 2839 2631 2845 2632
rect 2839 2627 2840 2631
rect 2844 2630 2845 2631
rect 2883 2631 2889 2632
rect 2883 2630 2884 2631
rect 2844 2628 2884 2630
rect 2844 2627 2845 2628
rect 2839 2626 2845 2627
rect 2883 2627 2884 2628
rect 2888 2627 2889 2631
rect 2883 2626 2889 2627
rect 2951 2631 2957 2632
rect 2951 2627 2952 2631
rect 2956 2630 2957 2631
rect 2995 2631 3001 2632
rect 2995 2630 2996 2631
rect 2956 2628 2996 2630
rect 2956 2627 2957 2628
rect 2951 2626 2957 2627
rect 2995 2627 2996 2628
rect 3000 2627 3001 2631
rect 2995 2626 3001 2627
rect 3063 2631 3069 2632
rect 3063 2627 3064 2631
rect 3068 2630 3069 2631
rect 3107 2631 3113 2632
rect 3107 2630 3108 2631
rect 3068 2628 3108 2630
rect 3068 2627 3069 2628
rect 3063 2626 3069 2627
rect 3107 2627 3108 2628
rect 3112 2627 3113 2631
rect 3107 2626 3113 2627
rect 250 2619 257 2620
rect 250 2615 251 2619
rect 256 2615 257 2619
rect 250 2614 257 2615
rect 335 2619 341 2620
rect 335 2615 336 2619
rect 340 2618 341 2619
rect 379 2619 385 2620
rect 379 2618 380 2619
rect 340 2616 380 2618
rect 340 2615 341 2616
rect 335 2614 341 2615
rect 379 2615 380 2616
rect 384 2615 385 2619
rect 379 2614 385 2615
rect 439 2619 445 2620
rect 439 2615 440 2619
rect 444 2618 445 2619
rect 523 2619 529 2620
rect 523 2618 524 2619
rect 444 2616 524 2618
rect 444 2615 445 2616
rect 439 2614 445 2615
rect 523 2615 524 2616
rect 528 2615 529 2619
rect 523 2614 529 2615
rect 691 2619 697 2620
rect 691 2615 692 2619
rect 696 2618 697 2619
rect 758 2619 764 2620
rect 758 2618 759 2619
rect 696 2616 759 2618
rect 696 2615 697 2616
rect 691 2614 697 2615
rect 758 2615 759 2616
rect 763 2615 764 2619
rect 758 2614 764 2615
rect 867 2619 873 2620
rect 867 2615 868 2619
rect 872 2618 873 2619
rect 906 2619 912 2620
rect 906 2618 907 2619
rect 872 2616 907 2618
rect 872 2615 873 2616
rect 867 2614 873 2615
rect 906 2615 907 2616
rect 911 2615 912 2619
rect 906 2614 912 2615
rect 966 2619 972 2620
rect 966 2615 967 2619
rect 971 2618 972 2619
rect 1051 2619 1057 2620
rect 1051 2618 1052 2619
rect 971 2616 1052 2618
rect 971 2615 972 2616
rect 966 2614 972 2615
rect 1051 2615 1052 2616
rect 1056 2615 1057 2619
rect 1051 2614 1057 2615
rect 1243 2619 1252 2620
rect 1243 2615 1244 2619
rect 1251 2615 1252 2619
rect 1243 2614 1252 2615
rect 1327 2619 1333 2620
rect 1327 2615 1328 2619
rect 1332 2618 1333 2619
rect 1435 2619 1441 2620
rect 1435 2618 1436 2619
rect 1332 2616 1436 2618
rect 1332 2615 1333 2616
rect 1327 2614 1333 2615
rect 1435 2615 1436 2616
rect 1440 2615 1441 2619
rect 1435 2614 1441 2615
rect 1527 2619 1533 2620
rect 1527 2615 1528 2619
rect 1532 2618 1533 2619
rect 1635 2619 1641 2620
rect 1635 2618 1636 2619
rect 1532 2616 1636 2618
rect 1532 2615 1533 2616
rect 1527 2614 1533 2615
rect 1635 2615 1636 2616
rect 1640 2615 1641 2619
rect 1635 2614 1641 2615
rect 1923 2615 1929 2616
rect 1923 2611 1924 2615
rect 1928 2614 1929 2615
rect 1958 2615 1964 2616
rect 1958 2614 1959 2615
rect 1928 2612 1959 2614
rect 1928 2611 1929 2612
rect 1923 2610 1929 2611
rect 1958 2611 1959 2612
rect 1963 2611 1964 2615
rect 1958 2610 1964 2611
rect 1999 2615 2005 2616
rect 1999 2611 2000 2615
rect 2004 2614 2005 2615
rect 2099 2615 2105 2616
rect 2099 2614 2100 2615
rect 2004 2612 2100 2614
rect 2004 2611 2005 2612
rect 1999 2610 2005 2611
rect 2099 2611 2100 2612
rect 2104 2611 2105 2615
rect 2099 2610 2105 2611
rect 2183 2615 2189 2616
rect 2183 2611 2184 2615
rect 2188 2614 2189 2615
rect 2291 2615 2297 2616
rect 2291 2614 2292 2615
rect 2188 2612 2292 2614
rect 2188 2611 2189 2612
rect 2183 2610 2189 2611
rect 2291 2611 2292 2612
rect 2296 2611 2297 2615
rect 2291 2610 2297 2611
rect 2490 2615 2497 2616
rect 2490 2611 2491 2615
rect 2496 2611 2497 2615
rect 2490 2610 2497 2611
rect 2583 2615 2589 2616
rect 2583 2611 2584 2615
rect 2588 2614 2589 2615
rect 2691 2615 2697 2616
rect 2691 2614 2692 2615
rect 2588 2612 2692 2614
rect 2588 2611 2589 2612
rect 2583 2610 2589 2611
rect 2691 2611 2692 2612
rect 2696 2611 2697 2615
rect 2691 2610 2697 2611
rect 2899 2615 2905 2616
rect 2899 2611 2900 2615
rect 2904 2614 2905 2615
rect 2958 2615 2964 2616
rect 2958 2614 2959 2615
rect 2904 2612 2959 2614
rect 2904 2611 2905 2612
rect 2899 2610 2905 2611
rect 2958 2611 2959 2612
rect 2963 2611 2964 2615
rect 2958 2610 2964 2611
rect 3107 2615 3113 2616
rect 3107 2611 3108 2615
rect 3112 2614 3113 2615
rect 3151 2615 3157 2616
rect 3151 2614 3152 2615
rect 3112 2612 3152 2614
rect 3112 2611 3113 2612
rect 3107 2610 3113 2611
rect 3151 2611 3152 2612
rect 3156 2611 3157 2615
rect 3151 2610 3157 2611
rect 3271 2615 3277 2616
rect 3271 2611 3272 2615
rect 3276 2614 3277 2615
rect 3323 2615 3329 2616
rect 3323 2614 3324 2615
rect 3276 2612 3324 2614
rect 3276 2611 3277 2612
rect 3271 2610 3277 2611
rect 3323 2611 3324 2612
rect 3328 2611 3329 2615
rect 3323 2610 3329 2611
rect 3515 2615 3524 2616
rect 3515 2611 3516 2615
rect 3523 2611 3524 2615
rect 3515 2610 3524 2611
rect 222 2609 228 2610
rect 222 2605 223 2609
rect 227 2605 228 2609
rect 222 2604 228 2605
rect 350 2609 356 2610
rect 350 2605 351 2609
rect 355 2605 356 2609
rect 350 2604 356 2605
rect 494 2609 500 2610
rect 494 2605 495 2609
rect 499 2605 500 2609
rect 494 2604 500 2605
rect 662 2609 668 2610
rect 662 2605 663 2609
rect 667 2605 668 2609
rect 662 2604 668 2605
rect 838 2609 844 2610
rect 838 2605 839 2609
rect 843 2605 844 2609
rect 838 2604 844 2605
rect 1022 2609 1028 2610
rect 1022 2605 1023 2609
rect 1027 2605 1028 2609
rect 1022 2604 1028 2605
rect 1214 2609 1220 2610
rect 1214 2605 1215 2609
rect 1219 2605 1220 2609
rect 1214 2604 1220 2605
rect 1406 2609 1412 2610
rect 1406 2605 1407 2609
rect 1411 2605 1412 2609
rect 1406 2604 1412 2605
rect 1606 2609 1612 2610
rect 1606 2605 1607 2609
rect 1611 2605 1612 2609
rect 1606 2604 1612 2605
rect 1894 2605 1900 2606
rect 1894 2601 1895 2605
rect 1899 2601 1900 2605
rect 1894 2600 1900 2601
rect 2070 2605 2076 2606
rect 2070 2601 2071 2605
rect 2075 2601 2076 2605
rect 2070 2600 2076 2601
rect 2262 2605 2268 2606
rect 2262 2601 2263 2605
rect 2267 2601 2268 2605
rect 2262 2600 2268 2601
rect 2462 2605 2468 2606
rect 2462 2601 2463 2605
rect 2467 2601 2468 2605
rect 2462 2600 2468 2601
rect 2662 2605 2668 2606
rect 2662 2601 2663 2605
rect 2667 2601 2668 2605
rect 2662 2600 2668 2601
rect 2870 2605 2876 2606
rect 2870 2601 2871 2605
rect 2875 2601 2876 2605
rect 2870 2600 2876 2601
rect 3078 2605 3084 2606
rect 3078 2601 3079 2605
rect 3083 2601 3084 2605
rect 3078 2600 3084 2601
rect 3294 2605 3300 2606
rect 3294 2601 3295 2605
rect 3299 2601 3300 2605
rect 3294 2600 3300 2601
rect 3486 2605 3492 2606
rect 3486 2601 3487 2605
rect 3491 2601 3492 2605
rect 3486 2600 3492 2601
rect 110 2596 116 2597
rect 1822 2596 1828 2597
rect 110 2592 111 2596
rect 115 2592 116 2596
rect 335 2595 341 2596
rect 335 2594 336 2595
rect 277 2592 336 2594
rect 110 2591 116 2592
rect 335 2591 336 2592
rect 340 2591 341 2595
rect 439 2595 445 2596
rect 439 2594 440 2595
rect 405 2592 440 2594
rect 335 2590 341 2591
rect 439 2591 440 2592
rect 444 2591 445 2595
rect 1327 2595 1333 2596
rect 1327 2594 1328 2595
rect 1269 2592 1328 2594
rect 439 2590 445 2591
rect 654 2591 660 2592
rect 654 2587 655 2591
rect 659 2590 660 2591
rect 758 2591 764 2592
rect 659 2588 681 2590
rect 659 2587 660 2588
rect 654 2586 660 2587
rect 758 2587 759 2591
rect 763 2590 764 2591
rect 906 2591 912 2592
rect 763 2588 857 2590
rect 763 2587 764 2588
rect 758 2586 764 2587
rect 906 2587 907 2591
rect 911 2590 912 2591
rect 1327 2591 1328 2592
rect 1332 2591 1333 2595
rect 1527 2595 1533 2596
rect 1527 2594 1528 2595
rect 1461 2592 1528 2594
rect 1327 2590 1333 2591
rect 1527 2591 1528 2592
rect 1532 2591 1533 2595
rect 1822 2592 1823 2596
rect 1827 2592 1828 2596
rect 1822 2591 1828 2592
rect 1862 2592 1868 2593
rect 3574 2592 3580 2593
rect 1527 2590 1533 2591
rect 911 2588 1041 2590
rect 1862 2588 1863 2592
rect 1867 2588 1868 2592
rect 1999 2591 2005 2592
rect 1999 2590 2000 2591
rect 1949 2588 2000 2590
rect 911 2587 912 2588
rect 1862 2587 1868 2588
rect 1999 2587 2000 2588
rect 2004 2587 2005 2591
rect 2183 2591 2189 2592
rect 2183 2590 2184 2591
rect 2125 2588 2184 2590
rect 906 2586 912 2587
rect 1999 2586 2005 2587
rect 2183 2587 2184 2588
rect 2188 2587 2189 2591
rect 2583 2591 2589 2592
rect 2583 2590 2584 2591
rect 2517 2588 2584 2590
rect 2183 2586 2189 2587
rect 2238 2587 2244 2588
rect 2238 2583 2239 2587
rect 2243 2586 2244 2587
rect 2583 2587 2584 2588
rect 2588 2587 2589 2591
rect 3574 2588 3575 2592
rect 3579 2588 3580 2592
rect 2583 2586 2589 2587
rect 2958 2587 2964 2588
rect 2243 2584 2281 2586
rect 2243 2583 2244 2584
rect 2238 2582 2244 2583
rect 2958 2583 2959 2587
rect 2963 2586 2964 2587
rect 3151 2587 3157 2588
rect 3574 2587 3580 2588
rect 2963 2584 3097 2586
rect 2963 2583 2964 2584
rect 2958 2582 2964 2583
rect 3151 2583 3152 2587
rect 3156 2586 3157 2587
rect 3156 2584 3313 2586
rect 3156 2583 3157 2584
rect 3151 2582 3157 2583
rect 110 2579 116 2580
rect 110 2575 111 2579
rect 115 2575 116 2579
rect 110 2574 116 2575
rect 494 2579 500 2580
rect 494 2575 495 2579
rect 499 2578 500 2579
rect 1762 2579 1768 2580
rect 1762 2578 1763 2579
rect 499 2576 505 2578
rect 1657 2576 1763 2578
rect 499 2575 500 2576
rect 494 2574 500 2575
rect 1762 2575 1763 2576
rect 1767 2575 1768 2579
rect 1762 2574 1768 2575
rect 1822 2579 1828 2580
rect 1822 2575 1823 2579
rect 1827 2575 1828 2579
rect 1822 2574 1828 2575
rect 1862 2575 1868 2576
rect 1862 2571 1863 2575
rect 1867 2571 1868 2575
rect 1862 2570 1868 2571
rect 2530 2575 2536 2576
rect 2530 2571 2531 2575
rect 2535 2574 2536 2575
rect 2782 2575 2788 2576
rect 2535 2572 2673 2574
rect 2535 2571 2536 2572
rect 2530 2570 2536 2571
rect 2782 2571 2783 2575
rect 2787 2574 2788 2575
rect 3574 2575 3580 2576
rect 2787 2572 2881 2574
rect 2787 2571 2788 2572
rect 2782 2570 2788 2571
rect 3574 2571 3575 2575
rect 3579 2571 3580 2575
rect 3574 2570 3580 2571
rect 214 2569 220 2570
rect 214 2565 215 2569
rect 219 2565 220 2569
rect 214 2564 220 2565
rect 342 2569 348 2570
rect 342 2565 343 2569
rect 347 2565 348 2569
rect 342 2564 348 2565
rect 486 2569 492 2570
rect 486 2565 487 2569
rect 491 2565 492 2569
rect 486 2564 492 2565
rect 654 2569 660 2570
rect 654 2565 655 2569
rect 659 2565 660 2569
rect 654 2564 660 2565
rect 830 2569 836 2570
rect 830 2565 831 2569
rect 835 2565 836 2569
rect 830 2564 836 2565
rect 1014 2569 1020 2570
rect 1014 2565 1015 2569
rect 1019 2565 1020 2569
rect 1014 2564 1020 2565
rect 1206 2569 1212 2570
rect 1206 2565 1207 2569
rect 1211 2565 1212 2569
rect 1206 2564 1212 2565
rect 1398 2569 1404 2570
rect 1398 2565 1399 2569
rect 1403 2565 1404 2569
rect 1398 2564 1404 2565
rect 1598 2569 1604 2570
rect 1598 2565 1599 2569
rect 1603 2565 1604 2569
rect 1598 2564 1604 2565
rect 1886 2565 1892 2566
rect 1886 2561 1887 2565
rect 1891 2561 1892 2565
rect 1886 2560 1892 2561
rect 2062 2565 2068 2566
rect 2062 2561 2063 2565
rect 2067 2561 2068 2565
rect 2062 2560 2068 2561
rect 2254 2565 2260 2566
rect 2254 2561 2255 2565
rect 2259 2561 2260 2565
rect 2254 2560 2260 2561
rect 2454 2565 2460 2566
rect 2454 2561 2455 2565
rect 2459 2561 2460 2565
rect 2454 2560 2460 2561
rect 2654 2565 2660 2566
rect 2654 2561 2655 2565
rect 2659 2561 2660 2565
rect 2654 2560 2660 2561
rect 2862 2565 2868 2566
rect 2862 2561 2863 2565
rect 2867 2561 2868 2565
rect 2862 2560 2868 2561
rect 3070 2565 3076 2566
rect 3070 2561 3071 2565
rect 3075 2561 3076 2565
rect 3070 2560 3076 2561
rect 3286 2565 3292 2566
rect 3286 2561 3287 2565
rect 3291 2561 3292 2565
rect 3286 2560 3292 2561
rect 3478 2565 3484 2566
rect 3478 2561 3479 2565
rect 3483 2561 3484 2565
rect 3478 2560 3484 2561
rect 3518 2559 3524 2560
rect 3518 2555 3519 2559
rect 3523 2558 3524 2559
rect 3527 2559 3533 2560
rect 3527 2558 3528 2559
rect 3523 2556 3528 2558
rect 3523 2555 3524 2556
rect 3518 2554 3524 2555
rect 3527 2555 3528 2556
rect 3532 2555 3533 2559
rect 3527 2554 3533 2555
rect 270 2547 276 2548
rect 270 2543 271 2547
rect 275 2543 276 2547
rect 270 2542 276 2543
rect 470 2547 476 2548
rect 470 2543 471 2547
rect 475 2543 476 2547
rect 470 2542 476 2543
rect 670 2547 676 2548
rect 670 2543 671 2547
rect 675 2543 676 2547
rect 670 2542 676 2543
rect 854 2547 860 2548
rect 854 2543 855 2547
rect 859 2543 860 2547
rect 854 2542 860 2543
rect 1022 2547 1028 2548
rect 1022 2543 1023 2547
rect 1027 2543 1028 2547
rect 1022 2542 1028 2543
rect 1174 2547 1180 2548
rect 1174 2543 1175 2547
rect 1179 2543 1180 2547
rect 1174 2542 1180 2543
rect 1318 2547 1324 2548
rect 1318 2543 1319 2547
rect 1323 2543 1324 2547
rect 1318 2542 1324 2543
rect 1454 2547 1460 2548
rect 1454 2543 1455 2547
rect 1459 2543 1460 2547
rect 1454 2542 1460 2543
rect 1590 2547 1596 2548
rect 1590 2543 1591 2547
rect 1595 2543 1596 2547
rect 1590 2542 1596 2543
rect 1726 2547 1732 2548
rect 1726 2543 1727 2547
rect 1731 2543 1732 2547
rect 1726 2542 1732 2543
rect 1886 2543 1892 2544
rect 966 2539 972 2540
rect 966 2538 967 2539
rect 110 2537 116 2538
rect 110 2533 111 2537
rect 115 2533 116 2537
rect 913 2536 967 2538
rect 966 2535 967 2536
rect 971 2535 972 2539
rect 966 2534 972 2535
rect 1246 2539 1252 2540
rect 1246 2535 1247 2539
rect 1251 2538 1252 2539
rect 1886 2539 1887 2543
rect 1891 2539 1892 2543
rect 1886 2538 1892 2539
rect 2038 2543 2044 2544
rect 2038 2539 2039 2543
rect 2043 2539 2044 2543
rect 2038 2538 2044 2539
rect 2214 2543 2220 2544
rect 2214 2539 2215 2543
rect 2219 2539 2220 2543
rect 2214 2538 2220 2539
rect 2398 2543 2404 2544
rect 2398 2539 2399 2543
rect 2403 2539 2404 2543
rect 2398 2538 2404 2539
rect 2574 2543 2580 2544
rect 2574 2539 2575 2543
rect 2579 2539 2580 2543
rect 2574 2538 2580 2539
rect 2742 2543 2748 2544
rect 2742 2539 2743 2543
rect 2747 2539 2748 2543
rect 2742 2538 2748 2539
rect 2902 2543 2908 2544
rect 2902 2539 2903 2543
rect 2907 2539 2908 2543
rect 2902 2538 2908 2539
rect 3054 2543 3060 2544
rect 3054 2539 3055 2543
rect 3059 2539 3060 2543
rect 3054 2538 3060 2539
rect 3198 2543 3204 2544
rect 3198 2539 3199 2543
rect 3203 2539 3204 2543
rect 3198 2538 3204 2539
rect 3342 2543 3348 2544
rect 3342 2539 3343 2543
rect 3347 2539 3348 2543
rect 3342 2538 3348 2539
rect 3478 2543 3484 2544
rect 3478 2539 3479 2543
rect 3483 2539 3484 2543
rect 3478 2538 3484 2539
rect 1251 2536 1337 2538
rect 1822 2537 1828 2538
rect 1251 2535 1252 2536
rect 1246 2534 1252 2535
rect 110 2532 116 2533
rect 1822 2533 1823 2537
rect 1827 2533 1828 2537
rect 1958 2535 1964 2536
rect 1958 2534 1959 2535
rect 1822 2532 1828 2533
rect 1862 2533 1868 2534
rect 1862 2529 1863 2533
rect 1867 2529 1868 2533
rect 1945 2532 1959 2534
rect 1958 2531 1959 2532
rect 1963 2531 1964 2535
rect 3271 2535 3277 2536
rect 3271 2534 3272 2535
rect 3257 2532 3272 2534
rect 1958 2530 1964 2531
rect 3271 2531 3272 2532
rect 3276 2531 3277 2535
rect 3271 2530 3277 2531
rect 3574 2533 3580 2534
rect 1862 2528 1868 2529
rect 3574 2529 3575 2533
rect 3579 2529 3580 2533
rect 3574 2528 3580 2529
rect 214 2523 220 2524
rect 110 2520 116 2521
rect 110 2516 111 2520
rect 115 2516 116 2520
rect 214 2519 215 2523
rect 219 2522 220 2523
rect 338 2523 344 2524
rect 219 2520 297 2522
rect 219 2519 220 2520
rect 214 2518 220 2519
rect 338 2519 339 2523
rect 343 2522 344 2523
rect 847 2523 853 2524
rect 847 2522 848 2523
rect 343 2520 497 2522
rect 733 2520 848 2522
rect 343 2519 344 2520
rect 338 2518 344 2519
rect 847 2519 848 2520
rect 852 2519 853 2523
rect 1158 2523 1164 2524
rect 1158 2522 1159 2523
rect 1085 2520 1159 2522
rect 847 2518 853 2519
rect 1158 2519 1159 2520
rect 1163 2519 1164 2523
rect 1311 2523 1317 2524
rect 1311 2522 1312 2523
rect 1237 2520 1312 2522
rect 1158 2518 1164 2519
rect 1311 2519 1312 2520
rect 1316 2519 1317 2523
rect 1311 2518 1317 2519
rect 1386 2523 1392 2524
rect 1386 2519 1387 2523
rect 1391 2522 1392 2523
rect 1522 2523 1528 2524
rect 1391 2520 1481 2522
rect 1391 2519 1392 2520
rect 1386 2518 1392 2519
rect 1522 2519 1523 2523
rect 1527 2522 1528 2523
rect 1658 2523 1664 2524
rect 1527 2520 1617 2522
rect 1527 2519 1528 2520
rect 1522 2518 1528 2519
rect 1658 2519 1659 2523
rect 1663 2522 1664 2523
rect 1663 2520 1753 2522
rect 1822 2520 1828 2521
rect 1663 2519 1664 2520
rect 1658 2518 1664 2519
rect 110 2515 116 2516
rect 1822 2516 1823 2520
rect 1827 2516 1828 2520
rect 1954 2519 1960 2520
rect 1822 2515 1828 2516
rect 1862 2516 1868 2517
rect 1862 2512 1863 2516
rect 1867 2512 1868 2516
rect 1954 2515 1955 2519
rect 1959 2518 1960 2519
rect 2106 2519 2112 2520
rect 1959 2516 2065 2518
rect 1959 2515 1960 2516
rect 1954 2514 1960 2515
rect 2106 2515 2107 2519
rect 2111 2518 2112 2519
rect 2567 2519 2573 2520
rect 2567 2518 2568 2519
rect 2111 2516 2241 2518
rect 2461 2516 2568 2518
rect 2111 2515 2112 2516
rect 2106 2514 2112 2515
rect 2567 2515 2568 2516
rect 2572 2515 2573 2519
rect 2642 2519 2648 2520
rect 2642 2518 2643 2519
rect 2637 2516 2643 2518
rect 2567 2514 2573 2515
rect 2642 2515 2643 2516
rect 2647 2515 2648 2519
rect 2895 2519 2901 2520
rect 2895 2518 2896 2519
rect 2805 2516 2896 2518
rect 2642 2514 2648 2515
rect 2895 2515 2896 2516
rect 2900 2515 2901 2519
rect 3047 2519 3053 2520
rect 3047 2518 3048 2519
rect 2965 2516 3048 2518
rect 2895 2514 2901 2515
rect 3047 2515 3048 2516
rect 3052 2515 3053 2519
rect 3146 2519 3152 2520
rect 3146 2518 3147 2519
rect 3117 2516 3147 2518
rect 3047 2514 3053 2515
rect 3146 2515 3147 2516
rect 3151 2515 3152 2519
rect 3146 2514 3152 2515
rect 3266 2519 3272 2520
rect 3266 2515 3267 2519
rect 3271 2518 3272 2519
rect 3546 2519 3552 2520
rect 3546 2518 3547 2519
rect 3271 2516 3369 2518
rect 3541 2516 3547 2518
rect 3271 2515 3272 2516
rect 3266 2514 3272 2515
rect 3546 2515 3547 2516
rect 3551 2515 3552 2519
rect 3546 2514 3552 2515
rect 3574 2516 3580 2517
rect 1862 2511 1868 2512
rect 3574 2512 3575 2516
rect 3579 2512 3580 2516
rect 3574 2511 3580 2512
rect 278 2507 284 2508
rect 278 2503 279 2507
rect 283 2503 284 2507
rect 278 2502 284 2503
rect 478 2507 484 2508
rect 478 2503 479 2507
rect 483 2503 484 2507
rect 478 2502 484 2503
rect 678 2507 684 2508
rect 678 2503 679 2507
rect 683 2503 684 2507
rect 678 2502 684 2503
rect 862 2507 868 2508
rect 862 2503 863 2507
rect 867 2503 868 2507
rect 862 2502 868 2503
rect 1030 2507 1036 2508
rect 1030 2503 1031 2507
rect 1035 2503 1036 2507
rect 1030 2502 1036 2503
rect 1182 2507 1188 2508
rect 1182 2503 1183 2507
rect 1187 2503 1188 2507
rect 1182 2502 1188 2503
rect 1326 2507 1332 2508
rect 1326 2503 1327 2507
rect 1331 2503 1332 2507
rect 1326 2502 1332 2503
rect 1462 2507 1468 2508
rect 1462 2503 1463 2507
rect 1467 2503 1468 2507
rect 1462 2502 1468 2503
rect 1598 2507 1604 2508
rect 1598 2503 1599 2507
rect 1603 2503 1604 2507
rect 1598 2502 1604 2503
rect 1734 2507 1740 2508
rect 1734 2503 1735 2507
rect 1739 2503 1740 2507
rect 1734 2502 1740 2503
rect 1894 2503 1900 2504
rect 1894 2499 1895 2503
rect 1899 2499 1900 2503
rect 1894 2498 1900 2499
rect 2046 2503 2052 2504
rect 2046 2499 2047 2503
rect 2051 2499 2052 2503
rect 2046 2498 2052 2499
rect 2222 2503 2228 2504
rect 2222 2499 2223 2503
rect 2227 2499 2228 2503
rect 2222 2498 2228 2499
rect 2406 2503 2412 2504
rect 2406 2499 2407 2503
rect 2411 2499 2412 2503
rect 2406 2498 2412 2499
rect 2582 2503 2588 2504
rect 2582 2499 2583 2503
rect 2587 2499 2588 2503
rect 2582 2498 2588 2499
rect 2750 2503 2756 2504
rect 2750 2499 2751 2503
rect 2755 2499 2756 2503
rect 2750 2498 2756 2499
rect 2910 2503 2916 2504
rect 2910 2499 2911 2503
rect 2915 2499 2916 2503
rect 2910 2498 2916 2499
rect 3062 2503 3068 2504
rect 3062 2499 3063 2503
rect 3067 2499 3068 2503
rect 3062 2498 3068 2499
rect 3206 2503 3212 2504
rect 3206 2499 3207 2503
rect 3211 2499 3212 2503
rect 3206 2498 3212 2499
rect 3350 2503 3356 2504
rect 3350 2499 3351 2503
rect 3355 2499 3356 2503
rect 3350 2498 3356 2499
rect 3486 2503 3492 2504
rect 3486 2499 3487 2503
rect 3491 2499 3492 2503
rect 3486 2498 3492 2499
rect 307 2495 313 2496
rect 307 2491 308 2495
rect 312 2494 313 2495
rect 338 2495 344 2496
rect 338 2494 339 2495
rect 312 2492 339 2494
rect 312 2491 313 2492
rect 307 2490 313 2491
rect 338 2491 339 2492
rect 343 2491 344 2495
rect 338 2490 344 2491
rect 494 2495 500 2496
rect 494 2491 495 2495
rect 499 2494 500 2495
rect 507 2495 513 2496
rect 507 2494 508 2495
rect 499 2492 508 2494
rect 499 2491 500 2492
rect 494 2490 500 2491
rect 507 2491 508 2492
rect 512 2491 513 2495
rect 507 2490 513 2491
rect 707 2495 713 2496
rect 707 2491 708 2495
rect 712 2494 713 2495
rect 839 2495 845 2496
rect 839 2494 840 2495
rect 712 2492 840 2494
rect 712 2491 713 2492
rect 707 2490 713 2491
rect 839 2491 840 2492
rect 844 2491 845 2495
rect 839 2490 845 2491
rect 847 2495 853 2496
rect 847 2491 848 2495
rect 852 2494 853 2495
rect 891 2495 897 2496
rect 891 2494 892 2495
rect 852 2492 892 2494
rect 852 2491 853 2492
rect 847 2490 853 2491
rect 891 2491 892 2492
rect 896 2491 897 2495
rect 891 2490 897 2491
rect 1059 2495 1068 2496
rect 1059 2491 1060 2495
rect 1067 2491 1068 2495
rect 1059 2490 1068 2491
rect 1158 2495 1164 2496
rect 1158 2491 1159 2495
rect 1163 2494 1164 2495
rect 1211 2495 1217 2496
rect 1211 2494 1212 2495
rect 1163 2492 1212 2494
rect 1163 2491 1164 2492
rect 1158 2490 1164 2491
rect 1211 2491 1212 2492
rect 1216 2491 1217 2495
rect 1211 2490 1217 2491
rect 1311 2495 1317 2496
rect 1311 2491 1312 2495
rect 1316 2494 1317 2495
rect 1355 2495 1361 2496
rect 1355 2494 1356 2495
rect 1316 2492 1356 2494
rect 1316 2491 1317 2492
rect 1311 2490 1317 2491
rect 1355 2491 1356 2492
rect 1360 2491 1361 2495
rect 1355 2490 1361 2491
rect 1491 2495 1497 2496
rect 1491 2491 1492 2495
rect 1496 2494 1497 2495
rect 1522 2495 1528 2496
rect 1522 2494 1523 2495
rect 1496 2492 1523 2494
rect 1496 2491 1497 2492
rect 1491 2490 1497 2491
rect 1522 2491 1523 2492
rect 1527 2491 1528 2495
rect 1522 2490 1528 2491
rect 1627 2495 1633 2496
rect 1627 2491 1628 2495
rect 1632 2494 1633 2495
rect 1658 2495 1664 2496
rect 1658 2494 1659 2495
rect 1632 2492 1659 2494
rect 1632 2491 1633 2492
rect 1627 2490 1633 2491
rect 1658 2491 1659 2492
rect 1663 2491 1664 2495
rect 1658 2490 1664 2491
rect 1762 2495 1769 2496
rect 1762 2491 1763 2495
rect 1768 2491 1769 2495
rect 1762 2490 1769 2491
rect 1923 2491 1929 2492
rect 1386 2487 1392 2488
rect 1386 2486 1387 2487
rect 1268 2484 1387 2486
rect 1268 2482 1270 2484
rect 1386 2483 1387 2484
rect 1391 2483 1392 2487
rect 1923 2487 1924 2491
rect 1928 2490 1929 2491
rect 1954 2491 1960 2492
rect 1954 2490 1955 2491
rect 1928 2488 1955 2490
rect 1928 2487 1929 2488
rect 1923 2486 1929 2487
rect 1954 2487 1955 2488
rect 1959 2487 1960 2491
rect 1954 2486 1960 2487
rect 2075 2491 2081 2492
rect 2075 2487 2076 2491
rect 2080 2490 2081 2491
rect 2106 2491 2112 2492
rect 2106 2490 2107 2491
rect 2080 2488 2107 2490
rect 2080 2487 2081 2488
rect 2075 2486 2081 2487
rect 2106 2487 2107 2488
rect 2111 2487 2112 2491
rect 2106 2486 2112 2487
rect 2251 2491 2257 2492
rect 2251 2487 2252 2491
rect 2256 2490 2257 2491
rect 2270 2491 2276 2492
rect 2270 2490 2271 2491
rect 2256 2488 2271 2490
rect 2256 2487 2257 2488
rect 2251 2486 2257 2487
rect 2270 2487 2271 2488
rect 2275 2487 2276 2491
rect 2270 2486 2276 2487
rect 2435 2491 2441 2492
rect 2435 2487 2436 2491
rect 2440 2490 2441 2491
rect 2530 2491 2536 2492
rect 2530 2490 2531 2491
rect 2440 2488 2531 2490
rect 2440 2487 2441 2488
rect 2435 2486 2441 2487
rect 2530 2487 2531 2488
rect 2535 2487 2536 2491
rect 2530 2486 2536 2487
rect 2567 2491 2573 2492
rect 2567 2487 2568 2491
rect 2572 2490 2573 2491
rect 2611 2491 2617 2492
rect 2611 2490 2612 2491
rect 2572 2488 2612 2490
rect 2572 2487 2573 2488
rect 2567 2486 2573 2487
rect 2611 2487 2612 2488
rect 2616 2487 2617 2491
rect 2611 2486 2617 2487
rect 2779 2491 2788 2492
rect 2779 2487 2780 2491
rect 2787 2487 2788 2491
rect 2779 2486 2788 2487
rect 2895 2491 2901 2492
rect 2895 2487 2896 2491
rect 2900 2490 2901 2491
rect 2939 2491 2945 2492
rect 2939 2490 2940 2491
rect 2900 2488 2940 2490
rect 2900 2487 2901 2488
rect 2895 2486 2901 2487
rect 2939 2487 2940 2488
rect 2944 2487 2945 2491
rect 2939 2486 2945 2487
rect 3047 2491 3053 2492
rect 3047 2487 3048 2491
rect 3052 2490 3053 2491
rect 3091 2491 3097 2492
rect 3091 2490 3092 2491
rect 3052 2488 3092 2490
rect 3052 2487 3053 2488
rect 3047 2486 3053 2487
rect 3091 2487 3092 2488
rect 3096 2487 3097 2491
rect 3091 2486 3097 2487
rect 3235 2491 3241 2492
rect 3235 2487 3236 2491
rect 3240 2490 3241 2491
rect 3266 2491 3272 2492
rect 3266 2490 3267 2491
rect 3240 2488 3267 2490
rect 3240 2487 3241 2488
rect 3235 2486 3241 2487
rect 3266 2487 3267 2488
rect 3271 2487 3272 2491
rect 3266 2486 3272 2487
rect 3367 2491 3373 2492
rect 3367 2487 3368 2491
rect 3372 2490 3373 2491
rect 3379 2491 3385 2492
rect 3379 2490 3380 2491
rect 3372 2488 3380 2490
rect 3372 2487 3373 2488
rect 3367 2486 3373 2487
rect 3379 2487 3380 2488
rect 3384 2487 3385 2491
rect 3379 2486 3385 2487
rect 3515 2491 3524 2492
rect 3515 2487 3516 2491
rect 3523 2487 3524 2491
rect 3515 2486 3524 2487
rect 1386 2482 1392 2483
rect 1267 2481 1273 2482
rect 211 2479 220 2480
rect 211 2475 212 2479
rect 219 2475 220 2479
rect 211 2474 220 2475
rect 302 2479 308 2480
rect 302 2475 303 2479
rect 307 2478 308 2479
rect 347 2479 353 2480
rect 347 2478 348 2479
rect 307 2476 348 2478
rect 307 2475 308 2476
rect 302 2474 308 2475
rect 347 2475 348 2476
rect 352 2475 353 2479
rect 347 2474 353 2475
rect 407 2479 413 2480
rect 407 2475 408 2479
rect 412 2478 413 2479
rect 491 2479 497 2480
rect 491 2478 492 2479
rect 412 2476 492 2478
rect 412 2475 413 2476
rect 407 2474 413 2475
rect 491 2475 492 2476
rect 496 2475 497 2479
rect 491 2474 497 2475
rect 567 2479 573 2480
rect 567 2475 568 2479
rect 572 2478 573 2479
rect 635 2479 641 2480
rect 635 2478 636 2479
rect 572 2476 636 2478
rect 572 2475 573 2476
rect 567 2474 573 2475
rect 635 2475 636 2476
rect 640 2475 641 2479
rect 635 2474 641 2475
rect 695 2479 701 2480
rect 695 2475 696 2479
rect 700 2478 701 2479
rect 771 2479 777 2480
rect 771 2478 772 2479
rect 700 2476 772 2478
rect 700 2475 701 2476
rect 695 2474 701 2475
rect 771 2475 772 2476
rect 776 2475 777 2479
rect 771 2474 777 2475
rect 831 2479 837 2480
rect 831 2475 832 2479
rect 836 2478 837 2479
rect 907 2479 913 2480
rect 907 2478 908 2479
rect 836 2476 908 2478
rect 836 2475 837 2476
rect 831 2474 837 2475
rect 907 2475 908 2476
rect 912 2475 913 2479
rect 907 2474 913 2475
rect 1035 2479 1041 2480
rect 1035 2475 1036 2479
rect 1040 2478 1041 2479
rect 1074 2479 1080 2480
rect 1074 2478 1075 2479
rect 1040 2476 1075 2478
rect 1040 2475 1041 2476
rect 1035 2474 1041 2475
rect 1074 2475 1075 2476
rect 1079 2475 1080 2479
rect 1074 2474 1080 2475
rect 1155 2479 1164 2480
rect 1155 2475 1156 2479
rect 1163 2475 1164 2479
rect 1267 2477 1268 2481
rect 1272 2477 1273 2481
rect 1267 2476 1273 2477
rect 1311 2479 1317 2480
rect 1155 2474 1164 2475
rect 1311 2475 1312 2479
rect 1316 2478 1317 2479
rect 1371 2479 1377 2480
rect 1371 2478 1372 2479
rect 1316 2476 1372 2478
rect 1316 2475 1317 2476
rect 1311 2474 1317 2475
rect 1371 2475 1372 2476
rect 1376 2475 1377 2479
rect 1371 2474 1377 2475
rect 1415 2479 1421 2480
rect 1415 2475 1416 2479
rect 1420 2478 1421 2479
rect 1475 2479 1481 2480
rect 1475 2478 1476 2479
rect 1420 2476 1476 2478
rect 1420 2475 1421 2476
rect 1415 2474 1421 2475
rect 1475 2475 1476 2476
rect 1480 2475 1481 2479
rect 1475 2474 1481 2475
rect 1519 2479 1525 2480
rect 1519 2475 1520 2479
rect 1524 2478 1525 2479
rect 1579 2479 1585 2480
rect 1579 2478 1580 2479
rect 1524 2476 1580 2478
rect 1524 2475 1525 2476
rect 1519 2474 1525 2475
rect 1579 2475 1580 2476
rect 1584 2475 1585 2479
rect 1579 2474 1585 2475
rect 1615 2479 1621 2480
rect 1615 2475 1616 2479
rect 1620 2478 1621 2479
rect 1675 2479 1681 2480
rect 1675 2478 1676 2479
rect 1620 2476 1676 2478
rect 1620 2475 1621 2476
rect 1615 2474 1621 2475
rect 1675 2475 1676 2476
rect 1680 2475 1681 2479
rect 1675 2474 1681 2475
rect 1711 2479 1717 2480
rect 1711 2475 1712 2479
rect 1716 2478 1717 2479
rect 1763 2479 1769 2480
rect 1763 2478 1764 2479
rect 1716 2476 1764 2478
rect 1716 2475 1717 2476
rect 1711 2474 1717 2475
rect 1763 2475 1764 2476
rect 1768 2475 1769 2479
rect 1763 2474 1769 2475
rect 1807 2479 1813 2480
rect 1807 2475 1808 2479
rect 1812 2478 1813 2479
rect 1923 2479 1929 2480
rect 1923 2478 1924 2479
rect 1812 2476 1924 2478
rect 1812 2475 1813 2476
rect 1807 2474 1813 2475
rect 1923 2475 1924 2476
rect 1928 2475 1929 2479
rect 1923 2474 1929 2475
rect 1959 2479 1965 2480
rect 1959 2475 1960 2479
rect 1964 2478 1965 2479
rect 2019 2479 2025 2480
rect 2019 2478 2020 2479
rect 1964 2476 2020 2478
rect 1964 2475 1965 2476
rect 1959 2474 1965 2475
rect 2019 2475 2020 2476
rect 2024 2475 2025 2479
rect 2019 2474 2025 2475
rect 2079 2479 2085 2480
rect 2079 2475 2080 2479
rect 2084 2478 2085 2479
rect 2155 2479 2161 2480
rect 2155 2478 2156 2479
rect 2084 2476 2156 2478
rect 2084 2475 2085 2476
rect 2079 2474 2085 2475
rect 2155 2475 2156 2476
rect 2160 2475 2161 2479
rect 2155 2474 2161 2475
rect 2215 2479 2221 2480
rect 2215 2475 2216 2479
rect 2220 2478 2221 2479
rect 2307 2479 2313 2480
rect 2307 2478 2308 2479
rect 2220 2476 2308 2478
rect 2220 2475 2221 2476
rect 2215 2474 2221 2475
rect 2307 2475 2308 2476
rect 2312 2475 2313 2479
rect 2307 2474 2313 2475
rect 2467 2479 2473 2480
rect 2467 2475 2468 2479
rect 2472 2478 2473 2479
rect 2538 2479 2544 2480
rect 2538 2478 2539 2479
rect 2472 2476 2539 2478
rect 2472 2475 2473 2476
rect 2467 2474 2473 2475
rect 2538 2475 2539 2476
rect 2543 2475 2544 2479
rect 2538 2474 2544 2475
rect 2627 2479 2633 2480
rect 2627 2475 2628 2479
rect 2632 2478 2633 2479
rect 2642 2479 2648 2480
rect 2642 2478 2643 2479
rect 2632 2476 2643 2478
rect 2632 2475 2633 2476
rect 2627 2474 2633 2475
rect 2642 2475 2643 2476
rect 2647 2475 2648 2479
rect 2642 2474 2648 2475
rect 2795 2479 2801 2480
rect 2795 2475 2796 2479
rect 2800 2478 2801 2479
rect 2874 2479 2880 2480
rect 2874 2478 2875 2479
rect 2800 2476 2875 2478
rect 2800 2475 2801 2476
rect 2795 2474 2801 2475
rect 2874 2475 2875 2476
rect 2879 2475 2880 2479
rect 2874 2474 2880 2475
rect 2971 2479 2977 2480
rect 2971 2475 2972 2479
rect 2976 2478 2977 2479
rect 3050 2479 3056 2480
rect 3050 2478 3051 2479
rect 2976 2476 3051 2478
rect 2976 2475 2977 2476
rect 2971 2474 2977 2475
rect 3050 2475 3051 2476
rect 3055 2475 3056 2479
rect 3050 2474 3056 2475
rect 3146 2479 3153 2480
rect 3146 2475 3147 2479
rect 3152 2475 3153 2479
rect 3146 2474 3153 2475
rect 3310 2479 3316 2480
rect 3310 2475 3311 2479
rect 3315 2478 3316 2479
rect 3323 2479 3329 2480
rect 3323 2478 3324 2479
rect 3315 2476 3324 2478
rect 3315 2475 3316 2476
rect 3310 2474 3316 2475
rect 3323 2475 3324 2476
rect 3328 2475 3329 2479
rect 3323 2474 3329 2475
rect 3499 2479 3505 2480
rect 3499 2475 3500 2479
rect 3504 2478 3505 2479
rect 3546 2479 3552 2480
rect 3546 2478 3547 2479
rect 3504 2476 3547 2478
rect 3504 2475 3505 2476
rect 3499 2474 3505 2475
rect 3546 2475 3547 2476
rect 3551 2475 3552 2479
rect 3546 2474 3552 2475
rect 182 2469 188 2470
rect 182 2465 183 2469
rect 187 2465 188 2469
rect 182 2464 188 2465
rect 318 2469 324 2470
rect 318 2465 319 2469
rect 323 2465 324 2469
rect 318 2464 324 2465
rect 462 2469 468 2470
rect 462 2465 463 2469
rect 467 2465 468 2469
rect 462 2464 468 2465
rect 606 2469 612 2470
rect 606 2465 607 2469
rect 611 2465 612 2469
rect 606 2464 612 2465
rect 742 2469 748 2470
rect 742 2465 743 2469
rect 747 2465 748 2469
rect 742 2464 748 2465
rect 878 2469 884 2470
rect 878 2465 879 2469
rect 883 2465 884 2469
rect 878 2464 884 2465
rect 1006 2469 1012 2470
rect 1006 2465 1007 2469
rect 1011 2465 1012 2469
rect 1006 2464 1012 2465
rect 1126 2469 1132 2470
rect 1126 2465 1127 2469
rect 1131 2465 1132 2469
rect 1126 2464 1132 2465
rect 1238 2469 1244 2470
rect 1238 2465 1239 2469
rect 1243 2465 1244 2469
rect 1238 2464 1244 2465
rect 1342 2469 1348 2470
rect 1342 2465 1343 2469
rect 1347 2465 1348 2469
rect 1342 2464 1348 2465
rect 1446 2469 1452 2470
rect 1446 2465 1447 2469
rect 1451 2465 1452 2469
rect 1446 2464 1452 2465
rect 1550 2469 1556 2470
rect 1550 2465 1551 2469
rect 1555 2465 1556 2469
rect 1550 2464 1556 2465
rect 1646 2469 1652 2470
rect 1646 2465 1647 2469
rect 1651 2465 1652 2469
rect 1646 2464 1652 2465
rect 1734 2469 1740 2470
rect 1734 2465 1735 2469
rect 1739 2465 1740 2469
rect 1734 2464 1740 2465
rect 1894 2469 1900 2470
rect 1894 2465 1895 2469
rect 1899 2465 1900 2469
rect 1894 2464 1900 2465
rect 1990 2469 1996 2470
rect 1990 2465 1991 2469
rect 1995 2465 1996 2469
rect 1990 2464 1996 2465
rect 2126 2469 2132 2470
rect 2126 2465 2127 2469
rect 2131 2465 2132 2469
rect 2126 2464 2132 2465
rect 2278 2469 2284 2470
rect 2278 2465 2279 2469
rect 2283 2465 2284 2469
rect 2278 2464 2284 2465
rect 2438 2469 2444 2470
rect 2438 2465 2439 2469
rect 2443 2465 2444 2469
rect 2438 2464 2444 2465
rect 2598 2469 2604 2470
rect 2598 2465 2599 2469
rect 2603 2465 2604 2469
rect 2598 2464 2604 2465
rect 2766 2469 2772 2470
rect 2766 2465 2767 2469
rect 2771 2465 2772 2469
rect 2766 2464 2772 2465
rect 2942 2469 2948 2470
rect 2942 2465 2943 2469
rect 2947 2465 2948 2469
rect 2942 2464 2948 2465
rect 3118 2469 3124 2470
rect 3118 2465 3119 2469
rect 3123 2465 3124 2469
rect 3118 2464 3124 2465
rect 3294 2469 3300 2470
rect 3294 2465 3295 2469
rect 3299 2465 3300 2469
rect 3294 2464 3300 2465
rect 3470 2469 3476 2470
rect 3470 2465 3471 2469
rect 3475 2465 3476 2469
rect 3470 2464 3476 2465
rect 1062 2463 1068 2464
rect 1062 2462 1063 2463
rect 1060 2459 1063 2462
rect 1067 2459 1068 2463
rect 1060 2458 1068 2459
rect 110 2456 116 2457
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 302 2455 308 2456
rect 302 2454 303 2455
rect 237 2452 303 2454
rect 110 2451 116 2452
rect 302 2451 303 2452
rect 307 2451 308 2455
rect 407 2455 413 2456
rect 407 2454 408 2455
rect 373 2452 408 2454
rect 302 2450 308 2451
rect 407 2451 408 2452
rect 412 2451 413 2455
rect 695 2455 701 2456
rect 695 2454 696 2455
rect 661 2452 696 2454
rect 407 2450 413 2451
rect 695 2451 696 2452
rect 700 2451 701 2455
rect 831 2455 837 2456
rect 831 2454 832 2455
rect 797 2452 832 2454
rect 695 2450 701 2451
rect 831 2451 832 2452
rect 836 2451 837 2455
rect 1060 2453 1062 2458
rect 1822 2456 1828 2457
rect 1311 2455 1317 2456
rect 1311 2454 1312 2455
rect 1293 2452 1312 2454
rect 831 2450 837 2451
rect 839 2451 845 2452
rect 839 2447 840 2451
rect 844 2450 845 2451
rect 1074 2451 1080 2452
rect 844 2448 897 2450
rect 844 2447 845 2448
rect 839 2446 845 2447
rect 1074 2447 1075 2451
rect 1079 2450 1080 2451
rect 1311 2451 1312 2452
rect 1316 2451 1317 2455
rect 1415 2455 1421 2456
rect 1415 2454 1416 2455
rect 1397 2452 1416 2454
rect 1311 2450 1317 2451
rect 1415 2451 1416 2452
rect 1420 2451 1421 2455
rect 1519 2455 1525 2456
rect 1519 2454 1520 2455
rect 1501 2452 1520 2454
rect 1415 2450 1421 2451
rect 1519 2451 1520 2452
rect 1524 2451 1525 2455
rect 1615 2455 1621 2456
rect 1615 2454 1616 2455
rect 1605 2452 1616 2454
rect 1519 2450 1525 2451
rect 1615 2451 1616 2452
rect 1620 2451 1621 2455
rect 1711 2455 1717 2456
rect 1711 2454 1712 2455
rect 1701 2452 1712 2454
rect 1615 2450 1621 2451
rect 1711 2451 1712 2452
rect 1716 2451 1717 2455
rect 1807 2455 1813 2456
rect 1807 2454 1808 2455
rect 1789 2452 1808 2454
rect 1711 2450 1717 2451
rect 1807 2451 1808 2452
rect 1812 2451 1813 2455
rect 1822 2452 1823 2456
rect 1827 2452 1828 2456
rect 1822 2451 1828 2452
rect 1862 2456 1868 2457
rect 3574 2456 3580 2457
rect 1862 2452 1863 2456
rect 1867 2452 1868 2456
rect 1959 2455 1965 2456
rect 1959 2454 1960 2455
rect 1949 2452 1960 2454
rect 1862 2451 1868 2452
rect 1959 2451 1960 2452
rect 1964 2451 1965 2455
rect 2079 2455 2085 2456
rect 2079 2454 2080 2455
rect 2045 2452 2080 2454
rect 1807 2450 1813 2451
rect 1959 2450 1965 2451
rect 2079 2451 2080 2452
rect 2084 2451 2085 2455
rect 2215 2455 2221 2456
rect 2215 2454 2216 2455
rect 2181 2452 2216 2454
rect 2079 2450 2085 2451
rect 2215 2451 2216 2452
rect 2220 2451 2221 2455
rect 3367 2455 3373 2456
rect 3367 2454 3368 2455
rect 3349 2452 3368 2454
rect 2215 2450 2221 2451
rect 2270 2451 2276 2452
rect 1079 2448 1145 2450
rect 1079 2447 1080 2448
rect 1074 2446 1080 2447
rect 2270 2447 2271 2451
rect 2275 2450 2276 2451
rect 2538 2451 2544 2452
rect 2275 2448 2297 2450
rect 2275 2447 2276 2448
rect 2270 2446 2276 2447
rect 2538 2447 2539 2451
rect 2543 2450 2544 2451
rect 2874 2451 2880 2452
rect 2543 2448 2617 2450
rect 2543 2447 2544 2448
rect 2538 2446 2544 2447
rect 2874 2447 2875 2451
rect 2879 2450 2880 2451
rect 3050 2451 3056 2452
rect 2879 2448 2961 2450
rect 2879 2447 2880 2448
rect 2874 2446 2880 2447
rect 3050 2447 3051 2451
rect 3055 2450 3056 2451
rect 3367 2451 3368 2452
rect 3372 2451 3373 2455
rect 3574 2452 3575 2456
rect 3579 2452 3580 2456
rect 3574 2451 3580 2452
rect 3367 2450 3373 2451
rect 3055 2448 3137 2450
rect 3055 2447 3056 2448
rect 3050 2446 3056 2447
rect 110 2439 116 2440
rect 110 2435 111 2439
rect 115 2435 116 2439
rect 110 2434 116 2435
rect 386 2439 392 2440
rect 386 2435 387 2439
rect 391 2438 392 2439
rect 1822 2439 1828 2440
rect 391 2436 473 2438
rect 391 2435 392 2436
rect 386 2434 392 2435
rect 1822 2435 1823 2439
rect 1827 2435 1828 2439
rect 1822 2434 1828 2435
rect 1862 2439 1868 2440
rect 1862 2435 1863 2439
rect 1867 2435 1868 2439
rect 1862 2434 1868 2435
rect 2390 2439 2396 2440
rect 2390 2435 2391 2439
rect 2395 2438 2396 2439
rect 2694 2439 2700 2440
rect 2395 2436 2449 2438
rect 2395 2435 2396 2436
rect 2390 2434 2396 2435
rect 2694 2435 2695 2439
rect 2699 2438 2700 2439
rect 3574 2439 3580 2440
rect 2699 2436 2777 2438
rect 2699 2435 2700 2436
rect 2694 2434 2700 2435
rect 3574 2435 3575 2439
rect 3579 2435 3580 2439
rect 3574 2434 3580 2435
rect 174 2429 180 2430
rect 174 2425 175 2429
rect 179 2425 180 2429
rect 174 2424 180 2425
rect 310 2429 316 2430
rect 310 2425 311 2429
rect 315 2425 316 2429
rect 310 2424 316 2425
rect 454 2429 460 2430
rect 454 2425 455 2429
rect 459 2425 460 2429
rect 454 2424 460 2425
rect 598 2429 604 2430
rect 598 2425 599 2429
rect 603 2425 604 2429
rect 598 2424 604 2425
rect 734 2429 740 2430
rect 734 2425 735 2429
rect 739 2425 740 2429
rect 734 2424 740 2425
rect 870 2429 876 2430
rect 870 2425 871 2429
rect 875 2425 876 2429
rect 870 2424 876 2425
rect 998 2429 1004 2430
rect 998 2425 999 2429
rect 1003 2425 1004 2429
rect 998 2424 1004 2425
rect 1118 2429 1124 2430
rect 1118 2425 1119 2429
rect 1123 2425 1124 2429
rect 1118 2424 1124 2425
rect 1230 2429 1236 2430
rect 1230 2425 1231 2429
rect 1235 2425 1236 2429
rect 1230 2424 1236 2425
rect 1334 2429 1340 2430
rect 1334 2425 1335 2429
rect 1339 2425 1340 2429
rect 1334 2424 1340 2425
rect 1438 2429 1444 2430
rect 1438 2425 1439 2429
rect 1443 2425 1444 2429
rect 1438 2424 1444 2425
rect 1542 2429 1548 2430
rect 1542 2425 1543 2429
rect 1547 2425 1548 2429
rect 1542 2424 1548 2425
rect 1638 2429 1644 2430
rect 1638 2425 1639 2429
rect 1643 2425 1644 2429
rect 1638 2424 1644 2425
rect 1726 2429 1732 2430
rect 1726 2425 1727 2429
rect 1731 2425 1732 2429
rect 1726 2424 1732 2425
rect 1886 2429 1892 2430
rect 1886 2425 1887 2429
rect 1891 2425 1892 2429
rect 1886 2424 1892 2425
rect 1982 2429 1988 2430
rect 1982 2425 1983 2429
rect 1987 2425 1988 2429
rect 1982 2424 1988 2425
rect 2118 2429 2124 2430
rect 2118 2425 2119 2429
rect 2123 2425 2124 2429
rect 2118 2424 2124 2425
rect 2270 2429 2276 2430
rect 2270 2425 2271 2429
rect 2275 2425 2276 2429
rect 2270 2424 2276 2425
rect 2430 2429 2436 2430
rect 2430 2425 2431 2429
rect 2435 2425 2436 2429
rect 2430 2424 2436 2425
rect 2590 2429 2596 2430
rect 2590 2425 2591 2429
rect 2595 2425 2596 2429
rect 2590 2424 2596 2425
rect 2758 2429 2764 2430
rect 2758 2425 2759 2429
rect 2763 2425 2764 2429
rect 2758 2424 2764 2425
rect 2934 2429 2940 2430
rect 2934 2425 2935 2429
rect 2939 2425 2940 2429
rect 2934 2424 2940 2425
rect 3110 2429 3116 2430
rect 3110 2425 3111 2429
rect 3115 2425 3116 2429
rect 3110 2424 3116 2425
rect 3286 2429 3292 2430
rect 3286 2425 3287 2429
rect 3291 2425 3292 2429
rect 3286 2424 3292 2425
rect 3462 2429 3468 2430
rect 3462 2425 3463 2429
rect 3467 2425 3468 2429
rect 3462 2424 3468 2425
rect 3510 2423 3517 2424
rect 3510 2419 3511 2423
rect 3516 2419 3517 2423
rect 3510 2418 3517 2419
rect 1158 2407 1164 2408
rect 1158 2403 1159 2407
rect 1163 2406 1164 2407
rect 1163 2404 1374 2406
rect 1163 2403 1164 2404
rect 1158 2402 1164 2403
rect 150 2399 156 2400
rect 150 2395 151 2399
rect 155 2395 156 2399
rect 150 2394 156 2395
rect 318 2399 324 2400
rect 318 2395 319 2399
rect 323 2395 324 2399
rect 318 2394 324 2395
rect 478 2399 484 2400
rect 478 2395 479 2399
rect 483 2395 484 2399
rect 478 2394 484 2395
rect 638 2399 644 2400
rect 638 2395 639 2399
rect 643 2395 644 2399
rect 638 2394 644 2395
rect 782 2399 788 2400
rect 782 2395 783 2399
rect 787 2395 788 2399
rect 782 2394 788 2395
rect 918 2399 924 2400
rect 918 2395 919 2399
rect 923 2395 924 2399
rect 918 2394 924 2395
rect 1046 2399 1052 2400
rect 1046 2395 1047 2399
rect 1051 2395 1052 2399
rect 1046 2394 1052 2395
rect 1174 2399 1180 2400
rect 1174 2395 1175 2399
rect 1179 2395 1180 2399
rect 1174 2394 1180 2395
rect 1302 2399 1308 2400
rect 1302 2395 1303 2399
rect 1307 2395 1308 2399
rect 1302 2394 1308 2395
rect 567 2391 573 2392
rect 567 2390 568 2391
rect 110 2389 116 2390
rect 110 2385 111 2389
rect 115 2385 116 2389
rect 537 2388 568 2390
rect 567 2387 568 2388
rect 572 2387 573 2391
rect 1372 2390 1374 2404
rect 1430 2399 1436 2400
rect 1430 2395 1431 2399
rect 1435 2395 1436 2399
rect 1430 2394 1436 2395
rect 2350 2399 2356 2400
rect 2350 2395 2351 2399
rect 2355 2395 2356 2399
rect 2350 2394 2356 2395
rect 2502 2399 2508 2400
rect 2502 2395 2503 2399
rect 2507 2395 2508 2399
rect 2502 2394 2508 2395
rect 2654 2399 2660 2400
rect 2654 2395 2655 2399
rect 2659 2395 2660 2399
rect 2654 2394 2660 2395
rect 2806 2399 2812 2400
rect 2806 2395 2807 2399
rect 2811 2395 2812 2399
rect 2806 2394 2812 2395
rect 2966 2399 2972 2400
rect 2966 2395 2967 2399
rect 2971 2395 2972 2399
rect 2966 2394 2972 2395
rect 3134 2399 3140 2400
rect 3134 2395 3135 2399
rect 3139 2395 3140 2399
rect 3134 2394 3140 2395
rect 3302 2399 3308 2400
rect 3302 2395 3303 2399
rect 3307 2395 3308 2399
rect 3302 2394 3308 2395
rect 3470 2399 3476 2400
rect 3470 2395 3471 2399
rect 3475 2395 3476 2399
rect 3470 2394 3476 2395
rect 1372 2388 1449 2390
rect 1822 2389 1828 2390
rect 567 2386 573 2387
rect 110 2384 116 2385
rect 1822 2385 1823 2389
rect 1827 2385 1828 2389
rect 1822 2384 1828 2385
rect 1862 2389 1868 2390
rect 1862 2385 1863 2389
rect 1867 2385 1868 2389
rect 3312 2388 3321 2390
rect 3574 2389 3580 2390
rect 1862 2384 1868 2385
rect 3310 2387 3316 2388
rect 3310 2383 3311 2387
rect 3315 2383 3316 2387
rect 3574 2385 3575 2389
rect 3579 2385 3580 2389
rect 3574 2384 3580 2385
rect 3310 2382 3316 2383
rect 2510 2379 2516 2380
rect 218 2375 224 2376
rect 218 2374 219 2375
rect 110 2372 116 2373
rect 213 2372 219 2374
rect 110 2368 111 2372
rect 115 2368 116 2372
rect 218 2371 219 2372
rect 223 2371 224 2375
rect 218 2370 224 2371
rect 226 2375 232 2376
rect 226 2371 227 2375
rect 231 2374 232 2375
rect 546 2375 552 2376
rect 231 2372 345 2374
rect 231 2371 232 2372
rect 226 2370 232 2371
rect 546 2371 547 2375
rect 551 2374 552 2375
rect 706 2375 712 2376
rect 551 2372 665 2374
rect 551 2371 552 2372
rect 546 2370 552 2371
rect 706 2371 707 2375
rect 711 2374 712 2375
rect 1039 2375 1045 2376
rect 1039 2374 1040 2375
rect 711 2372 809 2374
rect 981 2372 1040 2374
rect 711 2371 712 2372
rect 706 2370 712 2371
rect 1039 2371 1040 2372
rect 1044 2371 1045 2375
rect 1166 2375 1172 2376
rect 1166 2374 1167 2375
rect 1109 2372 1167 2374
rect 1039 2370 1045 2371
rect 1166 2371 1167 2372
rect 1171 2371 1172 2375
rect 1295 2375 1301 2376
rect 1295 2374 1296 2375
rect 1237 2372 1296 2374
rect 1166 2370 1172 2371
rect 1295 2371 1296 2372
rect 1300 2371 1301 2375
rect 1423 2375 1429 2376
rect 1423 2374 1424 2375
rect 1365 2372 1424 2374
rect 1295 2370 1301 2371
rect 1423 2371 1424 2372
rect 1428 2371 1429 2375
rect 2510 2375 2511 2379
rect 2515 2375 2516 2379
rect 2510 2374 2516 2375
rect 2586 2375 2592 2376
rect 2586 2374 2587 2375
rect 1423 2370 1429 2371
rect 1822 2372 1828 2373
rect 110 2367 116 2368
rect 1822 2368 1823 2372
rect 1827 2368 1828 2372
rect 1822 2367 1828 2368
rect 1862 2372 1868 2373
rect 2413 2372 2514 2374
rect 2565 2372 2587 2374
rect 1862 2368 1863 2372
rect 1867 2368 1868 2372
rect 2586 2371 2587 2372
rect 2591 2371 2592 2375
rect 2799 2375 2805 2376
rect 2799 2374 2800 2375
rect 2717 2372 2800 2374
rect 2586 2370 2592 2371
rect 2799 2371 2800 2372
rect 2804 2371 2805 2375
rect 2959 2375 2965 2376
rect 2959 2374 2960 2375
rect 2869 2372 2960 2374
rect 2799 2370 2805 2371
rect 2959 2371 2960 2372
rect 2964 2371 2965 2375
rect 3127 2375 3133 2376
rect 3127 2374 3128 2375
rect 3029 2372 3128 2374
rect 2959 2370 2965 2371
rect 3127 2371 3128 2372
rect 3132 2371 3133 2375
rect 3294 2375 3300 2376
rect 3294 2374 3295 2375
rect 3197 2372 3295 2374
rect 3127 2370 3133 2371
rect 3294 2371 3295 2372
rect 3299 2371 3300 2375
rect 3538 2375 3544 2376
rect 3538 2374 3539 2375
rect 3533 2372 3539 2374
rect 3294 2370 3300 2371
rect 3538 2371 3539 2372
rect 3543 2371 3544 2375
rect 3538 2370 3544 2371
rect 3574 2372 3580 2373
rect 1862 2367 1868 2368
rect 3574 2368 3575 2372
rect 3579 2368 3580 2372
rect 3574 2367 3580 2368
rect 158 2359 164 2360
rect 158 2355 159 2359
rect 163 2355 164 2359
rect 158 2354 164 2355
rect 326 2359 332 2360
rect 326 2355 327 2359
rect 331 2355 332 2359
rect 326 2354 332 2355
rect 486 2359 492 2360
rect 486 2355 487 2359
rect 491 2355 492 2359
rect 486 2354 492 2355
rect 646 2359 652 2360
rect 646 2355 647 2359
rect 651 2355 652 2359
rect 646 2354 652 2355
rect 790 2359 796 2360
rect 790 2355 791 2359
rect 795 2355 796 2359
rect 790 2354 796 2355
rect 926 2359 932 2360
rect 926 2355 927 2359
rect 931 2355 932 2359
rect 926 2354 932 2355
rect 1054 2359 1060 2360
rect 1054 2355 1055 2359
rect 1059 2355 1060 2359
rect 1054 2354 1060 2355
rect 1182 2359 1188 2360
rect 1182 2355 1183 2359
rect 1187 2355 1188 2359
rect 1182 2354 1188 2355
rect 1310 2359 1316 2360
rect 1310 2355 1311 2359
rect 1315 2355 1316 2359
rect 1310 2354 1316 2355
rect 1438 2359 1444 2360
rect 1438 2355 1439 2359
rect 1443 2355 1444 2359
rect 1438 2354 1444 2355
rect 2358 2359 2364 2360
rect 2358 2355 2359 2359
rect 2363 2355 2364 2359
rect 2358 2354 2364 2355
rect 2510 2359 2516 2360
rect 2510 2355 2511 2359
rect 2515 2355 2516 2359
rect 2510 2354 2516 2355
rect 2662 2359 2668 2360
rect 2662 2355 2663 2359
rect 2667 2355 2668 2359
rect 2662 2354 2668 2355
rect 2814 2359 2820 2360
rect 2814 2355 2815 2359
rect 2819 2355 2820 2359
rect 2814 2354 2820 2355
rect 2974 2359 2980 2360
rect 2974 2355 2975 2359
rect 2979 2355 2980 2359
rect 2974 2354 2980 2355
rect 3142 2359 3148 2360
rect 3142 2355 3143 2359
rect 3147 2355 3148 2359
rect 3142 2354 3148 2355
rect 3310 2359 3316 2360
rect 3310 2355 3311 2359
rect 3315 2355 3316 2359
rect 3310 2354 3316 2355
rect 3478 2359 3484 2360
rect 3478 2355 3479 2359
rect 3483 2355 3484 2359
rect 3478 2354 3484 2355
rect 187 2347 193 2348
rect 187 2343 188 2347
rect 192 2346 193 2347
rect 226 2347 232 2348
rect 226 2346 227 2347
rect 192 2344 227 2346
rect 192 2343 193 2344
rect 187 2342 193 2343
rect 226 2343 227 2344
rect 231 2343 232 2347
rect 226 2342 232 2343
rect 355 2347 361 2348
rect 355 2343 356 2347
rect 360 2346 361 2347
rect 386 2347 392 2348
rect 386 2346 387 2347
rect 360 2344 387 2346
rect 360 2343 361 2344
rect 355 2342 361 2343
rect 386 2343 387 2344
rect 391 2343 392 2347
rect 386 2342 392 2343
rect 515 2347 521 2348
rect 515 2343 516 2347
rect 520 2346 521 2347
rect 546 2347 552 2348
rect 546 2346 547 2347
rect 520 2344 547 2346
rect 520 2343 521 2344
rect 515 2342 521 2343
rect 546 2343 547 2344
rect 551 2343 552 2347
rect 546 2342 552 2343
rect 675 2347 681 2348
rect 675 2343 676 2347
rect 680 2346 681 2347
rect 706 2347 712 2348
rect 706 2346 707 2347
rect 680 2344 707 2346
rect 680 2343 681 2344
rect 675 2342 681 2343
rect 706 2343 707 2344
rect 711 2343 712 2347
rect 706 2342 712 2343
rect 751 2347 757 2348
rect 751 2343 752 2347
rect 756 2346 757 2347
rect 819 2347 825 2348
rect 819 2346 820 2347
rect 756 2344 820 2346
rect 756 2343 757 2344
rect 751 2342 757 2343
rect 819 2343 820 2344
rect 824 2343 825 2347
rect 819 2342 825 2343
rect 955 2347 961 2348
rect 955 2343 956 2347
rect 960 2346 961 2347
rect 1026 2347 1032 2348
rect 1026 2346 1027 2347
rect 960 2344 1027 2346
rect 960 2343 961 2344
rect 955 2342 961 2343
rect 1026 2343 1027 2344
rect 1031 2343 1032 2347
rect 1026 2342 1032 2343
rect 1039 2347 1045 2348
rect 1039 2343 1040 2347
rect 1044 2346 1045 2347
rect 1083 2347 1089 2348
rect 1083 2346 1084 2347
rect 1044 2344 1084 2346
rect 1044 2343 1045 2344
rect 1039 2342 1045 2343
rect 1083 2343 1084 2344
rect 1088 2343 1089 2347
rect 1083 2342 1089 2343
rect 1166 2347 1172 2348
rect 1166 2343 1167 2347
rect 1171 2346 1172 2347
rect 1211 2347 1217 2348
rect 1211 2346 1212 2347
rect 1171 2344 1212 2346
rect 1171 2343 1172 2344
rect 1166 2342 1172 2343
rect 1211 2343 1212 2344
rect 1216 2343 1217 2347
rect 1211 2342 1217 2343
rect 1295 2347 1301 2348
rect 1295 2343 1296 2347
rect 1300 2346 1301 2347
rect 1339 2347 1345 2348
rect 1339 2346 1340 2347
rect 1300 2344 1340 2346
rect 1300 2343 1301 2344
rect 1295 2342 1301 2343
rect 1339 2343 1340 2344
rect 1344 2343 1345 2347
rect 1339 2342 1345 2343
rect 1423 2347 1429 2348
rect 1423 2343 1424 2347
rect 1428 2346 1429 2347
rect 1467 2347 1473 2348
rect 1467 2346 1468 2347
rect 1428 2344 1468 2346
rect 1428 2343 1429 2344
rect 1423 2342 1429 2343
rect 1467 2343 1468 2344
rect 1472 2343 1473 2347
rect 1467 2342 1473 2343
rect 2387 2347 2396 2348
rect 2387 2343 2388 2347
rect 2395 2343 2396 2347
rect 2387 2342 2396 2343
rect 2538 2347 2545 2348
rect 2538 2343 2539 2347
rect 2544 2343 2545 2347
rect 2538 2342 2545 2343
rect 2691 2347 2700 2348
rect 2691 2343 2692 2347
rect 2699 2343 2700 2347
rect 2691 2342 2700 2343
rect 2799 2347 2805 2348
rect 2799 2343 2800 2347
rect 2804 2346 2805 2347
rect 2843 2347 2849 2348
rect 2843 2346 2844 2347
rect 2804 2344 2844 2346
rect 2804 2343 2805 2344
rect 2799 2342 2805 2343
rect 2843 2343 2844 2344
rect 2848 2343 2849 2347
rect 2843 2342 2849 2343
rect 2959 2347 2965 2348
rect 2959 2343 2960 2347
rect 2964 2346 2965 2347
rect 3003 2347 3009 2348
rect 3003 2346 3004 2347
rect 2964 2344 3004 2346
rect 2964 2343 2965 2344
rect 2959 2342 2965 2343
rect 3003 2343 3004 2344
rect 3008 2343 3009 2347
rect 3003 2342 3009 2343
rect 3127 2347 3133 2348
rect 3127 2343 3128 2347
rect 3132 2346 3133 2347
rect 3171 2347 3177 2348
rect 3171 2346 3172 2347
rect 3132 2344 3172 2346
rect 3132 2343 3133 2344
rect 3127 2342 3133 2343
rect 3171 2343 3172 2344
rect 3176 2343 3177 2347
rect 3171 2342 3177 2343
rect 3339 2347 3345 2348
rect 3339 2343 3340 2347
rect 3344 2346 3345 2347
rect 3370 2347 3376 2348
rect 3370 2346 3371 2347
rect 3344 2344 3371 2346
rect 3344 2343 3345 2344
rect 3339 2342 3345 2343
rect 3370 2343 3371 2344
rect 3375 2343 3376 2347
rect 3370 2342 3376 2343
rect 3507 2347 3516 2348
rect 3507 2343 3508 2347
rect 3515 2343 3516 2347
rect 3507 2342 3516 2343
rect 2958 2339 2964 2340
rect 2958 2338 2959 2339
rect 2732 2336 2959 2338
rect 2732 2334 2734 2336
rect 2958 2335 2959 2336
rect 2963 2335 2964 2339
rect 2958 2334 2964 2335
rect 2731 2333 2737 2334
rect 171 2331 177 2332
rect 171 2327 172 2331
rect 176 2330 177 2331
rect 218 2331 224 2332
rect 218 2330 219 2331
rect 176 2328 219 2330
rect 176 2327 177 2328
rect 171 2326 177 2327
rect 218 2327 219 2328
rect 223 2327 224 2331
rect 218 2326 224 2327
rect 231 2331 237 2332
rect 231 2327 232 2331
rect 236 2330 237 2331
rect 291 2331 297 2332
rect 291 2330 292 2331
rect 236 2328 292 2330
rect 236 2327 237 2328
rect 231 2326 237 2327
rect 291 2327 292 2328
rect 296 2327 297 2331
rect 291 2326 297 2327
rect 435 2331 444 2332
rect 435 2327 436 2331
rect 443 2327 444 2331
rect 435 2326 444 2327
rect 495 2331 501 2332
rect 495 2327 496 2331
rect 500 2330 501 2331
rect 571 2331 577 2332
rect 571 2330 572 2331
rect 500 2328 572 2330
rect 500 2327 501 2328
rect 495 2326 501 2327
rect 571 2327 572 2328
rect 576 2327 577 2331
rect 571 2326 577 2327
rect 631 2331 637 2332
rect 631 2327 632 2331
rect 636 2330 637 2331
rect 707 2331 713 2332
rect 707 2330 708 2331
rect 636 2328 708 2330
rect 636 2327 637 2328
rect 631 2326 637 2327
rect 707 2327 708 2328
rect 712 2327 713 2331
rect 707 2326 713 2327
rect 783 2331 789 2332
rect 783 2327 784 2331
rect 788 2330 789 2331
rect 835 2331 841 2332
rect 835 2330 836 2331
rect 788 2328 836 2330
rect 788 2327 789 2328
rect 783 2326 789 2327
rect 835 2327 836 2328
rect 840 2327 841 2331
rect 835 2326 841 2327
rect 887 2331 893 2332
rect 887 2327 888 2331
rect 892 2330 893 2331
rect 955 2331 961 2332
rect 955 2330 956 2331
rect 892 2328 956 2330
rect 892 2327 893 2328
rect 887 2326 893 2327
rect 955 2327 956 2328
rect 960 2327 961 2331
rect 955 2326 961 2327
rect 999 2331 1005 2332
rect 999 2327 1000 2331
rect 1004 2330 1005 2331
rect 1067 2331 1073 2332
rect 1067 2330 1068 2331
rect 1004 2328 1068 2330
rect 1004 2327 1005 2328
rect 999 2326 1005 2327
rect 1067 2327 1068 2328
rect 1072 2327 1073 2331
rect 1067 2326 1073 2327
rect 1102 2331 1108 2332
rect 1102 2327 1103 2331
rect 1107 2330 1108 2331
rect 1187 2331 1193 2332
rect 1187 2330 1188 2331
rect 1107 2328 1188 2330
rect 1107 2327 1108 2328
rect 1102 2326 1108 2327
rect 1187 2327 1188 2328
rect 1192 2327 1193 2331
rect 1187 2326 1193 2327
rect 1218 2331 1224 2332
rect 1218 2327 1219 2331
rect 1223 2330 1224 2331
rect 1307 2331 1313 2332
rect 1307 2330 1308 2331
rect 1223 2328 1308 2330
rect 1223 2327 1224 2328
rect 1218 2326 1224 2327
rect 1307 2327 1308 2328
rect 1312 2327 1313 2331
rect 1307 2326 1313 2327
rect 2379 2331 2385 2332
rect 2379 2327 2380 2331
rect 2384 2330 2385 2331
rect 2418 2331 2424 2332
rect 2418 2330 2419 2331
rect 2384 2328 2419 2330
rect 2384 2327 2385 2328
rect 2379 2326 2385 2327
rect 2418 2327 2419 2328
rect 2423 2327 2424 2331
rect 2418 2326 2424 2327
rect 2475 2331 2481 2332
rect 2475 2327 2476 2331
rect 2480 2330 2481 2331
rect 2522 2331 2528 2332
rect 2522 2330 2523 2331
rect 2480 2328 2523 2330
rect 2480 2327 2481 2328
rect 2475 2326 2481 2327
rect 2522 2327 2523 2328
rect 2527 2327 2528 2331
rect 2522 2326 2528 2327
rect 2586 2331 2593 2332
rect 2586 2327 2587 2331
rect 2592 2327 2593 2331
rect 2731 2329 2732 2333
rect 2736 2329 2737 2333
rect 2731 2328 2737 2329
rect 2839 2331 2845 2332
rect 2586 2326 2593 2327
rect 2839 2327 2840 2331
rect 2844 2330 2845 2331
rect 2907 2331 2913 2332
rect 2907 2330 2908 2331
rect 2844 2328 2908 2330
rect 2844 2327 2845 2328
rect 2839 2326 2845 2327
rect 2907 2327 2908 2328
rect 2912 2327 2913 2331
rect 2907 2326 2913 2327
rect 3107 2331 3113 2332
rect 3107 2327 3108 2331
rect 3112 2330 3113 2331
rect 3150 2331 3156 2332
rect 3150 2330 3151 2331
rect 3112 2328 3151 2330
rect 3112 2327 3113 2328
rect 3107 2326 3113 2327
rect 3150 2327 3151 2328
rect 3155 2327 3156 2331
rect 3150 2326 3156 2327
rect 3294 2331 3300 2332
rect 3294 2327 3295 2331
rect 3299 2330 3300 2331
rect 3315 2331 3321 2332
rect 3315 2330 3316 2331
rect 3299 2328 3316 2330
rect 3299 2327 3300 2328
rect 3294 2326 3300 2327
rect 3315 2327 3316 2328
rect 3320 2327 3321 2331
rect 3315 2326 3321 2327
rect 3515 2331 3521 2332
rect 3515 2327 3516 2331
rect 3520 2330 3521 2331
rect 3538 2331 3544 2332
rect 3538 2330 3539 2331
rect 3520 2328 3539 2330
rect 3520 2327 3521 2328
rect 3515 2326 3521 2327
rect 3538 2327 3539 2328
rect 3543 2327 3544 2331
rect 3538 2326 3544 2327
rect 142 2321 148 2322
rect 142 2317 143 2321
rect 147 2317 148 2321
rect 142 2316 148 2317
rect 262 2321 268 2322
rect 262 2317 263 2321
rect 267 2317 268 2321
rect 262 2316 268 2317
rect 406 2321 412 2322
rect 406 2317 407 2321
rect 411 2317 412 2321
rect 406 2316 412 2317
rect 542 2321 548 2322
rect 542 2317 543 2321
rect 547 2317 548 2321
rect 542 2316 548 2317
rect 678 2321 684 2322
rect 678 2317 679 2321
rect 683 2317 684 2321
rect 678 2316 684 2317
rect 806 2321 812 2322
rect 806 2317 807 2321
rect 811 2317 812 2321
rect 806 2316 812 2317
rect 926 2321 932 2322
rect 926 2317 927 2321
rect 931 2317 932 2321
rect 926 2316 932 2317
rect 1038 2321 1044 2322
rect 1038 2317 1039 2321
rect 1043 2317 1044 2321
rect 1038 2316 1044 2317
rect 1158 2321 1164 2322
rect 1158 2317 1159 2321
rect 1163 2317 1164 2321
rect 1158 2316 1164 2317
rect 1278 2321 1284 2322
rect 1278 2317 1279 2321
rect 1283 2317 1284 2321
rect 1278 2316 1284 2317
rect 2350 2321 2356 2322
rect 2350 2317 2351 2321
rect 2355 2317 2356 2321
rect 2350 2316 2356 2317
rect 2446 2321 2452 2322
rect 2446 2317 2447 2321
rect 2451 2317 2452 2321
rect 2446 2316 2452 2317
rect 2558 2321 2564 2322
rect 2558 2317 2559 2321
rect 2563 2317 2564 2321
rect 2558 2316 2564 2317
rect 2702 2321 2708 2322
rect 2702 2317 2703 2321
rect 2707 2317 2708 2321
rect 2702 2316 2708 2317
rect 2878 2321 2884 2322
rect 2878 2317 2879 2321
rect 2883 2317 2884 2321
rect 2878 2316 2884 2317
rect 3078 2321 3084 2322
rect 3078 2317 3079 2321
rect 3083 2317 3084 2321
rect 3078 2316 3084 2317
rect 3286 2321 3292 2322
rect 3286 2317 3287 2321
rect 3291 2317 3292 2321
rect 3286 2316 3292 2317
rect 3486 2321 3492 2322
rect 3486 2317 3487 2321
rect 3491 2317 3492 2321
rect 3486 2316 3492 2317
rect 110 2308 116 2309
rect 1822 2308 1828 2309
rect 110 2304 111 2308
rect 115 2304 116 2308
rect 231 2307 237 2308
rect 231 2306 232 2307
rect 197 2304 232 2306
rect 110 2303 116 2304
rect 231 2303 232 2304
rect 236 2303 237 2307
rect 495 2307 501 2308
rect 495 2306 496 2307
rect 461 2304 496 2306
rect 231 2302 237 2303
rect 495 2303 496 2304
rect 500 2303 501 2307
rect 631 2307 637 2308
rect 631 2306 632 2307
rect 597 2304 632 2306
rect 495 2302 501 2303
rect 631 2303 632 2304
rect 636 2303 637 2307
rect 751 2307 757 2308
rect 751 2306 752 2307
rect 733 2304 752 2306
rect 631 2302 637 2303
rect 751 2303 752 2304
rect 756 2303 757 2307
rect 887 2307 893 2308
rect 887 2306 888 2307
rect 861 2304 888 2306
rect 751 2302 757 2303
rect 887 2303 888 2304
rect 892 2303 893 2307
rect 999 2307 1005 2308
rect 999 2306 1000 2307
rect 981 2304 1000 2306
rect 887 2302 893 2303
rect 999 2303 1000 2304
rect 1004 2303 1005 2307
rect 1102 2307 1108 2308
rect 1102 2306 1103 2307
rect 1093 2304 1103 2306
rect 999 2302 1005 2303
rect 1102 2303 1103 2304
rect 1107 2303 1108 2307
rect 1218 2307 1224 2308
rect 1218 2306 1219 2307
rect 1213 2304 1219 2306
rect 1102 2302 1108 2303
rect 1218 2303 1219 2304
rect 1223 2303 1224 2307
rect 1822 2304 1823 2308
rect 1827 2304 1828 2308
rect 1218 2302 1224 2303
rect 1226 2303 1232 2304
rect 1822 2303 1828 2304
rect 1862 2308 1868 2309
rect 3574 2308 3580 2309
rect 1862 2304 1863 2308
rect 1867 2304 1868 2308
rect 2839 2307 2845 2308
rect 2839 2306 2840 2307
rect 2757 2304 2840 2306
rect 1862 2303 1868 2304
rect 2418 2303 2424 2304
rect 1226 2299 1227 2303
rect 1231 2302 1232 2303
rect 1231 2300 1297 2302
rect 1231 2299 1232 2300
rect 1226 2298 1232 2299
rect 2418 2299 2419 2303
rect 2423 2302 2424 2303
rect 2522 2303 2528 2304
rect 2423 2300 2465 2302
rect 2423 2299 2424 2300
rect 2418 2298 2424 2299
rect 2522 2299 2523 2303
rect 2527 2302 2528 2303
rect 2839 2303 2840 2304
rect 2844 2303 2845 2307
rect 3574 2304 3575 2308
rect 3579 2304 3580 2308
rect 2839 2302 2845 2303
rect 2958 2303 2964 2304
rect 2527 2300 2577 2302
rect 2527 2299 2528 2300
rect 2522 2298 2528 2299
rect 2958 2299 2959 2303
rect 2963 2302 2964 2303
rect 3150 2303 3156 2304
rect 3574 2303 3580 2304
rect 2963 2300 3097 2302
rect 2963 2299 2964 2300
rect 2958 2298 2964 2299
rect 3150 2299 3151 2303
rect 3155 2302 3156 2303
rect 3155 2300 3305 2302
rect 3155 2299 3156 2300
rect 3150 2298 3156 2299
rect 110 2291 116 2292
rect 110 2287 111 2291
rect 115 2287 116 2291
rect 386 2291 392 2292
rect 386 2290 387 2291
rect 313 2288 387 2290
rect 110 2286 116 2287
rect 386 2287 387 2288
rect 391 2287 392 2291
rect 386 2286 392 2287
rect 1822 2291 1828 2292
rect 1822 2287 1823 2291
rect 1827 2287 1828 2291
rect 1822 2286 1828 2287
rect 1862 2291 1868 2292
rect 1862 2287 1863 2291
rect 1867 2287 1868 2291
rect 2946 2291 2952 2292
rect 2946 2290 2947 2291
rect 2929 2288 2947 2290
rect 1862 2286 1868 2287
rect 2946 2287 2947 2288
rect 2951 2287 2952 2291
rect 2946 2286 2952 2287
rect 3574 2291 3580 2292
rect 3574 2287 3575 2291
rect 3579 2287 3580 2291
rect 3574 2286 3580 2287
rect 134 2281 140 2282
rect 134 2277 135 2281
rect 139 2277 140 2281
rect 134 2276 140 2277
rect 254 2281 260 2282
rect 254 2277 255 2281
rect 259 2277 260 2281
rect 254 2276 260 2277
rect 398 2281 404 2282
rect 398 2277 399 2281
rect 403 2277 404 2281
rect 398 2276 404 2277
rect 534 2281 540 2282
rect 534 2277 535 2281
rect 539 2277 540 2281
rect 534 2276 540 2277
rect 670 2281 676 2282
rect 670 2277 671 2281
rect 675 2277 676 2281
rect 670 2276 676 2277
rect 798 2281 804 2282
rect 798 2277 799 2281
rect 803 2277 804 2281
rect 798 2276 804 2277
rect 918 2281 924 2282
rect 918 2277 919 2281
rect 923 2277 924 2281
rect 918 2276 924 2277
rect 1030 2281 1036 2282
rect 1030 2277 1031 2281
rect 1035 2277 1036 2281
rect 1030 2276 1036 2277
rect 1150 2281 1156 2282
rect 1150 2277 1151 2281
rect 1155 2277 1156 2281
rect 1150 2276 1156 2277
rect 1270 2281 1276 2282
rect 1270 2277 1271 2281
rect 1275 2277 1276 2281
rect 1270 2276 1276 2277
rect 2342 2281 2348 2282
rect 2342 2277 2343 2281
rect 2347 2277 2348 2281
rect 2342 2276 2348 2277
rect 2438 2281 2444 2282
rect 2438 2277 2439 2281
rect 2443 2277 2444 2281
rect 2438 2276 2444 2277
rect 2550 2281 2556 2282
rect 2550 2277 2551 2281
rect 2555 2277 2556 2281
rect 2550 2276 2556 2277
rect 2694 2281 2700 2282
rect 2694 2277 2695 2281
rect 2699 2277 2700 2281
rect 2694 2276 2700 2277
rect 2870 2281 2876 2282
rect 2870 2277 2871 2281
rect 2875 2277 2876 2281
rect 2870 2276 2876 2277
rect 3070 2281 3076 2282
rect 3070 2277 3071 2281
rect 3075 2277 3076 2281
rect 3070 2276 3076 2277
rect 3278 2281 3284 2282
rect 3278 2277 3279 2281
rect 3283 2277 3284 2281
rect 3278 2276 3284 2277
rect 3478 2281 3484 2282
rect 3478 2277 3479 2281
rect 3483 2277 3484 2281
rect 3478 2276 3484 2277
rect 2374 2275 2380 2276
rect 2374 2271 2375 2275
rect 2379 2274 2380 2275
rect 2391 2275 2397 2276
rect 2391 2274 2392 2275
rect 2379 2272 2392 2274
rect 2379 2271 2380 2272
rect 2374 2270 2380 2271
rect 2391 2271 2392 2272
rect 2396 2271 2397 2275
rect 2391 2270 2397 2271
rect 3518 2275 3524 2276
rect 3518 2271 3519 2275
rect 3523 2274 3524 2275
rect 3527 2275 3533 2276
rect 3527 2274 3528 2275
rect 3523 2272 3528 2274
rect 3523 2271 3524 2272
rect 3518 2270 3524 2271
rect 3527 2271 3528 2272
rect 3532 2271 3533 2275
rect 3527 2270 3533 2271
rect 134 2259 140 2260
rect 134 2255 135 2259
rect 139 2255 140 2259
rect 134 2254 140 2255
rect 230 2259 236 2260
rect 230 2255 231 2259
rect 235 2255 236 2259
rect 230 2254 236 2255
rect 350 2259 356 2260
rect 350 2255 351 2259
rect 355 2255 356 2259
rect 350 2254 356 2255
rect 470 2259 476 2260
rect 470 2255 471 2259
rect 475 2255 476 2259
rect 470 2254 476 2255
rect 590 2259 596 2260
rect 590 2255 591 2259
rect 595 2255 596 2259
rect 590 2254 596 2255
rect 710 2259 716 2260
rect 710 2255 711 2259
rect 715 2255 716 2259
rect 710 2254 716 2255
rect 822 2259 828 2260
rect 822 2255 823 2259
rect 827 2255 828 2259
rect 822 2254 828 2255
rect 934 2259 940 2260
rect 934 2255 935 2259
rect 939 2255 940 2259
rect 934 2254 940 2255
rect 1054 2259 1060 2260
rect 1054 2255 1055 2259
rect 1059 2255 1060 2259
rect 1054 2254 1060 2255
rect 1174 2259 1180 2260
rect 1174 2255 1175 2259
rect 1179 2255 1180 2259
rect 1174 2254 1180 2255
rect 2334 2259 2340 2260
rect 2334 2255 2335 2259
rect 2339 2255 2340 2259
rect 2334 2254 2340 2255
rect 2446 2259 2452 2260
rect 2446 2255 2447 2259
rect 2451 2255 2452 2259
rect 2446 2254 2452 2255
rect 2582 2259 2588 2260
rect 2582 2255 2583 2259
rect 2587 2255 2588 2259
rect 2582 2254 2588 2255
rect 2734 2259 2740 2260
rect 2734 2255 2735 2259
rect 2739 2255 2740 2259
rect 2734 2254 2740 2255
rect 2910 2259 2916 2260
rect 2910 2255 2911 2259
rect 2915 2255 2916 2259
rect 2910 2254 2916 2255
rect 3102 2259 3108 2260
rect 3102 2255 3103 2259
rect 3107 2255 3108 2259
rect 3102 2254 3108 2255
rect 3302 2259 3308 2260
rect 3302 2255 3303 2259
rect 3307 2255 3308 2259
rect 3302 2254 3308 2255
rect 3478 2259 3484 2260
rect 3478 2255 3479 2259
rect 3483 2255 3484 2259
rect 3478 2254 3484 2255
rect 438 2251 444 2252
rect 110 2249 116 2250
rect 110 2245 111 2249
rect 115 2245 116 2249
rect 438 2247 439 2251
rect 443 2250 444 2251
rect 783 2251 789 2252
rect 783 2250 784 2251
rect 443 2248 489 2250
rect 769 2248 784 2250
rect 443 2247 444 2248
rect 438 2246 444 2247
rect 783 2247 784 2248
rect 788 2247 789 2251
rect 3370 2251 3376 2252
rect 3370 2250 3371 2251
rect 783 2246 789 2247
rect 1822 2249 1828 2250
rect 110 2244 116 2245
rect 1822 2245 1823 2249
rect 1827 2245 1828 2249
rect 1822 2244 1828 2245
rect 1862 2249 1868 2250
rect 1862 2245 1863 2249
rect 1867 2245 1868 2249
rect 3361 2248 3371 2250
rect 3370 2247 3371 2248
rect 3375 2247 3376 2251
rect 3370 2246 3376 2247
rect 3574 2249 3580 2250
rect 1862 2244 1868 2245
rect 3574 2245 3575 2249
rect 3579 2245 3580 2249
rect 3574 2244 3580 2245
rect 127 2235 133 2236
rect 110 2232 116 2233
rect 110 2228 111 2232
rect 115 2228 116 2232
rect 127 2231 128 2235
rect 132 2234 133 2235
rect 202 2235 208 2236
rect 132 2232 161 2234
rect 132 2231 133 2232
rect 127 2230 133 2231
rect 202 2231 203 2235
rect 207 2234 208 2235
rect 298 2235 304 2236
rect 207 2232 257 2234
rect 207 2231 208 2232
rect 202 2230 208 2231
rect 298 2231 299 2235
rect 303 2234 304 2235
rect 538 2235 544 2236
rect 303 2232 377 2234
rect 303 2231 304 2232
rect 298 2230 304 2231
rect 538 2231 539 2235
rect 543 2234 544 2235
rect 778 2235 784 2236
rect 543 2232 617 2234
rect 543 2231 544 2232
rect 538 2230 544 2231
rect 778 2231 779 2235
rect 783 2234 784 2235
rect 1047 2235 1053 2236
rect 1047 2234 1048 2235
rect 783 2232 849 2234
rect 997 2232 1048 2234
rect 783 2231 784 2232
rect 778 2230 784 2231
rect 1047 2231 1048 2232
rect 1052 2231 1053 2235
rect 1138 2235 1144 2236
rect 1138 2234 1139 2235
rect 1117 2232 1139 2234
rect 1047 2230 1053 2231
rect 1138 2231 1139 2232
rect 1143 2231 1144 2235
rect 1138 2230 1144 2231
rect 1146 2235 1152 2236
rect 1146 2231 1147 2235
rect 1151 2234 1152 2235
rect 2439 2235 2445 2236
rect 2439 2234 2440 2235
rect 1151 2232 1201 2234
rect 1822 2232 1828 2233
rect 1151 2231 1152 2232
rect 1146 2230 1152 2231
rect 110 2227 116 2228
rect 1822 2228 1823 2232
rect 1827 2228 1828 2232
rect 1822 2227 1828 2228
rect 1862 2232 1868 2233
rect 2397 2232 2440 2234
rect 1862 2228 1863 2232
rect 1867 2228 1868 2232
rect 2439 2231 2440 2232
rect 2444 2231 2445 2235
rect 2566 2235 2572 2236
rect 2566 2234 2567 2235
rect 2509 2232 2567 2234
rect 2439 2230 2445 2231
rect 2566 2231 2567 2232
rect 2571 2231 2572 2235
rect 2566 2230 2572 2231
rect 2574 2235 2580 2236
rect 2574 2231 2575 2235
rect 2579 2234 2580 2235
rect 2726 2235 2732 2236
rect 2579 2232 2609 2234
rect 2579 2231 2580 2232
rect 2574 2230 2580 2231
rect 2726 2231 2727 2235
rect 2731 2234 2732 2235
rect 3014 2235 3020 2236
rect 3014 2234 3015 2235
rect 2731 2232 2761 2234
rect 2973 2232 3015 2234
rect 2731 2231 2732 2232
rect 2726 2230 2732 2231
rect 3014 2231 3015 2232
rect 3019 2231 3020 2235
rect 3014 2230 3020 2231
rect 3022 2235 3028 2236
rect 3022 2231 3023 2235
rect 3027 2234 3028 2235
rect 3546 2235 3552 2236
rect 3546 2234 3547 2235
rect 3027 2232 3129 2234
rect 3541 2232 3547 2234
rect 3027 2231 3028 2232
rect 3022 2230 3028 2231
rect 3546 2231 3547 2232
rect 3551 2231 3552 2235
rect 3546 2230 3552 2231
rect 3574 2232 3580 2233
rect 1862 2227 1868 2228
rect 3574 2228 3575 2232
rect 3579 2228 3580 2232
rect 3574 2227 3580 2228
rect 142 2219 148 2220
rect 142 2215 143 2219
rect 147 2215 148 2219
rect 142 2214 148 2215
rect 238 2219 244 2220
rect 238 2215 239 2219
rect 243 2215 244 2219
rect 238 2214 244 2215
rect 358 2219 364 2220
rect 358 2215 359 2219
rect 363 2215 364 2219
rect 358 2214 364 2215
rect 478 2219 484 2220
rect 478 2215 479 2219
rect 483 2215 484 2219
rect 478 2214 484 2215
rect 598 2219 604 2220
rect 598 2215 599 2219
rect 603 2215 604 2219
rect 598 2214 604 2215
rect 718 2219 724 2220
rect 718 2215 719 2219
rect 723 2215 724 2219
rect 718 2214 724 2215
rect 830 2219 836 2220
rect 830 2215 831 2219
rect 835 2215 836 2219
rect 830 2214 836 2215
rect 942 2219 948 2220
rect 942 2215 943 2219
rect 947 2215 948 2219
rect 942 2214 948 2215
rect 1062 2219 1068 2220
rect 1062 2215 1063 2219
rect 1067 2215 1068 2219
rect 1182 2219 1188 2220
rect 1062 2214 1068 2215
rect 1146 2215 1152 2216
rect 1146 2214 1147 2215
rect 952 2212 1058 2214
rect 952 2210 954 2212
rect 859 2209 954 2210
rect 171 2207 177 2208
rect 171 2203 172 2207
rect 176 2206 177 2207
rect 202 2207 208 2208
rect 202 2206 203 2207
rect 176 2204 203 2206
rect 176 2203 177 2204
rect 171 2202 177 2203
rect 202 2203 203 2204
rect 207 2203 208 2207
rect 202 2202 208 2203
rect 267 2207 273 2208
rect 267 2203 268 2207
rect 272 2206 273 2207
rect 298 2207 304 2208
rect 298 2206 299 2207
rect 272 2204 299 2206
rect 272 2203 273 2204
rect 267 2202 273 2203
rect 298 2203 299 2204
rect 303 2203 304 2207
rect 298 2202 304 2203
rect 386 2207 393 2208
rect 386 2203 387 2207
rect 392 2203 393 2207
rect 386 2202 393 2203
rect 507 2207 513 2208
rect 507 2203 508 2207
rect 512 2206 513 2207
rect 538 2207 544 2208
rect 538 2206 539 2207
rect 512 2204 539 2206
rect 512 2203 513 2204
rect 507 2202 513 2203
rect 538 2203 539 2204
rect 543 2203 544 2207
rect 538 2202 544 2203
rect 627 2207 636 2208
rect 627 2203 628 2207
rect 635 2203 636 2207
rect 627 2202 636 2203
rect 747 2207 753 2208
rect 747 2203 748 2207
rect 752 2206 753 2207
rect 778 2207 784 2208
rect 778 2206 779 2207
rect 752 2204 779 2206
rect 752 2203 753 2204
rect 747 2202 753 2203
rect 778 2203 779 2204
rect 783 2203 784 2207
rect 859 2205 860 2209
rect 864 2208 954 2209
rect 1056 2210 1058 2212
rect 1072 2212 1147 2214
rect 1072 2210 1074 2212
rect 1146 2211 1147 2212
rect 1151 2211 1152 2215
rect 1182 2215 1183 2219
rect 1187 2215 1188 2219
rect 1182 2214 1188 2215
rect 2342 2219 2348 2220
rect 2342 2215 2343 2219
rect 2347 2215 2348 2219
rect 2342 2214 2348 2215
rect 2454 2219 2460 2220
rect 2454 2215 2455 2219
rect 2459 2215 2460 2219
rect 2454 2214 2460 2215
rect 2590 2219 2596 2220
rect 2590 2215 2591 2219
rect 2595 2215 2596 2219
rect 2590 2214 2596 2215
rect 2742 2219 2748 2220
rect 2742 2215 2743 2219
rect 2747 2215 2748 2219
rect 2742 2214 2748 2215
rect 2918 2219 2924 2220
rect 2918 2215 2919 2219
rect 2923 2215 2924 2219
rect 3110 2219 3116 2220
rect 2918 2214 2924 2215
rect 3022 2215 3028 2216
rect 3022 2214 3023 2215
rect 1146 2210 1152 2211
rect 2940 2212 3023 2214
rect 2940 2210 2942 2212
rect 3022 2211 3023 2212
rect 3027 2211 3028 2215
rect 3110 2215 3111 2219
rect 3115 2215 3116 2219
rect 3110 2214 3116 2215
rect 3310 2219 3316 2220
rect 3310 2215 3311 2219
rect 3315 2215 3316 2219
rect 3310 2214 3316 2215
rect 3486 2219 3492 2220
rect 3486 2215 3487 2219
rect 3491 2215 3492 2219
rect 3486 2214 3492 2215
rect 3022 2210 3028 2211
rect 1056 2208 1074 2210
rect 2771 2209 2942 2210
rect 864 2205 865 2208
rect 859 2204 865 2205
rect 970 2207 977 2208
rect 778 2202 784 2203
rect 970 2203 971 2207
rect 976 2203 977 2207
rect 970 2202 977 2203
rect 1047 2207 1053 2208
rect 1047 2203 1048 2207
rect 1052 2206 1053 2207
rect 1091 2207 1097 2208
rect 1091 2206 1092 2207
rect 1052 2204 1092 2206
rect 1052 2203 1053 2204
rect 1047 2202 1053 2203
rect 1091 2203 1092 2204
rect 1096 2203 1097 2207
rect 1091 2202 1097 2203
rect 1138 2207 1144 2208
rect 1138 2203 1139 2207
rect 1143 2206 1144 2207
rect 1211 2207 1217 2208
rect 1211 2206 1212 2207
rect 1143 2204 1212 2206
rect 1143 2203 1144 2204
rect 1138 2202 1144 2203
rect 1211 2203 1212 2204
rect 1216 2203 1217 2207
rect 1211 2202 1217 2203
rect 2371 2207 2380 2208
rect 2371 2203 2372 2207
rect 2379 2203 2380 2207
rect 2371 2202 2380 2203
rect 2439 2207 2445 2208
rect 2439 2203 2440 2207
rect 2444 2206 2445 2207
rect 2483 2207 2489 2208
rect 2483 2206 2484 2207
rect 2444 2204 2484 2206
rect 2444 2203 2445 2204
rect 2439 2202 2445 2203
rect 2483 2203 2484 2204
rect 2488 2203 2489 2207
rect 2483 2202 2489 2203
rect 2566 2207 2572 2208
rect 2566 2203 2567 2207
rect 2571 2206 2572 2207
rect 2619 2207 2625 2208
rect 2619 2206 2620 2207
rect 2571 2204 2620 2206
rect 2571 2203 2572 2204
rect 2566 2202 2572 2203
rect 2619 2203 2620 2204
rect 2624 2203 2625 2207
rect 2771 2205 2772 2209
rect 2776 2208 2942 2209
rect 2776 2205 2777 2208
rect 2771 2204 2777 2205
rect 2946 2207 2953 2208
rect 2619 2202 2625 2203
rect 2946 2203 2947 2207
rect 2952 2203 2953 2207
rect 2946 2202 2953 2203
rect 3014 2207 3020 2208
rect 3014 2203 3015 2207
rect 3019 2206 3020 2207
rect 3139 2207 3145 2208
rect 3139 2206 3140 2207
rect 3019 2204 3140 2206
rect 3019 2203 3020 2204
rect 3014 2202 3020 2203
rect 3139 2203 3140 2204
rect 3144 2203 3145 2207
rect 3139 2202 3145 2203
rect 3339 2207 3348 2208
rect 3339 2203 3340 2207
rect 3347 2203 3348 2207
rect 3339 2202 3348 2203
rect 3515 2207 3524 2208
rect 3515 2203 3516 2207
rect 3523 2203 3524 2207
rect 3515 2202 3524 2203
rect 978 2199 984 2200
rect 978 2198 979 2199
rect 812 2196 979 2198
rect 812 2194 814 2196
rect 978 2195 979 2196
rect 983 2195 984 2199
rect 978 2194 984 2195
rect 2283 2195 2289 2196
rect 811 2193 817 2194
rect 127 2191 133 2192
rect 127 2187 128 2191
rect 132 2190 133 2191
rect 171 2191 177 2192
rect 171 2190 172 2191
rect 132 2188 172 2190
rect 132 2187 133 2188
rect 127 2186 133 2187
rect 171 2187 172 2188
rect 176 2187 177 2191
rect 171 2186 177 2187
rect 207 2191 213 2192
rect 207 2187 208 2191
rect 212 2190 213 2191
rect 275 2191 281 2192
rect 275 2190 276 2191
rect 212 2188 276 2190
rect 212 2187 213 2188
rect 207 2186 213 2187
rect 275 2187 276 2188
rect 280 2187 281 2191
rect 275 2186 281 2187
rect 411 2191 417 2192
rect 411 2187 412 2191
rect 416 2190 417 2191
rect 426 2191 432 2192
rect 426 2190 427 2191
rect 416 2188 427 2190
rect 416 2187 417 2188
rect 411 2186 417 2187
rect 426 2187 427 2188
rect 431 2187 432 2191
rect 426 2186 432 2187
rect 471 2191 477 2192
rect 471 2187 472 2191
rect 476 2190 477 2191
rect 547 2191 553 2192
rect 547 2190 548 2191
rect 476 2188 548 2190
rect 476 2187 477 2188
rect 471 2186 477 2187
rect 547 2187 548 2188
rect 552 2187 553 2191
rect 547 2186 553 2187
rect 607 2191 613 2192
rect 607 2187 608 2191
rect 612 2190 613 2191
rect 683 2191 689 2192
rect 683 2190 684 2191
rect 612 2188 684 2190
rect 612 2187 613 2188
rect 607 2186 613 2187
rect 683 2187 684 2188
rect 688 2187 689 2191
rect 811 2189 812 2193
rect 816 2189 817 2193
rect 811 2188 817 2189
rect 863 2191 869 2192
rect 683 2186 689 2187
rect 863 2187 864 2191
rect 868 2190 869 2191
rect 939 2191 945 2192
rect 939 2190 940 2191
rect 868 2188 940 2190
rect 868 2187 869 2188
rect 863 2186 869 2187
rect 939 2187 940 2188
rect 944 2187 945 2191
rect 939 2186 945 2187
rect 1059 2191 1065 2192
rect 1059 2187 1060 2191
rect 1064 2190 1065 2191
rect 1119 2191 1125 2192
rect 1119 2190 1120 2191
rect 1064 2188 1120 2190
rect 1064 2187 1065 2188
rect 1059 2186 1065 2187
rect 1119 2187 1120 2188
rect 1124 2187 1125 2191
rect 1119 2186 1125 2187
rect 1187 2191 1193 2192
rect 1187 2187 1188 2191
rect 1192 2190 1193 2191
rect 1230 2191 1236 2192
rect 1230 2190 1231 2191
rect 1192 2188 1231 2190
rect 1192 2187 1193 2188
rect 1187 2186 1193 2187
rect 1230 2187 1231 2188
rect 1235 2187 1236 2191
rect 1230 2186 1236 2187
rect 1255 2191 1261 2192
rect 1255 2187 1256 2191
rect 1260 2190 1261 2191
rect 1315 2191 1321 2192
rect 1315 2190 1316 2191
rect 1260 2188 1316 2190
rect 1260 2187 1261 2188
rect 1255 2186 1261 2187
rect 1315 2187 1316 2188
rect 1320 2187 1321 2191
rect 2283 2191 2284 2195
rect 2288 2194 2289 2195
rect 2322 2195 2328 2196
rect 2322 2194 2323 2195
rect 2288 2192 2323 2194
rect 2288 2191 2289 2192
rect 2283 2190 2289 2191
rect 2322 2191 2323 2192
rect 2327 2191 2328 2195
rect 2322 2190 2328 2191
rect 2371 2195 2377 2196
rect 2371 2191 2372 2195
rect 2376 2194 2377 2195
rect 2410 2195 2416 2196
rect 2410 2194 2411 2195
rect 2376 2192 2411 2194
rect 2376 2191 2377 2192
rect 2371 2190 2377 2191
rect 2410 2191 2411 2192
rect 2415 2191 2416 2195
rect 2410 2190 2416 2191
rect 2467 2195 2473 2196
rect 2467 2191 2468 2195
rect 2472 2194 2473 2195
rect 2514 2195 2520 2196
rect 2514 2194 2515 2195
rect 2472 2192 2515 2194
rect 2472 2191 2473 2192
rect 2467 2190 2473 2191
rect 2514 2191 2515 2192
rect 2519 2191 2520 2195
rect 2514 2190 2520 2191
rect 2574 2195 2585 2196
rect 2574 2191 2575 2195
rect 2579 2191 2580 2195
rect 2584 2191 2585 2195
rect 2574 2190 2585 2191
rect 2723 2195 2732 2196
rect 2723 2191 2724 2195
rect 2731 2191 2732 2195
rect 2723 2190 2732 2191
rect 2822 2195 2828 2196
rect 2822 2191 2823 2195
rect 2827 2194 2828 2195
rect 2899 2195 2905 2196
rect 2899 2194 2900 2195
rect 2827 2192 2900 2194
rect 2827 2191 2828 2192
rect 2822 2190 2828 2191
rect 2899 2191 2900 2192
rect 2904 2191 2905 2195
rect 2899 2190 2905 2191
rect 2943 2195 2949 2196
rect 2943 2191 2944 2195
rect 2948 2194 2949 2195
rect 3099 2195 3105 2196
rect 3099 2194 3100 2195
rect 2948 2192 3100 2194
rect 2948 2191 2949 2192
rect 2943 2190 2949 2191
rect 3099 2191 3100 2192
rect 3104 2191 3105 2195
rect 3099 2190 3105 2191
rect 3199 2195 3205 2196
rect 3199 2191 3200 2195
rect 3204 2194 3205 2195
rect 3315 2195 3321 2196
rect 3315 2194 3316 2195
rect 3204 2192 3316 2194
rect 3204 2191 3205 2192
rect 3199 2190 3205 2191
rect 3315 2191 3316 2192
rect 3320 2191 3321 2195
rect 3315 2190 3321 2191
rect 3515 2195 3521 2196
rect 3515 2191 3516 2195
rect 3520 2194 3521 2195
rect 3546 2195 3552 2196
rect 3546 2194 3547 2195
rect 3520 2192 3547 2194
rect 3520 2191 3521 2192
rect 3515 2190 3521 2191
rect 3546 2191 3547 2192
rect 3551 2191 3552 2195
rect 3546 2190 3552 2191
rect 1315 2186 1321 2187
rect 2254 2185 2260 2186
rect 142 2181 148 2182
rect 142 2177 143 2181
rect 147 2177 148 2181
rect 142 2176 148 2177
rect 246 2181 252 2182
rect 246 2177 247 2181
rect 251 2177 252 2181
rect 246 2176 252 2177
rect 382 2181 388 2182
rect 382 2177 383 2181
rect 387 2177 388 2181
rect 382 2176 388 2177
rect 518 2181 524 2182
rect 518 2177 519 2181
rect 523 2177 524 2181
rect 518 2176 524 2177
rect 654 2181 660 2182
rect 654 2177 655 2181
rect 659 2177 660 2181
rect 654 2176 660 2177
rect 782 2181 788 2182
rect 782 2177 783 2181
rect 787 2177 788 2181
rect 782 2176 788 2177
rect 910 2181 916 2182
rect 910 2177 911 2181
rect 915 2177 916 2181
rect 910 2176 916 2177
rect 1030 2181 1036 2182
rect 1030 2177 1031 2181
rect 1035 2177 1036 2181
rect 1030 2176 1036 2177
rect 1158 2181 1164 2182
rect 1158 2177 1159 2181
rect 1163 2177 1164 2181
rect 1158 2176 1164 2177
rect 1286 2181 1292 2182
rect 1286 2177 1287 2181
rect 1291 2177 1292 2181
rect 2254 2181 2255 2185
rect 2259 2181 2260 2185
rect 2254 2180 2260 2181
rect 2342 2185 2348 2186
rect 2342 2181 2343 2185
rect 2347 2181 2348 2185
rect 2342 2180 2348 2181
rect 2438 2185 2444 2186
rect 2438 2181 2439 2185
rect 2443 2181 2444 2185
rect 2438 2180 2444 2181
rect 2550 2185 2556 2186
rect 2550 2181 2551 2185
rect 2555 2181 2556 2185
rect 2550 2180 2556 2181
rect 2694 2185 2700 2186
rect 2694 2181 2695 2185
rect 2699 2181 2700 2185
rect 2694 2180 2700 2181
rect 2870 2185 2876 2186
rect 2870 2181 2871 2185
rect 2875 2181 2876 2185
rect 2870 2180 2876 2181
rect 3070 2185 3076 2186
rect 3070 2181 3071 2185
rect 3075 2181 3076 2185
rect 3070 2180 3076 2181
rect 3286 2185 3292 2186
rect 3286 2181 3287 2185
rect 3291 2181 3292 2185
rect 3286 2180 3292 2181
rect 3486 2185 3492 2186
rect 3486 2181 3487 2185
rect 3491 2181 3492 2185
rect 3486 2180 3492 2181
rect 1286 2176 1292 2177
rect 1862 2172 1868 2173
rect 3574 2172 3580 2173
rect 110 2168 116 2169
rect 1822 2168 1828 2169
rect 110 2164 111 2168
rect 115 2164 116 2168
rect 207 2167 213 2168
rect 207 2166 208 2167
rect 197 2164 208 2166
rect 110 2163 116 2164
rect 207 2163 208 2164
rect 212 2163 213 2167
rect 471 2167 477 2168
rect 471 2166 472 2167
rect 437 2164 472 2166
rect 207 2162 213 2163
rect 471 2163 472 2164
rect 476 2163 477 2167
rect 607 2167 613 2168
rect 607 2166 608 2167
rect 573 2164 608 2166
rect 471 2162 477 2163
rect 607 2163 608 2164
rect 612 2163 613 2167
rect 863 2167 869 2168
rect 863 2166 864 2167
rect 837 2164 864 2166
rect 607 2162 613 2163
rect 630 2163 636 2164
rect 630 2159 631 2163
rect 635 2162 636 2163
rect 863 2163 864 2164
rect 868 2163 869 2167
rect 970 2167 976 2168
rect 970 2166 971 2167
rect 965 2164 971 2166
rect 863 2162 869 2163
rect 970 2163 971 2164
rect 975 2163 976 2167
rect 1822 2164 1823 2168
rect 1827 2164 1828 2168
rect 1862 2168 1863 2172
rect 1867 2168 1868 2172
rect 2822 2171 2828 2172
rect 2822 2170 2823 2171
rect 2749 2168 2823 2170
rect 1862 2167 1868 2168
rect 2322 2167 2328 2168
rect 970 2162 976 2163
rect 978 2163 984 2164
rect 635 2160 673 2162
rect 635 2159 636 2160
rect 630 2158 636 2159
rect 978 2159 979 2163
rect 983 2162 984 2163
rect 1119 2163 1125 2164
rect 983 2160 1049 2162
rect 983 2159 984 2160
rect 978 2158 984 2159
rect 1119 2159 1120 2163
rect 1124 2162 1125 2163
rect 1230 2163 1236 2164
rect 1822 2163 1828 2164
rect 2322 2163 2323 2167
rect 2327 2166 2328 2167
rect 2410 2167 2416 2168
rect 2327 2164 2361 2166
rect 2327 2163 2328 2164
rect 1124 2160 1177 2162
rect 1124 2159 1125 2160
rect 1119 2158 1125 2159
rect 1230 2159 1231 2163
rect 1235 2162 1236 2163
rect 2322 2162 2328 2163
rect 2410 2163 2411 2167
rect 2415 2166 2416 2167
rect 2514 2167 2520 2168
rect 2415 2164 2457 2166
rect 2415 2163 2416 2164
rect 2410 2162 2416 2163
rect 2514 2163 2515 2167
rect 2519 2166 2520 2167
rect 2822 2167 2823 2168
rect 2827 2167 2828 2171
rect 2943 2171 2949 2172
rect 2943 2170 2944 2171
rect 2925 2168 2944 2170
rect 2822 2166 2828 2167
rect 2943 2167 2944 2168
rect 2948 2167 2949 2171
rect 3199 2171 3205 2172
rect 3199 2170 3200 2171
rect 3125 2168 3200 2170
rect 2943 2166 2949 2167
rect 3199 2167 3200 2168
rect 3204 2167 3205 2171
rect 3574 2168 3575 2172
rect 3579 2168 3580 2172
rect 3574 2167 3580 2168
rect 3199 2166 3205 2167
rect 2519 2164 2569 2166
rect 2519 2163 2520 2164
rect 2514 2162 2520 2163
rect 1235 2160 1305 2162
rect 1235 2159 1236 2160
rect 1230 2158 1236 2159
rect 1862 2155 1868 2156
rect 110 2151 116 2152
rect 110 2147 111 2151
rect 115 2147 116 2151
rect 110 2146 116 2147
rect 1822 2151 1828 2152
rect 1822 2147 1823 2151
rect 1827 2147 1828 2151
rect 1862 2151 1863 2155
rect 1867 2151 1868 2155
rect 2342 2155 2348 2156
rect 2342 2154 2343 2155
rect 2305 2152 2343 2154
rect 1862 2150 1868 2151
rect 2342 2151 2343 2152
rect 2347 2151 2348 2155
rect 2342 2150 2348 2151
rect 3198 2155 3204 2156
rect 3198 2151 3199 2155
rect 3203 2154 3204 2155
rect 3574 2155 3580 2156
rect 3203 2152 3297 2154
rect 3203 2151 3204 2152
rect 3198 2150 3204 2151
rect 3574 2151 3575 2155
rect 3579 2151 3580 2155
rect 3574 2150 3580 2151
rect 1822 2146 1828 2147
rect 2246 2145 2252 2146
rect 134 2141 140 2142
rect 134 2137 135 2141
rect 139 2137 140 2141
rect 134 2136 140 2137
rect 238 2141 244 2142
rect 238 2137 239 2141
rect 243 2137 244 2141
rect 238 2136 244 2137
rect 374 2141 380 2142
rect 374 2137 375 2141
rect 379 2137 380 2141
rect 374 2136 380 2137
rect 510 2141 516 2142
rect 510 2137 511 2141
rect 515 2137 516 2141
rect 510 2136 516 2137
rect 646 2141 652 2142
rect 646 2137 647 2141
rect 651 2137 652 2141
rect 646 2136 652 2137
rect 774 2141 780 2142
rect 774 2137 775 2141
rect 779 2137 780 2141
rect 774 2136 780 2137
rect 902 2141 908 2142
rect 902 2137 903 2141
rect 907 2137 908 2141
rect 902 2136 908 2137
rect 1022 2141 1028 2142
rect 1022 2137 1023 2141
rect 1027 2137 1028 2141
rect 1022 2136 1028 2137
rect 1150 2141 1156 2142
rect 1150 2137 1151 2141
rect 1155 2137 1156 2141
rect 1150 2136 1156 2137
rect 1278 2141 1284 2142
rect 1278 2137 1279 2141
rect 1283 2137 1284 2141
rect 2246 2141 2247 2145
rect 2251 2141 2252 2145
rect 2246 2140 2252 2141
rect 2334 2145 2340 2146
rect 2334 2141 2335 2145
rect 2339 2141 2340 2145
rect 2334 2140 2340 2141
rect 2430 2145 2436 2146
rect 2430 2141 2431 2145
rect 2435 2141 2436 2145
rect 2430 2140 2436 2141
rect 2542 2145 2548 2146
rect 2542 2141 2543 2145
rect 2547 2141 2548 2145
rect 2542 2140 2548 2141
rect 2686 2145 2692 2146
rect 2686 2141 2687 2145
rect 2691 2141 2692 2145
rect 2686 2140 2692 2141
rect 2862 2145 2868 2146
rect 2862 2141 2863 2145
rect 2867 2141 2868 2145
rect 2862 2140 2868 2141
rect 3062 2145 3068 2146
rect 3062 2141 3063 2145
rect 3067 2141 3068 2145
rect 3062 2140 3068 2141
rect 3278 2145 3284 2146
rect 3278 2141 3279 2145
rect 3283 2141 3284 2145
rect 3278 2140 3284 2141
rect 3478 2145 3484 2146
rect 3478 2141 3479 2145
rect 3483 2141 3484 2145
rect 3478 2140 3484 2141
rect 1278 2136 1284 2137
rect 3518 2139 3524 2140
rect 270 2135 276 2136
rect 270 2131 271 2135
rect 275 2134 276 2135
rect 287 2135 293 2136
rect 287 2134 288 2135
rect 275 2132 288 2134
rect 275 2131 276 2132
rect 270 2130 276 2131
rect 287 2131 288 2132
rect 292 2131 293 2135
rect 3518 2135 3519 2139
rect 3523 2138 3524 2139
rect 3527 2139 3533 2140
rect 3527 2138 3528 2139
rect 3523 2136 3528 2138
rect 3523 2135 3524 2136
rect 3518 2134 3524 2135
rect 3527 2135 3528 2136
rect 3532 2135 3533 2139
rect 3527 2134 3533 2135
rect 287 2130 293 2131
rect 2150 2115 2156 2116
rect 134 2111 140 2112
rect 134 2107 135 2111
rect 139 2107 140 2111
rect 134 2106 140 2107
rect 230 2111 236 2112
rect 230 2107 231 2111
rect 235 2107 236 2111
rect 230 2106 236 2107
rect 358 2111 364 2112
rect 358 2107 359 2111
rect 363 2107 364 2111
rect 358 2106 364 2107
rect 478 2111 484 2112
rect 478 2107 479 2111
rect 483 2107 484 2111
rect 478 2106 484 2107
rect 598 2111 604 2112
rect 598 2107 599 2111
rect 603 2107 604 2111
rect 598 2106 604 2107
rect 718 2111 724 2112
rect 718 2107 719 2111
rect 723 2107 724 2111
rect 718 2106 724 2107
rect 830 2111 836 2112
rect 830 2107 831 2111
rect 835 2107 836 2111
rect 830 2106 836 2107
rect 942 2111 948 2112
rect 942 2107 943 2111
rect 947 2107 948 2111
rect 942 2106 948 2107
rect 1054 2111 1060 2112
rect 1054 2107 1055 2111
rect 1059 2107 1060 2111
rect 1054 2106 1060 2107
rect 1174 2111 1180 2112
rect 1174 2107 1175 2111
rect 1179 2107 1180 2111
rect 2150 2111 2151 2115
rect 2155 2111 2156 2115
rect 2150 2110 2156 2111
rect 2238 2115 2244 2116
rect 2238 2111 2239 2115
rect 2243 2111 2244 2115
rect 2238 2110 2244 2111
rect 2326 2115 2332 2116
rect 2326 2111 2327 2115
rect 2331 2111 2332 2115
rect 2326 2110 2332 2111
rect 2414 2115 2420 2116
rect 2414 2111 2415 2115
rect 2419 2111 2420 2115
rect 2414 2110 2420 2111
rect 2502 2115 2508 2116
rect 2502 2111 2503 2115
rect 2507 2111 2508 2115
rect 2502 2110 2508 2111
rect 2614 2115 2620 2116
rect 2614 2111 2615 2115
rect 2619 2111 2620 2115
rect 2614 2110 2620 2111
rect 2750 2115 2756 2116
rect 2750 2111 2751 2115
rect 2755 2111 2756 2115
rect 2750 2110 2756 2111
rect 2918 2115 2924 2116
rect 2918 2111 2919 2115
rect 2923 2111 2924 2115
rect 2918 2110 2924 2111
rect 3102 2115 3108 2116
rect 3102 2111 3103 2115
rect 3107 2111 3108 2115
rect 3102 2110 3108 2111
rect 3302 2115 3308 2116
rect 3302 2111 3303 2115
rect 3307 2111 3308 2115
rect 3302 2110 3308 2111
rect 3478 2115 3484 2116
rect 3478 2111 3479 2115
rect 3483 2111 3484 2115
rect 3478 2110 3484 2111
rect 1174 2106 1180 2107
rect 2482 2107 2488 2108
rect 1862 2105 1868 2106
rect 426 2103 432 2104
rect 426 2102 427 2103
rect 110 2101 116 2102
rect 110 2097 111 2101
rect 115 2097 116 2101
rect 417 2100 427 2102
rect 426 2099 427 2100
rect 431 2099 432 2103
rect 1255 2103 1261 2104
rect 1255 2102 1256 2103
rect 1233 2100 1256 2102
rect 426 2098 432 2099
rect 1255 2099 1256 2100
rect 1260 2099 1261 2103
rect 1255 2098 1261 2099
rect 1822 2101 1828 2102
rect 110 2096 116 2097
rect 1822 2097 1823 2101
rect 1827 2097 1828 2101
rect 1862 2101 1863 2105
rect 1867 2101 1868 2105
rect 2482 2103 2483 2107
rect 2487 2106 2488 2107
rect 3199 2107 3205 2108
rect 2487 2104 2521 2106
rect 2487 2103 2488 2104
rect 2482 2102 2488 2103
rect 3199 2103 3200 2107
rect 3204 2106 3205 2107
rect 3204 2104 3321 2106
rect 3574 2105 3580 2106
rect 3204 2103 3205 2104
rect 3199 2102 3205 2103
rect 1862 2100 1868 2101
rect 3574 2101 3575 2105
rect 3579 2101 3580 2105
rect 3574 2100 3580 2101
rect 1822 2096 1828 2097
rect 2231 2091 2237 2092
rect 2231 2090 2232 2091
rect 1862 2088 1868 2089
rect 2213 2088 2232 2090
rect 202 2087 208 2088
rect 110 2084 116 2085
rect 110 2080 111 2084
rect 115 2080 116 2084
rect 110 2079 116 2080
rect 196 2078 198 2085
rect 202 2083 203 2087
rect 207 2086 208 2087
rect 426 2087 432 2088
rect 207 2084 257 2086
rect 207 2083 208 2084
rect 202 2082 208 2083
rect 426 2083 427 2087
rect 431 2086 432 2087
rect 546 2087 552 2088
rect 431 2084 505 2086
rect 431 2083 432 2084
rect 426 2082 432 2083
rect 546 2083 547 2087
rect 551 2086 552 2087
rect 823 2087 829 2088
rect 823 2086 824 2087
rect 551 2084 625 2086
rect 781 2084 824 2086
rect 551 2083 552 2084
rect 546 2082 552 2083
rect 823 2083 824 2084
rect 828 2083 829 2087
rect 935 2087 941 2088
rect 935 2086 936 2087
rect 893 2084 936 2086
rect 823 2082 829 2083
rect 935 2083 936 2084
rect 940 2083 941 2087
rect 1047 2087 1053 2088
rect 1047 2086 1048 2087
rect 1005 2084 1048 2086
rect 935 2082 941 2083
rect 1047 2083 1048 2084
rect 1052 2083 1053 2087
rect 1167 2087 1173 2088
rect 1167 2086 1168 2087
rect 1117 2084 1168 2086
rect 1047 2082 1053 2083
rect 1167 2083 1168 2084
rect 1172 2083 1173 2087
rect 1167 2082 1173 2083
rect 1822 2084 1828 2085
rect 1822 2080 1823 2084
rect 1827 2080 1828 2084
rect 1862 2084 1863 2088
rect 1867 2084 1868 2088
rect 2231 2087 2232 2088
rect 2236 2087 2237 2091
rect 2306 2091 2312 2092
rect 2306 2090 2307 2091
rect 2301 2088 2307 2090
rect 2231 2086 2237 2087
rect 2306 2087 2307 2088
rect 2311 2087 2312 2091
rect 2407 2091 2413 2092
rect 2407 2090 2408 2091
rect 2389 2088 2408 2090
rect 2306 2086 2312 2087
rect 2407 2087 2408 2088
rect 2412 2087 2413 2091
rect 2495 2091 2501 2092
rect 2495 2090 2496 2091
rect 2477 2088 2496 2090
rect 2407 2086 2413 2087
rect 2495 2087 2496 2088
rect 2500 2087 2501 2091
rect 2743 2091 2749 2092
rect 2743 2090 2744 2091
rect 2677 2088 2744 2090
rect 2495 2086 2501 2087
rect 2743 2087 2744 2088
rect 2748 2087 2749 2091
rect 2911 2091 2917 2092
rect 2911 2090 2912 2091
rect 2813 2088 2912 2090
rect 2743 2086 2749 2087
rect 2911 2087 2912 2088
rect 2916 2087 2917 2091
rect 3094 2091 3100 2092
rect 3094 2090 3095 2091
rect 2981 2088 3095 2090
rect 2911 2086 2917 2087
rect 3094 2087 3095 2088
rect 3099 2087 3100 2091
rect 3295 2091 3301 2092
rect 3295 2090 3296 2091
rect 3165 2088 3296 2090
rect 3094 2086 3100 2087
rect 3295 2087 3296 2088
rect 3300 2087 3301 2091
rect 3554 2091 3560 2092
rect 3554 2090 3555 2091
rect 3541 2088 3555 2090
rect 3295 2086 3301 2087
rect 3554 2087 3555 2088
rect 3559 2087 3560 2091
rect 3554 2086 3560 2087
rect 3574 2088 3580 2089
rect 1862 2083 1868 2084
rect 3574 2084 3575 2088
rect 3579 2084 3580 2088
rect 3574 2083 3580 2084
rect 207 2079 213 2080
rect 1822 2079 1828 2080
rect 207 2078 208 2079
rect 196 2076 208 2078
rect 207 2075 208 2076
rect 212 2075 213 2079
rect 207 2074 213 2075
rect 2158 2075 2164 2076
rect 142 2071 148 2072
rect 142 2067 143 2071
rect 147 2067 148 2071
rect 142 2066 148 2067
rect 238 2071 244 2072
rect 238 2067 239 2071
rect 243 2067 244 2071
rect 238 2066 244 2067
rect 366 2071 372 2072
rect 366 2067 367 2071
rect 371 2067 372 2071
rect 366 2066 372 2067
rect 486 2071 492 2072
rect 486 2067 487 2071
rect 491 2067 492 2071
rect 486 2066 492 2067
rect 606 2071 612 2072
rect 606 2067 607 2071
rect 611 2067 612 2071
rect 606 2066 612 2067
rect 726 2071 732 2072
rect 726 2067 727 2071
rect 731 2067 732 2071
rect 726 2066 732 2067
rect 838 2071 844 2072
rect 838 2067 839 2071
rect 843 2067 844 2071
rect 838 2066 844 2067
rect 950 2071 956 2072
rect 950 2067 951 2071
rect 955 2067 956 2071
rect 950 2066 956 2067
rect 1062 2071 1068 2072
rect 1062 2067 1063 2071
rect 1067 2067 1068 2071
rect 1062 2066 1068 2067
rect 1182 2071 1188 2072
rect 1182 2067 1183 2071
rect 1187 2067 1188 2071
rect 2158 2071 2159 2075
rect 2163 2071 2164 2075
rect 2158 2070 2164 2071
rect 2246 2075 2252 2076
rect 2246 2071 2247 2075
rect 2251 2071 2252 2075
rect 2246 2070 2252 2071
rect 2334 2075 2340 2076
rect 2334 2071 2335 2075
rect 2339 2071 2340 2075
rect 2334 2070 2340 2071
rect 2422 2075 2428 2076
rect 2422 2071 2423 2075
rect 2427 2071 2428 2075
rect 2422 2070 2428 2071
rect 2510 2075 2516 2076
rect 2510 2071 2511 2075
rect 2515 2071 2516 2075
rect 2510 2070 2516 2071
rect 2622 2075 2628 2076
rect 2622 2071 2623 2075
rect 2627 2071 2628 2075
rect 2622 2070 2628 2071
rect 2758 2075 2764 2076
rect 2758 2071 2759 2075
rect 2763 2071 2764 2075
rect 2758 2070 2764 2071
rect 2926 2075 2932 2076
rect 2926 2071 2927 2075
rect 2931 2071 2932 2075
rect 2926 2070 2932 2071
rect 3110 2075 3116 2076
rect 3110 2071 3111 2075
rect 3115 2071 3116 2075
rect 3110 2070 3116 2071
rect 3310 2075 3316 2076
rect 3310 2071 3311 2075
rect 3315 2071 3316 2075
rect 3310 2070 3316 2071
rect 3486 2075 3492 2076
rect 3486 2071 3487 2075
rect 3491 2071 3492 2075
rect 3486 2070 3492 2071
rect 1182 2066 1188 2067
rect 2187 2063 2196 2064
rect 171 2059 177 2060
rect 171 2055 172 2059
rect 176 2058 177 2059
rect 202 2059 208 2060
rect 202 2058 203 2059
rect 176 2056 203 2058
rect 176 2055 177 2056
rect 171 2054 177 2055
rect 202 2055 203 2056
rect 207 2055 208 2059
rect 202 2054 208 2055
rect 267 2059 276 2060
rect 267 2055 268 2059
rect 275 2055 276 2059
rect 267 2054 276 2055
rect 395 2059 401 2060
rect 395 2055 396 2059
rect 400 2058 401 2059
rect 426 2059 432 2060
rect 426 2058 427 2059
rect 400 2056 427 2058
rect 400 2055 401 2056
rect 395 2054 401 2055
rect 426 2055 427 2056
rect 431 2055 432 2059
rect 426 2054 432 2055
rect 515 2059 521 2060
rect 515 2055 516 2059
rect 520 2058 521 2059
rect 546 2059 552 2060
rect 546 2058 547 2059
rect 520 2056 547 2058
rect 520 2055 521 2056
rect 515 2054 521 2055
rect 546 2055 547 2056
rect 551 2055 552 2059
rect 546 2054 552 2055
rect 634 2059 641 2060
rect 634 2055 635 2059
rect 640 2055 641 2059
rect 634 2054 641 2055
rect 755 2059 764 2060
rect 755 2055 756 2059
rect 763 2055 764 2059
rect 755 2054 764 2055
rect 823 2059 829 2060
rect 823 2055 824 2059
rect 828 2058 829 2059
rect 867 2059 873 2060
rect 867 2058 868 2059
rect 828 2056 868 2058
rect 828 2055 829 2056
rect 823 2054 829 2055
rect 867 2055 868 2056
rect 872 2055 873 2059
rect 867 2054 873 2055
rect 935 2059 941 2060
rect 935 2055 936 2059
rect 940 2058 941 2059
rect 979 2059 985 2060
rect 979 2058 980 2059
rect 940 2056 980 2058
rect 940 2055 941 2056
rect 935 2054 941 2055
rect 979 2055 980 2056
rect 984 2055 985 2059
rect 979 2054 985 2055
rect 1047 2059 1053 2060
rect 1047 2055 1048 2059
rect 1052 2058 1053 2059
rect 1091 2059 1097 2060
rect 1091 2058 1092 2059
rect 1052 2056 1092 2058
rect 1052 2055 1053 2056
rect 1047 2054 1053 2055
rect 1091 2055 1092 2056
rect 1096 2055 1097 2059
rect 1091 2054 1097 2055
rect 1167 2059 1173 2060
rect 1167 2055 1168 2059
rect 1172 2058 1173 2059
rect 1211 2059 1217 2060
rect 1211 2058 1212 2059
rect 1172 2056 1212 2058
rect 1172 2055 1173 2056
rect 1167 2054 1173 2055
rect 1211 2055 1212 2056
rect 1216 2055 1217 2059
rect 2187 2059 2188 2063
rect 2195 2059 2196 2063
rect 2187 2058 2196 2059
rect 2231 2063 2237 2064
rect 2231 2059 2232 2063
rect 2236 2062 2237 2063
rect 2275 2063 2281 2064
rect 2275 2062 2276 2063
rect 2236 2060 2276 2062
rect 2236 2059 2237 2060
rect 2231 2058 2237 2059
rect 2275 2059 2276 2060
rect 2280 2059 2281 2063
rect 2275 2058 2281 2059
rect 2342 2063 2348 2064
rect 2342 2059 2343 2063
rect 2347 2062 2348 2063
rect 2363 2063 2369 2064
rect 2363 2062 2364 2063
rect 2347 2060 2364 2062
rect 2347 2059 2348 2060
rect 2342 2058 2348 2059
rect 2363 2059 2364 2060
rect 2368 2059 2369 2063
rect 2363 2058 2369 2059
rect 2407 2063 2413 2064
rect 2407 2059 2408 2063
rect 2412 2062 2413 2063
rect 2451 2063 2457 2064
rect 2451 2062 2452 2063
rect 2412 2060 2452 2062
rect 2412 2059 2413 2060
rect 2407 2058 2413 2059
rect 2451 2059 2452 2060
rect 2456 2059 2457 2063
rect 2451 2058 2457 2059
rect 2495 2063 2501 2064
rect 2495 2059 2496 2063
rect 2500 2062 2501 2063
rect 2539 2063 2545 2064
rect 2539 2062 2540 2063
rect 2500 2060 2540 2062
rect 2500 2059 2501 2060
rect 2495 2058 2501 2059
rect 2539 2059 2540 2060
rect 2544 2059 2545 2063
rect 2539 2058 2545 2059
rect 2651 2063 2657 2064
rect 2651 2059 2652 2063
rect 2656 2062 2657 2063
rect 2662 2063 2668 2064
rect 2662 2062 2663 2063
rect 2656 2060 2663 2062
rect 2656 2059 2657 2060
rect 2651 2058 2657 2059
rect 2662 2059 2663 2060
rect 2667 2059 2668 2063
rect 2662 2058 2668 2059
rect 2743 2063 2749 2064
rect 2743 2059 2744 2063
rect 2748 2062 2749 2063
rect 2787 2063 2793 2064
rect 2787 2062 2788 2063
rect 2748 2060 2788 2062
rect 2748 2059 2749 2060
rect 2743 2058 2749 2059
rect 2787 2059 2788 2060
rect 2792 2059 2793 2063
rect 2787 2058 2793 2059
rect 2911 2063 2917 2064
rect 2911 2059 2912 2063
rect 2916 2062 2917 2063
rect 2955 2063 2961 2064
rect 2955 2062 2956 2063
rect 2916 2060 2956 2062
rect 2916 2059 2917 2060
rect 2911 2058 2917 2059
rect 2955 2059 2956 2060
rect 2960 2059 2961 2063
rect 2955 2058 2961 2059
rect 3094 2063 3100 2064
rect 3094 2059 3095 2063
rect 3099 2062 3100 2063
rect 3139 2063 3145 2064
rect 3139 2062 3140 2063
rect 3099 2060 3140 2062
rect 3099 2059 3100 2060
rect 3094 2058 3100 2059
rect 3139 2059 3140 2060
rect 3144 2059 3145 2063
rect 3139 2058 3145 2059
rect 3295 2063 3301 2064
rect 3295 2059 3296 2063
rect 3300 2062 3301 2063
rect 3339 2063 3345 2064
rect 3339 2062 3340 2063
rect 3300 2060 3340 2062
rect 3300 2059 3301 2060
rect 3295 2058 3301 2059
rect 3339 2059 3340 2060
rect 3344 2059 3345 2063
rect 3339 2058 3345 2059
rect 3515 2063 3524 2064
rect 3515 2059 3516 2063
rect 3523 2059 3524 2063
rect 3515 2058 3524 2059
rect 1211 2054 1217 2055
rect 3199 2055 3205 2056
rect 3199 2054 3200 2055
rect 2740 2052 3200 2054
rect 2740 2050 2742 2052
rect 3199 2051 3200 2052
rect 3204 2051 3205 2055
rect 3199 2050 3205 2051
rect 2739 2049 2745 2050
rect 2027 2047 2033 2048
rect 2027 2043 2028 2047
rect 2032 2046 2033 2047
rect 2070 2047 2076 2048
rect 2070 2046 2071 2047
rect 2032 2044 2071 2046
rect 2032 2043 2033 2044
rect 2027 2042 2033 2043
rect 2070 2043 2071 2044
rect 2075 2043 2076 2047
rect 2070 2042 2076 2043
rect 2079 2047 2085 2048
rect 2079 2043 2080 2047
rect 2084 2046 2085 2047
rect 2155 2047 2161 2048
rect 2155 2046 2156 2047
rect 2084 2044 2156 2046
rect 2084 2043 2085 2044
rect 2079 2042 2085 2043
rect 2155 2043 2156 2044
rect 2160 2043 2161 2047
rect 2155 2042 2161 2043
rect 2283 2047 2289 2048
rect 2283 2043 2284 2047
rect 2288 2046 2289 2047
rect 2306 2047 2312 2048
rect 2306 2046 2307 2047
rect 2288 2044 2307 2046
rect 2288 2043 2289 2044
rect 2283 2042 2289 2043
rect 2306 2043 2307 2044
rect 2311 2043 2312 2047
rect 2306 2042 2312 2043
rect 2366 2047 2372 2048
rect 2366 2043 2367 2047
rect 2371 2046 2372 2047
rect 2427 2047 2433 2048
rect 2427 2046 2428 2047
rect 2371 2044 2428 2046
rect 2371 2043 2372 2044
rect 2366 2042 2372 2043
rect 2427 2043 2428 2044
rect 2432 2043 2433 2047
rect 2427 2042 2433 2043
rect 2463 2047 2469 2048
rect 2463 2043 2464 2047
rect 2468 2046 2469 2047
rect 2579 2047 2585 2048
rect 2579 2046 2580 2047
rect 2468 2044 2580 2046
rect 2468 2043 2469 2044
rect 2463 2042 2469 2043
rect 2579 2043 2580 2044
rect 2584 2043 2585 2047
rect 2739 2045 2740 2049
rect 2744 2045 2745 2049
rect 2739 2044 2745 2045
rect 2830 2047 2836 2048
rect 2579 2042 2585 2043
rect 2830 2043 2831 2047
rect 2835 2046 2836 2047
rect 2907 2047 2913 2048
rect 2907 2046 2908 2047
rect 2835 2044 2908 2046
rect 2835 2043 2836 2044
rect 2830 2042 2836 2043
rect 2907 2043 2908 2044
rect 2912 2043 2913 2047
rect 2907 2042 2913 2043
rect 2990 2047 2996 2048
rect 2990 2043 2991 2047
rect 2995 2046 2996 2047
rect 3091 2047 3097 2048
rect 3091 2046 3092 2047
rect 2995 2044 3092 2046
rect 2995 2043 2996 2044
rect 2990 2042 2996 2043
rect 3091 2043 3092 2044
rect 3096 2043 3097 2047
rect 3091 2042 3097 2043
rect 3174 2047 3180 2048
rect 3174 2043 3175 2047
rect 3179 2046 3180 2047
rect 3275 2047 3281 2048
rect 3275 2046 3276 2047
rect 3179 2044 3276 2046
rect 3179 2043 3180 2044
rect 3174 2042 3180 2043
rect 3275 2043 3276 2044
rect 3280 2043 3281 2047
rect 3275 2042 3281 2043
rect 3418 2047 3424 2048
rect 3418 2043 3419 2047
rect 3423 2046 3424 2047
rect 3467 2047 3473 2048
rect 3467 2046 3468 2047
rect 3423 2044 3468 2046
rect 3423 2043 3424 2044
rect 3418 2042 3424 2043
rect 3467 2043 3468 2044
rect 3472 2043 3473 2047
rect 3467 2042 3473 2043
rect 1998 2037 2004 2038
rect 195 2035 201 2036
rect 195 2031 196 2035
rect 200 2034 201 2035
rect 207 2035 213 2036
rect 207 2034 208 2035
rect 200 2032 208 2034
rect 200 2031 201 2032
rect 195 2030 201 2031
rect 207 2031 208 2032
rect 212 2031 213 2035
rect 207 2030 213 2031
rect 339 2035 345 2036
rect 339 2031 340 2035
rect 344 2034 345 2035
rect 386 2035 392 2036
rect 386 2034 387 2035
rect 344 2032 387 2034
rect 344 2031 345 2032
rect 339 2030 345 2031
rect 386 2031 387 2032
rect 391 2031 392 2035
rect 386 2030 392 2031
rect 398 2035 404 2036
rect 398 2031 399 2035
rect 403 2034 404 2035
rect 475 2035 481 2036
rect 475 2034 476 2035
rect 403 2032 476 2034
rect 403 2031 404 2032
rect 398 2030 404 2031
rect 475 2031 476 2032
rect 480 2031 481 2035
rect 475 2030 481 2031
rect 527 2035 533 2036
rect 527 2031 528 2035
rect 532 2034 533 2035
rect 603 2035 609 2036
rect 603 2034 604 2035
rect 532 2032 604 2034
rect 532 2031 533 2032
rect 527 2030 533 2031
rect 603 2031 604 2032
rect 608 2031 609 2035
rect 603 2030 609 2031
rect 723 2035 729 2036
rect 723 2031 724 2035
rect 728 2034 729 2035
rect 754 2035 760 2036
rect 728 2032 730 2034
rect 728 2031 732 2032
rect 723 2030 727 2031
rect 726 2027 727 2030
rect 731 2027 732 2031
rect 754 2031 755 2035
rect 759 2034 760 2035
rect 835 2035 841 2036
rect 835 2034 836 2035
rect 759 2032 836 2034
rect 759 2031 760 2032
rect 754 2030 760 2031
rect 835 2031 836 2032
rect 840 2031 841 2035
rect 835 2030 841 2031
rect 939 2035 945 2036
rect 939 2031 940 2035
rect 944 2034 945 2035
rect 982 2035 988 2036
rect 982 2034 983 2035
rect 944 2032 983 2034
rect 944 2031 945 2032
rect 939 2030 945 2031
rect 982 2031 983 2032
rect 987 2031 988 2035
rect 982 2030 988 2031
rect 1043 2035 1049 2036
rect 1043 2031 1044 2035
rect 1048 2034 1049 2035
rect 1082 2035 1088 2036
rect 1082 2034 1083 2035
rect 1048 2032 1083 2034
rect 1048 2031 1049 2032
rect 1043 2030 1049 2031
rect 1082 2031 1083 2032
rect 1087 2031 1088 2035
rect 1082 2030 1088 2031
rect 1147 2035 1153 2036
rect 1147 2031 1148 2035
rect 1152 2034 1153 2035
rect 1190 2035 1196 2036
rect 1190 2034 1191 2035
rect 1152 2032 1191 2034
rect 1152 2031 1153 2032
rect 1147 2030 1153 2031
rect 1190 2031 1191 2032
rect 1195 2031 1196 2035
rect 1190 2030 1196 2031
rect 1251 2035 1257 2036
rect 1251 2031 1252 2035
rect 1256 2034 1257 2035
rect 1295 2035 1301 2036
rect 1295 2034 1296 2035
rect 1256 2032 1296 2034
rect 1256 2031 1257 2032
rect 1251 2030 1257 2031
rect 1295 2031 1296 2032
rect 1300 2031 1301 2035
rect 1295 2030 1301 2031
rect 1310 2035 1316 2036
rect 1310 2031 1311 2035
rect 1315 2034 1316 2035
rect 1355 2035 1361 2036
rect 1355 2034 1356 2035
rect 1315 2032 1356 2034
rect 1315 2031 1316 2032
rect 1310 2030 1316 2031
rect 1355 2031 1356 2032
rect 1360 2031 1361 2035
rect 1998 2033 1999 2037
rect 2003 2033 2004 2037
rect 1998 2032 2004 2033
rect 2126 2037 2132 2038
rect 2126 2033 2127 2037
rect 2131 2033 2132 2037
rect 2126 2032 2132 2033
rect 2254 2037 2260 2038
rect 2254 2033 2255 2037
rect 2259 2033 2260 2037
rect 2254 2032 2260 2033
rect 2398 2037 2404 2038
rect 2398 2033 2399 2037
rect 2403 2033 2404 2037
rect 2398 2032 2404 2033
rect 2550 2037 2556 2038
rect 2550 2033 2551 2037
rect 2555 2033 2556 2037
rect 2550 2032 2556 2033
rect 2710 2037 2716 2038
rect 2710 2033 2711 2037
rect 2715 2033 2716 2037
rect 2710 2032 2716 2033
rect 2878 2037 2884 2038
rect 2878 2033 2879 2037
rect 2883 2033 2884 2037
rect 2878 2032 2884 2033
rect 3062 2037 3068 2038
rect 3062 2033 3063 2037
rect 3067 2033 3068 2037
rect 3062 2032 3068 2033
rect 3246 2037 3252 2038
rect 3246 2033 3247 2037
rect 3251 2033 3252 2037
rect 3246 2032 3252 2033
rect 3438 2037 3444 2038
rect 3438 2033 3439 2037
rect 3443 2033 3444 2037
rect 3438 2032 3444 2033
rect 1355 2030 1361 2031
rect 726 2026 732 2027
rect 166 2025 172 2026
rect 166 2021 167 2025
rect 171 2021 172 2025
rect 166 2020 172 2021
rect 310 2025 316 2026
rect 310 2021 311 2025
rect 315 2021 316 2025
rect 310 2020 316 2021
rect 446 2025 452 2026
rect 446 2021 447 2025
rect 451 2021 452 2025
rect 446 2020 452 2021
rect 574 2025 580 2026
rect 574 2021 575 2025
rect 579 2021 580 2025
rect 574 2020 580 2021
rect 694 2025 700 2026
rect 694 2021 695 2025
rect 699 2021 700 2025
rect 694 2020 700 2021
rect 806 2025 812 2026
rect 806 2021 807 2025
rect 811 2021 812 2025
rect 806 2020 812 2021
rect 910 2025 916 2026
rect 910 2021 911 2025
rect 915 2021 916 2025
rect 910 2020 916 2021
rect 1014 2025 1020 2026
rect 1014 2021 1015 2025
rect 1019 2021 1020 2025
rect 1014 2020 1020 2021
rect 1118 2025 1124 2026
rect 1118 2021 1119 2025
rect 1123 2021 1124 2025
rect 1118 2020 1124 2021
rect 1222 2025 1228 2026
rect 1222 2021 1223 2025
rect 1227 2021 1228 2025
rect 1222 2020 1228 2021
rect 1326 2025 1332 2026
rect 1326 2021 1327 2025
rect 1331 2021 1332 2025
rect 1326 2020 1332 2021
rect 1862 2024 1868 2025
rect 3574 2024 3580 2025
rect 1862 2020 1863 2024
rect 1867 2020 1868 2024
rect 2079 2023 2085 2024
rect 2079 2022 2080 2023
rect 2053 2020 2080 2022
rect 1862 2019 1868 2020
rect 2079 2019 2080 2020
rect 2084 2019 2085 2023
rect 2366 2023 2372 2024
rect 2366 2022 2367 2023
rect 2309 2020 2367 2022
rect 2079 2018 2085 2019
rect 2366 2019 2367 2020
rect 2371 2019 2372 2023
rect 2463 2023 2469 2024
rect 2463 2022 2464 2023
rect 2453 2020 2464 2022
rect 2366 2018 2372 2019
rect 2463 2019 2464 2020
rect 2468 2019 2469 2023
rect 2830 2023 2836 2024
rect 2830 2022 2831 2023
rect 2765 2020 2831 2022
rect 2463 2018 2469 2019
rect 2478 2019 2484 2020
rect 2478 2015 2479 2019
rect 2483 2018 2484 2019
rect 2830 2019 2831 2020
rect 2835 2019 2836 2023
rect 2990 2023 2996 2024
rect 2990 2022 2991 2023
rect 2933 2020 2991 2022
rect 2830 2018 2836 2019
rect 2990 2019 2991 2020
rect 2995 2019 2996 2023
rect 3174 2023 3180 2024
rect 3174 2022 3175 2023
rect 3117 2020 3175 2022
rect 2990 2018 2996 2019
rect 3174 2019 3175 2020
rect 3179 2019 3180 2023
rect 3574 2020 3575 2024
rect 3579 2020 3580 2024
rect 3174 2018 3180 2019
rect 3342 2019 3348 2020
rect 3574 2019 3580 2020
rect 2483 2016 2569 2018
rect 2483 2015 2484 2016
rect 2478 2014 2484 2015
rect 3342 2015 3343 2019
rect 3347 2018 3348 2019
rect 3347 2016 3457 2018
rect 3347 2015 3348 2016
rect 3342 2014 3348 2015
rect 110 2012 116 2013
rect 1822 2012 1828 2013
rect 110 2008 111 2012
rect 115 2008 116 2012
rect 398 2011 404 2012
rect 398 2010 399 2011
rect 365 2008 399 2010
rect 110 2007 116 2008
rect 398 2007 399 2008
rect 403 2007 404 2011
rect 527 2011 533 2012
rect 527 2010 528 2011
rect 501 2008 528 2010
rect 398 2006 404 2007
rect 527 2007 528 2008
rect 532 2007 533 2011
rect 634 2011 640 2012
rect 634 2010 635 2011
rect 629 2008 635 2010
rect 527 2006 533 2007
rect 634 2007 635 2008
rect 639 2007 640 2011
rect 754 2011 760 2012
rect 754 2010 755 2011
rect 749 2008 755 2010
rect 634 2006 640 2007
rect 754 2007 755 2008
rect 759 2007 760 2011
rect 1822 2008 1823 2012
rect 1827 2008 1828 2012
rect 754 2006 760 2007
rect 762 2007 768 2008
rect 762 2003 763 2007
rect 767 2006 768 2007
rect 982 2007 988 2008
rect 767 2004 825 2006
rect 767 2003 768 2004
rect 762 2002 768 2003
rect 982 2003 983 2007
rect 987 2006 988 2007
rect 1082 2007 1088 2008
rect 987 2004 1033 2006
rect 987 2003 988 2004
rect 982 2002 988 2003
rect 1082 2003 1083 2007
rect 1087 2006 1088 2007
rect 1190 2007 1196 2008
rect 1087 2004 1137 2006
rect 1087 2003 1088 2004
rect 1082 2002 1088 2003
rect 1190 2003 1191 2007
rect 1195 2006 1196 2007
rect 1295 2007 1301 2008
rect 1822 2007 1828 2008
rect 1862 2007 1868 2008
rect 1195 2004 1241 2006
rect 1195 2003 1196 2004
rect 1190 2002 1196 2003
rect 1295 2003 1296 2007
rect 1300 2006 1301 2007
rect 1300 2004 1345 2006
rect 1300 2003 1301 2004
rect 1295 2002 1301 2003
rect 1862 2003 1863 2007
rect 1867 2003 1868 2007
rect 2194 2007 2200 2008
rect 2194 2006 2195 2007
rect 2177 2004 2195 2006
rect 1862 2002 1868 2003
rect 2194 2003 2195 2004
rect 2199 2003 2200 2007
rect 2194 2002 2200 2003
rect 3150 2007 3156 2008
rect 3150 2003 3151 2007
rect 3155 2006 3156 2007
rect 3574 2007 3580 2008
rect 3155 2004 3257 2006
rect 3155 2003 3156 2004
rect 3150 2002 3156 2003
rect 3574 2003 3575 2007
rect 3579 2003 3580 2007
rect 3574 2002 3580 2003
rect 1990 1997 1996 1998
rect 110 1995 116 1996
rect 110 1991 111 1995
rect 115 1991 116 1995
rect 1014 1995 1020 1996
rect 1014 1994 1015 1995
rect 961 1992 1015 1994
rect 110 1990 116 1991
rect 1014 1991 1015 1992
rect 1019 1991 1020 1995
rect 1014 1990 1020 1991
rect 1822 1995 1828 1996
rect 1822 1991 1823 1995
rect 1827 1991 1828 1995
rect 1990 1993 1991 1997
rect 1995 1993 1996 1997
rect 1990 1992 1996 1993
rect 2118 1997 2124 1998
rect 2118 1993 2119 1997
rect 2123 1993 2124 1997
rect 2118 1992 2124 1993
rect 2246 1997 2252 1998
rect 2246 1993 2247 1997
rect 2251 1993 2252 1997
rect 2246 1992 2252 1993
rect 2390 1997 2396 1998
rect 2390 1993 2391 1997
rect 2395 1993 2396 1997
rect 2390 1992 2396 1993
rect 2542 1997 2548 1998
rect 2542 1993 2543 1997
rect 2547 1993 2548 1997
rect 2542 1992 2548 1993
rect 2702 1997 2708 1998
rect 2702 1993 2703 1997
rect 2707 1993 2708 1997
rect 2702 1992 2708 1993
rect 2870 1997 2876 1998
rect 2870 1993 2871 1997
rect 2875 1993 2876 1997
rect 2870 1992 2876 1993
rect 3054 1997 3060 1998
rect 3054 1993 3055 1997
rect 3059 1993 3060 1997
rect 3054 1992 3060 1993
rect 3238 1997 3244 1998
rect 3238 1993 3239 1997
rect 3243 1993 3244 1997
rect 3238 1992 3244 1993
rect 3430 1997 3436 1998
rect 3430 1993 3431 1997
rect 3435 1993 3436 1997
rect 3430 1992 3436 1993
rect 1822 1990 1828 1991
rect 158 1985 164 1986
rect 158 1981 159 1985
rect 163 1981 164 1985
rect 158 1980 164 1981
rect 302 1985 308 1986
rect 302 1981 303 1985
rect 307 1981 308 1985
rect 302 1980 308 1981
rect 438 1985 444 1986
rect 438 1981 439 1985
rect 443 1981 444 1985
rect 438 1980 444 1981
rect 566 1985 572 1986
rect 566 1981 567 1985
rect 571 1981 572 1985
rect 566 1980 572 1981
rect 686 1985 692 1986
rect 686 1981 687 1985
rect 691 1981 692 1985
rect 686 1980 692 1981
rect 798 1985 804 1986
rect 798 1981 799 1985
rect 803 1981 804 1985
rect 798 1980 804 1981
rect 902 1985 908 1986
rect 902 1981 903 1985
rect 907 1981 908 1985
rect 902 1980 908 1981
rect 1006 1985 1012 1986
rect 1006 1981 1007 1985
rect 1011 1981 1012 1985
rect 1006 1980 1012 1981
rect 1110 1985 1116 1986
rect 1110 1981 1111 1985
rect 1115 1981 1116 1985
rect 1110 1980 1116 1981
rect 1214 1985 1220 1986
rect 1214 1981 1215 1985
rect 1219 1981 1220 1985
rect 1214 1980 1220 1981
rect 1318 1985 1324 1986
rect 1318 1981 1319 1985
rect 1323 1981 1324 1985
rect 1318 1980 1324 1981
rect 206 1979 213 1980
rect 206 1975 207 1979
rect 212 1975 213 1979
rect 206 1974 213 1975
rect 1902 1967 1908 1968
rect 158 1963 164 1964
rect 158 1959 159 1963
rect 163 1959 164 1963
rect 158 1958 164 1959
rect 294 1963 300 1964
rect 294 1959 295 1963
rect 299 1959 300 1963
rect 294 1958 300 1959
rect 438 1963 444 1964
rect 438 1959 439 1963
rect 443 1959 444 1963
rect 438 1958 444 1959
rect 582 1963 588 1964
rect 582 1959 583 1963
rect 587 1959 588 1963
rect 582 1958 588 1959
rect 718 1963 724 1964
rect 718 1959 719 1963
rect 723 1959 724 1963
rect 718 1958 724 1959
rect 854 1963 860 1964
rect 854 1959 855 1963
rect 859 1959 860 1963
rect 854 1958 860 1959
rect 990 1963 996 1964
rect 990 1959 991 1963
rect 995 1959 996 1963
rect 990 1958 996 1959
rect 1118 1963 1124 1964
rect 1118 1959 1119 1963
rect 1123 1959 1124 1963
rect 1118 1958 1124 1959
rect 1238 1963 1244 1964
rect 1238 1959 1239 1963
rect 1243 1959 1244 1963
rect 1238 1958 1244 1959
rect 1358 1963 1364 1964
rect 1358 1959 1359 1963
rect 1363 1959 1364 1963
rect 1358 1958 1364 1959
rect 1478 1963 1484 1964
rect 1478 1959 1479 1963
rect 1483 1959 1484 1963
rect 1478 1958 1484 1959
rect 1598 1963 1604 1964
rect 1598 1959 1599 1963
rect 1603 1959 1604 1963
rect 1902 1963 1903 1967
rect 1907 1963 1908 1967
rect 1902 1962 1908 1963
rect 2158 1967 2164 1968
rect 2158 1963 2159 1967
rect 2163 1963 2164 1967
rect 2158 1962 2164 1963
rect 2398 1967 2404 1968
rect 2398 1963 2399 1967
rect 2403 1963 2404 1967
rect 2398 1962 2404 1963
rect 2614 1967 2620 1968
rect 2614 1963 2615 1967
rect 2619 1963 2620 1967
rect 2614 1962 2620 1963
rect 2814 1967 2820 1968
rect 2814 1963 2815 1967
rect 2819 1963 2820 1967
rect 2814 1962 2820 1963
rect 2998 1967 3004 1968
rect 2998 1963 2999 1967
rect 3003 1963 3004 1967
rect 2998 1962 3004 1963
rect 3166 1967 3172 1968
rect 3166 1963 3167 1967
rect 3171 1963 3172 1967
rect 3166 1962 3172 1963
rect 3334 1967 3340 1968
rect 3334 1963 3335 1967
rect 3339 1963 3340 1967
rect 3334 1962 3340 1963
rect 3478 1967 3484 1968
rect 3478 1963 3479 1967
rect 3483 1963 3484 1967
rect 3478 1962 3484 1963
rect 1598 1958 1604 1959
rect 3258 1959 3264 1960
rect 1862 1957 1868 1958
rect 386 1955 392 1956
rect 110 1953 116 1954
rect 110 1949 111 1953
rect 115 1949 116 1953
rect 386 1951 387 1955
rect 391 1954 392 1955
rect 1310 1955 1316 1956
rect 1310 1954 1311 1955
rect 391 1952 457 1954
rect 728 1952 737 1954
rect 1297 1952 1311 1954
rect 391 1951 392 1952
rect 386 1950 392 1951
rect 726 1951 732 1952
rect 110 1948 116 1949
rect 726 1947 727 1951
rect 731 1947 732 1951
rect 1310 1951 1311 1952
rect 1315 1951 1316 1955
rect 1310 1950 1316 1951
rect 1822 1953 1828 1954
rect 1822 1949 1823 1953
rect 1827 1949 1828 1953
rect 1862 1953 1863 1957
rect 1867 1953 1868 1957
rect 3258 1955 3259 1959
rect 3263 1958 3264 1959
rect 3263 1956 3353 1958
rect 3574 1957 3580 1958
rect 3263 1955 3264 1956
rect 3258 1954 3264 1955
rect 1862 1952 1868 1953
rect 3574 1953 3575 1957
rect 3579 1953 3580 1957
rect 3574 1952 3580 1953
rect 1822 1948 1828 1949
rect 726 1946 732 1947
rect 2010 1943 2016 1944
rect 2010 1942 2011 1943
rect 1862 1940 1868 1941
rect 1965 1940 2011 1942
rect 287 1939 293 1940
rect 287 1938 288 1939
rect 110 1936 116 1937
rect 221 1936 288 1938
rect 110 1932 111 1936
rect 115 1932 116 1936
rect 287 1935 288 1936
rect 292 1935 293 1939
rect 431 1939 437 1940
rect 431 1938 432 1939
rect 357 1936 432 1938
rect 287 1934 293 1935
rect 431 1935 432 1936
rect 436 1935 437 1939
rect 431 1934 437 1935
rect 506 1939 512 1940
rect 506 1935 507 1939
rect 511 1938 512 1939
rect 786 1939 792 1940
rect 511 1936 609 1938
rect 511 1935 512 1936
rect 506 1934 512 1935
rect 786 1935 787 1939
rect 791 1938 792 1939
rect 922 1939 928 1940
rect 791 1936 881 1938
rect 791 1935 792 1936
rect 786 1934 792 1935
rect 922 1935 923 1939
rect 927 1938 928 1939
rect 1231 1939 1237 1940
rect 1231 1938 1232 1939
rect 927 1936 1017 1938
rect 1181 1936 1232 1938
rect 927 1935 928 1936
rect 922 1934 928 1935
rect 1231 1935 1232 1936
rect 1236 1935 1237 1939
rect 1231 1934 1237 1935
rect 1306 1939 1312 1940
rect 1306 1935 1307 1939
rect 1311 1938 1312 1939
rect 1426 1939 1432 1940
rect 1311 1936 1385 1938
rect 1311 1935 1312 1936
rect 1306 1934 1312 1935
rect 1426 1935 1427 1939
rect 1431 1938 1432 1939
rect 1546 1939 1552 1940
rect 1431 1936 1505 1938
rect 1431 1935 1432 1936
rect 1426 1934 1432 1935
rect 1546 1935 1547 1939
rect 1551 1938 1552 1939
rect 1551 1936 1625 1938
rect 1822 1936 1828 1937
rect 1551 1935 1552 1936
rect 1546 1934 1552 1935
rect 110 1931 116 1932
rect 1822 1932 1823 1936
rect 1827 1932 1828 1936
rect 1862 1936 1863 1940
rect 1867 1936 1868 1940
rect 2010 1939 2011 1940
rect 2015 1939 2016 1943
rect 2391 1943 2397 1944
rect 2391 1942 2392 1943
rect 2221 1940 2392 1942
rect 2010 1938 2016 1939
rect 2391 1939 2392 1940
rect 2396 1939 2397 1943
rect 2607 1943 2613 1944
rect 2607 1942 2608 1943
rect 2461 1940 2608 1942
rect 2391 1938 2397 1939
rect 2607 1939 2608 1940
rect 2612 1939 2613 1943
rect 2807 1943 2813 1944
rect 2807 1942 2808 1943
rect 2677 1940 2808 1942
rect 2607 1938 2613 1939
rect 2807 1939 2808 1940
rect 2812 1939 2813 1943
rect 2991 1943 2997 1944
rect 2991 1942 2992 1943
rect 2877 1940 2992 1942
rect 2807 1938 2813 1939
rect 2991 1939 2992 1940
rect 2996 1939 2997 1943
rect 3159 1943 3165 1944
rect 3159 1942 3160 1943
rect 3061 1940 3160 1942
rect 2991 1938 2997 1939
rect 3159 1939 3160 1940
rect 3164 1939 3165 1943
rect 3327 1943 3333 1944
rect 3327 1942 3328 1943
rect 3229 1940 3328 1942
rect 3159 1938 3165 1939
rect 3327 1939 3328 1940
rect 3332 1939 3333 1943
rect 3546 1943 3552 1944
rect 3546 1942 3547 1943
rect 3541 1940 3547 1942
rect 3327 1938 3333 1939
rect 3546 1939 3547 1940
rect 3551 1939 3552 1943
rect 3546 1938 3552 1939
rect 3574 1940 3580 1941
rect 1862 1935 1868 1936
rect 3574 1936 3575 1940
rect 3579 1936 3580 1940
rect 3574 1935 3580 1936
rect 1822 1931 1828 1932
rect 1910 1927 1916 1928
rect 166 1923 172 1924
rect 166 1919 167 1923
rect 171 1919 172 1923
rect 166 1918 172 1919
rect 302 1923 308 1924
rect 302 1919 303 1923
rect 307 1919 308 1923
rect 302 1918 308 1919
rect 446 1923 452 1924
rect 446 1919 447 1923
rect 451 1919 452 1923
rect 446 1918 452 1919
rect 590 1923 596 1924
rect 590 1919 591 1923
rect 595 1919 596 1923
rect 590 1918 596 1919
rect 726 1923 732 1924
rect 726 1919 727 1923
rect 731 1919 732 1923
rect 862 1923 868 1924
rect 726 1918 732 1919
rect 786 1919 792 1920
rect 786 1918 787 1919
rect 736 1916 787 1918
rect 736 1914 738 1916
rect 786 1915 787 1916
rect 791 1915 792 1919
rect 862 1919 863 1923
rect 867 1919 868 1923
rect 862 1918 868 1919
rect 998 1923 1004 1924
rect 998 1919 999 1923
rect 1003 1919 1004 1923
rect 998 1918 1004 1919
rect 1126 1923 1132 1924
rect 1126 1919 1127 1923
rect 1131 1919 1132 1923
rect 1126 1918 1132 1919
rect 1246 1923 1252 1924
rect 1246 1919 1247 1923
rect 1251 1919 1252 1923
rect 1246 1918 1252 1919
rect 1366 1923 1372 1924
rect 1366 1919 1367 1923
rect 1371 1919 1372 1923
rect 1366 1918 1372 1919
rect 1486 1923 1492 1924
rect 1486 1919 1487 1923
rect 1491 1919 1492 1923
rect 1486 1918 1492 1919
rect 1606 1923 1612 1924
rect 1606 1919 1607 1923
rect 1611 1919 1612 1923
rect 1910 1923 1911 1927
rect 1915 1923 1916 1927
rect 1910 1922 1916 1923
rect 2166 1927 2172 1928
rect 2166 1923 2167 1927
rect 2171 1923 2172 1927
rect 2166 1922 2172 1923
rect 2406 1927 2412 1928
rect 2406 1923 2407 1927
rect 2411 1923 2412 1927
rect 2406 1922 2412 1923
rect 2622 1927 2628 1928
rect 2622 1923 2623 1927
rect 2627 1923 2628 1927
rect 2622 1922 2628 1923
rect 2822 1927 2828 1928
rect 2822 1923 2823 1927
rect 2827 1923 2828 1927
rect 2822 1922 2828 1923
rect 3006 1927 3012 1928
rect 3006 1923 3007 1927
rect 3011 1923 3012 1927
rect 3006 1922 3012 1923
rect 3174 1927 3180 1928
rect 3174 1923 3175 1927
rect 3179 1923 3180 1927
rect 3174 1922 3180 1923
rect 3342 1927 3348 1928
rect 3342 1923 3343 1927
rect 3347 1923 3348 1927
rect 3342 1922 3348 1923
rect 3486 1927 3492 1928
rect 3486 1923 3487 1927
rect 3491 1923 3492 1927
rect 3486 1922 3492 1923
rect 1606 1918 1612 1919
rect 786 1914 792 1915
rect 1939 1915 1948 1916
rect 619 1913 738 1914
rect 195 1911 201 1912
rect 195 1907 196 1911
rect 200 1910 201 1911
rect 206 1911 212 1912
rect 206 1910 207 1911
rect 200 1908 207 1910
rect 200 1907 201 1908
rect 195 1906 201 1907
rect 206 1907 207 1908
rect 211 1907 212 1911
rect 206 1906 212 1907
rect 287 1911 293 1912
rect 287 1907 288 1911
rect 292 1910 293 1911
rect 331 1911 337 1912
rect 331 1910 332 1911
rect 292 1908 332 1910
rect 292 1907 293 1908
rect 287 1906 293 1907
rect 331 1907 332 1908
rect 336 1907 337 1911
rect 331 1906 337 1907
rect 475 1911 481 1912
rect 475 1907 476 1911
rect 480 1910 481 1911
rect 506 1911 512 1912
rect 506 1910 507 1911
rect 480 1908 507 1910
rect 480 1907 481 1908
rect 475 1906 481 1907
rect 506 1907 507 1908
rect 511 1907 512 1911
rect 619 1909 620 1913
rect 624 1912 738 1913
rect 624 1909 625 1912
rect 619 1908 625 1909
rect 755 1911 761 1912
rect 506 1906 512 1907
rect 755 1907 756 1911
rect 760 1910 761 1911
rect 778 1911 784 1912
rect 778 1910 779 1911
rect 760 1908 779 1910
rect 760 1907 761 1908
rect 755 1906 761 1907
rect 778 1907 779 1908
rect 783 1907 784 1911
rect 778 1906 784 1907
rect 891 1911 897 1912
rect 891 1907 892 1911
rect 896 1910 897 1911
rect 922 1911 928 1912
rect 922 1910 923 1911
rect 896 1908 923 1910
rect 896 1907 897 1908
rect 891 1906 897 1907
rect 922 1907 923 1908
rect 927 1907 928 1911
rect 922 1906 928 1907
rect 1014 1911 1020 1912
rect 1014 1907 1015 1911
rect 1019 1910 1020 1911
rect 1027 1911 1033 1912
rect 1027 1910 1028 1911
rect 1019 1908 1028 1910
rect 1019 1907 1020 1908
rect 1014 1906 1020 1907
rect 1027 1907 1028 1908
rect 1032 1907 1033 1911
rect 1027 1906 1033 1907
rect 1155 1911 1161 1912
rect 1155 1907 1156 1911
rect 1160 1910 1161 1911
rect 1231 1911 1237 1912
rect 1160 1908 1226 1910
rect 1160 1907 1161 1908
rect 1155 1906 1161 1907
rect 1224 1902 1226 1908
rect 1231 1907 1232 1911
rect 1236 1910 1237 1911
rect 1275 1911 1281 1912
rect 1275 1910 1276 1911
rect 1236 1908 1276 1910
rect 1236 1907 1237 1908
rect 1231 1906 1237 1907
rect 1275 1907 1276 1908
rect 1280 1907 1281 1911
rect 1275 1906 1281 1907
rect 1395 1911 1401 1912
rect 1395 1907 1396 1911
rect 1400 1910 1401 1911
rect 1426 1911 1432 1912
rect 1426 1910 1427 1911
rect 1400 1908 1427 1910
rect 1400 1907 1401 1908
rect 1395 1906 1401 1907
rect 1426 1907 1427 1908
rect 1431 1907 1432 1911
rect 1426 1906 1432 1907
rect 1515 1911 1521 1912
rect 1515 1907 1516 1911
rect 1520 1910 1521 1911
rect 1546 1911 1552 1912
rect 1546 1910 1547 1911
rect 1520 1908 1547 1910
rect 1520 1907 1521 1908
rect 1515 1906 1521 1907
rect 1546 1907 1547 1908
rect 1551 1907 1552 1911
rect 1546 1906 1552 1907
rect 1635 1911 1641 1912
rect 1635 1907 1636 1911
rect 1640 1910 1641 1911
rect 1666 1911 1672 1912
rect 1666 1910 1667 1911
rect 1640 1908 1667 1910
rect 1640 1907 1641 1908
rect 1635 1906 1641 1907
rect 1666 1907 1667 1908
rect 1671 1907 1672 1911
rect 1939 1911 1940 1915
rect 1947 1911 1948 1915
rect 2194 1915 2201 1916
rect 1939 1910 1948 1911
rect 2055 1911 2061 1912
rect 2055 1910 2056 1911
rect 1666 1906 1672 1907
rect 2004 1908 2056 1910
rect 2004 1906 2006 1908
rect 2055 1907 2056 1908
rect 2060 1907 2061 1911
rect 2194 1911 2195 1915
rect 2200 1911 2201 1915
rect 2194 1910 2201 1911
rect 2391 1915 2397 1916
rect 2391 1911 2392 1915
rect 2396 1914 2397 1915
rect 2435 1915 2441 1916
rect 2435 1914 2436 1915
rect 2396 1912 2436 1914
rect 2396 1911 2397 1912
rect 2391 1910 2397 1911
rect 2435 1911 2436 1912
rect 2440 1911 2441 1915
rect 2435 1910 2441 1911
rect 2651 1915 2660 1916
rect 2651 1911 2652 1915
rect 2659 1911 2660 1915
rect 2651 1910 2660 1911
rect 2807 1915 2813 1916
rect 2807 1911 2808 1915
rect 2812 1914 2813 1915
rect 2851 1915 2857 1916
rect 2851 1914 2852 1915
rect 2812 1912 2852 1914
rect 2812 1911 2813 1912
rect 2807 1910 2813 1911
rect 2851 1911 2852 1912
rect 2856 1911 2857 1915
rect 2851 1910 2857 1911
rect 2991 1915 2997 1916
rect 2991 1911 2992 1915
rect 2996 1914 2997 1915
rect 3035 1915 3041 1916
rect 3035 1914 3036 1915
rect 2996 1912 3036 1914
rect 2996 1911 2997 1912
rect 2991 1910 2997 1911
rect 3035 1911 3036 1912
rect 3040 1911 3041 1915
rect 3035 1910 3041 1911
rect 3159 1915 3165 1916
rect 3159 1911 3160 1915
rect 3164 1914 3165 1915
rect 3203 1915 3209 1916
rect 3203 1914 3204 1915
rect 3164 1912 3204 1914
rect 3164 1911 3165 1912
rect 3159 1910 3165 1911
rect 3203 1911 3204 1912
rect 3208 1911 3209 1915
rect 3203 1910 3209 1911
rect 3327 1915 3333 1916
rect 3327 1911 3328 1915
rect 3332 1914 3333 1915
rect 3371 1915 3377 1916
rect 3371 1914 3372 1915
rect 3332 1912 3372 1914
rect 3332 1911 3333 1912
rect 3327 1910 3333 1911
rect 3371 1911 3372 1912
rect 3376 1911 3377 1915
rect 3371 1910 3377 1911
rect 3515 1915 3521 1916
rect 3515 1911 3516 1915
rect 3520 1914 3521 1915
rect 3554 1915 3560 1916
rect 3554 1914 3555 1915
rect 3520 1912 3555 1914
rect 3520 1911 3521 1912
rect 3515 1910 3521 1911
rect 3554 1911 3555 1912
rect 3559 1911 3560 1915
rect 3554 1910 3560 1911
rect 2055 1906 2061 1907
rect 1923 1905 2006 1906
rect 1306 1903 1312 1904
rect 1306 1902 1307 1903
rect 1224 1900 1307 1902
rect 1306 1899 1307 1900
rect 1311 1899 1312 1903
rect 1923 1901 1924 1905
rect 1928 1904 2006 1905
rect 1928 1901 1929 1904
rect 1923 1900 1929 1901
rect 2010 1903 2017 1904
rect 1306 1898 1312 1899
rect 2010 1899 2011 1903
rect 2016 1899 2017 1903
rect 2010 1898 2017 1899
rect 2047 1903 2053 1904
rect 2047 1899 2048 1903
rect 2052 1902 2053 1903
rect 2099 1903 2105 1904
rect 2099 1902 2100 1903
rect 2052 1900 2100 1902
rect 2052 1899 2053 1900
rect 2047 1898 2053 1899
rect 2099 1899 2100 1900
rect 2104 1899 2105 1903
rect 2099 1898 2105 1899
rect 2110 1903 2116 1904
rect 2110 1899 2111 1903
rect 2115 1902 2116 1903
rect 2195 1903 2201 1904
rect 2195 1902 2196 1903
rect 2115 1900 2196 1902
rect 2115 1899 2116 1900
rect 2110 1898 2116 1899
rect 2195 1899 2196 1900
rect 2200 1899 2201 1903
rect 2195 1898 2201 1899
rect 2247 1903 2253 1904
rect 2247 1899 2248 1903
rect 2252 1902 2253 1903
rect 2323 1903 2329 1904
rect 2323 1902 2324 1903
rect 2252 1900 2324 1902
rect 2252 1899 2253 1900
rect 2247 1898 2253 1899
rect 2323 1899 2324 1900
rect 2328 1899 2329 1903
rect 2323 1898 2329 1899
rect 2391 1903 2397 1904
rect 2391 1899 2392 1903
rect 2396 1902 2397 1903
rect 2475 1903 2481 1904
rect 2475 1902 2476 1903
rect 2396 1900 2476 1902
rect 2396 1899 2397 1900
rect 2391 1898 2397 1899
rect 2475 1899 2476 1900
rect 2480 1899 2481 1903
rect 2475 1898 2481 1899
rect 2607 1903 2613 1904
rect 2607 1899 2608 1903
rect 2612 1902 2613 1903
rect 2635 1903 2641 1904
rect 2635 1902 2636 1903
rect 2612 1900 2636 1902
rect 2612 1899 2613 1900
rect 2607 1898 2613 1899
rect 2635 1899 2636 1900
rect 2640 1899 2641 1903
rect 2635 1898 2641 1899
rect 2695 1903 2701 1904
rect 2695 1899 2696 1903
rect 2700 1902 2701 1903
rect 2795 1903 2801 1904
rect 2795 1902 2796 1903
rect 2700 1900 2796 1902
rect 2700 1899 2701 1900
rect 2695 1898 2701 1899
rect 2795 1899 2796 1900
rect 2800 1899 2801 1903
rect 2795 1898 2801 1899
rect 2947 1903 2956 1904
rect 2947 1899 2948 1903
rect 2955 1899 2956 1903
rect 2947 1898 2956 1899
rect 3015 1903 3021 1904
rect 3015 1899 3016 1903
rect 3020 1902 3021 1903
rect 3099 1903 3105 1904
rect 3099 1902 3100 1903
rect 3020 1900 3100 1902
rect 3020 1899 3021 1900
rect 3015 1898 3021 1899
rect 3099 1899 3100 1900
rect 3104 1899 3105 1903
rect 3099 1898 3105 1899
rect 3159 1903 3165 1904
rect 3159 1899 3160 1903
rect 3164 1902 3165 1903
rect 3243 1903 3249 1904
rect 3243 1902 3244 1903
rect 3164 1900 3244 1902
rect 3164 1899 3165 1900
rect 3159 1898 3165 1899
rect 3243 1899 3244 1900
rect 3248 1899 3249 1903
rect 3243 1898 3249 1899
rect 3387 1903 3393 1904
rect 3387 1899 3388 1903
rect 3392 1902 3393 1903
rect 3426 1903 3432 1904
rect 3426 1902 3427 1903
rect 3392 1900 3427 1902
rect 3392 1899 3393 1900
rect 3387 1898 3393 1899
rect 3426 1899 3427 1900
rect 3431 1899 3432 1903
rect 3426 1898 3432 1899
rect 3515 1903 3521 1904
rect 3515 1899 3516 1903
rect 3520 1902 3521 1903
rect 3546 1903 3552 1904
rect 3546 1902 3547 1903
rect 3520 1900 3547 1902
rect 3520 1899 3521 1900
rect 3515 1898 3521 1899
rect 3546 1899 3547 1900
rect 3551 1899 3552 1903
rect 3546 1898 3552 1899
rect 1894 1893 1900 1894
rect 251 1891 257 1892
rect 251 1887 252 1891
rect 256 1890 257 1891
rect 319 1891 325 1892
rect 319 1890 320 1891
rect 256 1888 320 1890
rect 256 1887 257 1888
rect 251 1886 257 1887
rect 319 1887 320 1888
rect 324 1887 325 1891
rect 319 1886 325 1887
rect 431 1891 437 1892
rect 431 1887 432 1891
rect 436 1890 437 1891
rect 507 1891 513 1892
rect 507 1890 508 1891
rect 436 1888 508 1890
rect 436 1887 437 1888
rect 431 1886 437 1887
rect 507 1887 508 1888
rect 512 1887 513 1891
rect 507 1886 513 1887
rect 747 1891 756 1892
rect 747 1887 748 1891
rect 755 1887 756 1891
rect 747 1886 756 1887
rect 963 1891 969 1892
rect 963 1887 964 1891
rect 968 1890 969 1891
rect 1030 1891 1036 1892
rect 1030 1890 1031 1891
rect 968 1888 1031 1890
rect 968 1887 969 1888
rect 963 1886 969 1887
rect 1030 1887 1031 1888
rect 1035 1887 1036 1891
rect 1030 1886 1036 1887
rect 1039 1891 1045 1892
rect 1039 1887 1040 1891
rect 1044 1890 1045 1891
rect 1155 1891 1161 1892
rect 1155 1890 1156 1891
rect 1044 1888 1156 1890
rect 1044 1887 1045 1888
rect 1039 1886 1045 1887
rect 1155 1887 1156 1888
rect 1160 1887 1161 1891
rect 1155 1886 1161 1887
rect 1231 1891 1237 1892
rect 1231 1887 1232 1891
rect 1236 1890 1237 1891
rect 1323 1891 1329 1892
rect 1323 1890 1324 1891
rect 1236 1888 1324 1890
rect 1236 1887 1237 1888
rect 1231 1886 1237 1887
rect 1323 1887 1324 1888
rect 1328 1887 1329 1891
rect 1323 1886 1329 1887
rect 1391 1891 1397 1892
rect 1391 1887 1392 1891
rect 1396 1890 1397 1891
rect 1483 1891 1489 1892
rect 1483 1890 1484 1891
rect 1396 1888 1484 1890
rect 1396 1887 1397 1888
rect 1391 1886 1397 1887
rect 1483 1887 1484 1888
rect 1488 1887 1489 1891
rect 1483 1886 1489 1887
rect 1551 1891 1557 1892
rect 1551 1887 1552 1891
rect 1556 1890 1557 1891
rect 1635 1891 1641 1892
rect 1635 1890 1636 1891
rect 1556 1888 1636 1890
rect 1556 1887 1557 1888
rect 1551 1886 1557 1887
rect 1635 1887 1636 1888
rect 1640 1887 1641 1891
rect 1635 1886 1641 1887
rect 1763 1891 1769 1892
rect 1763 1887 1764 1891
rect 1768 1890 1769 1891
rect 1768 1888 1874 1890
rect 1894 1889 1895 1893
rect 1899 1889 1900 1893
rect 1894 1888 1900 1889
rect 1982 1893 1988 1894
rect 1982 1889 1983 1893
rect 1987 1889 1988 1893
rect 1982 1888 1988 1889
rect 2070 1893 2076 1894
rect 2070 1889 2071 1893
rect 2075 1889 2076 1893
rect 2070 1888 2076 1889
rect 2166 1893 2172 1894
rect 2166 1889 2167 1893
rect 2171 1889 2172 1893
rect 2166 1888 2172 1889
rect 2294 1893 2300 1894
rect 2294 1889 2295 1893
rect 2299 1889 2300 1893
rect 2294 1888 2300 1889
rect 2446 1893 2452 1894
rect 2446 1889 2447 1893
rect 2451 1889 2452 1893
rect 2446 1888 2452 1889
rect 2606 1893 2612 1894
rect 2606 1889 2607 1893
rect 2611 1889 2612 1893
rect 2606 1888 2612 1889
rect 2766 1893 2772 1894
rect 2766 1889 2767 1893
rect 2771 1889 2772 1893
rect 2766 1888 2772 1889
rect 2918 1893 2924 1894
rect 2918 1889 2919 1893
rect 2923 1889 2924 1893
rect 2918 1888 2924 1889
rect 3070 1893 3076 1894
rect 3070 1889 3071 1893
rect 3075 1889 3076 1893
rect 3070 1888 3076 1889
rect 3214 1893 3220 1894
rect 3214 1889 3215 1893
rect 3219 1889 3220 1893
rect 3214 1888 3220 1889
rect 3358 1893 3364 1894
rect 3358 1889 3359 1893
rect 3363 1889 3364 1893
rect 3358 1888 3364 1889
rect 3486 1893 3492 1894
rect 3486 1889 3487 1893
rect 3491 1889 3492 1893
rect 3486 1888 3492 1889
rect 1768 1887 1769 1888
rect 1763 1886 1769 1887
rect 222 1881 228 1882
rect 222 1877 223 1881
rect 227 1877 228 1881
rect 222 1876 228 1877
rect 478 1881 484 1882
rect 478 1877 479 1881
rect 483 1877 484 1881
rect 478 1876 484 1877
rect 718 1881 724 1882
rect 718 1877 719 1881
rect 723 1877 724 1881
rect 718 1876 724 1877
rect 934 1881 940 1882
rect 934 1877 935 1881
rect 939 1877 940 1881
rect 934 1876 940 1877
rect 1126 1881 1132 1882
rect 1126 1877 1127 1881
rect 1131 1877 1132 1881
rect 1126 1876 1132 1877
rect 1294 1881 1300 1882
rect 1294 1877 1295 1881
rect 1299 1877 1300 1881
rect 1294 1876 1300 1877
rect 1454 1881 1460 1882
rect 1454 1877 1455 1881
rect 1459 1877 1460 1881
rect 1454 1876 1460 1877
rect 1606 1881 1612 1882
rect 1606 1877 1607 1881
rect 1611 1877 1612 1881
rect 1606 1876 1612 1877
rect 1734 1881 1740 1882
rect 1734 1877 1735 1881
rect 1739 1877 1740 1881
rect 1734 1876 1740 1877
rect 1862 1880 1868 1881
rect 1862 1876 1863 1880
rect 1867 1876 1868 1880
rect 1862 1875 1868 1876
rect 1872 1874 1874 1888
rect 3574 1880 3580 1881
rect 2047 1879 2053 1880
rect 2047 1878 2048 1879
rect 2037 1876 2048 1878
rect 2047 1875 2048 1876
rect 2052 1875 2053 1879
rect 2247 1879 2253 1880
rect 2247 1878 2248 1879
rect 2221 1876 2248 1878
rect 2047 1874 2053 1875
rect 2055 1875 2061 1876
rect 1872 1872 1913 1874
rect 2055 1871 2056 1875
rect 2060 1874 2061 1875
rect 2247 1875 2248 1876
rect 2252 1875 2253 1879
rect 2391 1879 2397 1880
rect 2391 1878 2392 1879
rect 2349 1876 2392 1878
rect 2247 1874 2253 1875
rect 2391 1875 2392 1876
rect 2396 1875 2397 1879
rect 2695 1879 2701 1880
rect 2695 1878 2696 1879
rect 2661 1876 2696 1878
rect 2391 1874 2397 1875
rect 2402 1875 2408 1876
rect 2060 1872 2089 1874
rect 2060 1871 2061 1872
rect 2055 1870 2061 1871
rect 2402 1871 2403 1875
rect 2407 1874 2408 1875
rect 2695 1875 2696 1876
rect 2700 1875 2701 1879
rect 3015 1879 3021 1880
rect 3015 1878 3016 1879
rect 2973 1876 3016 1878
rect 2695 1874 2701 1875
rect 3015 1875 3016 1876
rect 3020 1875 3021 1879
rect 3159 1879 3165 1880
rect 3159 1878 3160 1879
rect 3125 1876 3160 1878
rect 3015 1874 3021 1875
rect 3159 1875 3160 1876
rect 3164 1875 3165 1879
rect 3418 1879 3424 1880
rect 3418 1878 3419 1879
rect 3413 1876 3419 1878
rect 3159 1874 3165 1875
rect 3418 1875 3419 1876
rect 3423 1875 3424 1879
rect 3574 1876 3575 1880
rect 3579 1876 3580 1880
rect 3418 1874 3424 1875
rect 3426 1875 3432 1876
rect 3574 1875 3580 1876
rect 2407 1872 2465 1874
rect 2407 1871 2408 1872
rect 2402 1870 2408 1871
rect 3426 1871 3427 1875
rect 3431 1874 3432 1875
rect 3431 1872 3505 1874
rect 3431 1871 3432 1872
rect 3426 1870 3432 1871
rect 110 1868 116 1869
rect 1822 1868 1828 1869
rect 110 1864 111 1868
rect 115 1864 116 1868
rect 778 1867 784 1868
rect 778 1866 779 1867
rect 773 1864 779 1866
rect 110 1863 116 1864
rect 319 1863 325 1864
rect 319 1859 320 1863
rect 324 1862 325 1863
rect 778 1863 779 1864
rect 783 1863 784 1867
rect 1039 1867 1045 1868
rect 1039 1866 1040 1867
rect 989 1864 1040 1866
rect 778 1862 784 1863
rect 1039 1863 1040 1864
rect 1044 1863 1045 1867
rect 1231 1867 1237 1868
rect 1231 1866 1232 1867
rect 1181 1864 1232 1866
rect 1039 1862 1045 1863
rect 1231 1863 1232 1864
rect 1236 1863 1237 1867
rect 1391 1867 1397 1868
rect 1391 1866 1392 1867
rect 1349 1864 1392 1866
rect 1231 1862 1237 1863
rect 1391 1863 1392 1864
rect 1396 1863 1397 1867
rect 1551 1867 1557 1868
rect 1551 1866 1552 1867
rect 1509 1864 1552 1866
rect 1391 1862 1397 1863
rect 1551 1863 1552 1864
rect 1556 1863 1557 1867
rect 1666 1867 1672 1868
rect 1666 1866 1667 1867
rect 1661 1864 1667 1866
rect 1551 1862 1557 1863
rect 1666 1863 1667 1864
rect 1671 1863 1672 1867
rect 1822 1864 1823 1868
rect 1827 1864 1828 1868
rect 1822 1863 1828 1864
rect 1862 1863 1868 1864
rect 1666 1862 1672 1863
rect 324 1860 497 1862
rect 324 1859 325 1860
rect 319 1858 325 1859
rect 1862 1859 1863 1863
rect 1867 1859 1868 1863
rect 1862 1858 1868 1859
rect 2674 1863 2680 1864
rect 2674 1859 2675 1863
rect 2679 1862 2680 1863
rect 3335 1863 3341 1864
rect 3335 1862 3336 1863
rect 2679 1860 2777 1862
rect 3265 1860 3336 1862
rect 2679 1859 2680 1860
rect 2674 1858 2680 1859
rect 3335 1859 3336 1860
rect 3340 1859 3341 1863
rect 3335 1858 3341 1859
rect 3574 1863 3580 1864
rect 3574 1859 3575 1863
rect 3579 1859 3580 1863
rect 3574 1858 3580 1859
rect 1886 1853 1892 1854
rect 110 1851 116 1852
rect 110 1847 111 1851
rect 115 1847 116 1851
rect 110 1846 116 1847
rect 1822 1851 1828 1852
rect 1822 1847 1823 1851
rect 1827 1847 1828 1851
rect 1886 1849 1887 1853
rect 1891 1849 1892 1853
rect 1886 1848 1892 1849
rect 1974 1853 1980 1854
rect 1974 1849 1975 1853
rect 1979 1849 1980 1853
rect 1974 1848 1980 1849
rect 2062 1853 2068 1854
rect 2062 1849 2063 1853
rect 2067 1849 2068 1853
rect 2062 1848 2068 1849
rect 2158 1853 2164 1854
rect 2158 1849 2159 1853
rect 2163 1849 2164 1853
rect 2158 1848 2164 1849
rect 2286 1853 2292 1854
rect 2286 1849 2287 1853
rect 2291 1849 2292 1853
rect 2286 1848 2292 1849
rect 2438 1853 2444 1854
rect 2438 1849 2439 1853
rect 2443 1849 2444 1853
rect 2438 1848 2444 1849
rect 2598 1853 2604 1854
rect 2598 1849 2599 1853
rect 2603 1849 2604 1853
rect 2598 1848 2604 1849
rect 2758 1853 2764 1854
rect 2758 1849 2759 1853
rect 2763 1849 2764 1853
rect 2758 1848 2764 1849
rect 2910 1853 2916 1854
rect 2910 1849 2911 1853
rect 2915 1849 2916 1853
rect 2910 1848 2916 1849
rect 3062 1853 3068 1854
rect 3062 1849 3063 1853
rect 3067 1849 3068 1853
rect 3062 1848 3068 1849
rect 3206 1853 3212 1854
rect 3206 1849 3207 1853
rect 3211 1849 3212 1853
rect 3206 1848 3212 1849
rect 3350 1853 3356 1854
rect 3350 1849 3351 1853
rect 3355 1849 3356 1853
rect 3350 1848 3356 1849
rect 3478 1853 3484 1854
rect 3478 1849 3479 1853
rect 3483 1849 3484 1853
rect 3478 1848 3484 1849
rect 1822 1846 1828 1847
rect 214 1841 220 1842
rect 214 1837 215 1841
rect 219 1837 220 1841
rect 214 1836 220 1837
rect 470 1841 476 1842
rect 470 1837 471 1841
rect 475 1837 476 1841
rect 470 1836 476 1837
rect 710 1841 716 1842
rect 710 1837 711 1841
rect 715 1837 716 1841
rect 710 1836 716 1837
rect 926 1841 932 1842
rect 926 1837 927 1841
rect 931 1837 932 1841
rect 926 1836 932 1837
rect 1118 1841 1124 1842
rect 1118 1837 1119 1841
rect 1123 1837 1124 1841
rect 1118 1836 1124 1837
rect 1286 1841 1292 1842
rect 1286 1837 1287 1841
rect 1291 1837 1292 1841
rect 1286 1836 1292 1837
rect 1446 1841 1452 1842
rect 1446 1837 1447 1841
rect 1451 1837 1452 1841
rect 1446 1836 1452 1837
rect 1598 1841 1604 1842
rect 1598 1837 1599 1841
rect 1603 1837 1604 1841
rect 1598 1836 1604 1837
rect 1726 1841 1732 1842
rect 1726 1837 1727 1841
rect 1731 1837 1732 1841
rect 1726 1836 1732 1837
rect 263 1835 269 1836
rect 263 1831 264 1835
rect 268 1834 269 1835
rect 282 1835 288 1836
rect 282 1834 283 1835
rect 268 1832 283 1834
rect 268 1831 269 1832
rect 263 1830 269 1831
rect 282 1831 283 1832
rect 287 1831 288 1835
rect 282 1830 288 1831
rect 1766 1835 1772 1836
rect 1766 1831 1767 1835
rect 1771 1834 1772 1835
rect 1775 1835 1781 1836
rect 1775 1834 1776 1835
rect 1771 1832 1776 1834
rect 1771 1831 1772 1832
rect 1766 1830 1772 1831
rect 1775 1831 1776 1832
rect 1780 1831 1781 1835
rect 1775 1830 1781 1831
rect 1998 1827 2004 1828
rect 1998 1823 1999 1827
rect 2003 1823 2004 1827
rect 1998 1822 2004 1823
rect 2222 1827 2228 1828
rect 2222 1823 2223 1827
rect 2227 1823 2228 1827
rect 2222 1822 2228 1823
rect 2438 1827 2444 1828
rect 2438 1823 2439 1827
rect 2443 1823 2444 1827
rect 2438 1822 2444 1823
rect 2638 1827 2644 1828
rect 2638 1823 2639 1827
rect 2643 1823 2644 1827
rect 2638 1822 2644 1823
rect 2830 1827 2836 1828
rect 2830 1823 2831 1827
rect 2835 1823 2836 1827
rect 2830 1822 2836 1823
rect 3014 1827 3020 1828
rect 3014 1823 3015 1827
rect 3019 1823 3020 1827
rect 3014 1822 3020 1823
rect 3198 1827 3204 1828
rect 3198 1823 3199 1827
rect 3203 1823 3204 1827
rect 3198 1822 3204 1823
rect 3390 1827 3396 1828
rect 3390 1823 3391 1827
rect 3395 1823 3396 1827
rect 3390 1822 3396 1823
rect 246 1819 252 1820
rect 246 1815 247 1819
rect 251 1815 252 1819
rect 246 1814 252 1815
rect 414 1819 420 1820
rect 414 1815 415 1819
rect 419 1815 420 1819
rect 414 1814 420 1815
rect 590 1819 596 1820
rect 590 1815 591 1819
rect 595 1815 596 1819
rect 590 1814 596 1815
rect 758 1819 764 1820
rect 758 1815 759 1819
rect 763 1815 764 1819
rect 758 1814 764 1815
rect 926 1819 932 1820
rect 926 1815 927 1819
rect 931 1815 932 1819
rect 926 1814 932 1815
rect 1078 1819 1084 1820
rect 1078 1815 1079 1819
rect 1083 1815 1084 1819
rect 1078 1814 1084 1815
rect 1222 1819 1228 1820
rect 1222 1815 1223 1819
rect 1227 1815 1228 1819
rect 1222 1814 1228 1815
rect 1358 1819 1364 1820
rect 1358 1815 1359 1819
rect 1363 1815 1364 1819
rect 1358 1814 1364 1815
rect 1486 1819 1492 1820
rect 1486 1815 1487 1819
rect 1491 1815 1492 1819
rect 1486 1814 1492 1815
rect 1614 1819 1620 1820
rect 1614 1815 1615 1819
rect 1619 1815 1620 1819
rect 1614 1814 1620 1815
rect 1726 1819 1732 1820
rect 1726 1815 1727 1819
rect 1731 1815 1732 1819
rect 2110 1819 2116 1820
rect 2110 1818 2111 1819
rect 1726 1814 1732 1815
rect 1862 1817 1868 1818
rect 1862 1813 1863 1817
rect 1867 1813 1868 1817
rect 2057 1816 2111 1818
rect 2110 1815 2111 1816
rect 2115 1815 2116 1819
rect 2110 1814 2116 1815
rect 2718 1819 2724 1820
rect 2718 1815 2719 1819
rect 2723 1818 2724 1819
rect 2723 1816 2849 1818
rect 3574 1817 3580 1818
rect 2723 1815 2724 1816
rect 2718 1814 2724 1815
rect 1862 1812 1868 1813
rect 3574 1813 3575 1817
rect 3579 1813 3580 1817
rect 3574 1812 3580 1813
rect 750 1811 756 1812
rect 110 1809 116 1810
rect 110 1805 111 1809
rect 115 1805 116 1809
rect 750 1807 751 1811
rect 755 1810 756 1811
rect 1030 1811 1036 1812
rect 755 1808 777 1810
rect 755 1807 756 1808
rect 750 1806 756 1807
rect 1030 1807 1031 1811
rect 1035 1810 1036 1811
rect 1035 1808 1097 1810
rect 1822 1809 1828 1810
rect 1035 1807 1036 1808
rect 1030 1806 1036 1807
rect 110 1804 116 1805
rect 1822 1805 1823 1809
rect 1827 1805 1828 1809
rect 1822 1804 1828 1805
rect 2431 1803 2437 1804
rect 2431 1802 2432 1803
rect 1862 1800 1868 1801
rect 2285 1800 2432 1802
rect 1862 1796 1863 1800
rect 1867 1796 1868 1800
rect 2431 1799 2432 1800
rect 2436 1799 2437 1803
rect 2631 1803 2637 1804
rect 2631 1802 2632 1803
rect 2501 1800 2632 1802
rect 2431 1798 2437 1799
rect 2631 1799 2632 1800
rect 2636 1799 2637 1803
rect 2818 1803 2824 1804
rect 2818 1802 2819 1803
rect 2701 1800 2819 1802
rect 2631 1798 2637 1799
rect 2818 1799 2819 1800
rect 2823 1799 2824 1803
rect 2818 1798 2824 1799
rect 2898 1803 2904 1804
rect 2898 1799 2899 1803
rect 2903 1802 2904 1803
rect 3082 1803 3088 1804
rect 2903 1800 3041 1802
rect 2903 1799 2904 1800
rect 2898 1798 2904 1799
rect 3082 1799 3083 1803
rect 3087 1802 3088 1803
rect 3458 1803 3464 1804
rect 3458 1802 3459 1803
rect 3087 1800 3225 1802
rect 3453 1800 3459 1802
rect 3087 1799 3088 1800
rect 3082 1798 3088 1799
rect 3458 1799 3459 1800
rect 3463 1799 3464 1803
rect 3458 1798 3464 1799
rect 3574 1800 3580 1801
rect 407 1795 413 1796
rect 407 1794 408 1795
rect 110 1792 116 1793
rect 309 1792 408 1794
rect 110 1788 111 1792
rect 115 1788 116 1792
rect 407 1791 408 1792
rect 412 1791 413 1795
rect 574 1795 580 1796
rect 574 1794 575 1795
rect 477 1792 575 1794
rect 407 1790 413 1791
rect 574 1791 575 1792
rect 579 1791 580 1795
rect 658 1795 664 1796
rect 658 1794 659 1795
rect 653 1792 659 1794
rect 574 1790 580 1791
rect 658 1791 659 1792
rect 663 1791 664 1795
rect 658 1790 664 1791
rect 826 1795 832 1796
rect 826 1791 827 1795
rect 831 1794 832 1795
rect 1146 1795 1152 1796
rect 831 1792 953 1794
rect 831 1791 832 1792
rect 826 1790 832 1791
rect 1146 1791 1147 1795
rect 1151 1794 1152 1795
rect 1290 1795 1296 1796
rect 1151 1792 1249 1794
rect 1151 1791 1152 1792
rect 1146 1790 1152 1791
rect 1290 1791 1291 1795
rect 1295 1794 1296 1795
rect 1554 1795 1560 1796
rect 1295 1792 1385 1794
rect 1295 1791 1296 1792
rect 1290 1790 1296 1791
rect 110 1787 116 1788
rect 1548 1786 1550 1793
rect 1554 1791 1555 1795
rect 1559 1794 1560 1795
rect 1682 1795 1688 1796
rect 1862 1795 1868 1796
rect 3574 1796 3575 1800
rect 3579 1796 3580 1800
rect 3574 1795 3580 1796
rect 1559 1792 1641 1794
rect 1559 1791 1560 1792
rect 1554 1790 1560 1791
rect 1682 1791 1683 1795
rect 1687 1794 1688 1795
rect 1687 1792 1753 1794
rect 1822 1792 1828 1793
rect 1687 1791 1688 1792
rect 1682 1790 1688 1791
rect 1822 1788 1823 1792
rect 1827 1788 1828 1792
rect 1562 1787 1568 1788
rect 1822 1787 1828 1788
rect 2006 1787 2012 1788
rect 1562 1786 1563 1787
rect 1548 1784 1563 1786
rect 1562 1783 1563 1784
rect 1567 1783 1568 1787
rect 1562 1782 1568 1783
rect 2006 1783 2007 1787
rect 2011 1783 2012 1787
rect 2006 1782 2012 1783
rect 2230 1787 2236 1788
rect 2230 1783 2231 1787
rect 2235 1783 2236 1787
rect 2230 1782 2236 1783
rect 2446 1787 2452 1788
rect 2446 1783 2447 1787
rect 2451 1783 2452 1787
rect 2446 1782 2452 1783
rect 2646 1787 2652 1788
rect 2646 1783 2647 1787
rect 2651 1783 2652 1787
rect 2646 1782 2652 1783
rect 2838 1787 2844 1788
rect 2838 1783 2839 1787
rect 2843 1783 2844 1787
rect 2838 1782 2844 1783
rect 3022 1787 3028 1788
rect 3022 1783 3023 1787
rect 3027 1783 3028 1787
rect 3022 1782 3028 1783
rect 3206 1787 3212 1788
rect 3206 1783 3207 1787
rect 3211 1783 3212 1787
rect 3206 1782 3212 1783
rect 3398 1787 3404 1788
rect 3398 1783 3399 1787
rect 3403 1783 3404 1787
rect 3398 1782 3404 1783
rect 254 1779 260 1780
rect 254 1775 255 1779
rect 259 1775 260 1779
rect 254 1774 260 1775
rect 422 1779 428 1780
rect 422 1775 423 1779
rect 427 1775 428 1779
rect 422 1774 428 1775
rect 598 1779 604 1780
rect 598 1775 599 1779
rect 603 1775 604 1779
rect 598 1774 604 1775
rect 766 1779 772 1780
rect 766 1775 767 1779
rect 771 1775 772 1779
rect 766 1774 772 1775
rect 934 1779 940 1780
rect 934 1775 935 1779
rect 939 1775 940 1779
rect 934 1774 940 1775
rect 1086 1779 1092 1780
rect 1086 1775 1087 1779
rect 1091 1775 1092 1779
rect 1086 1774 1092 1775
rect 1230 1779 1236 1780
rect 1230 1775 1231 1779
rect 1235 1775 1236 1779
rect 1230 1774 1236 1775
rect 1366 1779 1372 1780
rect 1366 1775 1367 1779
rect 1371 1775 1372 1779
rect 1366 1774 1372 1775
rect 1494 1779 1500 1780
rect 1494 1775 1495 1779
rect 1499 1775 1500 1779
rect 1494 1774 1500 1775
rect 1622 1779 1628 1780
rect 1622 1775 1623 1779
rect 1627 1775 1628 1779
rect 1622 1774 1628 1775
rect 1734 1779 1740 1780
rect 1734 1775 1735 1779
rect 1739 1775 1740 1779
rect 1734 1774 1740 1775
rect 2007 1775 2013 1776
rect 2007 1771 2008 1775
rect 2012 1774 2013 1775
rect 2035 1775 2041 1776
rect 2035 1774 2036 1775
rect 2012 1772 2036 1774
rect 2012 1771 2013 1772
rect 2007 1770 2013 1771
rect 2035 1771 2036 1772
rect 2040 1771 2041 1775
rect 2035 1770 2041 1771
rect 2259 1775 2268 1776
rect 2259 1771 2260 1775
rect 2267 1771 2268 1775
rect 2259 1770 2268 1771
rect 2475 1775 2484 1776
rect 2475 1771 2476 1775
rect 2483 1771 2484 1775
rect 2475 1770 2484 1771
rect 2631 1775 2637 1776
rect 2631 1771 2632 1775
rect 2636 1774 2637 1775
rect 2675 1775 2681 1776
rect 2675 1774 2676 1775
rect 2636 1772 2676 1774
rect 2636 1771 2637 1772
rect 2631 1770 2637 1771
rect 2675 1771 2676 1772
rect 2680 1771 2681 1775
rect 2675 1770 2681 1771
rect 2867 1775 2873 1776
rect 2867 1771 2868 1775
rect 2872 1774 2873 1775
rect 2898 1775 2904 1776
rect 2898 1774 2899 1775
rect 2872 1772 2899 1774
rect 2872 1771 2873 1772
rect 2867 1770 2873 1771
rect 2898 1771 2899 1772
rect 2903 1771 2904 1775
rect 2898 1770 2904 1771
rect 3051 1775 3057 1776
rect 3051 1771 3052 1775
rect 3056 1774 3057 1775
rect 3082 1775 3088 1776
rect 3082 1774 3083 1775
rect 3056 1772 3083 1774
rect 3056 1771 3057 1772
rect 3051 1770 3057 1771
rect 3082 1771 3083 1772
rect 3087 1771 3088 1775
rect 3082 1770 3088 1771
rect 3235 1775 3241 1776
rect 3235 1771 3236 1775
rect 3240 1774 3241 1775
rect 3258 1775 3264 1776
rect 3258 1774 3259 1775
rect 3240 1772 3259 1774
rect 3240 1771 3241 1772
rect 3235 1770 3241 1771
rect 3258 1771 3259 1772
rect 3263 1771 3264 1775
rect 3258 1770 3264 1771
rect 3335 1775 3341 1776
rect 3335 1771 3336 1775
rect 3340 1774 3341 1775
rect 3427 1775 3433 1776
rect 3427 1774 3428 1775
rect 3340 1772 3428 1774
rect 3340 1771 3341 1772
rect 3335 1770 3341 1771
rect 3427 1771 3428 1772
rect 3432 1771 3433 1775
rect 3427 1770 3433 1771
rect 282 1767 289 1768
rect 282 1763 283 1767
rect 288 1763 289 1767
rect 282 1762 289 1763
rect 407 1767 413 1768
rect 407 1763 408 1767
rect 412 1766 413 1767
rect 451 1767 457 1768
rect 451 1766 452 1767
rect 412 1764 452 1766
rect 412 1763 413 1764
rect 407 1762 413 1763
rect 451 1763 452 1764
rect 456 1763 457 1767
rect 451 1762 457 1763
rect 574 1767 580 1768
rect 574 1763 575 1767
rect 579 1766 580 1767
rect 627 1767 633 1768
rect 627 1766 628 1767
rect 579 1764 628 1766
rect 579 1763 580 1764
rect 574 1762 580 1763
rect 627 1763 628 1764
rect 632 1763 633 1767
rect 627 1762 633 1763
rect 795 1767 801 1768
rect 795 1763 796 1767
rect 800 1766 801 1767
rect 826 1767 832 1768
rect 826 1766 827 1767
rect 800 1764 827 1766
rect 800 1763 801 1764
rect 795 1762 801 1763
rect 826 1763 827 1764
rect 831 1763 832 1767
rect 826 1762 832 1763
rect 963 1767 969 1768
rect 963 1763 964 1767
rect 968 1766 969 1767
rect 978 1767 984 1768
rect 978 1766 979 1767
rect 968 1764 979 1766
rect 968 1763 969 1764
rect 963 1762 969 1763
rect 978 1763 979 1764
rect 983 1763 984 1767
rect 978 1762 984 1763
rect 1115 1767 1121 1768
rect 1115 1763 1116 1767
rect 1120 1766 1121 1767
rect 1146 1767 1152 1768
rect 1146 1766 1147 1767
rect 1120 1764 1147 1766
rect 1120 1763 1121 1764
rect 1115 1762 1121 1763
rect 1146 1763 1147 1764
rect 1151 1763 1152 1767
rect 1146 1762 1152 1763
rect 1259 1767 1265 1768
rect 1259 1763 1260 1767
rect 1264 1766 1265 1767
rect 1290 1767 1296 1768
rect 1290 1766 1291 1767
rect 1264 1764 1291 1766
rect 1264 1763 1265 1764
rect 1259 1762 1265 1763
rect 1290 1763 1291 1764
rect 1295 1763 1296 1767
rect 1290 1762 1296 1763
rect 1395 1767 1401 1768
rect 1395 1763 1396 1767
rect 1400 1766 1401 1767
rect 1434 1767 1440 1768
rect 1434 1766 1435 1767
rect 1400 1764 1435 1766
rect 1400 1763 1401 1764
rect 1395 1762 1401 1763
rect 1434 1763 1435 1764
rect 1439 1763 1440 1767
rect 1434 1762 1440 1763
rect 1523 1767 1529 1768
rect 1523 1763 1524 1767
rect 1528 1766 1529 1767
rect 1554 1767 1560 1768
rect 1554 1766 1555 1767
rect 1528 1764 1555 1766
rect 1528 1763 1529 1764
rect 1523 1762 1529 1763
rect 1554 1763 1555 1764
rect 1559 1763 1560 1767
rect 1554 1762 1560 1763
rect 1651 1767 1657 1768
rect 1651 1763 1652 1767
rect 1656 1766 1657 1767
rect 1682 1767 1688 1768
rect 1682 1766 1683 1767
rect 1656 1764 1683 1766
rect 1656 1763 1657 1764
rect 1651 1762 1657 1763
rect 1682 1763 1683 1764
rect 1687 1763 1688 1767
rect 1682 1762 1688 1763
rect 1763 1767 1772 1768
rect 1763 1763 1764 1767
rect 1771 1763 1772 1767
rect 1763 1762 1772 1763
rect 538 1759 544 1760
rect 538 1758 539 1759
rect 356 1756 539 1758
rect 356 1754 358 1756
rect 538 1755 539 1756
rect 543 1755 544 1759
rect 1971 1759 1977 1760
rect 538 1754 544 1755
rect 1562 1755 1568 1756
rect 1562 1754 1563 1755
rect 355 1753 361 1754
rect 355 1749 356 1753
rect 360 1749 361 1753
rect 1555 1753 1563 1754
rect 355 1748 361 1749
rect 415 1751 421 1752
rect 415 1747 416 1751
rect 420 1750 421 1751
rect 499 1751 505 1752
rect 499 1750 500 1751
rect 420 1748 500 1750
rect 420 1747 421 1748
rect 415 1746 421 1747
rect 499 1747 500 1748
rect 504 1747 505 1751
rect 499 1746 505 1747
rect 643 1751 649 1752
rect 643 1747 644 1751
rect 648 1750 649 1751
rect 658 1751 664 1752
rect 658 1750 659 1751
rect 648 1748 659 1750
rect 648 1747 649 1748
rect 643 1746 649 1747
rect 658 1747 659 1748
rect 663 1747 664 1751
rect 658 1746 664 1747
rect 795 1751 801 1752
rect 795 1747 796 1751
rect 800 1750 801 1751
rect 838 1751 844 1752
rect 838 1750 839 1751
rect 800 1748 839 1750
rect 800 1747 801 1748
rect 795 1746 801 1747
rect 838 1747 839 1748
rect 843 1747 844 1751
rect 838 1746 844 1747
rect 863 1751 869 1752
rect 863 1747 864 1751
rect 868 1750 869 1751
rect 947 1751 953 1752
rect 947 1750 948 1751
rect 868 1748 948 1750
rect 868 1747 869 1748
rect 863 1746 869 1747
rect 947 1747 948 1748
rect 952 1747 953 1751
rect 947 1746 953 1747
rect 1099 1751 1105 1752
rect 1099 1747 1100 1751
rect 1104 1750 1105 1751
rect 1110 1751 1116 1752
rect 1110 1750 1111 1751
rect 1104 1748 1111 1750
rect 1104 1747 1105 1748
rect 1099 1746 1105 1747
rect 1110 1747 1111 1748
rect 1115 1747 1116 1751
rect 1110 1746 1116 1747
rect 1207 1751 1213 1752
rect 1207 1747 1208 1751
rect 1212 1750 1213 1751
rect 1251 1751 1257 1752
rect 1251 1750 1252 1751
rect 1212 1748 1252 1750
rect 1212 1747 1213 1748
rect 1207 1746 1213 1747
rect 1251 1747 1252 1748
rect 1256 1747 1257 1751
rect 1251 1746 1257 1747
rect 1319 1751 1325 1752
rect 1319 1747 1320 1751
rect 1324 1750 1325 1751
rect 1403 1751 1409 1752
rect 1403 1750 1404 1751
rect 1324 1748 1404 1750
rect 1324 1747 1325 1748
rect 1319 1746 1325 1747
rect 1403 1747 1404 1748
rect 1408 1747 1409 1751
rect 1555 1749 1556 1753
rect 1560 1751 1563 1753
rect 1567 1751 1568 1755
rect 1971 1755 1972 1759
rect 1976 1758 1977 1759
rect 2034 1759 2040 1760
rect 2034 1758 2035 1759
rect 1976 1756 2035 1758
rect 1976 1755 1977 1756
rect 1971 1754 1977 1755
rect 2034 1755 2035 1756
rect 2039 1755 2040 1759
rect 2034 1754 2040 1755
rect 2115 1759 2121 1760
rect 2115 1755 2116 1759
rect 2120 1758 2121 1759
rect 2186 1759 2192 1760
rect 2186 1758 2187 1759
rect 2120 1756 2187 1758
rect 2120 1755 2121 1756
rect 2115 1754 2121 1755
rect 2186 1755 2187 1756
rect 2191 1755 2192 1759
rect 2186 1754 2192 1755
rect 2223 1759 2229 1760
rect 2223 1755 2224 1759
rect 2228 1758 2229 1759
rect 2275 1759 2281 1760
rect 2275 1758 2276 1759
rect 2228 1756 2276 1758
rect 2228 1755 2229 1756
rect 2223 1754 2229 1755
rect 2275 1755 2276 1756
rect 2280 1755 2281 1759
rect 2275 1754 2281 1755
rect 2431 1759 2437 1760
rect 2431 1755 2432 1759
rect 2436 1758 2437 1759
rect 2443 1759 2449 1760
rect 2443 1758 2444 1759
rect 2436 1756 2444 1758
rect 2436 1755 2437 1756
rect 2431 1754 2437 1755
rect 2443 1755 2444 1756
rect 2448 1755 2449 1759
rect 2443 1754 2449 1755
rect 2527 1759 2533 1760
rect 2527 1755 2528 1759
rect 2532 1758 2533 1759
rect 2627 1759 2633 1760
rect 2627 1758 2628 1759
rect 2532 1756 2628 1758
rect 2532 1755 2533 1756
rect 2527 1754 2533 1755
rect 2627 1755 2628 1756
rect 2632 1755 2633 1759
rect 2627 1754 2633 1755
rect 2818 1759 2825 1760
rect 2818 1755 2819 1759
rect 2824 1755 2825 1759
rect 2818 1754 2825 1755
rect 2911 1759 2917 1760
rect 2911 1755 2912 1759
rect 2916 1758 2917 1759
rect 3019 1759 3025 1760
rect 3019 1758 3020 1759
rect 2916 1756 3020 1758
rect 2916 1755 2917 1756
rect 2911 1754 2917 1755
rect 3019 1755 3020 1756
rect 3024 1755 3025 1759
rect 3019 1754 3025 1755
rect 3227 1759 3236 1760
rect 3227 1755 3228 1759
rect 3235 1755 3236 1759
rect 3227 1754 3236 1755
rect 3443 1759 3449 1760
rect 3443 1755 3444 1759
rect 3448 1758 3449 1759
rect 3458 1759 3464 1760
rect 3458 1758 3459 1759
rect 3448 1756 3459 1758
rect 3448 1755 3449 1756
rect 3443 1754 3449 1755
rect 3458 1755 3459 1756
rect 3463 1755 3464 1759
rect 3458 1754 3464 1755
rect 1560 1750 1568 1751
rect 1623 1751 1629 1752
rect 1560 1749 1561 1750
rect 1555 1748 1561 1749
rect 1403 1746 1409 1747
rect 1623 1747 1624 1751
rect 1628 1750 1629 1751
rect 1715 1751 1721 1752
rect 1715 1750 1716 1751
rect 1628 1748 1716 1750
rect 1628 1747 1629 1748
rect 1623 1746 1629 1747
rect 1715 1747 1716 1748
rect 1720 1747 1721 1751
rect 1715 1746 1721 1747
rect 1942 1749 1948 1750
rect 1942 1745 1943 1749
rect 1947 1745 1948 1749
rect 1942 1744 1948 1745
rect 2086 1749 2092 1750
rect 2086 1745 2087 1749
rect 2091 1745 2092 1749
rect 2086 1744 2092 1745
rect 2246 1749 2252 1750
rect 2246 1745 2247 1749
rect 2251 1745 2252 1749
rect 2246 1744 2252 1745
rect 2414 1749 2420 1750
rect 2414 1745 2415 1749
rect 2419 1745 2420 1749
rect 2414 1744 2420 1745
rect 2598 1749 2604 1750
rect 2598 1745 2599 1749
rect 2603 1745 2604 1749
rect 2598 1744 2604 1745
rect 2790 1749 2796 1750
rect 2790 1745 2791 1749
rect 2795 1745 2796 1749
rect 2790 1744 2796 1745
rect 2990 1749 2996 1750
rect 2990 1745 2991 1749
rect 2995 1745 2996 1749
rect 2990 1744 2996 1745
rect 3198 1749 3204 1750
rect 3198 1745 3199 1749
rect 3203 1745 3204 1749
rect 3198 1744 3204 1745
rect 3414 1749 3420 1750
rect 3414 1745 3415 1749
rect 3419 1745 3420 1749
rect 3414 1744 3420 1745
rect 326 1741 332 1742
rect 326 1737 327 1741
rect 331 1737 332 1741
rect 326 1736 332 1737
rect 470 1741 476 1742
rect 470 1737 471 1741
rect 475 1737 476 1741
rect 470 1736 476 1737
rect 614 1741 620 1742
rect 614 1737 615 1741
rect 619 1737 620 1741
rect 614 1736 620 1737
rect 766 1741 772 1742
rect 766 1737 767 1741
rect 771 1737 772 1741
rect 766 1736 772 1737
rect 918 1741 924 1742
rect 918 1737 919 1741
rect 923 1737 924 1741
rect 918 1736 924 1737
rect 1070 1741 1076 1742
rect 1070 1737 1071 1741
rect 1075 1737 1076 1741
rect 1070 1736 1076 1737
rect 1222 1741 1228 1742
rect 1222 1737 1223 1741
rect 1227 1737 1228 1741
rect 1222 1736 1228 1737
rect 1374 1741 1380 1742
rect 1374 1737 1375 1741
rect 1379 1737 1380 1741
rect 1374 1736 1380 1737
rect 1526 1741 1532 1742
rect 1526 1737 1527 1741
rect 1531 1737 1532 1741
rect 1526 1736 1532 1737
rect 1686 1741 1692 1742
rect 1686 1737 1687 1741
rect 1691 1737 1692 1741
rect 1686 1736 1692 1737
rect 1862 1736 1868 1737
rect 3574 1736 3580 1737
rect 1862 1732 1863 1736
rect 1867 1732 1868 1736
rect 2007 1735 2013 1736
rect 2007 1734 2008 1735
rect 1997 1732 2008 1734
rect 1862 1731 1868 1732
rect 2007 1731 2008 1732
rect 2012 1731 2013 1735
rect 2527 1735 2533 1736
rect 2527 1734 2528 1735
rect 2469 1732 2528 1734
rect 2007 1730 2013 1731
rect 2034 1731 2040 1732
rect 110 1728 116 1729
rect 1822 1728 1828 1729
rect 110 1724 111 1728
rect 115 1724 116 1728
rect 415 1727 421 1728
rect 415 1726 416 1727
rect 381 1724 416 1726
rect 110 1723 116 1724
rect 415 1723 416 1724
rect 420 1723 421 1727
rect 863 1727 869 1728
rect 863 1726 864 1727
rect 821 1724 864 1726
rect 415 1722 421 1723
rect 538 1723 544 1724
rect 538 1719 539 1723
rect 543 1722 544 1723
rect 863 1723 864 1724
rect 868 1723 869 1727
rect 978 1727 984 1728
rect 978 1726 979 1727
rect 973 1724 979 1726
rect 863 1722 869 1723
rect 978 1723 979 1724
rect 983 1723 984 1727
rect 1207 1727 1213 1728
rect 1207 1726 1208 1727
rect 1125 1724 1208 1726
rect 978 1722 984 1723
rect 1207 1723 1208 1724
rect 1212 1723 1213 1727
rect 1319 1727 1325 1728
rect 1319 1726 1320 1727
rect 1277 1724 1320 1726
rect 1207 1722 1213 1723
rect 1319 1723 1320 1724
rect 1324 1723 1325 1727
rect 1434 1727 1440 1728
rect 1434 1726 1435 1727
rect 1429 1724 1435 1726
rect 1319 1722 1325 1723
rect 1434 1723 1435 1724
rect 1439 1723 1440 1727
rect 1623 1727 1629 1728
rect 1623 1726 1624 1727
rect 1581 1724 1624 1726
rect 1434 1722 1440 1723
rect 1623 1723 1624 1724
rect 1628 1723 1629 1727
rect 1822 1724 1823 1728
rect 1827 1724 1828 1728
rect 2034 1727 2035 1731
rect 2039 1730 2040 1731
rect 2186 1731 2192 1732
rect 2039 1728 2105 1730
rect 2039 1727 2040 1728
rect 2034 1726 2040 1727
rect 2186 1727 2187 1731
rect 2191 1730 2192 1731
rect 2527 1731 2528 1732
rect 2532 1731 2533 1735
rect 2911 1735 2917 1736
rect 2911 1734 2912 1735
rect 2845 1732 2912 1734
rect 2527 1730 2533 1731
rect 2911 1731 2912 1732
rect 2916 1731 2917 1735
rect 3258 1735 3264 1736
rect 3258 1734 3259 1735
rect 3253 1732 3259 1734
rect 2911 1730 2917 1731
rect 3258 1731 3259 1732
rect 3263 1731 3264 1735
rect 3574 1732 3575 1736
rect 3579 1732 3580 1736
rect 3574 1731 3580 1732
rect 3258 1730 3264 1731
rect 2191 1728 2265 1730
rect 2191 1727 2192 1728
rect 2186 1726 2192 1727
rect 1822 1723 1828 1724
rect 1623 1722 1629 1723
rect 543 1720 633 1722
rect 543 1719 544 1720
rect 538 1718 544 1719
rect 1862 1719 1868 1720
rect 1862 1715 1863 1719
rect 1867 1715 1868 1719
rect 3082 1719 3088 1720
rect 3082 1718 3083 1719
rect 1862 1714 1868 1715
rect 2476 1716 2609 1718
rect 3041 1716 3083 1718
rect 110 1711 116 1712
rect 110 1707 111 1711
rect 115 1707 116 1711
rect 614 1711 620 1712
rect 614 1710 615 1711
rect 521 1708 615 1710
rect 110 1706 116 1707
rect 614 1707 615 1708
rect 619 1707 620 1711
rect 614 1706 620 1707
rect 1686 1711 1692 1712
rect 1686 1707 1687 1711
rect 1691 1710 1692 1711
rect 1822 1711 1828 1712
rect 1691 1708 1697 1710
rect 1691 1707 1692 1708
rect 1686 1706 1692 1707
rect 1822 1707 1823 1711
rect 1827 1707 1828 1711
rect 1822 1706 1828 1707
rect 1934 1709 1940 1710
rect 1934 1705 1935 1709
rect 1939 1705 1940 1709
rect 1934 1704 1940 1705
rect 2078 1709 2084 1710
rect 2078 1705 2079 1709
rect 2083 1705 2084 1709
rect 2078 1704 2084 1705
rect 2238 1709 2244 1710
rect 2238 1705 2239 1709
rect 2243 1705 2244 1709
rect 2238 1704 2244 1705
rect 2406 1709 2412 1710
rect 2406 1705 2407 1709
rect 2411 1705 2412 1709
rect 2406 1704 2412 1705
rect 2310 1703 2316 1704
rect 318 1701 324 1702
rect 318 1697 319 1701
rect 323 1697 324 1701
rect 318 1696 324 1697
rect 462 1701 468 1702
rect 462 1697 463 1701
rect 467 1697 468 1701
rect 462 1696 468 1697
rect 606 1701 612 1702
rect 606 1697 607 1701
rect 611 1697 612 1701
rect 606 1696 612 1697
rect 758 1701 764 1702
rect 758 1697 759 1701
rect 763 1697 764 1701
rect 758 1696 764 1697
rect 910 1701 916 1702
rect 910 1697 911 1701
rect 915 1697 916 1701
rect 910 1696 916 1697
rect 1062 1701 1068 1702
rect 1062 1697 1063 1701
rect 1067 1697 1068 1701
rect 1062 1696 1068 1697
rect 1214 1701 1220 1702
rect 1214 1697 1215 1701
rect 1219 1697 1220 1701
rect 1214 1696 1220 1697
rect 1366 1701 1372 1702
rect 1366 1697 1367 1701
rect 1371 1697 1372 1701
rect 1366 1696 1372 1697
rect 1518 1701 1524 1702
rect 1518 1697 1519 1701
rect 1523 1697 1524 1701
rect 1518 1696 1524 1697
rect 1678 1701 1684 1702
rect 1678 1697 1679 1701
rect 1683 1697 1684 1701
rect 2310 1699 2311 1703
rect 2315 1702 2316 1703
rect 2476 1702 2478 1716
rect 3082 1715 3083 1716
rect 3087 1715 3088 1719
rect 3082 1714 3088 1715
rect 3574 1719 3580 1720
rect 3574 1715 3575 1719
rect 3579 1715 3580 1719
rect 3574 1714 3580 1715
rect 2590 1709 2596 1710
rect 2590 1705 2591 1709
rect 2595 1705 2596 1709
rect 2590 1704 2596 1705
rect 2782 1709 2788 1710
rect 2782 1705 2783 1709
rect 2787 1705 2788 1709
rect 2782 1704 2788 1705
rect 2982 1709 2988 1710
rect 2982 1705 2983 1709
rect 2987 1705 2988 1709
rect 2982 1704 2988 1705
rect 3190 1709 3196 1710
rect 3190 1705 3191 1709
rect 3195 1705 3196 1709
rect 3190 1704 3196 1705
rect 3406 1709 3412 1710
rect 3406 1705 3407 1709
rect 3411 1705 3412 1709
rect 3406 1704 3412 1705
rect 2315 1700 2478 1702
rect 3455 1703 3461 1704
rect 2315 1699 2316 1700
rect 2310 1698 2316 1699
rect 3455 1699 3456 1703
rect 3460 1702 3461 1703
rect 3466 1703 3472 1704
rect 3466 1702 3467 1703
rect 3460 1700 3467 1702
rect 3460 1699 3461 1700
rect 3455 1698 3461 1699
rect 3466 1699 3467 1700
rect 3471 1699 3472 1703
rect 3466 1698 3472 1699
rect 1678 1696 1684 1697
rect 1910 1683 1916 1684
rect 1910 1679 1911 1683
rect 1915 1679 1916 1683
rect 1910 1678 1916 1679
rect 2030 1683 2036 1684
rect 2030 1679 2031 1683
rect 2035 1679 2036 1683
rect 2030 1678 2036 1679
rect 2150 1683 2156 1684
rect 2150 1679 2151 1683
rect 2155 1679 2156 1683
rect 2150 1678 2156 1679
rect 2270 1683 2276 1684
rect 2270 1679 2271 1683
rect 2275 1679 2276 1683
rect 2270 1678 2276 1679
rect 2398 1683 2404 1684
rect 2398 1679 2399 1683
rect 2403 1679 2404 1683
rect 2398 1678 2404 1679
rect 2542 1683 2548 1684
rect 2542 1679 2543 1683
rect 2547 1679 2548 1683
rect 2542 1678 2548 1679
rect 2694 1683 2700 1684
rect 2694 1679 2695 1683
rect 2699 1679 2700 1683
rect 2694 1678 2700 1679
rect 2862 1683 2868 1684
rect 2862 1679 2863 1683
rect 2867 1679 2868 1683
rect 2862 1678 2868 1679
rect 3046 1683 3052 1684
rect 3046 1679 3047 1683
rect 3051 1679 3052 1683
rect 3046 1678 3052 1679
rect 3238 1683 3244 1684
rect 3238 1679 3239 1683
rect 3243 1679 3244 1683
rect 3238 1678 3244 1679
rect 3430 1683 3436 1684
rect 3430 1679 3431 1683
rect 3435 1679 3436 1683
rect 3430 1678 3436 1679
rect 310 1675 316 1676
rect 310 1671 311 1675
rect 315 1671 316 1675
rect 310 1670 316 1671
rect 446 1675 452 1676
rect 446 1671 447 1675
rect 451 1671 452 1675
rect 446 1670 452 1671
rect 590 1675 596 1676
rect 590 1671 591 1675
rect 595 1671 596 1675
rect 590 1670 596 1671
rect 734 1675 740 1676
rect 734 1671 735 1675
rect 739 1671 740 1675
rect 734 1670 740 1671
rect 886 1675 892 1676
rect 886 1671 887 1675
rect 891 1671 892 1675
rect 886 1670 892 1671
rect 1038 1675 1044 1676
rect 1038 1671 1039 1675
rect 1043 1671 1044 1675
rect 1038 1670 1044 1671
rect 1190 1675 1196 1676
rect 1190 1671 1191 1675
rect 1195 1671 1196 1675
rect 1190 1670 1196 1671
rect 1342 1675 1348 1676
rect 1342 1671 1343 1675
rect 1347 1671 1348 1675
rect 1342 1670 1348 1671
rect 1494 1675 1500 1676
rect 1494 1671 1495 1675
rect 1499 1671 1500 1675
rect 1494 1670 1500 1671
rect 1646 1675 1652 1676
rect 1646 1671 1647 1675
rect 1651 1671 1652 1675
rect 2223 1675 2229 1676
rect 2223 1674 2224 1675
rect 1646 1670 1652 1671
rect 1862 1673 1868 1674
rect 1862 1669 1863 1673
rect 1867 1669 1868 1673
rect 2209 1672 2224 1674
rect 2223 1671 2224 1672
rect 2228 1671 2229 1675
rect 2223 1670 2229 1671
rect 3230 1675 3236 1676
rect 3230 1671 3231 1675
rect 3235 1674 3236 1675
rect 3235 1672 3257 1674
rect 3574 1673 3580 1674
rect 3235 1671 3236 1672
rect 3230 1670 3236 1671
rect 1862 1668 1868 1669
rect 3574 1669 3575 1673
rect 3579 1669 3580 1673
rect 3574 1668 3580 1669
rect 838 1667 844 1668
rect 110 1665 116 1666
rect 110 1661 111 1665
rect 115 1661 116 1665
rect 838 1663 839 1667
rect 843 1666 844 1667
rect 1110 1667 1116 1668
rect 1110 1666 1111 1667
rect 843 1664 905 1666
rect 1097 1664 1111 1666
rect 843 1663 844 1664
rect 838 1662 844 1663
rect 1110 1663 1111 1664
rect 1115 1663 1116 1667
rect 1110 1662 1116 1663
rect 1822 1665 1828 1666
rect 110 1660 116 1661
rect 1822 1661 1823 1665
rect 1827 1661 1828 1665
rect 1822 1660 1828 1661
rect 2023 1659 2029 1660
rect 2023 1658 2024 1659
rect 1862 1656 1868 1657
rect 1973 1656 2024 1658
rect 1862 1652 1863 1656
rect 1867 1652 1868 1656
rect 2023 1655 2024 1656
rect 2028 1655 2029 1659
rect 2143 1659 2149 1660
rect 2143 1658 2144 1659
rect 2093 1656 2144 1658
rect 2023 1654 2029 1655
rect 2143 1655 2144 1656
rect 2148 1655 2149 1659
rect 2391 1659 2397 1660
rect 2391 1658 2392 1659
rect 2333 1656 2392 1658
rect 2143 1654 2149 1655
rect 2391 1655 2392 1656
rect 2396 1655 2397 1659
rect 2466 1659 2472 1660
rect 2466 1658 2467 1659
rect 2461 1656 2467 1658
rect 2391 1654 2397 1655
rect 2466 1655 2467 1656
rect 2471 1655 2472 1659
rect 2610 1659 2616 1660
rect 2466 1654 2472 1655
rect 254 1651 260 1652
rect 110 1648 116 1649
rect 110 1644 111 1648
rect 115 1644 116 1648
rect 254 1647 255 1651
rect 259 1650 260 1651
rect 378 1651 384 1652
rect 259 1648 337 1650
rect 259 1647 260 1648
rect 254 1646 260 1647
rect 378 1647 379 1651
rect 383 1650 384 1651
rect 514 1651 520 1652
rect 383 1648 473 1650
rect 383 1647 384 1648
rect 378 1646 384 1647
rect 514 1647 515 1651
rect 519 1650 520 1651
rect 879 1651 885 1652
rect 879 1650 880 1651
rect 519 1648 617 1650
rect 797 1648 880 1650
rect 519 1647 520 1648
rect 514 1646 520 1647
rect 879 1647 880 1648
rect 884 1647 885 1651
rect 879 1646 885 1647
rect 1142 1651 1148 1652
rect 1142 1647 1143 1651
rect 1147 1650 1148 1651
rect 1410 1651 1416 1652
rect 1147 1648 1217 1650
rect 1147 1647 1148 1648
rect 1142 1646 1148 1647
rect 110 1643 116 1644
rect 1404 1642 1406 1649
rect 1410 1647 1411 1651
rect 1415 1650 1416 1651
rect 1562 1651 1568 1652
rect 1862 1651 1868 1652
rect 1415 1648 1521 1650
rect 1415 1647 1416 1648
rect 1410 1646 1416 1647
rect 1562 1647 1563 1651
rect 1567 1650 1568 1651
rect 2604 1650 2606 1657
rect 2610 1655 2611 1659
rect 2615 1658 2616 1659
rect 2762 1659 2768 1660
rect 2615 1656 2721 1658
rect 2615 1655 2616 1656
rect 2610 1654 2616 1655
rect 2762 1655 2763 1659
rect 2767 1658 2768 1659
rect 2930 1659 2936 1660
rect 2767 1656 2889 1658
rect 2767 1655 2768 1656
rect 2762 1654 2768 1655
rect 2930 1655 2931 1659
rect 2935 1658 2936 1659
rect 3498 1659 3504 1660
rect 3498 1658 3499 1659
rect 2935 1656 3073 1658
rect 3493 1656 3499 1658
rect 2935 1655 2936 1656
rect 2930 1654 2936 1655
rect 3498 1655 3499 1656
rect 3503 1655 3504 1659
rect 3498 1654 3504 1655
rect 3574 1656 3580 1657
rect 3574 1652 3575 1656
rect 3579 1652 3580 1656
rect 2618 1651 2624 1652
rect 3574 1651 3580 1652
rect 2618 1650 2619 1651
rect 1567 1648 1673 1650
rect 1822 1648 1828 1649
rect 2604 1648 2619 1650
rect 1567 1647 1568 1648
rect 1562 1646 1568 1647
rect 1822 1644 1823 1648
rect 1827 1644 1828 1648
rect 2618 1647 2619 1648
rect 2623 1647 2624 1651
rect 2618 1646 2624 1647
rect 1415 1643 1421 1644
rect 1822 1643 1828 1644
rect 1918 1643 1924 1644
rect 1415 1642 1416 1643
rect 1404 1640 1416 1642
rect 1415 1639 1416 1640
rect 1420 1639 1421 1643
rect 1415 1638 1421 1639
rect 1918 1639 1919 1643
rect 1923 1639 1924 1643
rect 1918 1638 1924 1639
rect 2038 1643 2044 1644
rect 2038 1639 2039 1643
rect 2043 1639 2044 1643
rect 2038 1638 2044 1639
rect 2158 1643 2164 1644
rect 2158 1639 2159 1643
rect 2163 1639 2164 1643
rect 2158 1638 2164 1639
rect 2278 1643 2284 1644
rect 2278 1639 2279 1643
rect 2283 1639 2284 1643
rect 2278 1638 2284 1639
rect 2406 1643 2412 1644
rect 2406 1639 2407 1643
rect 2411 1639 2412 1643
rect 2406 1638 2412 1639
rect 2550 1643 2556 1644
rect 2550 1639 2551 1643
rect 2555 1639 2556 1643
rect 2550 1638 2556 1639
rect 2702 1643 2708 1644
rect 2702 1639 2703 1643
rect 2707 1639 2708 1643
rect 2702 1638 2708 1639
rect 2870 1643 2876 1644
rect 2870 1639 2871 1643
rect 2875 1639 2876 1643
rect 2870 1638 2876 1639
rect 3054 1643 3060 1644
rect 3054 1639 3055 1643
rect 3059 1639 3060 1643
rect 3054 1638 3060 1639
rect 3246 1643 3252 1644
rect 3246 1639 3247 1643
rect 3251 1639 3252 1643
rect 3246 1638 3252 1639
rect 3438 1643 3444 1644
rect 3438 1639 3439 1643
rect 3443 1639 3444 1643
rect 3438 1638 3444 1639
rect 318 1635 324 1636
rect 318 1631 319 1635
rect 323 1631 324 1635
rect 318 1630 324 1631
rect 454 1635 460 1636
rect 454 1631 455 1635
rect 459 1631 460 1635
rect 454 1630 460 1631
rect 598 1635 604 1636
rect 598 1631 599 1635
rect 603 1631 604 1635
rect 598 1630 604 1631
rect 742 1635 748 1636
rect 742 1631 743 1635
rect 747 1631 748 1635
rect 742 1630 748 1631
rect 894 1635 900 1636
rect 894 1631 895 1635
rect 899 1631 900 1635
rect 894 1630 900 1631
rect 1046 1635 1052 1636
rect 1046 1631 1047 1635
rect 1051 1631 1052 1635
rect 1046 1630 1052 1631
rect 1198 1635 1204 1636
rect 1198 1631 1199 1635
rect 1203 1631 1204 1635
rect 1198 1630 1204 1631
rect 1350 1635 1356 1636
rect 1350 1631 1351 1635
rect 1355 1631 1356 1635
rect 1350 1630 1356 1631
rect 1502 1635 1508 1636
rect 1502 1631 1503 1635
rect 1507 1631 1508 1635
rect 1502 1630 1508 1631
rect 1654 1635 1660 1636
rect 1654 1631 1655 1635
rect 1659 1631 1660 1635
rect 1654 1630 1660 1631
rect 1947 1631 1953 1632
rect 1947 1627 1948 1631
rect 1952 1630 1953 1631
rect 1958 1631 1964 1632
rect 1958 1630 1959 1631
rect 1952 1628 1959 1630
rect 1952 1627 1953 1628
rect 1947 1626 1953 1627
rect 1958 1627 1959 1628
rect 1963 1627 1964 1631
rect 1958 1626 1964 1627
rect 2023 1631 2029 1632
rect 2023 1627 2024 1631
rect 2028 1630 2029 1631
rect 2067 1631 2073 1632
rect 2067 1630 2068 1631
rect 2028 1628 2068 1630
rect 2028 1627 2029 1628
rect 2023 1626 2029 1627
rect 2067 1627 2068 1628
rect 2072 1627 2073 1631
rect 2067 1626 2073 1627
rect 2143 1631 2149 1632
rect 2143 1627 2144 1631
rect 2148 1630 2149 1631
rect 2187 1631 2193 1632
rect 2187 1630 2188 1631
rect 2148 1628 2188 1630
rect 2148 1627 2149 1628
rect 2143 1626 2149 1627
rect 2187 1627 2188 1628
rect 2192 1627 2193 1631
rect 2187 1626 2193 1627
rect 2307 1631 2316 1632
rect 2307 1627 2308 1631
rect 2315 1627 2316 1631
rect 2307 1626 2316 1627
rect 2391 1631 2397 1632
rect 2391 1627 2392 1631
rect 2396 1630 2397 1631
rect 2435 1631 2441 1632
rect 2435 1630 2436 1631
rect 2396 1628 2436 1630
rect 2396 1627 2397 1628
rect 2391 1626 2397 1627
rect 2435 1627 2436 1628
rect 2440 1627 2441 1631
rect 2435 1626 2441 1627
rect 2579 1631 2585 1632
rect 2579 1627 2580 1631
rect 2584 1630 2585 1631
rect 2610 1631 2616 1632
rect 2610 1630 2611 1631
rect 2584 1628 2611 1630
rect 2584 1627 2585 1628
rect 2579 1626 2585 1627
rect 2610 1627 2611 1628
rect 2615 1627 2616 1631
rect 2610 1626 2616 1627
rect 2731 1631 2737 1632
rect 2731 1627 2732 1631
rect 2736 1630 2737 1631
rect 2762 1631 2768 1632
rect 2762 1630 2763 1631
rect 2736 1628 2763 1630
rect 2736 1627 2737 1628
rect 2731 1626 2737 1627
rect 2762 1627 2763 1628
rect 2767 1627 2768 1631
rect 2762 1626 2768 1627
rect 2899 1631 2905 1632
rect 2899 1627 2900 1631
rect 2904 1630 2905 1631
rect 2930 1631 2936 1632
rect 2930 1630 2931 1631
rect 2904 1628 2931 1630
rect 2904 1627 2905 1628
rect 2899 1626 2905 1627
rect 2930 1627 2931 1628
rect 2935 1627 2936 1631
rect 2930 1626 2936 1627
rect 3082 1631 3089 1632
rect 3082 1627 3083 1631
rect 3088 1627 3089 1631
rect 3082 1626 3089 1627
rect 3270 1631 3281 1632
rect 3270 1627 3271 1631
rect 3275 1627 3276 1631
rect 3280 1627 3281 1631
rect 3270 1626 3281 1627
rect 3466 1631 3473 1632
rect 3466 1627 3467 1631
rect 3472 1627 3473 1631
rect 3466 1626 3473 1627
rect 347 1623 353 1624
rect 347 1619 348 1623
rect 352 1622 353 1623
rect 378 1623 384 1624
rect 378 1622 379 1623
rect 352 1620 379 1622
rect 352 1619 353 1620
rect 347 1618 353 1619
rect 378 1619 379 1620
rect 383 1619 384 1623
rect 378 1618 384 1619
rect 483 1623 489 1624
rect 483 1619 484 1623
rect 488 1622 489 1623
rect 514 1623 520 1624
rect 514 1622 515 1623
rect 488 1620 515 1622
rect 488 1619 489 1620
rect 483 1618 489 1619
rect 514 1619 515 1620
rect 519 1619 520 1623
rect 514 1618 520 1619
rect 614 1623 620 1624
rect 614 1619 615 1623
rect 619 1622 620 1623
rect 627 1623 633 1624
rect 627 1622 628 1623
rect 619 1620 628 1622
rect 619 1619 620 1620
rect 614 1618 620 1619
rect 627 1619 628 1620
rect 632 1619 633 1623
rect 627 1618 633 1619
rect 750 1623 756 1624
rect 750 1619 751 1623
rect 755 1622 756 1623
rect 771 1623 777 1624
rect 771 1622 772 1623
rect 755 1620 772 1622
rect 755 1619 756 1620
rect 750 1618 756 1619
rect 771 1619 772 1620
rect 776 1619 777 1623
rect 771 1618 777 1619
rect 879 1623 885 1624
rect 879 1619 880 1623
rect 884 1622 885 1623
rect 923 1623 929 1624
rect 923 1622 924 1623
rect 884 1620 924 1622
rect 884 1619 885 1620
rect 879 1618 885 1619
rect 923 1619 924 1620
rect 928 1619 929 1623
rect 923 1618 929 1619
rect 1075 1623 1081 1624
rect 1075 1619 1076 1623
rect 1080 1622 1081 1623
rect 1142 1623 1148 1624
rect 1142 1622 1143 1623
rect 1080 1620 1143 1622
rect 1080 1619 1081 1620
rect 1075 1618 1081 1619
rect 1142 1619 1143 1620
rect 1147 1619 1148 1623
rect 1142 1618 1148 1619
rect 1206 1623 1212 1624
rect 1206 1619 1207 1623
rect 1211 1622 1212 1623
rect 1227 1623 1233 1624
rect 1227 1622 1228 1623
rect 1211 1620 1228 1622
rect 1211 1619 1212 1620
rect 1206 1618 1212 1619
rect 1227 1619 1228 1620
rect 1232 1619 1233 1623
rect 1227 1618 1233 1619
rect 1379 1623 1385 1624
rect 1379 1619 1380 1623
rect 1384 1622 1385 1623
rect 1410 1623 1416 1624
rect 1410 1622 1411 1623
rect 1384 1620 1411 1622
rect 1384 1619 1385 1620
rect 1379 1618 1385 1619
rect 1410 1619 1411 1620
rect 1415 1619 1416 1623
rect 1410 1618 1416 1619
rect 1531 1623 1537 1624
rect 1531 1619 1532 1623
rect 1536 1622 1537 1623
rect 1562 1623 1568 1624
rect 1562 1622 1563 1623
rect 1536 1620 1563 1622
rect 1536 1619 1537 1620
rect 1531 1618 1537 1619
rect 1562 1619 1563 1620
rect 1567 1619 1568 1623
rect 1562 1618 1568 1619
rect 1683 1623 1692 1624
rect 1683 1619 1684 1623
rect 1691 1619 1692 1623
rect 1683 1618 1692 1619
rect 2618 1615 2624 1616
rect 2618 1614 2619 1615
rect 2611 1613 2619 1614
rect 1923 1611 1929 1612
rect 1923 1607 1924 1611
rect 1928 1610 1929 1611
rect 1974 1611 1980 1612
rect 1974 1610 1975 1611
rect 1928 1608 1975 1610
rect 1928 1607 1929 1608
rect 1923 1606 1929 1607
rect 1974 1607 1975 1608
rect 1979 1607 1980 1611
rect 1974 1606 1980 1607
rect 2043 1611 2049 1612
rect 2043 1607 2044 1611
rect 2048 1610 2049 1611
rect 2082 1611 2088 1612
rect 2082 1610 2083 1611
rect 2048 1608 2083 1610
rect 2048 1607 2049 1608
rect 2043 1606 2049 1607
rect 2082 1607 2083 1608
rect 2087 1607 2088 1611
rect 2082 1606 2088 1607
rect 2111 1611 2117 1612
rect 2111 1607 2112 1611
rect 2116 1610 2117 1611
rect 2179 1611 2185 1612
rect 2179 1610 2180 1611
rect 2116 1608 2180 1610
rect 2116 1607 2117 1608
rect 2111 1606 2117 1607
rect 2179 1607 2180 1608
rect 2184 1607 2185 1611
rect 2179 1606 2185 1607
rect 2315 1611 2321 1612
rect 2315 1607 2316 1611
rect 2320 1610 2321 1611
rect 2359 1611 2365 1612
rect 2359 1610 2360 1611
rect 2320 1608 2360 1610
rect 2320 1607 2321 1608
rect 2315 1606 2321 1607
rect 2359 1607 2360 1608
rect 2364 1607 2365 1611
rect 2359 1606 2365 1607
rect 2459 1611 2468 1612
rect 2459 1607 2460 1611
rect 2467 1607 2468 1611
rect 2611 1609 2612 1613
rect 2616 1611 2619 1613
rect 2623 1611 2624 1615
rect 2616 1610 2624 1611
rect 2679 1611 2685 1612
rect 2616 1609 2617 1610
rect 2611 1608 2617 1609
rect 2459 1606 2468 1607
rect 2679 1607 2680 1611
rect 2684 1610 2685 1611
rect 2771 1611 2777 1612
rect 2771 1610 2772 1611
rect 2684 1608 2772 1610
rect 2684 1607 2685 1608
rect 2679 1606 2685 1607
rect 2771 1607 2772 1608
rect 2776 1607 2777 1611
rect 2771 1606 2777 1607
rect 2863 1611 2869 1612
rect 2863 1607 2864 1611
rect 2868 1610 2869 1611
rect 2939 1611 2945 1612
rect 2939 1610 2940 1611
rect 2868 1608 2940 1610
rect 2868 1607 2869 1608
rect 2863 1606 2869 1607
rect 2939 1607 2940 1608
rect 2944 1607 2945 1611
rect 2939 1606 2945 1607
rect 3023 1611 3029 1612
rect 3023 1607 3024 1611
rect 3028 1610 3029 1611
rect 3123 1611 3129 1612
rect 3123 1610 3124 1611
rect 3028 1608 3124 1610
rect 3028 1607 3029 1608
rect 3023 1606 3029 1607
rect 3123 1607 3124 1608
rect 3128 1607 3129 1611
rect 3123 1606 3129 1607
rect 3307 1611 3316 1612
rect 3307 1607 3308 1611
rect 3315 1607 3316 1611
rect 3307 1606 3316 1607
rect 3498 1611 3505 1612
rect 3498 1607 3499 1611
rect 3504 1607 3505 1611
rect 3498 1606 3505 1607
rect 251 1603 260 1604
rect 251 1599 252 1603
rect 259 1599 260 1603
rect 251 1598 260 1599
rect 327 1603 333 1604
rect 327 1599 328 1603
rect 332 1602 333 1603
rect 379 1603 385 1604
rect 379 1602 380 1603
rect 332 1600 380 1602
rect 332 1599 333 1600
rect 327 1598 333 1599
rect 379 1599 380 1600
rect 384 1599 385 1603
rect 379 1598 385 1599
rect 439 1603 445 1604
rect 439 1599 440 1603
rect 444 1602 445 1603
rect 515 1603 521 1604
rect 515 1602 516 1603
rect 444 1600 516 1602
rect 444 1599 445 1600
rect 439 1598 445 1599
rect 515 1599 516 1600
rect 520 1599 521 1603
rect 515 1598 521 1599
rect 650 1603 657 1604
rect 650 1599 651 1603
rect 656 1599 657 1603
rect 650 1598 657 1599
rect 711 1603 717 1604
rect 711 1599 712 1603
rect 716 1602 717 1603
rect 787 1603 793 1604
rect 787 1602 788 1603
rect 716 1600 788 1602
rect 716 1599 717 1600
rect 711 1598 717 1599
rect 787 1599 788 1600
rect 792 1599 793 1603
rect 787 1598 793 1599
rect 931 1603 937 1604
rect 931 1599 932 1603
rect 936 1602 937 1603
rect 954 1603 960 1604
rect 954 1602 955 1603
rect 936 1600 955 1602
rect 936 1599 937 1600
rect 931 1598 937 1599
rect 954 1599 955 1600
rect 959 1599 960 1603
rect 954 1598 960 1599
rect 999 1603 1005 1604
rect 999 1599 1000 1603
rect 1004 1602 1005 1603
rect 1083 1603 1089 1604
rect 1083 1602 1084 1603
rect 1004 1600 1084 1602
rect 1004 1599 1005 1600
rect 999 1598 1005 1599
rect 1083 1599 1084 1600
rect 1088 1599 1089 1603
rect 1083 1598 1089 1599
rect 1174 1603 1180 1604
rect 1174 1599 1175 1603
rect 1179 1602 1180 1603
rect 1243 1603 1249 1604
rect 1243 1602 1244 1603
rect 1179 1600 1244 1602
rect 1179 1599 1180 1600
rect 1174 1598 1180 1599
rect 1243 1599 1244 1600
rect 1248 1599 1249 1603
rect 1243 1598 1249 1599
rect 1403 1603 1409 1604
rect 1403 1599 1404 1603
rect 1408 1602 1409 1603
rect 1415 1603 1421 1604
rect 1415 1602 1416 1603
rect 1408 1600 1416 1602
rect 1408 1599 1409 1600
rect 1403 1598 1409 1599
rect 1415 1599 1416 1600
rect 1420 1599 1421 1603
rect 1415 1598 1421 1599
rect 1479 1603 1485 1604
rect 1479 1599 1480 1603
rect 1484 1602 1485 1603
rect 1571 1603 1577 1604
rect 1571 1602 1572 1603
rect 1484 1600 1572 1602
rect 1484 1599 1485 1600
rect 1479 1598 1485 1599
rect 1571 1599 1572 1600
rect 1576 1599 1577 1603
rect 1571 1598 1577 1599
rect 1894 1601 1900 1602
rect 1894 1597 1895 1601
rect 1899 1597 1900 1601
rect 1894 1596 1900 1597
rect 2014 1601 2020 1602
rect 2014 1597 2015 1601
rect 2019 1597 2020 1601
rect 2014 1596 2020 1597
rect 2150 1601 2156 1602
rect 2150 1597 2151 1601
rect 2155 1597 2156 1601
rect 2150 1596 2156 1597
rect 2286 1601 2292 1602
rect 2286 1597 2287 1601
rect 2291 1597 2292 1601
rect 2286 1596 2292 1597
rect 2430 1601 2436 1602
rect 2430 1597 2431 1601
rect 2435 1597 2436 1601
rect 2430 1596 2436 1597
rect 2582 1601 2588 1602
rect 2582 1597 2583 1601
rect 2587 1597 2588 1601
rect 2582 1596 2588 1597
rect 2742 1601 2748 1602
rect 2742 1597 2743 1601
rect 2747 1597 2748 1601
rect 2742 1596 2748 1597
rect 2910 1601 2916 1602
rect 2910 1597 2911 1601
rect 2915 1597 2916 1601
rect 2910 1596 2916 1597
rect 3094 1601 3100 1602
rect 3094 1597 3095 1601
rect 3099 1597 3100 1601
rect 3094 1596 3100 1597
rect 3278 1601 3284 1602
rect 3278 1597 3279 1601
rect 3283 1597 3284 1601
rect 3278 1596 3284 1597
rect 3470 1601 3476 1602
rect 3470 1597 3471 1601
rect 3475 1597 3476 1601
rect 3470 1596 3476 1597
rect 222 1593 228 1594
rect 222 1589 223 1593
rect 227 1589 228 1593
rect 222 1588 228 1589
rect 350 1593 356 1594
rect 350 1589 351 1593
rect 355 1589 356 1593
rect 350 1588 356 1589
rect 486 1593 492 1594
rect 486 1589 487 1593
rect 491 1589 492 1593
rect 486 1588 492 1589
rect 622 1593 628 1594
rect 622 1589 623 1593
rect 627 1589 628 1593
rect 622 1588 628 1589
rect 758 1593 764 1594
rect 758 1589 759 1593
rect 763 1589 764 1593
rect 758 1588 764 1589
rect 902 1593 908 1594
rect 902 1589 903 1593
rect 907 1589 908 1593
rect 902 1588 908 1589
rect 1054 1593 1060 1594
rect 1054 1589 1055 1593
rect 1059 1589 1060 1593
rect 1054 1588 1060 1589
rect 1214 1593 1220 1594
rect 1214 1589 1215 1593
rect 1219 1589 1220 1593
rect 1214 1588 1220 1589
rect 1374 1593 1380 1594
rect 1374 1589 1375 1593
rect 1379 1589 1380 1593
rect 1374 1588 1380 1589
rect 1542 1593 1548 1594
rect 1542 1589 1543 1593
rect 1547 1589 1548 1593
rect 1542 1588 1548 1589
rect 1862 1588 1868 1589
rect 3574 1588 3580 1589
rect 1862 1584 1863 1588
rect 1867 1584 1868 1588
rect 1958 1587 1964 1588
rect 1958 1586 1959 1587
rect 1949 1584 1959 1586
rect 1862 1583 1868 1584
rect 1958 1583 1959 1584
rect 1963 1583 1964 1587
rect 2679 1587 2685 1588
rect 2679 1586 2680 1587
rect 2637 1584 2680 1586
rect 1958 1582 1964 1583
rect 1974 1583 1980 1584
rect 110 1580 116 1581
rect 1822 1580 1828 1581
rect 110 1576 111 1580
rect 115 1576 116 1580
rect 327 1579 333 1580
rect 327 1578 328 1579
rect 277 1576 328 1578
rect 110 1575 116 1576
rect 327 1575 328 1576
rect 332 1575 333 1579
rect 439 1579 445 1580
rect 439 1578 440 1579
rect 405 1576 440 1578
rect 327 1574 333 1575
rect 439 1575 440 1576
rect 444 1575 445 1579
rect 711 1579 717 1580
rect 711 1578 712 1579
rect 677 1576 712 1578
rect 439 1574 445 1575
rect 711 1575 712 1576
rect 716 1575 717 1579
rect 999 1579 1005 1580
rect 999 1578 1000 1579
rect 957 1576 1000 1578
rect 711 1574 717 1575
rect 750 1575 756 1576
rect 750 1571 751 1575
rect 755 1574 756 1575
rect 999 1575 1000 1576
rect 1004 1575 1005 1579
rect 1174 1579 1180 1580
rect 1174 1578 1175 1579
rect 1109 1576 1175 1578
rect 999 1574 1005 1575
rect 1174 1575 1175 1576
rect 1179 1575 1180 1579
rect 1479 1579 1485 1580
rect 1479 1578 1480 1579
rect 1429 1576 1480 1578
rect 1174 1574 1180 1575
rect 1206 1575 1212 1576
rect 755 1572 777 1574
rect 755 1571 756 1572
rect 750 1570 756 1571
rect 1206 1571 1207 1575
rect 1211 1574 1212 1575
rect 1479 1575 1480 1576
rect 1484 1575 1485 1579
rect 1822 1576 1823 1580
rect 1827 1576 1828 1580
rect 1974 1579 1975 1583
rect 1979 1582 1980 1583
rect 2082 1583 2088 1584
rect 1979 1580 2033 1582
rect 1979 1579 1980 1580
rect 1974 1578 1980 1579
rect 2082 1579 2083 1583
rect 2087 1582 2088 1583
rect 2359 1583 2365 1584
rect 2087 1580 2169 1582
rect 2087 1579 2088 1580
rect 2082 1578 2088 1579
rect 2359 1579 2360 1583
rect 2364 1582 2365 1583
rect 2679 1583 2680 1584
rect 2684 1583 2685 1587
rect 2863 1587 2869 1588
rect 2863 1586 2864 1587
rect 2797 1584 2864 1586
rect 2679 1582 2685 1583
rect 2863 1583 2864 1584
rect 2868 1583 2869 1587
rect 3023 1587 3029 1588
rect 3023 1586 3024 1587
rect 2965 1584 3024 1586
rect 2863 1582 2869 1583
rect 3023 1583 3024 1584
rect 3028 1583 3029 1587
rect 3574 1584 3575 1588
rect 3579 1584 3580 1588
rect 3023 1582 3029 1583
rect 3270 1583 3276 1584
rect 3574 1583 3580 1584
rect 2364 1580 2449 1582
rect 2364 1579 2365 1580
rect 2359 1578 2365 1579
rect 3270 1579 3271 1583
rect 3275 1582 3276 1583
rect 3275 1580 3297 1582
rect 3275 1579 3276 1580
rect 3270 1578 3276 1579
rect 1822 1575 1828 1576
rect 1479 1574 1485 1575
rect 1211 1572 1233 1574
rect 1211 1571 1212 1572
rect 1206 1570 1212 1571
rect 1862 1571 1868 1572
rect 1862 1567 1863 1571
rect 1867 1567 1868 1571
rect 1862 1566 1868 1567
rect 2222 1571 2228 1572
rect 2222 1567 2223 1571
rect 2227 1570 2228 1571
rect 3018 1571 3024 1572
rect 2227 1568 2297 1570
rect 2227 1567 2228 1568
rect 2222 1566 2228 1567
rect 3018 1567 3019 1571
rect 3023 1570 3024 1571
rect 3574 1571 3580 1572
rect 3023 1568 3105 1570
rect 3023 1567 3024 1568
rect 3018 1566 3024 1567
rect 3574 1567 3575 1571
rect 3579 1567 3580 1571
rect 3574 1566 3580 1567
rect 110 1563 116 1564
rect 110 1559 111 1563
rect 115 1559 116 1563
rect 110 1558 116 1559
rect 462 1563 468 1564
rect 462 1559 463 1563
rect 467 1562 468 1563
rect 1542 1563 1548 1564
rect 467 1560 497 1562
rect 467 1559 468 1560
rect 462 1558 468 1559
rect 1542 1559 1543 1563
rect 1547 1562 1548 1563
rect 1822 1563 1828 1564
rect 1547 1560 1553 1562
rect 1547 1559 1548 1560
rect 1542 1558 1548 1559
rect 1822 1559 1823 1563
rect 1827 1559 1828 1563
rect 1822 1558 1828 1559
rect 1886 1561 1892 1562
rect 1886 1557 1887 1561
rect 1891 1557 1892 1561
rect 1886 1556 1892 1557
rect 2006 1561 2012 1562
rect 2006 1557 2007 1561
rect 2011 1557 2012 1561
rect 2006 1556 2012 1557
rect 2142 1561 2148 1562
rect 2142 1557 2143 1561
rect 2147 1557 2148 1561
rect 2142 1556 2148 1557
rect 2278 1561 2284 1562
rect 2278 1557 2279 1561
rect 2283 1557 2284 1561
rect 2278 1556 2284 1557
rect 2422 1561 2428 1562
rect 2422 1557 2423 1561
rect 2427 1557 2428 1561
rect 2422 1556 2428 1557
rect 2574 1561 2580 1562
rect 2574 1557 2575 1561
rect 2579 1557 2580 1561
rect 2574 1556 2580 1557
rect 2734 1561 2740 1562
rect 2734 1557 2735 1561
rect 2739 1557 2740 1561
rect 2734 1556 2740 1557
rect 2902 1561 2908 1562
rect 2902 1557 2903 1561
rect 2907 1557 2908 1561
rect 2902 1556 2908 1557
rect 3086 1561 3092 1562
rect 3086 1557 3087 1561
rect 3091 1557 3092 1561
rect 3086 1556 3092 1557
rect 3270 1561 3276 1562
rect 3270 1557 3271 1561
rect 3275 1557 3276 1561
rect 3270 1556 3276 1557
rect 3462 1561 3468 1562
rect 3462 1557 3463 1561
rect 3467 1557 3468 1561
rect 3462 1556 3468 1557
rect 3511 1555 3520 1556
rect 214 1553 220 1554
rect 214 1549 215 1553
rect 219 1549 220 1553
rect 214 1548 220 1549
rect 342 1553 348 1554
rect 342 1549 343 1553
rect 347 1549 348 1553
rect 342 1548 348 1549
rect 478 1553 484 1554
rect 478 1549 479 1553
rect 483 1549 484 1553
rect 478 1548 484 1549
rect 614 1553 620 1554
rect 614 1549 615 1553
rect 619 1549 620 1553
rect 614 1548 620 1549
rect 750 1553 756 1554
rect 750 1549 751 1553
rect 755 1549 756 1553
rect 750 1548 756 1549
rect 894 1553 900 1554
rect 894 1549 895 1553
rect 899 1549 900 1553
rect 894 1548 900 1549
rect 1046 1553 1052 1554
rect 1046 1549 1047 1553
rect 1051 1549 1052 1553
rect 1046 1548 1052 1549
rect 1206 1553 1212 1554
rect 1206 1549 1207 1553
rect 1211 1549 1212 1553
rect 1206 1548 1212 1549
rect 1366 1553 1372 1554
rect 1366 1549 1367 1553
rect 1371 1549 1372 1553
rect 1366 1548 1372 1549
rect 1534 1553 1540 1554
rect 1534 1549 1535 1553
rect 1539 1549 1540 1553
rect 3511 1551 3512 1555
rect 3519 1551 3520 1555
rect 3511 1550 3520 1551
rect 1534 1548 1540 1549
rect 1886 1531 1892 1532
rect 134 1527 140 1528
rect 134 1523 135 1527
rect 139 1523 140 1527
rect 134 1522 140 1523
rect 270 1527 276 1528
rect 270 1523 271 1527
rect 275 1523 276 1527
rect 270 1522 276 1523
rect 422 1527 428 1528
rect 422 1523 423 1527
rect 427 1523 428 1527
rect 422 1522 428 1523
rect 582 1527 588 1528
rect 582 1523 583 1527
rect 587 1523 588 1527
rect 582 1522 588 1523
rect 734 1527 740 1528
rect 734 1523 735 1527
rect 739 1523 740 1527
rect 734 1522 740 1523
rect 886 1527 892 1528
rect 886 1523 887 1527
rect 891 1523 892 1527
rect 886 1522 892 1523
rect 1038 1527 1044 1528
rect 1038 1523 1039 1527
rect 1043 1523 1044 1527
rect 1038 1522 1044 1523
rect 1190 1527 1196 1528
rect 1190 1523 1191 1527
rect 1195 1523 1196 1527
rect 1190 1522 1196 1523
rect 1342 1527 1348 1528
rect 1342 1523 1343 1527
rect 1347 1523 1348 1527
rect 1342 1522 1348 1523
rect 1494 1527 1500 1528
rect 1494 1523 1495 1527
rect 1499 1523 1500 1527
rect 1886 1527 1887 1531
rect 1891 1527 1892 1531
rect 1886 1526 1892 1527
rect 2022 1531 2028 1532
rect 2022 1527 2023 1531
rect 2027 1527 2028 1531
rect 2022 1526 2028 1527
rect 2182 1531 2188 1532
rect 2182 1527 2183 1531
rect 2187 1527 2188 1531
rect 2182 1526 2188 1527
rect 2342 1531 2348 1532
rect 2342 1527 2343 1531
rect 2347 1527 2348 1531
rect 2342 1526 2348 1527
rect 2502 1531 2508 1532
rect 2502 1527 2503 1531
rect 2507 1527 2508 1531
rect 2502 1526 2508 1527
rect 2662 1531 2668 1532
rect 2662 1527 2663 1531
rect 2667 1527 2668 1531
rect 2662 1526 2668 1527
rect 2822 1531 2828 1532
rect 2822 1527 2823 1531
rect 2827 1527 2828 1531
rect 2822 1526 2828 1527
rect 2982 1531 2988 1532
rect 2982 1527 2983 1531
rect 2987 1527 2988 1531
rect 2982 1526 2988 1527
rect 3150 1531 3156 1532
rect 3150 1527 3151 1531
rect 3155 1527 3156 1531
rect 3150 1526 3156 1527
rect 3318 1531 3324 1532
rect 3318 1527 3319 1531
rect 3323 1527 3324 1531
rect 3318 1526 3324 1527
rect 3478 1531 3484 1532
rect 3478 1527 3479 1531
rect 3483 1527 3484 1531
rect 3478 1526 3484 1527
rect 1494 1522 1500 1523
rect 2111 1523 2117 1524
rect 2111 1522 2112 1523
rect 1862 1521 1868 1522
rect 650 1519 656 1520
rect 650 1518 651 1519
rect 110 1517 116 1518
rect 110 1513 111 1517
rect 115 1513 116 1517
rect 641 1516 651 1518
rect 650 1515 651 1516
rect 655 1515 656 1519
rect 954 1519 960 1520
rect 954 1518 955 1519
rect 945 1516 955 1518
rect 650 1514 656 1515
rect 954 1515 955 1516
rect 959 1515 960 1519
rect 954 1514 960 1515
rect 1822 1517 1828 1518
rect 110 1512 116 1513
rect 1822 1513 1823 1517
rect 1827 1513 1828 1517
rect 1862 1517 1863 1521
rect 1867 1517 1868 1521
rect 2081 1520 2112 1522
rect 2111 1519 2112 1520
rect 2116 1519 2117 1523
rect 2111 1518 2117 1519
rect 3078 1523 3084 1524
rect 3078 1519 3079 1523
rect 3083 1522 3084 1523
rect 3310 1523 3316 1524
rect 3083 1520 3169 1522
rect 3083 1519 3084 1520
rect 3078 1518 3084 1519
rect 3310 1519 3311 1523
rect 3315 1522 3316 1523
rect 3315 1520 3337 1522
rect 3574 1521 3580 1522
rect 3315 1519 3316 1520
rect 3310 1518 3316 1519
rect 1862 1516 1868 1517
rect 3574 1517 3575 1521
rect 3579 1517 3580 1521
rect 3574 1516 3580 1517
rect 1822 1512 1828 1513
rect 2015 1507 2021 1508
rect 2015 1506 2016 1507
rect 1862 1504 1868 1505
rect 1949 1504 2016 1506
rect 207 1503 213 1504
rect 110 1500 116 1501
rect 110 1496 111 1500
rect 115 1496 116 1500
rect 110 1495 116 1496
rect 196 1496 198 1501
rect 207 1499 208 1503
rect 212 1502 213 1503
rect 338 1503 344 1504
rect 212 1500 297 1502
rect 212 1499 213 1500
rect 207 1498 213 1499
rect 338 1499 339 1503
rect 343 1502 344 1503
rect 650 1503 656 1504
rect 343 1500 449 1502
rect 343 1499 344 1500
rect 338 1498 344 1499
rect 650 1499 651 1503
rect 655 1502 656 1503
rect 954 1503 960 1504
rect 655 1500 761 1502
rect 655 1499 656 1500
rect 650 1498 656 1499
rect 954 1499 955 1503
rect 959 1502 960 1503
rect 1335 1503 1341 1504
rect 1335 1502 1336 1503
rect 959 1500 1065 1502
rect 1253 1500 1336 1502
rect 959 1499 960 1500
rect 954 1498 960 1499
rect 1335 1499 1336 1500
rect 1340 1499 1341 1503
rect 1410 1503 1416 1504
rect 1410 1502 1411 1503
rect 1405 1500 1411 1502
rect 1335 1498 1341 1499
rect 1410 1499 1411 1500
rect 1415 1499 1416 1503
rect 1410 1498 1416 1499
rect 1418 1503 1424 1504
rect 1418 1499 1419 1503
rect 1423 1502 1424 1503
rect 1423 1500 1521 1502
rect 1822 1500 1828 1501
rect 1423 1499 1424 1500
rect 1418 1498 1424 1499
rect 1822 1496 1823 1500
rect 1827 1496 1828 1500
rect 1862 1500 1863 1504
rect 1867 1500 1868 1504
rect 2015 1503 2016 1504
rect 2020 1503 2021 1507
rect 2335 1507 2341 1508
rect 2335 1506 2336 1507
rect 2245 1504 2336 1506
rect 2015 1502 2021 1503
rect 2335 1503 2336 1504
rect 2340 1503 2341 1507
rect 2495 1507 2501 1508
rect 2495 1506 2496 1507
rect 2405 1504 2496 1506
rect 2335 1502 2341 1503
rect 2495 1503 2496 1504
rect 2500 1503 2501 1507
rect 2730 1507 2736 1508
rect 2730 1506 2731 1507
rect 2495 1502 2501 1503
rect 1862 1499 1868 1500
rect 2564 1500 2566 1505
rect 2725 1504 2731 1506
rect 2730 1503 2731 1504
rect 2735 1503 2736 1507
rect 2975 1507 2981 1508
rect 2975 1506 2976 1507
rect 2885 1504 2976 1506
rect 2730 1502 2736 1503
rect 2975 1503 2976 1504
rect 2980 1503 2981 1507
rect 3143 1507 3149 1508
rect 3143 1506 3144 1507
rect 3045 1504 3144 1506
rect 2975 1502 2981 1503
rect 3143 1503 3144 1504
rect 3148 1503 3149 1507
rect 3546 1507 3552 1508
rect 3546 1506 3547 1507
rect 3541 1504 3547 1506
rect 3143 1502 3149 1503
rect 3546 1503 3547 1504
rect 3551 1503 3552 1507
rect 3546 1502 3552 1503
rect 3574 1504 3580 1505
rect 3574 1500 3575 1504
rect 3579 1500 3580 1504
rect 2564 1499 2572 1500
rect 3574 1499 3580 1500
rect 2564 1496 2567 1499
rect 196 1495 204 1496
rect 1822 1495 1828 1496
rect 2566 1495 2567 1496
rect 2571 1495 2572 1499
rect 196 1492 199 1495
rect 198 1491 199 1492
rect 203 1491 204 1495
rect 2566 1494 2572 1495
rect 198 1490 204 1491
rect 1894 1491 1900 1492
rect 142 1487 148 1488
rect 142 1483 143 1487
rect 147 1483 148 1487
rect 142 1482 148 1483
rect 278 1487 284 1488
rect 278 1483 279 1487
rect 283 1483 284 1487
rect 278 1482 284 1483
rect 430 1487 436 1488
rect 430 1483 431 1487
rect 435 1483 436 1487
rect 430 1482 436 1483
rect 590 1487 596 1488
rect 590 1483 591 1487
rect 595 1483 596 1487
rect 590 1482 596 1483
rect 742 1487 748 1488
rect 742 1483 743 1487
rect 747 1483 748 1487
rect 742 1482 748 1483
rect 894 1487 900 1488
rect 894 1483 895 1487
rect 899 1483 900 1487
rect 894 1482 900 1483
rect 1046 1487 1052 1488
rect 1046 1483 1047 1487
rect 1051 1483 1052 1487
rect 1046 1482 1052 1483
rect 1198 1487 1204 1488
rect 1198 1483 1199 1487
rect 1203 1483 1204 1487
rect 1198 1482 1204 1483
rect 1350 1487 1356 1488
rect 1350 1483 1351 1487
rect 1355 1483 1356 1487
rect 1350 1482 1356 1483
rect 1502 1487 1508 1488
rect 1502 1483 1503 1487
rect 1507 1483 1508 1487
rect 1894 1487 1895 1491
rect 1899 1487 1900 1491
rect 1894 1486 1900 1487
rect 2030 1491 2036 1492
rect 2030 1487 2031 1491
rect 2035 1487 2036 1491
rect 2030 1486 2036 1487
rect 2190 1491 2196 1492
rect 2190 1487 2191 1491
rect 2195 1487 2196 1491
rect 2190 1486 2196 1487
rect 2350 1491 2356 1492
rect 2350 1487 2351 1491
rect 2355 1487 2356 1491
rect 2350 1486 2356 1487
rect 2510 1491 2516 1492
rect 2510 1487 2511 1491
rect 2515 1487 2516 1491
rect 2510 1486 2516 1487
rect 2670 1491 2676 1492
rect 2670 1487 2671 1491
rect 2675 1487 2676 1491
rect 2670 1486 2676 1487
rect 2830 1491 2836 1492
rect 2830 1487 2831 1491
rect 2835 1487 2836 1491
rect 2830 1486 2836 1487
rect 2990 1491 2996 1492
rect 2990 1487 2991 1491
rect 2995 1487 2996 1491
rect 2990 1486 2996 1487
rect 3158 1491 3164 1492
rect 3158 1487 3159 1491
rect 3163 1487 3164 1491
rect 3158 1486 3164 1487
rect 3326 1491 3332 1492
rect 3326 1487 3327 1491
rect 3331 1487 3332 1491
rect 3326 1486 3332 1487
rect 3486 1491 3492 1492
rect 3486 1487 3487 1491
rect 3491 1487 3492 1491
rect 3486 1486 3492 1487
rect 1502 1482 1508 1483
rect 1807 1479 1813 1480
rect 171 1475 177 1476
rect 171 1471 172 1475
rect 176 1474 177 1475
rect 207 1475 213 1476
rect 207 1474 208 1475
rect 176 1472 208 1474
rect 176 1471 177 1472
rect 171 1470 177 1471
rect 207 1471 208 1472
rect 212 1471 213 1475
rect 207 1470 213 1471
rect 307 1475 313 1476
rect 307 1471 308 1475
rect 312 1474 313 1475
rect 338 1475 344 1476
rect 338 1474 339 1475
rect 312 1472 339 1474
rect 312 1471 313 1472
rect 307 1470 313 1471
rect 338 1471 339 1472
rect 343 1471 344 1475
rect 338 1470 344 1471
rect 459 1475 468 1476
rect 459 1471 460 1475
rect 467 1471 468 1475
rect 459 1470 468 1471
rect 619 1475 625 1476
rect 619 1471 620 1475
rect 624 1474 625 1475
rect 650 1475 656 1476
rect 650 1474 651 1475
rect 624 1472 651 1474
rect 624 1471 625 1472
rect 619 1470 625 1471
rect 650 1471 651 1472
rect 655 1471 656 1475
rect 650 1470 656 1471
rect 727 1475 733 1476
rect 727 1471 728 1475
rect 732 1474 733 1475
rect 771 1475 777 1476
rect 771 1474 772 1475
rect 732 1472 772 1474
rect 732 1471 733 1472
rect 727 1470 733 1471
rect 771 1471 772 1472
rect 776 1471 777 1475
rect 771 1470 777 1471
rect 923 1475 929 1476
rect 923 1471 924 1475
rect 928 1474 929 1475
rect 954 1475 960 1476
rect 954 1474 955 1475
rect 928 1472 955 1474
rect 928 1471 929 1472
rect 923 1470 929 1471
rect 954 1471 955 1472
rect 959 1471 960 1475
rect 954 1470 960 1471
rect 1075 1475 1084 1476
rect 1075 1471 1076 1475
rect 1083 1471 1084 1475
rect 1075 1470 1084 1471
rect 1227 1475 1233 1476
rect 1227 1471 1228 1475
rect 1232 1474 1233 1475
rect 1335 1475 1341 1476
rect 1232 1472 1330 1474
rect 1232 1471 1233 1472
rect 1227 1470 1233 1471
rect 1328 1466 1330 1472
rect 1335 1471 1336 1475
rect 1340 1474 1341 1475
rect 1379 1475 1385 1476
rect 1379 1474 1380 1475
rect 1340 1472 1380 1474
rect 1340 1471 1341 1472
rect 1335 1470 1341 1471
rect 1379 1471 1380 1472
rect 1384 1471 1385 1475
rect 1379 1470 1385 1471
rect 1531 1475 1537 1476
rect 1531 1471 1532 1475
rect 1536 1474 1537 1475
rect 1542 1475 1548 1476
rect 1542 1474 1543 1475
rect 1536 1472 1543 1474
rect 1536 1471 1537 1472
rect 1531 1470 1537 1471
rect 1542 1471 1543 1472
rect 1547 1471 1548 1475
rect 1807 1475 1808 1479
rect 1812 1478 1813 1479
rect 1923 1479 1929 1480
rect 1923 1478 1924 1479
rect 1812 1476 1924 1478
rect 1812 1475 1813 1476
rect 1807 1474 1813 1475
rect 1923 1475 1924 1476
rect 1928 1475 1929 1479
rect 1923 1474 1929 1475
rect 2015 1479 2021 1480
rect 2015 1475 2016 1479
rect 2020 1478 2021 1479
rect 2059 1479 2065 1480
rect 2059 1478 2060 1479
rect 2020 1476 2060 1478
rect 2020 1475 2021 1476
rect 2015 1474 2021 1475
rect 2059 1475 2060 1476
rect 2064 1475 2065 1479
rect 2059 1474 2065 1475
rect 2219 1479 2228 1480
rect 2219 1475 2220 1479
rect 2227 1475 2228 1479
rect 2219 1474 2228 1475
rect 2335 1479 2341 1480
rect 2335 1475 2336 1479
rect 2340 1478 2341 1479
rect 2379 1479 2385 1480
rect 2379 1478 2380 1479
rect 2340 1476 2380 1478
rect 2340 1475 2341 1476
rect 2335 1474 2341 1475
rect 2379 1475 2380 1476
rect 2384 1475 2385 1479
rect 2379 1474 2385 1475
rect 2495 1479 2501 1480
rect 2495 1475 2496 1479
rect 2500 1478 2501 1479
rect 2539 1479 2545 1480
rect 2539 1478 2540 1479
rect 2500 1476 2540 1478
rect 2500 1475 2501 1476
rect 2495 1474 2501 1475
rect 2539 1475 2540 1476
rect 2544 1475 2545 1479
rect 2539 1474 2545 1475
rect 2699 1479 2708 1480
rect 2699 1475 2700 1479
rect 2707 1475 2708 1479
rect 2699 1474 2708 1475
rect 2730 1479 2736 1480
rect 2730 1475 2731 1479
rect 2735 1478 2736 1479
rect 2859 1479 2865 1480
rect 2859 1478 2860 1479
rect 2735 1476 2860 1478
rect 2735 1475 2736 1476
rect 2730 1474 2736 1475
rect 2859 1475 2860 1476
rect 2864 1475 2865 1479
rect 2859 1474 2865 1475
rect 2975 1479 2981 1480
rect 2975 1475 2976 1479
rect 2980 1478 2981 1479
rect 3019 1479 3025 1480
rect 3019 1478 3020 1479
rect 2980 1476 3020 1478
rect 2980 1475 2981 1476
rect 2975 1474 2981 1475
rect 3019 1475 3020 1476
rect 3024 1475 3025 1479
rect 3019 1474 3025 1475
rect 3143 1479 3149 1480
rect 3143 1475 3144 1479
rect 3148 1478 3149 1479
rect 3187 1479 3193 1480
rect 3187 1478 3188 1479
rect 3148 1476 3188 1478
rect 3148 1475 3149 1476
rect 3143 1474 3149 1475
rect 3187 1475 3188 1476
rect 3192 1475 3193 1479
rect 3187 1474 3193 1475
rect 3350 1479 3361 1480
rect 3350 1475 3351 1479
rect 3355 1475 3356 1479
rect 3360 1475 3361 1479
rect 3350 1474 3361 1475
rect 3514 1479 3521 1480
rect 3514 1475 3515 1479
rect 3520 1475 3521 1479
rect 3514 1474 3521 1475
rect 1542 1470 1548 1471
rect 1418 1467 1424 1468
rect 1418 1466 1419 1467
rect 1328 1464 1419 1466
rect 1090 1463 1096 1464
rect 1090 1462 1091 1463
rect 820 1460 1091 1462
rect 820 1458 822 1460
rect 1090 1459 1091 1460
rect 1095 1459 1096 1463
rect 1418 1463 1419 1464
rect 1423 1463 1424 1467
rect 1418 1462 1424 1463
rect 1090 1458 1096 1459
rect 2211 1459 2217 1460
rect 819 1457 825 1458
rect 171 1455 177 1456
rect 171 1451 172 1455
rect 176 1454 177 1455
rect 198 1455 204 1456
rect 198 1454 199 1455
rect 176 1452 199 1454
rect 176 1451 177 1452
rect 171 1450 177 1451
rect 198 1451 199 1452
rect 203 1451 204 1455
rect 198 1450 204 1451
rect 207 1455 213 1456
rect 207 1451 208 1455
rect 212 1454 213 1455
rect 291 1455 297 1456
rect 291 1454 292 1455
rect 212 1452 292 1454
rect 212 1451 213 1452
rect 207 1450 213 1451
rect 291 1451 292 1452
rect 296 1451 297 1455
rect 291 1450 297 1451
rect 351 1455 357 1456
rect 351 1451 352 1455
rect 356 1454 357 1455
rect 427 1455 433 1456
rect 427 1454 428 1455
rect 356 1452 428 1454
rect 356 1451 357 1452
rect 351 1450 357 1451
rect 427 1451 428 1452
rect 432 1451 433 1455
rect 427 1450 433 1451
rect 563 1455 569 1456
rect 563 1451 564 1455
rect 568 1454 569 1455
rect 615 1455 621 1456
rect 568 1452 610 1454
rect 568 1451 569 1452
rect 563 1450 569 1451
rect 608 1446 610 1452
rect 615 1451 616 1455
rect 620 1454 621 1455
rect 691 1455 697 1456
rect 691 1454 692 1455
rect 620 1452 692 1454
rect 620 1451 621 1452
rect 615 1450 621 1451
rect 691 1451 692 1452
rect 696 1451 697 1455
rect 819 1453 820 1457
rect 824 1453 825 1457
rect 819 1452 825 1453
rect 871 1455 877 1456
rect 691 1450 697 1451
rect 871 1451 872 1455
rect 876 1454 877 1455
rect 939 1455 945 1456
rect 939 1454 940 1455
rect 876 1452 940 1454
rect 876 1451 877 1452
rect 871 1450 877 1451
rect 939 1451 940 1452
rect 944 1451 945 1455
rect 939 1450 945 1451
rect 983 1455 989 1456
rect 983 1451 984 1455
rect 988 1454 989 1455
rect 1051 1455 1057 1456
rect 1051 1454 1052 1455
rect 988 1452 1052 1454
rect 988 1451 989 1452
rect 983 1450 989 1451
rect 1051 1451 1052 1452
rect 1056 1451 1057 1455
rect 1051 1450 1057 1451
rect 1171 1455 1177 1456
rect 1171 1451 1172 1455
rect 1176 1454 1177 1455
rect 1210 1455 1216 1456
rect 1210 1454 1211 1455
rect 1176 1452 1211 1454
rect 1176 1451 1177 1452
rect 1171 1450 1177 1451
rect 1210 1451 1211 1452
rect 1215 1451 1216 1455
rect 1210 1450 1216 1451
rect 1291 1455 1297 1456
rect 1291 1451 1292 1455
rect 1296 1454 1297 1455
rect 1402 1455 1408 1456
rect 1402 1454 1403 1455
rect 1296 1452 1403 1454
rect 1296 1451 1297 1452
rect 1291 1450 1297 1451
rect 1402 1451 1403 1452
rect 1407 1451 1408 1455
rect 1402 1450 1408 1451
rect 1410 1455 1417 1456
rect 1410 1451 1411 1455
rect 1416 1451 1417 1455
rect 1410 1450 1417 1451
rect 1463 1455 1469 1456
rect 1463 1451 1464 1455
rect 1468 1454 1469 1455
rect 1531 1455 1537 1456
rect 1531 1454 1532 1455
rect 1468 1452 1532 1454
rect 1468 1451 1469 1452
rect 1463 1450 1469 1451
rect 1531 1451 1532 1452
rect 1536 1451 1537 1455
rect 1531 1450 1537 1451
rect 1591 1455 1597 1456
rect 1591 1451 1592 1455
rect 1596 1454 1597 1455
rect 1659 1455 1665 1456
rect 1659 1454 1660 1455
rect 1596 1452 1660 1454
rect 1596 1451 1597 1452
rect 1591 1450 1597 1451
rect 1659 1451 1660 1452
rect 1664 1451 1665 1455
rect 1659 1450 1665 1451
rect 1703 1455 1709 1456
rect 1703 1451 1704 1455
rect 1708 1454 1709 1455
rect 1763 1455 1769 1456
rect 1763 1454 1764 1455
rect 1708 1452 1764 1454
rect 1708 1451 1709 1452
rect 1703 1450 1709 1451
rect 1763 1451 1764 1452
rect 1768 1451 1769 1455
rect 2211 1455 2212 1459
rect 2216 1458 2217 1459
rect 2222 1459 2228 1460
rect 2222 1458 2223 1459
rect 2216 1456 2223 1458
rect 2216 1455 2217 1456
rect 2211 1454 2217 1455
rect 2222 1455 2223 1456
rect 2227 1455 2228 1459
rect 2222 1454 2228 1455
rect 2287 1459 2293 1460
rect 2287 1455 2288 1459
rect 2292 1458 2293 1459
rect 2387 1459 2393 1460
rect 2387 1458 2388 1459
rect 2292 1456 2388 1458
rect 2292 1455 2293 1456
rect 2287 1454 2293 1455
rect 2387 1455 2388 1456
rect 2392 1455 2393 1459
rect 2387 1454 2393 1455
rect 2555 1459 2561 1460
rect 2555 1455 2556 1459
rect 2560 1458 2561 1459
rect 2566 1459 2572 1460
rect 2566 1458 2567 1459
rect 2560 1456 2567 1458
rect 2560 1455 2561 1456
rect 2555 1454 2561 1455
rect 2566 1455 2567 1456
rect 2571 1455 2572 1459
rect 2566 1454 2572 1455
rect 2715 1459 2724 1460
rect 2715 1455 2716 1459
rect 2723 1455 2724 1459
rect 2715 1454 2724 1455
rect 2823 1459 2829 1460
rect 2823 1455 2824 1459
rect 2828 1458 2829 1459
rect 2875 1459 2881 1460
rect 2875 1458 2876 1459
rect 2828 1456 2876 1458
rect 2828 1455 2829 1456
rect 2823 1454 2829 1455
rect 2875 1455 2876 1456
rect 2880 1455 2881 1459
rect 2875 1454 2881 1455
rect 2943 1459 2949 1460
rect 2943 1455 2944 1459
rect 2948 1458 2949 1459
rect 3035 1459 3041 1460
rect 3035 1458 3036 1459
rect 2948 1456 3036 1458
rect 2948 1455 2949 1456
rect 2943 1454 2949 1455
rect 3035 1455 3036 1456
rect 3040 1455 3041 1459
rect 3035 1454 3041 1455
rect 3111 1459 3117 1460
rect 3111 1455 3112 1459
rect 3116 1458 3117 1459
rect 3203 1459 3209 1460
rect 3203 1458 3204 1459
rect 3116 1456 3204 1458
rect 3116 1455 3117 1456
rect 3111 1454 3117 1455
rect 3203 1455 3204 1456
rect 3208 1455 3209 1459
rect 3203 1454 3209 1455
rect 3279 1459 3285 1460
rect 3279 1455 3280 1459
rect 3284 1458 3285 1459
rect 3371 1459 3377 1460
rect 3371 1458 3372 1459
rect 3284 1456 3372 1458
rect 3284 1455 3285 1456
rect 3279 1454 3285 1455
rect 3371 1455 3372 1456
rect 3376 1455 3377 1459
rect 3371 1454 3377 1455
rect 3515 1459 3521 1460
rect 3515 1455 3516 1459
rect 3520 1458 3521 1459
rect 3546 1459 3552 1460
rect 3546 1458 3547 1459
rect 3520 1456 3547 1458
rect 3520 1455 3521 1456
rect 3515 1454 3521 1455
rect 3546 1455 3547 1456
rect 3551 1455 3552 1459
rect 3546 1454 3552 1455
rect 1763 1450 1769 1451
rect 2182 1449 2188 1450
rect 622 1447 628 1448
rect 622 1446 623 1447
rect 142 1445 148 1446
rect 142 1441 143 1445
rect 147 1441 148 1445
rect 142 1440 148 1441
rect 262 1445 268 1446
rect 262 1441 263 1445
rect 267 1441 268 1445
rect 262 1440 268 1441
rect 398 1445 404 1446
rect 398 1441 399 1445
rect 403 1441 404 1445
rect 398 1440 404 1441
rect 534 1445 540 1446
rect 534 1441 535 1445
rect 539 1441 540 1445
rect 608 1444 623 1446
rect 622 1443 623 1444
rect 627 1443 628 1447
rect 622 1442 628 1443
rect 662 1445 668 1446
rect 534 1440 540 1441
rect 662 1441 663 1445
rect 667 1441 668 1445
rect 662 1440 668 1441
rect 790 1445 796 1446
rect 790 1441 791 1445
rect 795 1441 796 1445
rect 790 1440 796 1441
rect 910 1445 916 1446
rect 910 1441 911 1445
rect 915 1441 916 1445
rect 910 1440 916 1441
rect 1022 1445 1028 1446
rect 1022 1441 1023 1445
rect 1027 1441 1028 1445
rect 1022 1440 1028 1441
rect 1142 1445 1148 1446
rect 1142 1441 1143 1445
rect 1147 1441 1148 1445
rect 1142 1440 1148 1441
rect 1262 1445 1268 1446
rect 1262 1441 1263 1445
rect 1267 1441 1268 1445
rect 1262 1440 1268 1441
rect 1382 1445 1388 1446
rect 1382 1441 1383 1445
rect 1387 1441 1388 1445
rect 1382 1440 1388 1441
rect 1502 1445 1508 1446
rect 1502 1441 1503 1445
rect 1507 1441 1508 1445
rect 1502 1440 1508 1441
rect 1630 1445 1636 1446
rect 1630 1441 1631 1445
rect 1635 1441 1636 1445
rect 1630 1440 1636 1441
rect 1734 1445 1740 1446
rect 1734 1441 1735 1445
rect 1739 1441 1740 1445
rect 2182 1445 2183 1449
rect 2187 1445 2188 1449
rect 2182 1444 2188 1445
rect 2358 1449 2364 1450
rect 2358 1445 2359 1449
rect 2363 1445 2364 1449
rect 2358 1444 2364 1445
rect 2526 1449 2532 1450
rect 2526 1445 2527 1449
rect 2531 1445 2532 1449
rect 2526 1444 2532 1445
rect 2686 1449 2692 1450
rect 2686 1445 2687 1449
rect 2691 1445 2692 1449
rect 2686 1444 2692 1445
rect 2846 1449 2852 1450
rect 2846 1445 2847 1449
rect 2851 1445 2852 1449
rect 2846 1444 2852 1445
rect 3006 1449 3012 1450
rect 3006 1445 3007 1449
rect 3011 1445 3012 1449
rect 3006 1444 3012 1445
rect 3174 1449 3180 1450
rect 3174 1445 3175 1449
rect 3179 1445 3180 1449
rect 3174 1444 3180 1445
rect 3342 1449 3348 1450
rect 3342 1445 3343 1449
rect 3347 1445 3348 1449
rect 3342 1444 3348 1445
rect 3486 1449 3492 1450
rect 3486 1445 3487 1449
rect 3491 1445 3492 1449
rect 3486 1444 3492 1445
rect 1734 1440 1740 1441
rect 1078 1439 1084 1440
rect 1078 1438 1079 1439
rect 1076 1435 1079 1438
rect 1083 1435 1084 1439
rect 1076 1434 1084 1435
rect 1862 1436 1868 1437
rect 3574 1436 3580 1437
rect 110 1432 116 1433
rect 110 1428 111 1432
rect 115 1428 116 1432
rect 207 1431 213 1432
rect 207 1430 208 1431
rect 197 1428 208 1430
rect 110 1427 116 1428
rect 207 1427 208 1428
rect 212 1427 213 1431
rect 351 1431 357 1432
rect 351 1430 352 1431
rect 317 1428 352 1430
rect 207 1426 213 1427
rect 351 1427 352 1428
rect 356 1427 357 1431
rect 615 1431 621 1432
rect 615 1430 616 1431
rect 589 1428 616 1430
rect 351 1426 357 1427
rect 615 1427 616 1428
rect 620 1427 621 1431
rect 727 1431 733 1432
rect 727 1430 728 1431
rect 717 1428 728 1430
rect 615 1426 621 1427
rect 727 1427 728 1428
rect 732 1427 733 1431
rect 871 1431 877 1432
rect 871 1430 872 1431
rect 845 1428 872 1430
rect 727 1426 733 1427
rect 871 1427 872 1428
rect 876 1427 877 1431
rect 983 1431 989 1432
rect 983 1430 984 1431
rect 965 1428 984 1430
rect 871 1426 877 1427
rect 983 1427 984 1428
rect 988 1427 989 1431
rect 1076 1429 1078 1434
rect 1822 1432 1828 1433
rect 1463 1431 1469 1432
rect 1463 1430 1464 1431
rect 1437 1428 1464 1430
rect 983 1426 989 1427
rect 1090 1427 1096 1428
rect 1090 1423 1091 1427
rect 1095 1426 1096 1427
rect 1210 1427 1216 1428
rect 1095 1424 1161 1426
rect 1095 1423 1096 1424
rect 1090 1422 1096 1423
rect 1210 1423 1211 1427
rect 1215 1426 1216 1427
rect 1463 1427 1464 1428
rect 1468 1427 1469 1431
rect 1703 1431 1709 1432
rect 1703 1430 1704 1431
rect 1685 1428 1704 1430
rect 1463 1426 1469 1427
rect 1703 1427 1704 1428
rect 1708 1427 1709 1431
rect 1807 1431 1813 1432
rect 1807 1430 1808 1431
rect 1789 1428 1808 1430
rect 1703 1426 1709 1427
rect 1807 1427 1808 1428
rect 1812 1427 1813 1431
rect 1822 1428 1823 1432
rect 1827 1428 1828 1432
rect 1862 1432 1863 1436
rect 1867 1432 1868 1436
rect 2287 1435 2293 1436
rect 2287 1434 2288 1435
rect 2237 1432 2288 1434
rect 1862 1431 1868 1432
rect 2287 1431 2288 1432
rect 2292 1431 2293 1435
rect 2823 1435 2829 1436
rect 2823 1434 2824 1435
rect 2741 1432 2824 1434
rect 2287 1430 2293 1431
rect 2426 1431 2432 1432
rect 1822 1427 1828 1428
rect 2426 1427 2427 1431
rect 2431 1430 2432 1431
rect 2823 1431 2824 1432
rect 2828 1431 2829 1435
rect 2943 1435 2949 1436
rect 2943 1434 2944 1435
rect 2901 1432 2944 1434
rect 2823 1430 2829 1431
rect 2943 1431 2944 1432
rect 2948 1431 2949 1435
rect 3111 1435 3117 1436
rect 3111 1434 3112 1435
rect 3061 1432 3112 1434
rect 2943 1430 2949 1431
rect 3111 1431 3112 1432
rect 3116 1431 3117 1435
rect 3279 1435 3285 1436
rect 3279 1434 3280 1435
rect 3229 1432 3280 1434
rect 3111 1430 3117 1431
rect 3279 1431 3280 1432
rect 3284 1431 3285 1435
rect 3574 1432 3575 1436
rect 3579 1432 3580 1436
rect 3574 1431 3580 1432
rect 3279 1430 3285 1431
rect 2431 1428 2545 1430
rect 2431 1427 2432 1428
rect 1807 1426 1813 1427
rect 2426 1426 2432 1427
rect 1215 1424 1281 1426
rect 1215 1423 1216 1424
rect 1210 1422 1216 1423
rect 1862 1419 1868 1420
rect 110 1415 116 1416
rect 110 1411 111 1415
rect 115 1411 116 1415
rect 534 1415 540 1416
rect 534 1414 535 1415
rect 449 1412 535 1414
rect 110 1410 116 1411
rect 534 1411 535 1412
rect 539 1411 540 1415
rect 1822 1415 1828 1416
rect 534 1410 540 1411
rect 1444 1412 1513 1414
rect 134 1405 140 1406
rect 134 1401 135 1405
rect 139 1401 140 1405
rect 134 1400 140 1401
rect 254 1405 260 1406
rect 254 1401 255 1405
rect 259 1401 260 1405
rect 254 1400 260 1401
rect 390 1405 396 1406
rect 390 1401 391 1405
rect 395 1401 396 1405
rect 390 1400 396 1401
rect 526 1405 532 1406
rect 526 1401 527 1405
rect 531 1401 532 1405
rect 526 1400 532 1401
rect 654 1405 660 1406
rect 654 1401 655 1405
rect 659 1401 660 1405
rect 654 1400 660 1401
rect 782 1405 788 1406
rect 782 1401 783 1405
rect 787 1401 788 1405
rect 782 1400 788 1401
rect 902 1405 908 1406
rect 902 1401 903 1405
rect 907 1401 908 1405
rect 902 1400 908 1401
rect 1014 1405 1020 1406
rect 1014 1401 1015 1405
rect 1019 1401 1020 1405
rect 1014 1400 1020 1401
rect 1134 1405 1140 1406
rect 1134 1401 1135 1405
rect 1139 1401 1140 1405
rect 1134 1400 1140 1401
rect 1254 1405 1260 1406
rect 1254 1401 1255 1405
rect 1259 1401 1260 1405
rect 1254 1400 1260 1401
rect 1374 1405 1380 1406
rect 1374 1401 1375 1405
rect 1379 1401 1380 1405
rect 1374 1400 1380 1401
rect 1402 1399 1408 1400
rect 1402 1395 1403 1399
rect 1407 1398 1408 1399
rect 1444 1398 1446 1412
rect 1822 1411 1823 1415
rect 1827 1411 1828 1415
rect 1862 1415 1863 1419
rect 1867 1415 1868 1419
rect 2474 1419 2480 1420
rect 2474 1418 2475 1419
rect 2409 1416 2475 1418
rect 1862 1414 1868 1415
rect 2474 1415 2475 1416
rect 2479 1415 2480 1419
rect 2474 1414 2480 1415
rect 3258 1419 3264 1420
rect 3258 1415 3259 1419
rect 3263 1418 3264 1419
rect 3574 1419 3580 1420
rect 3263 1416 3353 1418
rect 3263 1415 3264 1416
rect 3258 1414 3264 1415
rect 3574 1415 3575 1419
rect 3579 1415 3580 1419
rect 3574 1414 3580 1415
rect 1822 1410 1828 1411
rect 2174 1409 2180 1410
rect 1494 1405 1500 1406
rect 1494 1401 1495 1405
rect 1499 1401 1500 1405
rect 1494 1400 1500 1401
rect 1622 1405 1628 1406
rect 1622 1401 1623 1405
rect 1627 1401 1628 1405
rect 1622 1400 1628 1401
rect 1726 1405 1732 1406
rect 1726 1401 1727 1405
rect 1731 1401 1732 1405
rect 2174 1405 2175 1409
rect 2179 1405 2180 1409
rect 2174 1404 2180 1405
rect 2350 1409 2356 1410
rect 2350 1405 2351 1409
rect 2355 1405 2356 1409
rect 2350 1404 2356 1405
rect 2518 1409 2524 1410
rect 2518 1405 2519 1409
rect 2523 1405 2524 1409
rect 2518 1404 2524 1405
rect 2678 1409 2684 1410
rect 2678 1405 2679 1409
rect 2683 1405 2684 1409
rect 2678 1404 2684 1405
rect 2838 1409 2844 1410
rect 2838 1405 2839 1409
rect 2843 1405 2844 1409
rect 2838 1404 2844 1405
rect 2998 1409 3004 1410
rect 2998 1405 2999 1409
rect 3003 1405 3004 1409
rect 2998 1404 3004 1405
rect 3166 1409 3172 1410
rect 3166 1405 3167 1409
rect 3171 1405 3172 1409
rect 3166 1404 3172 1405
rect 3334 1409 3340 1410
rect 3334 1405 3335 1409
rect 3339 1405 3340 1409
rect 3334 1404 3340 1405
rect 3478 1409 3484 1410
rect 3478 1405 3479 1409
rect 3483 1405 3484 1409
rect 3478 1404 3484 1405
rect 1726 1400 1732 1401
rect 3518 1403 3524 1404
rect 3518 1399 3519 1403
rect 3523 1402 3524 1403
rect 3527 1403 3533 1404
rect 3527 1402 3528 1403
rect 3523 1400 3528 1402
rect 3523 1399 3524 1400
rect 3518 1398 3524 1399
rect 3527 1399 3528 1400
rect 3532 1399 3533 1403
rect 3527 1398 3533 1399
rect 1407 1396 1446 1398
rect 1407 1395 1408 1396
rect 1402 1394 1408 1395
rect 134 1383 140 1384
rect 134 1379 135 1383
rect 139 1379 140 1383
rect 134 1378 140 1379
rect 326 1383 332 1384
rect 326 1379 327 1383
rect 331 1379 332 1383
rect 326 1378 332 1379
rect 550 1383 556 1384
rect 550 1379 551 1383
rect 555 1379 556 1383
rect 550 1378 556 1379
rect 782 1383 788 1384
rect 782 1379 783 1383
rect 787 1379 788 1383
rect 782 1378 788 1379
rect 1022 1383 1028 1384
rect 1022 1379 1023 1383
rect 1027 1379 1028 1383
rect 1022 1378 1028 1379
rect 1262 1383 1268 1384
rect 1262 1379 1263 1383
rect 1267 1379 1268 1383
rect 1262 1378 1268 1379
rect 1502 1383 1508 1384
rect 1502 1379 1503 1383
rect 1507 1379 1508 1383
rect 1502 1378 1508 1379
rect 1726 1383 1732 1384
rect 1726 1379 1727 1383
rect 1731 1379 1732 1383
rect 1726 1378 1732 1379
rect 2078 1379 2084 1380
rect 622 1375 628 1376
rect 110 1373 116 1374
rect 110 1369 111 1373
rect 115 1369 116 1373
rect 622 1371 623 1375
rect 627 1374 628 1375
rect 1591 1375 1597 1376
rect 1591 1374 1592 1375
rect 627 1372 801 1374
rect 1561 1372 1592 1374
rect 627 1371 628 1372
rect 622 1370 628 1371
rect 1591 1371 1592 1372
rect 1596 1371 1597 1375
rect 2078 1375 2079 1379
rect 2083 1375 2084 1379
rect 2078 1374 2084 1375
rect 2262 1379 2268 1380
rect 2262 1375 2263 1379
rect 2267 1375 2268 1379
rect 2262 1374 2268 1375
rect 2438 1379 2444 1380
rect 2438 1375 2439 1379
rect 2443 1375 2444 1379
rect 2438 1374 2444 1375
rect 2614 1379 2620 1380
rect 2614 1375 2615 1379
rect 2619 1375 2620 1379
rect 2614 1374 2620 1375
rect 2782 1379 2788 1380
rect 2782 1375 2783 1379
rect 2787 1375 2788 1379
rect 2782 1374 2788 1375
rect 2934 1379 2940 1380
rect 2934 1375 2935 1379
rect 2939 1375 2940 1379
rect 2934 1374 2940 1375
rect 3078 1379 3084 1380
rect 3078 1375 3079 1379
rect 3083 1375 3084 1379
rect 3078 1374 3084 1375
rect 3222 1379 3228 1380
rect 3222 1375 3223 1379
rect 3227 1375 3228 1379
rect 3222 1374 3228 1375
rect 3358 1379 3364 1380
rect 3358 1375 3359 1379
rect 3363 1375 3364 1379
rect 3358 1374 3364 1375
rect 3478 1379 3484 1380
rect 3478 1375 3479 1379
rect 3483 1375 3484 1379
rect 3478 1374 3484 1375
rect 1591 1370 1597 1371
rect 1822 1373 1828 1374
rect 110 1368 116 1369
rect 1822 1369 1823 1373
rect 1827 1369 1828 1373
rect 2538 1371 2544 1372
rect 1822 1368 1828 1369
rect 1862 1369 1868 1370
rect 1862 1365 1863 1369
rect 1867 1365 1868 1369
rect 2538 1367 2539 1371
rect 2543 1370 2544 1371
rect 3350 1371 3356 1372
rect 2543 1368 2633 1370
rect 2543 1367 2544 1368
rect 2538 1366 2544 1367
rect 3350 1367 3351 1371
rect 3355 1370 3356 1371
rect 3355 1368 3377 1370
rect 3574 1369 3580 1370
rect 3355 1367 3356 1368
rect 3350 1366 3356 1367
rect 1862 1364 1868 1365
rect 3574 1365 3575 1369
rect 3579 1365 3580 1369
rect 3574 1364 3580 1365
rect 207 1359 213 1360
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 110 1351 116 1352
rect 196 1352 198 1357
rect 207 1355 208 1359
rect 212 1358 213 1359
rect 394 1359 400 1360
rect 212 1356 353 1358
rect 212 1355 213 1356
rect 207 1354 213 1355
rect 394 1355 395 1359
rect 399 1358 400 1359
rect 850 1359 856 1360
rect 399 1356 577 1358
rect 399 1355 400 1356
rect 394 1354 400 1355
rect 850 1355 851 1359
rect 855 1358 856 1359
rect 1495 1359 1501 1360
rect 1495 1358 1496 1359
rect 855 1356 1049 1358
rect 1325 1356 1496 1358
rect 855 1355 856 1356
rect 850 1354 856 1355
rect 1495 1355 1496 1356
rect 1500 1355 1501 1359
rect 1495 1354 1501 1355
rect 1638 1359 1644 1360
rect 1638 1355 1639 1359
rect 1643 1358 1644 1359
rect 1643 1356 1753 1358
rect 1822 1356 1828 1357
rect 1643 1355 1644 1356
rect 1638 1354 1644 1355
rect 1822 1352 1823 1356
rect 1827 1352 1828 1356
rect 2255 1355 2261 1356
rect 2255 1354 2256 1355
rect 196 1351 204 1352
rect 1822 1351 1828 1352
rect 1862 1352 1868 1353
rect 2141 1352 2256 1354
rect 196 1348 199 1351
rect 198 1347 199 1348
rect 203 1347 204 1351
rect 1862 1348 1863 1352
rect 1867 1348 1868 1352
rect 2255 1351 2256 1352
rect 2260 1351 2261 1355
rect 2338 1355 2344 1356
rect 2338 1354 2339 1355
rect 2325 1352 2339 1354
rect 2255 1350 2261 1351
rect 2338 1351 2339 1352
rect 2343 1351 2344 1355
rect 2607 1355 2613 1356
rect 2607 1354 2608 1355
rect 2501 1352 2608 1354
rect 2338 1350 2344 1351
rect 2607 1351 2608 1352
rect 2612 1351 2613 1355
rect 2927 1355 2933 1356
rect 2927 1354 2928 1355
rect 2845 1352 2928 1354
rect 2607 1350 2613 1351
rect 2927 1351 2928 1352
rect 2932 1351 2933 1355
rect 3071 1355 3077 1356
rect 3071 1354 3072 1355
rect 2997 1352 3072 1354
rect 2927 1350 2933 1351
rect 3071 1351 3072 1352
rect 3076 1351 3077 1355
rect 3215 1355 3221 1356
rect 3215 1354 3216 1355
rect 3141 1352 3216 1354
rect 3071 1350 3077 1351
rect 3215 1351 3216 1352
rect 3220 1351 3221 1355
rect 3351 1355 3357 1356
rect 3351 1354 3352 1355
rect 3285 1352 3352 1354
rect 3215 1350 3221 1351
rect 3351 1351 3352 1352
rect 3356 1351 3357 1355
rect 3546 1355 3552 1356
rect 3546 1354 3547 1355
rect 3541 1352 3547 1354
rect 3351 1350 3357 1351
rect 3546 1351 3547 1352
rect 3551 1351 3552 1355
rect 3546 1350 3552 1351
rect 3574 1352 3580 1353
rect 1862 1347 1868 1348
rect 3574 1348 3575 1352
rect 3579 1348 3580 1352
rect 3574 1347 3580 1348
rect 198 1346 204 1347
rect 142 1343 148 1344
rect 142 1339 143 1343
rect 147 1339 148 1343
rect 142 1338 148 1339
rect 334 1343 340 1344
rect 334 1339 335 1343
rect 339 1339 340 1343
rect 334 1338 340 1339
rect 558 1343 564 1344
rect 558 1339 559 1343
rect 563 1339 564 1343
rect 558 1338 564 1339
rect 790 1343 796 1344
rect 790 1339 791 1343
rect 795 1339 796 1343
rect 790 1338 796 1339
rect 1030 1343 1036 1344
rect 1030 1339 1031 1343
rect 1035 1339 1036 1343
rect 1030 1338 1036 1339
rect 1270 1343 1276 1344
rect 1270 1339 1271 1343
rect 1275 1339 1276 1343
rect 1270 1338 1276 1339
rect 1510 1343 1516 1344
rect 1510 1339 1511 1343
rect 1515 1339 1516 1343
rect 1510 1338 1516 1339
rect 1734 1343 1740 1344
rect 1734 1339 1735 1343
rect 1739 1339 1740 1343
rect 1734 1338 1740 1339
rect 2086 1339 2092 1340
rect 2086 1335 2087 1339
rect 2091 1335 2092 1339
rect 2086 1334 2092 1335
rect 2270 1339 2276 1340
rect 2270 1335 2271 1339
rect 2275 1335 2276 1339
rect 2270 1334 2276 1335
rect 2446 1339 2452 1340
rect 2446 1335 2447 1339
rect 2451 1335 2452 1339
rect 2446 1334 2452 1335
rect 2622 1339 2628 1340
rect 2622 1335 2623 1339
rect 2627 1335 2628 1339
rect 2622 1334 2628 1335
rect 2790 1339 2796 1340
rect 2790 1335 2791 1339
rect 2795 1335 2796 1339
rect 2790 1334 2796 1335
rect 2942 1339 2948 1340
rect 2942 1335 2943 1339
rect 2947 1335 2948 1339
rect 2942 1334 2948 1335
rect 3086 1339 3092 1340
rect 3086 1335 3087 1339
rect 3091 1335 3092 1339
rect 3086 1334 3092 1335
rect 3230 1339 3236 1340
rect 3230 1335 3231 1339
rect 3235 1335 3236 1339
rect 3230 1334 3236 1335
rect 3366 1339 3372 1340
rect 3366 1335 3367 1339
rect 3371 1335 3372 1339
rect 3366 1334 3372 1335
rect 3486 1339 3492 1340
rect 3486 1335 3487 1339
rect 3491 1335 3492 1339
rect 3486 1334 3492 1335
rect 171 1331 177 1332
rect 171 1327 172 1331
rect 176 1330 177 1331
rect 207 1331 213 1332
rect 207 1330 208 1331
rect 176 1328 208 1330
rect 176 1327 177 1328
rect 171 1326 177 1327
rect 207 1327 208 1328
rect 212 1327 213 1331
rect 207 1326 213 1327
rect 363 1331 369 1332
rect 363 1327 364 1331
rect 368 1330 369 1331
rect 394 1331 400 1332
rect 394 1330 395 1331
rect 368 1328 395 1330
rect 368 1327 369 1328
rect 363 1326 369 1327
rect 394 1327 395 1328
rect 399 1327 400 1331
rect 394 1326 400 1327
rect 534 1331 540 1332
rect 534 1327 535 1331
rect 539 1330 540 1331
rect 587 1331 593 1332
rect 587 1330 588 1331
rect 539 1328 588 1330
rect 539 1327 540 1328
rect 534 1326 540 1327
rect 587 1327 588 1328
rect 592 1327 593 1331
rect 587 1326 593 1327
rect 819 1331 825 1332
rect 819 1327 820 1331
rect 824 1330 825 1331
rect 850 1331 856 1332
rect 850 1330 851 1331
rect 824 1328 851 1330
rect 824 1327 825 1328
rect 819 1326 825 1327
rect 850 1327 851 1328
rect 855 1327 856 1331
rect 850 1326 856 1327
rect 983 1331 989 1332
rect 983 1327 984 1331
rect 988 1330 989 1331
rect 1059 1331 1065 1332
rect 1059 1330 1060 1331
rect 988 1328 1060 1330
rect 988 1327 989 1328
rect 983 1326 989 1327
rect 1059 1327 1060 1328
rect 1064 1327 1065 1331
rect 1059 1326 1065 1327
rect 1299 1331 1308 1332
rect 1299 1327 1300 1331
rect 1307 1327 1308 1331
rect 1299 1326 1308 1327
rect 1495 1331 1501 1332
rect 1495 1327 1496 1331
rect 1500 1330 1501 1331
rect 1539 1331 1545 1332
rect 1539 1330 1540 1331
rect 1500 1328 1540 1330
rect 1500 1327 1501 1328
rect 1495 1326 1501 1327
rect 1539 1327 1540 1328
rect 1544 1327 1545 1331
rect 1539 1326 1545 1327
rect 1751 1331 1757 1332
rect 1751 1327 1752 1331
rect 1756 1330 1757 1331
rect 1763 1331 1769 1332
rect 1763 1330 1764 1331
rect 1756 1328 1764 1330
rect 1756 1327 1757 1328
rect 1751 1326 1757 1327
rect 1763 1327 1764 1328
rect 1768 1327 1769 1331
rect 1763 1326 1769 1327
rect 2115 1327 2124 1328
rect 2115 1323 2116 1327
rect 2123 1323 2124 1327
rect 2115 1322 2124 1323
rect 2255 1327 2261 1328
rect 2255 1323 2256 1327
rect 2260 1326 2261 1327
rect 2299 1327 2305 1328
rect 2299 1326 2300 1327
rect 2260 1324 2300 1326
rect 2260 1323 2261 1324
rect 2255 1322 2261 1323
rect 2299 1323 2300 1324
rect 2304 1323 2305 1327
rect 2299 1322 2305 1323
rect 2474 1327 2481 1328
rect 2474 1323 2475 1327
rect 2480 1323 2481 1327
rect 2474 1322 2481 1323
rect 2607 1327 2613 1328
rect 2607 1323 2608 1327
rect 2612 1326 2613 1327
rect 2651 1327 2657 1328
rect 2651 1326 2652 1327
rect 2612 1324 2652 1326
rect 2612 1323 2613 1324
rect 2607 1322 2613 1323
rect 2651 1323 2652 1324
rect 2656 1323 2657 1327
rect 2651 1322 2657 1323
rect 2819 1327 2828 1328
rect 2819 1323 2820 1327
rect 2827 1323 2828 1327
rect 2819 1322 2828 1323
rect 2927 1327 2933 1328
rect 2927 1323 2928 1327
rect 2932 1326 2933 1327
rect 2971 1327 2977 1328
rect 2971 1326 2972 1327
rect 2932 1324 2972 1326
rect 2932 1323 2933 1324
rect 2927 1322 2933 1323
rect 2971 1323 2972 1324
rect 2976 1323 2977 1327
rect 2971 1322 2977 1323
rect 3071 1327 3077 1328
rect 3071 1323 3072 1327
rect 3076 1326 3077 1327
rect 3115 1327 3121 1328
rect 3115 1326 3116 1327
rect 3076 1324 3116 1326
rect 3076 1323 3077 1324
rect 3071 1322 3077 1323
rect 3115 1323 3116 1324
rect 3120 1323 3121 1327
rect 3115 1322 3121 1323
rect 3215 1327 3221 1328
rect 3215 1323 3216 1327
rect 3220 1326 3221 1327
rect 3259 1327 3265 1328
rect 3259 1326 3260 1327
rect 3220 1324 3260 1326
rect 3220 1323 3221 1324
rect 3215 1322 3221 1323
rect 3259 1323 3260 1324
rect 3264 1323 3265 1327
rect 3259 1322 3265 1323
rect 3395 1327 3401 1328
rect 3395 1323 3396 1327
rect 3400 1326 3401 1327
rect 3418 1327 3424 1328
rect 3418 1326 3419 1327
rect 3400 1324 3419 1326
rect 3400 1323 3401 1324
rect 3395 1322 3401 1323
rect 3418 1323 3419 1324
rect 3423 1323 3424 1327
rect 3418 1322 3424 1323
rect 3515 1327 3524 1328
rect 3515 1323 3516 1327
rect 3523 1323 3524 1327
rect 3515 1322 3524 1323
rect 1458 1319 1464 1320
rect 1458 1318 1459 1319
rect 1100 1316 1459 1318
rect 1100 1314 1102 1316
rect 1458 1315 1459 1316
rect 1463 1315 1464 1319
rect 1458 1314 1464 1315
rect 2115 1315 2121 1316
rect 1099 1313 1105 1314
rect 171 1311 177 1312
rect 171 1307 172 1311
rect 176 1310 177 1311
rect 198 1311 204 1312
rect 198 1310 199 1311
rect 176 1308 199 1310
rect 176 1307 177 1308
rect 171 1306 177 1307
rect 198 1307 199 1308
rect 203 1307 204 1311
rect 198 1306 204 1307
rect 207 1311 213 1312
rect 207 1307 208 1311
rect 212 1310 213 1311
rect 355 1311 361 1312
rect 355 1310 356 1311
rect 212 1308 356 1310
rect 212 1307 213 1308
rect 207 1306 213 1307
rect 355 1307 356 1308
rect 360 1307 361 1311
rect 355 1306 361 1307
rect 555 1311 561 1312
rect 555 1307 556 1311
rect 560 1310 561 1311
rect 614 1311 620 1312
rect 614 1310 615 1311
rect 560 1308 615 1310
rect 560 1307 561 1308
rect 555 1306 561 1307
rect 614 1307 615 1308
rect 619 1307 620 1311
rect 614 1306 620 1307
rect 639 1311 645 1312
rect 639 1307 640 1311
rect 644 1310 645 1311
rect 747 1311 753 1312
rect 747 1310 748 1311
rect 644 1308 748 1310
rect 644 1307 645 1308
rect 639 1306 645 1307
rect 747 1307 748 1308
rect 752 1307 753 1311
rect 747 1306 753 1307
rect 831 1311 837 1312
rect 831 1307 832 1311
rect 836 1310 837 1311
rect 931 1311 937 1312
rect 931 1310 932 1311
rect 836 1308 932 1310
rect 836 1307 837 1308
rect 831 1306 837 1307
rect 931 1307 932 1308
rect 936 1307 937 1311
rect 1099 1309 1100 1313
rect 1104 1309 1105 1313
rect 1099 1308 1105 1309
rect 1214 1311 1220 1312
rect 931 1306 937 1307
rect 1214 1307 1215 1311
rect 1219 1310 1220 1311
rect 1259 1311 1265 1312
rect 1259 1310 1260 1311
rect 1219 1308 1260 1310
rect 1219 1307 1220 1308
rect 1214 1306 1220 1307
rect 1259 1307 1260 1308
rect 1264 1307 1265 1311
rect 1259 1306 1265 1307
rect 1327 1311 1333 1312
rect 1327 1307 1328 1311
rect 1332 1310 1333 1311
rect 1411 1311 1417 1312
rect 1411 1310 1412 1311
rect 1332 1308 1412 1310
rect 1332 1307 1333 1308
rect 1327 1306 1333 1307
rect 1411 1307 1412 1308
rect 1416 1307 1417 1311
rect 1411 1306 1417 1307
rect 1479 1311 1485 1312
rect 1479 1307 1480 1311
rect 1484 1310 1485 1311
rect 1563 1311 1569 1312
rect 1563 1310 1564 1311
rect 1484 1308 1564 1310
rect 1484 1307 1485 1308
rect 1479 1306 1485 1307
rect 1563 1307 1564 1308
rect 1568 1307 1569 1311
rect 1563 1306 1569 1307
rect 1631 1311 1637 1312
rect 1631 1307 1632 1311
rect 1636 1310 1637 1311
rect 1715 1311 1721 1312
rect 1715 1310 1716 1311
rect 1636 1308 1716 1310
rect 1636 1307 1637 1308
rect 1631 1306 1637 1307
rect 1715 1307 1716 1308
rect 1720 1307 1721 1311
rect 2115 1311 2116 1315
rect 2120 1314 2121 1315
rect 2294 1315 2300 1316
rect 2294 1314 2295 1315
rect 2120 1312 2295 1314
rect 2120 1311 2121 1312
rect 2115 1310 2121 1311
rect 2294 1311 2295 1312
rect 2299 1311 2300 1315
rect 2294 1310 2300 1311
rect 2338 1315 2345 1316
rect 2338 1311 2339 1315
rect 2344 1311 2345 1315
rect 2338 1310 2345 1311
rect 2431 1315 2437 1316
rect 2431 1311 2432 1315
rect 2436 1314 2437 1315
rect 2547 1315 2553 1316
rect 2547 1314 2548 1315
rect 2436 1312 2548 1314
rect 2436 1311 2437 1312
rect 2431 1310 2437 1311
rect 2547 1311 2548 1312
rect 2552 1311 2553 1315
rect 2547 1310 2553 1311
rect 2739 1315 2745 1316
rect 2739 1311 2740 1315
rect 2744 1314 2745 1315
rect 2762 1315 2768 1316
rect 2762 1314 2763 1315
rect 2744 1312 2763 1314
rect 2744 1311 2745 1312
rect 2739 1310 2745 1311
rect 2762 1311 2763 1312
rect 2767 1311 2768 1315
rect 2762 1310 2768 1311
rect 2815 1315 2821 1316
rect 2815 1311 2816 1315
rect 2820 1314 2821 1315
rect 2915 1315 2921 1316
rect 2915 1314 2916 1315
rect 2820 1312 2916 1314
rect 2820 1311 2821 1312
rect 2815 1310 2821 1311
rect 2915 1311 2916 1312
rect 2920 1311 2921 1315
rect 2915 1310 2921 1311
rect 3075 1315 3081 1316
rect 3075 1311 3076 1315
rect 3080 1314 3081 1315
rect 3114 1315 3120 1316
rect 3114 1314 3115 1315
rect 3080 1312 3115 1314
rect 3080 1311 3081 1312
rect 3075 1310 3081 1311
rect 3114 1311 3115 1312
rect 3119 1311 3120 1315
rect 3114 1310 3120 1311
rect 3227 1315 3233 1316
rect 3227 1311 3228 1315
rect 3232 1314 3233 1315
rect 3287 1315 3293 1316
rect 3287 1314 3288 1315
rect 3232 1312 3288 1314
rect 3232 1311 3233 1312
rect 3227 1310 3233 1311
rect 3287 1311 3288 1312
rect 3292 1311 3293 1315
rect 3287 1310 3293 1311
rect 3351 1315 3357 1316
rect 3351 1311 3352 1315
rect 3356 1314 3357 1315
rect 3379 1315 3385 1316
rect 3379 1314 3380 1315
rect 3356 1312 3380 1314
rect 3356 1311 3357 1312
rect 3351 1310 3357 1311
rect 3379 1311 3380 1312
rect 3384 1311 3385 1315
rect 3379 1310 3385 1311
rect 3515 1315 3521 1316
rect 3515 1311 3516 1315
rect 3520 1314 3521 1315
rect 3546 1315 3552 1316
rect 3546 1314 3547 1315
rect 3520 1312 3547 1314
rect 3520 1311 3521 1312
rect 3515 1310 3521 1311
rect 3546 1311 3547 1312
rect 3551 1311 3552 1315
rect 3546 1310 3552 1311
rect 1715 1306 1721 1307
rect 2086 1305 2092 1306
rect 142 1301 148 1302
rect 142 1297 143 1301
rect 147 1297 148 1301
rect 142 1296 148 1297
rect 326 1301 332 1302
rect 326 1297 327 1301
rect 331 1297 332 1301
rect 326 1296 332 1297
rect 526 1301 532 1302
rect 526 1297 527 1301
rect 531 1297 532 1301
rect 526 1296 532 1297
rect 718 1301 724 1302
rect 718 1297 719 1301
rect 723 1297 724 1301
rect 718 1296 724 1297
rect 902 1301 908 1302
rect 902 1297 903 1301
rect 907 1297 908 1301
rect 902 1296 908 1297
rect 1070 1301 1076 1302
rect 1070 1297 1071 1301
rect 1075 1297 1076 1301
rect 1070 1296 1076 1297
rect 1230 1301 1236 1302
rect 1230 1297 1231 1301
rect 1235 1297 1236 1301
rect 1230 1296 1236 1297
rect 1382 1301 1388 1302
rect 1382 1297 1383 1301
rect 1387 1297 1388 1301
rect 1382 1296 1388 1297
rect 1534 1301 1540 1302
rect 1534 1297 1535 1301
rect 1539 1297 1540 1301
rect 1534 1296 1540 1297
rect 1686 1301 1692 1302
rect 1686 1297 1687 1301
rect 1691 1297 1692 1301
rect 2086 1301 2087 1305
rect 2091 1301 2092 1305
rect 2086 1300 2092 1301
rect 2310 1305 2316 1306
rect 2310 1301 2311 1305
rect 2315 1301 2316 1305
rect 2310 1300 2316 1301
rect 2518 1305 2524 1306
rect 2518 1301 2519 1305
rect 2523 1301 2524 1305
rect 2518 1300 2524 1301
rect 2710 1305 2716 1306
rect 2710 1301 2711 1305
rect 2715 1301 2716 1305
rect 2710 1300 2716 1301
rect 2886 1305 2892 1306
rect 2886 1301 2887 1305
rect 2891 1301 2892 1305
rect 2886 1300 2892 1301
rect 3046 1305 3052 1306
rect 3046 1301 3047 1305
rect 3051 1301 3052 1305
rect 3046 1300 3052 1301
rect 3198 1305 3204 1306
rect 3198 1301 3199 1305
rect 3203 1301 3204 1305
rect 3198 1300 3204 1301
rect 3350 1305 3356 1306
rect 3350 1301 3351 1305
rect 3355 1301 3356 1305
rect 3350 1300 3356 1301
rect 3486 1305 3492 1306
rect 3486 1301 3487 1305
rect 3491 1301 3492 1305
rect 3486 1300 3492 1301
rect 1686 1296 1692 1297
rect 1862 1292 1868 1293
rect 3574 1292 3580 1293
rect 110 1288 116 1289
rect 1822 1288 1828 1289
rect 110 1284 111 1288
rect 115 1284 116 1288
rect 207 1287 213 1288
rect 207 1286 208 1287
rect 197 1284 208 1286
rect 110 1283 116 1284
rect 207 1283 208 1284
rect 212 1283 213 1287
rect 639 1287 645 1288
rect 639 1286 640 1287
rect 581 1284 640 1286
rect 207 1282 213 1283
rect 639 1283 640 1284
rect 644 1283 645 1287
rect 831 1287 837 1288
rect 831 1286 832 1287
rect 773 1284 832 1286
rect 639 1282 645 1283
rect 831 1283 832 1284
rect 836 1283 837 1287
rect 983 1287 989 1288
rect 983 1286 984 1287
rect 957 1284 984 1286
rect 831 1282 837 1283
rect 983 1283 984 1284
rect 988 1283 989 1287
rect 1214 1287 1220 1288
rect 1214 1286 1215 1287
rect 1125 1284 1215 1286
rect 983 1282 989 1283
rect 1214 1283 1215 1284
rect 1219 1283 1220 1287
rect 1327 1287 1333 1288
rect 1327 1286 1328 1287
rect 1285 1284 1328 1286
rect 1214 1282 1220 1283
rect 1327 1283 1328 1284
rect 1332 1283 1333 1287
rect 1479 1287 1485 1288
rect 1479 1286 1480 1287
rect 1437 1284 1480 1286
rect 1327 1282 1333 1283
rect 1479 1283 1480 1284
rect 1484 1283 1485 1287
rect 1631 1287 1637 1288
rect 1631 1286 1632 1287
rect 1589 1284 1632 1286
rect 1479 1282 1485 1283
rect 1631 1283 1632 1284
rect 1636 1283 1637 1287
rect 1751 1287 1757 1288
rect 1751 1286 1752 1287
rect 1741 1284 1752 1286
rect 1631 1282 1637 1283
rect 1751 1283 1752 1284
rect 1756 1283 1757 1287
rect 1822 1284 1823 1288
rect 1827 1284 1828 1288
rect 1862 1288 1863 1292
rect 1867 1288 1868 1292
rect 2431 1291 2437 1292
rect 2431 1290 2432 1291
rect 2365 1288 2432 1290
rect 1862 1287 1868 1288
rect 2431 1287 2432 1288
rect 2436 1287 2437 1291
rect 2815 1291 2821 1292
rect 2815 1290 2816 1291
rect 2765 1288 2816 1290
rect 2431 1286 2437 1287
rect 2442 1287 2448 1288
rect 1822 1283 1828 1284
rect 2442 1283 2443 1287
rect 2447 1286 2448 1287
rect 2815 1287 2816 1288
rect 2820 1287 2821 1291
rect 3574 1288 3575 1292
rect 3579 1288 3580 1292
rect 2815 1286 2821 1287
rect 3114 1287 3120 1288
rect 2447 1284 2537 1286
rect 2447 1283 2448 1284
rect 1751 1282 1757 1283
rect 2442 1282 2448 1283
rect 3114 1283 3115 1287
rect 3119 1286 3120 1287
rect 3287 1287 3293 1288
rect 3574 1287 3580 1288
rect 3119 1284 3217 1286
rect 3119 1283 3120 1284
rect 3114 1282 3120 1283
rect 3287 1283 3288 1287
rect 3292 1286 3293 1287
rect 3292 1284 3369 1286
rect 3292 1283 3293 1284
rect 3287 1282 3293 1283
rect 1862 1275 1868 1276
rect 110 1271 116 1272
rect 110 1267 111 1271
rect 115 1267 116 1271
rect 110 1266 116 1267
rect 210 1271 216 1272
rect 210 1267 211 1271
rect 215 1270 216 1271
rect 1822 1271 1828 1272
rect 215 1268 337 1270
rect 215 1267 216 1268
rect 210 1266 216 1267
rect 1822 1267 1823 1271
rect 1827 1267 1828 1271
rect 1862 1271 1863 1275
rect 1867 1271 1868 1275
rect 1862 1270 1868 1271
rect 2958 1275 2964 1276
rect 2958 1271 2959 1275
rect 2963 1274 2964 1275
rect 3574 1275 3580 1276
rect 2963 1272 3057 1274
rect 2963 1271 2964 1272
rect 2958 1270 2964 1271
rect 3574 1271 3575 1275
rect 3579 1271 3580 1275
rect 3574 1270 3580 1271
rect 1822 1266 1828 1267
rect 2078 1265 2084 1266
rect 134 1261 140 1262
rect 134 1257 135 1261
rect 139 1257 140 1261
rect 134 1256 140 1257
rect 318 1261 324 1262
rect 318 1257 319 1261
rect 323 1257 324 1261
rect 318 1256 324 1257
rect 518 1261 524 1262
rect 518 1257 519 1261
rect 523 1257 524 1261
rect 518 1256 524 1257
rect 710 1261 716 1262
rect 710 1257 711 1261
rect 715 1257 716 1261
rect 710 1256 716 1257
rect 894 1261 900 1262
rect 894 1257 895 1261
rect 899 1257 900 1261
rect 894 1256 900 1257
rect 1062 1261 1068 1262
rect 1062 1257 1063 1261
rect 1067 1257 1068 1261
rect 1062 1256 1068 1257
rect 1222 1261 1228 1262
rect 1222 1257 1223 1261
rect 1227 1257 1228 1261
rect 1222 1256 1228 1257
rect 1374 1261 1380 1262
rect 1374 1257 1375 1261
rect 1379 1257 1380 1261
rect 1374 1256 1380 1257
rect 1526 1261 1532 1262
rect 1526 1257 1527 1261
rect 1531 1257 1532 1261
rect 1526 1256 1532 1257
rect 1678 1261 1684 1262
rect 1678 1257 1679 1261
rect 1683 1257 1684 1261
rect 2078 1261 2079 1265
rect 2083 1261 2084 1265
rect 2078 1260 2084 1261
rect 2302 1265 2308 1266
rect 2302 1261 2303 1265
rect 2307 1261 2308 1265
rect 2302 1260 2308 1261
rect 2510 1265 2516 1266
rect 2510 1261 2511 1265
rect 2515 1261 2516 1265
rect 2510 1260 2516 1261
rect 2702 1265 2708 1266
rect 2702 1261 2703 1265
rect 2707 1261 2708 1265
rect 2702 1260 2708 1261
rect 2878 1265 2884 1266
rect 2878 1261 2879 1265
rect 2883 1261 2884 1265
rect 2878 1260 2884 1261
rect 3038 1265 3044 1266
rect 3038 1261 3039 1265
rect 3043 1261 3044 1265
rect 3038 1260 3044 1261
rect 3190 1265 3196 1266
rect 3190 1261 3191 1265
rect 3195 1261 3196 1265
rect 3190 1260 3196 1261
rect 3342 1265 3348 1266
rect 3342 1261 3343 1265
rect 3347 1261 3348 1265
rect 3342 1260 3348 1261
rect 3478 1265 3484 1266
rect 3478 1261 3479 1265
rect 3483 1261 3484 1265
rect 3478 1260 3484 1261
rect 1678 1256 1684 1257
rect 2127 1259 2136 1260
rect 2127 1255 2128 1259
rect 2135 1255 2136 1259
rect 2127 1254 2136 1255
rect 2927 1259 2933 1260
rect 2927 1255 2928 1259
rect 2932 1258 2933 1259
rect 2950 1259 2956 1260
rect 2950 1258 2951 1259
rect 2932 1256 2951 1258
rect 2932 1255 2933 1256
rect 2927 1254 2933 1255
rect 2950 1255 2951 1256
rect 2955 1255 2956 1259
rect 2950 1254 2956 1255
rect 3518 1259 3524 1260
rect 3518 1255 3519 1259
rect 3523 1258 3524 1259
rect 3527 1259 3533 1260
rect 3527 1258 3528 1259
rect 3523 1256 3528 1258
rect 3523 1255 3524 1256
rect 3518 1254 3524 1255
rect 3527 1255 3528 1256
rect 3532 1255 3533 1259
rect 3527 1254 3533 1255
rect 2762 1251 2768 1252
rect 2762 1247 2763 1251
rect 2767 1250 2768 1251
rect 2958 1251 2964 1252
rect 2958 1250 2959 1251
rect 2767 1248 2959 1250
rect 2767 1247 2768 1248
rect 2762 1246 2768 1247
rect 2958 1247 2959 1248
rect 2963 1247 2964 1251
rect 2958 1246 2964 1247
rect 1902 1239 1908 1240
rect 134 1235 140 1236
rect 134 1231 135 1235
rect 139 1231 140 1235
rect 134 1230 140 1231
rect 294 1235 300 1236
rect 294 1231 295 1235
rect 299 1231 300 1235
rect 294 1230 300 1231
rect 478 1235 484 1236
rect 478 1231 479 1235
rect 483 1231 484 1235
rect 478 1230 484 1231
rect 654 1235 660 1236
rect 654 1231 655 1235
rect 659 1231 660 1235
rect 654 1230 660 1231
rect 814 1235 820 1236
rect 814 1231 815 1235
rect 819 1231 820 1235
rect 814 1230 820 1231
rect 966 1235 972 1236
rect 966 1231 967 1235
rect 971 1231 972 1235
rect 966 1230 972 1231
rect 1110 1235 1116 1236
rect 1110 1231 1111 1235
rect 1115 1231 1116 1235
rect 1110 1230 1116 1231
rect 1246 1235 1252 1236
rect 1246 1231 1247 1235
rect 1251 1231 1252 1235
rect 1246 1230 1252 1231
rect 1382 1235 1388 1236
rect 1382 1231 1383 1235
rect 1387 1231 1388 1235
rect 1382 1230 1388 1231
rect 1526 1235 1532 1236
rect 1526 1231 1527 1235
rect 1531 1231 1532 1235
rect 1902 1235 1903 1239
rect 1907 1235 1908 1239
rect 1902 1234 1908 1235
rect 1990 1239 1996 1240
rect 1990 1235 1991 1239
rect 1995 1235 1996 1239
rect 1990 1234 1996 1235
rect 2094 1239 2100 1240
rect 2094 1235 2095 1239
rect 2099 1235 2100 1239
rect 2094 1234 2100 1235
rect 2214 1239 2220 1240
rect 2214 1235 2215 1239
rect 2219 1235 2220 1239
rect 2214 1234 2220 1235
rect 2350 1239 2356 1240
rect 2350 1235 2351 1239
rect 2355 1235 2356 1239
rect 2350 1234 2356 1235
rect 2486 1239 2492 1240
rect 2486 1235 2487 1239
rect 2491 1235 2492 1239
rect 2486 1234 2492 1235
rect 2630 1239 2636 1240
rect 2630 1235 2631 1239
rect 2635 1235 2636 1239
rect 2630 1234 2636 1235
rect 2774 1239 2780 1240
rect 2774 1235 2775 1239
rect 2779 1235 2780 1239
rect 2774 1234 2780 1235
rect 2918 1239 2924 1240
rect 2918 1235 2919 1239
rect 2923 1235 2924 1239
rect 2918 1234 2924 1235
rect 3062 1239 3068 1240
rect 3062 1235 3063 1239
rect 3067 1235 3068 1239
rect 3062 1234 3068 1235
rect 3206 1239 3212 1240
rect 3206 1235 3207 1239
rect 3211 1235 3212 1239
rect 3206 1234 3212 1235
rect 3350 1239 3356 1240
rect 3350 1235 3351 1239
rect 3355 1235 3356 1239
rect 3350 1234 3356 1235
rect 3478 1239 3484 1240
rect 3478 1235 3479 1239
rect 3483 1235 3484 1239
rect 3478 1234 3484 1235
rect 1526 1230 1532 1231
rect 2554 1231 2560 1232
rect 1862 1229 1868 1230
rect 614 1227 620 1228
rect 110 1225 116 1226
rect 110 1221 111 1225
rect 115 1221 116 1225
rect 614 1223 615 1227
rect 619 1226 620 1227
rect 1458 1227 1464 1228
rect 619 1224 673 1226
rect 619 1223 620 1224
rect 614 1222 620 1223
rect 1458 1223 1459 1227
rect 1463 1226 1464 1227
rect 1463 1224 1545 1226
rect 1822 1225 1828 1226
rect 1463 1223 1464 1224
rect 1458 1222 1464 1223
rect 110 1220 116 1221
rect 1822 1221 1823 1225
rect 1827 1221 1828 1225
rect 1862 1225 1863 1229
rect 1867 1225 1868 1229
rect 2554 1227 2555 1231
rect 2559 1230 2560 1231
rect 3138 1231 3144 1232
rect 2559 1228 2649 1230
rect 2559 1227 2560 1228
rect 2554 1226 2560 1227
rect 3138 1227 3139 1231
rect 3143 1230 3144 1231
rect 3418 1231 3424 1232
rect 3418 1230 3419 1231
rect 3143 1228 3225 1230
rect 3409 1228 3419 1230
rect 3143 1227 3144 1228
rect 3138 1226 3144 1227
rect 3418 1227 3419 1228
rect 3423 1227 3424 1231
rect 3418 1226 3424 1227
rect 3574 1229 3580 1230
rect 1862 1224 1868 1225
rect 3574 1225 3575 1229
rect 3579 1225 3580 1229
rect 3574 1224 3580 1225
rect 1822 1220 1828 1221
rect 1970 1215 1976 1216
rect 1970 1214 1971 1215
rect 1862 1212 1868 1213
rect 1965 1212 1971 1214
rect 287 1211 293 1212
rect 287 1210 288 1211
rect 110 1208 116 1209
rect 197 1208 288 1210
rect 110 1204 111 1208
rect 115 1204 116 1208
rect 287 1207 288 1208
rect 292 1207 293 1211
rect 471 1211 477 1212
rect 471 1210 472 1211
rect 357 1208 472 1210
rect 287 1206 293 1207
rect 471 1207 472 1208
rect 476 1207 477 1211
rect 546 1211 552 1212
rect 546 1210 547 1211
rect 541 1208 547 1210
rect 471 1206 477 1207
rect 546 1207 547 1208
rect 551 1207 552 1211
rect 546 1206 552 1207
rect 722 1211 728 1212
rect 722 1207 723 1211
rect 727 1210 728 1211
rect 1103 1211 1109 1212
rect 1103 1210 1104 1211
rect 727 1208 841 1210
rect 1029 1208 1104 1210
rect 727 1207 728 1208
rect 722 1206 728 1207
rect 1103 1207 1104 1208
rect 1108 1207 1109 1211
rect 1239 1211 1245 1212
rect 1239 1210 1240 1211
rect 1173 1208 1240 1210
rect 1103 1206 1109 1207
rect 1239 1207 1240 1208
rect 1244 1207 1245 1211
rect 1375 1211 1381 1212
rect 1375 1210 1376 1211
rect 1309 1208 1376 1210
rect 1239 1206 1245 1207
rect 1375 1207 1376 1208
rect 1380 1207 1381 1211
rect 1519 1211 1525 1212
rect 1519 1210 1520 1211
rect 1445 1208 1520 1210
rect 1375 1206 1381 1207
rect 1519 1207 1520 1208
rect 1524 1207 1525 1211
rect 1519 1206 1525 1207
rect 1822 1208 1828 1209
rect 110 1203 116 1204
rect 1822 1204 1823 1208
rect 1827 1204 1828 1208
rect 1862 1208 1863 1212
rect 1867 1208 1868 1212
rect 1970 1211 1971 1212
rect 1975 1211 1976 1215
rect 1970 1210 1976 1211
rect 1978 1215 1984 1216
rect 1978 1211 1979 1215
rect 1983 1214 1984 1215
rect 2086 1215 2092 1216
rect 1983 1212 2017 1214
rect 1983 1211 1984 1212
rect 1978 1210 1984 1211
rect 2086 1211 2087 1215
rect 2091 1214 2092 1215
rect 2162 1215 2168 1216
rect 2091 1212 2121 1214
rect 2091 1211 2092 1212
rect 2086 1210 2092 1211
rect 2162 1211 2163 1215
rect 2167 1214 2168 1215
rect 2282 1215 2288 1216
rect 2167 1212 2241 1214
rect 2167 1211 2168 1212
rect 2162 1210 2168 1211
rect 2282 1211 2283 1215
rect 2287 1214 2288 1215
rect 2623 1215 2629 1216
rect 2623 1214 2624 1215
rect 2287 1212 2377 1214
rect 2549 1212 2624 1214
rect 2287 1211 2288 1212
rect 2282 1210 2288 1211
rect 2623 1211 2624 1212
rect 2628 1211 2629 1215
rect 2623 1210 2629 1211
rect 2698 1215 2704 1216
rect 2698 1211 2699 1215
rect 2703 1214 2704 1215
rect 3055 1215 3061 1216
rect 3055 1214 3056 1215
rect 2703 1212 2801 1214
rect 2981 1212 3056 1214
rect 2703 1211 2704 1212
rect 2698 1210 2704 1211
rect 3055 1211 3056 1212
rect 3060 1211 3061 1215
rect 3199 1215 3205 1216
rect 3199 1214 3200 1215
rect 3125 1212 3200 1214
rect 3055 1210 3061 1211
rect 3199 1211 3200 1212
rect 3204 1211 3205 1215
rect 3546 1215 3552 1216
rect 3546 1214 3547 1215
rect 3541 1212 3547 1214
rect 3199 1210 3205 1211
rect 3546 1211 3547 1212
rect 3551 1211 3552 1215
rect 3546 1210 3552 1211
rect 3574 1212 3580 1213
rect 1862 1207 1868 1208
rect 3574 1208 3575 1212
rect 3579 1208 3580 1212
rect 3574 1207 3580 1208
rect 1822 1203 1828 1204
rect 1910 1199 1916 1200
rect 142 1195 148 1196
rect 142 1191 143 1195
rect 147 1191 148 1195
rect 142 1190 148 1191
rect 302 1195 308 1196
rect 302 1191 303 1195
rect 307 1191 308 1195
rect 302 1190 308 1191
rect 486 1195 492 1196
rect 486 1191 487 1195
rect 491 1191 492 1195
rect 486 1190 492 1191
rect 662 1195 668 1196
rect 662 1191 663 1195
rect 667 1191 668 1195
rect 662 1190 668 1191
rect 822 1195 828 1196
rect 822 1191 823 1195
rect 827 1191 828 1195
rect 822 1190 828 1191
rect 974 1195 980 1196
rect 974 1191 975 1195
rect 979 1191 980 1195
rect 974 1190 980 1191
rect 1118 1195 1124 1196
rect 1118 1191 1119 1195
rect 1123 1191 1124 1195
rect 1118 1190 1124 1191
rect 1254 1195 1260 1196
rect 1254 1191 1255 1195
rect 1259 1191 1260 1195
rect 1254 1190 1260 1191
rect 1390 1195 1396 1196
rect 1390 1191 1391 1195
rect 1395 1191 1396 1195
rect 1390 1190 1396 1191
rect 1534 1195 1540 1196
rect 1534 1191 1535 1195
rect 1539 1191 1540 1195
rect 1910 1195 1911 1199
rect 1915 1195 1916 1199
rect 1910 1194 1916 1195
rect 1998 1199 2004 1200
rect 1998 1195 1999 1199
rect 2003 1195 2004 1199
rect 1998 1194 2004 1195
rect 2102 1199 2108 1200
rect 2102 1195 2103 1199
rect 2107 1195 2108 1199
rect 2222 1199 2228 1200
rect 2102 1194 2108 1195
rect 2162 1195 2168 1196
rect 2162 1194 2163 1195
rect 1534 1190 1540 1191
rect 2112 1192 2163 1194
rect 2112 1190 2114 1192
rect 2162 1191 2163 1192
rect 2167 1191 2168 1195
rect 2222 1195 2223 1199
rect 2227 1195 2228 1199
rect 2222 1194 2228 1195
rect 2358 1199 2364 1200
rect 2358 1195 2359 1199
rect 2363 1195 2364 1199
rect 2358 1194 2364 1195
rect 2494 1199 2500 1200
rect 2494 1195 2495 1199
rect 2499 1195 2500 1199
rect 2638 1199 2644 1200
rect 2494 1194 2500 1195
rect 2554 1195 2560 1196
rect 2554 1194 2555 1195
rect 2162 1190 2168 1191
rect 2504 1192 2555 1194
rect 2504 1190 2506 1192
rect 2554 1191 2555 1192
rect 2559 1191 2560 1195
rect 2638 1195 2639 1199
rect 2643 1195 2644 1199
rect 2638 1194 2644 1195
rect 2782 1199 2788 1200
rect 2782 1195 2783 1199
rect 2787 1195 2788 1199
rect 2782 1194 2788 1195
rect 2926 1199 2932 1200
rect 2926 1195 2927 1199
rect 2931 1195 2932 1199
rect 2926 1194 2932 1195
rect 3070 1199 3076 1200
rect 3070 1195 3071 1199
rect 3075 1195 3076 1199
rect 3070 1194 3076 1195
rect 3214 1199 3220 1200
rect 3214 1195 3215 1199
rect 3219 1195 3220 1199
rect 3214 1194 3220 1195
rect 3358 1199 3364 1200
rect 3358 1195 3359 1199
rect 3363 1195 3364 1199
rect 3358 1194 3364 1195
rect 3486 1199 3492 1200
rect 3486 1195 3487 1199
rect 3491 1195 3492 1199
rect 3486 1194 3492 1195
rect 2554 1190 2560 1191
rect 2027 1189 2114 1190
rect 1939 1187 1945 1188
rect 171 1183 177 1184
rect 171 1179 172 1183
rect 176 1182 177 1183
rect 210 1183 216 1184
rect 210 1182 211 1183
rect 176 1180 211 1182
rect 176 1179 177 1180
rect 171 1178 177 1179
rect 210 1179 211 1180
rect 215 1179 216 1183
rect 210 1178 216 1179
rect 287 1183 293 1184
rect 287 1179 288 1183
rect 292 1182 293 1183
rect 331 1183 337 1184
rect 331 1182 332 1183
rect 292 1180 332 1182
rect 292 1179 293 1180
rect 287 1178 293 1179
rect 331 1179 332 1180
rect 336 1179 337 1183
rect 331 1178 337 1179
rect 471 1183 477 1184
rect 471 1179 472 1183
rect 476 1182 477 1183
rect 515 1183 521 1184
rect 515 1182 516 1183
rect 476 1180 516 1182
rect 476 1179 477 1180
rect 471 1178 477 1179
rect 515 1179 516 1180
rect 520 1179 521 1183
rect 515 1178 521 1179
rect 691 1183 697 1184
rect 691 1179 692 1183
rect 696 1182 697 1183
rect 722 1183 728 1184
rect 722 1182 723 1183
rect 696 1180 723 1182
rect 696 1179 697 1180
rect 691 1178 697 1179
rect 722 1179 723 1180
rect 727 1179 728 1183
rect 722 1178 728 1179
rect 823 1183 829 1184
rect 823 1179 824 1183
rect 828 1182 829 1183
rect 851 1183 857 1184
rect 851 1182 852 1183
rect 828 1180 852 1182
rect 828 1179 829 1180
rect 823 1178 829 1179
rect 851 1179 852 1180
rect 856 1179 857 1183
rect 851 1178 857 1179
rect 1003 1183 1009 1184
rect 1003 1179 1004 1183
rect 1008 1182 1009 1183
rect 1050 1183 1056 1184
rect 1050 1182 1051 1183
rect 1008 1180 1051 1182
rect 1008 1179 1009 1180
rect 1003 1178 1009 1179
rect 1050 1179 1051 1180
rect 1055 1179 1056 1183
rect 1050 1178 1056 1179
rect 1103 1183 1109 1184
rect 1103 1179 1104 1183
rect 1108 1182 1109 1183
rect 1147 1183 1153 1184
rect 1147 1182 1148 1183
rect 1108 1180 1148 1182
rect 1108 1179 1109 1180
rect 1103 1178 1109 1179
rect 1147 1179 1148 1180
rect 1152 1179 1153 1183
rect 1147 1178 1153 1179
rect 1239 1183 1245 1184
rect 1239 1179 1240 1183
rect 1244 1182 1245 1183
rect 1283 1183 1289 1184
rect 1283 1182 1284 1183
rect 1244 1180 1284 1182
rect 1244 1179 1245 1180
rect 1239 1178 1245 1179
rect 1283 1179 1284 1180
rect 1288 1179 1289 1183
rect 1283 1178 1289 1179
rect 1375 1183 1381 1184
rect 1375 1179 1376 1183
rect 1380 1182 1381 1183
rect 1419 1183 1425 1184
rect 1419 1182 1420 1183
rect 1380 1180 1420 1182
rect 1380 1179 1381 1180
rect 1375 1178 1381 1179
rect 1419 1179 1420 1180
rect 1424 1179 1425 1183
rect 1419 1178 1425 1179
rect 1519 1183 1525 1184
rect 1519 1179 1520 1183
rect 1524 1182 1525 1183
rect 1563 1183 1569 1184
rect 1563 1182 1564 1183
rect 1524 1180 1564 1182
rect 1524 1179 1525 1180
rect 1519 1178 1525 1179
rect 1563 1179 1564 1180
rect 1568 1179 1569 1183
rect 1939 1183 1940 1187
rect 1944 1186 1945 1187
rect 1978 1187 1984 1188
rect 1978 1186 1979 1187
rect 1944 1184 1979 1186
rect 1944 1183 1945 1184
rect 1939 1182 1945 1183
rect 1978 1183 1979 1184
rect 1983 1183 1984 1187
rect 2027 1185 2028 1189
rect 2032 1188 2114 1189
rect 2387 1189 2506 1190
rect 2032 1185 2033 1188
rect 2027 1184 2033 1185
rect 2130 1187 2137 1188
rect 1978 1182 1984 1183
rect 2130 1183 2131 1187
rect 2136 1183 2137 1187
rect 2130 1182 2137 1183
rect 2251 1187 2257 1188
rect 2251 1183 2252 1187
rect 2256 1186 2257 1187
rect 2282 1187 2288 1188
rect 2282 1186 2283 1187
rect 2256 1184 2283 1186
rect 2256 1183 2257 1184
rect 2251 1182 2257 1183
rect 2282 1183 2283 1184
rect 2287 1183 2288 1187
rect 2387 1185 2388 1189
rect 2392 1188 2506 1189
rect 2392 1185 2393 1188
rect 2387 1184 2393 1185
rect 2511 1187 2517 1188
rect 2282 1182 2288 1183
rect 2511 1183 2512 1187
rect 2516 1186 2517 1187
rect 2523 1187 2529 1188
rect 2523 1186 2524 1187
rect 2516 1184 2524 1186
rect 2516 1183 2517 1184
rect 2511 1182 2517 1183
rect 2523 1183 2524 1184
rect 2528 1183 2529 1187
rect 2523 1182 2529 1183
rect 2623 1187 2629 1188
rect 2623 1183 2624 1187
rect 2628 1186 2629 1187
rect 2667 1187 2673 1188
rect 2667 1186 2668 1187
rect 2628 1184 2668 1186
rect 2628 1183 2629 1184
rect 2623 1182 2629 1183
rect 2667 1183 2668 1184
rect 2672 1183 2673 1187
rect 2667 1182 2673 1183
rect 2811 1187 2820 1188
rect 2811 1183 2812 1187
rect 2819 1183 2820 1187
rect 2811 1182 2820 1183
rect 2950 1187 2961 1188
rect 2950 1183 2951 1187
rect 2955 1183 2956 1187
rect 2960 1183 2961 1187
rect 2950 1182 2961 1183
rect 3055 1187 3061 1188
rect 3055 1183 3056 1187
rect 3060 1186 3061 1187
rect 3099 1187 3105 1188
rect 3099 1186 3100 1187
rect 3060 1184 3100 1186
rect 3060 1183 3061 1184
rect 3055 1182 3061 1183
rect 3099 1183 3100 1184
rect 3104 1183 3105 1187
rect 3099 1182 3105 1183
rect 3199 1187 3205 1188
rect 3199 1183 3200 1187
rect 3204 1186 3205 1187
rect 3243 1187 3249 1188
rect 3243 1186 3244 1187
rect 3204 1184 3244 1186
rect 3204 1183 3205 1184
rect 3199 1182 3205 1183
rect 3243 1183 3244 1184
rect 3248 1183 3249 1187
rect 3243 1182 3249 1183
rect 3386 1187 3393 1188
rect 3386 1183 3387 1187
rect 3392 1183 3393 1187
rect 3386 1182 3393 1183
rect 3515 1187 3524 1188
rect 3515 1183 3516 1187
rect 3523 1183 3524 1187
rect 3515 1182 3524 1183
rect 1563 1178 1569 1179
rect 1923 1171 1929 1172
rect 195 1167 201 1168
rect 195 1163 196 1167
rect 200 1166 201 1167
rect 234 1167 240 1168
rect 234 1166 235 1167
rect 200 1164 235 1166
rect 200 1163 201 1164
rect 195 1162 201 1163
rect 234 1163 235 1164
rect 239 1163 240 1167
rect 234 1162 240 1163
rect 347 1167 353 1168
rect 347 1163 348 1167
rect 352 1166 353 1167
rect 390 1167 396 1168
rect 390 1166 391 1167
rect 352 1164 391 1166
rect 352 1163 353 1164
rect 347 1162 353 1163
rect 390 1163 391 1164
rect 395 1163 396 1167
rect 390 1162 396 1163
rect 499 1167 505 1168
rect 499 1163 500 1167
rect 504 1166 505 1167
rect 546 1167 552 1168
rect 546 1166 547 1167
rect 504 1164 547 1166
rect 504 1163 505 1164
rect 499 1162 505 1163
rect 546 1163 547 1164
rect 551 1163 552 1167
rect 546 1162 552 1163
rect 643 1167 652 1168
rect 643 1163 644 1167
rect 651 1163 652 1167
rect 643 1162 652 1163
rect 703 1167 709 1168
rect 703 1163 704 1167
rect 708 1166 709 1167
rect 787 1167 793 1168
rect 787 1166 788 1167
rect 708 1164 788 1166
rect 708 1163 709 1164
rect 703 1162 709 1163
rect 787 1163 788 1164
rect 792 1163 793 1167
rect 787 1162 793 1163
rect 939 1167 945 1168
rect 939 1163 940 1167
rect 944 1166 945 1167
rect 998 1167 1004 1168
rect 998 1166 999 1167
rect 944 1164 999 1166
rect 944 1163 945 1164
rect 939 1162 945 1163
rect 998 1163 999 1164
rect 1003 1163 1004 1167
rect 998 1162 1004 1163
rect 1007 1167 1013 1168
rect 1007 1163 1008 1167
rect 1012 1166 1013 1167
rect 1091 1167 1097 1168
rect 1091 1166 1092 1167
rect 1012 1164 1092 1166
rect 1012 1163 1013 1164
rect 1007 1162 1013 1163
rect 1091 1163 1092 1164
rect 1096 1163 1097 1167
rect 1091 1162 1097 1163
rect 1167 1167 1173 1168
rect 1167 1163 1168 1167
rect 1172 1166 1173 1167
rect 1259 1167 1265 1168
rect 1259 1166 1260 1167
rect 1172 1164 1260 1166
rect 1172 1163 1173 1164
rect 1167 1162 1173 1163
rect 1259 1163 1260 1164
rect 1264 1163 1265 1167
rect 1259 1162 1265 1163
rect 1335 1167 1341 1168
rect 1335 1163 1336 1167
rect 1340 1166 1341 1167
rect 1427 1167 1433 1168
rect 1427 1166 1428 1167
rect 1340 1164 1428 1166
rect 1340 1163 1341 1164
rect 1335 1162 1341 1163
rect 1427 1163 1428 1164
rect 1432 1163 1433 1167
rect 1427 1162 1433 1163
rect 1527 1167 1533 1168
rect 1527 1163 1528 1167
rect 1532 1166 1533 1167
rect 1603 1167 1609 1168
rect 1603 1166 1604 1167
rect 1532 1164 1604 1166
rect 1532 1163 1533 1164
rect 1527 1162 1533 1163
rect 1603 1163 1604 1164
rect 1608 1163 1609 1167
rect 1603 1162 1609 1163
rect 1763 1167 1769 1168
rect 1763 1163 1764 1167
rect 1768 1166 1769 1167
rect 1870 1167 1876 1168
rect 1870 1166 1871 1167
rect 1768 1164 1871 1166
rect 1768 1163 1769 1164
rect 1763 1162 1769 1163
rect 1870 1163 1871 1164
rect 1875 1163 1876 1167
rect 1923 1167 1924 1171
rect 1928 1170 1929 1171
rect 1970 1171 1976 1172
rect 1970 1170 1971 1171
rect 1928 1168 1971 1170
rect 1928 1167 1929 1168
rect 1923 1166 1929 1167
rect 1970 1167 1971 1168
rect 1975 1167 1976 1171
rect 1970 1166 1976 1167
rect 2086 1171 2097 1172
rect 2086 1167 2087 1171
rect 2091 1167 2092 1171
rect 2096 1167 2097 1171
rect 2086 1166 2097 1167
rect 2175 1171 2181 1172
rect 2175 1167 2176 1171
rect 2180 1170 2181 1171
rect 2283 1171 2289 1172
rect 2283 1170 2284 1171
rect 2180 1168 2284 1170
rect 2180 1167 2181 1168
rect 2175 1166 2181 1167
rect 2283 1167 2284 1168
rect 2288 1167 2289 1171
rect 2283 1166 2289 1167
rect 2467 1171 2473 1172
rect 2467 1167 2468 1171
rect 2472 1170 2473 1171
rect 2478 1171 2484 1172
rect 2478 1170 2479 1171
rect 2472 1168 2479 1170
rect 2472 1167 2473 1168
rect 2467 1166 2473 1167
rect 2478 1167 2479 1168
rect 2483 1167 2484 1171
rect 2478 1166 2484 1167
rect 2643 1171 2649 1172
rect 2643 1167 2644 1171
rect 2648 1170 2649 1171
rect 2698 1171 2704 1172
rect 2698 1170 2699 1171
rect 2648 1168 2699 1170
rect 2648 1167 2649 1168
rect 2643 1166 2649 1167
rect 2698 1167 2699 1168
rect 2703 1167 2704 1171
rect 2698 1166 2704 1167
rect 2719 1171 2725 1172
rect 2719 1167 2720 1171
rect 2724 1170 2725 1171
rect 2819 1171 2825 1172
rect 2819 1170 2820 1171
rect 2724 1168 2820 1170
rect 2724 1167 2725 1168
rect 2719 1166 2725 1167
rect 2819 1167 2820 1168
rect 2824 1167 2825 1171
rect 2819 1166 2825 1167
rect 2895 1171 2901 1172
rect 2895 1167 2896 1171
rect 2900 1170 2901 1171
rect 2995 1171 3001 1172
rect 2995 1170 2996 1171
rect 2900 1168 2996 1170
rect 2900 1167 2901 1168
rect 2895 1166 2901 1167
rect 2995 1167 2996 1168
rect 3000 1167 3001 1171
rect 2995 1166 3001 1167
rect 3055 1171 3061 1172
rect 3055 1167 3056 1171
rect 3060 1170 3061 1171
rect 3171 1171 3177 1172
rect 3171 1170 3172 1171
rect 3060 1168 3172 1170
rect 3060 1167 3061 1168
rect 3055 1166 3061 1167
rect 3171 1167 3172 1168
rect 3176 1167 3177 1171
rect 3355 1171 3361 1172
rect 3355 1168 3356 1171
rect 3171 1166 3177 1167
rect 3354 1167 3356 1168
rect 3360 1167 3361 1171
rect 1870 1162 1876 1163
rect 3354 1163 3355 1167
rect 3359 1166 3361 1167
rect 3515 1171 3521 1172
rect 3515 1167 3516 1171
rect 3520 1170 3521 1171
rect 3546 1171 3552 1172
rect 3546 1170 3547 1171
rect 3520 1168 3547 1170
rect 3520 1167 3521 1168
rect 3515 1166 3521 1167
rect 3546 1167 3547 1168
rect 3551 1167 3552 1171
rect 3546 1166 3552 1167
rect 3359 1163 3360 1166
rect 3354 1162 3360 1163
rect 1894 1161 1900 1162
rect 166 1157 172 1158
rect 166 1153 167 1157
rect 171 1153 172 1157
rect 166 1152 172 1153
rect 318 1157 324 1158
rect 318 1153 319 1157
rect 323 1153 324 1157
rect 318 1152 324 1153
rect 470 1157 476 1158
rect 470 1153 471 1157
rect 475 1153 476 1157
rect 470 1152 476 1153
rect 614 1157 620 1158
rect 614 1153 615 1157
rect 619 1153 620 1157
rect 614 1152 620 1153
rect 758 1157 764 1158
rect 758 1153 759 1157
rect 763 1153 764 1157
rect 758 1152 764 1153
rect 910 1157 916 1158
rect 910 1153 911 1157
rect 915 1153 916 1157
rect 910 1152 916 1153
rect 1062 1157 1068 1158
rect 1062 1153 1063 1157
rect 1067 1153 1068 1157
rect 1062 1152 1068 1153
rect 1230 1157 1236 1158
rect 1230 1153 1231 1157
rect 1235 1153 1236 1157
rect 1230 1152 1236 1153
rect 1398 1157 1404 1158
rect 1398 1153 1399 1157
rect 1403 1153 1404 1157
rect 1398 1152 1404 1153
rect 1574 1157 1580 1158
rect 1574 1153 1575 1157
rect 1579 1153 1580 1157
rect 1574 1152 1580 1153
rect 1734 1157 1740 1158
rect 1734 1153 1735 1157
rect 1739 1153 1740 1157
rect 1894 1157 1895 1161
rect 1899 1157 1900 1161
rect 1894 1156 1900 1157
rect 2062 1161 2068 1162
rect 2062 1157 2063 1161
rect 2067 1157 2068 1161
rect 2062 1156 2068 1157
rect 2254 1161 2260 1162
rect 2254 1157 2255 1161
rect 2259 1157 2260 1161
rect 2254 1156 2260 1157
rect 2438 1161 2444 1162
rect 2438 1157 2439 1161
rect 2443 1157 2444 1161
rect 2438 1156 2444 1157
rect 2614 1161 2620 1162
rect 2614 1157 2615 1161
rect 2619 1157 2620 1161
rect 2614 1156 2620 1157
rect 2790 1161 2796 1162
rect 2790 1157 2791 1161
rect 2795 1157 2796 1161
rect 2790 1156 2796 1157
rect 2966 1161 2972 1162
rect 2966 1157 2967 1161
rect 2971 1157 2972 1161
rect 2966 1156 2972 1157
rect 3142 1161 3148 1162
rect 3142 1157 3143 1161
rect 3147 1157 3148 1161
rect 3142 1156 3148 1157
rect 3326 1161 3332 1162
rect 3326 1157 3327 1161
rect 3331 1157 3332 1161
rect 3326 1156 3332 1157
rect 3486 1161 3492 1162
rect 3486 1157 3487 1161
rect 3491 1157 3492 1161
rect 3486 1156 3492 1157
rect 1734 1152 1740 1153
rect 1862 1148 1868 1149
rect 3574 1148 3580 1149
rect 110 1144 116 1145
rect 1822 1144 1828 1145
rect 110 1140 111 1144
rect 115 1140 116 1144
rect 703 1143 709 1144
rect 703 1142 704 1143
rect 669 1140 704 1142
rect 110 1139 116 1140
rect 234 1139 240 1140
rect 234 1135 235 1139
rect 239 1138 240 1139
rect 390 1139 396 1140
rect 239 1136 337 1138
rect 239 1135 240 1136
rect 234 1134 240 1135
rect 390 1135 391 1139
rect 395 1138 396 1139
rect 703 1139 704 1140
rect 708 1139 709 1143
rect 823 1143 829 1144
rect 823 1142 824 1143
rect 813 1140 824 1142
rect 703 1138 709 1139
rect 823 1139 824 1140
rect 828 1139 829 1143
rect 1007 1143 1013 1144
rect 1007 1142 1008 1143
rect 965 1140 1008 1142
rect 823 1138 829 1139
rect 1007 1139 1008 1140
rect 1012 1139 1013 1143
rect 1167 1143 1173 1144
rect 1167 1142 1168 1143
rect 1117 1140 1168 1142
rect 1007 1138 1013 1139
rect 1167 1139 1168 1140
rect 1172 1139 1173 1143
rect 1335 1143 1341 1144
rect 1335 1142 1336 1143
rect 1285 1140 1336 1142
rect 1167 1138 1173 1139
rect 1335 1139 1336 1140
rect 1340 1139 1341 1143
rect 1527 1143 1533 1144
rect 1527 1142 1528 1143
rect 1453 1140 1528 1142
rect 1335 1138 1341 1139
rect 1527 1139 1528 1140
rect 1532 1139 1533 1143
rect 1822 1140 1823 1144
rect 1827 1140 1828 1144
rect 1862 1144 1863 1148
rect 1867 1144 1868 1148
rect 2175 1147 2181 1148
rect 2175 1146 2176 1147
rect 2117 1144 2176 1146
rect 1862 1143 1868 1144
rect 1870 1143 1876 1144
rect 1527 1138 1533 1139
rect 1538 1139 1544 1140
rect 1822 1139 1828 1140
rect 1870 1139 1871 1143
rect 1875 1142 1876 1143
rect 2175 1143 2176 1144
rect 2180 1143 2181 1147
rect 2511 1147 2517 1148
rect 2511 1146 2512 1147
rect 2493 1144 2512 1146
rect 2175 1142 2181 1143
rect 2511 1143 2512 1144
rect 2516 1143 2517 1147
rect 2719 1147 2725 1148
rect 2719 1146 2720 1147
rect 2669 1144 2720 1146
rect 2511 1142 2517 1143
rect 2719 1143 2720 1144
rect 2724 1143 2725 1147
rect 2895 1147 2901 1148
rect 2895 1146 2896 1147
rect 2845 1144 2896 1146
rect 2719 1142 2725 1143
rect 2895 1143 2896 1144
rect 2900 1143 2901 1147
rect 3055 1147 3061 1148
rect 3055 1146 3056 1147
rect 3021 1144 3056 1146
rect 2895 1142 2901 1143
rect 3055 1143 3056 1144
rect 3060 1143 3061 1147
rect 3386 1147 3392 1148
rect 3386 1146 3387 1147
rect 3381 1144 3387 1146
rect 3055 1142 3061 1143
rect 3386 1143 3387 1144
rect 3391 1143 3392 1147
rect 3574 1144 3575 1148
rect 3579 1144 3580 1148
rect 3574 1143 3580 1144
rect 3386 1142 3392 1143
rect 1875 1140 1913 1142
rect 1875 1139 1876 1140
rect 395 1136 489 1138
rect 395 1135 396 1136
rect 390 1134 396 1135
rect 1538 1135 1539 1139
rect 1543 1138 1544 1139
rect 1870 1138 1876 1139
rect 1543 1136 1593 1138
rect 1543 1135 1544 1136
rect 1538 1134 1544 1135
rect 1862 1131 1868 1132
rect 110 1127 116 1128
rect 110 1123 111 1127
rect 115 1123 116 1127
rect 250 1127 256 1128
rect 250 1126 251 1127
rect 217 1124 251 1126
rect 110 1122 116 1123
rect 250 1123 251 1124
rect 255 1123 256 1127
rect 250 1122 256 1123
rect 1822 1127 1828 1128
rect 1822 1123 1823 1127
rect 1827 1123 1828 1127
rect 1862 1127 1863 1131
rect 1867 1127 1868 1131
rect 1862 1126 1868 1127
rect 2134 1131 2140 1132
rect 2134 1127 2135 1131
rect 2139 1130 2140 1131
rect 3142 1131 3148 1132
rect 2139 1128 2265 1130
rect 2139 1127 2140 1128
rect 2134 1126 2140 1127
rect 3142 1127 3143 1131
rect 3147 1130 3148 1131
rect 3574 1131 3580 1132
rect 3147 1128 3153 1130
rect 3147 1127 3148 1128
rect 3142 1126 3148 1127
rect 3574 1127 3575 1131
rect 3579 1127 3580 1131
rect 3574 1126 3580 1127
rect 1822 1122 1828 1123
rect 1886 1121 1892 1122
rect 158 1117 164 1118
rect 158 1113 159 1117
rect 163 1113 164 1117
rect 158 1112 164 1113
rect 310 1117 316 1118
rect 310 1113 311 1117
rect 315 1113 316 1117
rect 310 1112 316 1113
rect 462 1117 468 1118
rect 462 1113 463 1117
rect 467 1113 468 1117
rect 462 1112 468 1113
rect 606 1117 612 1118
rect 606 1113 607 1117
rect 611 1113 612 1117
rect 606 1112 612 1113
rect 750 1117 756 1118
rect 750 1113 751 1117
rect 755 1113 756 1117
rect 750 1112 756 1113
rect 902 1117 908 1118
rect 902 1113 903 1117
rect 907 1113 908 1117
rect 902 1112 908 1113
rect 1054 1117 1060 1118
rect 1054 1113 1055 1117
rect 1059 1113 1060 1117
rect 1054 1112 1060 1113
rect 1222 1117 1228 1118
rect 1222 1113 1223 1117
rect 1227 1113 1228 1117
rect 1222 1112 1228 1113
rect 1390 1117 1396 1118
rect 1390 1113 1391 1117
rect 1395 1113 1396 1117
rect 1390 1112 1396 1113
rect 1566 1117 1572 1118
rect 1566 1113 1567 1117
rect 1571 1113 1572 1117
rect 1566 1112 1572 1113
rect 1726 1117 1732 1118
rect 1726 1113 1727 1117
rect 1731 1113 1732 1117
rect 1886 1117 1887 1121
rect 1891 1117 1892 1121
rect 1886 1116 1892 1117
rect 2054 1121 2060 1122
rect 2054 1117 2055 1121
rect 2059 1117 2060 1121
rect 2054 1116 2060 1117
rect 2246 1121 2252 1122
rect 2246 1117 2247 1121
rect 2251 1117 2252 1121
rect 2246 1116 2252 1117
rect 2430 1121 2436 1122
rect 2430 1117 2431 1121
rect 2435 1117 2436 1121
rect 2430 1116 2436 1117
rect 2606 1121 2612 1122
rect 2606 1117 2607 1121
rect 2611 1117 2612 1121
rect 2606 1116 2612 1117
rect 2782 1121 2788 1122
rect 2782 1117 2783 1121
rect 2787 1117 2788 1121
rect 2782 1116 2788 1117
rect 2958 1121 2964 1122
rect 2958 1117 2959 1121
rect 2963 1117 2964 1121
rect 2958 1116 2964 1117
rect 3134 1121 3140 1122
rect 3134 1117 3135 1121
rect 3139 1117 3140 1121
rect 3134 1116 3140 1117
rect 3318 1121 3324 1122
rect 3318 1117 3319 1121
rect 3323 1117 3324 1121
rect 3318 1116 3324 1117
rect 3478 1121 3484 1122
rect 3478 1117 3479 1121
rect 3483 1117 3484 1121
rect 3478 1116 3484 1117
rect 1726 1112 1732 1113
rect 3518 1115 3524 1116
rect 1766 1111 1772 1112
rect 1766 1107 1767 1111
rect 1771 1110 1772 1111
rect 1775 1111 1781 1112
rect 1775 1110 1776 1111
rect 1771 1108 1776 1110
rect 1771 1107 1772 1108
rect 1766 1106 1772 1107
rect 1775 1107 1776 1108
rect 1780 1107 1781 1111
rect 3518 1111 3519 1115
rect 3523 1114 3524 1115
rect 3527 1115 3533 1116
rect 3527 1114 3528 1115
rect 3523 1112 3528 1114
rect 3523 1111 3524 1112
rect 3518 1110 3524 1111
rect 3527 1111 3528 1112
rect 3532 1111 3533 1115
rect 3527 1110 3533 1111
rect 1775 1106 1781 1107
rect 214 1091 220 1092
rect 214 1087 215 1091
rect 219 1087 220 1091
rect 214 1086 220 1087
rect 326 1091 332 1092
rect 326 1087 327 1091
rect 331 1087 332 1091
rect 326 1086 332 1087
rect 438 1091 444 1092
rect 438 1087 439 1091
rect 443 1087 444 1091
rect 438 1086 444 1087
rect 558 1091 564 1092
rect 558 1087 559 1091
rect 563 1087 564 1091
rect 558 1086 564 1087
rect 678 1091 684 1092
rect 678 1087 679 1091
rect 683 1087 684 1091
rect 678 1086 684 1087
rect 806 1091 812 1092
rect 806 1087 807 1091
rect 811 1087 812 1091
rect 806 1086 812 1087
rect 942 1091 948 1092
rect 942 1087 943 1091
rect 947 1087 948 1091
rect 942 1086 948 1087
rect 1086 1091 1092 1092
rect 1086 1087 1087 1091
rect 1091 1087 1092 1091
rect 1086 1086 1092 1087
rect 1246 1091 1252 1092
rect 1246 1087 1247 1091
rect 1251 1087 1252 1091
rect 1246 1086 1252 1087
rect 1406 1091 1412 1092
rect 1406 1087 1407 1091
rect 1411 1087 1412 1091
rect 1406 1086 1412 1087
rect 1574 1091 1580 1092
rect 1574 1087 1575 1091
rect 1579 1087 1580 1091
rect 1574 1086 1580 1087
rect 1726 1091 1732 1092
rect 1726 1087 1727 1091
rect 1731 1087 1732 1091
rect 1726 1086 1732 1087
rect 1934 1087 1940 1088
rect 646 1083 652 1084
rect 110 1081 116 1082
rect 110 1077 111 1081
rect 115 1077 116 1081
rect 646 1079 647 1083
rect 651 1082 652 1083
rect 1338 1083 1344 1084
rect 651 1080 697 1082
rect 651 1079 652 1080
rect 646 1078 652 1079
rect 1338 1079 1339 1083
rect 1343 1082 1344 1083
rect 1934 1083 1935 1087
rect 1939 1083 1940 1087
rect 1934 1082 1940 1083
rect 2094 1087 2100 1088
rect 2094 1083 2095 1087
rect 2099 1083 2100 1087
rect 2094 1082 2100 1083
rect 2246 1087 2252 1088
rect 2246 1083 2247 1087
rect 2251 1083 2252 1087
rect 2246 1082 2252 1083
rect 2406 1087 2412 1088
rect 2406 1083 2407 1087
rect 2411 1083 2412 1087
rect 2406 1082 2412 1083
rect 2566 1087 2572 1088
rect 2566 1083 2567 1087
rect 2571 1083 2572 1087
rect 2566 1082 2572 1083
rect 2734 1087 2740 1088
rect 2734 1083 2735 1087
rect 2739 1083 2740 1087
rect 2734 1082 2740 1083
rect 2910 1087 2916 1088
rect 2910 1083 2911 1087
rect 2915 1083 2916 1087
rect 2910 1082 2916 1083
rect 3094 1087 3100 1088
rect 3094 1083 3095 1087
rect 3099 1083 3100 1087
rect 3094 1082 3100 1083
rect 3286 1087 3292 1088
rect 3286 1083 3287 1087
rect 3291 1083 3292 1087
rect 3286 1082 3292 1083
rect 3478 1087 3484 1088
rect 3478 1083 3479 1087
rect 3483 1083 3484 1087
rect 3478 1082 3484 1083
rect 1343 1080 1425 1082
rect 1822 1081 1828 1082
rect 1343 1079 1344 1080
rect 1338 1078 1344 1079
rect 110 1076 116 1077
rect 1822 1077 1823 1081
rect 1827 1077 1828 1081
rect 2010 1079 2016 1080
rect 2010 1078 2011 1079
rect 1822 1076 1828 1077
rect 1862 1077 1868 1078
rect 1862 1073 1863 1077
rect 1867 1073 1868 1077
rect 1993 1076 2011 1078
rect 2010 1075 2011 1076
rect 2015 1075 2016 1079
rect 2478 1079 2484 1080
rect 2478 1078 2479 1079
rect 2465 1076 2479 1078
rect 2010 1074 2016 1075
rect 2478 1075 2479 1076
rect 2483 1075 2484 1079
rect 2642 1079 2648 1080
rect 2642 1078 2643 1079
rect 2625 1076 2643 1078
rect 2478 1074 2484 1075
rect 2642 1075 2643 1076
rect 2647 1075 2648 1079
rect 3354 1079 3360 1080
rect 3354 1078 3355 1079
rect 3345 1076 3355 1078
rect 2642 1074 2648 1075
rect 3354 1075 3355 1076
rect 3359 1075 3360 1079
rect 3354 1074 3360 1075
rect 3574 1077 3580 1078
rect 1862 1072 1868 1073
rect 3574 1073 3575 1077
rect 3579 1073 3580 1077
rect 3574 1072 3580 1073
rect 319 1067 325 1068
rect 319 1066 320 1067
rect 110 1064 116 1065
rect 277 1064 320 1066
rect 110 1060 111 1064
rect 115 1060 116 1064
rect 319 1063 320 1064
rect 324 1063 325 1067
rect 431 1067 437 1068
rect 431 1066 432 1067
rect 389 1064 432 1066
rect 319 1062 325 1063
rect 431 1063 432 1064
rect 436 1063 437 1067
rect 543 1067 549 1068
rect 543 1066 544 1067
rect 501 1064 544 1066
rect 431 1062 437 1063
rect 543 1063 544 1064
rect 548 1063 549 1067
rect 543 1062 549 1063
rect 551 1067 557 1068
rect 551 1063 552 1067
rect 556 1066 557 1067
rect 935 1067 941 1068
rect 935 1066 936 1067
rect 556 1064 585 1066
rect 869 1064 936 1066
rect 556 1063 557 1064
rect 551 1062 557 1063
rect 935 1063 936 1064
rect 940 1063 941 1067
rect 1031 1067 1037 1068
rect 1031 1066 1032 1067
rect 1005 1064 1032 1066
rect 935 1062 941 1063
rect 1031 1063 1032 1064
rect 1036 1063 1037 1067
rect 1239 1067 1245 1068
rect 1239 1066 1240 1067
rect 1149 1064 1240 1066
rect 1031 1062 1037 1063
rect 1239 1063 1240 1064
rect 1244 1063 1245 1067
rect 1399 1067 1405 1068
rect 1399 1066 1400 1067
rect 1309 1064 1400 1066
rect 1239 1062 1245 1063
rect 1399 1063 1400 1064
rect 1404 1063 1405 1067
rect 1399 1062 1405 1063
rect 1566 1067 1572 1068
rect 1566 1063 1567 1067
rect 1571 1066 1572 1067
rect 1642 1067 1648 1068
rect 1571 1064 1601 1066
rect 1571 1063 1572 1064
rect 1566 1062 1572 1063
rect 1642 1063 1643 1067
rect 1647 1066 1648 1067
rect 1647 1064 1753 1066
rect 1822 1064 1828 1065
rect 1647 1063 1648 1064
rect 1642 1062 1648 1063
rect 110 1059 116 1060
rect 1822 1060 1823 1064
rect 1827 1060 1828 1064
rect 2002 1063 2008 1064
rect 1822 1059 1828 1060
rect 1862 1060 1868 1061
rect 1862 1056 1863 1060
rect 1867 1056 1868 1060
rect 2002 1059 2003 1063
rect 2007 1062 2008 1063
rect 2399 1063 2405 1064
rect 2399 1062 2400 1063
rect 2007 1060 2121 1062
rect 2309 1060 2400 1062
rect 2007 1059 2008 1060
rect 2002 1058 2008 1059
rect 2399 1059 2400 1060
rect 2404 1059 2405 1063
rect 2399 1058 2405 1059
rect 2634 1063 2640 1064
rect 2634 1059 2635 1063
rect 2639 1062 2640 1063
rect 2855 1063 2861 1064
rect 2639 1060 2761 1062
rect 2639 1059 2640 1060
rect 2634 1058 2640 1059
rect 2855 1059 2856 1063
rect 2860 1062 2861 1063
rect 2978 1063 2984 1064
rect 2860 1060 2937 1062
rect 2860 1059 2861 1060
rect 2855 1058 2861 1059
rect 2978 1059 2979 1063
rect 2983 1062 2984 1063
rect 3546 1063 3552 1064
rect 3546 1062 3547 1063
rect 2983 1060 3121 1062
rect 3541 1060 3547 1062
rect 2983 1059 2984 1060
rect 2978 1058 2984 1059
rect 3546 1059 3547 1060
rect 3551 1059 3552 1063
rect 3546 1058 3552 1059
rect 3574 1060 3580 1061
rect 1862 1055 1868 1056
rect 3574 1056 3575 1060
rect 3579 1056 3580 1060
rect 3574 1055 3580 1056
rect 222 1051 228 1052
rect 222 1047 223 1051
rect 227 1047 228 1051
rect 222 1046 228 1047
rect 334 1051 340 1052
rect 334 1047 335 1051
rect 339 1047 340 1051
rect 334 1046 340 1047
rect 446 1051 452 1052
rect 446 1047 447 1051
rect 451 1047 452 1051
rect 446 1046 452 1047
rect 566 1051 572 1052
rect 566 1047 567 1051
rect 571 1047 572 1051
rect 566 1046 572 1047
rect 686 1051 692 1052
rect 686 1047 687 1051
rect 691 1047 692 1051
rect 686 1046 692 1047
rect 814 1051 820 1052
rect 814 1047 815 1051
rect 819 1047 820 1051
rect 814 1046 820 1047
rect 950 1051 956 1052
rect 950 1047 951 1051
rect 955 1047 956 1051
rect 950 1046 956 1047
rect 1094 1051 1100 1052
rect 1094 1047 1095 1051
rect 1099 1047 1100 1051
rect 1094 1046 1100 1047
rect 1254 1051 1260 1052
rect 1254 1047 1255 1051
rect 1259 1047 1260 1051
rect 1254 1046 1260 1047
rect 1414 1051 1420 1052
rect 1414 1047 1415 1051
rect 1419 1047 1420 1051
rect 1414 1046 1420 1047
rect 1582 1051 1588 1052
rect 1582 1047 1583 1051
rect 1587 1047 1588 1051
rect 1582 1046 1588 1047
rect 1734 1051 1740 1052
rect 1734 1047 1735 1051
rect 1739 1047 1740 1051
rect 1734 1046 1740 1047
rect 1942 1047 1948 1048
rect 1942 1043 1943 1047
rect 1947 1043 1948 1047
rect 1942 1042 1948 1043
rect 2102 1047 2108 1048
rect 2102 1043 2103 1047
rect 2107 1043 2108 1047
rect 2102 1042 2108 1043
rect 2254 1047 2260 1048
rect 2254 1043 2255 1047
rect 2259 1043 2260 1047
rect 2254 1042 2260 1043
rect 2414 1047 2420 1048
rect 2414 1043 2415 1047
rect 2419 1043 2420 1047
rect 2414 1042 2420 1043
rect 2574 1047 2580 1048
rect 2574 1043 2575 1047
rect 2579 1043 2580 1047
rect 2574 1042 2580 1043
rect 2742 1047 2748 1048
rect 2742 1043 2743 1047
rect 2747 1043 2748 1047
rect 2742 1042 2748 1043
rect 2918 1047 2924 1048
rect 2918 1043 2919 1047
rect 2923 1043 2924 1047
rect 2918 1042 2924 1043
rect 3102 1047 3108 1048
rect 3102 1043 3103 1047
rect 3107 1043 3108 1047
rect 3102 1042 3108 1043
rect 3294 1047 3300 1048
rect 3294 1043 3295 1047
rect 3299 1043 3300 1047
rect 3294 1042 3300 1043
rect 3486 1047 3492 1048
rect 3486 1043 3487 1047
rect 3491 1043 3492 1047
rect 3486 1042 3492 1043
rect 250 1039 257 1040
rect 250 1035 251 1039
rect 256 1035 257 1039
rect 250 1034 257 1035
rect 319 1039 325 1040
rect 319 1035 320 1039
rect 324 1038 325 1039
rect 363 1039 369 1040
rect 363 1038 364 1039
rect 324 1036 364 1038
rect 324 1035 325 1036
rect 319 1034 325 1035
rect 363 1035 364 1036
rect 368 1035 369 1039
rect 363 1034 369 1035
rect 431 1039 437 1040
rect 431 1035 432 1039
rect 436 1038 437 1039
rect 475 1039 481 1040
rect 475 1038 476 1039
rect 436 1036 476 1038
rect 436 1035 437 1036
rect 431 1034 437 1035
rect 475 1035 476 1036
rect 480 1035 481 1039
rect 475 1034 481 1035
rect 543 1039 549 1040
rect 543 1035 544 1039
rect 548 1038 549 1039
rect 595 1039 601 1040
rect 595 1038 596 1039
rect 548 1036 596 1038
rect 548 1035 549 1036
rect 543 1034 549 1035
rect 595 1035 596 1036
rect 600 1035 601 1039
rect 595 1034 601 1035
rect 714 1039 721 1040
rect 714 1035 715 1039
rect 720 1035 721 1039
rect 714 1034 721 1035
rect 843 1039 849 1040
rect 843 1035 844 1039
rect 848 1038 849 1039
rect 858 1039 864 1040
rect 858 1038 859 1039
rect 848 1036 859 1038
rect 848 1035 849 1036
rect 843 1034 849 1035
rect 858 1035 859 1036
rect 863 1035 864 1039
rect 858 1034 864 1035
rect 935 1039 941 1040
rect 935 1035 936 1039
rect 940 1038 941 1039
rect 979 1039 985 1040
rect 979 1038 980 1039
rect 940 1036 980 1038
rect 940 1035 941 1036
rect 935 1034 941 1035
rect 979 1035 980 1036
rect 984 1035 985 1039
rect 979 1034 985 1035
rect 1031 1039 1037 1040
rect 1031 1035 1032 1039
rect 1036 1038 1037 1039
rect 1123 1039 1129 1040
rect 1123 1038 1124 1039
rect 1036 1036 1124 1038
rect 1036 1035 1037 1036
rect 1031 1034 1037 1035
rect 1123 1035 1124 1036
rect 1128 1035 1129 1039
rect 1123 1034 1129 1035
rect 1239 1039 1245 1040
rect 1239 1035 1240 1039
rect 1244 1038 1245 1039
rect 1283 1039 1289 1040
rect 1283 1038 1284 1039
rect 1244 1036 1284 1038
rect 1244 1035 1245 1036
rect 1239 1034 1245 1035
rect 1283 1035 1284 1036
rect 1288 1035 1289 1039
rect 1283 1034 1289 1035
rect 1399 1039 1405 1040
rect 1399 1035 1400 1039
rect 1404 1038 1405 1039
rect 1443 1039 1449 1040
rect 1443 1038 1444 1039
rect 1404 1036 1444 1038
rect 1404 1035 1405 1036
rect 1399 1034 1405 1035
rect 1443 1035 1444 1036
rect 1448 1035 1449 1039
rect 1443 1034 1449 1035
rect 1611 1039 1617 1040
rect 1611 1035 1612 1039
rect 1616 1038 1617 1039
rect 1642 1039 1648 1040
rect 1642 1038 1643 1039
rect 1616 1036 1643 1038
rect 1616 1035 1617 1036
rect 1611 1034 1617 1035
rect 1642 1035 1643 1036
rect 1647 1035 1648 1039
rect 1642 1034 1648 1035
rect 1763 1039 1772 1040
rect 1763 1035 1764 1039
rect 1771 1035 1772 1039
rect 1763 1034 1772 1035
rect 1971 1035 1977 1036
rect 1971 1031 1972 1035
rect 1976 1034 1977 1035
rect 2002 1035 2008 1036
rect 2002 1034 2003 1035
rect 1976 1032 2003 1034
rect 1976 1031 1977 1032
rect 1971 1030 1977 1031
rect 2002 1031 2003 1032
rect 2007 1031 2008 1035
rect 2002 1030 2008 1031
rect 2131 1035 2140 1036
rect 2131 1031 2132 1035
rect 2139 1031 2140 1035
rect 2131 1030 2140 1031
rect 2283 1035 2289 1036
rect 2283 1031 2284 1035
rect 2288 1034 2289 1035
rect 2378 1035 2384 1036
rect 2378 1034 2379 1035
rect 2288 1032 2379 1034
rect 2288 1031 2289 1032
rect 2283 1030 2289 1031
rect 2378 1031 2379 1032
rect 2383 1031 2384 1035
rect 2378 1030 2384 1031
rect 2399 1035 2405 1036
rect 2399 1031 2400 1035
rect 2404 1034 2405 1035
rect 2443 1035 2449 1036
rect 2443 1034 2444 1035
rect 2404 1032 2444 1034
rect 2404 1031 2405 1032
rect 2399 1030 2405 1031
rect 2443 1031 2444 1032
rect 2448 1031 2449 1035
rect 2443 1030 2449 1031
rect 2603 1035 2609 1036
rect 2603 1031 2604 1035
rect 2608 1034 2609 1035
rect 2634 1035 2640 1036
rect 2634 1034 2635 1035
rect 2608 1032 2635 1034
rect 2608 1031 2609 1032
rect 2603 1030 2609 1031
rect 2634 1031 2635 1032
rect 2639 1031 2640 1035
rect 2634 1030 2640 1031
rect 2771 1035 2777 1036
rect 2771 1031 2772 1035
rect 2776 1034 2777 1035
rect 2855 1035 2861 1036
rect 2855 1034 2856 1035
rect 2776 1032 2856 1034
rect 2776 1031 2777 1032
rect 2771 1030 2777 1031
rect 2855 1031 2856 1032
rect 2860 1031 2861 1035
rect 2855 1030 2861 1031
rect 2947 1035 2953 1036
rect 2947 1031 2948 1035
rect 2952 1034 2953 1035
rect 2978 1035 2984 1036
rect 2978 1034 2979 1035
rect 2952 1032 2979 1034
rect 2952 1031 2953 1032
rect 2947 1030 2953 1031
rect 2978 1031 2979 1032
rect 2983 1031 2984 1035
rect 2978 1030 2984 1031
rect 3131 1035 3137 1036
rect 3131 1031 3132 1035
rect 3136 1034 3137 1035
rect 3142 1035 3148 1036
rect 3142 1034 3143 1035
rect 3136 1032 3143 1034
rect 3136 1031 3137 1032
rect 3131 1030 3137 1031
rect 3142 1031 3143 1032
rect 3147 1031 3148 1035
rect 3142 1030 3148 1031
rect 3263 1035 3269 1036
rect 3263 1031 3264 1035
rect 3268 1034 3269 1035
rect 3323 1035 3329 1036
rect 3323 1034 3324 1035
rect 3268 1032 3324 1034
rect 3268 1031 3269 1032
rect 3263 1030 3269 1031
rect 3323 1031 3324 1032
rect 3328 1031 3329 1035
rect 3323 1030 3329 1031
rect 3515 1035 3524 1036
rect 3515 1031 3516 1035
rect 3523 1031 3524 1035
rect 3515 1030 3524 1031
rect 371 1019 377 1020
rect 371 1015 372 1019
rect 376 1018 377 1019
rect 410 1019 416 1020
rect 410 1018 411 1019
rect 376 1016 411 1018
rect 376 1015 377 1016
rect 371 1014 377 1015
rect 410 1015 411 1016
rect 415 1015 416 1019
rect 410 1014 416 1015
rect 459 1019 465 1020
rect 459 1015 460 1019
rect 464 1018 465 1019
rect 502 1019 508 1020
rect 502 1018 503 1019
rect 464 1016 503 1018
rect 464 1015 465 1016
rect 459 1014 465 1015
rect 502 1015 503 1016
rect 507 1015 508 1019
rect 502 1014 508 1015
rect 551 1019 557 1020
rect 551 1015 552 1019
rect 556 1018 557 1019
rect 563 1019 569 1020
rect 563 1018 564 1019
rect 556 1016 564 1018
rect 556 1015 557 1016
rect 551 1014 557 1015
rect 563 1015 564 1016
rect 568 1015 569 1019
rect 563 1014 569 1015
rect 683 1019 689 1020
rect 683 1015 684 1019
rect 688 1018 689 1019
rect 722 1019 728 1020
rect 722 1018 723 1019
rect 688 1016 723 1018
rect 688 1015 689 1016
rect 683 1014 689 1015
rect 722 1015 723 1016
rect 727 1015 728 1019
rect 722 1014 728 1015
rect 819 1019 828 1020
rect 819 1015 820 1019
rect 827 1015 828 1019
rect 819 1014 828 1015
rect 979 1019 985 1020
rect 979 1015 980 1019
rect 984 1018 985 1019
rect 1038 1019 1044 1020
rect 1038 1018 1039 1019
rect 984 1016 1039 1018
rect 984 1015 985 1016
rect 979 1014 985 1015
rect 1038 1015 1039 1016
rect 1043 1015 1044 1019
rect 1038 1014 1044 1015
rect 1163 1019 1169 1020
rect 1163 1015 1164 1019
rect 1168 1018 1169 1019
rect 1202 1019 1208 1020
rect 1202 1018 1203 1019
rect 1168 1016 1203 1018
rect 1168 1015 1169 1016
rect 1163 1014 1169 1015
rect 1202 1015 1203 1016
rect 1207 1015 1208 1019
rect 1202 1014 1208 1015
rect 1278 1019 1284 1020
rect 1278 1015 1279 1019
rect 1283 1018 1284 1019
rect 1355 1019 1361 1020
rect 1355 1018 1356 1019
rect 1283 1016 1356 1018
rect 1283 1015 1284 1016
rect 1278 1014 1284 1015
rect 1355 1015 1356 1016
rect 1360 1015 1361 1019
rect 1355 1014 1361 1015
rect 1563 1019 1572 1020
rect 1563 1015 1564 1019
rect 1571 1015 1572 1019
rect 1563 1014 1572 1015
rect 1623 1019 1629 1020
rect 1623 1015 1624 1019
rect 1628 1018 1629 1019
rect 1763 1019 1769 1020
rect 1763 1018 1764 1019
rect 1628 1016 1764 1018
rect 1628 1015 1629 1016
rect 1623 1014 1629 1015
rect 1763 1015 1764 1016
rect 1768 1015 1769 1019
rect 1763 1014 1769 1015
rect 1971 1019 1977 1020
rect 1971 1015 1972 1019
rect 1976 1018 1977 1019
rect 2010 1019 2016 1020
rect 2010 1018 2011 1019
rect 1976 1016 2011 1018
rect 1976 1015 1977 1016
rect 1971 1014 1977 1015
rect 2010 1015 2011 1016
rect 2015 1015 2016 1019
rect 2010 1014 2016 1015
rect 2099 1019 2105 1020
rect 2099 1015 2100 1019
rect 2104 1018 2105 1019
rect 2114 1019 2120 1020
rect 2114 1018 2115 1019
rect 2104 1016 2115 1018
rect 2104 1015 2105 1016
rect 2099 1014 2105 1015
rect 2114 1015 2115 1016
rect 2119 1015 2120 1019
rect 2114 1014 2120 1015
rect 2151 1019 2157 1020
rect 2151 1015 2152 1019
rect 2156 1018 2157 1019
rect 2219 1019 2225 1020
rect 2219 1018 2220 1019
rect 2156 1016 2220 1018
rect 2156 1015 2157 1016
rect 2151 1014 2157 1015
rect 2219 1015 2220 1016
rect 2224 1015 2225 1019
rect 2219 1014 2225 1015
rect 2271 1019 2277 1020
rect 2271 1015 2272 1019
rect 2276 1018 2277 1019
rect 2339 1019 2345 1020
rect 2339 1018 2340 1019
rect 2276 1016 2340 1018
rect 2276 1015 2277 1016
rect 2271 1014 2277 1015
rect 2339 1015 2340 1016
rect 2344 1015 2345 1019
rect 2339 1014 2345 1015
rect 2391 1019 2397 1020
rect 2391 1015 2392 1019
rect 2396 1018 2397 1019
rect 2467 1019 2473 1020
rect 2467 1018 2468 1019
rect 2396 1016 2468 1018
rect 2396 1015 2397 1016
rect 2391 1014 2397 1015
rect 2467 1015 2468 1016
rect 2472 1015 2473 1019
rect 2467 1014 2473 1015
rect 2603 1019 2609 1020
rect 2603 1015 2604 1019
rect 2608 1018 2609 1019
rect 2642 1019 2648 1020
rect 2642 1018 2643 1019
rect 2608 1016 2643 1018
rect 2608 1015 2609 1016
rect 2603 1014 2609 1015
rect 2642 1015 2643 1016
rect 2647 1015 2648 1019
rect 2642 1014 2648 1015
rect 2663 1019 2669 1020
rect 2663 1015 2664 1019
rect 2668 1018 2669 1019
rect 2747 1019 2753 1020
rect 2747 1018 2748 1019
rect 2668 1016 2748 1018
rect 2668 1015 2669 1016
rect 2663 1014 2669 1015
rect 2747 1015 2748 1016
rect 2752 1015 2753 1019
rect 2747 1014 2753 1015
rect 2823 1019 2829 1020
rect 2823 1015 2824 1019
rect 2828 1018 2829 1019
rect 2899 1019 2905 1020
rect 2899 1018 2900 1019
rect 2828 1016 2900 1018
rect 2828 1015 2829 1016
rect 2823 1014 2829 1015
rect 2899 1015 2900 1016
rect 2904 1015 2905 1019
rect 2899 1014 2905 1015
rect 2967 1019 2973 1020
rect 2967 1015 2968 1019
rect 2972 1018 2973 1019
rect 3059 1019 3065 1020
rect 3059 1018 3060 1019
rect 2972 1016 3060 1018
rect 2972 1015 2973 1016
rect 2967 1014 2973 1015
rect 3059 1015 3060 1016
rect 3064 1015 3065 1019
rect 3059 1014 3065 1015
rect 3219 1019 3225 1020
rect 3219 1015 3220 1019
rect 3224 1018 3225 1019
rect 3287 1019 3293 1020
rect 3287 1018 3288 1019
rect 3224 1016 3288 1018
rect 3224 1015 3225 1016
rect 3219 1014 3225 1015
rect 3287 1015 3288 1016
rect 3292 1015 3293 1019
rect 3287 1014 3293 1015
rect 3379 1019 3385 1020
rect 3379 1015 3380 1019
rect 3384 1018 3385 1019
rect 3418 1019 3424 1020
rect 3418 1018 3419 1019
rect 3384 1016 3419 1018
rect 3384 1015 3385 1016
rect 3379 1014 3385 1015
rect 3418 1015 3419 1016
rect 3423 1015 3424 1019
rect 3418 1014 3424 1015
rect 3515 1019 3521 1020
rect 3515 1015 3516 1019
rect 3520 1018 3521 1019
rect 3546 1019 3552 1020
rect 3546 1018 3547 1019
rect 3520 1016 3547 1018
rect 3520 1015 3521 1016
rect 3515 1014 3521 1015
rect 3546 1015 3547 1016
rect 3551 1015 3552 1019
rect 3546 1014 3552 1015
rect 342 1009 348 1010
rect 342 1005 343 1009
rect 347 1005 348 1009
rect 342 1004 348 1005
rect 430 1009 436 1010
rect 430 1005 431 1009
rect 435 1005 436 1009
rect 430 1004 436 1005
rect 534 1009 540 1010
rect 534 1005 535 1009
rect 539 1005 540 1009
rect 534 1004 540 1005
rect 654 1009 660 1010
rect 654 1005 655 1009
rect 659 1005 660 1009
rect 654 1004 660 1005
rect 790 1009 796 1010
rect 790 1005 791 1009
rect 795 1005 796 1009
rect 790 1004 796 1005
rect 950 1009 956 1010
rect 950 1005 951 1009
rect 955 1005 956 1009
rect 950 1004 956 1005
rect 1134 1009 1140 1010
rect 1134 1005 1135 1009
rect 1139 1005 1140 1009
rect 1134 1004 1140 1005
rect 1326 1009 1332 1010
rect 1326 1005 1327 1009
rect 1331 1005 1332 1009
rect 1326 1004 1332 1005
rect 1534 1009 1540 1010
rect 1534 1005 1535 1009
rect 1539 1005 1540 1009
rect 1534 1004 1540 1005
rect 1734 1009 1740 1010
rect 1734 1005 1735 1009
rect 1739 1005 1740 1009
rect 1734 1004 1740 1005
rect 1942 1009 1948 1010
rect 1942 1005 1943 1009
rect 1947 1005 1948 1009
rect 1942 1004 1948 1005
rect 2070 1009 2076 1010
rect 2070 1005 2071 1009
rect 2075 1005 2076 1009
rect 2070 1004 2076 1005
rect 2190 1009 2196 1010
rect 2190 1005 2191 1009
rect 2195 1005 2196 1009
rect 2190 1004 2196 1005
rect 2310 1009 2316 1010
rect 2310 1005 2311 1009
rect 2315 1005 2316 1009
rect 2310 1004 2316 1005
rect 2438 1009 2444 1010
rect 2438 1005 2439 1009
rect 2443 1005 2444 1009
rect 2438 1004 2444 1005
rect 2574 1009 2580 1010
rect 2574 1005 2575 1009
rect 2579 1005 2580 1009
rect 2574 1004 2580 1005
rect 2718 1009 2724 1010
rect 2718 1005 2719 1009
rect 2723 1005 2724 1009
rect 2718 1004 2724 1005
rect 2870 1009 2876 1010
rect 2870 1005 2871 1009
rect 2875 1005 2876 1009
rect 2870 1004 2876 1005
rect 3030 1009 3036 1010
rect 3030 1005 3031 1009
rect 3035 1005 3036 1009
rect 3030 1004 3036 1005
rect 3190 1009 3196 1010
rect 3190 1005 3191 1009
rect 3195 1005 3196 1009
rect 3190 1004 3196 1005
rect 3350 1009 3356 1010
rect 3350 1005 3351 1009
rect 3355 1005 3356 1009
rect 3350 1004 3356 1005
rect 3486 1009 3492 1010
rect 3486 1005 3487 1009
rect 3491 1005 3492 1009
rect 3486 1004 3492 1005
rect 110 996 116 997
rect 1822 996 1828 997
rect 110 992 111 996
rect 115 992 116 996
rect 714 995 720 996
rect 714 994 715 995
rect 709 992 715 994
rect 110 991 116 992
rect 410 991 416 992
rect 410 987 411 991
rect 415 990 416 991
rect 502 991 508 992
rect 415 988 449 990
rect 415 987 416 988
rect 410 986 416 987
rect 502 987 503 991
rect 507 990 508 991
rect 714 991 715 992
rect 719 991 720 995
rect 1623 995 1629 996
rect 1623 994 1624 995
rect 1589 992 1624 994
rect 714 990 720 991
rect 722 991 728 992
rect 507 988 553 990
rect 507 987 508 988
rect 502 986 508 987
rect 722 987 723 991
rect 727 990 728 991
rect 858 991 864 992
rect 727 988 809 990
rect 727 987 728 988
rect 722 986 728 987
rect 858 987 859 991
rect 863 990 864 991
rect 1038 991 1044 992
rect 863 988 969 990
rect 863 987 864 988
rect 858 986 864 987
rect 1038 987 1039 991
rect 1043 990 1044 991
rect 1202 991 1208 992
rect 1043 988 1153 990
rect 1043 987 1044 988
rect 1038 986 1044 987
rect 1202 987 1203 991
rect 1207 990 1208 991
rect 1623 991 1624 992
rect 1628 991 1629 995
rect 1822 992 1823 996
rect 1827 992 1828 996
rect 1822 991 1828 992
rect 1862 996 1868 997
rect 3574 996 3580 997
rect 1862 992 1863 996
rect 1867 992 1868 996
rect 2151 995 2157 996
rect 2151 994 2152 995
rect 2125 992 2152 994
rect 1862 991 1868 992
rect 2151 991 2152 992
rect 2156 991 2157 995
rect 2271 995 2277 996
rect 2271 994 2272 995
rect 2245 992 2272 994
rect 1623 990 1629 991
rect 2151 990 2157 991
rect 2271 991 2272 992
rect 2276 991 2277 995
rect 2391 995 2397 996
rect 2391 994 2392 995
rect 2365 992 2392 994
rect 2271 990 2277 991
rect 2391 991 2392 992
rect 2396 991 2397 995
rect 2663 995 2669 996
rect 2663 994 2664 995
rect 2629 992 2664 994
rect 2391 990 2397 991
rect 2663 991 2664 992
rect 2668 991 2669 995
rect 2823 995 2829 996
rect 2823 994 2824 995
rect 2773 992 2824 994
rect 2663 990 2669 991
rect 2823 991 2824 992
rect 2828 991 2829 995
rect 2967 995 2973 996
rect 2967 994 2968 995
rect 2925 992 2968 994
rect 2823 990 2829 991
rect 2967 991 2968 992
rect 2972 991 2973 995
rect 3263 995 3269 996
rect 3263 994 3264 995
rect 3245 992 3264 994
rect 2967 990 2973 991
rect 3263 991 3264 992
rect 3268 991 3269 995
rect 3574 992 3575 996
rect 3579 992 3580 996
rect 3263 990 3269 991
rect 3287 991 3293 992
rect 1207 988 1345 990
rect 1207 987 1208 988
rect 1202 986 1208 987
rect 3287 987 3288 991
rect 3292 990 3293 991
rect 3418 991 3424 992
rect 3574 991 3580 992
rect 3292 988 3369 990
rect 3292 987 3293 988
rect 3287 986 3293 987
rect 3418 987 3419 991
rect 3423 990 3424 991
rect 3423 988 3505 990
rect 3423 987 3424 988
rect 3418 986 3424 987
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 110 974 116 975
rect 1734 979 1740 980
rect 1734 975 1735 979
rect 1739 978 1740 979
rect 1822 979 1828 980
rect 1739 976 1745 978
rect 1739 975 1740 976
rect 1734 974 1740 975
rect 1822 975 1823 979
rect 1827 975 1828 979
rect 1822 974 1828 975
rect 1862 979 1868 980
rect 1862 975 1863 979
rect 1867 975 1868 979
rect 1862 974 1868 975
rect 1942 979 1948 980
rect 1942 975 1943 979
rect 1947 978 1948 979
rect 2378 979 2384 980
rect 1947 976 1953 978
rect 1947 975 1948 976
rect 1942 974 1948 975
rect 2378 975 2379 979
rect 2383 978 2384 979
rect 2958 979 2964 980
rect 2383 976 2449 978
rect 2383 975 2384 976
rect 2378 974 2384 975
rect 2958 975 2959 979
rect 2963 978 2964 979
rect 3574 979 3580 980
rect 2963 976 3041 978
rect 2963 975 2964 976
rect 2958 974 2964 975
rect 3574 975 3575 979
rect 3579 975 3580 979
rect 3574 974 3580 975
rect 334 969 340 970
rect 334 965 335 969
rect 339 965 340 969
rect 334 964 340 965
rect 422 969 428 970
rect 422 965 423 969
rect 427 965 428 969
rect 422 964 428 965
rect 526 969 532 970
rect 526 965 527 969
rect 531 965 532 969
rect 526 964 532 965
rect 646 969 652 970
rect 646 965 647 969
rect 651 965 652 969
rect 646 964 652 965
rect 782 969 788 970
rect 782 965 783 969
rect 787 965 788 969
rect 782 964 788 965
rect 942 969 948 970
rect 942 965 943 969
rect 947 965 948 969
rect 942 964 948 965
rect 1126 969 1132 970
rect 1126 965 1127 969
rect 1131 965 1132 969
rect 1126 964 1132 965
rect 1318 969 1324 970
rect 1318 965 1319 969
rect 1323 965 1324 969
rect 1318 964 1324 965
rect 1526 969 1532 970
rect 1526 965 1527 969
rect 1531 965 1532 969
rect 1526 964 1532 965
rect 1726 969 1732 970
rect 1726 965 1727 969
rect 1731 965 1732 969
rect 1726 964 1732 965
rect 1934 969 1940 970
rect 1934 965 1935 969
rect 1939 965 1940 969
rect 1934 964 1940 965
rect 2062 969 2068 970
rect 2062 965 2063 969
rect 2067 965 2068 969
rect 2062 964 2068 965
rect 2182 969 2188 970
rect 2182 965 2183 969
rect 2187 965 2188 969
rect 2182 964 2188 965
rect 2302 969 2308 970
rect 2302 965 2303 969
rect 2307 965 2308 969
rect 2302 964 2308 965
rect 2430 969 2436 970
rect 2430 965 2431 969
rect 2435 965 2436 969
rect 2430 964 2436 965
rect 2566 969 2572 970
rect 2566 965 2567 969
rect 2571 965 2572 969
rect 2566 964 2572 965
rect 2710 969 2716 970
rect 2710 965 2711 969
rect 2715 965 2716 969
rect 2710 964 2716 965
rect 2862 969 2868 970
rect 2862 965 2863 969
rect 2867 965 2868 969
rect 2862 964 2868 965
rect 3022 969 3028 970
rect 3022 965 3023 969
rect 3027 965 3028 969
rect 3022 964 3028 965
rect 3182 969 3188 970
rect 3182 965 3183 969
rect 3187 965 3188 969
rect 3182 964 3188 965
rect 3342 969 3348 970
rect 3342 965 3343 969
rect 3347 965 3348 969
rect 3342 964 3348 965
rect 3478 969 3484 970
rect 3478 965 3479 969
rect 3483 965 3484 969
rect 3478 964 3484 965
rect 383 963 389 964
rect 383 959 384 963
rect 388 962 389 963
rect 402 963 408 964
rect 402 962 403 963
rect 388 960 403 962
rect 388 959 389 960
rect 383 958 389 959
rect 402 959 403 960
rect 407 959 408 963
rect 402 958 408 959
rect 2534 955 2540 956
rect 2534 951 2535 955
rect 2539 954 2540 955
rect 2958 955 2964 956
rect 2958 954 2959 955
rect 2539 952 2959 954
rect 2539 951 2540 952
rect 2534 950 2540 951
rect 2958 951 2959 952
rect 2963 951 2964 955
rect 2958 950 2964 951
rect 366 943 372 944
rect 366 939 367 943
rect 371 939 372 943
rect 366 938 372 939
rect 462 943 468 944
rect 462 939 463 943
rect 467 939 468 943
rect 462 938 468 939
rect 574 943 580 944
rect 574 939 575 943
rect 579 939 580 943
rect 574 938 580 939
rect 702 943 708 944
rect 702 939 703 943
rect 707 939 708 943
rect 702 938 708 939
rect 846 943 852 944
rect 846 939 847 943
rect 851 939 852 943
rect 846 938 852 939
rect 1006 943 1012 944
rect 1006 939 1007 943
rect 1011 939 1012 943
rect 1006 938 1012 939
rect 1174 943 1180 944
rect 1174 939 1175 943
rect 1179 939 1180 943
rect 1174 938 1180 939
rect 1350 943 1356 944
rect 1350 939 1351 943
rect 1355 939 1356 943
rect 1350 938 1356 939
rect 1526 943 1532 944
rect 1526 939 1527 943
rect 1531 939 1532 943
rect 1526 938 1532 939
rect 1710 943 1716 944
rect 1710 939 1711 943
rect 1715 939 1716 943
rect 1710 938 1716 939
rect 1886 943 1892 944
rect 1886 939 1887 943
rect 1891 939 1892 943
rect 1886 938 1892 939
rect 2046 943 2052 944
rect 2046 939 2047 943
rect 2051 939 2052 943
rect 2046 938 2052 939
rect 2198 943 2204 944
rect 2198 939 2199 943
rect 2203 939 2204 943
rect 2198 938 2204 939
rect 2350 943 2356 944
rect 2350 939 2351 943
rect 2355 939 2356 943
rect 2350 938 2356 939
rect 2494 943 2500 944
rect 2494 939 2495 943
rect 2499 939 2500 943
rect 2494 938 2500 939
rect 2630 943 2636 944
rect 2630 939 2631 943
rect 2635 939 2636 943
rect 2630 938 2636 939
rect 2758 943 2764 944
rect 2758 939 2759 943
rect 2763 939 2764 943
rect 2758 938 2764 939
rect 2886 943 2892 944
rect 2886 939 2887 943
rect 2891 939 2892 943
rect 2886 938 2892 939
rect 3022 943 3028 944
rect 3022 939 3023 943
rect 3027 939 3028 943
rect 3022 938 3028 939
rect 822 935 828 936
rect 110 933 116 934
rect 110 929 111 933
rect 115 929 116 933
rect 822 931 823 935
rect 827 934 828 935
rect 1278 935 1284 936
rect 1278 934 1279 935
rect 827 932 865 934
rect 1233 932 1279 934
rect 827 931 828 932
rect 822 930 828 931
rect 1278 931 1279 932
rect 1283 931 1284 935
rect 2114 935 2120 936
rect 1278 930 1284 931
rect 1822 933 1828 934
rect 110 928 116 929
rect 1822 929 1823 933
rect 1827 929 1828 933
rect 1822 928 1828 929
rect 1862 933 1868 934
rect 1862 929 1863 933
rect 1867 929 1868 933
rect 2114 931 2115 935
rect 2119 934 2120 935
rect 2119 932 2217 934
rect 3574 933 3580 934
rect 2119 931 2120 932
rect 2114 930 2120 931
rect 1862 928 1868 929
rect 3574 929 3575 933
rect 3579 929 3580 933
rect 3574 928 3580 929
rect 455 919 461 920
rect 455 918 456 919
rect 110 916 116 917
rect 429 916 456 918
rect 110 912 111 916
rect 115 912 116 916
rect 455 915 456 916
rect 460 915 461 919
rect 562 919 568 920
rect 562 918 563 919
rect 525 916 563 918
rect 455 914 461 915
rect 562 915 563 916
rect 567 915 568 919
rect 695 919 701 920
rect 695 918 696 919
rect 637 916 696 918
rect 562 914 568 915
rect 695 915 696 916
rect 700 915 701 919
rect 839 919 845 920
rect 839 918 840 919
rect 765 916 840 918
rect 695 914 701 915
rect 839 915 840 916
rect 844 915 845 919
rect 1166 919 1172 920
rect 1166 918 1167 919
rect 1069 916 1167 918
rect 839 914 845 915
rect 1166 915 1167 916
rect 1171 915 1172 919
rect 1519 919 1525 920
rect 1519 918 1520 919
rect 1413 916 1520 918
rect 1166 914 1172 915
rect 1519 915 1520 916
rect 1524 915 1525 919
rect 1658 919 1664 920
rect 1658 918 1659 919
rect 1589 916 1659 918
rect 1519 914 1525 915
rect 1658 915 1659 916
rect 1663 915 1664 919
rect 1658 914 1664 915
rect 1666 919 1672 920
rect 1666 915 1667 919
rect 1671 918 1672 919
rect 2015 919 2021 920
rect 2015 918 2016 919
rect 1671 916 1737 918
rect 1822 916 1828 917
rect 1671 915 1672 916
rect 1666 914 1672 915
rect 110 911 116 912
rect 1822 912 1823 916
rect 1827 912 1828 916
rect 1822 911 1828 912
rect 1862 916 1868 917
rect 1949 916 2016 918
rect 1862 912 1863 916
rect 1867 912 1868 916
rect 2015 915 2016 916
rect 2020 915 2021 919
rect 2015 914 2021 915
rect 2038 919 2044 920
rect 2038 915 2039 919
rect 2043 918 2044 919
rect 2266 919 2272 920
rect 2043 916 2073 918
rect 2043 915 2044 916
rect 2038 914 2044 915
rect 2266 915 2267 919
rect 2271 918 2272 919
rect 2623 919 2629 920
rect 2623 918 2624 919
rect 2271 916 2377 918
rect 2557 916 2624 918
rect 2271 915 2272 916
rect 2266 914 2272 915
rect 2623 915 2624 916
rect 2628 915 2629 919
rect 2714 919 2720 920
rect 2714 918 2715 919
rect 2693 916 2715 918
rect 2623 914 2629 915
rect 2714 915 2715 916
rect 2719 915 2720 919
rect 2854 919 2860 920
rect 2854 918 2855 919
rect 2821 916 2855 918
rect 2714 914 2720 915
rect 2854 915 2855 916
rect 2859 915 2860 919
rect 3015 919 3021 920
rect 3015 918 3016 919
rect 2949 916 3016 918
rect 2854 914 2860 915
rect 3015 915 3016 916
rect 3020 915 3021 919
rect 3090 919 3096 920
rect 3090 918 3091 919
rect 3085 916 3091 918
rect 3015 914 3021 915
rect 3090 915 3091 916
rect 3095 915 3096 919
rect 3090 914 3096 915
rect 3574 916 3580 917
rect 1862 911 1868 912
rect 3574 912 3575 916
rect 3579 912 3580 916
rect 3574 911 3580 912
rect 374 903 380 904
rect 374 899 375 903
rect 379 899 380 903
rect 374 898 380 899
rect 470 903 476 904
rect 470 899 471 903
rect 475 899 476 903
rect 470 898 476 899
rect 582 903 588 904
rect 582 899 583 903
rect 587 899 588 903
rect 582 898 588 899
rect 710 903 716 904
rect 710 899 711 903
rect 715 899 716 903
rect 710 898 716 899
rect 854 903 860 904
rect 854 899 855 903
rect 859 899 860 903
rect 854 898 860 899
rect 1014 903 1020 904
rect 1014 899 1015 903
rect 1019 899 1020 903
rect 1014 898 1020 899
rect 1182 903 1188 904
rect 1182 899 1183 903
rect 1187 899 1188 903
rect 1182 898 1188 899
rect 1358 903 1364 904
rect 1358 899 1359 903
rect 1363 899 1364 903
rect 1358 898 1364 899
rect 1534 903 1540 904
rect 1534 899 1535 903
rect 1539 899 1540 903
rect 1534 898 1540 899
rect 1718 903 1724 904
rect 1718 899 1719 903
rect 1723 899 1724 903
rect 1718 898 1724 899
rect 1894 903 1900 904
rect 1894 899 1895 903
rect 1899 899 1900 903
rect 1894 898 1900 899
rect 2054 903 2060 904
rect 2054 899 2055 903
rect 2059 899 2060 903
rect 2054 898 2060 899
rect 2206 903 2212 904
rect 2206 899 2207 903
rect 2211 899 2212 903
rect 2206 898 2212 899
rect 2358 903 2364 904
rect 2358 899 2359 903
rect 2363 899 2364 903
rect 2358 898 2364 899
rect 2502 903 2508 904
rect 2502 899 2503 903
rect 2507 899 2508 903
rect 2502 898 2508 899
rect 2638 903 2644 904
rect 2638 899 2639 903
rect 2643 899 2644 903
rect 2638 898 2644 899
rect 2766 903 2772 904
rect 2766 899 2767 903
rect 2771 899 2772 903
rect 2766 898 2772 899
rect 2894 903 2900 904
rect 2894 899 2895 903
rect 2899 899 2900 903
rect 2894 898 2900 899
rect 3030 903 3036 904
rect 3030 899 3031 903
rect 3035 899 3036 903
rect 3030 898 3036 899
rect 402 891 409 892
rect 402 887 403 891
rect 408 887 409 891
rect 402 886 409 887
rect 455 891 461 892
rect 455 887 456 891
rect 460 890 461 891
rect 499 891 505 892
rect 499 890 500 891
rect 460 888 500 890
rect 460 887 461 888
rect 455 886 461 887
rect 499 887 500 888
rect 504 887 505 891
rect 499 886 505 887
rect 611 891 617 892
rect 611 887 612 891
rect 616 890 617 891
rect 634 891 640 892
rect 634 890 635 891
rect 616 888 635 890
rect 616 887 617 888
rect 611 886 617 887
rect 634 887 635 888
rect 639 887 640 891
rect 634 886 640 887
rect 695 891 701 892
rect 695 887 696 891
rect 700 890 701 891
rect 739 891 745 892
rect 739 890 740 891
rect 700 888 740 890
rect 700 887 701 888
rect 695 886 701 887
rect 739 887 740 888
rect 744 887 745 891
rect 739 886 745 887
rect 839 891 845 892
rect 839 887 840 891
rect 844 890 845 891
rect 883 891 889 892
rect 883 890 884 891
rect 844 888 884 890
rect 844 887 845 888
rect 839 886 845 887
rect 883 887 884 888
rect 888 887 889 891
rect 883 886 889 887
rect 991 891 997 892
rect 991 887 992 891
rect 996 890 997 891
rect 1043 891 1049 892
rect 1043 890 1044 891
rect 996 888 1044 890
rect 996 887 997 888
rect 991 886 997 887
rect 1043 887 1044 888
rect 1048 887 1049 891
rect 1043 886 1049 887
rect 1166 891 1172 892
rect 1166 887 1167 891
rect 1171 890 1172 891
rect 1211 891 1217 892
rect 1211 890 1212 891
rect 1171 888 1212 890
rect 1171 887 1172 888
rect 1166 886 1172 887
rect 1211 887 1212 888
rect 1216 887 1217 891
rect 1211 886 1217 887
rect 1387 891 1396 892
rect 1387 887 1388 891
rect 1395 887 1396 891
rect 1387 886 1396 887
rect 1519 891 1525 892
rect 1519 887 1520 891
rect 1524 890 1525 891
rect 1563 891 1569 892
rect 1563 890 1564 891
rect 1524 888 1564 890
rect 1524 887 1525 888
rect 1519 886 1525 887
rect 1563 887 1564 888
rect 1568 887 1569 891
rect 1563 886 1569 887
rect 1734 891 1740 892
rect 1734 887 1735 891
rect 1739 890 1740 891
rect 1747 891 1753 892
rect 1747 890 1748 891
rect 1739 888 1748 890
rect 1739 887 1740 888
rect 1734 886 1740 887
rect 1747 887 1748 888
rect 1752 887 1753 891
rect 1747 886 1753 887
rect 1923 891 1929 892
rect 1923 887 1924 891
rect 1928 890 1929 891
rect 1942 891 1948 892
rect 1942 890 1943 891
rect 1928 888 1943 890
rect 1928 887 1929 888
rect 1923 886 1929 887
rect 1942 887 1943 888
rect 1947 887 1948 891
rect 1942 886 1948 887
rect 2015 891 2021 892
rect 2015 887 2016 891
rect 2020 890 2021 891
rect 2083 891 2089 892
rect 2083 890 2084 891
rect 2020 888 2084 890
rect 2020 887 2021 888
rect 2015 886 2021 887
rect 2083 887 2084 888
rect 2088 887 2089 891
rect 2083 886 2089 887
rect 2235 891 2241 892
rect 2235 887 2236 891
rect 2240 890 2241 891
rect 2266 891 2272 892
rect 2266 890 2267 891
rect 2240 888 2267 890
rect 2240 887 2241 888
rect 2235 886 2241 887
rect 2266 887 2267 888
rect 2271 887 2272 891
rect 2266 886 2272 887
rect 2387 891 2396 892
rect 2387 887 2388 891
rect 2395 887 2396 891
rect 2387 886 2396 887
rect 2531 891 2540 892
rect 2531 887 2532 891
rect 2539 887 2540 891
rect 2531 886 2540 887
rect 2623 891 2629 892
rect 2623 887 2624 891
rect 2628 890 2629 891
rect 2667 891 2673 892
rect 2667 890 2668 891
rect 2628 888 2668 890
rect 2628 887 2629 888
rect 2623 886 2629 887
rect 2667 887 2668 888
rect 2672 887 2673 891
rect 2667 886 2673 887
rect 2714 891 2720 892
rect 2714 887 2715 891
rect 2719 890 2720 891
rect 2795 891 2801 892
rect 2795 890 2796 891
rect 2719 888 2796 890
rect 2719 887 2720 888
rect 2714 886 2720 887
rect 2795 887 2796 888
rect 2800 887 2801 891
rect 2795 886 2801 887
rect 2854 891 2860 892
rect 2854 887 2855 891
rect 2859 890 2860 891
rect 2923 891 2929 892
rect 2923 890 2924 891
rect 2859 888 2924 890
rect 2859 887 2860 888
rect 2854 886 2860 887
rect 2923 887 2924 888
rect 2928 887 2929 891
rect 2923 886 2929 887
rect 3015 891 3021 892
rect 3015 887 3016 891
rect 3020 890 3021 891
rect 3059 891 3065 892
rect 3059 890 3060 891
rect 3020 888 3060 890
rect 3020 887 3021 888
rect 3015 886 3021 887
rect 3059 887 3060 888
rect 3064 887 3065 891
rect 3059 886 3065 887
rect 1923 879 1929 880
rect 371 875 377 876
rect 371 871 372 875
rect 376 874 377 875
rect 410 875 416 876
rect 410 874 411 875
rect 376 872 411 874
rect 376 871 377 872
rect 371 870 377 871
rect 410 871 411 872
rect 415 871 416 875
rect 410 870 416 871
rect 459 875 465 876
rect 459 871 460 875
rect 464 874 465 875
rect 502 875 508 876
rect 502 874 503 875
rect 464 872 503 874
rect 464 871 465 872
rect 459 870 465 871
rect 502 871 503 872
rect 507 871 508 875
rect 502 870 508 871
rect 562 875 569 876
rect 562 871 563 875
rect 568 871 569 875
rect 562 870 569 871
rect 675 875 681 876
rect 675 871 676 875
rect 680 874 681 875
rect 718 875 724 876
rect 718 874 719 875
rect 680 872 719 874
rect 680 871 681 872
rect 675 870 681 871
rect 718 871 719 872
rect 723 871 724 875
rect 718 870 724 871
rect 811 875 820 876
rect 811 871 812 875
rect 819 871 820 875
rect 811 870 820 871
rect 955 875 961 876
rect 955 871 956 875
rect 960 874 961 875
rect 1026 875 1032 876
rect 1026 874 1027 875
rect 960 872 1027 874
rect 960 871 961 872
rect 955 870 961 871
rect 1026 871 1027 872
rect 1031 871 1032 875
rect 1026 870 1032 871
rect 1115 875 1121 876
rect 1115 871 1116 875
rect 1120 874 1121 875
rect 1194 875 1200 876
rect 1194 874 1195 875
rect 1120 872 1195 874
rect 1120 871 1121 872
rect 1115 870 1121 871
rect 1194 871 1195 872
rect 1199 871 1200 875
rect 1194 870 1200 871
rect 1222 875 1228 876
rect 1222 871 1223 875
rect 1227 874 1228 875
rect 1291 875 1297 876
rect 1291 874 1292 875
rect 1227 872 1292 874
rect 1227 871 1228 872
rect 1222 870 1228 871
rect 1291 871 1292 872
rect 1296 871 1297 875
rect 1291 870 1297 871
rect 1475 875 1481 876
rect 1475 871 1476 875
rect 1480 874 1481 875
rect 1518 875 1524 876
rect 1518 874 1519 875
rect 1480 872 1519 874
rect 1480 871 1481 872
rect 1475 870 1481 871
rect 1518 871 1519 872
rect 1523 871 1524 875
rect 1518 870 1524 871
rect 1658 875 1665 876
rect 1658 871 1659 875
rect 1664 871 1665 875
rect 1923 875 1924 879
rect 1928 878 1929 879
rect 1966 879 1972 880
rect 1966 878 1967 879
rect 1928 876 1967 878
rect 1928 875 1929 876
rect 1923 874 1929 875
rect 1966 875 1967 876
rect 1971 875 1972 879
rect 1966 874 1972 875
rect 2038 879 2049 880
rect 2038 875 2039 879
rect 2043 875 2044 879
rect 2048 875 2049 879
rect 2038 874 2049 875
rect 2195 879 2201 880
rect 2195 875 2196 879
rect 2200 875 2201 879
rect 2263 879 2269 880
rect 2195 874 2201 875
rect 2206 875 2212 876
rect 2206 874 2207 875
rect 2197 872 2207 874
rect 1658 870 1665 871
rect 2206 871 2207 872
rect 2211 871 2212 875
rect 2263 875 2264 879
rect 2268 878 2269 879
rect 2347 879 2353 880
rect 2347 878 2348 879
rect 2268 876 2348 878
rect 2268 875 2269 876
rect 2263 874 2269 875
rect 2347 875 2348 876
rect 2352 875 2353 879
rect 2347 874 2353 875
rect 2382 879 2388 880
rect 2382 875 2383 879
rect 2387 878 2388 879
rect 2515 879 2521 880
rect 2515 878 2516 879
rect 2387 876 2516 878
rect 2387 875 2388 876
rect 2382 874 2388 875
rect 2515 875 2516 876
rect 2520 875 2521 879
rect 2515 874 2521 875
rect 2691 879 2697 880
rect 2691 875 2692 879
rect 2696 878 2697 879
rect 2759 879 2765 880
rect 2759 878 2760 879
rect 2696 876 2760 878
rect 2696 875 2697 876
rect 2691 874 2697 875
rect 2759 875 2760 876
rect 2764 875 2765 879
rect 2759 874 2765 875
rect 2875 879 2884 880
rect 2875 875 2876 879
rect 2883 875 2884 879
rect 2875 874 2884 875
rect 3067 879 3073 880
rect 3067 875 3068 879
rect 3072 878 3073 879
rect 3090 879 3096 880
rect 3090 878 3091 879
rect 3072 876 3091 878
rect 3072 875 3073 876
rect 3067 874 3073 875
rect 3090 875 3091 876
rect 3095 875 3096 879
rect 3090 874 3096 875
rect 3159 879 3165 880
rect 3159 875 3160 879
rect 3164 878 3165 879
rect 3267 879 3273 880
rect 3267 878 3268 879
rect 3164 876 3268 878
rect 3164 875 3165 876
rect 3159 874 3165 875
rect 3267 875 3268 876
rect 3272 875 3273 879
rect 3267 874 3273 875
rect 3406 879 3412 880
rect 3406 875 3407 879
rect 3411 878 3412 879
rect 3467 879 3473 880
rect 3467 878 3468 879
rect 3411 876 3468 878
rect 3411 875 3412 876
rect 3406 874 3412 875
rect 3467 875 3468 876
rect 3472 875 3473 879
rect 3467 874 3473 875
rect 2206 870 2212 871
rect 1894 869 1900 870
rect 342 865 348 866
rect 342 861 343 865
rect 347 861 348 865
rect 342 860 348 861
rect 430 865 436 866
rect 430 861 431 865
rect 435 861 436 865
rect 430 860 436 861
rect 534 865 540 866
rect 534 861 535 865
rect 539 861 540 865
rect 534 860 540 861
rect 646 865 652 866
rect 646 861 647 865
rect 651 861 652 865
rect 646 860 652 861
rect 782 865 788 866
rect 782 861 783 865
rect 787 861 788 865
rect 782 860 788 861
rect 926 865 932 866
rect 926 861 927 865
rect 931 861 932 865
rect 926 860 932 861
rect 1086 865 1092 866
rect 1086 861 1087 865
rect 1091 861 1092 865
rect 1086 860 1092 861
rect 1262 865 1268 866
rect 1262 861 1263 865
rect 1267 861 1268 865
rect 1262 860 1268 861
rect 1446 865 1452 866
rect 1446 861 1447 865
rect 1451 861 1452 865
rect 1446 860 1452 861
rect 1630 865 1636 866
rect 1630 861 1631 865
rect 1635 861 1636 865
rect 1894 865 1895 869
rect 1899 865 1900 869
rect 1894 864 1900 865
rect 2014 869 2020 870
rect 2014 865 2015 869
rect 2019 865 2020 869
rect 2014 864 2020 865
rect 2166 869 2172 870
rect 2166 865 2167 869
rect 2171 865 2172 869
rect 2166 864 2172 865
rect 2318 869 2324 870
rect 2318 865 2319 869
rect 2323 865 2324 869
rect 2318 864 2324 865
rect 2486 869 2492 870
rect 2486 865 2487 869
rect 2491 865 2492 869
rect 2486 864 2492 865
rect 2662 869 2668 870
rect 2662 865 2663 869
rect 2667 865 2668 869
rect 2662 864 2668 865
rect 2846 869 2852 870
rect 2846 865 2847 869
rect 2851 865 2852 869
rect 2846 864 2852 865
rect 3038 869 3044 870
rect 3038 865 3039 869
rect 3043 865 3044 869
rect 3038 864 3044 865
rect 3238 869 3244 870
rect 3238 865 3239 869
rect 3243 865 3244 869
rect 3238 864 3244 865
rect 3438 869 3444 870
rect 3438 865 3439 869
rect 3443 865 3444 869
rect 3438 864 3444 865
rect 1630 860 1636 861
rect 1862 856 1868 857
rect 3574 856 3580 857
rect 110 852 116 853
rect 1822 852 1828 853
rect 110 848 111 852
rect 115 848 116 852
rect 991 851 997 852
rect 991 850 992 851
rect 981 848 992 850
rect 110 847 116 848
rect 410 847 416 848
rect 410 843 411 847
rect 415 846 416 847
rect 502 847 508 848
rect 415 844 449 846
rect 415 843 416 844
rect 410 842 416 843
rect 502 843 503 847
rect 507 846 508 847
rect 634 847 640 848
rect 507 844 553 846
rect 507 843 508 844
rect 502 842 508 843
rect 634 843 635 847
rect 639 846 640 847
rect 718 847 724 848
rect 639 844 665 846
rect 639 843 640 844
rect 634 842 640 843
rect 718 843 719 847
rect 723 846 724 847
rect 991 847 992 848
rect 996 847 997 851
rect 1822 848 1823 852
rect 1827 848 1828 852
rect 1862 852 1863 856
rect 1867 852 1868 856
rect 2263 855 2269 856
rect 2263 854 2264 855
rect 2221 852 2264 854
rect 1862 851 1868 852
rect 1966 851 1972 852
rect 991 846 997 847
rect 1026 847 1032 848
rect 723 844 801 846
rect 723 843 724 844
rect 718 842 724 843
rect 1026 843 1027 847
rect 1031 846 1032 847
rect 1194 847 1200 848
rect 1031 844 1105 846
rect 1031 843 1032 844
rect 1026 842 1032 843
rect 1194 843 1195 847
rect 1199 846 1200 847
rect 1518 847 1524 848
rect 1822 847 1828 848
rect 1966 847 1967 851
rect 1971 850 1972 851
rect 2263 851 2264 852
rect 2268 851 2269 855
rect 2382 855 2388 856
rect 2382 854 2383 855
rect 2373 852 2383 854
rect 2263 850 2269 851
rect 2382 851 2383 852
rect 2387 851 2388 855
rect 3159 855 3165 856
rect 3159 854 3160 855
rect 3093 852 3160 854
rect 2382 850 2388 851
rect 2390 851 2396 852
rect 1971 848 2033 850
rect 1971 847 1972 848
rect 1199 844 1281 846
rect 1199 843 1200 844
rect 1194 842 1200 843
rect 1518 843 1519 847
rect 1523 846 1524 847
rect 1966 846 1972 847
rect 2390 847 2391 851
rect 2395 850 2396 851
rect 2759 851 2765 852
rect 2395 848 2505 850
rect 2395 847 2396 848
rect 2390 846 2396 847
rect 2759 847 2760 851
rect 2764 850 2765 851
rect 3159 851 3160 852
rect 3164 851 3165 855
rect 3574 852 3575 856
rect 3579 852 3580 856
rect 3574 851 3580 852
rect 3159 850 3165 851
rect 2764 848 2865 850
rect 2764 847 2765 848
rect 2759 846 2765 847
rect 1523 844 1649 846
rect 1523 843 1524 844
rect 1518 842 1524 843
rect 1862 839 1868 840
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 430 835 436 836
rect 430 834 431 835
rect 393 832 431 834
rect 110 830 116 831
rect 430 831 431 832
rect 435 831 436 835
rect 430 830 436 831
rect 1822 835 1828 836
rect 1822 831 1823 835
rect 1827 831 1828 835
rect 1862 835 1863 839
rect 1867 835 1868 839
rect 1862 834 1868 835
rect 2662 839 2668 840
rect 2662 835 2663 839
rect 2667 838 2668 839
rect 3514 839 3520 840
rect 3514 838 3515 839
rect 2667 836 2673 838
rect 3100 836 3249 838
rect 3489 836 3515 838
rect 2667 835 2668 836
rect 2662 834 2668 835
rect 1822 830 1828 831
rect 1886 829 1892 830
rect 334 825 340 826
rect 334 821 335 825
rect 339 821 340 825
rect 334 820 340 821
rect 422 825 428 826
rect 422 821 423 825
rect 427 821 428 825
rect 422 820 428 821
rect 526 825 532 826
rect 526 821 527 825
rect 531 821 532 825
rect 526 820 532 821
rect 638 825 644 826
rect 638 821 639 825
rect 643 821 644 825
rect 638 820 644 821
rect 774 825 780 826
rect 774 821 775 825
rect 779 821 780 825
rect 774 820 780 821
rect 918 825 924 826
rect 918 821 919 825
rect 923 821 924 825
rect 918 820 924 821
rect 1078 825 1084 826
rect 1078 821 1079 825
rect 1083 821 1084 825
rect 1078 820 1084 821
rect 1254 825 1260 826
rect 1254 821 1255 825
rect 1259 821 1260 825
rect 1254 820 1260 821
rect 1438 825 1444 826
rect 1438 821 1439 825
rect 1443 821 1444 825
rect 1438 820 1444 821
rect 1622 825 1628 826
rect 1622 821 1623 825
rect 1627 821 1628 825
rect 1886 825 1887 829
rect 1891 825 1892 829
rect 1886 824 1892 825
rect 2006 829 2012 830
rect 2006 825 2007 829
rect 2011 825 2012 829
rect 2006 824 2012 825
rect 2158 829 2164 830
rect 2158 825 2159 829
rect 2163 825 2164 829
rect 2158 824 2164 825
rect 2310 829 2316 830
rect 2310 825 2311 829
rect 2315 825 2316 829
rect 2310 824 2316 825
rect 2478 829 2484 830
rect 2478 825 2479 829
rect 2483 825 2484 829
rect 2478 824 2484 825
rect 2654 829 2660 830
rect 2654 825 2655 829
rect 2659 825 2660 829
rect 2654 824 2660 825
rect 2838 829 2844 830
rect 2838 825 2839 829
rect 2843 825 2844 829
rect 2838 824 2844 825
rect 3030 829 3036 830
rect 3030 825 3031 829
rect 3035 825 3036 829
rect 3030 824 3036 825
rect 1622 820 1628 821
rect 1926 823 1932 824
rect 1478 819 1484 820
rect 1478 815 1479 819
rect 1483 818 1484 819
rect 1487 819 1493 820
rect 1487 818 1488 819
rect 1483 816 1488 818
rect 1483 815 1484 816
rect 1478 814 1484 815
rect 1487 815 1488 816
rect 1492 815 1493 819
rect 1926 819 1927 823
rect 1931 822 1932 823
rect 1935 823 1941 824
rect 1935 822 1936 823
rect 1931 820 1936 822
rect 1931 819 1932 820
rect 1926 818 1932 819
rect 1935 819 1936 820
rect 1940 819 1941 823
rect 1935 818 1941 819
rect 2878 823 2884 824
rect 2878 819 2879 823
rect 2883 822 2884 823
rect 3100 822 3102 836
rect 3514 835 3515 836
rect 3519 835 3520 839
rect 3514 834 3520 835
rect 3574 839 3580 840
rect 3574 835 3575 839
rect 3579 835 3580 839
rect 3574 834 3580 835
rect 3230 829 3236 830
rect 3230 825 3231 829
rect 3235 825 3236 829
rect 3230 824 3236 825
rect 3430 829 3436 830
rect 3430 825 3431 829
rect 3435 825 3436 829
rect 3430 824 3436 825
rect 2883 820 3102 822
rect 2883 819 2884 820
rect 2878 818 2884 819
rect 1487 814 1493 815
rect 1886 807 1892 808
rect 286 803 292 804
rect 286 799 287 803
rect 291 799 292 803
rect 286 798 292 799
rect 406 803 412 804
rect 406 799 407 803
rect 411 799 412 803
rect 406 798 412 799
rect 534 803 540 804
rect 534 799 535 803
rect 539 799 540 803
rect 534 798 540 799
rect 678 803 684 804
rect 678 799 679 803
rect 683 799 684 803
rect 678 798 684 799
rect 822 803 828 804
rect 822 799 823 803
rect 827 799 828 803
rect 822 798 828 799
rect 974 803 980 804
rect 974 799 975 803
rect 979 799 980 803
rect 974 798 980 799
rect 1126 803 1132 804
rect 1126 799 1127 803
rect 1131 799 1132 803
rect 1126 798 1132 799
rect 1278 803 1284 804
rect 1278 799 1279 803
rect 1283 799 1284 803
rect 1278 798 1284 799
rect 1438 803 1444 804
rect 1438 799 1439 803
rect 1443 799 1444 803
rect 1438 798 1444 799
rect 1598 803 1604 804
rect 1598 799 1599 803
rect 1603 799 1604 803
rect 1886 803 1887 807
rect 1891 803 1892 807
rect 1886 802 1892 803
rect 1990 807 1996 808
rect 1990 803 1991 807
rect 1995 803 1996 807
rect 1990 802 1996 803
rect 2134 807 2140 808
rect 2134 803 2135 807
rect 2139 803 2140 807
rect 2134 802 2140 803
rect 2286 807 2292 808
rect 2286 803 2287 807
rect 2291 803 2292 807
rect 2286 802 2292 803
rect 2454 807 2460 808
rect 2454 803 2455 807
rect 2459 803 2460 807
rect 2454 802 2460 803
rect 2622 807 2628 808
rect 2622 803 2623 807
rect 2627 803 2628 807
rect 2622 802 2628 803
rect 2798 807 2804 808
rect 2798 803 2799 807
rect 2803 803 2804 807
rect 2798 802 2804 803
rect 2966 807 2972 808
rect 2966 803 2967 807
rect 2971 803 2972 807
rect 2966 802 2972 803
rect 3142 807 3148 808
rect 3142 803 3143 807
rect 3147 803 3148 807
rect 3142 802 3148 803
rect 3318 807 3324 808
rect 3318 803 3319 807
rect 3323 803 3324 807
rect 3318 802 3324 803
rect 3478 807 3484 808
rect 3478 803 3479 807
rect 3483 803 3484 807
rect 3478 802 3484 803
rect 1598 798 1604 799
rect 2206 799 2212 800
rect 2206 798 2207 799
rect 1862 797 1868 798
rect 474 795 480 796
rect 110 793 116 794
rect 110 789 111 793
rect 115 789 116 793
rect 474 791 475 795
rect 479 794 480 795
rect 814 795 820 796
rect 479 792 553 794
rect 479 791 480 792
rect 474 790 480 791
rect 814 791 815 795
rect 819 794 820 795
rect 1222 795 1228 796
rect 1222 794 1223 795
rect 819 792 841 794
rect 1185 792 1223 794
rect 819 791 820 792
rect 814 790 820 791
rect 1222 791 1223 792
rect 1227 791 1228 795
rect 1222 790 1228 791
rect 1518 795 1524 796
rect 1518 791 1519 795
rect 1523 794 1524 795
rect 1523 792 1617 794
rect 1822 793 1828 794
rect 1523 791 1524 792
rect 1518 790 1524 791
rect 110 788 116 789
rect 1822 789 1823 793
rect 1827 789 1828 793
rect 1862 793 1863 797
rect 1867 793 1868 797
rect 2193 796 2207 798
rect 2206 795 2207 796
rect 2211 795 2212 799
rect 3406 799 3412 800
rect 3406 798 3407 799
rect 3377 796 3407 798
rect 2206 794 2212 795
rect 3406 795 3407 796
rect 3411 795 3412 799
rect 3406 794 3412 795
rect 3574 797 3580 798
rect 1862 792 1868 793
rect 3574 793 3575 797
rect 3579 793 3580 797
rect 3574 792 3580 793
rect 1822 788 1828 789
rect 1954 783 1960 784
rect 1954 782 1955 783
rect 1862 780 1868 781
rect 1949 780 1955 782
rect 246 779 252 780
rect 110 776 116 777
rect 110 772 111 776
rect 115 772 116 776
rect 246 775 247 779
rect 251 778 252 779
rect 527 779 533 780
rect 527 778 528 779
rect 251 776 313 778
rect 469 776 528 778
rect 251 775 252 776
rect 246 774 252 775
rect 527 775 528 776
rect 532 775 533 779
rect 815 779 821 780
rect 815 778 816 779
rect 741 776 816 778
rect 527 774 533 775
rect 815 775 816 776
rect 820 775 821 779
rect 1119 779 1125 780
rect 1119 778 1120 779
rect 1037 776 1120 778
rect 815 774 821 775
rect 1119 775 1120 776
rect 1124 775 1125 779
rect 1431 779 1437 780
rect 1431 778 1432 779
rect 1341 776 1432 778
rect 1119 774 1125 775
rect 1431 775 1432 776
rect 1436 775 1437 779
rect 1591 779 1597 780
rect 1591 778 1592 779
rect 1501 776 1592 778
rect 1431 774 1437 775
rect 1591 775 1592 776
rect 1596 775 1597 779
rect 1591 774 1597 775
rect 1822 776 1828 777
rect 110 771 116 772
rect 1822 772 1823 776
rect 1827 772 1828 776
rect 1862 776 1863 780
rect 1867 776 1868 780
rect 1954 779 1955 780
rect 1959 779 1960 783
rect 2127 783 2133 784
rect 2127 782 2128 783
rect 2053 780 2128 782
rect 1954 778 1960 779
rect 2127 779 2128 780
rect 2132 779 2133 783
rect 2127 778 2133 779
rect 2202 783 2208 784
rect 2202 779 2203 783
rect 2207 782 2208 783
rect 2354 783 2360 784
rect 2207 780 2313 782
rect 2207 779 2208 780
rect 2202 778 2208 779
rect 2354 779 2355 783
rect 2359 782 2360 783
rect 2791 783 2797 784
rect 2791 782 2792 783
rect 2359 780 2481 782
rect 2685 780 2792 782
rect 2359 779 2360 780
rect 2354 778 2360 779
rect 2791 779 2792 780
rect 2796 779 2797 783
rect 2866 783 2872 784
rect 2791 778 2797 779
rect 1862 775 1868 776
rect 2860 774 2862 781
rect 2866 779 2867 783
rect 2871 782 2872 783
rect 3311 783 3317 784
rect 3311 782 3312 783
rect 2871 780 2993 782
rect 3205 780 3312 782
rect 2871 779 2872 780
rect 2866 778 2872 779
rect 3311 779 3312 780
rect 3316 779 3317 783
rect 3546 783 3552 784
rect 3546 782 3547 783
rect 3541 780 3547 782
rect 3311 778 3317 779
rect 3546 779 3547 780
rect 3551 779 3552 783
rect 3546 778 3552 779
rect 3574 780 3580 781
rect 3574 776 3575 780
rect 3579 776 3580 780
rect 2959 775 2965 776
rect 3574 775 3580 776
rect 2959 774 2960 775
rect 2860 772 2960 774
rect 1822 771 1828 772
rect 2959 771 2960 772
rect 2964 771 2965 775
rect 2959 770 2965 771
rect 1894 767 1900 768
rect 294 763 300 764
rect 294 759 295 763
rect 299 759 300 763
rect 294 758 300 759
rect 414 763 420 764
rect 414 759 415 763
rect 419 759 420 763
rect 542 763 548 764
rect 414 758 420 759
rect 474 759 480 760
rect 474 758 475 759
rect 424 756 475 758
rect 424 754 426 756
rect 474 755 475 756
rect 479 755 480 759
rect 542 759 543 763
rect 547 759 548 763
rect 542 758 548 759
rect 686 763 692 764
rect 686 759 687 763
rect 691 759 692 763
rect 686 758 692 759
rect 830 763 836 764
rect 830 759 831 763
rect 835 759 836 763
rect 830 758 836 759
rect 982 763 988 764
rect 982 759 983 763
rect 987 759 988 763
rect 982 758 988 759
rect 1134 763 1140 764
rect 1134 759 1135 763
rect 1139 759 1140 763
rect 1134 758 1140 759
rect 1286 763 1292 764
rect 1286 759 1287 763
rect 1291 759 1292 763
rect 1286 758 1292 759
rect 1446 763 1452 764
rect 1446 759 1447 763
rect 1451 759 1452 763
rect 1446 758 1452 759
rect 1606 763 1612 764
rect 1606 759 1607 763
rect 1611 759 1612 763
rect 1894 763 1895 767
rect 1899 763 1900 767
rect 1894 762 1900 763
rect 1998 767 2004 768
rect 1998 763 1999 767
rect 2003 763 2004 767
rect 1998 762 2004 763
rect 2142 767 2148 768
rect 2142 763 2143 767
rect 2147 763 2148 767
rect 2142 762 2148 763
rect 2294 767 2300 768
rect 2294 763 2295 767
rect 2299 763 2300 767
rect 2294 762 2300 763
rect 2462 767 2468 768
rect 2462 763 2463 767
rect 2467 763 2468 767
rect 2462 762 2468 763
rect 2630 767 2636 768
rect 2630 763 2631 767
rect 2635 763 2636 767
rect 2630 762 2636 763
rect 2806 767 2812 768
rect 2806 763 2807 767
rect 2811 763 2812 767
rect 2806 762 2812 763
rect 2974 767 2980 768
rect 2974 763 2975 767
rect 2979 763 2980 767
rect 2974 762 2980 763
rect 3150 767 3156 768
rect 3150 763 3151 767
rect 3155 763 3156 767
rect 3150 762 3156 763
rect 3326 767 3332 768
rect 3326 763 3327 767
rect 3331 763 3332 767
rect 3326 762 3332 763
rect 3486 767 3492 768
rect 3486 763 3487 767
rect 3491 763 3492 767
rect 3486 762 3492 763
rect 1606 758 1612 759
rect 474 754 480 755
rect 1923 755 1932 756
rect 323 753 426 754
rect 323 749 324 753
rect 328 752 426 753
rect 328 749 329 752
rect 323 748 329 749
rect 430 751 436 752
rect 430 747 431 751
rect 435 750 436 751
rect 443 751 449 752
rect 443 750 444 751
rect 435 748 444 750
rect 435 747 436 748
rect 430 746 436 747
rect 443 747 444 748
rect 448 747 449 751
rect 443 746 449 747
rect 527 751 533 752
rect 527 747 528 751
rect 532 750 533 751
rect 571 751 577 752
rect 571 750 572 751
rect 532 748 572 750
rect 532 747 533 748
rect 527 746 533 747
rect 571 747 572 748
rect 576 747 577 751
rect 571 746 577 747
rect 706 751 712 752
rect 706 747 707 751
rect 711 750 712 751
rect 715 751 721 752
rect 715 750 716 751
rect 711 748 716 750
rect 711 747 712 748
rect 706 746 712 747
rect 715 747 716 748
rect 720 747 721 751
rect 715 746 721 747
rect 815 751 821 752
rect 815 747 816 751
rect 820 750 821 751
rect 859 751 865 752
rect 859 750 860 751
rect 820 748 860 750
rect 820 747 821 748
rect 815 746 821 747
rect 859 747 860 748
rect 864 747 865 751
rect 859 746 865 747
rect 999 751 1005 752
rect 999 747 1000 751
rect 1004 750 1005 751
rect 1011 751 1017 752
rect 1011 750 1012 751
rect 1004 748 1012 750
rect 1004 747 1005 748
rect 999 746 1005 747
rect 1011 747 1012 748
rect 1016 747 1017 751
rect 1011 746 1017 747
rect 1119 751 1125 752
rect 1119 747 1120 751
rect 1124 750 1125 751
rect 1163 751 1169 752
rect 1163 750 1164 751
rect 1124 748 1164 750
rect 1124 747 1125 748
rect 1119 746 1125 747
rect 1163 747 1164 748
rect 1168 747 1169 751
rect 1163 746 1169 747
rect 1314 751 1321 752
rect 1314 747 1315 751
rect 1320 747 1321 751
rect 1314 746 1321 747
rect 1475 751 1484 752
rect 1475 747 1476 751
rect 1483 747 1484 751
rect 1475 746 1484 747
rect 1591 751 1597 752
rect 1591 747 1592 751
rect 1596 750 1597 751
rect 1635 751 1641 752
rect 1635 750 1636 751
rect 1596 748 1636 750
rect 1596 747 1597 748
rect 1591 746 1597 747
rect 1635 747 1636 748
rect 1640 747 1641 751
rect 1923 751 1924 755
rect 1931 751 1932 755
rect 1923 750 1932 751
rect 2027 755 2033 756
rect 2027 751 2028 755
rect 2032 754 2033 755
rect 2127 755 2133 756
rect 2032 752 2122 754
rect 2032 751 2033 752
rect 2027 750 2033 751
rect 1635 746 1641 747
rect 2120 746 2122 752
rect 2127 751 2128 755
rect 2132 754 2133 755
rect 2171 755 2177 756
rect 2171 754 2172 755
rect 2132 752 2172 754
rect 2132 751 2133 752
rect 2127 750 2133 751
rect 2171 751 2172 752
rect 2176 751 2177 755
rect 2171 750 2177 751
rect 2323 755 2329 756
rect 2323 751 2324 755
rect 2328 754 2329 755
rect 2354 755 2360 756
rect 2354 754 2355 755
rect 2328 752 2355 754
rect 2328 751 2329 752
rect 2323 750 2329 751
rect 2354 751 2355 752
rect 2359 751 2360 755
rect 2354 750 2360 751
rect 2491 755 2497 756
rect 2491 751 2492 755
rect 2496 754 2497 755
rect 2506 755 2512 756
rect 2506 754 2507 755
rect 2496 752 2507 754
rect 2496 751 2497 752
rect 2491 750 2497 751
rect 2506 751 2507 752
rect 2511 751 2512 755
rect 2506 750 2512 751
rect 2659 755 2668 756
rect 2659 751 2660 755
rect 2667 751 2668 755
rect 2659 750 2668 751
rect 2791 755 2797 756
rect 2791 751 2792 755
rect 2796 754 2797 755
rect 2835 755 2841 756
rect 2835 754 2836 755
rect 2796 752 2836 754
rect 2796 751 2797 752
rect 2791 750 2797 751
rect 2835 751 2836 752
rect 2840 751 2841 755
rect 2835 750 2841 751
rect 2959 755 2965 756
rect 2959 751 2960 755
rect 2964 754 2965 755
rect 3003 755 3009 756
rect 3003 754 3004 755
rect 2964 752 3004 754
rect 2964 751 2965 752
rect 2959 750 2965 751
rect 3003 751 3004 752
rect 3008 751 3009 755
rect 3003 750 3009 751
rect 3179 755 3185 756
rect 3179 751 3180 755
rect 3184 754 3185 755
rect 3234 755 3240 756
rect 3234 754 3235 755
rect 3184 752 3235 754
rect 3184 751 3185 752
rect 3179 750 3185 751
rect 3234 751 3235 752
rect 3239 751 3240 755
rect 3234 750 3240 751
rect 3311 755 3317 756
rect 3311 751 3312 755
rect 3316 754 3317 755
rect 3355 755 3361 756
rect 3355 754 3356 755
rect 3316 752 3356 754
rect 3316 751 3317 752
rect 3311 750 3317 751
rect 3355 751 3356 752
rect 3360 751 3361 755
rect 3355 750 3361 751
rect 3514 755 3521 756
rect 3514 751 3515 755
rect 3520 751 3521 755
rect 3514 750 3521 751
rect 2202 747 2208 748
rect 2202 746 2203 747
rect 2120 744 2203 746
rect 1162 743 1168 744
rect 1162 742 1163 743
rect 964 740 1163 742
rect 964 738 966 740
rect 1162 739 1163 740
rect 1167 739 1168 743
rect 2202 743 2203 744
rect 2207 743 2208 747
rect 2202 742 2208 743
rect 1162 738 1168 739
rect 1923 739 1929 740
rect 963 737 969 738
rect 243 735 252 736
rect 243 731 244 735
rect 251 731 252 735
rect 243 730 252 731
rect 326 735 332 736
rect 326 731 327 735
rect 331 734 332 735
rect 387 735 393 736
rect 387 734 388 735
rect 331 732 388 734
rect 331 731 332 732
rect 326 730 332 731
rect 387 731 388 732
rect 392 731 393 735
rect 387 730 393 731
rect 447 735 453 736
rect 447 731 448 735
rect 452 734 453 735
rect 531 735 537 736
rect 531 734 532 735
rect 452 732 532 734
rect 452 731 453 732
rect 447 730 453 731
rect 531 731 532 732
rect 536 731 537 735
rect 531 730 537 731
rect 675 735 681 736
rect 675 731 676 735
rect 680 734 681 735
rect 738 735 744 736
rect 738 734 739 735
rect 680 732 739 734
rect 680 731 681 732
rect 675 730 681 731
rect 738 731 739 732
rect 743 731 744 735
rect 738 730 744 731
rect 819 735 825 736
rect 819 731 820 735
rect 824 734 825 735
rect 842 735 848 736
rect 842 734 843 735
rect 824 732 843 734
rect 824 731 825 732
rect 819 730 825 731
rect 842 731 843 732
rect 847 731 848 735
rect 963 733 964 737
rect 968 733 969 737
rect 963 732 969 733
rect 1115 735 1121 736
rect 842 730 848 731
rect 1115 731 1116 735
rect 1120 734 1121 735
rect 1142 735 1148 736
rect 1142 734 1143 735
rect 1120 732 1143 734
rect 1120 731 1121 732
rect 1115 730 1121 731
rect 1142 731 1143 732
rect 1147 731 1148 735
rect 1142 730 1148 731
rect 1231 735 1237 736
rect 1231 731 1232 735
rect 1236 734 1237 735
rect 1275 735 1281 736
rect 1275 734 1276 735
rect 1236 732 1276 734
rect 1236 731 1237 732
rect 1231 730 1237 731
rect 1275 731 1276 732
rect 1280 731 1281 735
rect 1275 730 1281 731
rect 1431 735 1437 736
rect 1431 731 1432 735
rect 1436 734 1437 735
rect 1443 735 1449 736
rect 1443 734 1444 735
rect 1436 732 1444 734
rect 1436 731 1437 732
rect 1431 730 1437 731
rect 1443 731 1444 732
rect 1448 731 1449 735
rect 1443 730 1449 731
rect 1519 735 1525 736
rect 1519 731 1520 735
rect 1524 734 1525 735
rect 1611 735 1617 736
rect 1611 734 1612 735
rect 1524 732 1612 734
rect 1524 731 1525 732
rect 1519 730 1525 731
rect 1611 731 1612 732
rect 1616 731 1617 735
rect 1611 730 1617 731
rect 1763 735 1769 736
rect 1763 731 1764 735
rect 1768 734 1769 735
rect 1870 735 1876 736
rect 1870 734 1871 735
rect 1768 732 1871 734
rect 1768 731 1769 732
rect 1763 730 1769 731
rect 1870 731 1871 732
rect 1875 731 1876 735
rect 1923 735 1924 739
rect 1928 738 1929 739
rect 1954 739 1960 740
rect 1954 738 1955 739
rect 1928 736 1955 738
rect 1928 735 1929 736
rect 1923 734 1929 735
rect 1954 735 1955 736
rect 1959 735 1960 739
rect 1954 734 1960 735
rect 2091 739 2100 740
rect 2091 735 2092 739
rect 2099 735 2100 739
rect 2091 734 2100 735
rect 2175 739 2181 740
rect 2175 735 2176 739
rect 2180 738 2181 739
rect 2283 739 2289 740
rect 2283 738 2284 739
rect 2180 736 2284 738
rect 2180 735 2181 736
rect 2175 734 2181 735
rect 2283 735 2284 736
rect 2288 735 2289 739
rect 2283 734 2289 735
rect 2367 739 2373 740
rect 2367 735 2368 739
rect 2372 738 2373 739
rect 2475 739 2481 740
rect 2475 738 2476 739
rect 2372 736 2476 738
rect 2372 735 2373 736
rect 2367 734 2373 735
rect 2475 735 2476 736
rect 2480 735 2481 739
rect 2475 734 2481 735
rect 2667 739 2673 740
rect 2667 735 2668 739
rect 2672 738 2673 739
rect 2730 739 2736 740
rect 2730 738 2731 739
rect 2672 736 2731 738
rect 2672 735 2673 736
rect 2667 734 2673 735
rect 2730 735 2731 736
rect 2735 735 2736 739
rect 2730 734 2736 735
rect 2851 739 2857 740
rect 2851 735 2852 739
rect 2856 738 2857 739
rect 2866 739 2872 740
rect 2866 738 2867 739
rect 2856 736 2867 738
rect 2856 735 2857 736
rect 2851 734 2857 735
rect 2866 735 2867 736
rect 2871 735 2872 739
rect 2866 734 2872 735
rect 3027 739 3033 740
rect 3027 735 3028 739
rect 3032 738 3033 739
rect 3058 739 3064 740
rect 3058 738 3059 739
rect 3032 736 3059 738
rect 3032 735 3033 736
rect 3027 734 3033 735
rect 3058 735 3059 736
rect 3063 735 3064 739
rect 3058 734 3064 735
rect 3103 739 3109 740
rect 3103 735 3104 739
rect 3108 738 3109 739
rect 3195 739 3201 740
rect 3195 738 3196 739
rect 3108 736 3196 738
rect 3108 735 3109 736
rect 3103 734 3109 735
rect 3195 735 3196 736
rect 3200 735 3201 739
rect 3195 734 3201 735
rect 3226 739 3232 740
rect 3226 735 3227 739
rect 3231 738 3232 739
rect 3363 739 3369 740
rect 3363 738 3364 739
rect 3231 736 3364 738
rect 3231 735 3232 736
rect 3226 734 3232 735
rect 3363 735 3364 736
rect 3368 735 3369 739
rect 3363 734 3369 735
rect 3515 739 3521 740
rect 3515 735 3516 739
rect 3520 738 3521 739
rect 3546 739 3552 740
rect 3546 738 3547 739
rect 3520 736 3547 738
rect 3520 735 3521 736
rect 3515 734 3521 735
rect 3546 735 3547 736
rect 3551 735 3552 739
rect 3546 734 3552 735
rect 1870 730 1876 731
rect 1894 729 1900 730
rect 214 725 220 726
rect 214 721 215 725
rect 219 721 220 725
rect 214 720 220 721
rect 358 725 364 726
rect 358 721 359 725
rect 363 721 364 725
rect 358 720 364 721
rect 502 725 508 726
rect 502 721 503 725
rect 507 721 508 725
rect 502 720 508 721
rect 646 725 652 726
rect 646 721 647 725
rect 651 721 652 725
rect 646 720 652 721
rect 790 725 796 726
rect 790 721 791 725
rect 795 721 796 725
rect 790 720 796 721
rect 934 725 940 726
rect 934 721 935 725
rect 939 721 940 725
rect 934 720 940 721
rect 1086 725 1092 726
rect 1086 721 1087 725
rect 1091 721 1092 725
rect 1086 720 1092 721
rect 1246 725 1252 726
rect 1246 721 1247 725
rect 1251 721 1252 725
rect 1246 720 1252 721
rect 1414 725 1420 726
rect 1414 721 1415 725
rect 1419 721 1420 725
rect 1414 720 1420 721
rect 1582 725 1588 726
rect 1582 721 1583 725
rect 1587 721 1588 725
rect 1582 720 1588 721
rect 1734 725 1740 726
rect 1734 721 1735 725
rect 1739 721 1740 725
rect 1894 725 1895 729
rect 1899 725 1900 729
rect 1894 724 1900 725
rect 2062 729 2068 730
rect 2062 725 2063 729
rect 2067 725 2068 729
rect 2062 724 2068 725
rect 2254 729 2260 730
rect 2254 725 2255 729
rect 2259 725 2260 729
rect 2254 724 2260 725
rect 2446 729 2452 730
rect 2446 725 2447 729
rect 2451 725 2452 729
rect 2446 724 2452 725
rect 2638 729 2644 730
rect 2638 725 2639 729
rect 2643 725 2644 729
rect 2638 724 2644 725
rect 2822 729 2828 730
rect 2822 725 2823 729
rect 2827 725 2828 729
rect 2822 724 2828 725
rect 2998 729 3004 730
rect 2998 725 2999 729
rect 3003 725 3004 729
rect 2998 724 3004 725
rect 3166 729 3172 730
rect 3166 725 3167 729
rect 3171 725 3172 729
rect 3166 724 3172 725
rect 3334 729 3340 730
rect 3334 725 3335 729
rect 3339 725 3340 729
rect 3334 724 3340 725
rect 3486 729 3492 730
rect 3486 725 3487 729
rect 3491 725 3492 729
rect 3486 724 3492 725
rect 1734 720 1740 721
rect 1862 716 1868 717
rect 3574 716 3580 717
rect 110 712 116 713
rect 1822 712 1828 713
rect 110 708 111 712
rect 115 708 116 712
rect 326 711 332 712
rect 326 710 327 711
rect 269 708 327 710
rect 110 707 116 708
rect 326 707 327 708
rect 331 707 332 711
rect 447 711 453 712
rect 447 710 448 711
rect 413 708 448 710
rect 326 706 332 707
rect 447 707 448 708
rect 452 707 453 711
rect 706 711 712 712
rect 706 710 707 711
rect 701 708 707 710
rect 447 706 453 707
rect 706 707 707 708
rect 711 707 712 711
rect 999 711 1005 712
rect 999 710 1000 711
rect 989 708 1000 710
rect 706 706 712 707
rect 738 707 744 708
rect 738 703 739 707
rect 743 706 744 707
rect 999 707 1000 708
rect 1004 707 1005 711
rect 1231 711 1237 712
rect 1231 710 1232 711
rect 1141 708 1232 710
rect 999 706 1005 707
rect 1231 707 1232 708
rect 1236 707 1237 711
rect 1519 711 1525 712
rect 1519 710 1520 711
rect 1469 708 1520 710
rect 1231 706 1237 707
rect 1519 707 1520 708
rect 1524 707 1525 711
rect 1822 708 1823 712
rect 1827 708 1828 712
rect 1862 712 1863 716
rect 1867 712 1868 716
rect 2175 715 2181 716
rect 2175 714 2176 715
rect 2117 712 2176 714
rect 1862 711 1868 712
rect 1870 711 1876 712
rect 1822 707 1828 708
rect 1870 707 1871 711
rect 1875 710 1876 711
rect 2175 711 2176 712
rect 2180 711 2181 715
rect 2367 715 2373 716
rect 2367 714 2368 715
rect 2309 712 2368 714
rect 2175 710 2181 711
rect 2367 711 2368 712
rect 2372 711 2373 715
rect 2506 715 2512 716
rect 2506 714 2507 715
rect 2501 712 2507 714
rect 2367 710 2373 711
rect 2506 711 2507 712
rect 2511 711 2512 715
rect 3103 715 3109 716
rect 3103 714 3104 715
rect 3053 712 3104 714
rect 2506 710 2512 711
rect 2730 711 2736 712
rect 1875 708 1913 710
rect 1875 707 1876 708
rect 1519 706 1525 707
rect 1870 706 1876 707
rect 2730 707 2731 711
rect 2735 710 2736 711
rect 3103 711 3104 712
rect 3108 711 3109 715
rect 3226 715 3232 716
rect 3226 714 3227 715
rect 3221 712 3227 714
rect 3103 710 3109 711
rect 3226 711 3227 712
rect 3231 711 3232 715
rect 3574 712 3575 716
rect 3579 712 3580 716
rect 3226 710 3232 711
rect 3234 711 3240 712
rect 3574 711 3580 712
rect 2735 708 2841 710
rect 2735 707 2736 708
rect 2730 706 2736 707
rect 3234 707 3235 711
rect 3239 710 3240 711
rect 3239 708 3353 710
rect 3239 707 3240 708
rect 3234 706 3240 707
rect 743 704 809 706
rect 743 703 744 704
rect 738 702 744 703
rect 1862 699 1868 700
rect 110 695 116 696
rect 110 691 111 695
rect 115 691 116 695
rect 110 690 116 691
rect 502 695 508 696
rect 502 691 503 695
rect 507 694 508 695
rect 1162 695 1168 696
rect 507 692 513 694
rect 507 691 508 692
rect 502 690 508 691
rect 1162 691 1163 695
rect 1167 694 1168 695
rect 1518 695 1524 696
rect 1167 692 1257 694
rect 1167 691 1168 692
rect 1162 690 1168 691
rect 1518 691 1519 695
rect 1523 694 1524 695
rect 1822 695 1828 696
rect 1523 692 1593 694
rect 1523 691 1524 692
rect 1518 690 1524 691
rect 1822 691 1823 695
rect 1827 691 1828 695
rect 1862 695 1863 699
rect 1867 695 1868 699
rect 2706 699 2712 700
rect 2706 698 2707 699
rect 2689 696 2707 698
rect 1862 694 1868 695
rect 2706 695 2707 696
rect 2711 695 2712 699
rect 2706 694 2712 695
rect 3574 699 3580 700
rect 3574 695 3575 699
rect 3579 695 3580 699
rect 3574 694 3580 695
rect 1822 690 1828 691
rect 1886 689 1892 690
rect 206 685 212 686
rect 206 681 207 685
rect 211 681 212 685
rect 206 680 212 681
rect 350 685 356 686
rect 350 681 351 685
rect 355 681 356 685
rect 350 680 356 681
rect 494 685 500 686
rect 494 681 495 685
rect 499 681 500 685
rect 494 680 500 681
rect 638 685 644 686
rect 638 681 639 685
rect 643 681 644 685
rect 638 680 644 681
rect 782 685 788 686
rect 782 681 783 685
rect 787 681 788 685
rect 782 680 788 681
rect 926 685 932 686
rect 926 681 927 685
rect 931 681 932 685
rect 926 680 932 681
rect 1078 685 1084 686
rect 1078 681 1079 685
rect 1083 681 1084 685
rect 1078 680 1084 681
rect 1238 685 1244 686
rect 1238 681 1239 685
rect 1243 681 1244 685
rect 1238 680 1244 681
rect 1406 685 1412 686
rect 1406 681 1407 685
rect 1411 681 1412 685
rect 1406 680 1412 681
rect 1574 685 1580 686
rect 1574 681 1575 685
rect 1579 681 1580 685
rect 1574 680 1580 681
rect 1726 685 1732 686
rect 1726 681 1727 685
rect 1731 681 1732 685
rect 1886 685 1887 689
rect 1891 685 1892 689
rect 1886 684 1892 685
rect 2054 689 2060 690
rect 2054 685 2055 689
rect 2059 685 2060 689
rect 2054 684 2060 685
rect 2246 689 2252 690
rect 2246 685 2247 689
rect 2251 685 2252 689
rect 2246 684 2252 685
rect 2438 689 2444 690
rect 2438 685 2439 689
rect 2443 685 2444 689
rect 2438 684 2444 685
rect 2630 689 2636 690
rect 2630 685 2631 689
rect 2635 685 2636 689
rect 2630 684 2636 685
rect 2814 689 2820 690
rect 2814 685 2815 689
rect 2819 685 2820 689
rect 2814 684 2820 685
rect 2990 689 2996 690
rect 2990 685 2991 689
rect 2995 685 2996 689
rect 2990 684 2996 685
rect 3158 689 3164 690
rect 3158 685 3159 689
rect 3163 685 3164 689
rect 3158 684 3164 685
rect 3326 689 3332 690
rect 3326 685 3327 689
rect 3331 685 3332 689
rect 3326 684 3332 685
rect 3478 689 3484 690
rect 3478 685 3479 689
rect 3483 685 3484 689
rect 3478 684 3484 685
rect 1726 680 1732 681
rect 3518 683 3524 684
rect 1766 679 1772 680
rect 1766 675 1767 679
rect 1771 678 1772 679
rect 1775 679 1781 680
rect 1775 678 1776 679
rect 1771 676 1776 678
rect 1771 675 1772 676
rect 1766 674 1772 675
rect 1775 675 1776 676
rect 1780 675 1781 679
rect 3518 679 3519 683
rect 3523 682 3524 683
rect 3527 683 3533 684
rect 3527 682 3528 683
rect 3523 680 3528 682
rect 3523 679 3524 680
rect 3518 678 3524 679
rect 3527 679 3528 680
rect 3532 679 3533 683
rect 3527 678 3533 679
rect 1775 674 1781 675
rect 134 663 140 664
rect 134 659 135 663
rect 139 659 140 663
rect 134 658 140 659
rect 294 663 300 664
rect 294 659 295 663
rect 299 659 300 663
rect 294 658 300 659
rect 462 663 468 664
rect 462 659 463 663
rect 467 659 468 663
rect 462 658 468 659
rect 622 663 628 664
rect 622 659 623 663
rect 627 659 628 663
rect 622 658 628 659
rect 774 663 780 664
rect 774 659 775 663
rect 779 659 780 663
rect 774 658 780 659
rect 926 663 932 664
rect 926 659 927 663
rect 931 659 932 663
rect 926 658 932 659
rect 1070 663 1076 664
rect 1070 659 1071 663
rect 1075 659 1076 663
rect 1070 658 1076 659
rect 1206 663 1212 664
rect 1206 659 1207 663
rect 1211 659 1212 663
rect 1206 658 1212 659
rect 1342 663 1348 664
rect 1342 659 1343 663
rect 1347 659 1348 663
rect 1342 658 1348 659
rect 1478 663 1484 664
rect 1478 659 1479 663
rect 1483 659 1484 663
rect 1478 658 1484 659
rect 1614 663 1620 664
rect 1614 659 1615 663
rect 1619 659 1620 663
rect 1614 658 1620 659
rect 1726 663 1732 664
rect 1726 659 1727 663
rect 1731 659 1732 663
rect 1726 658 1732 659
rect 2214 663 2220 664
rect 2214 659 2215 663
rect 2219 659 2220 663
rect 2214 658 2220 659
rect 2358 663 2364 664
rect 2358 659 2359 663
rect 2363 659 2364 663
rect 2358 658 2364 659
rect 2510 663 2516 664
rect 2510 659 2511 663
rect 2515 659 2516 663
rect 2510 658 2516 659
rect 2670 663 2676 664
rect 2670 659 2671 663
rect 2675 659 2676 663
rect 2670 658 2676 659
rect 2830 663 2836 664
rect 2830 659 2831 663
rect 2835 659 2836 663
rect 2830 658 2836 659
rect 2990 663 2996 664
rect 2990 659 2991 663
rect 2995 659 2996 663
rect 2990 658 2996 659
rect 3158 663 3164 664
rect 3158 659 3159 663
rect 3163 659 3164 663
rect 3158 658 3164 659
rect 3326 663 3332 664
rect 3326 659 3327 663
rect 3331 659 3332 663
rect 3326 658 3332 659
rect 3478 663 3484 664
rect 3478 659 3479 663
rect 3483 659 3484 663
rect 3478 658 3484 659
rect 842 655 848 656
rect 842 654 843 655
rect 110 653 116 654
rect 110 649 111 653
rect 115 649 116 653
rect 833 652 843 654
rect 842 651 843 652
rect 847 651 848 655
rect 1142 655 1148 656
rect 1142 654 1143 655
rect 1129 652 1143 654
rect 842 650 848 651
rect 1142 651 1143 652
rect 1147 651 1148 655
rect 2094 655 2100 656
rect 1142 650 1148 651
rect 1822 653 1828 654
rect 110 648 116 649
rect 1822 649 1823 653
rect 1827 649 1828 653
rect 1822 648 1828 649
rect 1862 653 1868 654
rect 1862 649 1863 653
rect 1867 649 1868 653
rect 2094 651 2095 655
rect 2099 654 2100 655
rect 3058 655 3064 656
rect 3058 654 3059 655
rect 2099 652 2233 654
rect 3049 652 3059 654
rect 2099 651 2100 652
rect 2094 650 2100 651
rect 3058 651 3059 652
rect 3063 651 3064 655
rect 3058 650 3064 651
rect 3574 653 3580 654
rect 1862 648 1868 649
rect 3574 649 3575 653
rect 3579 649 3580 653
rect 3574 648 3580 649
rect 202 639 208 640
rect 110 636 116 637
rect 110 632 111 636
rect 115 632 116 636
rect 110 631 116 632
rect 197 632 199 638
rect 202 635 203 639
rect 207 638 208 639
rect 362 639 368 640
rect 207 636 321 638
rect 207 635 208 636
rect 202 634 208 635
rect 362 635 363 639
rect 367 638 368 639
rect 767 639 773 640
rect 767 638 768 639
rect 367 636 489 638
rect 685 636 768 638
rect 367 635 368 636
rect 362 634 368 635
rect 767 635 768 636
rect 772 635 773 639
rect 1023 639 1029 640
rect 1023 638 1024 639
rect 989 636 1024 638
rect 767 634 773 635
rect 1023 635 1024 636
rect 1028 635 1029 639
rect 1335 639 1341 640
rect 1335 638 1336 639
rect 1269 636 1336 638
rect 1023 634 1029 635
rect 1335 635 1336 636
rect 1340 635 1341 639
rect 1410 639 1416 640
rect 1410 638 1411 639
rect 1405 636 1411 638
rect 1335 634 1341 635
rect 1410 635 1411 636
rect 1415 635 1416 639
rect 1410 634 1416 635
rect 1418 639 1424 640
rect 1418 635 1419 639
rect 1423 638 1424 639
rect 1590 639 1596 640
rect 1423 636 1505 638
rect 1423 635 1424 636
rect 1418 634 1424 635
rect 1590 635 1591 639
rect 1595 638 1596 639
rect 1682 639 1688 640
rect 1595 636 1641 638
rect 1595 635 1596 636
rect 1590 634 1596 635
rect 1682 635 1683 639
rect 1687 638 1688 639
rect 2282 639 2288 640
rect 1687 636 1753 638
rect 1822 636 1828 637
rect 1687 635 1688 636
rect 1682 634 1688 635
rect 1822 632 1823 636
rect 1827 632 1828 636
rect 197 631 205 632
rect 1822 631 1828 632
rect 1862 636 1868 637
rect 1862 632 1863 636
rect 1867 632 1868 636
rect 2282 635 2283 639
rect 2287 638 2288 639
rect 2426 639 2432 640
rect 2287 636 2385 638
rect 2287 635 2288 636
rect 2282 634 2288 635
rect 2426 635 2427 639
rect 2431 638 2432 639
rect 2822 639 2828 640
rect 2822 638 2823 639
rect 2431 636 2537 638
rect 2733 636 2823 638
rect 2431 635 2432 636
rect 2426 634 2432 635
rect 2822 635 2823 636
rect 2827 635 2828 639
rect 2982 639 2988 640
rect 2982 638 2983 639
rect 2893 636 2983 638
rect 2822 634 2828 635
rect 2982 635 2983 636
rect 2987 635 2988 639
rect 2982 634 2988 635
rect 3058 639 3064 640
rect 3058 635 3059 639
rect 3063 638 3064 639
rect 3226 639 3232 640
rect 3063 636 3185 638
rect 3063 635 3064 636
rect 3058 634 3064 635
rect 3226 635 3227 639
rect 3231 638 3232 639
rect 3546 639 3552 640
rect 3546 638 3547 639
rect 3231 636 3353 638
rect 3541 636 3547 638
rect 3231 635 3232 636
rect 3226 634 3232 635
rect 3546 635 3547 636
rect 3551 635 3552 639
rect 3546 634 3552 635
rect 3574 636 3580 637
rect 1862 631 1868 632
rect 3574 632 3575 636
rect 3579 632 3580 636
rect 3574 631 3580 632
rect 197 628 200 631
rect 199 627 200 628
rect 204 627 205 631
rect 199 626 205 627
rect 142 623 148 624
rect 142 619 143 623
rect 147 619 148 623
rect 142 618 148 619
rect 302 623 308 624
rect 302 619 303 623
rect 307 619 308 623
rect 302 618 308 619
rect 470 623 476 624
rect 470 619 471 623
rect 475 619 476 623
rect 470 618 476 619
rect 630 623 636 624
rect 630 619 631 623
rect 635 619 636 623
rect 630 618 636 619
rect 782 623 788 624
rect 782 619 783 623
rect 787 619 788 623
rect 782 618 788 619
rect 934 623 940 624
rect 934 619 935 623
rect 939 619 940 623
rect 934 618 940 619
rect 1078 623 1084 624
rect 1078 619 1079 623
rect 1083 619 1084 623
rect 1078 618 1084 619
rect 1214 623 1220 624
rect 1214 619 1215 623
rect 1219 619 1220 623
rect 1214 618 1220 619
rect 1350 623 1356 624
rect 1350 619 1351 623
rect 1355 619 1356 623
rect 1486 623 1492 624
rect 1350 618 1356 619
rect 1418 619 1424 620
rect 1418 618 1419 619
rect 1244 616 1346 618
rect 1244 614 1246 616
rect 1344 614 1346 616
rect 1360 616 1419 618
rect 1360 614 1362 616
rect 1418 615 1419 616
rect 1423 615 1424 619
rect 1486 619 1487 623
rect 1491 619 1492 623
rect 1486 618 1492 619
rect 1622 623 1628 624
rect 1622 619 1623 623
rect 1627 619 1628 623
rect 1622 618 1628 619
rect 1734 623 1740 624
rect 1734 619 1735 623
rect 1739 619 1740 623
rect 1734 618 1740 619
rect 2222 623 2228 624
rect 2222 619 2223 623
rect 2227 619 2228 623
rect 2222 618 2228 619
rect 2366 623 2372 624
rect 2366 619 2367 623
rect 2371 619 2372 623
rect 2366 618 2372 619
rect 2518 623 2524 624
rect 2518 619 2519 623
rect 2523 619 2524 623
rect 2518 618 2524 619
rect 2678 623 2684 624
rect 2678 619 2679 623
rect 2683 619 2684 623
rect 2678 618 2684 619
rect 2838 623 2844 624
rect 2838 619 2839 623
rect 2843 619 2844 623
rect 2838 618 2844 619
rect 2998 623 3004 624
rect 2998 619 2999 623
rect 3003 619 3004 623
rect 2998 618 3004 619
rect 3166 623 3172 624
rect 3166 619 3167 623
rect 3171 619 3172 623
rect 3166 618 3172 619
rect 3334 623 3340 624
rect 3334 619 3335 623
rect 3339 619 3340 623
rect 3334 618 3340 619
rect 3486 623 3492 624
rect 3486 619 3487 623
rect 3491 619 3492 623
rect 3486 618 3492 619
rect 1418 614 1424 615
rect 1243 613 1249 614
rect 171 611 177 612
rect 171 607 172 611
rect 176 610 177 611
rect 202 611 208 612
rect 202 610 203 611
rect 176 608 203 610
rect 176 607 177 608
rect 171 606 177 607
rect 202 607 203 608
rect 207 607 208 611
rect 202 606 208 607
rect 331 611 337 612
rect 331 607 332 611
rect 336 610 337 611
rect 362 611 368 612
rect 362 610 363 611
rect 336 608 363 610
rect 336 607 337 608
rect 331 606 337 607
rect 362 607 363 608
rect 367 607 368 611
rect 362 606 368 607
rect 499 611 508 612
rect 499 607 500 611
rect 507 607 508 611
rect 499 606 508 607
rect 659 611 668 612
rect 659 607 660 611
rect 667 607 668 611
rect 659 606 668 607
rect 767 611 773 612
rect 767 607 768 611
rect 772 610 773 611
rect 811 611 817 612
rect 811 610 812 611
rect 772 608 812 610
rect 772 607 773 608
rect 767 606 773 607
rect 811 607 812 608
rect 816 607 817 611
rect 811 606 817 607
rect 963 611 969 612
rect 963 607 964 611
rect 968 610 969 611
rect 999 611 1005 612
rect 999 610 1000 611
rect 968 608 1000 610
rect 968 607 969 608
rect 963 606 969 607
rect 999 607 1000 608
rect 1004 607 1005 611
rect 999 606 1005 607
rect 1023 611 1029 612
rect 1023 607 1024 611
rect 1028 610 1029 611
rect 1107 611 1113 612
rect 1107 610 1108 611
rect 1028 608 1108 610
rect 1028 607 1029 608
rect 1023 606 1029 607
rect 1107 607 1108 608
rect 1112 607 1113 611
rect 1243 609 1244 613
rect 1248 609 1249 613
rect 1344 612 1362 614
rect 1243 608 1249 609
rect 1335 611 1341 612
rect 1107 606 1113 607
rect 1335 607 1336 611
rect 1340 610 1341 611
rect 1379 611 1385 612
rect 1379 610 1380 611
rect 1340 608 1380 610
rect 1340 607 1341 608
rect 1335 606 1341 607
rect 1379 607 1380 608
rect 1384 607 1385 611
rect 1379 606 1385 607
rect 1515 611 1524 612
rect 1515 607 1516 611
rect 1523 607 1524 611
rect 1515 606 1524 607
rect 1651 611 1657 612
rect 1651 607 1652 611
rect 1656 610 1657 611
rect 1682 611 1688 612
rect 1682 610 1683 611
rect 1656 608 1683 610
rect 1656 607 1657 608
rect 1651 606 1657 607
rect 1682 607 1683 608
rect 1687 607 1688 611
rect 1682 606 1688 607
rect 1763 611 1772 612
rect 1763 607 1764 611
rect 1771 607 1772 611
rect 1763 606 1772 607
rect 2251 611 2257 612
rect 2251 607 2252 611
rect 2256 610 2257 611
rect 2282 611 2288 612
rect 2282 610 2283 611
rect 2256 608 2283 610
rect 2256 607 2257 608
rect 2251 606 2257 607
rect 2282 607 2283 608
rect 2287 607 2288 611
rect 2282 606 2288 607
rect 2395 611 2401 612
rect 2395 607 2396 611
rect 2400 610 2401 611
rect 2426 611 2432 612
rect 2426 610 2427 611
rect 2400 608 2427 610
rect 2400 607 2401 608
rect 2395 606 2401 607
rect 2426 607 2427 608
rect 2431 607 2432 611
rect 2426 606 2432 607
rect 2535 611 2541 612
rect 2535 607 2536 611
rect 2540 610 2541 611
rect 2547 611 2553 612
rect 2547 610 2548 611
rect 2540 608 2548 610
rect 2540 607 2541 608
rect 2535 606 2541 607
rect 2547 607 2548 608
rect 2552 607 2553 611
rect 2547 606 2553 607
rect 2706 611 2713 612
rect 2706 607 2707 611
rect 2712 607 2713 611
rect 2706 606 2713 607
rect 2822 611 2828 612
rect 2822 607 2823 611
rect 2827 610 2828 611
rect 2867 611 2873 612
rect 2867 610 2868 611
rect 2827 608 2868 610
rect 2827 607 2828 608
rect 2822 606 2828 607
rect 2867 607 2868 608
rect 2872 607 2873 611
rect 2867 606 2873 607
rect 3027 611 3033 612
rect 3027 607 3028 611
rect 3032 610 3033 611
rect 3058 611 3064 612
rect 3058 610 3059 611
rect 3032 608 3059 610
rect 3032 607 3033 608
rect 3027 606 3033 607
rect 3058 607 3059 608
rect 3063 607 3064 611
rect 3058 606 3064 607
rect 3195 611 3201 612
rect 3195 607 3196 611
rect 3200 610 3201 611
rect 3226 611 3232 612
rect 3226 610 3227 611
rect 3200 608 3227 610
rect 3200 607 3201 608
rect 3195 606 3201 607
rect 3226 607 3227 608
rect 3231 607 3232 611
rect 3226 606 3232 607
rect 3363 611 3369 612
rect 3363 607 3364 611
rect 3368 610 3369 611
rect 3386 611 3392 612
rect 3386 610 3387 611
rect 3368 608 3387 610
rect 3368 607 3369 608
rect 3363 606 3369 607
rect 3386 607 3387 608
rect 3391 607 3392 611
rect 3386 606 3392 607
rect 3515 611 3524 612
rect 3515 607 3516 611
rect 3523 607 3524 611
rect 3515 606 3524 607
rect 2746 603 2752 604
rect 2746 602 2747 603
rect 2596 600 2747 602
rect 2596 598 2598 600
rect 2746 599 2747 600
rect 2751 599 2752 603
rect 2746 598 2752 599
rect 2595 597 2601 598
rect 171 595 177 596
rect 171 591 172 595
rect 176 594 177 595
rect 199 595 205 596
rect 199 594 200 595
rect 176 592 200 594
rect 176 591 177 592
rect 171 590 177 591
rect 199 591 200 592
rect 204 591 205 595
rect 199 590 205 591
rect 207 595 213 596
rect 207 591 208 595
rect 212 594 213 595
rect 331 595 337 596
rect 331 594 332 595
rect 212 592 332 594
rect 212 591 213 592
rect 207 590 213 591
rect 331 591 332 592
rect 336 591 337 595
rect 331 590 337 591
rect 415 595 421 596
rect 415 591 416 595
rect 420 594 421 595
rect 515 595 521 596
rect 515 594 516 595
rect 420 592 516 594
rect 420 591 421 592
rect 415 590 421 591
rect 515 591 516 592
rect 520 591 521 595
rect 515 590 521 591
rect 699 595 705 596
rect 699 591 700 595
rect 704 594 705 595
rect 754 595 760 596
rect 754 594 755 595
rect 704 592 755 594
rect 704 591 705 592
rect 699 590 705 591
rect 754 591 755 592
rect 759 591 760 595
rect 754 590 760 591
rect 790 595 796 596
rect 790 591 791 595
rect 795 594 796 595
rect 875 595 881 596
rect 875 594 876 595
rect 795 592 876 594
rect 795 591 796 592
rect 790 590 796 591
rect 875 591 876 592
rect 880 591 881 595
rect 875 590 881 591
rect 1038 595 1044 596
rect 1038 591 1039 595
rect 1043 594 1044 595
rect 1051 595 1057 596
rect 1051 594 1052 595
rect 1043 592 1052 594
rect 1043 591 1044 592
rect 1038 590 1044 591
rect 1051 591 1052 592
rect 1056 591 1057 595
rect 1051 590 1057 591
rect 1227 595 1233 596
rect 1227 591 1228 595
rect 1232 594 1233 595
rect 1306 595 1312 596
rect 1306 594 1307 595
rect 1232 592 1307 594
rect 1232 591 1233 592
rect 1227 590 1233 591
rect 1306 591 1307 592
rect 1311 591 1312 595
rect 1306 590 1312 591
rect 1403 595 1412 596
rect 1403 591 1404 595
rect 1411 591 1412 595
rect 1403 590 1412 591
rect 1587 595 1596 596
rect 1587 591 1588 595
rect 1595 591 1596 595
rect 1587 590 1596 591
rect 1663 595 1669 596
rect 1663 591 1664 595
rect 1668 594 1669 595
rect 1763 595 1769 596
rect 1763 594 1764 595
rect 1668 592 1764 594
rect 1668 591 1669 592
rect 1663 590 1669 591
rect 1763 591 1764 592
rect 1768 591 1769 595
rect 1763 590 1769 591
rect 2227 595 2236 596
rect 2227 591 2228 595
rect 2235 591 2236 595
rect 2227 590 2236 591
rect 2263 595 2269 596
rect 2263 591 2264 595
rect 2268 594 2269 595
rect 2315 595 2321 596
rect 2315 594 2316 595
rect 2268 592 2316 594
rect 2268 591 2269 592
rect 2263 590 2269 591
rect 2315 591 2316 592
rect 2320 591 2321 595
rect 2315 590 2321 591
rect 2351 595 2357 596
rect 2351 591 2352 595
rect 2356 594 2357 595
rect 2403 595 2409 596
rect 2403 594 2404 595
rect 2356 592 2404 594
rect 2356 591 2357 592
rect 2351 590 2357 591
rect 2403 591 2404 592
rect 2408 591 2409 595
rect 2403 590 2409 591
rect 2439 595 2445 596
rect 2439 591 2440 595
rect 2444 594 2445 595
rect 2491 595 2497 596
rect 2491 594 2492 595
rect 2444 592 2492 594
rect 2444 591 2445 592
rect 2439 590 2445 591
rect 2491 591 2492 592
rect 2496 591 2497 595
rect 2595 593 2596 597
rect 2600 593 2601 597
rect 2595 592 2601 593
rect 2639 595 2645 596
rect 2491 590 2497 591
rect 2639 591 2640 595
rect 2644 594 2645 595
rect 2707 595 2713 596
rect 2707 594 2708 595
rect 2644 592 2708 594
rect 2644 591 2645 592
rect 2639 590 2645 591
rect 2707 591 2708 592
rect 2712 591 2713 595
rect 2707 590 2713 591
rect 2843 595 2849 596
rect 2843 591 2844 595
rect 2848 594 2849 595
rect 2914 595 2920 596
rect 2914 594 2915 595
rect 2848 592 2915 594
rect 2848 591 2849 592
rect 2843 590 2849 591
rect 2914 591 2915 592
rect 2919 591 2920 595
rect 2914 590 2920 591
rect 2982 595 2988 596
rect 2982 591 2983 595
rect 2987 594 2988 595
rect 3003 595 3009 596
rect 3003 594 3004 595
rect 2987 592 3004 594
rect 2987 591 2988 592
rect 2982 590 2988 591
rect 3003 591 3004 592
rect 3008 591 3009 595
rect 3003 590 3009 591
rect 3171 595 3180 596
rect 3171 591 3172 595
rect 3179 591 3180 595
rect 3171 590 3180 591
rect 3255 595 3261 596
rect 3255 591 3256 595
rect 3260 594 3261 595
rect 3355 595 3361 596
rect 3355 594 3356 595
rect 3260 592 3356 594
rect 3260 591 3261 592
rect 3255 590 3261 591
rect 3355 591 3356 592
rect 3360 591 3361 595
rect 3355 590 3361 591
rect 3515 595 3521 596
rect 3515 591 3516 595
rect 3520 594 3521 595
rect 3546 595 3552 596
rect 3546 594 3547 595
rect 3520 592 3547 594
rect 3520 591 3521 592
rect 3515 590 3521 591
rect 3546 591 3547 592
rect 3551 591 3552 595
rect 3546 590 3552 591
rect 142 585 148 586
rect 142 581 143 585
rect 147 581 148 585
rect 142 580 148 581
rect 302 585 308 586
rect 302 581 303 585
rect 307 581 308 585
rect 302 580 308 581
rect 486 585 492 586
rect 486 581 487 585
rect 491 581 492 585
rect 486 580 492 581
rect 670 585 676 586
rect 670 581 671 585
rect 675 581 676 585
rect 670 580 676 581
rect 846 585 852 586
rect 846 581 847 585
rect 851 581 852 585
rect 846 580 852 581
rect 1022 585 1028 586
rect 1022 581 1023 585
rect 1027 581 1028 585
rect 1022 580 1028 581
rect 1198 585 1204 586
rect 1198 581 1199 585
rect 1203 581 1204 585
rect 1198 580 1204 581
rect 1374 585 1380 586
rect 1374 581 1375 585
rect 1379 581 1380 585
rect 1374 580 1380 581
rect 1558 585 1564 586
rect 1558 581 1559 585
rect 1563 581 1564 585
rect 1558 580 1564 581
rect 1734 585 1740 586
rect 1734 581 1735 585
rect 1739 581 1740 585
rect 1734 580 1740 581
rect 2198 585 2204 586
rect 2198 581 2199 585
rect 2203 581 2204 585
rect 2198 580 2204 581
rect 2286 585 2292 586
rect 2286 581 2287 585
rect 2291 581 2292 585
rect 2286 580 2292 581
rect 2374 585 2380 586
rect 2374 581 2375 585
rect 2379 581 2380 585
rect 2374 580 2380 581
rect 2462 585 2468 586
rect 2462 581 2463 585
rect 2467 581 2468 585
rect 2462 580 2468 581
rect 2566 585 2572 586
rect 2566 581 2567 585
rect 2571 581 2572 585
rect 2566 580 2572 581
rect 2678 585 2684 586
rect 2678 581 2679 585
rect 2683 581 2684 585
rect 2678 580 2684 581
rect 2814 585 2820 586
rect 2814 581 2815 585
rect 2819 581 2820 585
rect 2814 580 2820 581
rect 2974 585 2980 586
rect 2974 581 2975 585
rect 2979 581 2980 585
rect 2974 580 2980 581
rect 3142 585 3148 586
rect 3142 581 3143 585
rect 3147 581 3148 585
rect 3142 580 3148 581
rect 3326 585 3332 586
rect 3326 581 3327 585
rect 3331 581 3332 585
rect 3326 580 3332 581
rect 3486 585 3492 586
rect 3486 581 3487 585
rect 3491 581 3492 585
rect 3486 580 3492 581
rect 110 572 116 573
rect 1822 572 1828 573
rect 110 568 111 572
rect 115 568 116 572
rect 207 571 213 572
rect 207 570 208 571
rect 197 568 208 570
rect 110 567 116 568
rect 207 567 208 568
rect 212 567 213 571
rect 415 571 421 572
rect 415 570 416 571
rect 357 568 416 570
rect 207 566 213 567
rect 415 567 416 568
rect 420 567 421 571
rect 1663 571 1669 572
rect 1663 570 1664 571
rect 1613 568 1664 570
rect 415 566 421 567
rect 662 567 668 568
rect 662 563 663 567
rect 667 566 668 567
rect 754 567 760 568
rect 667 564 689 566
rect 667 563 668 564
rect 662 562 668 563
rect 754 563 755 567
rect 759 566 760 567
rect 999 567 1005 568
rect 759 564 865 566
rect 759 563 760 564
rect 754 562 760 563
rect 999 563 1000 567
rect 1004 566 1005 567
rect 1306 567 1312 568
rect 1004 564 1041 566
rect 1004 563 1005 564
rect 999 562 1005 563
rect 1306 563 1307 567
rect 1311 566 1312 567
rect 1663 567 1664 568
rect 1668 567 1669 571
rect 1822 568 1823 572
rect 1827 568 1828 572
rect 1822 567 1828 568
rect 1862 572 1868 573
rect 3574 572 3580 573
rect 1862 568 1863 572
rect 1867 568 1868 572
rect 2263 571 2269 572
rect 2263 570 2264 571
rect 2253 568 2264 570
rect 1862 567 1868 568
rect 2263 567 2264 568
rect 2268 567 2269 571
rect 2351 571 2357 572
rect 2351 570 2352 571
rect 2341 568 2352 570
rect 1663 566 1669 567
rect 2263 566 2269 567
rect 2351 567 2352 568
rect 2356 567 2357 571
rect 2439 571 2445 572
rect 2439 570 2440 571
rect 2429 568 2440 570
rect 2351 566 2357 567
rect 2439 567 2440 568
rect 2444 567 2445 571
rect 2535 571 2541 572
rect 2535 570 2536 571
rect 2517 568 2536 570
rect 2439 566 2445 567
rect 2535 567 2536 568
rect 2540 567 2541 571
rect 2639 571 2645 572
rect 2639 570 2640 571
rect 2621 568 2640 570
rect 2535 566 2541 567
rect 2639 567 2640 568
rect 2644 567 2645 571
rect 3255 571 3261 572
rect 3255 570 3256 571
rect 3197 568 3256 570
rect 2639 566 2645 567
rect 2746 567 2752 568
rect 1311 564 1393 566
rect 1311 563 1312 564
rect 1306 562 1312 563
rect 2746 563 2747 567
rect 2751 566 2752 567
rect 2914 567 2920 568
rect 2751 564 2833 566
rect 2751 563 2752 564
rect 2746 562 2752 563
rect 2914 563 2915 567
rect 2919 566 2920 567
rect 3255 567 3256 568
rect 3260 567 3261 571
rect 3386 571 3392 572
rect 3386 570 3387 571
rect 3381 568 3387 570
rect 3255 566 3261 567
rect 3386 567 3387 568
rect 3391 567 3392 571
rect 3574 568 3575 572
rect 3579 568 3580 572
rect 3574 567 3580 568
rect 3386 566 3392 567
rect 2919 564 2993 566
rect 2919 563 2920 564
rect 2914 562 2920 563
rect 110 555 116 556
rect 110 551 111 555
rect 115 551 116 555
rect 110 550 116 551
rect 1702 555 1708 556
rect 1702 551 1703 555
rect 1707 554 1708 555
rect 1822 555 1828 556
rect 1707 552 1745 554
rect 1707 551 1708 552
rect 1702 550 1708 551
rect 1822 551 1823 555
rect 1827 551 1828 555
rect 1822 550 1828 551
rect 1862 555 1868 556
rect 1862 551 1863 555
rect 1867 551 1868 555
rect 2754 555 2760 556
rect 2754 554 2755 555
rect 2729 552 2755 554
rect 1862 550 1868 551
rect 2754 551 2755 552
rect 2759 551 2760 555
rect 2754 550 2760 551
rect 3574 555 3580 556
rect 3574 551 3575 555
rect 3579 551 3580 555
rect 3574 550 3580 551
rect 134 545 140 546
rect 134 541 135 545
rect 139 541 140 545
rect 134 540 140 541
rect 294 545 300 546
rect 294 541 295 545
rect 299 541 300 545
rect 294 540 300 541
rect 478 545 484 546
rect 478 541 479 545
rect 483 541 484 545
rect 478 540 484 541
rect 662 545 668 546
rect 662 541 663 545
rect 667 541 668 545
rect 662 540 668 541
rect 838 545 844 546
rect 838 541 839 545
rect 843 541 844 545
rect 838 540 844 541
rect 1014 545 1020 546
rect 1014 541 1015 545
rect 1019 541 1020 545
rect 1014 540 1020 541
rect 1190 545 1196 546
rect 1190 541 1191 545
rect 1195 541 1196 545
rect 1190 540 1196 541
rect 1366 545 1372 546
rect 1366 541 1367 545
rect 1371 541 1372 545
rect 1366 540 1372 541
rect 1550 545 1556 546
rect 1550 541 1551 545
rect 1555 541 1556 545
rect 1550 540 1556 541
rect 1726 545 1732 546
rect 1726 541 1727 545
rect 1731 541 1732 545
rect 1726 540 1732 541
rect 2190 545 2196 546
rect 2190 541 2191 545
rect 2195 541 2196 545
rect 2190 540 2196 541
rect 2278 545 2284 546
rect 2278 541 2279 545
rect 2283 541 2284 545
rect 2278 540 2284 541
rect 2366 545 2372 546
rect 2366 541 2367 545
rect 2371 541 2372 545
rect 2366 540 2372 541
rect 2454 545 2460 546
rect 2454 541 2455 545
rect 2459 541 2460 545
rect 2454 540 2460 541
rect 2558 545 2564 546
rect 2558 541 2559 545
rect 2563 541 2564 545
rect 2558 540 2564 541
rect 2670 545 2676 546
rect 2670 541 2671 545
rect 2675 541 2676 545
rect 2670 540 2676 541
rect 2806 545 2812 546
rect 2806 541 2807 545
rect 2811 541 2812 545
rect 2806 540 2812 541
rect 2966 545 2972 546
rect 2966 541 2967 545
rect 2971 541 2972 545
rect 2966 540 2972 541
rect 3134 545 3140 546
rect 3134 541 3135 545
rect 3139 541 3140 545
rect 3134 540 3140 541
rect 3318 545 3324 546
rect 3318 541 3319 545
rect 3323 541 3324 545
rect 3318 540 3324 541
rect 3478 545 3484 546
rect 3478 541 3479 545
rect 3483 541 3484 545
rect 3478 540 3484 541
rect 527 539 536 540
rect 527 535 528 539
rect 535 535 536 539
rect 527 534 536 535
rect 1230 539 1236 540
rect 1230 535 1231 539
rect 1235 538 1236 539
rect 1239 539 1245 540
rect 1239 538 1240 539
rect 1235 536 1240 538
rect 1235 535 1236 536
rect 1230 534 1236 535
rect 1239 535 1240 536
rect 1244 535 1245 539
rect 1239 534 1245 535
rect 3518 539 3524 540
rect 3518 535 3519 539
rect 3523 538 3524 539
rect 3527 539 3533 540
rect 3527 538 3528 539
rect 3523 536 3528 538
rect 3523 535 3524 536
rect 3518 534 3524 535
rect 3527 535 3528 536
rect 3532 535 3533 539
rect 3527 534 3533 535
rect 134 519 140 520
rect 134 515 135 519
rect 139 515 140 519
rect 134 514 140 515
rect 302 519 308 520
rect 302 515 303 519
rect 307 515 308 519
rect 302 514 308 515
rect 494 519 500 520
rect 494 515 495 519
rect 499 515 500 519
rect 494 514 500 515
rect 678 519 684 520
rect 678 515 679 519
rect 683 515 684 519
rect 678 514 684 515
rect 862 519 868 520
rect 862 515 863 519
rect 867 515 868 519
rect 862 514 868 515
rect 1030 519 1036 520
rect 1030 515 1031 519
rect 1035 515 1036 519
rect 1030 514 1036 515
rect 1190 519 1196 520
rect 1190 515 1191 519
rect 1195 515 1196 519
rect 1190 514 1196 515
rect 1350 519 1356 520
rect 1350 515 1351 519
rect 1355 515 1356 519
rect 1350 514 1356 515
rect 1502 519 1508 520
rect 1502 515 1503 519
rect 1507 515 1508 519
rect 1502 514 1508 515
rect 1662 519 1668 520
rect 1662 515 1663 519
rect 1667 515 1668 519
rect 1662 514 1668 515
rect 2302 519 2308 520
rect 2302 515 2303 519
rect 2307 515 2308 519
rect 2302 514 2308 515
rect 2398 519 2404 520
rect 2398 515 2399 519
rect 2403 515 2404 519
rect 2398 514 2404 515
rect 2502 519 2508 520
rect 2502 515 2503 519
rect 2507 515 2508 519
rect 2502 514 2508 515
rect 2606 519 2612 520
rect 2606 515 2607 519
rect 2611 515 2612 519
rect 2606 514 2612 515
rect 2718 519 2724 520
rect 2718 515 2719 519
rect 2723 515 2724 519
rect 2718 514 2724 515
rect 2838 519 2844 520
rect 2838 515 2839 519
rect 2843 515 2844 519
rect 2838 514 2844 515
rect 2966 519 2972 520
rect 2966 515 2967 519
rect 2971 515 2972 519
rect 2966 514 2972 515
rect 3094 519 3100 520
rect 3094 515 3095 519
rect 3099 515 3100 519
rect 3094 514 3100 515
rect 3222 519 3228 520
rect 3222 515 3223 519
rect 3227 515 3228 519
rect 3222 514 3228 515
rect 3350 519 3356 520
rect 3350 515 3351 519
rect 3355 515 3356 519
rect 3350 514 3356 515
rect 3478 519 3484 520
rect 3478 515 3479 519
rect 3483 515 3484 519
rect 3478 514 3484 515
rect 790 511 796 512
rect 790 510 791 511
rect 110 509 116 510
rect 110 505 111 509
rect 115 505 116 509
rect 737 508 791 510
rect 790 507 791 508
rect 795 507 796 511
rect 2230 511 2236 512
rect 1040 508 1049 510
rect 1822 509 1828 510
rect 790 506 796 507
rect 1038 507 1044 508
rect 110 504 116 505
rect 1038 503 1039 507
rect 1043 503 1044 507
rect 1822 505 1823 509
rect 1827 505 1828 509
rect 1822 504 1828 505
rect 1862 509 1868 510
rect 1862 505 1863 509
rect 1867 505 1868 509
rect 2230 507 2231 511
rect 2235 510 2236 511
rect 3174 511 3180 512
rect 3174 510 3175 511
rect 2235 508 2321 510
rect 3153 508 3175 510
rect 2235 507 2236 508
rect 2230 506 2236 507
rect 3174 507 3175 508
rect 3179 507 3180 511
rect 3174 506 3180 507
rect 3290 511 3296 512
rect 3290 507 3291 511
rect 3295 510 3296 511
rect 3295 508 3369 510
rect 3574 509 3580 510
rect 3295 507 3296 508
rect 3290 506 3296 507
rect 1862 504 1868 505
rect 3574 505 3575 509
rect 3579 505 3580 509
rect 3574 504 3580 505
rect 1038 502 1044 503
rect 202 495 208 496
rect 110 492 116 493
rect 110 488 111 492
rect 115 488 116 492
rect 110 487 116 488
rect 197 488 199 494
rect 202 491 203 495
rect 207 494 208 495
rect 370 495 376 496
rect 207 492 329 494
rect 207 491 208 492
rect 202 490 208 491
rect 370 491 371 495
rect 375 494 376 495
rect 746 495 752 496
rect 375 492 521 494
rect 375 491 376 492
rect 370 490 376 491
rect 746 491 747 495
rect 751 494 752 495
rect 1343 495 1349 496
rect 1343 494 1344 495
rect 751 492 889 494
rect 1253 492 1344 494
rect 751 491 752 492
rect 746 490 752 491
rect 1343 491 1344 492
rect 1348 491 1349 495
rect 1418 495 1424 496
rect 1418 494 1419 495
rect 1413 492 1419 494
rect 1343 490 1349 491
rect 1418 491 1419 492
rect 1423 491 1424 495
rect 1570 495 1576 496
rect 1418 490 1424 491
rect 197 487 205 488
rect 197 484 200 487
rect 199 483 200 484
rect 204 483 205 487
rect 1564 486 1566 493
rect 1570 491 1571 495
rect 1575 494 1576 495
rect 2370 495 2376 496
rect 1575 492 1689 494
rect 1822 492 1828 493
rect 1575 491 1576 492
rect 1570 490 1576 491
rect 1822 488 1823 492
rect 1827 488 1828 492
rect 1586 487 1592 488
rect 1822 487 1828 488
rect 1862 492 1868 493
rect 1862 488 1863 492
rect 1867 488 1868 492
rect 2370 491 2371 495
rect 2375 494 2376 495
rect 2466 495 2472 496
rect 2375 492 2425 494
rect 2375 491 2376 492
rect 2370 490 2376 491
rect 2466 491 2467 495
rect 2471 494 2472 495
rect 2570 495 2576 496
rect 2471 492 2529 494
rect 2471 491 2472 492
rect 2466 490 2472 491
rect 2570 491 2571 495
rect 2575 494 2576 495
rect 2810 495 2816 496
rect 2810 494 2811 495
rect 2575 492 2633 494
rect 2781 492 2811 494
rect 2575 491 2576 492
rect 2570 490 2576 491
rect 2810 491 2811 492
rect 2815 491 2816 495
rect 2906 495 2912 496
rect 2906 494 2907 495
rect 2901 492 2907 494
rect 2810 490 2816 491
rect 2906 491 2907 492
rect 2911 491 2912 495
rect 3087 495 3093 496
rect 3087 494 3088 495
rect 3029 492 3088 494
rect 2906 490 2912 491
rect 3087 491 3088 492
rect 3092 491 3093 495
rect 3343 495 3349 496
rect 3343 494 3344 495
rect 3285 492 3344 494
rect 3087 490 3093 491
rect 3343 491 3344 492
rect 3348 491 3349 495
rect 3546 495 3552 496
rect 3546 494 3547 495
rect 3541 492 3547 494
rect 3343 490 3349 491
rect 3546 491 3547 492
rect 3551 491 3552 495
rect 3546 490 3552 491
rect 3574 492 3580 493
rect 1862 487 1868 488
rect 3574 488 3575 492
rect 3579 488 3580 492
rect 3574 487 3580 488
rect 1586 486 1587 487
rect 1564 484 1587 486
rect 199 482 205 483
rect 1586 483 1587 484
rect 1591 483 1592 487
rect 1586 482 1592 483
rect 142 479 148 480
rect 142 475 143 479
rect 147 475 148 479
rect 142 474 148 475
rect 310 479 316 480
rect 310 475 311 479
rect 315 475 316 479
rect 310 474 316 475
rect 502 479 508 480
rect 502 475 503 479
rect 507 475 508 479
rect 502 474 508 475
rect 686 479 692 480
rect 686 475 687 479
rect 691 475 692 479
rect 686 474 692 475
rect 870 479 876 480
rect 870 475 871 479
rect 875 475 876 479
rect 870 474 876 475
rect 1038 479 1044 480
rect 1038 475 1039 479
rect 1043 475 1044 479
rect 1038 474 1044 475
rect 1198 479 1204 480
rect 1198 475 1199 479
rect 1203 475 1204 479
rect 1198 474 1204 475
rect 1358 479 1364 480
rect 1358 475 1359 479
rect 1363 475 1364 479
rect 1358 474 1364 475
rect 1510 479 1516 480
rect 1510 475 1511 479
rect 1515 475 1516 479
rect 1510 474 1516 475
rect 1670 479 1676 480
rect 1670 475 1671 479
rect 1675 475 1676 479
rect 1670 474 1676 475
rect 2310 479 2316 480
rect 2310 475 2311 479
rect 2315 475 2316 479
rect 2310 474 2316 475
rect 2406 479 2412 480
rect 2406 475 2407 479
rect 2411 475 2412 479
rect 2406 474 2412 475
rect 2510 479 2516 480
rect 2510 475 2511 479
rect 2515 475 2516 479
rect 2510 474 2516 475
rect 2614 479 2620 480
rect 2614 475 2615 479
rect 2619 475 2620 479
rect 2614 474 2620 475
rect 2726 479 2732 480
rect 2726 475 2727 479
rect 2731 475 2732 479
rect 2726 474 2732 475
rect 2846 479 2852 480
rect 2846 475 2847 479
rect 2851 475 2852 479
rect 2846 474 2852 475
rect 2974 479 2980 480
rect 2974 475 2975 479
rect 2979 475 2980 479
rect 2974 474 2980 475
rect 3102 479 3108 480
rect 3102 475 3103 479
rect 3107 475 3108 479
rect 3102 474 3108 475
rect 3230 479 3236 480
rect 3230 475 3231 479
rect 3235 475 3236 479
rect 3230 474 3236 475
rect 3358 479 3364 480
rect 3358 475 3359 479
rect 3363 475 3364 479
rect 3358 474 3364 475
rect 3486 479 3492 480
rect 3486 475 3487 479
rect 3491 475 3492 479
rect 3486 474 3492 475
rect 171 467 177 468
rect 171 463 172 467
rect 176 466 177 467
rect 202 467 208 468
rect 202 466 203 467
rect 176 464 203 466
rect 176 463 177 464
rect 171 462 177 463
rect 202 463 203 464
rect 207 463 208 467
rect 202 462 208 463
rect 339 467 345 468
rect 339 463 340 467
rect 344 466 345 467
rect 370 467 376 468
rect 370 466 371 467
rect 344 464 371 466
rect 344 463 345 464
rect 339 462 345 463
rect 370 463 371 464
rect 375 463 376 467
rect 370 462 376 463
rect 530 467 537 468
rect 530 463 531 467
rect 536 463 537 467
rect 530 462 537 463
rect 715 467 721 468
rect 715 463 716 467
rect 720 466 721 467
rect 746 467 752 468
rect 746 466 747 467
rect 720 464 747 466
rect 720 463 721 464
rect 715 462 721 463
rect 746 463 747 464
rect 751 463 752 467
rect 746 462 752 463
rect 899 467 905 468
rect 899 463 900 467
rect 904 466 905 467
rect 938 467 944 468
rect 938 466 939 467
rect 904 464 939 466
rect 904 463 905 464
rect 899 462 905 463
rect 938 463 939 464
rect 943 463 944 467
rect 938 462 944 463
rect 1046 467 1052 468
rect 1046 463 1047 467
rect 1051 466 1052 467
rect 1067 467 1073 468
rect 1067 466 1068 467
rect 1051 464 1068 466
rect 1051 463 1052 464
rect 1046 462 1052 463
rect 1067 463 1068 464
rect 1072 463 1073 467
rect 1067 462 1073 463
rect 1227 467 1236 468
rect 1227 463 1228 467
rect 1235 463 1236 467
rect 1227 462 1236 463
rect 1343 467 1349 468
rect 1343 463 1344 467
rect 1348 466 1349 467
rect 1387 467 1393 468
rect 1387 466 1388 467
rect 1348 464 1388 466
rect 1348 463 1349 464
rect 1343 462 1349 463
rect 1387 463 1388 464
rect 1392 463 1393 467
rect 1387 462 1393 463
rect 1539 467 1545 468
rect 1539 463 1540 467
rect 1544 466 1545 467
rect 1570 467 1576 468
rect 1570 466 1571 467
rect 1544 464 1571 466
rect 1544 463 1545 464
rect 1539 462 1545 463
rect 1570 463 1571 464
rect 1575 463 1576 467
rect 1570 462 1576 463
rect 1699 467 1708 468
rect 1699 463 1700 467
rect 1707 463 1708 467
rect 1699 462 1708 463
rect 2339 467 2345 468
rect 2339 463 2340 467
rect 2344 466 2345 467
rect 2370 467 2376 468
rect 2370 466 2371 467
rect 2344 464 2371 466
rect 2344 463 2345 464
rect 2339 462 2345 463
rect 2370 463 2371 464
rect 2375 463 2376 467
rect 2370 462 2376 463
rect 2435 467 2441 468
rect 2435 463 2436 467
rect 2440 466 2441 467
rect 2466 467 2472 468
rect 2466 466 2467 467
rect 2440 464 2467 466
rect 2440 463 2441 464
rect 2435 462 2441 463
rect 2466 463 2467 464
rect 2471 463 2472 467
rect 2466 462 2472 463
rect 2539 467 2545 468
rect 2539 463 2540 467
rect 2544 466 2545 467
rect 2570 467 2576 468
rect 2570 466 2571 467
rect 2544 464 2571 466
rect 2544 463 2545 464
rect 2539 462 2545 463
rect 2570 463 2571 464
rect 2575 463 2576 467
rect 2570 462 2576 463
rect 2643 467 2652 468
rect 2643 463 2644 467
rect 2651 463 2652 467
rect 2643 462 2652 463
rect 2754 467 2761 468
rect 2754 463 2755 467
rect 2760 463 2761 467
rect 2754 462 2761 463
rect 2810 467 2816 468
rect 2810 463 2811 467
rect 2815 466 2816 467
rect 2875 467 2881 468
rect 2875 466 2876 467
rect 2815 464 2876 466
rect 2815 463 2816 464
rect 2810 462 2816 463
rect 2875 463 2876 464
rect 2880 463 2881 467
rect 2875 462 2881 463
rect 3003 467 3012 468
rect 3003 463 3004 467
rect 3011 463 3012 467
rect 3003 462 3012 463
rect 3087 467 3093 468
rect 3087 463 3088 467
rect 3092 466 3093 467
rect 3131 467 3137 468
rect 3131 466 3132 467
rect 3092 464 3132 466
rect 3092 463 3093 464
rect 3087 462 3093 463
rect 3131 463 3132 464
rect 3136 463 3137 467
rect 3131 462 3137 463
rect 3218 467 3224 468
rect 3218 463 3219 467
rect 3223 466 3224 467
rect 3259 467 3265 468
rect 3259 466 3260 467
rect 3223 464 3260 466
rect 3223 463 3224 464
rect 3218 462 3224 463
rect 3259 463 3260 464
rect 3264 463 3265 467
rect 3259 462 3265 463
rect 3343 467 3349 468
rect 3343 463 3344 467
rect 3348 466 3349 467
rect 3387 467 3393 468
rect 3387 466 3388 467
rect 3348 464 3388 466
rect 3348 463 3349 464
rect 3343 462 3349 463
rect 3387 463 3388 464
rect 3392 463 3393 467
rect 3387 462 3393 463
rect 3515 467 3524 468
rect 3515 463 3516 467
rect 3523 463 3524 467
rect 3515 462 3524 463
rect 2267 455 2276 456
rect 171 451 177 452
rect 171 447 172 451
rect 176 450 177 451
rect 199 451 205 452
rect 199 450 200 451
rect 176 448 200 450
rect 176 447 177 448
rect 171 446 177 447
rect 199 447 200 448
rect 204 447 205 451
rect 199 446 205 447
rect 207 451 213 452
rect 207 447 208 451
rect 212 450 213 451
rect 331 451 337 452
rect 331 450 332 451
rect 212 448 332 450
rect 212 447 213 448
rect 207 446 213 447
rect 331 447 332 448
rect 336 447 337 451
rect 331 446 337 447
rect 375 451 381 452
rect 375 447 376 451
rect 380 450 381 451
rect 523 451 529 452
rect 523 450 524 451
rect 380 448 524 450
rect 380 447 381 448
rect 375 446 381 447
rect 523 447 524 448
rect 528 447 529 451
rect 523 446 529 447
rect 663 451 669 452
rect 663 447 664 451
rect 668 450 669 451
rect 715 451 721 452
rect 715 450 716 451
rect 668 448 716 450
rect 668 447 669 448
rect 663 446 669 447
rect 715 447 716 448
rect 720 447 721 451
rect 715 446 721 447
rect 759 451 765 452
rect 759 447 760 451
rect 764 450 765 451
rect 907 451 913 452
rect 907 450 908 451
rect 764 448 908 450
rect 764 447 765 448
rect 759 446 765 447
rect 907 447 908 448
rect 912 447 913 451
rect 907 446 913 447
rect 1083 451 1089 452
rect 1083 447 1084 451
rect 1088 450 1089 451
rect 1094 451 1100 452
rect 1094 450 1095 451
rect 1088 448 1095 450
rect 1088 447 1089 448
rect 1083 446 1089 447
rect 1094 447 1095 448
rect 1099 447 1100 451
rect 1094 446 1100 447
rect 1251 451 1257 452
rect 1251 447 1252 451
rect 1256 450 1257 451
rect 1290 451 1296 452
rect 1290 450 1291 451
rect 1256 448 1291 450
rect 1256 447 1257 448
rect 1251 446 1257 447
rect 1290 447 1291 448
rect 1295 447 1296 451
rect 1290 446 1296 447
rect 1418 451 1425 452
rect 1418 447 1419 451
rect 1424 447 1425 451
rect 1418 446 1425 447
rect 1586 451 1593 452
rect 1586 447 1587 451
rect 1592 447 1593 451
rect 1586 446 1593 447
rect 1663 451 1669 452
rect 1663 447 1664 451
rect 1668 450 1669 451
rect 1755 451 1761 452
rect 1755 450 1756 451
rect 1668 448 1756 450
rect 1668 447 1669 448
rect 1663 446 1669 447
rect 1755 447 1756 448
rect 1760 447 1761 451
rect 2267 451 2268 455
rect 2275 451 2276 455
rect 2267 450 2276 451
rect 2303 455 2309 456
rect 2303 451 2304 455
rect 2308 454 2309 455
rect 2355 455 2361 456
rect 2355 454 2356 455
rect 2308 452 2356 454
rect 2308 451 2309 452
rect 2303 450 2309 451
rect 2355 451 2356 452
rect 2360 451 2361 455
rect 2355 450 2361 451
rect 2399 455 2405 456
rect 2399 451 2400 455
rect 2404 454 2405 455
rect 2459 455 2465 456
rect 2459 454 2460 455
rect 2404 452 2460 454
rect 2404 451 2405 452
rect 2399 450 2405 451
rect 2459 451 2460 452
rect 2464 451 2465 455
rect 2459 450 2465 451
rect 2511 455 2517 456
rect 2511 451 2512 455
rect 2516 454 2517 455
rect 2587 455 2593 456
rect 2587 454 2588 455
rect 2516 452 2588 454
rect 2516 451 2517 452
rect 2511 450 2517 451
rect 2587 451 2588 452
rect 2592 451 2593 455
rect 2587 450 2593 451
rect 2631 455 2637 456
rect 2631 451 2632 455
rect 2636 454 2637 455
rect 2723 455 2729 456
rect 2723 454 2724 455
rect 2636 452 2724 454
rect 2636 451 2637 452
rect 2631 450 2637 451
rect 2723 451 2724 452
rect 2728 451 2729 455
rect 2723 450 2729 451
rect 2875 455 2881 456
rect 2875 451 2876 455
rect 2880 454 2881 455
rect 2906 455 2912 456
rect 2906 454 2907 455
rect 2880 452 2907 454
rect 2880 451 2881 452
rect 2875 450 2881 451
rect 2906 451 2907 452
rect 2911 451 2912 455
rect 2906 450 2912 451
rect 2943 455 2949 456
rect 2943 451 2944 455
rect 2948 454 2949 455
rect 3027 455 3033 456
rect 3027 454 3028 455
rect 2948 452 3028 454
rect 2948 451 2949 452
rect 2943 450 2949 451
rect 3027 451 3028 452
rect 3032 451 3033 455
rect 3027 450 3033 451
rect 3187 455 3193 456
rect 3187 451 3188 455
rect 3192 454 3193 455
rect 3262 455 3268 456
rect 3262 454 3263 455
rect 3192 452 3263 454
rect 3192 451 3193 452
rect 3187 450 3193 451
rect 3262 451 3263 452
rect 3267 451 3268 455
rect 3262 450 3268 451
rect 3355 455 3361 456
rect 3355 451 3356 455
rect 3360 454 3361 455
rect 3407 455 3413 456
rect 3407 454 3408 455
rect 3360 452 3408 454
rect 3360 451 3361 452
rect 3355 450 3361 451
rect 3407 451 3408 452
rect 3412 451 3413 455
rect 3407 450 3413 451
rect 3515 455 3521 456
rect 3515 451 3516 455
rect 3520 454 3521 455
rect 3546 455 3552 456
rect 3546 454 3547 455
rect 3520 452 3547 454
rect 3520 451 3521 452
rect 3515 450 3521 451
rect 3546 451 3547 452
rect 3551 451 3552 455
rect 3546 450 3552 451
rect 1755 446 1761 447
rect 2238 445 2244 446
rect 142 441 148 442
rect 142 437 143 441
rect 147 437 148 441
rect 142 436 148 437
rect 302 441 308 442
rect 302 437 303 441
rect 307 437 308 441
rect 302 436 308 437
rect 494 441 500 442
rect 494 437 495 441
rect 499 437 500 441
rect 494 436 500 437
rect 686 441 692 442
rect 686 437 687 441
rect 691 437 692 441
rect 686 436 692 437
rect 878 441 884 442
rect 878 437 879 441
rect 883 437 884 441
rect 878 436 884 437
rect 1054 441 1060 442
rect 1054 437 1055 441
rect 1059 437 1060 441
rect 1054 436 1060 437
rect 1222 441 1228 442
rect 1222 437 1223 441
rect 1227 437 1228 441
rect 1222 436 1228 437
rect 1390 441 1396 442
rect 1390 437 1391 441
rect 1395 437 1396 441
rect 1390 436 1396 437
rect 1558 441 1564 442
rect 1558 437 1559 441
rect 1563 437 1564 441
rect 1558 436 1564 437
rect 1726 441 1732 442
rect 1726 437 1727 441
rect 1731 437 1732 441
rect 2238 441 2239 445
rect 2243 441 2244 445
rect 2238 440 2244 441
rect 2326 445 2332 446
rect 2326 441 2327 445
rect 2331 441 2332 445
rect 2326 440 2332 441
rect 2430 445 2436 446
rect 2430 441 2431 445
rect 2435 441 2436 445
rect 2430 440 2436 441
rect 2558 445 2564 446
rect 2558 441 2559 445
rect 2563 441 2564 445
rect 2558 440 2564 441
rect 2694 445 2700 446
rect 2694 441 2695 445
rect 2699 441 2700 445
rect 2694 440 2700 441
rect 2846 445 2852 446
rect 2846 441 2847 445
rect 2851 441 2852 445
rect 2846 440 2852 441
rect 2998 445 3004 446
rect 2998 441 2999 445
rect 3003 441 3004 445
rect 2998 440 3004 441
rect 3158 445 3164 446
rect 3158 441 3159 445
rect 3163 441 3164 445
rect 3158 440 3164 441
rect 3326 445 3332 446
rect 3326 441 3327 445
rect 3331 441 3332 445
rect 3326 440 3332 441
rect 3486 445 3492 446
rect 3486 441 3487 445
rect 3491 441 3492 445
rect 3486 440 3492 441
rect 1726 436 1732 437
rect 1862 432 1868 433
rect 3574 432 3580 433
rect 110 428 116 429
rect 1822 428 1828 429
rect 110 424 111 428
rect 115 424 116 428
rect 207 427 213 428
rect 207 426 208 427
rect 197 424 208 426
rect 110 423 116 424
rect 207 423 208 424
rect 212 423 213 427
rect 375 427 381 428
rect 375 426 376 427
rect 357 424 376 426
rect 207 422 213 423
rect 375 423 376 424
rect 380 423 381 427
rect 759 427 765 428
rect 759 426 760 427
rect 741 424 760 426
rect 375 422 381 423
rect 759 423 760 424
rect 764 423 765 427
rect 938 427 944 428
rect 938 426 939 427
rect 933 424 939 426
rect 759 422 765 423
rect 938 423 939 424
rect 943 423 944 427
rect 1663 427 1669 428
rect 1663 426 1664 427
rect 1613 424 1664 426
rect 938 422 944 423
rect 1046 423 1052 424
rect 1046 419 1047 423
rect 1051 422 1052 423
rect 1290 423 1296 424
rect 1051 420 1073 422
rect 1051 419 1052 420
rect 1046 418 1052 419
rect 1290 419 1291 423
rect 1295 422 1296 423
rect 1663 423 1664 424
rect 1668 423 1669 427
rect 1822 424 1823 428
rect 1827 424 1828 428
rect 1862 428 1863 432
rect 1867 428 1868 432
rect 2303 431 2309 432
rect 2303 430 2304 431
rect 2293 428 2304 430
rect 1862 427 1868 428
rect 2303 427 2304 428
rect 2308 427 2309 431
rect 2399 431 2405 432
rect 2399 430 2400 431
rect 2381 428 2400 430
rect 2303 426 2309 427
rect 2399 427 2400 428
rect 2404 427 2405 431
rect 2511 431 2517 432
rect 2511 430 2512 431
rect 2485 428 2512 430
rect 2399 426 2405 427
rect 2511 427 2512 428
rect 2516 427 2517 431
rect 2631 431 2637 432
rect 2631 430 2632 431
rect 2613 428 2632 430
rect 2511 426 2517 427
rect 2631 427 2632 428
rect 2636 427 2637 431
rect 2943 431 2949 432
rect 2943 430 2944 431
rect 2901 428 2944 430
rect 2631 426 2637 427
rect 2646 427 2652 428
rect 1822 423 1828 424
rect 2646 423 2647 427
rect 2651 426 2652 427
rect 2943 427 2944 428
rect 2948 427 2949 431
rect 3218 431 3224 432
rect 3218 430 3219 431
rect 3213 428 3219 430
rect 2943 426 2949 427
rect 3218 427 3219 428
rect 3223 427 3224 431
rect 3574 428 3575 432
rect 3579 428 3580 432
rect 3218 426 3224 427
rect 3262 427 3268 428
rect 3574 427 3580 428
rect 2651 424 2713 426
rect 2651 423 2652 424
rect 1663 422 1669 423
rect 2646 422 2652 423
rect 3262 423 3263 427
rect 3267 426 3268 427
rect 3267 424 3345 426
rect 3267 423 3268 424
rect 3262 422 3268 423
rect 1295 420 1409 422
rect 1295 419 1296 420
rect 1290 418 1296 419
rect 1862 415 1868 416
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 110 406 116 407
rect 462 411 468 412
rect 462 407 463 411
rect 467 410 468 411
rect 1298 411 1304 412
rect 1298 410 1299 411
rect 467 408 505 410
rect 1273 408 1299 410
rect 467 407 468 408
rect 462 406 468 407
rect 1298 407 1299 408
rect 1303 407 1304 411
rect 1298 406 1304 407
rect 1822 411 1828 412
rect 1822 407 1823 411
rect 1827 407 1828 411
rect 1862 411 1863 415
rect 1867 411 1868 415
rect 1862 410 1868 411
rect 2998 415 3004 416
rect 2998 411 2999 415
rect 3003 414 3004 415
rect 3574 415 3580 416
rect 3003 412 3009 414
rect 3003 411 3004 412
rect 2998 410 3004 411
rect 3574 411 3575 415
rect 3579 411 3580 415
rect 3574 410 3580 411
rect 1822 406 1828 407
rect 2230 405 2236 406
rect 134 401 140 402
rect 134 397 135 401
rect 139 397 140 401
rect 134 396 140 397
rect 294 401 300 402
rect 294 397 295 401
rect 299 397 300 401
rect 294 396 300 397
rect 486 401 492 402
rect 486 397 487 401
rect 491 397 492 401
rect 486 396 492 397
rect 678 401 684 402
rect 678 397 679 401
rect 683 397 684 401
rect 678 396 684 397
rect 870 401 876 402
rect 870 397 871 401
rect 875 397 876 401
rect 870 396 876 397
rect 1046 401 1052 402
rect 1046 397 1047 401
rect 1051 397 1052 401
rect 1046 396 1052 397
rect 1214 401 1220 402
rect 1214 397 1215 401
rect 1219 397 1220 401
rect 1214 396 1220 397
rect 1382 401 1388 402
rect 1382 397 1383 401
rect 1387 397 1388 401
rect 1382 396 1388 397
rect 1550 401 1556 402
rect 1550 397 1551 401
rect 1555 397 1556 401
rect 1550 396 1556 397
rect 1718 401 1724 402
rect 1718 397 1719 401
rect 1723 397 1724 401
rect 2230 401 2231 405
rect 2235 401 2236 405
rect 2230 400 2236 401
rect 2318 405 2324 406
rect 2318 401 2319 405
rect 2323 401 2324 405
rect 2318 400 2324 401
rect 2422 405 2428 406
rect 2422 401 2423 405
rect 2427 401 2428 405
rect 2422 400 2428 401
rect 2550 405 2556 406
rect 2550 401 2551 405
rect 2555 401 2556 405
rect 2550 400 2556 401
rect 2686 405 2692 406
rect 2686 401 2687 405
rect 2691 401 2692 405
rect 2686 400 2692 401
rect 2838 405 2844 406
rect 2838 401 2839 405
rect 2843 401 2844 405
rect 2838 400 2844 401
rect 2990 405 2996 406
rect 2990 401 2991 405
rect 2995 401 2996 405
rect 2990 400 2996 401
rect 3150 405 3156 406
rect 3150 401 3151 405
rect 3155 401 3156 405
rect 3150 400 3156 401
rect 3318 405 3324 406
rect 3318 401 3319 405
rect 3323 401 3324 405
rect 3318 400 3324 401
rect 3478 405 3484 406
rect 3478 401 3479 405
rect 3483 401 3484 405
rect 3478 400 3484 401
rect 1718 396 1724 397
rect 3518 399 3524 400
rect 1766 395 1773 396
rect 1766 391 1767 395
rect 1772 391 1773 395
rect 3518 395 3519 399
rect 3523 398 3524 399
rect 3527 399 3533 400
rect 3527 398 3528 399
rect 3523 396 3528 398
rect 3523 395 3524 396
rect 3518 394 3524 395
rect 3527 395 3528 396
rect 3532 395 3533 399
rect 3527 394 3533 395
rect 1766 390 1773 391
rect 2270 391 2276 392
rect 2270 387 2271 391
rect 2275 390 2276 391
rect 2275 388 2470 390
rect 2275 387 2276 388
rect 2270 386 2276 387
rect 2182 383 2188 384
rect 134 379 140 380
rect 134 375 135 379
rect 139 375 140 379
rect 134 374 140 375
rect 262 379 268 380
rect 262 375 263 379
rect 267 375 268 379
rect 262 374 268 375
rect 422 379 428 380
rect 422 375 423 379
rect 427 375 428 379
rect 422 374 428 375
rect 590 379 596 380
rect 590 375 591 379
rect 595 375 596 379
rect 590 374 596 375
rect 766 379 772 380
rect 766 375 767 379
rect 771 375 772 379
rect 766 374 772 375
rect 934 379 940 380
rect 934 375 935 379
rect 939 375 940 379
rect 934 374 940 375
rect 1102 379 1108 380
rect 1102 375 1103 379
rect 1107 375 1108 379
rect 1102 374 1108 375
rect 1262 379 1268 380
rect 1262 375 1263 379
rect 1267 375 1268 379
rect 1262 374 1268 375
rect 1422 379 1428 380
rect 1422 375 1423 379
rect 1427 375 1428 379
rect 1422 374 1428 375
rect 1582 379 1588 380
rect 1582 375 1583 379
rect 1587 375 1588 379
rect 1582 374 1588 375
rect 1726 379 1732 380
rect 1726 375 1727 379
rect 1731 375 1732 379
rect 2182 379 2183 383
rect 2187 379 2188 383
rect 2182 378 2188 379
rect 2286 383 2292 384
rect 2286 379 2287 383
rect 2291 379 2292 383
rect 2286 378 2292 379
rect 2398 383 2404 384
rect 2398 379 2399 383
rect 2403 379 2404 383
rect 2398 378 2404 379
rect 1726 374 1732 375
rect 2468 374 2470 388
rect 2526 383 2532 384
rect 2526 379 2527 383
rect 2531 379 2532 383
rect 2526 378 2532 379
rect 2670 383 2676 384
rect 2670 379 2671 383
rect 2675 379 2676 383
rect 2670 378 2676 379
rect 2814 383 2820 384
rect 2814 379 2815 383
rect 2819 379 2820 383
rect 2814 378 2820 379
rect 2966 383 2972 384
rect 2966 379 2967 383
rect 2971 379 2972 383
rect 2966 378 2972 379
rect 3126 383 3132 384
rect 3126 379 3127 383
rect 3131 379 3132 383
rect 3126 378 3132 379
rect 3294 383 3300 384
rect 3294 379 3295 383
rect 3299 379 3300 383
rect 3294 378 3300 379
rect 3462 383 3468 384
rect 3462 379 3463 383
rect 3467 379 3468 383
rect 3462 378 3468 379
rect 3407 375 3413 376
rect 1862 373 1868 374
rect 663 371 669 372
rect 663 370 664 371
rect 110 369 116 370
rect 110 365 111 369
rect 115 365 116 369
rect 649 368 664 370
rect 663 367 664 368
rect 668 367 669 371
rect 663 366 669 367
rect 1094 371 1100 372
rect 1094 367 1095 371
rect 1099 370 1100 371
rect 1099 368 1121 370
rect 1822 369 1828 370
rect 1099 367 1100 368
rect 1094 366 1100 367
rect 110 364 116 365
rect 1822 365 1823 369
rect 1827 365 1828 369
rect 1862 369 1863 373
rect 1867 369 1868 373
rect 2468 372 2545 374
rect 3407 371 3408 375
rect 3412 374 3413 375
rect 3412 372 3481 374
rect 3574 373 3580 374
rect 3412 371 3413 372
rect 3407 370 3413 371
rect 1862 368 1868 369
rect 3574 369 3575 373
rect 3579 369 3580 373
rect 3574 368 3580 369
rect 1822 364 1828 365
rect 2279 359 2285 360
rect 2279 358 2280 359
rect 1862 356 1868 357
rect 2245 356 2280 358
rect 207 355 213 356
rect 110 352 116 353
rect 110 348 111 352
rect 115 348 116 352
rect 110 347 116 348
rect 196 346 198 353
rect 207 351 208 355
rect 212 354 213 355
rect 330 355 336 356
rect 212 352 289 354
rect 212 351 213 352
rect 207 350 213 351
rect 330 351 331 355
rect 335 354 336 355
rect 658 355 664 356
rect 335 352 449 354
rect 335 351 336 352
rect 330 350 336 351
rect 658 351 659 355
rect 663 354 664 355
rect 1034 355 1040 356
rect 1034 354 1035 355
rect 663 352 793 354
rect 997 352 1035 354
rect 663 351 664 352
rect 658 350 664 351
rect 1034 351 1035 352
rect 1039 351 1040 355
rect 1034 350 1040 351
rect 1254 355 1260 356
rect 1254 351 1255 355
rect 1259 354 1260 355
rect 1575 355 1581 356
rect 1575 354 1576 355
rect 1259 352 1289 354
rect 1485 352 1576 354
rect 1259 351 1260 352
rect 1254 350 1260 351
rect 1575 351 1576 352
rect 1580 351 1581 355
rect 1650 355 1656 356
rect 1650 354 1651 355
rect 1645 352 1651 354
rect 1575 350 1581 351
rect 1650 351 1651 352
rect 1655 351 1656 355
rect 1650 350 1656 351
rect 1658 355 1664 356
rect 1658 351 1659 355
rect 1663 354 1664 355
rect 1663 352 1753 354
rect 1822 352 1828 353
rect 1663 351 1664 352
rect 1658 350 1664 351
rect 1822 348 1823 352
rect 1827 348 1828 352
rect 1862 352 1863 356
rect 1867 352 1868 356
rect 2279 355 2280 356
rect 2284 355 2285 359
rect 2391 359 2397 360
rect 2391 358 2392 359
rect 2349 356 2392 358
rect 2279 354 2285 355
rect 2391 355 2392 356
rect 2396 355 2397 359
rect 2519 359 2525 360
rect 2519 358 2520 359
rect 2461 356 2520 358
rect 2391 354 2397 355
rect 2519 355 2520 356
rect 2524 355 2525 359
rect 2519 354 2525 355
rect 2594 359 2600 360
rect 2594 355 2595 359
rect 2599 358 2600 359
rect 2743 359 2749 360
rect 2599 356 2697 358
rect 2599 355 2600 356
rect 2594 354 2600 355
rect 2743 355 2744 359
rect 2748 358 2749 359
rect 2882 359 2888 360
rect 2748 356 2841 358
rect 2748 355 2749 356
rect 2743 354 2749 355
rect 2882 355 2883 359
rect 2887 358 2888 359
rect 3287 359 3293 360
rect 3287 358 3288 359
rect 2887 356 2993 358
rect 3189 356 3288 358
rect 2887 355 2888 356
rect 2882 354 2888 355
rect 3287 355 3288 356
rect 3292 355 3293 359
rect 3455 359 3461 360
rect 3455 358 3456 359
rect 3357 356 3456 358
rect 3287 354 3293 355
rect 3455 355 3456 356
rect 3460 355 3461 359
rect 3455 354 3461 355
rect 3574 356 3580 357
rect 1862 351 1868 352
rect 3574 352 3575 356
rect 3579 352 3580 356
rect 3574 351 3580 352
rect 242 347 248 348
rect 1822 347 1828 348
rect 242 346 243 347
rect 196 344 243 346
rect 242 343 243 344
rect 247 343 248 347
rect 242 342 248 343
rect 2190 343 2196 344
rect 142 339 148 340
rect 142 335 143 339
rect 147 335 148 339
rect 142 334 148 335
rect 270 339 276 340
rect 270 335 271 339
rect 275 335 276 339
rect 270 334 276 335
rect 430 339 436 340
rect 430 335 431 339
rect 435 335 436 339
rect 430 334 436 335
rect 598 339 604 340
rect 598 335 599 339
rect 603 335 604 339
rect 598 334 604 335
rect 774 339 780 340
rect 774 335 775 339
rect 779 335 780 339
rect 774 334 780 335
rect 942 339 948 340
rect 942 335 943 339
rect 947 335 948 339
rect 942 334 948 335
rect 1110 339 1116 340
rect 1110 335 1111 339
rect 1115 335 1116 339
rect 1110 334 1116 335
rect 1270 339 1276 340
rect 1270 335 1271 339
rect 1275 335 1276 339
rect 1270 334 1276 335
rect 1430 339 1436 340
rect 1430 335 1431 339
rect 1435 335 1436 339
rect 1430 334 1436 335
rect 1590 339 1596 340
rect 1590 335 1591 339
rect 1595 335 1596 339
rect 1734 339 1740 340
rect 1590 334 1596 335
rect 1658 335 1664 336
rect 1658 334 1659 335
rect 1460 332 1586 334
rect 1460 330 1462 332
rect 1584 330 1586 332
rect 1600 332 1659 334
rect 1600 330 1602 332
rect 1658 331 1659 332
rect 1663 331 1664 335
rect 1734 335 1735 339
rect 1739 335 1740 339
rect 2190 339 2191 343
rect 2195 339 2196 343
rect 2190 338 2196 339
rect 2294 343 2300 344
rect 2294 339 2295 343
rect 2299 339 2300 343
rect 2294 338 2300 339
rect 2406 343 2412 344
rect 2406 339 2407 343
rect 2411 339 2412 343
rect 2406 338 2412 339
rect 2534 343 2540 344
rect 2534 339 2535 343
rect 2539 339 2540 343
rect 2534 338 2540 339
rect 2678 343 2684 344
rect 2678 339 2679 343
rect 2683 339 2684 343
rect 2678 338 2684 339
rect 2822 343 2828 344
rect 2822 339 2823 343
rect 2827 339 2828 343
rect 2822 338 2828 339
rect 2974 343 2980 344
rect 2974 339 2975 343
rect 2979 339 2980 343
rect 2974 338 2980 339
rect 3134 343 3140 344
rect 3134 339 3135 343
rect 3139 339 3140 343
rect 3134 338 3140 339
rect 3302 343 3308 344
rect 3302 339 3303 343
rect 3307 339 3308 343
rect 3302 338 3308 339
rect 3470 343 3476 344
rect 3470 339 3471 343
rect 3475 339 3476 343
rect 3470 338 3476 339
rect 1734 334 1740 335
rect 1658 330 1664 331
rect 2159 331 2165 332
rect 1459 329 1465 330
rect 171 327 177 328
rect 171 323 172 327
rect 176 326 177 327
rect 207 327 213 328
rect 207 326 208 327
rect 176 324 208 326
rect 176 323 177 324
rect 171 322 177 323
rect 207 323 208 324
rect 212 323 213 327
rect 207 322 213 323
rect 299 327 305 328
rect 299 323 300 327
rect 304 326 305 327
rect 330 327 336 328
rect 330 326 331 327
rect 304 324 331 326
rect 304 323 305 324
rect 299 322 305 323
rect 330 323 331 324
rect 335 323 336 327
rect 330 322 336 323
rect 459 327 468 328
rect 459 323 460 327
rect 467 323 468 327
rect 459 322 468 323
rect 627 327 633 328
rect 627 323 628 327
rect 632 326 633 327
rect 658 327 664 328
rect 658 326 659 327
rect 632 324 659 326
rect 632 323 633 324
rect 627 322 633 323
rect 658 323 659 324
rect 663 323 664 327
rect 658 322 664 323
rect 782 327 788 328
rect 782 323 783 327
rect 787 326 788 327
rect 803 327 809 328
rect 803 326 804 327
rect 787 324 804 326
rect 787 323 788 324
rect 782 322 788 323
rect 803 323 804 324
rect 808 323 809 327
rect 803 322 809 323
rect 971 327 977 328
rect 971 323 972 327
rect 976 326 977 327
rect 994 327 1000 328
rect 994 326 995 327
rect 976 324 995 326
rect 976 323 977 324
rect 971 322 977 323
rect 994 323 995 324
rect 999 323 1000 327
rect 994 322 1000 323
rect 1034 327 1040 328
rect 1034 323 1035 327
rect 1039 326 1040 327
rect 1139 327 1145 328
rect 1139 326 1140 327
rect 1039 324 1140 326
rect 1039 323 1040 324
rect 1034 322 1040 323
rect 1139 323 1140 324
rect 1144 323 1145 327
rect 1139 322 1145 323
rect 1298 327 1305 328
rect 1298 323 1299 327
rect 1304 323 1305 327
rect 1459 325 1460 329
rect 1464 325 1465 329
rect 1584 328 1602 330
rect 1459 324 1465 325
rect 1575 327 1581 328
rect 1298 322 1305 323
rect 1575 323 1576 327
rect 1580 326 1581 327
rect 1619 327 1625 328
rect 1619 326 1620 327
rect 1580 324 1620 326
rect 1580 323 1581 324
rect 1575 322 1581 323
rect 1619 323 1620 324
rect 1624 323 1625 327
rect 1619 322 1625 323
rect 1763 327 1772 328
rect 1763 323 1764 327
rect 1771 323 1772 327
rect 2159 327 2160 331
rect 2164 330 2165 331
rect 2219 331 2225 332
rect 2219 330 2220 331
rect 2164 328 2220 330
rect 2164 327 2165 328
rect 2159 326 2165 327
rect 2219 327 2220 328
rect 2224 327 2225 331
rect 2219 326 2225 327
rect 2279 331 2285 332
rect 2279 327 2280 331
rect 2284 330 2285 331
rect 2323 331 2329 332
rect 2323 330 2324 331
rect 2284 328 2324 330
rect 2284 327 2285 328
rect 2279 326 2285 327
rect 2323 327 2324 328
rect 2328 327 2329 331
rect 2323 326 2329 327
rect 2391 331 2397 332
rect 2391 327 2392 331
rect 2396 330 2397 331
rect 2435 331 2441 332
rect 2435 330 2436 331
rect 2396 328 2436 330
rect 2396 327 2397 328
rect 2391 326 2397 327
rect 2435 327 2436 328
rect 2440 327 2441 331
rect 2435 326 2441 327
rect 2519 331 2525 332
rect 2519 327 2520 331
rect 2524 330 2525 331
rect 2563 331 2569 332
rect 2563 330 2564 331
rect 2524 328 2564 330
rect 2524 327 2525 328
rect 2519 326 2525 327
rect 2563 327 2564 328
rect 2568 327 2569 331
rect 2563 326 2569 327
rect 2707 331 2713 332
rect 2707 327 2708 331
rect 2712 330 2713 331
rect 2743 331 2749 332
rect 2743 330 2744 331
rect 2712 328 2744 330
rect 2712 327 2713 328
rect 2707 326 2713 327
rect 2743 327 2744 328
rect 2748 327 2749 331
rect 2743 326 2749 327
rect 2851 331 2857 332
rect 2851 327 2852 331
rect 2856 330 2857 331
rect 2882 331 2888 332
rect 2882 330 2883 331
rect 2856 328 2883 330
rect 2856 327 2857 328
rect 2851 326 2857 327
rect 2882 327 2883 328
rect 2887 327 2888 331
rect 2882 326 2888 327
rect 2998 331 3009 332
rect 2998 327 2999 331
rect 3003 327 3004 331
rect 3008 327 3009 331
rect 2998 326 3009 327
rect 3154 331 3160 332
rect 3154 327 3155 331
rect 3159 330 3160 331
rect 3163 331 3169 332
rect 3163 330 3164 331
rect 3159 328 3164 330
rect 3159 327 3160 328
rect 3154 326 3160 327
rect 3163 327 3164 328
rect 3168 327 3169 331
rect 3163 326 3169 327
rect 3287 331 3293 332
rect 3287 327 3288 331
rect 3292 330 3293 331
rect 3331 331 3337 332
rect 3331 330 3332 331
rect 3292 328 3332 330
rect 3292 327 3293 328
rect 3287 326 3293 327
rect 3331 327 3332 328
rect 3336 327 3337 331
rect 3331 326 3337 327
rect 3455 331 3461 332
rect 3455 327 3456 331
rect 3460 330 3461 331
rect 3499 331 3505 332
rect 3499 330 3500 331
rect 3460 328 3500 330
rect 3460 327 3461 328
rect 3455 326 3461 327
rect 3499 327 3500 328
rect 3504 327 3505 331
rect 3499 326 3505 327
rect 1763 322 1772 323
rect 242 315 249 316
rect 242 311 243 315
rect 248 311 249 315
rect 242 310 249 311
rect 303 315 309 316
rect 303 311 304 315
rect 308 314 309 315
rect 379 315 385 316
rect 379 314 380 315
rect 308 312 380 314
rect 308 311 309 312
rect 303 310 309 311
rect 379 311 380 312
rect 384 311 385 315
rect 379 310 385 311
rect 523 315 529 316
rect 523 311 524 315
rect 528 314 529 315
rect 554 315 560 316
rect 554 314 555 315
rect 528 312 555 314
rect 528 311 529 312
rect 523 310 529 311
rect 554 311 555 312
rect 559 311 560 315
rect 554 310 560 311
rect 567 315 573 316
rect 567 311 568 315
rect 572 314 573 315
rect 667 315 673 316
rect 667 314 668 315
rect 572 312 668 314
rect 572 311 573 312
rect 567 310 573 311
rect 667 311 668 312
rect 672 311 673 315
rect 667 310 673 311
rect 735 315 741 316
rect 735 311 736 315
rect 740 314 741 315
rect 819 315 825 316
rect 819 314 820 315
rect 740 312 820 314
rect 740 311 741 312
rect 735 310 741 311
rect 819 311 820 312
rect 824 311 825 315
rect 819 310 825 311
rect 963 315 969 316
rect 963 311 964 315
rect 968 314 969 315
rect 1023 315 1029 316
rect 1023 314 1024 315
rect 968 312 1024 314
rect 968 311 969 312
rect 963 310 969 311
rect 1023 311 1024 312
rect 1028 311 1029 315
rect 1023 310 1029 311
rect 1098 315 1104 316
rect 1098 311 1099 315
rect 1103 314 1104 315
rect 1107 315 1113 316
rect 1107 314 1108 315
rect 1103 312 1108 314
rect 1103 311 1104 312
rect 1098 310 1104 311
rect 1107 311 1108 312
rect 1112 311 1113 315
rect 1107 310 1113 311
rect 1251 315 1260 316
rect 1251 311 1252 315
rect 1259 311 1260 315
rect 1251 310 1260 311
rect 1311 315 1317 316
rect 1311 311 1312 315
rect 1316 314 1317 315
rect 1387 315 1393 316
rect 1387 314 1388 315
rect 1316 312 1388 314
rect 1316 311 1317 312
rect 1311 310 1317 311
rect 1387 311 1388 312
rect 1392 311 1393 315
rect 1387 310 1393 311
rect 1423 315 1429 316
rect 1423 311 1424 315
rect 1428 314 1429 315
rect 1515 315 1521 316
rect 1515 314 1516 315
rect 1428 312 1516 314
rect 1428 311 1429 312
rect 1423 310 1429 311
rect 1515 311 1516 312
rect 1520 311 1521 315
rect 1515 310 1521 311
rect 1650 315 1657 316
rect 1650 311 1651 315
rect 1656 311 1657 315
rect 1650 310 1657 311
rect 1695 315 1701 316
rect 1695 311 1696 315
rect 1700 314 1701 315
rect 1763 315 1769 316
rect 1763 314 1764 315
rect 1700 312 1764 314
rect 1700 311 1701 312
rect 1695 310 1701 311
rect 1763 311 1764 312
rect 1768 311 1769 315
rect 1763 310 1769 311
rect 1807 311 1813 312
rect 1807 307 1808 311
rect 1812 310 1813 311
rect 1923 311 1929 312
rect 1923 310 1924 311
rect 1812 308 1924 310
rect 1812 307 1813 308
rect 1807 306 1813 307
rect 1923 307 1924 308
rect 1928 307 1929 311
rect 1923 306 1929 307
rect 2115 311 2121 312
rect 2115 307 2116 311
rect 2120 310 2121 311
rect 2154 311 2160 312
rect 2154 310 2155 311
rect 2120 308 2155 310
rect 2120 307 2121 308
rect 2115 306 2121 307
rect 2154 307 2155 308
rect 2159 307 2160 311
rect 2154 306 2160 307
rect 2331 311 2337 312
rect 2331 307 2332 311
rect 2336 310 2337 311
rect 2362 311 2368 312
rect 2362 310 2363 311
rect 2336 308 2363 310
rect 2336 307 2337 308
rect 2331 306 2337 307
rect 2362 307 2363 308
rect 2367 307 2368 311
rect 2362 306 2368 307
rect 2539 311 2545 312
rect 2539 307 2540 311
rect 2544 310 2545 311
rect 2594 311 2600 312
rect 2594 310 2595 311
rect 2544 308 2595 310
rect 2544 307 2545 308
rect 2539 306 2545 307
rect 2594 307 2595 308
rect 2599 307 2600 311
rect 2594 306 2600 307
rect 2631 311 2637 312
rect 2631 307 2632 311
rect 2636 310 2637 311
rect 2739 311 2745 312
rect 2739 310 2740 311
rect 2636 308 2740 310
rect 2636 307 2637 308
rect 2631 306 2637 307
rect 2739 307 2740 308
rect 2744 307 2745 311
rect 2739 306 2745 307
rect 2854 311 2860 312
rect 2854 307 2855 311
rect 2859 310 2860 311
rect 2931 311 2937 312
rect 2931 310 2932 311
rect 2859 308 2932 310
rect 2859 307 2860 308
rect 2854 306 2860 307
rect 2931 307 2932 308
rect 2936 307 2937 311
rect 2931 306 2937 307
rect 3123 311 3129 312
rect 3123 307 3124 311
rect 3128 310 3129 311
rect 3215 311 3221 312
rect 3215 310 3216 311
rect 3128 308 3216 310
rect 3128 307 3129 308
rect 3123 306 3129 307
rect 3215 307 3216 308
rect 3220 307 3221 311
rect 3215 306 3221 307
rect 3238 311 3244 312
rect 3238 307 3239 311
rect 3243 310 3244 311
rect 3323 311 3329 312
rect 3323 310 3324 311
rect 3243 308 3324 310
rect 3243 307 3244 308
rect 3238 306 3244 307
rect 3323 307 3324 308
rect 3328 307 3329 311
rect 3323 306 3329 307
rect 3515 311 3524 312
rect 3515 307 3516 311
rect 3523 307 3524 311
rect 3515 306 3524 307
rect 214 305 220 306
rect 214 301 215 305
rect 219 301 220 305
rect 214 300 220 301
rect 350 305 356 306
rect 350 301 351 305
rect 355 301 356 305
rect 350 300 356 301
rect 494 305 500 306
rect 494 301 495 305
rect 499 301 500 305
rect 494 300 500 301
rect 638 305 644 306
rect 638 301 639 305
rect 643 301 644 305
rect 638 300 644 301
rect 790 305 796 306
rect 790 301 791 305
rect 795 301 796 305
rect 790 300 796 301
rect 934 305 940 306
rect 934 301 935 305
rect 939 301 940 305
rect 934 300 940 301
rect 1078 305 1084 306
rect 1078 301 1079 305
rect 1083 301 1084 305
rect 1078 300 1084 301
rect 1222 305 1228 306
rect 1222 301 1223 305
rect 1227 301 1228 305
rect 1222 300 1228 301
rect 1358 305 1364 306
rect 1358 301 1359 305
rect 1363 301 1364 305
rect 1358 300 1364 301
rect 1486 305 1492 306
rect 1486 301 1487 305
rect 1491 301 1492 305
rect 1486 300 1492 301
rect 1622 305 1628 306
rect 1622 301 1623 305
rect 1627 301 1628 305
rect 1622 300 1628 301
rect 1734 305 1740 306
rect 1734 301 1735 305
rect 1739 301 1740 305
rect 1734 300 1740 301
rect 1894 301 1900 302
rect 1894 297 1895 301
rect 1899 297 1900 301
rect 1894 296 1900 297
rect 2086 301 2092 302
rect 2086 297 2087 301
rect 2091 297 2092 301
rect 2086 296 2092 297
rect 2302 301 2308 302
rect 2302 297 2303 301
rect 2307 297 2308 301
rect 2302 296 2308 297
rect 2510 301 2516 302
rect 2510 297 2511 301
rect 2515 297 2516 301
rect 2510 296 2516 297
rect 2710 301 2716 302
rect 2710 297 2711 301
rect 2715 297 2716 301
rect 2710 296 2716 297
rect 2902 301 2908 302
rect 2902 297 2903 301
rect 2907 297 2908 301
rect 2902 296 2908 297
rect 3094 301 3100 302
rect 3094 297 3095 301
rect 3099 297 3100 301
rect 3094 296 3100 297
rect 3294 301 3300 302
rect 3294 297 3295 301
rect 3299 297 3300 301
rect 3294 296 3300 297
rect 3486 301 3492 302
rect 3486 297 3487 301
rect 3491 297 3492 301
rect 3486 296 3492 297
rect 110 292 116 293
rect 1822 292 1828 293
rect 110 288 111 292
rect 115 288 116 292
rect 303 291 309 292
rect 303 290 304 291
rect 269 288 304 290
rect 110 287 116 288
rect 303 287 304 288
rect 308 287 309 291
rect 559 291 565 292
rect 559 290 560 291
rect 549 288 560 290
rect 303 286 309 287
rect 559 287 560 288
rect 564 287 565 291
rect 735 291 741 292
rect 735 290 736 291
rect 693 288 736 290
rect 559 286 565 287
rect 735 287 736 288
rect 740 287 741 291
rect 994 291 1000 292
rect 994 290 995 291
rect 989 288 995 290
rect 735 286 741 287
rect 782 287 788 288
rect 782 283 783 287
rect 787 286 788 287
rect 994 287 995 288
rect 999 287 1000 291
rect 1311 291 1317 292
rect 1311 290 1312 291
rect 1277 288 1312 290
rect 994 286 1000 287
rect 1023 287 1029 288
rect 787 284 809 286
rect 787 283 788 284
rect 782 282 788 283
rect 1023 283 1024 287
rect 1028 286 1029 287
rect 1311 287 1312 288
rect 1316 287 1317 291
rect 1423 291 1429 292
rect 1423 290 1424 291
rect 1413 288 1424 290
rect 1311 286 1317 287
rect 1423 287 1424 288
rect 1428 287 1429 291
rect 1695 291 1701 292
rect 1695 290 1696 291
rect 1677 288 1696 290
rect 1423 286 1429 287
rect 1695 287 1696 288
rect 1700 287 1701 291
rect 1807 291 1813 292
rect 1807 290 1808 291
rect 1789 288 1808 290
rect 1695 286 1701 287
rect 1807 287 1808 288
rect 1812 287 1813 291
rect 1822 288 1823 292
rect 1827 288 1828 292
rect 2159 291 2165 292
rect 2159 290 2160 291
rect 1822 287 1828 288
rect 1862 288 1868 289
rect 1807 286 1813 287
rect 1028 284 1097 286
rect 1862 284 1863 288
rect 1867 284 1868 288
rect 2140 288 2160 290
rect 2140 285 2142 288
rect 2159 287 2160 288
rect 2164 287 2165 291
rect 3574 288 3580 289
rect 2159 286 2165 287
rect 2631 287 2637 288
rect 2631 286 2632 287
rect 2565 284 2632 286
rect 1028 283 1029 284
rect 1862 283 1868 284
rect 2154 283 2160 284
rect 1023 282 1029 283
rect 2154 279 2155 283
rect 2159 282 2160 283
rect 2631 283 2632 284
rect 2636 283 2637 287
rect 2854 287 2860 288
rect 2854 286 2855 287
rect 2765 284 2855 286
rect 2631 282 2637 283
rect 2854 283 2855 284
rect 2859 283 2860 287
rect 3154 287 3160 288
rect 3154 286 3155 287
rect 3149 284 3155 286
rect 2854 282 2860 283
rect 3154 283 3155 284
rect 3159 283 3160 287
rect 3574 284 3575 288
rect 3579 284 3580 288
rect 3154 282 3160 283
rect 3215 283 3221 284
rect 3574 283 3580 284
rect 2159 280 2321 282
rect 2159 279 2160 280
rect 2154 278 2160 279
rect 3215 279 3216 283
rect 3220 282 3221 283
rect 3220 280 3313 282
rect 3220 279 3221 280
rect 3215 278 3221 279
rect 110 275 116 276
rect 110 271 111 275
rect 115 271 116 275
rect 110 270 116 271
rect 1470 275 1476 276
rect 1470 271 1471 275
rect 1475 274 1476 275
rect 1822 275 1828 276
rect 1475 272 1497 274
rect 1475 271 1476 272
rect 1470 270 1476 271
rect 1822 271 1823 275
rect 1827 271 1828 275
rect 1822 270 1828 271
rect 1862 271 1868 272
rect 1862 267 1863 271
rect 1867 267 1868 271
rect 2986 271 2992 272
rect 2986 270 2987 271
rect 2953 268 2987 270
rect 1862 266 1868 267
rect 2986 267 2987 268
rect 2991 267 2992 271
rect 2986 266 2992 267
rect 3574 271 3580 272
rect 3574 267 3575 271
rect 3579 267 3580 271
rect 3574 266 3580 267
rect 206 265 212 266
rect 206 261 207 265
rect 211 261 212 265
rect 206 260 212 261
rect 342 265 348 266
rect 342 261 343 265
rect 347 261 348 265
rect 342 260 348 261
rect 486 265 492 266
rect 486 261 487 265
rect 491 261 492 265
rect 486 260 492 261
rect 630 265 636 266
rect 630 261 631 265
rect 635 261 636 265
rect 630 260 636 261
rect 782 265 788 266
rect 782 261 783 265
rect 787 261 788 265
rect 782 260 788 261
rect 926 265 932 266
rect 926 261 927 265
rect 931 261 932 265
rect 926 260 932 261
rect 1070 265 1076 266
rect 1070 261 1071 265
rect 1075 261 1076 265
rect 1070 260 1076 261
rect 1214 265 1220 266
rect 1214 261 1215 265
rect 1219 261 1220 265
rect 1214 260 1220 261
rect 1350 265 1356 266
rect 1350 261 1351 265
rect 1355 261 1356 265
rect 1350 260 1356 261
rect 1478 265 1484 266
rect 1478 261 1479 265
rect 1483 261 1484 265
rect 1478 260 1484 261
rect 1614 265 1620 266
rect 1614 261 1615 265
rect 1619 261 1620 265
rect 1614 260 1620 261
rect 1726 265 1732 266
rect 1726 261 1727 265
rect 1731 261 1732 265
rect 1726 260 1732 261
rect 1886 261 1892 262
rect 391 259 400 260
rect 391 255 392 259
rect 399 255 400 259
rect 1886 257 1887 261
rect 1891 257 1892 261
rect 1886 256 1892 257
rect 2078 261 2084 262
rect 2078 257 2079 261
rect 2083 257 2084 261
rect 2078 256 2084 257
rect 2294 261 2300 262
rect 2294 257 2295 261
rect 2299 257 2300 261
rect 2294 256 2300 257
rect 2502 261 2508 262
rect 2502 257 2503 261
rect 2507 257 2508 261
rect 2502 256 2508 257
rect 2702 261 2708 262
rect 2702 257 2703 261
rect 2707 257 2708 261
rect 2702 256 2708 257
rect 2894 261 2900 262
rect 2894 257 2895 261
rect 2899 257 2900 261
rect 2894 256 2900 257
rect 3086 261 3092 262
rect 3086 257 3087 261
rect 3091 257 3092 261
rect 3086 256 3092 257
rect 3286 261 3292 262
rect 3286 257 3287 261
rect 3291 257 3292 261
rect 3286 256 3292 257
rect 3478 261 3484 262
rect 3478 257 3479 261
rect 3483 257 3484 261
rect 3478 256 3484 257
rect 391 254 400 255
rect 1926 255 1932 256
rect 1926 251 1927 255
rect 1931 254 1932 255
rect 1935 255 1941 256
rect 1935 254 1936 255
rect 1931 252 1936 254
rect 1931 251 1932 252
rect 1926 250 1932 251
rect 1935 251 1936 252
rect 1940 251 1941 255
rect 1935 250 1941 251
rect 3518 255 3524 256
rect 3518 251 3519 255
rect 3523 254 3524 255
rect 3527 255 3533 256
rect 3527 254 3528 255
rect 3523 252 3528 254
rect 3523 251 3524 252
rect 3518 250 3524 251
rect 3527 251 3528 252
rect 3532 251 3533 255
rect 3527 250 3533 251
rect 1886 239 1892 240
rect 230 235 236 236
rect 230 231 231 235
rect 235 231 236 235
rect 230 230 236 231
rect 358 235 364 236
rect 358 231 359 235
rect 363 231 364 235
rect 358 230 364 231
rect 486 235 492 236
rect 486 231 487 235
rect 491 231 492 235
rect 486 230 492 231
rect 622 235 628 236
rect 622 231 623 235
rect 627 231 628 235
rect 622 230 628 231
rect 758 235 764 236
rect 758 231 759 235
rect 763 231 764 235
rect 758 230 764 231
rect 894 235 900 236
rect 894 231 895 235
rect 899 231 900 235
rect 894 230 900 231
rect 1030 235 1036 236
rect 1030 231 1031 235
rect 1035 231 1036 235
rect 1030 230 1036 231
rect 1158 235 1164 236
rect 1158 231 1159 235
rect 1163 231 1164 235
rect 1158 230 1164 231
rect 1294 235 1300 236
rect 1294 231 1295 235
rect 1299 231 1300 235
rect 1294 230 1300 231
rect 1430 235 1436 236
rect 1430 231 1431 235
rect 1435 231 1436 235
rect 1886 235 1887 239
rect 1891 235 1892 239
rect 1886 234 1892 235
rect 1998 239 2004 240
rect 1998 235 1999 239
rect 2003 235 2004 239
rect 1998 234 2004 235
rect 2142 239 2148 240
rect 2142 235 2143 239
rect 2147 235 2148 239
rect 2142 234 2148 235
rect 2294 239 2300 240
rect 2294 235 2295 239
rect 2299 235 2300 239
rect 2294 234 2300 235
rect 2454 239 2460 240
rect 2454 235 2455 239
rect 2459 235 2460 239
rect 2454 234 2460 235
rect 2614 239 2620 240
rect 2614 235 2615 239
rect 2619 235 2620 239
rect 2614 234 2620 235
rect 2782 239 2788 240
rect 2782 235 2783 239
rect 2787 235 2788 239
rect 2782 234 2788 235
rect 2950 239 2956 240
rect 2950 235 2951 239
rect 2955 235 2956 239
rect 2950 234 2956 235
rect 3126 239 3132 240
rect 3126 235 3127 239
rect 3131 235 3132 239
rect 3126 234 3132 235
rect 3310 239 3316 240
rect 3310 235 3311 239
rect 3315 235 3316 239
rect 3310 234 3316 235
rect 3478 239 3484 240
rect 3478 235 3479 239
rect 3483 235 3484 239
rect 3478 234 3484 235
rect 1430 230 1436 231
rect 2078 231 2084 232
rect 1862 229 1868 230
rect 426 227 432 228
rect 110 225 116 226
rect 110 221 111 225
rect 115 221 116 225
rect 426 223 427 227
rect 431 226 432 227
rect 554 227 560 228
rect 431 224 505 226
rect 431 223 432 224
rect 426 222 432 223
rect 554 223 555 227
rect 559 226 560 227
rect 1098 227 1104 228
rect 1098 226 1099 227
rect 559 224 641 226
rect 1089 224 1099 226
rect 559 223 560 224
rect 554 222 560 223
rect 1098 223 1099 224
rect 1103 223 1104 227
rect 1098 222 1104 223
rect 1822 225 1828 226
rect 110 220 116 221
rect 1822 221 1823 225
rect 1827 221 1828 225
rect 1862 225 1863 229
rect 1867 225 1868 229
rect 2078 227 2079 231
rect 2083 230 2084 231
rect 2362 231 2368 232
rect 2362 230 2363 231
rect 2083 228 2161 230
rect 2353 228 2363 230
rect 2083 227 2084 228
rect 2078 226 2084 227
rect 2362 227 2363 228
rect 2367 227 2368 231
rect 3238 231 3244 232
rect 3238 230 3239 231
rect 3185 228 3239 230
rect 2362 226 2368 227
rect 3238 227 3239 228
rect 3243 227 3244 231
rect 3238 226 3244 227
rect 3574 229 3580 230
rect 1862 224 1868 225
rect 3574 225 3575 229
rect 3579 225 3580 229
rect 3574 224 3580 225
rect 1822 220 1828 221
rect 1991 215 1997 216
rect 1991 214 1992 215
rect 1862 212 1868 213
rect 1949 212 1992 214
rect 206 211 212 212
rect 110 208 116 209
rect 110 204 111 208
rect 115 204 116 208
rect 206 207 207 211
rect 211 210 212 211
rect 479 211 485 212
rect 479 210 480 211
rect 211 208 257 210
rect 421 208 480 210
rect 211 207 212 208
rect 206 206 212 207
rect 479 207 480 208
rect 484 207 485 211
rect 479 206 485 207
rect 690 211 696 212
rect 690 207 691 211
rect 695 210 696 211
rect 1023 211 1029 212
rect 1023 210 1024 211
rect 695 208 785 210
rect 957 208 1024 210
rect 695 207 696 208
rect 690 206 696 207
rect 1023 207 1024 208
rect 1028 207 1029 211
rect 1287 211 1293 212
rect 1287 210 1288 211
rect 1221 208 1288 210
rect 1023 206 1029 207
rect 1287 207 1288 208
rect 1292 207 1293 211
rect 1362 211 1368 212
rect 1362 210 1363 211
rect 1357 208 1363 210
rect 1287 206 1293 207
rect 1362 207 1363 208
rect 1367 207 1368 211
rect 1362 206 1368 207
rect 1370 211 1376 212
rect 1370 207 1371 211
rect 1375 210 1376 211
rect 1375 208 1457 210
rect 1822 208 1828 209
rect 1375 207 1376 208
rect 1370 206 1376 207
rect 110 203 116 204
rect 1822 204 1823 208
rect 1827 204 1828 208
rect 1862 208 1863 212
rect 1867 208 1868 212
rect 1991 211 1992 212
rect 1996 211 1997 215
rect 2135 215 2141 216
rect 2135 214 2136 215
rect 2061 212 2136 214
rect 1991 210 1997 211
rect 2135 211 2136 212
rect 2140 211 2141 215
rect 2135 210 2141 211
rect 2362 215 2368 216
rect 2362 211 2363 215
rect 2367 214 2368 215
rect 2682 215 2688 216
rect 2367 212 2481 214
rect 2367 211 2368 212
rect 2362 210 2368 211
rect 1862 207 1868 208
rect 2676 206 2678 213
rect 2682 211 2683 215
rect 2687 214 2688 215
rect 2850 215 2856 216
rect 2687 212 2809 214
rect 2687 211 2688 212
rect 2682 210 2688 211
rect 2850 211 2851 215
rect 2855 214 2856 215
rect 3194 215 3200 216
rect 2855 212 2977 214
rect 2855 211 2856 212
rect 2850 210 2856 211
rect 3194 211 3195 215
rect 3199 214 3200 215
rect 3546 215 3552 216
rect 3546 214 3547 215
rect 3199 212 3337 214
rect 3541 212 3547 214
rect 3199 211 3200 212
rect 3194 210 3200 211
rect 3546 211 3547 212
rect 3551 211 3552 215
rect 3546 210 3552 211
rect 3574 212 3580 213
rect 3574 208 3575 212
rect 3579 208 3580 212
rect 2687 207 2693 208
rect 3574 207 3580 208
rect 2687 206 2688 207
rect 2676 204 2688 206
rect 1822 203 1828 204
rect 2687 203 2688 204
rect 2692 203 2693 207
rect 2687 202 2693 203
rect 1894 199 1900 200
rect 238 195 244 196
rect 238 191 239 195
rect 243 191 244 195
rect 238 190 244 191
rect 366 195 372 196
rect 366 191 367 195
rect 371 191 372 195
rect 494 195 500 196
rect 366 190 372 191
rect 426 191 432 192
rect 426 190 427 191
rect 376 188 427 190
rect 376 186 378 188
rect 426 187 427 188
rect 431 187 432 191
rect 494 191 495 195
rect 499 191 500 195
rect 494 190 500 191
rect 630 195 636 196
rect 630 191 631 195
rect 635 191 636 195
rect 630 190 636 191
rect 766 195 772 196
rect 766 191 767 195
rect 771 191 772 195
rect 766 190 772 191
rect 902 195 908 196
rect 902 191 903 195
rect 907 191 908 195
rect 902 190 908 191
rect 1038 195 1044 196
rect 1038 191 1039 195
rect 1043 191 1044 195
rect 1038 190 1044 191
rect 1166 195 1172 196
rect 1166 191 1167 195
rect 1171 191 1172 195
rect 1166 190 1172 191
rect 1302 195 1308 196
rect 1302 191 1303 195
rect 1307 191 1308 195
rect 1302 190 1308 191
rect 1438 195 1444 196
rect 1438 191 1439 195
rect 1443 191 1444 195
rect 1894 195 1895 199
rect 1899 195 1900 199
rect 1894 194 1900 195
rect 2006 199 2012 200
rect 2006 195 2007 199
rect 2011 195 2012 199
rect 2006 194 2012 195
rect 2150 199 2156 200
rect 2150 195 2151 199
rect 2155 195 2156 199
rect 2150 194 2156 195
rect 2302 199 2308 200
rect 2302 195 2303 199
rect 2307 195 2308 199
rect 2302 194 2308 195
rect 2462 199 2468 200
rect 2462 195 2463 199
rect 2467 195 2468 199
rect 2462 194 2468 195
rect 2622 199 2628 200
rect 2622 195 2623 199
rect 2627 195 2628 199
rect 2622 194 2628 195
rect 2790 199 2796 200
rect 2790 195 2791 199
rect 2795 195 2796 199
rect 2790 194 2796 195
rect 2958 199 2964 200
rect 2958 195 2959 199
rect 2963 195 2964 199
rect 2958 194 2964 195
rect 3134 199 3140 200
rect 3134 195 3135 199
rect 3139 195 3140 199
rect 3134 194 3140 195
rect 3318 199 3324 200
rect 3318 195 3319 199
rect 3323 195 3324 199
rect 3318 194 3324 195
rect 3486 199 3492 200
rect 3486 195 3487 199
rect 3491 195 3492 199
rect 3486 194 3492 195
rect 1438 190 1444 191
rect 426 186 432 187
rect 1923 187 1932 188
rect 267 185 378 186
rect 267 181 268 185
rect 272 184 378 185
rect 272 181 273 184
rect 267 180 273 181
rect 394 183 401 184
rect 394 179 395 183
rect 400 179 401 183
rect 394 178 401 179
rect 479 183 485 184
rect 479 179 480 183
rect 484 182 485 183
rect 523 183 529 184
rect 523 182 524 183
rect 484 180 524 182
rect 484 179 485 180
rect 479 178 485 179
rect 523 179 524 180
rect 528 179 529 183
rect 523 178 529 179
rect 659 183 665 184
rect 659 179 660 183
rect 664 182 665 183
rect 690 183 696 184
rect 690 182 691 183
rect 664 180 691 182
rect 664 179 665 180
rect 659 178 665 179
rect 690 179 691 180
rect 695 179 696 183
rect 690 178 696 179
rect 782 183 788 184
rect 782 179 783 183
rect 787 182 788 183
rect 795 183 801 184
rect 795 182 796 183
rect 787 180 796 182
rect 787 179 788 180
rect 782 178 788 179
rect 795 179 796 180
rect 800 179 801 183
rect 795 178 801 179
rect 931 183 940 184
rect 931 179 932 183
rect 939 179 940 183
rect 931 178 940 179
rect 1023 183 1029 184
rect 1023 179 1024 183
rect 1028 182 1029 183
rect 1067 183 1073 184
rect 1067 182 1068 183
rect 1028 180 1068 182
rect 1028 179 1029 180
rect 1023 178 1029 179
rect 1067 179 1068 180
rect 1072 179 1073 183
rect 1067 178 1073 179
rect 1195 183 1201 184
rect 1195 179 1196 183
rect 1200 182 1201 183
rect 1287 183 1293 184
rect 1200 180 1278 182
rect 1200 179 1201 180
rect 1195 178 1201 179
rect 1276 174 1278 180
rect 1287 179 1288 183
rect 1292 182 1293 183
rect 1331 183 1337 184
rect 1331 182 1332 183
rect 1292 180 1332 182
rect 1292 179 1293 180
rect 1287 178 1293 179
rect 1331 179 1332 180
rect 1336 179 1337 183
rect 1331 178 1337 179
rect 1467 183 1476 184
rect 1467 179 1468 183
rect 1475 179 1476 183
rect 1923 183 1924 187
rect 1931 183 1932 187
rect 1923 182 1932 183
rect 1991 187 1997 188
rect 1991 183 1992 187
rect 1996 186 1997 187
rect 2035 187 2041 188
rect 2035 186 2036 187
rect 1996 184 2036 186
rect 1996 183 1997 184
rect 1991 182 1997 183
rect 2035 183 2036 184
rect 2040 183 2041 187
rect 2035 182 2041 183
rect 2135 187 2141 188
rect 2135 183 2136 187
rect 2140 186 2141 187
rect 2179 187 2185 188
rect 2179 186 2180 187
rect 2140 184 2180 186
rect 2140 183 2141 184
rect 2135 182 2141 183
rect 2179 183 2180 184
rect 2184 183 2185 187
rect 2179 182 2185 183
rect 2331 187 2337 188
rect 2331 183 2332 187
rect 2336 186 2337 187
rect 2362 187 2368 188
rect 2362 186 2363 187
rect 2336 184 2363 186
rect 2336 183 2337 184
rect 2331 182 2337 183
rect 2362 183 2363 184
rect 2367 183 2368 187
rect 2362 182 2368 183
rect 2491 187 2497 188
rect 2491 183 2492 187
rect 2496 186 2497 187
rect 2506 187 2512 188
rect 2506 186 2507 187
rect 2496 184 2507 186
rect 2496 183 2497 184
rect 2491 182 2497 183
rect 2506 183 2507 184
rect 2511 183 2512 187
rect 2506 182 2512 183
rect 2651 187 2657 188
rect 2651 183 2652 187
rect 2656 186 2657 187
rect 2682 187 2688 188
rect 2682 186 2683 187
rect 2656 184 2683 186
rect 2656 183 2657 184
rect 2651 182 2657 183
rect 2682 183 2683 184
rect 2687 183 2688 187
rect 2682 182 2688 183
rect 2819 187 2825 188
rect 2819 183 2820 187
rect 2824 186 2825 187
rect 2850 187 2856 188
rect 2850 186 2851 187
rect 2824 184 2851 186
rect 2824 183 2825 184
rect 2819 182 2825 183
rect 2850 183 2851 184
rect 2855 183 2856 187
rect 2850 182 2856 183
rect 2986 187 2993 188
rect 2986 183 2987 187
rect 2992 183 2993 187
rect 2986 182 2993 183
rect 3163 187 3169 188
rect 3163 183 3164 187
rect 3168 186 3169 187
rect 3194 187 3200 188
rect 3194 186 3195 187
rect 3168 184 3195 186
rect 3168 183 3169 184
rect 3163 182 3169 183
rect 3194 183 3195 184
rect 3199 183 3200 187
rect 3194 182 3200 183
rect 3347 187 3353 188
rect 3347 183 3348 187
rect 3352 186 3353 187
rect 3370 187 3376 188
rect 3370 186 3371 187
rect 3352 184 3371 186
rect 3352 183 3353 184
rect 3347 182 3353 183
rect 3370 183 3371 184
rect 3375 183 3376 187
rect 3370 182 3376 183
rect 3515 187 3524 188
rect 3515 183 3516 187
rect 3523 183 3524 187
rect 3515 182 3524 183
rect 1467 178 1476 179
rect 1370 175 1376 176
rect 1370 174 1371 175
rect 1276 172 1371 174
rect 1370 171 1371 172
rect 1375 171 1376 175
rect 1370 170 1376 171
rect 1479 155 1485 156
rect 1479 154 1480 155
rect 1260 152 1480 154
rect 1260 150 1262 152
rect 1479 151 1480 152
rect 1484 151 1485 155
rect 2078 155 2084 156
rect 2078 154 2079 155
rect 1479 150 1485 151
rect 1924 152 2079 154
rect 1924 150 1926 152
rect 2078 151 2079 152
rect 2083 151 2084 155
rect 2078 150 2084 151
rect 1259 149 1265 150
rect 203 147 212 148
rect 203 143 204 147
rect 211 143 212 147
rect 203 142 212 143
rect 239 147 245 148
rect 239 143 240 147
rect 244 146 245 147
rect 291 147 297 148
rect 291 146 292 147
rect 244 144 292 146
rect 244 143 245 144
rect 239 142 245 143
rect 291 143 292 144
rect 296 143 297 147
rect 291 142 297 143
rect 327 147 333 148
rect 327 143 328 147
rect 332 146 333 147
rect 379 147 385 148
rect 379 146 380 147
rect 332 144 380 146
rect 332 143 333 144
rect 327 142 333 143
rect 379 143 380 144
rect 384 143 385 147
rect 379 142 385 143
rect 415 147 421 148
rect 415 143 416 147
rect 420 146 421 147
rect 467 147 473 148
rect 467 146 468 147
rect 420 144 468 146
rect 420 143 421 144
rect 415 142 421 143
rect 467 143 468 144
rect 472 143 473 147
rect 467 142 473 143
rect 503 147 509 148
rect 503 143 504 147
rect 508 146 509 147
rect 555 147 561 148
rect 555 146 556 147
rect 508 144 556 146
rect 508 143 509 144
rect 503 142 509 143
rect 555 143 556 144
rect 560 143 561 147
rect 555 142 561 143
rect 591 147 597 148
rect 591 143 592 147
rect 596 146 597 147
rect 643 147 649 148
rect 643 146 644 147
rect 596 144 644 146
rect 596 143 597 144
rect 591 142 597 143
rect 643 143 644 144
rect 648 143 649 147
rect 643 142 649 143
rect 679 147 685 148
rect 679 143 680 147
rect 684 146 685 147
rect 731 147 737 148
rect 731 146 732 147
rect 684 144 732 146
rect 684 143 685 144
rect 679 142 685 143
rect 731 143 732 144
rect 736 143 737 147
rect 731 142 737 143
rect 767 147 773 148
rect 767 143 768 147
rect 772 146 773 147
rect 819 147 825 148
rect 819 146 820 147
rect 772 144 820 146
rect 772 143 773 144
rect 767 142 773 143
rect 819 143 820 144
rect 824 143 825 147
rect 819 142 825 143
rect 907 147 913 148
rect 907 143 908 147
rect 912 146 913 147
rect 946 147 952 148
rect 946 146 947 147
rect 912 144 947 146
rect 912 143 913 144
rect 907 142 913 143
rect 946 143 947 144
rect 951 143 952 147
rect 946 142 952 143
rect 995 147 1001 148
rect 995 143 996 147
rect 1000 146 1001 147
rect 1039 147 1045 148
rect 1039 146 1040 147
rect 1000 144 1040 146
rect 1000 143 1001 144
rect 995 142 1001 143
rect 1039 143 1040 144
rect 1044 143 1045 147
rect 1039 142 1045 143
rect 1083 147 1089 148
rect 1083 143 1084 147
rect 1088 146 1089 147
rect 1122 147 1128 148
rect 1122 146 1123 147
rect 1088 144 1123 146
rect 1088 143 1089 144
rect 1083 142 1089 143
rect 1122 143 1123 144
rect 1127 143 1128 147
rect 1122 142 1128 143
rect 1171 147 1177 148
rect 1171 143 1172 147
rect 1176 146 1177 147
rect 1210 147 1216 148
rect 1210 146 1211 147
rect 1176 144 1211 146
rect 1176 143 1177 144
rect 1171 142 1177 143
rect 1210 143 1211 144
rect 1215 143 1216 147
rect 1259 145 1260 149
rect 1264 145 1265 149
rect 1923 149 1929 150
rect 1259 144 1265 145
rect 1347 147 1353 148
rect 1210 142 1216 143
rect 1347 143 1348 147
rect 1352 146 1353 147
rect 1362 147 1368 148
rect 1362 146 1363 147
rect 1352 144 1363 146
rect 1352 143 1353 144
rect 1347 142 1353 143
rect 1362 143 1363 144
rect 1367 143 1368 147
rect 1362 142 1368 143
rect 1383 147 1389 148
rect 1383 143 1384 147
rect 1388 146 1389 147
rect 1435 147 1441 148
rect 1435 146 1436 147
rect 1388 144 1436 146
rect 1388 143 1389 144
rect 1383 142 1389 143
rect 1435 143 1436 144
rect 1440 143 1441 147
rect 1435 142 1441 143
rect 1471 147 1477 148
rect 1471 143 1472 147
rect 1476 146 1477 147
rect 1531 147 1537 148
rect 1531 146 1532 147
rect 1476 144 1532 146
rect 1476 143 1477 144
rect 1471 142 1477 143
rect 1531 143 1532 144
rect 1536 143 1537 147
rect 1923 145 1924 149
rect 1928 145 1929 149
rect 1923 144 1929 145
rect 1967 147 1973 148
rect 1531 142 1537 143
rect 1967 143 1968 147
rect 1972 146 1973 147
rect 2011 147 2017 148
rect 2011 146 2012 147
rect 1972 144 2012 146
rect 1972 143 1973 144
rect 1967 142 1973 143
rect 2011 143 2012 144
rect 2016 143 2017 147
rect 2011 142 2017 143
rect 2047 147 2053 148
rect 2047 143 2048 147
rect 2052 146 2053 147
rect 2099 147 2105 148
rect 2099 146 2100 147
rect 2052 144 2100 146
rect 2052 143 2053 144
rect 2047 142 2053 143
rect 2099 143 2100 144
rect 2104 143 2105 147
rect 2099 142 2105 143
rect 2135 147 2141 148
rect 2135 143 2136 147
rect 2140 146 2141 147
rect 2187 147 2193 148
rect 2187 146 2188 147
rect 2140 144 2188 146
rect 2140 143 2141 144
rect 2135 142 2141 143
rect 2187 143 2188 144
rect 2192 143 2193 147
rect 2187 142 2193 143
rect 2223 147 2229 148
rect 2223 143 2224 147
rect 2228 146 2229 147
rect 2275 147 2281 148
rect 2275 146 2276 147
rect 2228 144 2276 146
rect 2228 143 2229 144
rect 2223 142 2229 143
rect 2275 143 2276 144
rect 2280 143 2281 147
rect 2275 142 2281 143
rect 2311 147 2317 148
rect 2311 143 2312 147
rect 2316 146 2317 147
rect 2363 147 2369 148
rect 2363 146 2364 147
rect 2316 144 2364 146
rect 2316 143 2317 144
rect 2311 142 2317 143
rect 2363 143 2364 144
rect 2368 143 2369 147
rect 2363 142 2369 143
rect 2407 147 2413 148
rect 2407 143 2408 147
rect 2412 146 2413 147
rect 2467 147 2473 148
rect 2467 146 2468 147
rect 2412 144 2468 146
rect 2412 143 2413 144
rect 2407 142 2413 143
rect 2467 143 2468 144
rect 2472 143 2473 147
rect 2467 142 2473 143
rect 2498 147 2504 148
rect 2498 143 2499 147
rect 2503 146 2504 147
rect 2571 147 2577 148
rect 2571 146 2572 147
rect 2503 144 2572 146
rect 2503 143 2504 144
rect 2498 142 2504 143
rect 2571 143 2572 144
rect 2576 143 2577 147
rect 2571 142 2577 143
rect 2675 147 2681 148
rect 2675 143 2676 147
rect 2680 146 2681 147
rect 2687 147 2693 148
rect 2687 146 2688 147
rect 2680 144 2688 146
rect 2680 143 2681 144
rect 2675 142 2681 143
rect 2687 143 2688 144
rect 2692 143 2693 147
rect 2687 142 2693 143
rect 2711 147 2717 148
rect 2711 143 2712 147
rect 2716 146 2717 147
rect 2771 147 2777 148
rect 2771 146 2772 147
rect 2716 144 2772 146
rect 2716 143 2717 144
rect 2711 142 2717 143
rect 2771 143 2772 144
rect 2776 143 2777 147
rect 2771 142 2777 143
rect 2823 147 2829 148
rect 2823 143 2824 147
rect 2828 146 2829 147
rect 2867 147 2873 148
rect 2867 146 2868 147
rect 2828 144 2868 146
rect 2828 143 2829 144
rect 2823 142 2829 143
rect 2867 143 2868 144
rect 2872 143 2873 147
rect 2867 142 2873 143
rect 2903 147 2909 148
rect 2903 143 2904 147
rect 2908 146 2909 147
rect 2963 147 2969 148
rect 2963 146 2964 147
rect 2908 144 2964 146
rect 2908 143 2909 144
rect 2903 142 2909 143
rect 2963 143 2964 144
rect 2968 143 2969 147
rect 2963 142 2969 143
rect 2999 147 3005 148
rect 2999 143 3000 147
rect 3004 146 3005 147
rect 3059 147 3065 148
rect 3059 146 3060 147
rect 3004 144 3060 146
rect 3004 143 3005 144
rect 2999 142 3005 143
rect 3059 143 3060 144
rect 3064 143 3065 147
rect 3059 142 3065 143
rect 3095 147 3101 148
rect 3095 143 3096 147
rect 3100 146 3101 147
rect 3155 147 3161 148
rect 3155 146 3156 147
rect 3100 144 3156 146
rect 3100 143 3101 144
rect 3095 142 3101 143
rect 3155 143 3156 144
rect 3160 143 3161 147
rect 3155 142 3161 143
rect 3191 147 3197 148
rect 3191 143 3192 147
rect 3196 146 3197 147
rect 3251 147 3257 148
rect 3251 146 3252 147
rect 3196 144 3252 146
rect 3196 143 3197 144
rect 3191 142 3197 143
rect 3251 143 3252 144
rect 3256 143 3257 147
rect 3251 142 3257 143
rect 3287 147 3293 148
rect 3287 143 3288 147
rect 3292 146 3293 147
rect 3339 147 3345 148
rect 3339 146 3340 147
rect 3292 144 3340 146
rect 3292 143 3293 144
rect 3287 142 3293 143
rect 3339 143 3340 144
rect 3344 143 3345 147
rect 3339 142 3345 143
rect 3427 147 3433 148
rect 3427 143 3428 147
rect 3432 146 3433 147
rect 3466 147 3472 148
rect 3466 146 3467 147
rect 3432 144 3467 146
rect 3432 143 3433 144
rect 3427 142 3433 143
rect 3466 143 3467 144
rect 3471 143 3472 147
rect 3466 142 3472 143
rect 3515 147 3521 148
rect 3515 143 3516 147
rect 3520 146 3521 147
rect 3546 147 3552 148
rect 3546 146 3547 147
rect 3520 144 3547 146
rect 3520 143 3521 144
rect 3515 142 3521 143
rect 3546 143 3547 144
rect 3551 143 3552 147
rect 3546 142 3552 143
rect 174 137 180 138
rect 174 133 175 137
rect 179 133 180 137
rect 174 132 180 133
rect 262 137 268 138
rect 262 133 263 137
rect 267 133 268 137
rect 262 132 268 133
rect 350 137 356 138
rect 350 133 351 137
rect 355 133 356 137
rect 350 132 356 133
rect 438 137 444 138
rect 438 133 439 137
rect 443 133 444 137
rect 438 132 444 133
rect 526 137 532 138
rect 526 133 527 137
rect 531 133 532 137
rect 526 132 532 133
rect 614 137 620 138
rect 614 133 615 137
rect 619 133 620 137
rect 614 132 620 133
rect 702 137 708 138
rect 702 133 703 137
rect 707 133 708 137
rect 702 132 708 133
rect 790 137 796 138
rect 790 133 791 137
rect 795 133 796 137
rect 790 132 796 133
rect 878 137 884 138
rect 878 133 879 137
rect 883 133 884 137
rect 878 132 884 133
rect 966 137 972 138
rect 966 133 967 137
rect 971 133 972 137
rect 966 132 972 133
rect 1054 137 1060 138
rect 1054 133 1055 137
rect 1059 133 1060 137
rect 1054 132 1060 133
rect 1142 137 1148 138
rect 1142 133 1143 137
rect 1147 133 1148 137
rect 1142 132 1148 133
rect 1230 137 1236 138
rect 1230 133 1231 137
rect 1235 133 1236 137
rect 1230 132 1236 133
rect 1318 137 1324 138
rect 1318 133 1319 137
rect 1323 133 1324 137
rect 1318 132 1324 133
rect 1406 137 1412 138
rect 1406 133 1407 137
rect 1411 133 1412 137
rect 1406 132 1412 133
rect 1502 137 1508 138
rect 1502 133 1503 137
rect 1507 133 1508 137
rect 1502 132 1508 133
rect 1894 137 1900 138
rect 1894 133 1895 137
rect 1899 133 1900 137
rect 1894 132 1900 133
rect 1982 137 1988 138
rect 1982 133 1983 137
rect 1987 133 1988 137
rect 1982 132 1988 133
rect 2070 137 2076 138
rect 2070 133 2071 137
rect 2075 133 2076 137
rect 2070 132 2076 133
rect 2158 137 2164 138
rect 2158 133 2159 137
rect 2163 133 2164 137
rect 2158 132 2164 133
rect 2246 137 2252 138
rect 2246 133 2247 137
rect 2251 133 2252 137
rect 2246 132 2252 133
rect 2334 137 2340 138
rect 2334 133 2335 137
rect 2339 133 2340 137
rect 2334 132 2340 133
rect 2438 137 2444 138
rect 2438 133 2439 137
rect 2443 133 2444 137
rect 2438 132 2444 133
rect 2542 137 2548 138
rect 2542 133 2543 137
rect 2547 133 2548 137
rect 2542 132 2548 133
rect 2646 137 2652 138
rect 2646 133 2647 137
rect 2651 133 2652 137
rect 2646 132 2652 133
rect 2742 137 2748 138
rect 2742 133 2743 137
rect 2747 133 2748 137
rect 2742 132 2748 133
rect 2838 137 2844 138
rect 2838 133 2839 137
rect 2843 133 2844 137
rect 2838 132 2844 133
rect 2934 137 2940 138
rect 2934 133 2935 137
rect 2939 133 2940 137
rect 2934 132 2940 133
rect 3030 137 3036 138
rect 3030 133 3031 137
rect 3035 133 3036 137
rect 3030 132 3036 133
rect 3126 137 3132 138
rect 3126 133 3127 137
rect 3131 133 3132 137
rect 3126 132 3132 133
rect 3222 137 3228 138
rect 3222 133 3223 137
rect 3227 133 3228 137
rect 3222 132 3228 133
rect 3310 137 3316 138
rect 3310 133 3311 137
rect 3315 133 3316 137
rect 3310 132 3316 133
rect 3398 137 3404 138
rect 3398 133 3399 137
rect 3403 133 3404 137
rect 3398 132 3404 133
rect 3486 137 3492 138
rect 3486 133 3487 137
rect 3491 133 3492 137
rect 3486 132 3492 133
rect 934 131 940 132
rect 934 130 935 131
rect 932 127 935 130
rect 939 127 940 131
rect 932 126 940 127
rect 110 124 116 125
rect 110 120 111 124
rect 115 120 116 124
rect 239 123 245 124
rect 239 122 240 123
rect 229 120 240 122
rect 110 119 116 120
rect 239 119 240 120
rect 244 119 245 123
rect 327 123 333 124
rect 327 122 328 123
rect 317 120 328 122
rect 239 118 245 119
rect 327 119 328 120
rect 332 119 333 123
rect 415 123 421 124
rect 415 122 416 123
rect 405 120 416 122
rect 327 118 333 119
rect 415 119 416 120
rect 420 119 421 123
rect 503 123 509 124
rect 503 122 504 123
rect 493 120 504 122
rect 415 118 421 119
rect 503 119 504 120
rect 508 119 509 123
rect 591 123 597 124
rect 591 122 592 123
rect 581 120 592 122
rect 503 118 509 119
rect 591 119 592 120
rect 596 119 597 123
rect 679 123 685 124
rect 679 122 680 123
rect 669 120 680 122
rect 591 118 597 119
rect 679 119 680 120
rect 684 119 685 123
rect 767 123 773 124
rect 767 122 768 123
rect 757 120 768 122
rect 679 118 685 119
rect 767 119 768 120
rect 772 119 773 123
rect 932 121 934 126
rect 1822 124 1828 125
rect 1383 123 1389 124
rect 1383 122 1384 123
rect 1373 120 1384 122
rect 767 118 773 119
rect 782 119 788 120
rect 782 115 783 119
rect 787 118 788 119
rect 946 119 952 120
rect 787 116 809 118
rect 787 115 788 116
rect 782 114 788 115
rect 946 115 947 119
rect 951 118 952 119
rect 1039 119 1045 120
rect 951 116 985 118
rect 951 115 952 116
rect 946 114 952 115
rect 1039 115 1040 119
rect 1044 118 1045 119
rect 1122 119 1128 120
rect 1044 116 1073 118
rect 1044 115 1045 116
rect 1039 114 1045 115
rect 1122 115 1123 119
rect 1127 118 1128 119
rect 1210 119 1216 120
rect 1127 116 1161 118
rect 1127 115 1128 116
rect 1122 114 1128 115
rect 1210 115 1211 119
rect 1215 118 1216 119
rect 1383 119 1384 120
rect 1388 119 1389 123
rect 1471 123 1477 124
rect 1471 122 1472 123
rect 1461 120 1472 122
rect 1383 118 1389 119
rect 1471 119 1472 120
rect 1476 119 1477 123
rect 1822 120 1823 124
rect 1827 120 1828 124
rect 1471 118 1477 119
rect 1479 119 1485 120
rect 1822 119 1828 120
rect 1862 124 1868 125
rect 3574 124 3580 125
rect 1862 120 1863 124
rect 1867 120 1868 124
rect 1967 123 1973 124
rect 1967 122 1968 123
rect 1949 120 1968 122
rect 1862 119 1868 120
rect 1967 119 1968 120
rect 1972 119 1973 123
rect 2047 123 2053 124
rect 2047 122 2048 123
rect 2037 120 2048 122
rect 1215 116 1249 118
rect 1215 115 1216 116
rect 1210 114 1216 115
rect 1479 115 1480 119
rect 1484 118 1485 119
rect 1967 118 1973 119
rect 2047 119 2048 120
rect 2052 119 2053 123
rect 2135 123 2141 124
rect 2135 122 2136 123
rect 2125 120 2136 122
rect 2047 118 2053 119
rect 2135 119 2136 120
rect 2140 119 2141 123
rect 2223 123 2229 124
rect 2223 122 2224 123
rect 2213 120 2224 122
rect 2135 118 2141 119
rect 2223 119 2224 120
rect 2228 119 2229 123
rect 2311 123 2317 124
rect 2311 122 2312 123
rect 2301 120 2312 122
rect 2223 118 2229 119
rect 2311 119 2312 120
rect 2316 119 2317 123
rect 2407 123 2413 124
rect 2407 122 2408 123
rect 2389 120 2408 122
rect 2311 118 2317 119
rect 2407 119 2408 120
rect 2412 119 2413 123
rect 2498 123 2504 124
rect 2498 122 2499 123
rect 2493 120 2499 122
rect 2407 118 2413 119
rect 2498 119 2499 120
rect 2503 119 2504 123
rect 2711 123 2717 124
rect 2711 122 2712 123
rect 2701 120 2712 122
rect 2498 118 2504 119
rect 2506 119 2512 120
rect 1484 116 1521 118
rect 1484 115 1485 116
rect 1479 114 1485 115
rect 2506 115 2507 119
rect 2511 118 2512 119
rect 2711 119 2712 120
rect 2716 119 2717 123
rect 2823 123 2829 124
rect 2823 122 2824 123
rect 2797 120 2824 122
rect 2711 118 2717 119
rect 2823 119 2824 120
rect 2828 119 2829 123
rect 2903 123 2909 124
rect 2903 122 2904 123
rect 2893 120 2904 122
rect 2823 118 2829 119
rect 2903 119 2904 120
rect 2908 119 2909 123
rect 2999 123 3005 124
rect 2999 122 3000 123
rect 2989 120 3000 122
rect 2903 118 2909 119
rect 2999 119 3000 120
rect 3004 119 3005 123
rect 3095 123 3101 124
rect 3095 122 3096 123
rect 3085 120 3096 122
rect 2999 118 3005 119
rect 3095 119 3096 120
rect 3100 119 3101 123
rect 3191 123 3197 124
rect 3191 122 3192 123
rect 3181 120 3192 122
rect 3095 118 3101 119
rect 3191 119 3192 120
rect 3196 119 3197 123
rect 3287 123 3293 124
rect 3287 122 3288 123
rect 3277 120 3288 122
rect 3191 118 3197 119
rect 3287 119 3288 120
rect 3292 119 3293 123
rect 3370 123 3376 124
rect 3370 122 3371 123
rect 3365 120 3371 122
rect 3287 118 3293 119
rect 3370 119 3371 120
rect 3375 119 3376 123
rect 3574 120 3575 124
rect 3579 120 3580 124
rect 3370 118 3376 119
rect 3466 119 3472 120
rect 3574 119 3580 120
rect 2511 116 2561 118
rect 2511 115 2512 116
rect 2506 114 2512 115
rect 3466 115 3467 119
rect 3471 118 3472 119
rect 3471 116 3505 118
rect 3471 115 3472 116
rect 3466 114 3472 115
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 110 102 116 103
rect 1822 107 1828 108
rect 1822 103 1823 107
rect 1827 103 1828 107
rect 1822 102 1828 103
rect 1862 107 1868 108
rect 1862 103 1863 107
rect 1867 103 1868 107
rect 1862 102 1868 103
rect 3574 107 3580 108
rect 3574 103 3575 107
rect 3579 103 3580 107
rect 3574 102 3580 103
rect 166 97 172 98
rect 166 93 167 97
rect 171 93 172 97
rect 166 92 172 93
rect 254 97 260 98
rect 254 93 255 97
rect 259 93 260 97
rect 254 92 260 93
rect 342 97 348 98
rect 342 93 343 97
rect 347 93 348 97
rect 342 92 348 93
rect 430 97 436 98
rect 430 93 431 97
rect 435 93 436 97
rect 430 92 436 93
rect 518 97 524 98
rect 518 93 519 97
rect 523 93 524 97
rect 518 92 524 93
rect 606 97 612 98
rect 606 93 607 97
rect 611 93 612 97
rect 606 92 612 93
rect 694 97 700 98
rect 694 93 695 97
rect 699 93 700 97
rect 694 92 700 93
rect 782 97 788 98
rect 782 93 783 97
rect 787 93 788 97
rect 782 92 788 93
rect 870 97 876 98
rect 870 93 871 97
rect 875 93 876 97
rect 870 92 876 93
rect 958 97 964 98
rect 958 93 959 97
rect 963 93 964 97
rect 958 92 964 93
rect 1046 97 1052 98
rect 1046 93 1047 97
rect 1051 93 1052 97
rect 1046 92 1052 93
rect 1134 97 1140 98
rect 1134 93 1135 97
rect 1139 93 1140 97
rect 1134 92 1140 93
rect 1222 97 1228 98
rect 1222 93 1223 97
rect 1227 93 1228 97
rect 1222 92 1228 93
rect 1310 97 1316 98
rect 1310 93 1311 97
rect 1315 93 1316 97
rect 1310 92 1316 93
rect 1398 97 1404 98
rect 1398 93 1399 97
rect 1403 93 1404 97
rect 1398 92 1404 93
rect 1494 97 1500 98
rect 1494 93 1495 97
rect 1499 93 1500 97
rect 1494 92 1500 93
rect 1886 97 1892 98
rect 1886 93 1887 97
rect 1891 93 1892 97
rect 1886 92 1892 93
rect 1974 97 1980 98
rect 1974 93 1975 97
rect 1979 93 1980 97
rect 1974 92 1980 93
rect 2062 97 2068 98
rect 2062 93 2063 97
rect 2067 93 2068 97
rect 2062 92 2068 93
rect 2150 97 2156 98
rect 2150 93 2151 97
rect 2155 93 2156 97
rect 2150 92 2156 93
rect 2238 97 2244 98
rect 2238 93 2239 97
rect 2243 93 2244 97
rect 2238 92 2244 93
rect 2326 97 2332 98
rect 2326 93 2327 97
rect 2331 93 2332 97
rect 2326 92 2332 93
rect 2430 97 2436 98
rect 2430 93 2431 97
rect 2435 93 2436 97
rect 2430 92 2436 93
rect 2534 97 2540 98
rect 2534 93 2535 97
rect 2539 93 2540 97
rect 2534 92 2540 93
rect 2638 97 2644 98
rect 2638 93 2639 97
rect 2643 93 2644 97
rect 2638 92 2644 93
rect 2734 97 2740 98
rect 2734 93 2735 97
rect 2739 93 2740 97
rect 2734 92 2740 93
rect 2830 97 2836 98
rect 2830 93 2831 97
rect 2835 93 2836 97
rect 2830 92 2836 93
rect 2926 97 2932 98
rect 2926 93 2927 97
rect 2931 93 2932 97
rect 2926 92 2932 93
rect 3022 97 3028 98
rect 3022 93 3023 97
rect 3027 93 3028 97
rect 3022 92 3028 93
rect 3118 97 3124 98
rect 3118 93 3119 97
rect 3123 93 3124 97
rect 3118 92 3124 93
rect 3214 97 3220 98
rect 3214 93 3215 97
rect 3219 93 3220 97
rect 3214 92 3220 93
rect 3302 97 3308 98
rect 3302 93 3303 97
rect 3307 93 3308 97
rect 3302 92 3308 93
rect 3390 97 3396 98
rect 3390 93 3391 97
rect 3395 93 3396 97
rect 3390 92 3396 93
rect 3478 97 3484 98
rect 3478 93 3479 97
rect 3483 93 3484 97
rect 3478 92 3484 93
<< m3c >>
rect 307 3639 311 3643
rect 395 3639 399 3643
rect 483 3639 487 3643
rect 571 3639 575 3643
rect 659 3639 663 3643
rect 239 3629 243 3633
rect 327 3629 331 3633
rect 415 3629 419 3633
rect 503 3629 507 3633
rect 591 3629 595 3633
rect 679 3629 683 3633
rect 111 3616 115 3620
rect 1823 3616 1827 3620
rect 307 3611 311 3615
rect 395 3611 399 3615
rect 483 3611 487 3615
rect 571 3611 575 3615
rect 659 3611 663 3615
rect 111 3599 115 3603
rect 1823 3599 1827 3603
rect 231 3589 235 3593
rect 319 3589 323 3593
rect 407 3589 411 3593
rect 495 3589 499 3593
rect 583 3589 587 3593
rect 671 3589 675 3593
rect 283 3583 284 3587
rect 284 3583 287 3587
rect 1887 3571 1891 3575
rect 1975 3571 1979 3575
rect 2063 3571 2067 3575
rect 2151 3571 2155 3575
rect 2239 3571 2243 3575
rect 2327 3571 2331 3575
rect 2415 3571 2419 3575
rect 2503 3571 2507 3575
rect 2591 3571 2595 3575
rect 2679 3571 2683 3575
rect 2767 3571 2771 3575
rect 2855 3571 2859 3575
rect 2943 3571 2947 3575
rect 3031 3571 3035 3575
rect 3119 3571 3123 3575
rect 3207 3571 3211 3575
rect 3295 3571 3299 3575
rect 247 3559 251 3563
rect 399 3559 403 3563
rect 543 3559 547 3563
rect 687 3559 691 3563
rect 823 3559 827 3563
rect 951 3559 955 3563
rect 1079 3559 1083 3563
rect 1199 3559 1203 3563
rect 1311 3559 1315 3563
rect 1423 3559 1427 3563
rect 1543 3559 1547 3563
rect 1863 3561 1867 3565
rect 3275 3563 3279 3567
rect 3575 3561 3579 3565
rect 111 3549 115 3553
rect 1491 3551 1495 3555
rect 1823 3549 1827 3553
rect 1863 3544 1867 3548
rect 2571 3547 2575 3551
rect 3575 3544 3579 3548
rect 111 3532 115 3536
rect 755 3535 759 3539
rect 1035 3535 1039 3539
rect 1823 3532 1827 3536
rect 1895 3531 1899 3535
rect 1983 3531 1987 3535
rect 2071 3531 2075 3535
rect 2159 3531 2163 3535
rect 2247 3531 2251 3535
rect 2335 3531 2339 3535
rect 2423 3531 2427 3535
rect 2511 3531 2515 3535
rect 2599 3531 2603 3535
rect 2687 3531 2691 3535
rect 2775 3531 2779 3535
rect 2863 3531 2867 3535
rect 2951 3531 2955 3535
rect 3039 3531 3043 3535
rect 3127 3531 3131 3535
rect 3215 3531 3219 3535
rect 3303 3531 3307 3535
rect 255 3519 259 3523
rect 407 3519 411 3523
rect 551 3519 555 3523
rect 695 3519 699 3523
rect 831 3519 835 3523
rect 959 3519 963 3523
rect 1087 3519 1091 3523
rect 1207 3519 1211 3523
rect 1319 3519 1323 3523
rect 1431 3519 1435 3523
rect 1551 3519 1555 3523
rect 1903 3519 1907 3523
rect 2631 3519 2632 3523
rect 2632 3519 2635 3523
rect 283 3507 284 3511
rect 284 3507 287 3511
rect 891 3507 895 3511
rect 1035 3507 1039 3511
rect 455 3495 459 3499
rect 755 3495 759 3499
rect 979 3495 983 3499
rect 1007 3495 1011 3499
rect 1247 3495 1248 3499
rect 1248 3495 1251 3499
rect 2083 3499 2087 3503
rect 2143 3499 2147 3503
rect 2351 3499 2355 3503
rect 2459 3499 2463 3503
rect 2571 3499 2575 3503
rect 2703 3499 2707 3503
rect 2891 3499 2895 3503
rect 3275 3499 3279 3503
rect 183 3485 187 3489
rect 351 3485 355 3489
rect 519 3485 523 3489
rect 679 3485 683 3489
rect 831 3485 835 3489
rect 967 3485 971 3489
rect 1095 3485 1099 3489
rect 1215 3485 1219 3489
rect 1335 3485 1339 3489
rect 1455 3485 1459 3489
rect 1575 3485 1579 3489
rect 1911 3489 1915 3493
rect 2015 3489 2019 3493
rect 2135 3489 2139 3493
rect 2263 3489 2267 3493
rect 2391 3489 2395 3493
rect 2527 3489 2531 3493
rect 2663 3489 2667 3493
rect 2799 3489 2803 3493
rect 2943 3489 2947 3493
rect 3087 3489 3091 3493
rect 111 3472 115 3476
rect 455 3467 459 3471
rect 891 3471 895 3475
rect 1823 3472 1827 3476
rect 1863 3476 1867 3480
rect 3575 3476 3579 3480
rect 1903 3471 1907 3475
rect 2083 3471 2087 3475
rect 2351 3471 2355 3475
rect 2459 3471 2463 3475
rect 2631 3471 2635 3475
rect 2891 3471 2895 3475
rect 111 3455 115 3459
rect 271 3455 275 3459
rect 175 3445 179 3449
rect 343 3445 347 3449
rect 511 3445 515 3449
rect 671 3445 675 3449
rect 823 3445 827 3449
rect 959 3445 963 3449
rect 979 3439 983 3443
rect 1087 3445 1091 3449
rect 1207 3445 1211 3449
rect 1327 3445 1331 3449
rect 1447 3445 1451 3449
rect 1335 3439 1339 3443
rect 1823 3455 1827 3459
rect 1863 3459 1867 3463
rect 2391 3459 2395 3463
rect 2799 3459 2803 3463
rect 3575 3459 3579 3463
rect 1567 3445 1571 3449
rect 1903 3449 1907 3453
rect 2007 3449 2011 3453
rect 2127 3449 2131 3453
rect 2255 3449 2259 3453
rect 2383 3449 2387 3453
rect 2519 3449 2523 3453
rect 2655 3449 2659 3453
rect 2791 3449 2795 3453
rect 2935 3449 2939 3453
rect 3079 3449 3083 3453
rect 135 3423 139 3427
rect 255 3423 259 3427
rect 415 3423 419 3427
rect 583 3423 587 3427
rect 759 3423 763 3427
rect 935 3423 939 3427
rect 1111 3423 1115 3427
rect 1295 3423 1299 3427
rect 1479 3423 1483 3427
rect 111 3413 115 3417
rect 679 3415 683 3419
rect 1007 3415 1011 3419
rect 1911 3419 1915 3423
rect 2071 3419 2075 3423
rect 2223 3419 2227 3423
rect 2367 3419 2371 3423
rect 2503 3419 2507 3423
rect 2631 3419 2635 3423
rect 2759 3419 2763 3423
rect 2887 3419 2891 3423
rect 3023 3419 3027 3423
rect 1823 3413 1827 3417
rect 1863 3409 1867 3413
rect 2143 3411 2147 3415
rect 2703 3411 2707 3415
rect 3575 3409 3579 3413
rect 111 3396 115 3400
rect 219 3399 223 3403
rect 1003 3399 1007 3403
rect 1587 3399 1591 3403
rect 1823 3396 1827 3400
rect 1863 3392 1867 3396
rect 2215 3395 2219 3399
rect 2291 3395 2295 3399
rect 2843 3395 2847 3399
rect 3091 3395 3095 3399
rect 3575 3392 3579 3396
rect 143 3383 147 3387
rect 263 3383 267 3387
rect 423 3383 427 3387
rect 591 3383 595 3387
rect 767 3383 771 3387
rect 943 3383 947 3387
rect 1119 3383 1123 3387
rect 1303 3383 1307 3387
rect 1487 3383 1491 3387
rect 1919 3379 1923 3383
rect 2079 3379 2083 3383
rect 2231 3379 2235 3383
rect 2375 3379 2379 3383
rect 2511 3379 2515 3383
rect 2639 3379 2643 3383
rect 2767 3379 2771 3383
rect 2895 3379 2899 3383
rect 3031 3379 3035 3383
rect 271 3371 275 3375
rect 219 3363 223 3367
rect 1003 3371 1007 3375
rect 1135 3371 1139 3375
rect 1335 3371 1336 3375
rect 1336 3371 1339 3375
rect 1951 3367 1952 3371
rect 1952 3367 1955 3371
rect 2291 3367 2295 3371
rect 2391 3367 2395 3371
rect 2603 3367 2607 3371
rect 2799 3367 2800 3371
rect 2800 3367 2803 3371
rect 2843 3367 2847 3371
rect 679 3359 683 3363
rect 951 3351 955 3355
rect 1587 3351 1588 3355
rect 1588 3351 1591 3355
rect 1991 3351 1995 3355
rect 2071 3351 2075 3355
rect 2215 3351 2219 3355
rect 2711 3351 2715 3355
rect 2987 3351 2991 3355
rect 3087 3351 3088 3355
rect 3088 3351 3091 3355
rect 207 3341 211 3345
rect 367 3341 371 3345
rect 535 3341 539 3345
rect 695 3341 699 3345
rect 855 3341 859 3345
rect 999 3341 1003 3345
rect 1143 3341 1147 3345
rect 1279 3341 1283 3345
rect 1415 3341 1419 3345
rect 1559 3341 1563 3345
rect 1895 3341 1899 3345
rect 2047 3341 2051 3345
rect 2207 3341 2211 3345
rect 2367 3341 2371 3345
rect 2535 3341 2539 3345
rect 2703 3341 2707 3345
rect 2879 3341 2883 3345
rect 3055 3341 3059 3345
rect 1951 3335 1955 3339
rect 111 3328 115 3332
rect 1823 3328 1827 3332
rect 1135 3323 1139 3327
rect 1863 3328 1867 3332
rect 1991 3323 1995 3327
rect 3575 3328 3579 3332
rect 2603 3323 2607 3327
rect 2987 3323 2991 3327
rect 111 3311 115 3315
rect 619 3311 623 3315
rect 1379 3311 1383 3315
rect 1823 3311 1827 3315
rect 1863 3311 1867 3315
rect 2495 3311 2499 3315
rect 2855 3311 2859 3315
rect 3575 3311 3579 3315
rect 199 3301 203 3305
rect 359 3301 363 3305
rect 527 3301 531 3305
rect 687 3301 691 3305
rect 847 3301 851 3305
rect 991 3301 995 3305
rect 1135 3301 1139 3305
rect 1271 3301 1275 3305
rect 1407 3301 1411 3305
rect 1551 3301 1555 3305
rect 1887 3301 1891 3305
rect 2039 3301 2043 3305
rect 2199 3301 2203 3305
rect 2359 3301 2363 3305
rect 2527 3301 2531 3305
rect 2695 3301 2699 3305
rect 2871 3301 2875 3305
rect 3047 3301 3051 3305
rect 255 3275 259 3279
rect 375 3275 379 3279
rect 511 3275 515 3279
rect 663 3275 667 3279
rect 823 3275 827 3279
rect 991 3275 995 3279
rect 1167 3275 1171 3279
rect 1343 3275 1347 3279
rect 1519 3275 1523 3279
rect 1887 3275 1891 3279
rect 2063 3275 2067 3279
rect 2263 3275 2267 3279
rect 2455 3275 2459 3279
rect 2639 3275 2643 3279
rect 2815 3275 2819 3279
rect 2983 3275 2987 3279
rect 3151 3275 3155 3279
rect 3319 3275 3323 3279
rect 3479 3275 3483 3279
rect 111 3265 115 3269
rect 739 3267 743 3271
rect 951 3267 955 3271
rect 1823 3265 1827 3269
rect 1863 3265 1867 3269
rect 2071 3263 2075 3267
rect 2711 3267 2715 3271
rect 3575 3265 3579 3269
rect 111 3248 115 3252
rect 1059 3251 1063 3255
rect 1587 3251 1591 3255
rect 1823 3248 1827 3252
rect 1863 3248 1867 3252
rect 2331 3251 2335 3255
rect 2339 3251 2343 3255
rect 3063 3251 3067 3255
rect 3071 3251 3075 3255
rect 3547 3251 3551 3255
rect 3575 3248 3579 3252
rect 263 3235 267 3239
rect 383 3235 387 3239
rect 519 3235 523 3239
rect 671 3235 675 3239
rect 831 3235 835 3239
rect 999 3235 1003 3239
rect 1175 3235 1179 3239
rect 1351 3235 1355 3239
rect 1527 3235 1531 3239
rect 1895 3235 1899 3239
rect 2071 3235 2075 3239
rect 2271 3235 2275 3239
rect 2463 3235 2467 3239
rect 2647 3235 2651 3239
rect 2823 3235 2827 3239
rect 2991 3235 2995 3239
rect 3159 3235 3163 3239
rect 3327 3235 3331 3239
rect 3487 3235 3491 3239
rect 295 3223 296 3227
rect 296 3223 299 3227
rect 1059 3223 1063 3227
rect 1207 3223 1208 3227
rect 1208 3223 1211 3227
rect 1379 3223 1380 3227
rect 1380 3223 1383 3227
rect 1955 3223 1959 3227
rect 2339 3223 2343 3227
rect 2495 3223 2496 3227
rect 2496 3223 2499 3227
rect 2679 3223 2680 3227
rect 2680 3223 2683 3227
rect 2855 3223 2856 3227
rect 2856 3223 2859 3227
rect 3063 3223 3067 3227
rect 463 3207 464 3211
rect 464 3207 467 3211
rect 1587 3207 1591 3211
rect 1963 3211 1967 3215
rect 2147 3211 2151 3215
rect 2331 3211 2332 3215
rect 2332 3211 2335 3215
rect 2763 3211 2767 3215
rect 2979 3211 2983 3215
rect 3071 3211 3072 3215
rect 3072 3211 3075 3215
rect 3411 3211 3415 3215
rect 3547 3211 3551 3215
rect 431 3197 435 3201
rect 551 3197 555 3201
rect 671 3197 675 3201
rect 799 3197 803 3201
rect 935 3197 939 3201
rect 1035 3199 1039 3203
rect 1079 3197 1083 3201
rect 1231 3197 1235 3201
rect 1383 3197 1387 3201
rect 1535 3197 1539 3201
rect 1895 3201 1899 3205
rect 2087 3201 2091 3205
rect 2303 3201 2307 3205
rect 2511 3201 2515 3205
rect 2703 3201 2707 3205
rect 2879 3201 2883 3205
rect 3039 3201 3043 3205
rect 3199 3201 3203 3205
rect 3351 3201 3355 3205
rect 3487 3201 3491 3205
rect 111 3184 115 3188
rect 1823 3184 1827 3188
rect 1863 3188 1867 3192
rect 1955 3187 1959 3191
rect 1207 3179 1211 3183
rect 1963 3183 1967 3187
rect 2679 3183 2683 3187
rect 2979 3183 2983 3187
rect 3575 3188 3579 3192
rect 111 3167 115 3171
rect 423 3157 427 3161
rect 543 3157 547 3161
rect 663 3157 667 3161
rect 503 3151 507 3155
rect 1823 3167 1827 3171
rect 1863 3171 1867 3175
rect 3575 3171 3579 3175
rect 791 3157 795 3161
rect 927 3157 931 3161
rect 1071 3157 1075 3161
rect 1223 3157 1227 3161
rect 1375 3157 1379 3161
rect 1527 3157 1531 3161
rect 1887 3161 1891 3165
rect 2079 3161 2083 3165
rect 2295 3161 2299 3165
rect 2503 3161 2507 3165
rect 2695 3161 2699 3165
rect 2871 3161 2875 3165
rect 3031 3161 3035 3165
rect 3191 3161 3195 3165
rect 3343 3161 3347 3165
rect 3479 3161 3483 3165
rect 1415 3151 1419 3155
rect 2543 3155 2547 3159
rect 2911 3155 2915 3159
rect 3519 3155 3523 3159
rect 463 3131 467 3135
rect 551 3131 555 3135
rect 639 3131 643 3135
rect 735 3131 739 3135
rect 847 3131 851 3135
rect 967 3131 971 3135
rect 1095 3131 1099 3135
rect 1231 3131 1235 3135
rect 1375 3131 1379 3135
rect 1519 3131 1523 3135
rect 1887 3135 1891 3139
rect 2079 3135 2083 3139
rect 2295 3135 2299 3139
rect 2503 3135 2507 3139
rect 2695 3135 2699 3139
rect 2871 3135 2875 3139
rect 3039 3135 3043 3139
rect 3191 3135 3195 3139
rect 3343 3135 3347 3139
rect 3479 3135 3483 3139
rect 111 3121 115 3125
rect 915 3123 919 3127
rect 1035 3123 1039 3127
rect 1823 3121 1827 3125
rect 1863 3125 1867 3129
rect 2147 3127 2151 3131
rect 2763 3127 2767 3131
rect 3411 3127 3415 3131
rect 3575 3125 3579 3129
rect 111 3104 115 3108
rect 1163 3107 1167 3111
rect 1587 3107 1591 3111
rect 1823 3104 1827 3108
rect 1863 3108 1867 3112
rect 2287 3111 2291 3115
rect 2363 3111 2367 3115
rect 3555 3111 3559 3115
rect 3575 3108 3579 3112
rect 471 3091 475 3095
rect 559 3091 563 3095
rect 647 3091 651 3095
rect 743 3091 747 3095
rect 855 3091 859 3095
rect 975 3091 979 3095
rect 1103 3091 1107 3095
rect 1239 3091 1243 3095
rect 1383 3091 1387 3095
rect 1527 3091 1531 3095
rect 1895 3095 1899 3099
rect 2087 3095 2091 3099
rect 2303 3095 2307 3099
rect 2511 3095 2515 3099
rect 2703 3095 2707 3099
rect 2879 3095 2883 3099
rect 3047 3095 3051 3099
rect 3199 3095 3203 3099
rect 3351 3095 3355 3099
rect 3487 3095 3491 3099
rect 503 3079 504 3083
rect 504 3079 507 3083
rect 1163 3079 1167 3083
rect 1415 3079 1416 3083
rect 1416 3079 1419 3083
rect 2363 3083 2367 3087
rect 2543 3083 2544 3087
rect 2544 3083 2547 3087
rect 2911 3083 2912 3087
rect 2912 3083 2915 3087
rect 3519 3083 3520 3087
rect 3520 3083 3523 3087
rect 223 3059 227 3063
rect 231 3059 235 3063
rect 1091 3059 1095 3063
rect 1539 3059 1543 3063
rect 1587 3059 1588 3063
rect 1588 3059 1591 3063
rect 1699 3059 1703 3063
rect 2287 3059 2288 3063
rect 2288 3059 2291 3063
rect 2783 3059 2784 3063
rect 2784 3059 2787 3063
rect 2931 3059 2935 3063
rect 151 3049 155 3053
rect 239 3049 243 3053
rect 327 3049 331 3053
rect 415 3049 419 3053
rect 503 3049 507 3053
rect 591 3049 595 3053
rect 679 3049 683 3053
rect 767 3049 771 3053
rect 855 3049 859 3053
rect 943 3049 947 3053
rect 1031 3049 1035 3053
rect 1119 3049 1123 3053
rect 1207 3049 1211 3053
rect 1295 3049 1299 3053
rect 1383 3049 1387 3053
rect 1471 3049 1475 3053
rect 1559 3049 1563 3053
rect 1647 3049 1651 3053
rect 1735 3049 1739 3053
rect 2255 3049 2259 3053
rect 2423 3049 2427 3053
rect 2591 3049 2595 3053
rect 2751 3049 2755 3053
rect 2919 3049 2923 3053
rect 3087 3049 3091 3053
rect 111 3036 115 3040
rect 231 3031 235 3035
rect 1091 3035 1095 3039
rect 1539 3031 1543 3035
rect 1823 3036 1827 3040
rect 1863 3036 1867 3040
rect 3575 3036 3579 3040
rect 3035 3031 3039 3035
rect 111 3019 115 3023
rect 1543 3019 1547 3023
rect 1823 3019 1827 3023
rect 1863 3019 1867 3023
rect 2499 3019 2503 3023
rect 3575 3019 3579 3023
rect 143 3009 147 3013
rect 231 3009 235 3013
rect 319 3009 323 3013
rect 407 3009 411 3013
rect 495 3009 499 3013
rect 583 3009 587 3013
rect 671 3009 675 3013
rect 759 3009 763 3013
rect 847 3009 851 3013
rect 935 3009 939 3013
rect 1023 3009 1027 3013
rect 1111 3009 1115 3013
rect 1199 3009 1203 3013
rect 1287 3009 1291 3013
rect 1375 3009 1379 3013
rect 1463 3009 1467 3013
rect 1551 3009 1555 3013
rect 1639 3009 1643 3013
rect 1727 3009 1731 3013
rect 2247 3009 2251 3013
rect 2415 3009 2419 3013
rect 2583 3009 2587 3013
rect 2743 3009 2747 3013
rect 2911 3009 2915 3013
rect 3079 3009 3083 3013
rect 1407 2979 1411 2983
rect 1519 2979 1523 2983
rect 1631 2979 1635 2983
rect 1727 2979 1731 2983
rect 2239 2983 2243 2987
rect 2463 2983 2467 2987
rect 2671 2983 2675 2987
rect 2863 2983 2867 2987
rect 3031 2983 3035 2987
rect 3191 2983 3195 2987
rect 3343 2983 3347 2987
rect 3479 2983 3483 2987
rect 111 2969 115 2973
rect 1699 2971 1703 2975
rect 1823 2969 1827 2973
rect 1863 2973 1867 2977
rect 2931 2975 2935 2979
rect 3575 2973 3579 2977
rect 111 2952 115 2956
rect 1479 2955 1483 2959
rect 1823 2952 1827 2956
rect 1863 2956 1867 2960
rect 2307 2959 2311 2963
rect 2351 2959 2355 2963
rect 2959 2959 2963 2963
rect 3099 2959 3103 2963
rect 3259 2959 3263 2963
rect 3547 2959 3551 2963
rect 3575 2956 3579 2960
rect 1499 2947 1503 2951
rect 1415 2939 1419 2943
rect 1527 2939 1531 2943
rect 1639 2939 1643 2943
rect 1735 2939 1739 2943
rect 2247 2943 2251 2947
rect 2471 2943 2475 2947
rect 2679 2943 2683 2947
rect 2871 2943 2875 2947
rect 3039 2943 3043 2947
rect 3199 2943 3203 2947
rect 3351 2943 3355 2947
rect 3487 2943 3491 2947
rect 1479 2927 1483 2931
rect 1535 2923 1539 2927
rect 1543 2927 1547 2931
rect 1763 2927 1764 2931
rect 1764 2927 1767 2931
rect 2351 2931 2355 2935
rect 2499 2931 2500 2935
rect 2500 2931 2503 2935
rect 2711 2931 2712 2935
rect 2712 2931 2715 2935
rect 3099 2931 3103 2935
rect 3259 2931 3263 2935
rect 3395 2931 3399 2935
rect 3555 2931 3559 2935
rect 1499 2915 1500 2919
rect 1500 2915 1503 2919
rect 1711 2915 1715 2919
rect 1359 2905 1363 2909
rect 1471 2905 1475 2909
rect 1583 2905 1587 2909
rect 1703 2905 1707 2909
rect 2307 2903 2311 2907
rect 2395 2903 2399 2907
rect 2751 2903 2755 2907
rect 3547 2903 3551 2907
rect 111 2892 115 2896
rect 1763 2891 1767 2895
rect 1823 2892 1827 2896
rect 2239 2893 2243 2897
rect 2463 2893 2467 2897
rect 2671 2893 2675 2897
rect 2855 2893 2859 2897
rect 3023 2893 3027 2897
rect 3183 2893 3187 2897
rect 3335 2893 3339 2897
rect 3487 2893 3491 2897
rect 1863 2880 1867 2884
rect 111 2875 115 2879
rect 1539 2875 1543 2879
rect 2395 2879 2399 2883
rect 1823 2875 1827 2879
rect 3395 2879 3399 2883
rect 3575 2880 3579 2884
rect 1351 2865 1355 2869
rect 1463 2865 1467 2869
rect 1575 2865 1579 2869
rect 1695 2865 1699 2869
rect 1419 2859 1423 2863
rect 1863 2863 1867 2867
rect 2547 2863 2551 2867
rect 3575 2863 3579 2867
rect 2231 2853 2235 2857
rect 2455 2853 2459 2857
rect 2663 2853 2667 2857
rect 2847 2853 2851 2857
rect 3015 2853 3019 2857
rect 3175 2853 3179 2857
rect 3327 2853 3331 2857
rect 3479 2853 3483 2857
rect 3519 2847 3523 2851
rect 135 2839 139 2843
rect 223 2839 227 2843
rect 311 2839 315 2843
rect 399 2839 403 2843
rect 487 2839 491 2843
rect 599 2839 603 2843
rect 727 2839 731 2843
rect 863 2839 867 2843
rect 999 2839 1003 2843
rect 1135 2839 1139 2843
rect 1263 2839 1267 2843
rect 1383 2839 1387 2843
rect 1503 2839 1507 2843
rect 1623 2839 1627 2843
rect 1727 2839 1731 2843
rect 111 2829 115 2833
rect 931 2831 935 2835
rect 1711 2831 1715 2835
rect 1823 2829 1827 2833
rect 1895 2827 1899 2831
rect 1983 2827 1987 2831
rect 2071 2827 2075 2831
rect 2159 2827 2163 2831
rect 2247 2827 2251 2831
rect 2335 2827 2339 2831
rect 2423 2827 2427 2831
rect 2511 2827 2515 2831
rect 2599 2827 2603 2831
rect 2687 2827 2691 2831
rect 2791 2827 2795 2831
rect 2903 2827 2907 2831
rect 3031 2827 3035 2831
rect 3175 2827 3179 2831
rect 3327 2827 3331 2831
rect 3479 2827 3483 2831
rect 111 2812 115 2816
rect 203 2815 207 2819
rect 379 2815 383 2819
rect 467 2815 471 2819
rect 559 2815 563 2819
rect 667 2815 671 2819
rect 1067 2815 1071 2819
rect 1331 2815 1335 2819
rect 1579 2815 1583 2819
rect 1691 2815 1695 2819
rect 1863 2817 1867 2821
rect 2499 2819 2503 2823
rect 3099 2819 3103 2823
rect 3575 2817 3579 2821
rect 1823 2812 1827 2816
rect 143 2799 147 2803
rect 231 2799 235 2803
rect 319 2799 323 2803
rect 407 2799 411 2803
rect 495 2799 499 2803
rect 607 2799 611 2803
rect 735 2799 739 2803
rect 871 2799 875 2803
rect 931 2795 935 2799
rect 1007 2799 1011 2803
rect 1143 2799 1147 2803
rect 1271 2799 1275 2803
rect 1391 2799 1395 2803
rect 1511 2799 1515 2803
rect 1631 2799 1635 2803
rect 1691 2795 1695 2799
rect 1735 2799 1739 2803
rect 1863 2800 1867 2804
rect 2491 2803 2495 2807
rect 3099 2803 3103 2807
rect 3243 2803 3247 2807
rect 3547 2803 3551 2807
rect 3575 2800 3579 2804
rect 203 2787 207 2791
rect 379 2787 383 2791
rect 467 2787 471 2791
rect 559 2787 563 2791
rect 667 2787 671 2791
rect 1331 2787 1335 2791
rect 1419 2787 1420 2791
rect 1420 2787 1423 2791
rect 1579 2787 1583 2791
rect 1795 2787 1799 2791
rect 1903 2787 1907 2791
rect 1991 2787 1995 2791
rect 2079 2787 2083 2791
rect 2167 2787 2171 2791
rect 2255 2787 2259 2791
rect 2343 2787 2347 2791
rect 2431 2787 2435 2791
rect 2519 2787 2523 2791
rect 2607 2787 2611 2791
rect 2695 2787 2699 2791
rect 2799 2787 2803 2791
rect 2911 2787 2915 2791
rect 3039 2787 3043 2791
rect 3183 2787 3187 2791
rect 3335 2787 3339 2791
rect 3487 2787 3491 2791
rect 571 2775 575 2779
rect 1191 2775 1195 2779
rect 191 2765 195 2769
rect 295 2765 299 2769
rect 415 2765 419 2769
rect 551 2765 555 2769
rect 687 2765 691 2769
rect 823 2765 827 2769
rect 959 2765 963 2769
rect 1067 2767 1071 2771
rect 2491 2775 2495 2779
rect 2547 2775 2548 2779
rect 2548 2775 2551 2779
rect 1087 2765 1091 2769
rect 1207 2765 1211 2769
rect 1319 2765 1323 2769
rect 1431 2765 1435 2769
rect 1535 2765 1539 2769
rect 1647 2765 1651 2769
rect 1735 2765 1739 2769
rect 3243 2775 3247 2779
rect 3519 2775 3520 2779
rect 3520 2775 3523 2779
rect 111 2752 115 2756
rect 1191 2751 1195 2755
rect 1795 2751 1799 2755
rect 1823 2752 1827 2756
rect 2023 2751 2027 2755
rect 2499 2751 2503 2755
rect 2707 2751 2711 2755
rect 3099 2751 3103 2755
rect 3199 2751 3203 2755
rect 3547 2751 3551 2755
rect 2047 2741 2051 2745
rect 2167 2741 2171 2745
rect 2295 2741 2299 2745
rect 2447 2741 2451 2745
rect 2623 2741 2627 2745
rect 2823 2741 2827 2745
rect 3039 2741 3043 2745
rect 3271 2741 3275 2745
rect 3487 2741 3491 2745
rect 111 2735 115 2739
rect 415 2735 419 2739
rect 1823 2735 1827 2739
rect 183 2725 187 2729
rect 287 2725 291 2729
rect 407 2725 411 2729
rect 543 2725 547 2729
rect 679 2725 683 2729
rect 815 2725 819 2729
rect 951 2725 955 2729
rect 1079 2725 1083 2729
rect 1199 2725 1203 2729
rect 1311 2725 1315 2729
rect 1423 2725 1427 2729
rect 1527 2725 1531 2729
rect 1639 2725 1643 2729
rect 1727 2725 1731 2729
rect 1863 2728 1867 2732
rect 2707 2723 2711 2727
rect 3575 2728 3579 2732
rect 1863 2711 1867 2715
rect 2371 2711 2375 2715
rect 2559 2711 2563 2715
rect 3575 2711 3579 2715
rect 2039 2701 2043 2705
rect 2159 2701 2163 2705
rect 2287 2701 2291 2705
rect 2439 2701 2443 2705
rect 2615 2701 2619 2705
rect 2815 2701 2819 2705
rect 3031 2701 3035 2705
rect 3263 2701 3267 2705
rect 3479 2701 3483 2705
rect 167 2695 171 2699
rect 279 2695 283 2699
rect 391 2695 395 2699
rect 503 2695 507 2699
rect 615 2695 619 2699
rect 3519 2695 3523 2699
rect 111 2685 115 2689
rect 571 2687 575 2691
rect 1823 2685 1827 2689
rect 1943 2679 1947 2683
rect 2055 2679 2059 2683
rect 2167 2679 2171 2683
rect 2287 2679 2291 2683
rect 2407 2679 2411 2683
rect 2519 2679 2523 2683
rect 2631 2679 2635 2683
rect 2735 2679 2739 2683
rect 2847 2679 2851 2683
rect 2959 2679 2963 2683
rect 3071 2679 3075 2683
rect 111 2668 115 2672
rect 235 2671 239 2675
rect 347 2671 351 2675
rect 571 2671 575 2675
rect 1823 2668 1827 2672
rect 1863 2669 1867 2673
rect 2023 2671 2027 2675
rect 3199 2671 3203 2675
rect 3575 2669 3579 2673
rect 251 2663 255 2667
rect 175 2655 179 2659
rect 287 2655 291 2659
rect 399 2655 403 2659
rect 511 2655 515 2659
rect 623 2655 627 2659
rect 1863 2652 1867 2656
rect 2011 2655 2015 2659
rect 2123 2655 2127 2659
rect 2491 2655 2495 2659
rect 3575 2652 3579 2656
rect 235 2643 239 2647
rect 347 2643 351 2647
rect 415 2643 419 2647
rect 571 2643 575 2647
rect 655 2643 656 2647
rect 656 2643 659 2647
rect 1951 2639 1955 2643
rect 2063 2639 2067 2643
rect 2175 2639 2179 2643
rect 2295 2639 2299 2643
rect 2415 2639 2419 2643
rect 2527 2639 2531 2643
rect 2639 2639 2643 2643
rect 2743 2639 2747 2643
rect 2855 2639 2859 2643
rect 2967 2639 2971 2643
rect 3079 2639 3083 2643
rect 2011 2627 2015 2631
rect 2123 2627 2127 2631
rect 2239 2627 2243 2631
rect 2371 2627 2375 2631
rect 2559 2627 2560 2631
rect 2560 2627 2563 2631
rect 251 2615 252 2619
rect 252 2615 255 2619
rect 759 2615 763 2619
rect 907 2615 911 2619
rect 967 2615 971 2619
rect 1247 2615 1248 2619
rect 1248 2615 1251 2619
rect 1959 2611 1963 2615
rect 2491 2611 2492 2615
rect 2492 2611 2495 2615
rect 2959 2611 2963 2615
rect 3519 2611 3520 2615
rect 3520 2611 3523 2615
rect 223 2605 227 2609
rect 351 2605 355 2609
rect 495 2605 499 2609
rect 663 2605 667 2609
rect 839 2605 843 2609
rect 1023 2605 1027 2609
rect 1215 2605 1219 2609
rect 1407 2605 1411 2609
rect 1607 2605 1611 2609
rect 1895 2601 1899 2605
rect 2071 2601 2075 2605
rect 2263 2601 2267 2605
rect 2463 2601 2467 2605
rect 2663 2601 2667 2605
rect 2871 2601 2875 2605
rect 3079 2601 3083 2605
rect 3295 2601 3299 2605
rect 3487 2601 3491 2605
rect 111 2592 115 2596
rect 655 2587 659 2591
rect 759 2587 763 2591
rect 907 2587 911 2591
rect 1823 2592 1827 2596
rect 1863 2588 1867 2592
rect 2239 2583 2243 2587
rect 3575 2588 3579 2592
rect 2959 2583 2963 2587
rect 111 2575 115 2579
rect 495 2575 499 2579
rect 1763 2575 1767 2579
rect 1823 2575 1827 2579
rect 1863 2571 1867 2575
rect 2531 2571 2535 2575
rect 2783 2571 2787 2575
rect 3575 2571 3579 2575
rect 215 2565 219 2569
rect 343 2565 347 2569
rect 487 2565 491 2569
rect 655 2565 659 2569
rect 831 2565 835 2569
rect 1015 2565 1019 2569
rect 1207 2565 1211 2569
rect 1399 2565 1403 2569
rect 1599 2565 1603 2569
rect 1887 2561 1891 2565
rect 2063 2561 2067 2565
rect 2255 2561 2259 2565
rect 2455 2561 2459 2565
rect 2655 2561 2659 2565
rect 2863 2561 2867 2565
rect 3071 2561 3075 2565
rect 3287 2561 3291 2565
rect 3479 2561 3483 2565
rect 3519 2555 3523 2559
rect 271 2543 275 2547
rect 471 2543 475 2547
rect 671 2543 675 2547
rect 855 2543 859 2547
rect 1023 2543 1027 2547
rect 1175 2543 1179 2547
rect 1319 2543 1323 2547
rect 1455 2543 1459 2547
rect 1591 2543 1595 2547
rect 1727 2543 1731 2547
rect 111 2533 115 2537
rect 967 2535 971 2539
rect 1247 2535 1251 2539
rect 1887 2539 1891 2543
rect 2039 2539 2043 2543
rect 2215 2539 2219 2543
rect 2399 2539 2403 2543
rect 2575 2539 2579 2543
rect 2743 2539 2747 2543
rect 2903 2539 2907 2543
rect 3055 2539 3059 2543
rect 3199 2539 3203 2543
rect 3343 2539 3347 2543
rect 3479 2539 3483 2543
rect 1823 2533 1827 2537
rect 1863 2529 1867 2533
rect 1959 2531 1963 2535
rect 3575 2529 3579 2533
rect 111 2516 115 2520
rect 215 2519 219 2523
rect 339 2519 343 2523
rect 1159 2519 1163 2523
rect 1387 2519 1391 2523
rect 1523 2519 1527 2523
rect 1659 2519 1663 2523
rect 1823 2516 1827 2520
rect 1863 2512 1867 2516
rect 1955 2515 1959 2519
rect 2107 2515 2111 2519
rect 2643 2515 2647 2519
rect 3147 2515 3151 2519
rect 3267 2515 3271 2519
rect 3547 2515 3551 2519
rect 3575 2512 3579 2516
rect 279 2503 283 2507
rect 479 2503 483 2507
rect 679 2503 683 2507
rect 863 2503 867 2507
rect 1031 2503 1035 2507
rect 1183 2503 1187 2507
rect 1327 2503 1331 2507
rect 1463 2503 1467 2507
rect 1599 2503 1603 2507
rect 1735 2503 1739 2507
rect 1895 2499 1899 2503
rect 2047 2499 2051 2503
rect 2223 2499 2227 2503
rect 2407 2499 2411 2503
rect 2583 2499 2587 2503
rect 2751 2499 2755 2503
rect 2911 2499 2915 2503
rect 3063 2499 3067 2503
rect 3207 2499 3211 2503
rect 3351 2499 3355 2503
rect 3487 2499 3491 2503
rect 339 2491 343 2495
rect 495 2491 499 2495
rect 1063 2491 1064 2495
rect 1064 2491 1067 2495
rect 1159 2491 1163 2495
rect 1523 2491 1527 2495
rect 1659 2491 1663 2495
rect 1763 2491 1764 2495
rect 1764 2491 1767 2495
rect 1387 2483 1391 2487
rect 1955 2487 1959 2491
rect 2107 2487 2111 2491
rect 2271 2487 2275 2491
rect 2531 2487 2535 2491
rect 2783 2487 2784 2491
rect 2784 2487 2787 2491
rect 3267 2487 3271 2491
rect 3519 2487 3520 2491
rect 3520 2487 3523 2491
rect 215 2475 216 2479
rect 216 2475 219 2479
rect 303 2475 307 2479
rect 1075 2475 1079 2479
rect 1159 2475 1160 2479
rect 1160 2475 1163 2479
rect 2539 2475 2543 2479
rect 2643 2475 2647 2479
rect 2875 2475 2879 2479
rect 3051 2475 3055 2479
rect 3147 2475 3148 2479
rect 3148 2475 3151 2479
rect 3311 2475 3315 2479
rect 3547 2475 3551 2479
rect 183 2465 187 2469
rect 319 2465 323 2469
rect 463 2465 467 2469
rect 607 2465 611 2469
rect 743 2465 747 2469
rect 879 2465 883 2469
rect 1007 2465 1011 2469
rect 1127 2465 1131 2469
rect 1239 2465 1243 2469
rect 1343 2465 1347 2469
rect 1447 2465 1451 2469
rect 1551 2465 1555 2469
rect 1647 2465 1651 2469
rect 1735 2465 1739 2469
rect 1895 2465 1899 2469
rect 1991 2465 1995 2469
rect 2127 2465 2131 2469
rect 2279 2465 2283 2469
rect 2439 2465 2443 2469
rect 2599 2465 2603 2469
rect 2767 2465 2771 2469
rect 2943 2465 2947 2469
rect 3119 2465 3123 2469
rect 3295 2465 3299 2469
rect 3471 2465 3475 2469
rect 1063 2459 1067 2463
rect 111 2452 115 2456
rect 303 2451 307 2455
rect 1075 2447 1079 2451
rect 1823 2452 1827 2456
rect 1863 2452 1867 2456
rect 2271 2447 2275 2451
rect 2539 2447 2543 2451
rect 2875 2447 2879 2451
rect 3051 2447 3055 2451
rect 3575 2452 3579 2456
rect 111 2435 115 2439
rect 387 2435 391 2439
rect 1823 2435 1827 2439
rect 1863 2435 1867 2439
rect 2391 2435 2395 2439
rect 2695 2435 2699 2439
rect 3575 2435 3579 2439
rect 175 2425 179 2429
rect 311 2425 315 2429
rect 455 2425 459 2429
rect 599 2425 603 2429
rect 735 2425 739 2429
rect 871 2425 875 2429
rect 999 2425 1003 2429
rect 1119 2425 1123 2429
rect 1231 2425 1235 2429
rect 1335 2425 1339 2429
rect 1439 2425 1443 2429
rect 1543 2425 1547 2429
rect 1639 2425 1643 2429
rect 1727 2425 1731 2429
rect 1887 2425 1891 2429
rect 1983 2425 1987 2429
rect 2119 2425 2123 2429
rect 2271 2425 2275 2429
rect 2431 2425 2435 2429
rect 2591 2425 2595 2429
rect 2759 2425 2763 2429
rect 2935 2425 2939 2429
rect 3111 2425 3115 2429
rect 3287 2425 3291 2429
rect 3463 2425 3467 2429
rect 3511 2419 3512 2423
rect 3512 2419 3515 2423
rect 1159 2403 1163 2407
rect 151 2395 155 2399
rect 319 2395 323 2399
rect 479 2395 483 2399
rect 639 2395 643 2399
rect 783 2395 787 2399
rect 919 2395 923 2399
rect 1047 2395 1051 2399
rect 1175 2395 1179 2399
rect 1303 2395 1307 2399
rect 111 2385 115 2389
rect 1431 2395 1435 2399
rect 2351 2395 2355 2399
rect 2503 2395 2507 2399
rect 2655 2395 2659 2399
rect 2807 2395 2811 2399
rect 2967 2395 2971 2399
rect 3135 2395 3139 2399
rect 3303 2395 3307 2399
rect 3471 2395 3475 2399
rect 1823 2385 1827 2389
rect 1863 2385 1867 2389
rect 3311 2383 3315 2387
rect 3575 2385 3579 2389
rect 111 2368 115 2372
rect 219 2371 223 2375
rect 227 2371 231 2375
rect 547 2371 551 2375
rect 707 2371 711 2375
rect 1167 2371 1171 2375
rect 2511 2375 2515 2379
rect 1823 2368 1827 2372
rect 1863 2368 1867 2372
rect 2587 2371 2591 2375
rect 3295 2371 3299 2375
rect 3539 2371 3543 2375
rect 3575 2368 3579 2372
rect 159 2355 163 2359
rect 327 2355 331 2359
rect 487 2355 491 2359
rect 647 2355 651 2359
rect 791 2355 795 2359
rect 927 2355 931 2359
rect 1055 2355 1059 2359
rect 1183 2355 1187 2359
rect 1311 2355 1315 2359
rect 1439 2355 1443 2359
rect 2359 2355 2363 2359
rect 2511 2355 2515 2359
rect 2663 2355 2667 2359
rect 2815 2355 2819 2359
rect 2975 2355 2979 2359
rect 3143 2355 3147 2359
rect 3311 2355 3315 2359
rect 3479 2355 3483 2359
rect 227 2343 231 2347
rect 387 2343 391 2347
rect 547 2343 551 2347
rect 707 2343 711 2347
rect 1027 2343 1031 2347
rect 1167 2343 1171 2347
rect 2391 2343 2392 2347
rect 2392 2343 2395 2347
rect 2539 2343 2540 2347
rect 2540 2343 2543 2347
rect 2695 2343 2696 2347
rect 2696 2343 2699 2347
rect 3371 2343 3375 2347
rect 3511 2343 3512 2347
rect 3512 2343 3515 2347
rect 2959 2335 2963 2339
rect 219 2327 223 2331
rect 439 2327 440 2331
rect 440 2327 443 2331
rect 1103 2327 1107 2331
rect 1219 2327 1223 2331
rect 2419 2327 2423 2331
rect 2523 2327 2527 2331
rect 2587 2327 2588 2331
rect 2588 2327 2591 2331
rect 3151 2327 3155 2331
rect 3295 2327 3299 2331
rect 3539 2327 3543 2331
rect 143 2317 147 2321
rect 263 2317 267 2321
rect 407 2317 411 2321
rect 543 2317 547 2321
rect 679 2317 683 2321
rect 807 2317 811 2321
rect 927 2317 931 2321
rect 1039 2317 1043 2321
rect 1159 2317 1163 2321
rect 1279 2317 1283 2321
rect 2351 2317 2355 2321
rect 2447 2317 2451 2321
rect 2559 2317 2563 2321
rect 2703 2317 2707 2321
rect 2879 2317 2883 2321
rect 3079 2317 3083 2321
rect 3287 2317 3291 2321
rect 3487 2317 3491 2321
rect 111 2304 115 2308
rect 1103 2303 1107 2307
rect 1219 2303 1223 2307
rect 1823 2304 1827 2308
rect 1863 2304 1867 2308
rect 1227 2299 1231 2303
rect 2419 2299 2423 2303
rect 2523 2299 2527 2303
rect 3575 2304 3579 2308
rect 2959 2299 2963 2303
rect 3151 2299 3155 2303
rect 111 2287 115 2291
rect 387 2287 391 2291
rect 1823 2287 1827 2291
rect 1863 2287 1867 2291
rect 2947 2287 2951 2291
rect 3575 2287 3579 2291
rect 135 2277 139 2281
rect 255 2277 259 2281
rect 399 2277 403 2281
rect 535 2277 539 2281
rect 671 2277 675 2281
rect 799 2277 803 2281
rect 919 2277 923 2281
rect 1031 2277 1035 2281
rect 1151 2277 1155 2281
rect 1271 2277 1275 2281
rect 2343 2277 2347 2281
rect 2439 2277 2443 2281
rect 2551 2277 2555 2281
rect 2695 2277 2699 2281
rect 2871 2277 2875 2281
rect 3071 2277 3075 2281
rect 3279 2277 3283 2281
rect 3479 2277 3483 2281
rect 2375 2271 2379 2275
rect 3519 2271 3523 2275
rect 135 2255 139 2259
rect 231 2255 235 2259
rect 351 2255 355 2259
rect 471 2255 475 2259
rect 591 2255 595 2259
rect 711 2255 715 2259
rect 823 2255 827 2259
rect 935 2255 939 2259
rect 1055 2255 1059 2259
rect 1175 2255 1179 2259
rect 2335 2255 2339 2259
rect 2447 2255 2451 2259
rect 2583 2255 2587 2259
rect 2735 2255 2739 2259
rect 2911 2255 2915 2259
rect 3103 2255 3107 2259
rect 3303 2255 3307 2259
rect 3479 2255 3483 2259
rect 111 2245 115 2249
rect 439 2247 443 2251
rect 1823 2245 1827 2249
rect 1863 2245 1867 2249
rect 3371 2247 3375 2251
rect 3575 2245 3579 2249
rect 111 2228 115 2232
rect 203 2231 207 2235
rect 299 2231 303 2235
rect 539 2231 543 2235
rect 779 2231 783 2235
rect 1139 2231 1143 2235
rect 1147 2231 1151 2235
rect 1823 2228 1827 2232
rect 1863 2228 1867 2232
rect 2567 2231 2571 2235
rect 2575 2231 2579 2235
rect 2727 2231 2731 2235
rect 3015 2231 3019 2235
rect 3023 2231 3027 2235
rect 3547 2231 3551 2235
rect 3575 2228 3579 2232
rect 143 2215 147 2219
rect 239 2215 243 2219
rect 359 2215 363 2219
rect 479 2215 483 2219
rect 599 2215 603 2219
rect 719 2215 723 2219
rect 831 2215 835 2219
rect 943 2215 947 2219
rect 1063 2215 1067 2219
rect 203 2203 207 2207
rect 299 2203 303 2207
rect 387 2203 388 2207
rect 388 2203 391 2207
rect 539 2203 543 2207
rect 631 2203 632 2207
rect 632 2203 635 2207
rect 779 2203 783 2207
rect 1147 2211 1151 2215
rect 1183 2215 1187 2219
rect 2343 2215 2347 2219
rect 2455 2215 2459 2219
rect 2591 2215 2595 2219
rect 2743 2215 2747 2219
rect 2919 2215 2923 2219
rect 3023 2211 3027 2215
rect 3111 2215 3115 2219
rect 3311 2215 3315 2219
rect 3487 2215 3491 2219
rect 971 2203 972 2207
rect 972 2203 975 2207
rect 1139 2203 1143 2207
rect 2375 2203 2376 2207
rect 2376 2203 2379 2207
rect 2567 2203 2571 2207
rect 2947 2203 2948 2207
rect 2948 2203 2951 2207
rect 3015 2203 3019 2207
rect 3343 2203 3344 2207
rect 3344 2203 3347 2207
rect 3519 2203 3520 2207
rect 3520 2203 3523 2207
rect 979 2195 983 2199
rect 427 2187 431 2191
rect 1231 2187 1235 2191
rect 2323 2191 2327 2195
rect 2411 2191 2415 2195
rect 2515 2191 2519 2195
rect 2575 2191 2579 2195
rect 2727 2191 2728 2195
rect 2728 2191 2731 2195
rect 2823 2191 2827 2195
rect 3547 2191 3551 2195
rect 143 2177 147 2181
rect 247 2177 251 2181
rect 383 2177 387 2181
rect 519 2177 523 2181
rect 655 2177 659 2181
rect 783 2177 787 2181
rect 911 2177 915 2181
rect 1031 2177 1035 2181
rect 1159 2177 1163 2181
rect 1287 2177 1291 2181
rect 2255 2181 2259 2185
rect 2343 2181 2347 2185
rect 2439 2181 2443 2185
rect 2551 2181 2555 2185
rect 2695 2181 2699 2185
rect 2871 2181 2875 2185
rect 3071 2181 3075 2185
rect 3287 2181 3291 2185
rect 3487 2181 3491 2185
rect 111 2164 115 2168
rect 631 2159 635 2163
rect 971 2163 975 2167
rect 1823 2164 1827 2168
rect 1863 2168 1867 2172
rect 979 2159 983 2163
rect 2323 2163 2327 2167
rect 1231 2159 1235 2163
rect 2411 2163 2415 2167
rect 2515 2163 2519 2167
rect 2823 2167 2827 2171
rect 3575 2168 3579 2172
rect 111 2147 115 2151
rect 1823 2147 1827 2151
rect 1863 2151 1867 2155
rect 2343 2151 2347 2155
rect 3199 2151 3203 2155
rect 3575 2151 3579 2155
rect 135 2137 139 2141
rect 239 2137 243 2141
rect 375 2137 379 2141
rect 511 2137 515 2141
rect 647 2137 651 2141
rect 775 2137 779 2141
rect 903 2137 907 2141
rect 1023 2137 1027 2141
rect 1151 2137 1155 2141
rect 1279 2137 1283 2141
rect 2247 2141 2251 2145
rect 2335 2141 2339 2145
rect 2431 2141 2435 2145
rect 2543 2141 2547 2145
rect 2687 2141 2691 2145
rect 2863 2141 2867 2145
rect 3063 2141 3067 2145
rect 3279 2141 3283 2145
rect 3479 2141 3483 2145
rect 271 2131 275 2135
rect 3519 2135 3523 2139
rect 135 2107 139 2111
rect 231 2107 235 2111
rect 359 2107 363 2111
rect 479 2107 483 2111
rect 599 2107 603 2111
rect 719 2107 723 2111
rect 831 2107 835 2111
rect 943 2107 947 2111
rect 1055 2107 1059 2111
rect 1175 2107 1179 2111
rect 2151 2111 2155 2115
rect 2239 2111 2243 2115
rect 2327 2111 2331 2115
rect 2415 2111 2419 2115
rect 2503 2111 2507 2115
rect 2615 2111 2619 2115
rect 2751 2111 2755 2115
rect 2919 2111 2923 2115
rect 3103 2111 3107 2115
rect 3303 2111 3307 2115
rect 3479 2111 3483 2115
rect 111 2097 115 2101
rect 427 2099 431 2103
rect 1823 2097 1827 2101
rect 1863 2101 1867 2105
rect 2483 2103 2487 2107
rect 3575 2101 3579 2105
rect 111 2080 115 2084
rect 203 2083 207 2087
rect 427 2083 431 2087
rect 547 2083 551 2087
rect 1823 2080 1827 2084
rect 1863 2084 1867 2088
rect 2307 2087 2311 2091
rect 3095 2087 3099 2091
rect 3555 2087 3559 2091
rect 3575 2084 3579 2088
rect 143 2067 147 2071
rect 239 2067 243 2071
rect 367 2067 371 2071
rect 487 2067 491 2071
rect 607 2067 611 2071
rect 727 2067 731 2071
rect 839 2067 843 2071
rect 951 2067 955 2071
rect 1063 2067 1067 2071
rect 1183 2067 1187 2071
rect 2159 2071 2163 2075
rect 2247 2071 2251 2075
rect 2335 2071 2339 2075
rect 2423 2071 2427 2075
rect 2511 2071 2515 2075
rect 2623 2071 2627 2075
rect 2759 2071 2763 2075
rect 2927 2071 2931 2075
rect 3111 2071 3115 2075
rect 3311 2071 3315 2075
rect 3487 2071 3491 2075
rect 203 2055 207 2059
rect 271 2055 272 2059
rect 272 2055 275 2059
rect 427 2055 431 2059
rect 547 2055 551 2059
rect 635 2055 636 2059
rect 636 2055 639 2059
rect 759 2055 760 2059
rect 760 2055 763 2059
rect 2191 2059 2192 2063
rect 2192 2059 2195 2063
rect 2343 2059 2347 2063
rect 2663 2059 2667 2063
rect 3095 2059 3099 2063
rect 3519 2059 3520 2063
rect 3520 2059 3523 2063
rect 2071 2043 2075 2047
rect 2307 2043 2311 2047
rect 2367 2043 2371 2047
rect 2831 2043 2835 2047
rect 2991 2043 2995 2047
rect 3175 2043 3179 2047
rect 3419 2043 3423 2047
rect 387 2031 391 2035
rect 399 2031 403 2035
rect 727 2027 731 2031
rect 755 2031 759 2035
rect 983 2031 987 2035
rect 1083 2031 1087 2035
rect 1191 2031 1195 2035
rect 1311 2031 1315 2035
rect 1999 2033 2003 2037
rect 2127 2033 2131 2037
rect 2255 2033 2259 2037
rect 2399 2033 2403 2037
rect 2551 2033 2555 2037
rect 2711 2033 2715 2037
rect 2879 2033 2883 2037
rect 3063 2033 3067 2037
rect 3247 2033 3251 2037
rect 3439 2033 3443 2037
rect 167 2021 171 2025
rect 311 2021 315 2025
rect 447 2021 451 2025
rect 575 2021 579 2025
rect 695 2021 699 2025
rect 807 2021 811 2025
rect 911 2021 915 2025
rect 1015 2021 1019 2025
rect 1119 2021 1123 2025
rect 1223 2021 1227 2025
rect 1327 2021 1331 2025
rect 1863 2020 1867 2024
rect 2367 2019 2371 2023
rect 2479 2015 2483 2019
rect 2831 2019 2835 2023
rect 2991 2019 2995 2023
rect 3175 2019 3179 2023
rect 3575 2020 3579 2024
rect 3343 2015 3347 2019
rect 111 2008 115 2012
rect 399 2007 403 2011
rect 635 2007 639 2011
rect 755 2007 759 2011
rect 1823 2008 1827 2012
rect 763 2003 767 2007
rect 983 2003 987 2007
rect 1083 2003 1087 2007
rect 1191 2003 1195 2007
rect 1863 2003 1867 2007
rect 2195 2003 2199 2007
rect 3151 2003 3155 2007
rect 3575 2003 3579 2007
rect 111 1991 115 1995
rect 1015 1991 1019 1995
rect 1823 1991 1827 1995
rect 1991 1993 1995 1997
rect 2119 1993 2123 1997
rect 2247 1993 2251 1997
rect 2391 1993 2395 1997
rect 2543 1993 2547 1997
rect 2703 1993 2707 1997
rect 2871 1993 2875 1997
rect 3055 1993 3059 1997
rect 3239 1993 3243 1997
rect 3431 1993 3435 1997
rect 159 1981 163 1985
rect 303 1981 307 1985
rect 439 1981 443 1985
rect 567 1981 571 1985
rect 687 1981 691 1985
rect 799 1981 803 1985
rect 903 1981 907 1985
rect 1007 1981 1011 1985
rect 1111 1981 1115 1985
rect 1215 1981 1219 1985
rect 1319 1981 1323 1985
rect 207 1975 208 1979
rect 208 1975 211 1979
rect 159 1959 163 1963
rect 295 1959 299 1963
rect 439 1959 443 1963
rect 583 1959 587 1963
rect 719 1959 723 1963
rect 855 1959 859 1963
rect 991 1959 995 1963
rect 1119 1959 1123 1963
rect 1239 1959 1243 1963
rect 1359 1959 1363 1963
rect 1479 1959 1483 1963
rect 1599 1959 1603 1963
rect 1903 1963 1907 1967
rect 2159 1963 2163 1967
rect 2399 1963 2403 1967
rect 2615 1963 2619 1967
rect 2815 1963 2819 1967
rect 2999 1963 3003 1967
rect 3167 1963 3171 1967
rect 3335 1963 3339 1967
rect 3479 1963 3483 1967
rect 111 1949 115 1953
rect 387 1951 391 1955
rect 727 1947 731 1951
rect 1311 1951 1315 1955
rect 1823 1949 1827 1953
rect 1863 1953 1867 1957
rect 3259 1955 3263 1959
rect 3575 1953 3579 1957
rect 111 1932 115 1936
rect 507 1935 511 1939
rect 787 1935 791 1939
rect 923 1935 927 1939
rect 1307 1935 1311 1939
rect 1427 1935 1431 1939
rect 1547 1935 1551 1939
rect 1823 1932 1827 1936
rect 1863 1936 1867 1940
rect 2011 1939 2015 1943
rect 3547 1939 3551 1943
rect 3575 1936 3579 1940
rect 167 1919 171 1923
rect 303 1919 307 1923
rect 447 1919 451 1923
rect 591 1919 595 1923
rect 727 1919 731 1923
rect 787 1915 791 1919
rect 863 1919 867 1923
rect 999 1919 1003 1923
rect 1127 1919 1131 1923
rect 1247 1919 1251 1923
rect 1367 1919 1371 1923
rect 1487 1919 1491 1923
rect 1607 1919 1611 1923
rect 1911 1923 1915 1927
rect 2167 1923 2171 1927
rect 2407 1923 2411 1927
rect 2623 1923 2627 1927
rect 2823 1923 2827 1927
rect 3007 1923 3011 1927
rect 3175 1923 3179 1927
rect 3343 1923 3347 1927
rect 3487 1923 3491 1927
rect 207 1907 211 1911
rect 507 1907 511 1911
rect 779 1907 783 1911
rect 923 1907 927 1911
rect 1015 1907 1019 1911
rect 1427 1907 1431 1911
rect 1547 1907 1551 1911
rect 1667 1907 1671 1911
rect 1943 1911 1944 1915
rect 1944 1911 1947 1915
rect 2195 1911 2196 1915
rect 2196 1911 2199 1915
rect 2655 1911 2656 1915
rect 2656 1911 2659 1915
rect 3555 1911 3559 1915
rect 1307 1899 1311 1903
rect 2011 1899 2012 1903
rect 2012 1899 2015 1903
rect 2111 1899 2115 1903
rect 2951 1899 2952 1903
rect 2952 1899 2955 1903
rect 3427 1899 3431 1903
rect 3547 1899 3551 1903
rect 751 1887 752 1891
rect 752 1887 755 1891
rect 1031 1887 1035 1891
rect 1895 1889 1899 1893
rect 1983 1889 1987 1893
rect 2071 1889 2075 1893
rect 2167 1889 2171 1893
rect 2295 1889 2299 1893
rect 2447 1889 2451 1893
rect 2607 1889 2611 1893
rect 2767 1889 2771 1893
rect 2919 1889 2923 1893
rect 3071 1889 3075 1893
rect 3215 1889 3219 1893
rect 3359 1889 3363 1893
rect 3487 1889 3491 1893
rect 223 1877 227 1881
rect 479 1877 483 1881
rect 719 1877 723 1881
rect 935 1877 939 1881
rect 1127 1877 1131 1881
rect 1295 1877 1299 1881
rect 1455 1877 1459 1881
rect 1607 1877 1611 1881
rect 1735 1877 1739 1881
rect 1863 1876 1867 1880
rect 2403 1871 2407 1875
rect 3419 1875 3423 1879
rect 3575 1876 3579 1880
rect 3427 1871 3431 1875
rect 111 1864 115 1868
rect 779 1863 783 1867
rect 1667 1863 1671 1867
rect 1823 1864 1827 1868
rect 1863 1859 1867 1863
rect 2675 1859 2679 1863
rect 3575 1859 3579 1863
rect 111 1847 115 1851
rect 1823 1847 1827 1851
rect 1887 1849 1891 1853
rect 1975 1849 1979 1853
rect 2063 1849 2067 1853
rect 2159 1849 2163 1853
rect 2287 1849 2291 1853
rect 2439 1849 2443 1853
rect 2599 1849 2603 1853
rect 2759 1849 2763 1853
rect 2911 1849 2915 1853
rect 3063 1849 3067 1853
rect 3207 1849 3211 1853
rect 3351 1849 3355 1853
rect 3479 1849 3483 1853
rect 215 1837 219 1841
rect 471 1837 475 1841
rect 711 1837 715 1841
rect 927 1837 931 1841
rect 1119 1837 1123 1841
rect 1287 1837 1291 1841
rect 1447 1837 1451 1841
rect 1599 1837 1603 1841
rect 1727 1837 1731 1841
rect 283 1831 287 1835
rect 1767 1831 1771 1835
rect 1999 1823 2003 1827
rect 2223 1823 2227 1827
rect 2439 1823 2443 1827
rect 2639 1823 2643 1827
rect 2831 1823 2835 1827
rect 3015 1823 3019 1827
rect 3199 1823 3203 1827
rect 3391 1823 3395 1827
rect 247 1815 251 1819
rect 415 1815 419 1819
rect 591 1815 595 1819
rect 759 1815 763 1819
rect 927 1815 931 1819
rect 1079 1815 1083 1819
rect 1223 1815 1227 1819
rect 1359 1815 1363 1819
rect 1487 1815 1491 1819
rect 1615 1815 1619 1819
rect 1727 1815 1731 1819
rect 1863 1813 1867 1817
rect 2111 1815 2115 1819
rect 2719 1815 2723 1819
rect 3575 1813 3579 1817
rect 111 1805 115 1809
rect 751 1807 755 1811
rect 1031 1807 1035 1811
rect 1823 1805 1827 1809
rect 1863 1796 1867 1800
rect 2819 1799 2823 1803
rect 2899 1799 2903 1803
rect 3083 1799 3087 1803
rect 3459 1799 3463 1803
rect 111 1788 115 1792
rect 575 1791 579 1795
rect 659 1791 663 1795
rect 827 1791 831 1795
rect 1147 1791 1151 1795
rect 1291 1791 1295 1795
rect 1555 1791 1559 1795
rect 3575 1796 3579 1800
rect 1683 1791 1687 1795
rect 1823 1788 1827 1792
rect 1563 1783 1567 1787
rect 2007 1783 2011 1787
rect 2231 1783 2235 1787
rect 2447 1783 2451 1787
rect 2647 1783 2651 1787
rect 2839 1783 2843 1787
rect 3023 1783 3027 1787
rect 3207 1783 3211 1787
rect 3399 1783 3403 1787
rect 255 1775 259 1779
rect 423 1775 427 1779
rect 599 1775 603 1779
rect 767 1775 771 1779
rect 935 1775 939 1779
rect 1087 1775 1091 1779
rect 1231 1775 1235 1779
rect 1367 1775 1371 1779
rect 1495 1775 1499 1779
rect 1623 1775 1627 1779
rect 1735 1775 1739 1779
rect 2263 1771 2264 1775
rect 2264 1771 2267 1775
rect 2479 1771 2480 1775
rect 2480 1771 2483 1775
rect 2899 1771 2903 1775
rect 3083 1771 3087 1775
rect 3259 1771 3263 1775
rect 283 1763 284 1767
rect 284 1763 287 1767
rect 575 1763 579 1767
rect 827 1763 831 1767
rect 979 1763 983 1767
rect 1147 1763 1151 1767
rect 1291 1763 1295 1767
rect 1435 1763 1439 1767
rect 1555 1763 1559 1767
rect 1683 1763 1687 1767
rect 1767 1763 1768 1767
rect 1768 1763 1771 1767
rect 539 1755 543 1759
rect 659 1747 663 1751
rect 839 1747 843 1751
rect 1111 1747 1115 1751
rect 1563 1751 1567 1755
rect 2035 1755 2039 1759
rect 2187 1755 2191 1759
rect 2819 1755 2820 1759
rect 2820 1755 2823 1759
rect 3231 1755 3232 1759
rect 3232 1755 3235 1759
rect 3459 1755 3463 1759
rect 1943 1745 1947 1749
rect 2087 1745 2091 1749
rect 2247 1745 2251 1749
rect 2415 1745 2419 1749
rect 2599 1745 2603 1749
rect 2791 1745 2795 1749
rect 2991 1745 2995 1749
rect 3199 1745 3203 1749
rect 3415 1745 3419 1749
rect 327 1737 331 1741
rect 471 1737 475 1741
rect 615 1737 619 1741
rect 767 1737 771 1741
rect 919 1737 923 1741
rect 1071 1737 1075 1741
rect 1223 1737 1227 1741
rect 1375 1737 1379 1741
rect 1527 1737 1531 1741
rect 1687 1737 1691 1741
rect 1863 1732 1867 1736
rect 111 1724 115 1728
rect 539 1719 543 1723
rect 979 1723 983 1727
rect 1435 1723 1439 1727
rect 1823 1724 1827 1728
rect 2035 1727 2039 1731
rect 2187 1727 2191 1731
rect 3259 1731 3263 1735
rect 3575 1732 3579 1736
rect 1863 1715 1867 1719
rect 111 1707 115 1711
rect 615 1707 619 1711
rect 1687 1707 1691 1711
rect 1823 1707 1827 1711
rect 1935 1705 1939 1709
rect 2079 1705 2083 1709
rect 2239 1705 2243 1709
rect 2407 1705 2411 1709
rect 319 1697 323 1701
rect 463 1697 467 1701
rect 607 1697 611 1701
rect 759 1697 763 1701
rect 911 1697 915 1701
rect 1063 1697 1067 1701
rect 1215 1697 1219 1701
rect 1367 1697 1371 1701
rect 1519 1697 1523 1701
rect 1679 1697 1683 1701
rect 2311 1699 2315 1703
rect 3083 1715 3087 1719
rect 3575 1715 3579 1719
rect 2591 1705 2595 1709
rect 2783 1705 2787 1709
rect 2983 1705 2987 1709
rect 3191 1705 3195 1709
rect 3407 1705 3411 1709
rect 3467 1699 3471 1703
rect 1911 1679 1915 1683
rect 2031 1679 2035 1683
rect 2151 1679 2155 1683
rect 2271 1679 2275 1683
rect 2399 1679 2403 1683
rect 2543 1679 2547 1683
rect 2695 1679 2699 1683
rect 2863 1679 2867 1683
rect 3047 1679 3051 1683
rect 3239 1679 3243 1683
rect 3431 1679 3435 1683
rect 311 1671 315 1675
rect 447 1671 451 1675
rect 591 1671 595 1675
rect 735 1671 739 1675
rect 887 1671 891 1675
rect 1039 1671 1043 1675
rect 1191 1671 1195 1675
rect 1343 1671 1347 1675
rect 1495 1671 1499 1675
rect 1647 1671 1651 1675
rect 1863 1669 1867 1673
rect 3231 1671 3235 1675
rect 3575 1669 3579 1673
rect 111 1661 115 1665
rect 839 1663 843 1667
rect 1111 1663 1115 1667
rect 1823 1661 1827 1665
rect 1863 1652 1867 1656
rect 2467 1655 2471 1659
rect 111 1644 115 1648
rect 255 1647 259 1651
rect 379 1647 383 1651
rect 515 1647 519 1651
rect 1143 1647 1147 1651
rect 1411 1647 1415 1651
rect 1563 1647 1567 1651
rect 2611 1655 2615 1659
rect 2763 1655 2767 1659
rect 2931 1655 2935 1659
rect 3499 1655 3503 1659
rect 3575 1652 3579 1656
rect 1823 1644 1827 1648
rect 2619 1647 2623 1651
rect 1919 1639 1923 1643
rect 2039 1639 2043 1643
rect 2159 1639 2163 1643
rect 2279 1639 2283 1643
rect 2407 1639 2411 1643
rect 2551 1639 2555 1643
rect 2703 1639 2707 1643
rect 2871 1639 2875 1643
rect 3055 1639 3059 1643
rect 3247 1639 3251 1643
rect 3439 1639 3443 1643
rect 319 1631 323 1635
rect 455 1631 459 1635
rect 599 1631 603 1635
rect 743 1631 747 1635
rect 895 1631 899 1635
rect 1047 1631 1051 1635
rect 1199 1631 1203 1635
rect 1351 1631 1355 1635
rect 1503 1631 1507 1635
rect 1655 1631 1659 1635
rect 1959 1627 1963 1631
rect 2311 1627 2312 1631
rect 2312 1627 2315 1631
rect 2611 1627 2615 1631
rect 2763 1627 2767 1631
rect 2931 1627 2935 1631
rect 3083 1627 3084 1631
rect 3084 1627 3087 1631
rect 3271 1627 3275 1631
rect 3467 1627 3468 1631
rect 3468 1627 3471 1631
rect 379 1619 383 1623
rect 515 1619 519 1623
rect 615 1619 619 1623
rect 751 1619 755 1623
rect 1143 1619 1147 1623
rect 1207 1619 1211 1623
rect 1411 1619 1415 1623
rect 1563 1619 1567 1623
rect 1687 1619 1688 1623
rect 1688 1619 1691 1623
rect 1975 1607 1979 1611
rect 2083 1607 2087 1611
rect 2463 1607 2464 1611
rect 2464 1607 2467 1611
rect 2619 1611 2623 1615
rect 3311 1607 3312 1611
rect 3312 1607 3315 1611
rect 3499 1607 3500 1611
rect 3500 1607 3503 1611
rect 255 1599 256 1603
rect 256 1599 259 1603
rect 651 1599 652 1603
rect 652 1599 655 1603
rect 955 1599 959 1603
rect 1175 1599 1179 1603
rect 1895 1597 1899 1601
rect 2015 1597 2019 1601
rect 2151 1597 2155 1601
rect 2287 1597 2291 1601
rect 2431 1597 2435 1601
rect 2583 1597 2587 1601
rect 2743 1597 2747 1601
rect 2911 1597 2915 1601
rect 3095 1597 3099 1601
rect 3279 1597 3283 1601
rect 3471 1597 3475 1601
rect 223 1589 227 1593
rect 351 1589 355 1593
rect 487 1589 491 1593
rect 623 1589 627 1593
rect 759 1589 763 1593
rect 903 1589 907 1593
rect 1055 1589 1059 1593
rect 1215 1589 1219 1593
rect 1375 1589 1379 1593
rect 1543 1589 1547 1593
rect 1863 1584 1867 1588
rect 1959 1583 1963 1587
rect 111 1576 115 1580
rect 751 1571 755 1575
rect 1175 1575 1179 1579
rect 1207 1571 1211 1575
rect 1823 1576 1827 1580
rect 1975 1579 1979 1583
rect 2083 1579 2087 1583
rect 3575 1584 3579 1588
rect 3271 1579 3275 1583
rect 1863 1567 1867 1571
rect 2223 1567 2227 1571
rect 3019 1567 3023 1571
rect 3575 1567 3579 1571
rect 111 1559 115 1563
rect 463 1559 467 1563
rect 1543 1559 1547 1563
rect 1823 1559 1827 1563
rect 1887 1557 1891 1561
rect 2007 1557 2011 1561
rect 2143 1557 2147 1561
rect 2279 1557 2283 1561
rect 2423 1557 2427 1561
rect 2575 1557 2579 1561
rect 2735 1557 2739 1561
rect 2903 1557 2907 1561
rect 3087 1557 3091 1561
rect 3271 1557 3275 1561
rect 3463 1557 3467 1561
rect 215 1549 219 1553
rect 343 1549 347 1553
rect 479 1549 483 1553
rect 615 1549 619 1553
rect 751 1549 755 1553
rect 895 1549 899 1553
rect 1047 1549 1051 1553
rect 1207 1549 1211 1553
rect 1367 1549 1371 1553
rect 1535 1549 1539 1553
rect 3515 1551 3516 1555
rect 3516 1551 3519 1555
rect 135 1523 139 1527
rect 271 1523 275 1527
rect 423 1523 427 1527
rect 583 1523 587 1527
rect 735 1523 739 1527
rect 887 1523 891 1527
rect 1039 1523 1043 1527
rect 1191 1523 1195 1527
rect 1343 1523 1347 1527
rect 1495 1523 1499 1527
rect 1887 1527 1891 1531
rect 2023 1527 2027 1531
rect 2183 1527 2187 1531
rect 2343 1527 2347 1531
rect 2503 1527 2507 1531
rect 2663 1527 2667 1531
rect 2823 1527 2827 1531
rect 2983 1527 2987 1531
rect 3151 1527 3155 1531
rect 3319 1527 3323 1531
rect 3479 1527 3483 1531
rect 111 1513 115 1517
rect 651 1515 655 1519
rect 955 1515 959 1519
rect 1823 1513 1827 1517
rect 1863 1517 1867 1521
rect 3079 1519 3083 1523
rect 3311 1519 3315 1523
rect 3575 1517 3579 1521
rect 111 1496 115 1500
rect 339 1499 343 1503
rect 651 1499 655 1503
rect 955 1499 959 1503
rect 1411 1499 1415 1503
rect 1419 1499 1423 1503
rect 1823 1496 1827 1500
rect 1863 1500 1867 1504
rect 2731 1503 2735 1507
rect 3547 1503 3551 1507
rect 3575 1500 3579 1504
rect 2567 1495 2571 1499
rect 199 1491 203 1495
rect 143 1483 147 1487
rect 279 1483 283 1487
rect 431 1483 435 1487
rect 591 1483 595 1487
rect 743 1483 747 1487
rect 895 1483 899 1487
rect 1047 1483 1051 1487
rect 1199 1483 1203 1487
rect 1351 1483 1355 1487
rect 1503 1483 1507 1487
rect 1895 1487 1899 1491
rect 2031 1487 2035 1491
rect 2191 1487 2195 1491
rect 2351 1487 2355 1491
rect 2511 1487 2515 1491
rect 2671 1487 2675 1491
rect 2831 1487 2835 1491
rect 2991 1487 2995 1491
rect 3159 1487 3163 1491
rect 3327 1487 3331 1491
rect 3487 1487 3491 1491
rect 339 1471 343 1475
rect 463 1471 464 1475
rect 464 1471 467 1475
rect 651 1471 655 1475
rect 955 1471 959 1475
rect 1079 1471 1080 1475
rect 1080 1471 1083 1475
rect 1543 1471 1547 1475
rect 2223 1475 2224 1479
rect 2224 1475 2227 1479
rect 2703 1475 2704 1479
rect 2704 1475 2707 1479
rect 2731 1475 2735 1479
rect 3351 1475 3355 1479
rect 3515 1475 3516 1479
rect 3516 1475 3519 1479
rect 1091 1459 1095 1463
rect 1419 1463 1423 1467
rect 199 1451 203 1455
rect 1211 1451 1215 1455
rect 1403 1451 1407 1455
rect 1411 1451 1412 1455
rect 1412 1451 1415 1455
rect 2223 1455 2227 1459
rect 2567 1455 2571 1459
rect 2719 1455 2720 1459
rect 2720 1455 2723 1459
rect 3547 1455 3551 1459
rect 143 1441 147 1445
rect 263 1441 267 1445
rect 399 1441 403 1445
rect 535 1441 539 1445
rect 623 1443 627 1447
rect 663 1441 667 1445
rect 791 1441 795 1445
rect 911 1441 915 1445
rect 1023 1441 1027 1445
rect 1143 1441 1147 1445
rect 1263 1441 1267 1445
rect 1383 1441 1387 1445
rect 1503 1441 1507 1445
rect 1631 1441 1635 1445
rect 1735 1441 1739 1445
rect 2183 1445 2187 1449
rect 2359 1445 2363 1449
rect 2527 1445 2531 1449
rect 2687 1445 2691 1449
rect 2847 1445 2851 1449
rect 3007 1445 3011 1449
rect 3175 1445 3179 1449
rect 3343 1445 3347 1449
rect 3487 1445 3491 1449
rect 1079 1435 1083 1439
rect 111 1428 115 1432
rect 1091 1423 1095 1427
rect 1211 1423 1215 1427
rect 1823 1428 1827 1432
rect 1863 1432 1867 1436
rect 2427 1427 2431 1431
rect 3575 1432 3579 1436
rect 111 1411 115 1415
rect 535 1411 539 1415
rect 135 1401 139 1405
rect 255 1401 259 1405
rect 391 1401 395 1405
rect 527 1401 531 1405
rect 655 1401 659 1405
rect 783 1401 787 1405
rect 903 1401 907 1405
rect 1015 1401 1019 1405
rect 1135 1401 1139 1405
rect 1255 1401 1259 1405
rect 1375 1401 1379 1405
rect 1403 1395 1407 1399
rect 1823 1411 1827 1415
rect 1863 1415 1867 1419
rect 2475 1415 2479 1419
rect 3259 1415 3263 1419
rect 3575 1415 3579 1419
rect 1495 1401 1499 1405
rect 1623 1401 1627 1405
rect 1727 1401 1731 1405
rect 2175 1405 2179 1409
rect 2351 1405 2355 1409
rect 2519 1405 2523 1409
rect 2679 1405 2683 1409
rect 2839 1405 2843 1409
rect 2999 1405 3003 1409
rect 3167 1405 3171 1409
rect 3335 1405 3339 1409
rect 3479 1405 3483 1409
rect 3519 1399 3523 1403
rect 135 1379 139 1383
rect 327 1379 331 1383
rect 551 1379 555 1383
rect 783 1379 787 1383
rect 1023 1379 1027 1383
rect 1263 1379 1267 1383
rect 1503 1379 1507 1383
rect 1727 1379 1731 1383
rect 111 1369 115 1373
rect 623 1371 627 1375
rect 2079 1375 2083 1379
rect 2263 1375 2267 1379
rect 2439 1375 2443 1379
rect 2615 1375 2619 1379
rect 2783 1375 2787 1379
rect 2935 1375 2939 1379
rect 3079 1375 3083 1379
rect 3223 1375 3227 1379
rect 3359 1375 3363 1379
rect 3479 1375 3483 1379
rect 1823 1369 1827 1373
rect 1863 1365 1867 1369
rect 2539 1367 2543 1371
rect 3351 1367 3355 1371
rect 3575 1365 3579 1369
rect 111 1352 115 1356
rect 395 1355 399 1359
rect 851 1355 855 1359
rect 1639 1355 1643 1359
rect 1823 1352 1827 1356
rect 199 1347 203 1351
rect 1863 1348 1867 1352
rect 2339 1351 2343 1355
rect 3547 1351 3551 1355
rect 3575 1348 3579 1352
rect 143 1339 147 1343
rect 335 1339 339 1343
rect 559 1339 563 1343
rect 791 1339 795 1343
rect 1031 1339 1035 1343
rect 1271 1339 1275 1343
rect 1511 1339 1515 1343
rect 1735 1339 1739 1343
rect 2087 1335 2091 1339
rect 2271 1335 2275 1339
rect 2447 1335 2451 1339
rect 2623 1335 2627 1339
rect 2791 1335 2795 1339
rect 2943 1335 2947 1339
rect 3087 1335 3091 1339
rect 3231 1335 3235 1339
rect 3367 1335 3371 1339
rect 3487 1335 3491 1339
rect 395 1327 399 1331
rect 535 1327 539 1331
rect 851 1327 855 1331
rect 1303 1327 1304 1331
rect 1304 1327 1307 1331
rect 2119 1323 2120 1327
rect 2120 1323 2123 1327
rect 2475 1323 2476 1327
rect 2476 1323 2479 1327
rect 2823 1323 2824 1327
rect 2824 1323 2827 1327
rect 3419 1323 3423 1327
rect 3519 1323 3520 1327
rect 3520 1323 3523 1327
rect 1459 1315 1463 1319
rect 199 1307 203 1311
rect 615 1307 619 1311
rect 1215 1307 1219 1311
rect 2295 1311 2299 1315
rect 2339 1311 2340 1315
rect 2340 1311 2343 1315
rect 2763 1311 2767 1315
rect 3115 1311 3119 1315
rect 3547 1311 3551 1315
rect 143 1297 147 1301
rect 327 1297 331 1301
rect 527 1297 531 1301
rect 719 1297 723 1301
rect 903 1297 907 1301
rect 1071 1297 1075 1301
rect 1231 1297 1235 1301
rect 1383 1297 1387 1301
rect 1535 1297 1539 1301
rect 1687 1297 1691 1301
rect 2087 1301 2091 1305
rect 2311 1301 2315 1305
rect 2519 1301 2523 1305
rect 2711 1301 2715 1305
rect 2887 1301 2891 1305
rect 3047 1301 3051 1305
rect 3199 1301 3203 1305
rect 3351 1301 3355 1305
rect 3487 1301 3491 1305
rect 111 1284 115 1288
rect 1215 1283 1219 1287
rect 1823 1284 1827 1288
rect 1863 1288 1867 1292
rect 2443 1283 2447 1287
rect 3575 1288 3579 1292
rect 3115 1283 3119 1287
rect 111 1267 115 1271
rect 211 1267 215 1271
rect 1823 1267 1827 1271
rect 1863 1271 1867 1275
rect 2959 1271 2963 1275
rect 3575 1271 3579 1275
rect 135 1257 139 1261
rect 319 1257 323 1261
rect 519 1257 523 1261
rect 711 1257 715 1261
rect 895 1257 899 1261
rect 1063 1257 1067 1261
rect 1223 1257 1227 1261
rect 1375 1257 1379 1261
rect 1527 1257 1531 1261
rect 1679 1257 1683 1261
rect 2079 1261 2083 1265
rect 2303 1261 2307 1265
rect 2511 1261 2515 1265
rect 2703 1261 2707 1265
rect 2879 1261 2883 1265
rect 3039 1261 3043 1265
rect 3191 1261 3195 1265
rect 3343 1261 3347 1265
rect 3479 1261 3483 1265
rect 2131 1255 2132 1259
rect 2132 1255 2135 1259
rect 2951 1255 2955 1259
rect 3519 1255 3523 1259
rect 2763 1247 2767 1251
rect 2959 1247 2963 1251
rect 135 1231 139 1235
rect 295 1231 299 1235
rect 479 1231 483 1235
rect 655 1231 659 1235
rect 815 1231 819 1235
rect 967 1231 971 1235
rect 1111 1231 1115 1235
rect 1247 1231 1251 1235
rect 1383 1231 1387 1235
rect 1527 1231 1531 1235
rect 1903 1235 1907 1239
rect 1991 1235 1995 1239
rect 2095 1235 2099 1239
rect 2215 1235 2219 1239
rect 2351 1235 2355 1239
rect 2487 1235 2491 1239
rect 2631 1235 2635 1239
rect 2775 1235 2779 1239
rect 2919 1235 2923 1239
rect 3063 1235 3067 1239
rect 3207 1235 3211 1239
rect 3351 1235 3355 1239
rect 3479 1235 3483 1239
rect 111 1221 115 1225
rect 615 1223 619 1227
rect 1459 1223 1463 1227
rect 1823 1221 1827 1225
rect 1863 1225 1867 1229
rect 2555 1227 2559 1231
rect 3139 1227 3143 1231
rect 3419 1227 3423 1231
rect 3575 1225 3579 1229
rect 111 1204 115 1208
rect 547 1207 551 1211
rect 723 1207 727 1211
rect 1823 1204 1827 1208
rect 1863 1208 1867 1212
rect 1971 1211 1975 1215
rect 1979 1211 1983 1215
rect 2087 1211 2091 1215
rect 2163 1211 2167 1215
rect 2283 1211 2287 1215
rect 2699 1211 2703 1215
rect 3547 1211 3551 1215
rect 3575 1208 3579 1212
rect 143 1191 147 1195
rect 303 1191 307 1195
rect 487 1191 491 1195
rect 663 1191 667 1195
rect 823 1191 827 1195
rect 975 1191 979 1195
rect 1119 1191 1123 1195
rect 1255 1191 1259 1195
rect 1391 1191 1395 1195
rect 1535 1191 1539 1195
rect 1911 1195 1915 1199
rect 1999 1195 2003 1199
rect 2103 1195 2107 1199
rect 2163 1191 2167 1195
rect 2223 1195 2227 1199
rect 2359 1195 2363 1199
rect 2495 1195 2499 1199
rect 2555 1191 2559 1195
rect 2639 1195 2643 1199
rect 2783 1195 2787 1199
rect 2927 1195 2931 1199
rect 3071 1195 3075 1199
rect 3215 1195 3219 1199
rect 3359 1195 3363 1199
rect 3487 1195 3491 1199
rect 211 1179 215 1183
rect 723 1179 727 1183
rect 1051 1179 1055 1183
rect 1979 1183 1983 1187
rect 2131 1183 2132 1187
rect 2132 1183 2135 1187
rect 2283 1183 2287 1187
rect 2815 1183 2816 1187
rect 2816 1183 2819 1187
rect 2951 1183 2955 1187
rect 3387 1183 3388 1187
rect 3388 1183 3391 1187
rect 3519 1183 3520 1187
rect 3520 1183 3523 1187
rect 235 1163 239 1167
rect 391 1163 395 1167
rect 547 1163 551 1167
rect 647 1163 648 1167
rect 648 1163 651 1167
rect 999 1163 1003 1167
rect 1871 1163 1875 1167
rect 1971 1167 1975 1171
rect 2087 1167 2091 1171
rect 2479 1167 2483 1171
rect 2699 1167 2703 1171
rect 3355 1163 3359 1167
rect 3547 1167 3551 1171
rect 167 1153 171 1157
rect 319 1153 323 1157
rect 471 1153 475 1157
rect 615 1153 619 1157
rect 759 1153 763 1157
rect 911 1153 915 1157
rect 1063 1153 1067 1157
rect 1231 1153 1235 1157
rect 1399 1153 1403 1157
rect 1575 1153 1579 1157
rect 1735 1153 1739 1157
rect 1895 1157 1899 1161
rect 2063 1157 2067 1161
rect 2255 1157 2259 1161
rect 2439 1157 2443 1161
rect 2615 1157 2619 1161
rect 2791 1157 2795 1161
rect 2967 1157 2971 1161
rect 3143 1157 3147 1161
rect 3327 1157 3331 1161
rect 3487 1157 3491 1161
rect 111 1140 115 1144
rect 235 1135 239 1139
rect 391 1135 395 1139
rect 1823 1140 1827 1144
rect 1863 1144 1867 1148
rect 1871 1139 1875 1143
rect 3387 1143 3391 1147
rect 3575 1144 3579 1148
rect 1539 1135 1543 1139
rect 111 1123 115 1127
rect 251 1123 255 1127
rect 1823 1123 1827 1127
rect 1863 1127 1867 1131
rect 2135 1127 2139 1131
rect 3143 1127 3147 1131
rect 3575 1127 3579 1131
rect 159 1113 163 1117
rect 311 1113 315 1117
rect 463 1113 467 1117
rect 607 1113 611 1117
rect 751 1113 755 1117
rect 903 1113 907 1117
rect 1055 1113 1059 1117
rect 1223 1113 1227 1117
rect 1391 1113 1395 1117
rect 1567 1113 1571 1117
rect 1727 1113 1731 1117
rect 1887 1117 1891 1121
rect 2055 1117 2059 1121
rect 2247 1117 2251 1121
rect 2431 1117 2435 1121
rect 2607 1117 2611 1121
rect 2783 1117 2787 1121
rect 2959 1117 2963 1121
rect 3135 1117 3139 1121
rect 3319 1117 3323 1121
rect 3479 1117 3483 1121
rect 1767 1107 1771 1111
rect 3519 1111 3523 1115
rect 215 1087 219 1091
rect 327 1087 331 1091
rect 439 1087 443 1091
rect 559 1087 563 1091
rect 679 1087 683 1091
rect 807 1087 811 1091
rect 943 1087 947 1091
rect 1087 1087 1091 1091
rect 1247 1087 1251 1091
rect 1407 1087 1411 1091
rect 1575 1087 1579 1091
rect 1727 1087 1731 1091
rect 111 1077 115 1081
rect 647 1079 651 1083
rect 1339 1079 1343 1083
rect 1935 1083 1939 1087
rect 2095 1083 2099 1087
rect 2247 1083 2251 1087
rect 2407 1083 2411 1087
rect 2567 1083 2571 1087
rect 2735 1083 2739 1087
rect 2911 1083 2915 1087
rect 3095 1083 3099 1087
rect 3287 1083 3291 1087
rect 3479 1083 3483 1087
rect 1823 1077 1827 1081
rect 1863 1073 1867 1077
rect 2011 1075 2015 1079
rect 2479 1075 2483 1079
rect 2643 1075 2647 1079
rect 3355 1075 3359 1079
rect 3575 1073 3579 1077
rect 111 1060 115 1064
rect 1567 1063 1571 1067
rect 1643 1063 1647 1067
rect 1823 1060 1827 1064
rect 1863 1056 1867 1060
rect 2003 1059 2007 1063
rect 2635 1059 2639 1063
rect 2979 1059 2983 1063
rect 3547 1059 3551 1063
rect 3575 1056 3579 1060
rect 223 1047 227 1051
rect 335 1047 339 1051
rect 447 1047 451 1051
rect 567 1047 571 1051
rect 687 1047 691 1051
rect 815 1047 819 1051
rect 951 1047 955 1051
rect 1095 1047 1099 1051
rect 1255 1047 1259 1051
rect 1415 1047 1419 1051
rect 1583 1047 1587 1051
rect 1735 1047 1739 1051
rect 1943 1043 1947 1047
rect 2103 1043 2107 1047
rect 2255 1043 2259 1047
rect 2415 1043 2419 1047
rect 2575 1043 2579 1047
rect 2743 1043 2747 1047
rect 2919 1043 2923 1047
rect 3103 1043 3107 1047
rect 3295 1043 3299 1047
rect 3487 1043 3491 1047
rect 251 1035 252 1039
rect 252 1035 255 1039
rect 715 1035 716 1039
rect 716 1035 719 1039
rect 859 1035 863 1039
rect 1643 1035 1647 1039
rect 1767 1035 1768 1039
rect 1768 1035 1771 1039
rect 2003 1031 2007 1035
rect 2135 1031 2136 1035
rect 2136 1031 2139 1035
rect 2379 1031 2383 1035
rect 2635 1031 2639 1035
rect 2979 1031 2983 1035
rect 3143 1031 3147 1035
rect 3519 1031 3520 1035
rect 3520 1031 3523 1035
rect 411 1015 415 1019
rect 503 1015 507 1019
rect 723 1015 727 1019
rect 823 1015 824 1019
rect 824 1015 827 1019
rect 1039 1015 1043 1019
rect 1203 1015 1207 1019
rect 1279 1015 1283 1019
rect 1567 1015 1568 1019
rect 1568 1015 1571 1019
rect 2011 1015 2015 1019
rect 2115 1015 2119 1019
rect 2643 1015 2647 1019
rect 3419 1015 3423 1019
rect 3547 1015 3551 1019
rect 343 1005 347 1009
rect 431 1005 435 1009
rect 535 1005 539 1009
rect 655 1005 659 1009
rect 791 1005 795 1009
rect 951 1005 955 1009
rect 1135 1005 1139 1009
rect 1327 1005 1331 1009
rect 1535 1005 1539 1009
rect 1735 1005 1739 1009
rect 1943 1005 1947 1009
rect 2071 1005 2075 1009
rect 2191 1005 2195 1009
rect 2311 1005 2315 1009
rect 2439 1005 2443 1009
rect 2575 1005 2579 1009
rect 2719 1005 2723 1009
rect 2871 1005 2875 1009
rect 3031 1005 3035 1009
rect 3191 1005 3195 1009
rect 3351 1005 3355 1009
rect 3487 1005 3491 1009
rect 111 992 115 996
rect 411 987 415 991
rect 503 987 507 991
rect 715 991 719 995
rect 723 987 727 991
rect 859 987 863 991
rect 1039 987 1043 991
rect 1203 987 1207 991
rect 1823 992 1827 996
rect 1863 992 1867 996
rect 3575 992 3579 996
rect 3419 987 3423 991
rect 111 975 115 979
rect 1735 975 1739 979
rect 1823 975 1827 979
rect 1863 975 1867 979
rect 1943 975 1947 979
rect 2379 975 2383 979
rect 2959 975 2963 979
rect 3575 975 3579 979
rect 335 965 339 969
rect 423 965 427 969
rect 527 965 531 969
rect 647 965 651 969
rect 783 965 787 969
rect 943 965 947 969
rect 1127 965 1131 969
rect 1319 965 1323 969
rect 1527 965 1531 969
rect 1727 965 1731 969
rect 1935 965 1939 969
rect 2063 965 2067 969
rect 2183 965 2187 969
rect 2303 965 2307 969
rect 2431 965 2435 969
rect 2567 965 2571 969
rect 2711 965 2715 969
rect 2863 965 2867 969
rect 3023 965 3027 969
rect 3183 965 3187 969
rect 3343 965 3347 969
rect 3479 965 3483 969
rect 403 959 407 963
rect 2535 951 2539 955
rect 2959 951 2963 955
rect 367 939 371 943
rect 463 939 467 943
rect 575 939 579 943
rect 703 939 707 943
rect 847 939 851 943
rect 1007 939 1011 943
rect 1175 939 1179 943
rect 1351 939 1355 943
rect 1527 939 1531 943
rect 1711 939 1715 943
rect 1887 939 1891 943
rect 2047 939 2051 943
rect 2199 939 2203 943
rect 2351 939 2355 943
rect 2495 939 2499 943
rect 2631 939 2635 943
rect 2759 939 2763 943
rect 2887 939 2891 943
rect 3023 939 3027 943
rect 111 929 115 933
rect 823 931 827 935
rect 1279 931 1283 935
rect 1823 929 1827 933
rect 1863 929 1867 933
rect 2115 931 2119 935
rect 3575 929 3579 933
rect 111 912 115 916
rect 563 915 567 919
rect 1167 915 1171 919
rect 1659 915 1663 919
rect 1667 915 1671 919
rect 1823 912 1827 916
rect 1863 912 1867 916
rect 2039 915 2043 919
rect 2267 915 2271 919
rect 2715 915 2719 919
rect 2855 915 2859 919
rect 3091 915 3095 919
rect 3575 912 3579 916
rect 375 899 379 903
rect 471 899 475 903
rect 583 899 587 903
rect 711 899 715 903
rect 855 899 859 903
rect 1015 899 1019 903
rect 1183 899 1187 903
rect 1359 899 1363 903
rect 1535 899 1539 903
rect 1719 899 1723 903
rect 1895 899 1899 903
rect 2055 899 2059 903
rect 2207 899 2211 903
rect 2359 899 2363 903
rect 2503 899 2507 903
rect 2639 899 2643 903
rect 2767 899 2771 903
rect 2895 899 2899 903
rect 3031 899 3035 903
rect 403 887 404 891
rect 404 887 407 891
rect 635 887 639 891
rect 1167 887 1171 891
rect 1391 887 1392 891
rect 1392 887 1395 891
rect 1735 887 1739 891
rect 1943 887 1947 891
rect 2267 887 2271 891
rect 2391 887 2392 891
rect 2392 887 2395 891
rect 2535 887 2536 891
rect 2536 887 2539 891
rect 2715 887 2719 891
rect 2855 887 2859 891
rect 411 871 415 875
rect 503 871 507 875
rect 563 871 564 875
rect 564 871 567 875
rect 719 871 723 875
rect 815 871 816 875
rect 816 871 819 875
rect 1027 871 1031 875
rect 1195 871 1199 875
rect 1223 871 1227 875
rect 1519 871 1523 875
rect 1659 871 1660 875
rect 1660 871 1663 875
rect 1967 875 1971 879
rect 2039 875 2043 879
rect 2207 871 2211 875
rect 2383 875 2387 879
rect 2879 875 2880 879
rect 2880 875 2883 879
rect 3091 875 3095 879
rect 3407 875 3411 879
rect 343 861 347 865
rect 431 861 435 865
rect 535 861 539 865
rect 647 861 651 865
rect 783 861 787 865
rect 927 861 931 865
rect 1087 861 1091 865
rect 1263 861 1267 865
rect 1447 861 1451 865
rect 1631 861 1635 865
rect 1895 865 1899 869
rect 2015 865 2019 869
rect 2167 865 2171 869
rect 2319 865 2323 869
rect 2487 865 2491 869
rect 2663 865 2667 869
rect 2847 865 2851 869
rect 3039 865 3043 869
rect 3239 865 3243 869
rect 3439 865 3443 869
rect 111 848 115 852
rect 411 843 415 847
rect 503 843 507 847
rect 635 843 639 847
rect 719 843 723 847
rect 1823 848 1827 852
rect 1863 852 1867 856
rect 1027 843 1031 847
rect 1195 843 1199 847
rect 1967 847 1971 851
rect 2383 851 2387 855
rect 1519 843 1523 847
rect 2391 847 2395 851
rect 3575 852 3579 856
rect 111 831 115 835
rect 431 831 435 835
rect 1823 831 1827 835
rect 1863 835 1867 839
rect 2663 835 2667 839
rect 335 821 339 825
rect 423 821 427 825
rect 527 821 531 825
rect 639 821 643 825
rect 775 821 779 825
rect 919 821 923 825
rect 1079 821 1083 825
rect 1255 821 1259 825
rect 1439 821 1443 825
rect 1623 821 1627 825
rect 1887 825 1891 829
rect 2007 825 2011 829
rect 2159 825 2163 829
rect 2311 825 2315 829
rect 2479 825 2483 829
rect 2655 825 2659 829
rect 2839 825 2843 829
rect 3031 825 3035 829
rect 1479 815 1483 819
rect 1927 819 1931 823
rect 2879 819 2883 823
rect 3515 835 3519 839
rect 3575 835 3579 839
rect 3231 825 3235 829
rect 3431 825 3435 829
rect 287 799 291 803
rect 407 799 411 803
rect 535 799 539 803
rect 679 799 683 803
rect 823 799 827 803
rect 975 799 979 803
rect 1127 799 1131 803
rect 1279 799 1283 803
rect 1439 799 1443 803
rect 1599 799 1603 803
rect 1887 803 1891 807
rect 1991 803 1995 807
rect 2135 803 2139 807
rect 2287 803 2291 807
rect 2455 803 2459 807
rect 2623 803 2627 807
rect 2799 803 2803 807
rect 2967 803 2971 807
rect 3143 803 3147 807
rect 3319 803 3323 807
rect 3479 803 3483 807
rect 111 789 115 793
rect 475 791 479 795
rect 815 791 819 795
rect 1223 791 1227 795
rect 1519 791 1523 795
rect 1823 789 1827 793
rect 1863 793 1867 797
rect 2207 795 2211 799
rect 3407 795 3411 799
rect 3575 793 3579 797
rect 111 772 115 776
rect 247 775 251 779
rect 1823 772 1827 776
rect 1863 776 1867 780
rect 1955 779 1959 783
rect 2203 779 2207 783
rect 2355 779 2359 783
rect 2867 779 2871 783
rect 3547 779 3551 783
rect 3575 776 3579 780
rect 295 759 299 763
rect 415 759 419 763
rect 475 755 479 759
rect 543 759 547 763
rect 687 759 691 763
rect 831 759 835 763
rect 983 759 987 763
rect 1135 759 1139 763
rect 1287 759 1291 763
rect 1447 759 1451 763
rect 1607 759 1611 763
rect 1895 763 1899 767
rect 1999 763 2003 767
rect 2143 763 2147 767
rect 2295 763 2299 767
rect 2463 763 2467 767
rect 2631 763 2635 767
rect 2807 763 2811 767
rect 2975 763 2979 767
rect 3151 763 3155 767
rect 3327 763 3331 767
rect 3487 763 3491 767
rect 431 747 435 751
rect 707 747 711 751
rect 1315 747 1316 751
rect 1316 747 1319 751
rect 1479 747 1480 751
rect 1480 747 1483 751
rect 1927 751 1928 755
rect 1928 751 1931 755
rect 2355 751 2359 755
rect 2507 751 2511 755
rect 2663 751 2664 755
rect 2664 751 2667 755
rect 3235 751 3239 755
rect 3515 751 3516 755
rect 3516 751 3519 755
rect 1163 739 1167 743
rect 2203 743 2207 747
rect 247 731 248 735
rect 248 731 251 735
rect 327 731 331 735
rect 739 731 743 735
rect 843 731 847 735
rect 1143 731 1147 735
rect 1871 731 1875 735
rect 1955 735 1959 739
rect 2095 735 2096 739
rect 2096 735 2099 739
rect 2731 735 2735 739
rect 2867 735 2871 739
rect 3059 735 3063 739
rect 3227 735 3231 739
rect 3547 735 3551 739
rect 215 721 219 725
rect 359 721 363 725
rect 503 721 507 725
rect 647 721 651 725
rect 791 721 795 725
rect 935 721 939 725
rect 1087 721 1091 725
rect 1247 721 1251 725
rect 1415 721 1419 725
rect 1583 721 1587 725
rect 1735 721 1739 725
rect 1895 725 1899 729
rect 2063 725 2067 729
rect 2255 725 2259 729
rect 2447 725 2451 729
rect 2639 725 2643 729
rect 2823 725 2827 729
rect 2999 725 3003 729
rect 3167 725 3171 729
rect 3335 725 3339 729
rect 3487 725 3491 729
rect 111 708 115 712
rect 327 707 331 711
rect 707 707 711 711
rect 739 703 743 707
rect 1823 708 1827 712
rect 1863 712 1867 716
rect 1871 707 1875 711
rect 2507 711 2511 715
rect 2731 707 2735 711
rect 3227 711 3231 715
rect 3575 712 3579 716
rect 3235 707 3239 711
rect 111 691 115 695
rect 503 691 507 695
rect 1163 691 1167 695
rect 1519 691 1523 695
rect 1823 691 1827 695
rect 1863 695 1867 699
rect 2707 695 2711 699
rect 3575 695 3579 699
rect 207 681 211 685
rect 351 681 355 685
rect 495 681 499 685
rect 639 681 643 685
rect 783 681 787 685
rect 927 681 931 685
rect 1079 681 1083 685
rect 1239 681 1243 685
rect 1407 681 1411 685
rect 1575 681 1579 685
rect 1727 681 1731 685
rect 1887 685 1891 689
rect 2055 685 2059 689
rect 2247 685 2251 689
rect 2439 685 2443 689
rect 2631 685 2635 689
rect 2815 685 2819 689
rect 2991 685 2995 689
rect 3159 685 3163 689
rect 3327 685 3331 689
rect 3479 685 3483 689
rect 1767 675 1771 679
rect 3519 679 3523 683
rect 135 659 139 663
rect 295 659 299 663
rect 463 659 467 663
rect 623 659 627 663
rect 775 659 779 663
rect 927 659 931 663
rect 1071 659 1075 663
rect 1207 659 1211 663
rect 1343 659 1347 663
rect 1479 659 1483 663
rect 1615 659 1619 663
rect 1727 659 1731 663
rect 2215 659 2219 663
rect 2359 659 2363 663
rect 2511 659 2515 663
rect 2671 659 2675 663
rect 2831 659 2835 663
rect 2991 659 2995 663
rect 3159 659 3163 663
rect 3327 659 3331 663
rect 3479 659 3483 663
rect 111 649 115 653
rect 843 651 847 655
rect 1143 651 1147 655
rect 1823 649 1827 653
rect 1863 649 1867 653
rect 2095 651 2099 655
rect 3059 651 3063 655
rect 3575 649 3579 653
rect 111 632 115 636
rect 203 635 207 639
rect 363 635 367 639
rect 1411 635 1415 639
rect 1419 635 1423 639
rect 1591 635 1595 639
rect 1683 635 1687 639
rect 1823 632 1827 636
rect 1863 632 1867 636
rect 2283 635 2287 639
rect 2427 635 2431 639
rect 2823 635 2827 639
rect 2983 635 2987 639
rect 3059 635 3063 639
rect 3227 635 3231 639
rect 3547 635 3551 639
rect 3575 632 3579 636
rect 143 619 147 623
rect 303 619 307 623
rect 471 619 475 623
rect 631 619 635 623
rect 783 619 787 623
rect 935 619 939 623
rect 1079 619 1083 623
rect 1215 619 1219 623
rect 1351 619 1355 623
rect 1419 615 1423 619
rect 1487 619 1491 623
rect 1623 619 1627 623
rect 1735 619 1739 623
rect 2223 619 2227 623
rect 2367 619 2371 623
rect 2519 619 2523 623
rect 2679 619 2683 623
rect 2839 619 2843 623
rect 2999 619 3003 623
rect 3167 619 3171 623
rect 3335 619 3339 623
rect 3487 619 3491 623
rect 203 607 207 611
rect 363 607 367 611
rect 503 607 504 611
rect 504 607 507 611
rect 663 607 664 611
rect 664 607 667 611
rect 1519 607 1520 611
rect 1520 607 1523 611
rect 1683 607 1687 611
rect 1767 607 1768 611
rect 1768 607 1771 611
rect 2283 607 2287 611
rect 2427 607 2431 611
rect 2707 607 2708 611
rect 2708 607 2711 611
rect 2823 607 2827 611
rect 3059 607 3063 611
rect 3227 607 3231 611
rect 3387 607 3391 611
rect 3519 607 3520 611
rect 3520 607 3523 611
rect 2747 599 2751 603
rect 755 591 759 595
rect 791 591 795 595
rect 1039 591 1043 595
rect 1307 591 1311 595
rect 1407 591 1408 595
rect 1408 591 1411 595
rect 1591 591 1592 595
rect 1592 591 1595 595
rect 2231 591 2232 595
rect 2232 591 2235 595
rect 2915 591 2919 595
rect 2983 591 2987 595
rect 3175 591 3176 595
rect 3176 591 3179 595
rect 3547 591 3551 595
rect 143 581 147 585
rect 303 581 307 585
rect 487 581 491 585
rect 671 581 675 585
rect 847 581 851 585
rect 1023 581 1027 585
rect 1199 581 1203 585
rect 1375 581 1379 585
rect 1559 581 1563 585
rect 1735 581 1739 585
rect 2199 581 2203 585
rect 2287 581 2291 585
rect 2375 581 2379 585
rect 2463 581 2467 585
rect 2567 581 2571 585
rect 2679 581 2683 585
rect 2815 581 2819 585
rect 2975 581 2979 585
rect 3143 581 3147 585
rect 3327 581 3331 585
rect 3487 581 3491 585
rect 111 568 115 572
rect 663 563 667 567
rect 755 563 759 567
rect 1307 563 1311 567
rect 1823 568 1827 572
rect 1863 568 1867 572
rect 2747 563 2751 567
rect 2915 563 2919 567
rect 3387 567 3391 571
rect 3575 568 3579 572
rect 111 551 115 555
rect 1703 551 1707 555
rect 1823 551 1827 555
rect 1863 551 1867 555
rect 2755 551 2759 555
rect 3575 551 3579 555
rect 135 541 139 545
rect 295 541 299 545
rect 479 541 483 545
rect 663 541 667 545
rect 839 541 843 545
rect 1015 541 1019 545
rect 1191 541 1195 545
rect 1367 541 1371 545
rect 1551 541 1555 545
rect 1727 541 1731 545
rect 2191 541 2195 545
rect 2279 541 2283 545
rect 2367 541 2371 545
rect 2455 541 2459 545
rect 2559 541 2563 545
rect 2671 541 2675 545
rect 2807 541 2811 545
rect 2967 541 2971 545
rect 3135 541 3139 545
rect 3319 541 3323 545
rect 3479 541 3483 545
rect 531 535 532 539
rect 532 535 535 539
rect 1231 535 1235 539
rect 3519 535 3523 539
rect 135 515 139 519
rect 303 515 307 519
rect 495 515 499 519
rect 679 515 683 519
rect 863 515 867 519
rect 1031 515 1035 519
rect 1191 515 1195 519
rect 1351 515 1355 519
rect 1503 515 1507 519
rect 1663 515 1667 519
rect 2303 515 2307 519
rect 2399 515 2403 519
rect 2503 515 2507 519
rect 2607 515 2611 519
rect 2719 515 2723 519
rect 2839 515 2843 519
rect 2967 515 2971 519
rect 3095 515 3099 519
rect 3223 515 3227 519
rect 3351 515 3355 519
rect 3479 515 3483 519
rect 111 505 115 509
rect 791 507 795 511
rect 1039 503 1043 507
rect 1823 505 1827 509
rect 1863 505 1867 509
rect 2231 507 2235 511
rect 3175 507 3179 511
rect 3291 507 3295 511
rect 3575 505 3579 509
rect 111 488 115 492
rect 203 491 207 495
rect 371 491 375 495
rect 747 491 751 495
rect 1419 491 1423 495
rect 1571 491 1575 495
rect 1823 488 1827 492
rect 1863 488 1867 492
rect 2371 491 2375 495
rect 2467 491 2471 495
rect 2571 491 2575 495
rect 2811 491 2815 495
rect 2907 491 2911 495
rect 3547 491 3551 495
rect 3575 488 3579 492
rect 1587 483 1591 487
rect 143 475 147 479
rect 311 475 315 479
rect 503 475 507 479
rect 687 475 691 479
rect 871 475 875 479
rect 1039 475 1043 479
rect 1199 475 1203 479
rect 1359 475 1363 479
rect 1511 475 1515 479
rect 1671 475 1675 479
rect 2311 475 2315 479
rect 2407 475 2411 479
rect 2511 475 2515 479
rect 2615 475 2619 479
rect 2727 475 2731 479
rect 2847 475 2851 479
rect 2975 475 2979 479
rect 3103 475 3107 479
rect 3231 475 3235 479
rect 3359 475 3363 479
rect 3487 475 3491 479
rect 203 463 207 467
rect 371 463 375 467
rect 531 463 532 467
rect 532 463 535 467
rect 747 463 751 467
rect 939 463 943 467
rect 1047 463 1051 467
rect 1231 463 1232 467
rect 1232 463 1235 467
rect 1571 463 1575 467
rect 1703 463 1704 467
rect 1704 463 1707 467
rect 2371 463 2375 467
rect 2467 463 2471 467
rect 2571 463 2575 467
rect 2647 463 2648 467
rect 2648 463 2651 467
rect 2755 463 2756 467
rect 2756 463 2759 467
rect 2811 463 2815 467
rect 3007 463 3008 467
rect 3008 463 3011 467
rect 3219 463 3223 467
rect 3519 463 3520 467
rect 3520 463 3523 467
rect 1095 447 1099 451
rect 1291 447 1295 451
rect 1419 447 1420 451
rect 1420 447 1423 451
rect 1587 447 1588 451
rect 1588 447 1591 451
rect 2271 451 2272 455
rect 2272 451 2275 455
rect 2907 451 2911 455
rect 3263 451 3267 455
rect 3547 451 3551 455
rect 143 437 147 441
rect 303 437 307 441
rect 495 437 499 441
rect 687 437 691 441
rect 879 437 883 441
rect 1055 437 1059 441
rect 1223 437 1227 441
rect 1391 437 1395 441
rect 1559 437 1563 441
rect 1727 437 1731 441
rect 2239 441 2243 445
rect 2327 441 2331 445
rect 2431 441 2435 445
rect 2559 441 2563 445
rect 2695 441 2699 445
rect 2847 441 2851 445
rect 2999 441 3003 445
rect 3159 441 3163 445
rect 3327 441 3331 445
rect 3487 441 3491 445
rect 111 424 115 428
rect 939 423 943 427
rect 1047 419 1051 423
rect 1291 419 1295 423
rect 1823 424 1827 428
rect 1863 428 1867 432
rect 2647 423 2651 427
rect 3219 427 3223 431
rect 3575 428 3579 432
rect 3263 423 3267 427
rect 111 407 115 411
rect 463 407 467 411
rect 1299 407 1303 411
rect 1823 407 1827 411
rect 1863 411 1867 415
rect 2999 411 3003 415
rect 3575 411 3579 415
rect 135 397 139 401
rect 295 397 299 401
rect 487 397 491 401
rect 679 397 683 401
rect 871 397 875 401
rect 1047 397 1051 401
rect 1215 397 1219 401
rect 1383 397 1387 401
rect 1551 397 1555 401
rect 1719 397 1723 401
rect 2231 401 2235 405
rect 2319 401 2323 405
rect 2423 401 2427 405
rect 2551 401 2555 405
rect 2687 401 2691 405
rect 2839 401 2843 405
rect 2991 401 2995 405
rect 3151 401 3155 405
rect 3319 401 3323 405
rect 3479 401 3483 405
rect 1767 391 1768 395
rect 1768 391 1771 395
rect 3519 395 3523 399
rect 2271 387 2275 391
rect 135 375 139 379
rect 263 375 267 379
rect 423 375 427 379
rect 591 375 595 379
rect 767 375 771 379
rect 935 375 939 379
rect 1103 375 1107 379
rect 1263 375 1267 379
rect 1423 375 1427 379
rect 1583 375 1587 379
rect 1727 375 1731 379
rect 2183 379 2187 383
rect 2287 379 2291 383
rect 2399 379 2403 383
rect 2527 379 2531 383
rect 2671 379 2675 383
rect 2815 379 2819 383
rect 2967 379 2971 383
rect 3127 379 3131 383
rect 3295 379 3299 383
rect 3463 379 3467 383
rect 111 365 115 369
rect 1095 367 1099 371
rect 1823 365 1827 369
rect 1863 369 1867 373
rect 3575 369 3579 373
rect 111 348 115 352
rect 331 351 335 355
rect 659 351 663 355
rect 1035 351 1039 355
rect 1255 351 1259 355
rect 1651 351 1655 355
rect 1659 351 1663 355
rect 1823 348 1827 352
rect 1863 352 1867 356
rect 2595 355 2599 359
rect 2883 355 2887 359
rect 3575 352 3579 356
rect 243 343 247 347
rect 143 335 147 339
rect 271 335 275 339
rect 431 335 435 339
rect 599 335 603 339
rect 775 335 779 339
rect 943 335 947 339
rect 1111 335 1115 339
rect 1271 335 1275 339
rect 1431 335 1435 339
rect 1591 335 1595 339
rect 1659 331 1663 335
rect 1735 335 1739 339
rect 2191 339 2195 343
rect 2295 339 2299 343
rect 2407 339 2411 343
rect 2535 339 2539 343
rect 2679 339 2683 343
rect 2823 339 2827 343
rect 2975 339 2979 343
rect 3135 339 3139 343
rect 3303 339 3307 343
rect 3471 339 3475 343
rect 331 323 335 327
rect 463 323 464 327
rect 464 323 467 327
rect 659 323 663 327
rect 783 323 787 327
rect 995 323 999 327
rect 1035 323 1039 327
rect 1299 323 1300 327
rect 1300 323 1303 327
rect 1767 323 1768 327
rect 1768 323 1771 327
rect 2883 327 2887 331
rect 2999 327 3003 331
rect 3155 327 3159 331
rect 243 311 244 315
rect 244 311 247 315
rect 555 311 559 315
rect 1099 311 1103 315
rect 1255 311 1256 315
rect 1256 311 1259 315
rect 1651 311 1652 315
rect 1652 311 1655 315
rect 2155 307 2159 311
rect 2363 307 2367 311
rect 2595 307 2599 311
rect 2855 307 2859 311
rect 3239 307 3243 311
rect 3519 307 3520 311
rect 3520 307 3523 311
rect 215 301 219 305
rect 351 301 355 305
rect 495 301 499 305
rect 639 301 643 305
rect 791 301 795 305
rect 935 301 939 305
rect 1079 301 1083 305
rect 1223 301 1227 305
rect 1359 301 1363 305
rect 1487 301 1491 305
rect 1623 301 1627 305
rect 1735 301 1739 305
rect 1895 297 1899 301
rect 2087 297 2091 301
rect 2303 297 2307 301
rect 2511 297 2515 301
rect 2711 297 2715 301
rect 2903 297 2907 301
rect 3095 297 3099 301
rect 3295 297 3299 301
rect 3487 297 3491 301
rect 111 288 115 292
rect 783 283 787 287
rect 995 287 999 291
rect 1823 288 1827 292
rect 1863 284 1867 288
rect 2155 279 2159 283
rect 2855 283 2859 287
rect 3155 283 3159 287
rect 3575 284 3579 288
rect 111 271 115 275
rect 1471 271 1475 275
rect 1823 271 1827 275
rect 1863 267 1867 271
rect 2987 267 2991 271
rect 3575 267 3579 271
rect 207 261 211 265
rect 343 261 347 265
rect 487 261 491 265
rect 631 261 635 265
rect 783 261 787 265
rect 927 261 931 265
rect 1071 261 1075 265
rect 1215 261 1219 265
rect 1351 261 1355 265
rect 1479 261 1483 265
rect 1615 261 1619 265
rect 1727 261 1731 265
rect 395 255 396 259
rect 396 255 399 259
rect 1887 257 1891 261
rect 2079 257 2083 261
rect 2295 257 2299 261
rect 2503 257 2507 261
rect 2703 257 2707 261
rect 2895 257 2899 261
rect 3087 257 3091 261
rect 3287 257 3291 261
rect 3479 257 3483 261
rect 1927 251 1931 255
rect 3519 251 3523 255
rect 231 231 235 235
rect 359 231 363 235
rect 487 231 491 235
rect 623 231 627 235
rect 759 231 763 235
rect 895 231 899 235
rect 1031 231 1035 235
rect 1159 231 1163 235
rect 1295 231 1299 235
rect 1431 231 1435 235
rect 1887 235 1891 239
rect 1999 235 2003 239
rect 2143 235 2147 239
rect 2295 235 2299 239
rect 2455 235 2459 239
rect 2615 235 2619 239
rect 2783 235 2787 239
rect 2951 235 2955 239
rect 3127 235 3131 239
rect 3311 235 3315 239
rect 3479 235 3483 239
rect 111 221 115 225
rect 427 223 431 227
rect 555 223 559 227
rect 1099 223 1103 227
rect 1823 221 1827 225
rect 1863 225 1867 229
rect 2079 227 2083 231
rect 2363 227 2367 231
rect 3239 227 3243 231
rect 3575 225 3579 229
rect 111 204 115 208
rect 207 207 211 211
rect 691 207 695 211
rect 1363 207 1367 211
rect 1371 207 1375 211
rect 1823 204 1827 208
rect 1863 208 1867 212
rect 2363 211 2367 215
rect 2683 211 2687 215
rect 2851 211 2855 215
rect 3195 211 3199 215
rect 3547 211 3551 215
rect 3575 208 3579 212
rect 239 191 243 195
rect 367 191 371 195
rect 427 187 431 191
rect 495 191 499 195
rect 631 191 635 195
rect 767 191 771 195
rect 903 191 907 195
rect 1039 191 1043 195
rect 1167 191 1171 195
rect 1303 191 1307 195
rect 1439 191 1443 195
rect 1895 195 1899 199
rect 2007 195 2011 199
rect 2151 195 2155 199
rect 2303 195 2307 199
rect 2463 195 2467 199
rect 2623 195 2627 199
rect 2791 195 2795 199
rect 2959 195 2963 199
rect 3135 195 3139 199
rect 3319 195 3323 199
rect 3487 195 3491 199
rect 395 179 396 183
rect 396 179 399 183
rect 691 179 695 183
rect 783 179 787 183
rect 935 179 936 183
rect 936 179 939 183
rect 1471 179 1472 183
rect 1472 179 1475 183
rect 1927 183 1928 187
rect 1928 183 1931 187
rect 2363 183 2367 187
rect 2507 183 2511 187
rect 2683 183 2687 187
rect 2851 183 2855 187
rect 2987 183 2988 187
rect 2988 183 2991 187
rect 3195 183 3199 187
rect 3371 183 3375 187
rect 3519 183 3520 187
rect 3520 183 3523 187
rect 1371 171 1375 175
rect 2079 151 2083 155
rect 207 143 208 147
rect 208 143 211 147
rect 947 143 951 147
rect 1123 143 1127 147
rect 1211 143 1215 147
rect 1363 143 1367 147
rect 2499 143 2503 147
rect 3467 143 3471 147
rect 3547 143 3551 147
rect 175 133 179 137
rect 263 133 267 137
rect 351 133 355 137
rect 439 133 443 137
rect 527 133 531 137
rect 615 133 619 137
rect 703 133 707 137
rect 791 133 795 137
rect 879 133 883 137
rect 967 133 971 137
rect 1055 133 1059 137
rect 1143 133 1147 137
rect 1231 133 1235 137
rect 1319 133 1323 137
rect 1407 133 1411 137
rect 1503 133 1507 137
rect 1895 133 1899 137
rect 1983 133 1987 137
rect 2071 133 2075 137
rect 2159 133 2163 137
rect 2247 133 2251 137
rect 2335 133 2339 137
rect 2439 133 2443 137
rect 2543 133 2547 137
rect 2647 133 2651 137
rect 2743 133 2747 137
rect 2839 133 2843 137
rect 2935 133 2939 137
rect 3031 133 3035 137
rect 3127 133 3131 137
rect 3223 133 3227 137
rect 3311 133 3315 137
rect 3399 133 3403 137
rect 3487 133 3491 137
rect 935 127 939 131
rect 111 120 115 124
rect 783 115 787 119
rect 947 115 951 119
rect 1123 115 1127 119
rect 1211 115 1215 119
rect 1823 120 1827 124
rect 1863 120 1867 124
rect 2499 119 2503 123
rect 2507 115 2511 119
rect 3371 119 3375 123
rect 3575 120 3579 124
rect 3467 115 3471 119
rect 111 103 115 107
rect 1823 103 1827 107
rect 1863 103 1867 107
rect 3575 103 3579 107
rect 167 93 171 97
rect 255 93 259 97
rect 343 93 347 97
rect 431 93 435 97
rect 519 93 523 97
rect 607 93 611 97
rect 695 93 699 97
rect 783 93 787 97
rect 871 93 875 97
rect 959 93 963 97
rect 1047 93 1051 97
rect 1135 93 1139 97
rect 1223 93 1227 97
rect 1311 93 1315 97
rect 1399 93 1403 97
rect 1495 93 1499 97
rect 1887 93 1891 97
rect 1975 93 1979 97
rect 2063 93 2067 97
rect 2151 93 2155 97
rect 2239 93 2243 97
rect 2327 93 2331 97
rect 2431 93 2435 97
rect 2535 93 2539 97
rect 2639 93 2643 97
rect 2735 93 2739 97
rect 2831 93 2835 97
rect 2927 93 2931 97
rect 3023 93 3027 97
rect 3119 93 3123 97
rect 3215 93 3219 97
rect 3303 93 3307 97
rect 3391 93 3395 97
rect 3479 93 3483 97
<< m3 >>
rect 111 3650 115 3651
rect 111 3645 115 3646
rect 239 3650 243 3651
rect 239 3645 243 3646
rect 327 3650 331 3651
rect 327 3645 331 3646
rect 415 3650 419 3651
rect 415 3645 419 3646
rect 503 3650 507 3651
rect 503 3645 507 3646
rect 591 3650 595 3651
rect 591 3645 595 3646
rect 679 3650 683 3651
rect 679 3645 683 3646
rect 1823 3650 1827 3651
rect 1823 3645 1827 3646
rect 112 3621 114 3645
rect 240 3634 242 3645
rect 306 3643 312 3644
rect 306 3639 307 3643
rect 311 3639 312 3643
rect 306 3638 312 3639
rect 238 3633 244 3634
rect 238 3629 239 3633
rect 243 3629 244 3633
rect 238 3628 244 3629
rect 110 3620 116 3621
rect 110 3616 111 3620
rect 115 3616 116 3620
rect 308 3616 310 3638
rect 328 3634 330 3645
rect 394 3643 400 3644
rect 394 3639 395 3643
rect 399 3639 400 3643
rect 394 3638 400 3639
rect 326 3633 332 3634
rect 326 3629 327 3633
rect 331 3629 332 3633
rect 326 3628 332 3629
rect 396 3616 398 3638
rect 416 3634 418 3645
rect 482 3643 488 3644
rect 482 3639 483 3643
rect 487 3639 488 3643
rect 482 3638 488 3639
rect 414 3633 420 3634
rect 414 3629 415 3633
rect 419 3629 420 3633
rect 414 3628 420 3629
rect 484 3616 486 3638
rect 504 3634 506 3645
rect 570 3643 576 3644
rect 570 3639 571 3643
rect 575 3639 576 3643
rect 570 3638 576 3639
rect 502 3633 508 3634
rect 502 3629 503 3633
rect 507 3629 508 3633
rect 502 3628 508 3629
rect 572 3616 574 3638
rect 592 3634 594 3645
rect 658 3643 664 3644
rect 658 3639 659 3643
rect 663 3639 664 3643
rect 658 3638 664 3639
rect 590 3633 596 3634
rect 590 3629 591 3633
rect 595 3629 596 3633
rect 590 3628 596 3629
rect 660 3616 662 3638
rect 680 3634 682 3645
rect 678 3633 684 3634
rect 678 3629 679 3633
rect 683 3629 684 3633
rect 678 3628 684 3629
rect 1824 3621 1826 3645
rect 1822 3620 1828 3621
rect 1822 3616 1823 3620
rect 1827 3616 1828 3620
rect 110 3615 116 3616
rect 306 3615 312 3616
rect 306 3611 307 3615
rect 311 3611 312 3615
rect 306 3610 312 3611
rect 394 3615 400 3616
rect 394 3611 395 3615
rect 399 3611 400 3615
rect 394 3610 400 3611
rect 482 3615 488 3616
rect 482 3611 483 3615
rect 487 3611 488 3615
rect 482 3610 488 3611
rect 570 3615 576 3616
rect 570 3611 571 3615
rect 575 3611 576 3615
rect 570 3610 576 3611
rect 658 3615 664 3616
rect 1822 3615 1828 3616
rect 658 3611 659 3615
rect 663 3611 664 3615
rect 658 3610 664 3611
rect 110 3603 116 3604
rect 110 3599 111 3603
rect 115 3599 116 3603
rect 110 3598 116 3599
rect 1822 3603 1828 3604
rect 1822 3599 1823 3603
rect 1827 3599 1828 3603
rect 1822 3598 1828 3599
rect 112 3575 114 3598
rect 230 3593 236 3594
rect 230 3589 231 3593
rect 235 3589 236 3593
rect 230 3588 236 3589
rect 318 3593 324 3594
rect 318 3589 319 3593
rect 323 3589 324 3593
rect 318 3588 324 3589
rect 406 3593 412 3594
rect 406 3589 407 3593
rect 411 3589 412 3593
rect 406 3588 412 3589
rect 494 3593 500 3594
rect 494 3589 495 3593
rect 499 3589 500 3593
rect 494 3588 500 3589
rect 582 3593 588 3594
rect 582 3589 583 3593
rect 587 3589 588 3593
rect 582 3588 588 3589
rect 670 3593 676 3594
rect 670 3589 671 3593
rect 675 3589 676 3593
rect 670 3588 676 3589
rect 232 3575 234 3588
rect 282 3587 288 3588
rect 282 3583 283 3587
rect 287 3583 288 3587
rect 282 3582 288 3583
rect 111 3574 115 3575
rect 111 3569 115 3570
rect 231 3574 235 3575
rect 231 3569 235 3570
rect 247 3574 251 3575
rect 247 3569 251 3570
rect 112 3554 114 3569
rect 248 3564 250 3569
rect 246 3563 252 3564
rect 246 3559 247 3563
rect 251 3559 252 3563
rect 246 3558 252 3559
rect 110 3553 116 3554
rect 110 3549 111 3553
rect 115 3549 116 3553
rect 110 3548 116 3549
rect 110 3536 116 3537
rect 110 3532 111 3536
rect 115 3532 116 3536
rect 110 3531 116 3532
rect 112 3507 114 3531
rect 254 3523 260 3524
rect 254 3519 255 3523
rect 259 3519 260 3523
rect 254 3518 260 3519
rect 256 3507 258 3518
rect 284 3512 286 3582
rect 320 3575 322 3588
rect 408 3575 410 3588
rect 496 3575 498 3588
rect 584 3575 586 3588
rect 672 3575 674 3588
rect 1824 3575 1826 3598
rect 1863 3586 1867 3587
rect 1863 3581 1867 3582
rect 1887 3586 1891 3587
rect 1887 3581 1891 3582
rect 1975 3586 1979 3587
rect 1975 3581 1979 3582
rect 2063 3586 2067 3587
rect 2063 3581 2067 3582
rect 2151 3586 2155 3587
rect 2151 3581 2155 3582
rect 2239 3586 2243 3587
rect 2239 3581 2243 3582
rect 2327 3586 2331 3587
rect 2327 3581 2331 3582
rect 2415 3586 2419 3587
rect 2415 3581 2419 3582
rect 2503 3586 2507 3587
rect 2503 3581 2507 3582
rect 2591 3586 2595 3587
rect 2591 3581 2595 3582
rect 2679 3586 2683 3587
rect 2679 3581 2683 3582
rect 2767 3586 2771 3587
rect 2767 3581 2771 3582
rect 2855 3586 2859 3587
rect 2855 3581 2859 3582
rect 2943 3586 2947 3587
rect 2943 3581 2947 3582
rect 3031 3586 3035 3587
rect 3031 3581 3035 3582
rect 3119 3586 3123 3587
rect 3119 3581 3123 3582
rect 3207 3586 3211 3587
rect 3207 3581 3211 3582
rect 3295 3586 3299 3587
rect 3295 3581 3299 3582
rect 3575 3586 3579 3587
rect 3575 3581 3579 3582
rect 319 3574 323 3575
rect 319 3569 323 3570
rect 399 3574 403 3575
rect 399 3569 403 3570
rect 407 3574 411 3575
rect 407 3569 411 3570
rect 495 3574 499 3575
rect 495 3569 499 3570
rect 543 3574 547 3575
rect 543 3569 547 3570
rect 583 3574 587 3575
rect 583 3569 587 3570
rect 671 3574 675 3575
rect 671 3569 675 3570
rect 687 3574 691 3575
rect 687 3569 691 3570
rect 823 3574 827 3575
rect 823 3569 827 3570
rect 951 3574 955 3575
rect 951 3569 955 3570
rect 1079 3574 1083 3575
rect 1079 3569 1083 3570
rect 1199 3574 1203 3575
rect 1199 3569 1203 3570
rect 1311 3574 1315 3575
rect 1311 3569 1315 3570
rect 1423 3574 1427 3575
rect 1423 3569 1427 3570
rect 1543 3574 1547 3575
rect 1543 3569 1547 3570
rect 1823 3574 1827 3575
rect 1823 3569 1827 3570
rect 400 3564 402 3569
rect 544 3564 546 3569
rect 688 3564 690 3569
rect 824 3564 826 3569
rect 952 3564 954 3569
rect 1080 3564 1082 3569
rect 1200 3564 1202 3569
rect 1312 3564 1314 3569
rect 1424 3564 1426 3569
rect 1544 3564 1546 3569
rect 398 3563 404 3564
rect 398 3559 399 3563
rect 403 3559 404 3563
rect 398 3558 404 3559
rect 542 3563 548 3564
rect 542 3559 543 3563
rect 547 3559 548 3563
rect 542 3558 548 3559
rect 686 3563 692 3564
rect 686 3559 687 3563
rect 691 3559 692 3563
rect 686 3558 692 3559
rect 822 3563 828 3564
rect 822 3559 823 3563
rect 827 3559 828 3563
rect 822 3558 828 3559
rect 950 3563 956 3564
rect 950 3559 951 3563
rect 955 3559 956 3563
rect 950 3558 956 3559
rect 1078 3563 1084 3564
rect 1078 3559 1079 3563
rect 1083 3559 1084 3563
rect 1078 3558 1084 3559
rect 1198 3563 1204 3564
rect 1198 3559 1199 3563
rect 1203 3559 1204 3563
rect 1198 3558 1204 3559
rect 1310 3563 1316 3564
rect 1310 3559 1311 3563
rect 1315 3559 1316 3563
rect 1310 3558 1316 3559
rect 1422 3563 1428 3564
rect 1422 3559 1423 3563
rect 1427 3559 1428 3563
rect 1422 3558 1428 3559
rect 1542 3563 1548 3564
rect 1542 3559 1543 3563
rect 1547 3559 1548 3563
rect 1542 3558 1548 3559
rect 1490 3555 1496 3556
rect 1490 3551 1491 3555
rect 1495 3551 1496 3555
rect 1824 3554 1826 3569
rect 1864 3566 1866 3581
rect 1888 3576 1890 3581
rect 1976 3576 1978 3581
rect 2064 3576 2066 3581
rect 2152 3576 2154 3581
rect 2240 3576 2242 3581
rect 2328 3576 2330 3581
rect 2416 3576 2418 3581
rect 2504 3576 2506 3581
rect 2592 3576 2594 3581
rect 2680 3576 2682 3581
rect 2768 3576 2770 3581
rect 2856 3576 2858 3581
rect 2944 3576 2946 3581
rect 3032 3576 3034 3581
rect 3120 3576 3122 3581
rect 3208 3576 3210 3581
rect 3296 3576 3298 3581
rect 1886 3575 1892 3576
rect 1886 3571 1887 3575
rect 1891 3571 1892 3575
rect 1886 3570 1892 3571
rect 1974 3575 1980 3576
rect 1974 3571 1975 3575
rect 1979 3571 1980 3575
rect 1974 3570 1980 3571
rect 2062 3575 2068 3576
rect 2062 3571 2063 3575
rect 2067 3571 2068 3575
rect 2062 3570 2068 3571
rect 2150 3575 2156 3576
rect 2150 3571 2151 3575
rect 2155 3571 2156 3575
rect 2150 3570 2156 3571
rect 2238 3575 2244 3576
rect 2238 3571 2239 3575
rect 2243 3571 2244 3575
rect 2238 3570 2244 3571
rect 2326 3575 2332 3576
rect 2326 3571 2327 3575
rect 2331 3571 2332 3575
rect 2326 3570 2332 3571
rect 2414 3575 2420 3576
rect 2414 3571 2415 3575
rect 2419 3571 2420 3575
rect 2414 3570 2420 3571
rect 2502 3575 2508 3576
rect 2502 3571 2503 3575
rect 2507 3571 2508 3575
rect 2502 3570 2508 3571
rect 2590 3575 2596 3576
rect 2590 3571 2591 3575
rect 2595 3571 2596 3575
rect 2590 3570 2596 3571
rect 2678 3575 2684 3576
rect 2678 3571 2679 3575
rect 2683 3571 2684 3575
rect 2678 3570 2684 3571
rect 2766 3575 2772 3576
rect 2766 3571 2767 3575
rect 2771 3571 2772 3575
rect 2766 3570 2772 3571
rect 2854 3575 2860 3576
rect 2854 3571 2855 3575
rect 2859 3571 2860 3575
rect 2854 3570 2860 3571
rect 2942 3575 2948 3576
rect 2942 3571 2943 3575
rect 2947 3571 2948 3575
rect 2942 3570 2948 3571
rect 3030 3575 3036 3576
rect 3030 3571 3031 3575
rect 3035 3571 3036 3575
rect 3030 3570 3036 3571
rect 3118 3575 3124 3576
rect 3118 3571 3119 3575
rect 3123 3571 3124 3575
rect 3118 3570 3124 3571
rect 3206 3575 3212 3576
rect 3206 3571 3207 3575
rect 3211 3571 3212 3575
rect 3206 3570 3212 3571
rect 3294 3575 3300 3576
rect 3294 3571 3295 3575
rect 3299 3571 3300 3575
rect 3294 3570 3300 3571
rect 3274 3567 3280 3568
rect 1862 3565 1868 3566
rect 1862 3561 1863 3565
rect 1867 3561 1868 3565
rect 3274 3563 3275 3567
rect 3279 3563 3280 3567
rect 3576 3566 3578 3581
rect 3274 3562 3280 3563
rect 3574 3565 3580 3566
rect 1862 3560 1868 3561
rect 1490 3550 1496 3551
rect 1822 3553 1828 3554
rect 754 3539 760 3540
rect 754 3535 755 3539
rect 759 3535 760 3539
rect 754 3534 760 3535
rect 1034 3539 1040 3540
rect 1034 3535 1035 3539
rect 1039 3535 1040 3539
rect 1034 3534 1040 3535
rect 406 3523 412 3524
rect 406 3519 407 3523
rect 411 3519 412 3523
rect 406 3518 412 3519
rect 550 3523 556 3524
rect 550 3519 551 3523
rect 555 3519 556 3523
rect 550 3518 556 3519
rect 694 3523 700 3524
rect 694 3519 695 3523
rect 699 3519 700 3523
rect 694 3518 700 3519
rect 282 3511 288 3512
rect 282 3507 283 3511
rect 287 3507 288 3511
rect 408 3507 410 3518
rect 552 3507 554 3518
rect 696 3507 698 3518
rect 111 3506 115 3507
rect 111 3501 115 3502
rect 183 3506 187 3507
rect 183 3501 187 3502
rect 255 3506 259 3507
rect 282 3506 288 3507
rect 351 3506 355 3507
rect 255 3501 259 3502
rect 351 3501 355 3502
rect 407 3506 411 3507
rect 407 3501 411 3502
rect 519 3506 523 3507
rect 519 3501 523 3502
rect 551 3506 555 3507
rect 551 3501 555 3502
rect 679 3506 683 3507
rect 679 3501 683 3502
rect 695 3506 699 3507
rect 695 3501 699 3502
rect 112 3477 114 3501
rect 184 3490 186 3501
rect 352 3490 354 3501
rect 454 3499 460 3500
rect 454 3495 455 3499
rect 459 3495 460 3499
rect 454 3494 460 3495
rect 182 3489 188 3490
rect 182 3485 183 3489
rect 187 3485 188 3489
rect 182 3484 188 3485
rect 350 3489 356 3490
rect 350 3485 351 3489
rect 355 3485 356 3489
rect 350 3484 356 3485
rect 110 3476 116 3477
rect 110 3472 111 3476
rect 115 3472 116 3476
rect 456 3472 458 3494
rect 520 3490 522 3501
rect 680 3490 682 3501
rect 756 3500 758 3534
rect 830 3523 836 3524
rect 830 3519 831 3523
rect 835 3519 836 3523
rect 830 3518 836 3519
rect 958 3523 964 3524
rect 958 3519 959 3523
rect 963 3519 964 3523
rect 958 3518 964 3519
rect 832 3507 834 3518
rect 890 3511 896 3512
rect 890 3507 891 3511
rect 895 3507 896 3511
rect 960 3507 962 3518
rect 1036 3512 1038 3534
rect 1086 3523 1092 3524
rect 1086 3519 1087 3523
rect 1091 3519 1092 3523
rect 1086 3518 1092 3519
rect 1206 3523 1212 3524
rect 1206 3519 1207 3523
rect 1211 3519 1212 3523
rect 1206 3518 1212 3519
rect 1318 3523 1324 3524
rect 1318 3519 1319 3523
rect 1323 3519 1324 3523
rect 1318 3518 1324 3519
rect 1430 3523 1436 3524
rect 1430 3519 1431 3523
rect 1435 3519 1436 3523
rect 1430 3518 1436 3519
rect 1034 3511 1040 3512
rect 1034 3507 1035 3511
rect 1039 3507 1040 3511
rect 1088 3507 1090 3518
rect 1208 3507 1210 3518
rect 1247 3516 1251 3517
rect 1247 3511 1251 3512
rect 831 3506 835 3507
rect 890 3506 896 3507
rect 959 3506 963 3507
rect 831 3501 835 3502
rect 754 3499 760 3500
rect 754 3495 755 3499
rect 759 3495 760 3499
rect 754 3494 760 3495
rect 832 3490 834 3501
rect 518 3489 524 3490
rect 518 3485 519 3489
rect 523 3485 524 3489
rect 518 3484 524 3485
rect 678 3489 684 3490
rect 678 3485 679 3489
rect 683 3485 684 3489
rect 678 3484 684 3485
rect 830 3489 836 3490
rect 830 3485 831 3489
rect 835 3485 836 3489
rect 830 3484 836 3485
rect 892 3476 894 3506
rect 959 3501 963 3502
rect 967 3506 971 3507
rect 1034 3506 1040 3507
rect 1087 3506 1091 3507
rect 967 3501 971 3502
rect 1087 3501 1091 3502
rect 1095 3506 1099 3507
rect 1095 3501 1099 3502
rect 1207 3506 1211 3507
rect 1207 3501 1211 3502
rect 1215 3506 1219 3507
rect 1215 3501 1219 3502
rect 968 3490 970 3501
rect 978 3499 984 3500
rect 978 3495 979 3499
rect 983 3495 984 3499
rect 978 3494 984 3495
rect 1006 3499 1012 3500
rect 1006 3495 1007 3499
rect 1011 3495 1012 3499
rect 1006 3494 1012 3495
rect 966 3489 972 3490
rect 966 3485 967 3489
rect 971 3485 972 3489
rect 966 3484 972 3485
rect 890 3475 896 3476
rect 110 3471 116 3472
rect 454 3471 460 3472
rect 454 3467 455 3471
rect 459 3467 460 3471
rect 890 3471 891 3475
rect 895 3471 896 3475
rect 890 3470 896 3471
rect 454 3466 460 3467
rect 110 3459 116 3460
rect 110 3455 111 3459
rect 115 3455 116 3459
rect 110 3454 116 3455
rect 270 3459 276 3460
rect 270 3455 271 3459
rect 275 3455 276 3459
rect 270 3454 276 3455
rect 112 3439 114 3454
rect 174 3449 180 3450
rect 174 3445 175 3449
rect 179 3445 180 3449
rect 174 3444 180 3445
rect 176 3439 178 3444
rect 111 3438 115 3439
rect 111 3433 115 3434
rect 135 3438 139 3439
rect 135 3433 139 3434
rect 175 3438 179 3439
rect 175 3433 179 3434
rect 255 3438 259 3439
rect 255 3433 259 3434
rect 112 3418 114 3433
rect 136 3428 138 3433
rect 256 3428 258 3433
rect 134 3427 140 3428
rect 134 3423 135 3427
rect 139 3423 140 3427
rect 134 3422 140 3423
rect 254 3427 260 3428
rect 254 3423 255 3427
rect 259 3423 260 3427
rect 254 3422 260 3423
rect 110 3417 116 3418
rect 110 3413 111 3417
rect 115 3413 116 3417
rect 110 3412 116 3413
rect 218 3403 224 3404
rect 110 3400 116 3401
rect 110 3396 111 3400
rect 115 3396 116 3400
rect 218 3399 219 3403
rect 223 3399 224 3403
rect 218 3398 224 3399
rect 110 3395 116 3396
rect 112 3363 114 3395
rect 142 3387 148 3388
rect 142 3383 143 3387
rect 147 3383 148 3387
rect 142 3382 148 3383
rect 144 3363 146 3382
rect 220 3368 222 3398
rect 262 3387 268 3388
rect 262 3383 263 3387
rect 267 3383 268 3387
rect 262 3382 268 3383
rect 218 3367 224 3368
rect 218 3363 219 3367
rect 223 3363 224 3367
rect 264 3363 266 3382
rect 272 3376 274 3454
rect 342 3449 348 3450
rect 342 3445 343 3449
rect 347 3445 348 3449
rect 342 3444 348 3445
rect 510 3449 516 3450
rect 510 3445 511 3449
rect 515 3445 516 3449
rect 510 3444 516 3445
rect 670 3449 676 3450
rect 670 3445 671 3449
rect 675 3445 676 3449
rect 670 3444 676 3445
rect 822 3449 828 3450
rect 822 3445 823 3449
rect 827 3445 828 3449
rect 822 3444 828 3445
rect 958 3449 964 3450
rect 958 3445 959 3449
rect 963 3445 964 3449
rect 958 3444 964 3445
rect 980 3444 982 3494
rect 344 3439 346 3444
rect 512 3439 514 3444
rect 672 3439 674 3444
rect 824 3439 826 3444
rect 960 3439 962 3444
rect 978 3443 984 3444
rect 978 3439 979 3443
rect 983 3439 984 3443
rect 343 3438 347 3439
rect 343 3433 347 3434
rect 415 3438 419 3439
rect 415 3433 419 3434
rect 511 3438 515 3439
rect 511 3433 515 3434
rect 583 3438 587 3439
rect 583 3433 587 3434
rect 671 3438 675 3439
rect 671 3433 675 3434
rect 759 3438 763 3439
rect 759 3433 763 3434
rect 823 3438 827 3439
rect 823 3433 827 3434
rect 935 3438 939 3439
rect 935 3433 939 3434
rect 959 3438 963 3439
rect 978 3438 984 3439
rect 959 3433 963 3434
rect 416 3428 418 3433
rect 584 3428 586 3433
rect 760 3428 762 3433
rect 936 3428 938 3433
rect 414 3427 420 3428
rect 414 3423 415 3427
rect 419 3423 420 3427
rect 414 3422 420 3423
rect 582 3427 588 3428
rect 582 3423 583 3427
rect 587 3423 588 3427
rect 582 3422 588 3423
rect 758 3427 764 3428
rect 758 3423 759 3427
rect 763 3423 764 3427
rect 758 3422 764 3423
rect 934 3427 940 3428
rect 934 3423 935 3427
rect 939 3423 940 3427
rect 934 3422 940 3423
rect 1008 3420 1010 3494
rect 1096 3490 1098 3501
rect 1216 3490 1218 3501
rect 1248 3500 1250 3511
rect 1320 3507 1322 3518
rect 1432 3507 1434 3518
rect 1492 3517 1494 3550
rect 1822 3549 1823 3553
rect 1827 3549 1828 3553
rect 2570 3551 2576 3552
rect 1822 3548 1828 3549
rect 1862 3548 1868 3549
rect 1862 3544 1863 3548
rect 1867 3544 1868 3548
rect 2570 3547 2571 3551
rect 2575 3547 2576 3551
rect 2570 3546 2576 3547
rect 1862 3543 1868 3544
rect 1822 3536 1828 3537
rect 1822 3532 1823 3536
rect 1827 3532 1828 3536
rect 1822 3531 1828 3532
rect 1550 3523 1556 3524
rect 1550 3519 1551 3523
rect 1555 3519 1556 3523
rect 1550 3518 1556 3519
rect 1491 3516 1495 3517
rect 1491 3511 1495 3512
rect 1552 3507 1554 3518
rect 1824 3507 1826 3531
rect 1864 3511 1866 3543
rect 1894 3535 1900 3536
rect 1894 3531 1895 3535
rect 1899 3531 1900 3535
rect 1894 3530 1900 3531
rect 1982 3535 1988 3536
rect 1982 3531 1983 3535
rect 1987 3531 1988 3535
rect 1982 3530 1988 3531
rect 2070 3535 2076 3536
rect 2070 3531 2071 3535
rect 2075 3531 2076 3535
rect 2070 3530 2076 3531
rect 2158 3535 2164 3536
rect 2158 3531 2159 3535
rect 2163 3531 2164 3535
rect 2158 3530 2164 3531
rect 2246 3535 2252 3536
rect 2246 3531 2247 3535
rect 2251 3531 2252 3535
rect 2246 3530 2252 3531
rect 2334 3535 2340 3536
rect 2334 3531 2335 3535
rect 2339 3531 2340 3535
rect 2334 3530 2340 3531
rect 2422 3535 2428 3536
rect 2422 3531 2423 3535
rect 2427 3531 2428 3535
rect 2422 3530 2428 3531
rect 2510 3535 2516 3536
rect 2510 3531 2511 3535
rect 2515 3531 2516 3535
rect 2510 3530 2516 3531
rect 1896 3511 1898 3530
rect 1902 3523 1908 3524
rect 1902 3519 1903 3523
rect 1907 3519 1908 3523
rect 1902 3518 1908 3519
rect 1863 3510 1867 3511
rect 1319 3506 1323 3507
rect 1319 3501 1323 3502
rect 1335 3506 1339 3507
rect 1335 3501 1339 3502
rect 1431 3506 1435 3507
rect 1431 3501 1435 3502
rect 1455 3506 1459 3507
rect 1455 3501 1459 3502
rect 1551 3506 1555 3507
rect 1551 3501 1555 3502
rect 1575 3506 1579 3507
rect 1575 3501 1579 3502
rect 1823 3506 1827 3507
rect 1863 3505 1867 3506
rect 1895 3510 1899 3511
rect 1895 3505 1899 3506
rect 1823 3501 1827 3502
rect 1246 3499 1252 3500
rect 1246 3495 1247 3499
rect 1251 3495 1252 3499
rect 1246 3494 1252 3495
rect 1336 3490 1338 3501
rect 1456 3490 1458 3501
rect 1576 3490 1578 3501
rect 1094 3489 1100 3490
rect 1094 3485 1095 3489
rect 1099 3485 1100 3489
rect 1094 3484 1100 3485
rect 1214 3489 1220 3490
rect 1214 3485 1215 3489
rect 1219 3485 1220 3489
rect 1214 3484 1220 3485
rect 1334 3489 1340 3490
rect 1334 3485 1335 3489
rect 1339 3485 1340 3489
rect 1334 3484 1340 3485
rect 1454 3489 1460 3490
rect 1454 3485 1455 3489
rect 1459 3485 1460 3489
rect 1454 3484 1460 3485
rect 1574 3489 1580 3490
rect 1574 3485 1575 3489
rect 1579 3485 1580 3489
rect 1574 3484 1580 3485
rect 1824 3477 1826 3501
rect 1864 3481 1866 3505
rect 1862 3480 1868 3481
rect 1822 3476 1828 3477
rect 1822 3472 1823 3476
rect 1827 3472 1828 3476
rect 1862 3476 1863 3480
rect 1867 3476 1868 3480
rect 1904 3476 1906 3518
rect 1984 3511 1986 3530
rect 2072 3511 2074 3530
rect 2160 3511 2162 3530
rect 2248 3511 2250 3530
rect 2336 3511 2338 3530
rect 2424 3511 2426 3530
rect 2512 3511 2514 3530
rect 1911 3510 1915 3511
rect 1911 3505 1915 3506
rect 1983 3510 1987 3511
rect 1983 3505 1987 3506
rect 2015 3510 2019 3511
rect 2015 3505 2019 3506
rect 2071 3510 2075 3511
rect 2071 3505 2075 3506
rect 2135 3510 2139 3511
rect 2135 3505 2139 3506
rect 2159 3510 2163 3511
rect 2159 3505 2163 3506
rect 2247 3510 2251 3511
rect 2247 3505 2251 3506
rect 2263 3510 2267 3511
rect 2263 3505 2267 3506
rect 2335 3510 2339 3511
rect 2335 3505 2339 3506
rect 2391 3510 2395 3511
rect 2391 3505 2395 3506
rect 2423 3510 2427 3511
rect 2423 3505 2427 3506
rect 2511 3510 2515 3511
rect 2511 3505 2515 3506
rect 2527 3510 2531 3511
rect 2527 3505 2531 3506
rect 1912 3494 1914 3505
rect 2016 3494 2018 3505
rect 2082 3503 2088 3504
rect 2082 3499 2083 3503
rect 2087 3499 2088 3503
rect 2082 3498 2088 3499
rect 1910 3493 1916 3494
rect 1910 3489 1911 3493
rect 1915 3489 1916 3493
rect 1910 3488 1916 3489
rect 2014 3493 2020 3494
rect 2014 3489 2015 3493
rect 2019 3489 2020 3493
rect 2014 3488 2020 3489
rect 2084 3476 2086 3498
rect 2136 3494 2138 3505
rect 2142 3503 2148 3504
rect 2142 3499 2143 3503
rect 2147 3499 2148 3503
rect 2142 3498 2148 3499
rect 2134 3493 2140 3494
rect 2134 3489 2135 3493
rect 2139 3489 2140 3493
rect 2134 3488 2140 3489
rect 1862 3475 1868 3476
rect 1902 3475 1908 3476
rect 1822 3471 1828 3472
rect 1902 3471 1903 3475
rect 1907 3471 1908 3475
rect 1902 3470 1908 3471
rect 2082 3475 2088 3476
rect 2082 3471 2083 3475
rect 2087 3471 2088 3475
rect 2082 3470 2088 3471
rect 1862 3463 1868 3464
rect 1822 3459 1828 3460
rect 1822 3455 1823 3459
rect 1827 3455 1828 3459
rect 1862 3459 1863 3463
rect 1867 3459 1868 3463
rect 1862 3458 1868 3459
rect 1822 3454 1828 3455
rect 1086 3449 1092 3450
rect 1086 3445 1087 3449
rect 1091 3445 1092 3449
rect 1086 3444 1092 3445
rect 1206 3449 1212 3450
rect 1206 3445 1207 3449
rect 1211 3445 1212 3449
rect 1206 3444 1212 3445
rect 1326 3449 1332 3450
rect 1326 3445 1327 3449
rect 1331 3445 1332 3449
rect 1326 3444 1332 3445
rect 1446 3449 1452 3450
rect 1446 3445 1447 3449
rect 1451 3445 1452 3449
rect 1446 3444 1452 3445
rect 1566 3449 1572 3450
rect 1566 3445 1567 3449
rect 1571 3445 1572 3449
rect 1566 3444 1572 3445
rect 1088 3439 1090 3444
rect 1208 3439 1210 3444
rect 1328 3439 1330 3444
rect 1334 3443 1340 3444
rect 1334 3439 1335 3443
rect 1339 3439 1340 3443
rect 1448 3439 1450 3444
rect 1568 3439 1570 3444
rect 1824 3439 1826 3454
rect 1087 3438 1091 3439
rect 1087 3433 1091 3434
rect 1111 3438 1115 3439
rect 1111 3433 1115 3434
rect 1207 3438 1211 3439
rect 1207 3433 1211 3434
rect 1295 3438 1299 3439
rect 1295 3433 1299 3434
rect 1327 3438 1331 3439
rect 1334 3438 1340 3439
rect 1447 3438 1451 3439
rect 1327 3433 1331 3434
rect 1112 3428 1114 3433
rect 1296 3428 1298 3433
rect 1110 3427 1116 3428
rect 1110 3423 1111 3427
rect 1115 3423 1116 3427
rect 1110 3422 1116 3423
rect 1294 3427 1300 3428
rect 1294 3423 1295 3427
rect 1299 3423 1300 3427
rect 1294 3422 1300 3423
rect 678 3419 684 3420
rect 678 3415 679 3419
rect 683 3415 684 3419
rect 678 3414 684 3415
rect 1006 3419 1012 3420
rect 1006 3415 1007 3419
rect 1011 3415 1012 3419
rect 1006 3414 1012 3415
rect 422 3387 428 3388
rect 422 3383 423 3387
rect 427 3383 428 3387
rect 422 3382 428 3383
rect 590 3387 596 3388
rect 590 3383 591 3387
rect 595 3383 596 3387
rect 590 3382 596 3383
rect 270 3375 276 3376
rect 270 3371 271 3375
rect 275 3371 276 3375
rect 270 3370 276 3371
rect 424 3363 426 3382
rect 592 3363 594 3382
rect 680 3364 682 3414
rect 1002 3403 1008 3404
rect 1002 3399 1003 3403
rect 1007 3399 1008 3403
rect 1002 3398 1008 3399
rect 766 3387 772 3388
rect 766 3383 767 3387
rect 771 3383 772 3387
rect 766 3382 772 3383
rect 942 3387 948 3388
rect 942 3383 943 3387
rect 947 3383 948 3387
rect 942 3382 948 3383
rect 678 3363 684 3364
rect 768 3363 770 3382
rect 944 3363 946 3382
rect 1004 3376 1006 3398
rect 1118 3387 1124 3388
rect 1118 3383 1119 3387
rect 1123 3383 1124 3387
rect 1118 3382 1124 3383
rect 1302 3387 1308 3388
rect 1302 3383 1303 3387
rect 1307 3383 1308 3387
rect 1302 3382 1308 3383
rect 1002 3375 1008 3376
rect 1002 3371 1003 3375
rect 1007 3371 1008 3375
rect 1002 3370 1008 3371
rect 1120 3363 1122 3382
rect 1134 3375 1140 3376
rect 1134 3371 1135 3375
rect 1139 3371 1140 3375
rect 1134 3370 1140 3371
rect 111 3362 115 3363
rect 111 3357 115 3358
rect 143 3362 147 3363
rect 143 3357 147 3358
rect 207 3362 211 3363
rect 218 3362 224 3363
rect 263 3362 267 3363
rect 207 3357 211 3358
rect 263 3357 267 3358
rect 367 3362 371 3363
rect 367 3357 371 3358
rect 423 3362 427 3363
rect 423 3357 427 3358
rect 535 3362 539 3363
rect 535 3357 539 3358
rect 591 3362 595 3363
rect 678 3359 679 3363
rect 683 3359 684 3363
rect 678 3358 684 3359
rect 695 3362 699 3363
rect 591 3357 595 3358
rect 695 3357 699 3358
rect 767 3362 771 3363
rect 767 3357 771 3358
rect 855 3362 859 3363
rect 855 3357 859 3358
rect 943 3362 947 3363
rect 943 3357 947 3358
rect 999 3362 1003 3363
rect 999 3357 1003 3358
rect 1119 3362 1123 3363
rect 1119 3357 1123 3358
rect 112 3333 114 3357
rect 208 3346 210 3357
rect 368 3346 370 3357
rect 536 3346 538 3357
rect 696 3346 698 3357
rect 856 3346 858 3357
rect 950 3355 956 3356
rect 950 3351 951 3355
rect 955 3351 956 3355
rect 950 3350 956 3351
rect 206 3345 212 3346
rect 206 3341 207 3345
rect 211 3341 212 3345
rect 206 3340 212 3341
rect 366 3345 372 3346
rect 366 3341 367 3345
rect 371 3341 372 3345
rect 366 3340 372 3341
rect 534 3345 540 3346
rect 534 3341 535 3345
rect 539 3341 540 3345
rect 534 3340 540 3341
rect 694 3345 700 3346
rect 694 3341 695 3345
rect 699 3341 700 3345
rect 694 3340 700 3341
rect 854 3345 860 3346
rect 854 3341 855 3345
rect 859 3341 860 3345
rect 854 3340 860 3341
rect 110 3332 116 3333
rect 110 3328 111 3332
rect 115 3328 116 3332
rect 110 3327 116 3328
rect 110 3315 116 3316
rect 110 3311 111 3315
rect 115 3311 116 3315
rect 110 3310 116 3311
rect 618 3315 624 3316
rect 618 3311 619 3315
rect 623 3311 624 3315
rect 618 3310 624 3311
rect 112 3291 114 3310
rect 198 3305 204 3306
rect 198 3301 199 3305
rect 203 3301 204 3305
rect 198 3300 204 3301
rect 358 3305 364 3306
rect 358 3301 359 3305
rect 363 3301 364 3305
rect 358 3300 364 3301
rect 526 3305 532 3306
rect 526 3301 527 3305
rect 531 3301 532 3305
rect 526 3300 532 3301
rect 200 3291 202 3300
rect 360 3291 362 3300
rect 528 3291 530 3300
rect 111 3290 115 3291
rect 111 3285 115 3286
rect 199 3290 203 3291
rect 199 3285 203 3286
rect 255 3290 259 3291
rect 255 3285 259 3286
rect 359 3290 363 3291
rect 359 3285 363 3286
rect 375 3290 379 3291
rect 375 3285 379 3286
rect 511 3290 515 3291
rect 511 3285 515 3286
rect 527 3290 531 3291
rect 527 3285 531 3286
rect 112 3270 114 3285
rect 256 3280 258 3285
rect 376 3280 378 3285
rect 512 3280 514 3285
rect 254 3279 260 3280
rect 254 3275 255 3279
rect 259 3275 260 3279
rect 254 3274 260 3275
rect 374 3279 380 3280
rect 374 3275 375 3279
rect 379 3275 380 3279
rect 374 3274 380 3275
rect 510 3279 516 3280
rect 510 3275 511 3279
rect 515 3275 516 3279
rect 510 3274 516 3275
rect 110 3269 116 3270
rect 620 3269 622 3310
rect 686 3305 692 3306
rect 686 3301 687 3305
rect 691 3301 692 3305
rect 686 3300 692 3301
rect 846 3305 852 3306
rect 846 3301 847 3305
rect 851 3301 852 3305
rect 846 3300 852 3301
rect 688 3291 690 3300
rect 848 3291 850 3300
rect 663 3290 667 3291
rect 663 3285 667 3286
rect 687 3290 691 3291
rect 687 3285 691 3286
rect 823 3290 827 3291
rect 823 3285 827 3286
rect 847 3290 851 3291
rect 847 3285 851 3286
rect 664 3280 666 3285
rect 824 3280 826 3285
rect 662 3279 668 3280
rect 662 3275 663 3279
rect 667 3275 668 3279
rect 662 3274 668 3275
rect 822 3279 828 3280
rect 822 3275 823 3279
rect 827 3275 828 3279
rect 822 3274 828 3275
rect 952 3272 954 3350
rect 1000 3346 1002 3357
rect 998 3345 1004 3346
rect 998 3341 999 3345
rect 1003 3341 1004 3345
rect 998 3340 1004 3341
rect 1136 3328 1138 3370
rect 1304 3363 1306 3382
rect 1336 3376 1338 3438
rect 1447 3433 1451 3434
rect 1479 3438 1483 3439
rect 1479 3433 1483 3434
rect 1567 3438 1571 3439
rect 1567 3433 1571 3434
rect 1823 3438 1827 3439
rect 1864 3435 1866 3458
rect 1902 3453 1908 3454
rect 1902 3449 1903 3453
rect 1907 3449 1908 3453
rect 1902 3448 1908 3449
rect 2006 3453 2012 3454
rect 2006 3449 2007 3453
rect 2011 3449 2012 3453
rect 2006 3448 2012 3449
rect 2126 3453 2132 3454
rect 2126 3449 2127 3453
rect 2131 3449 2132 3453
rect 2126 3448 2132 3449
rect 1904 3435 1906 3448
rect 2008 3435 2010 3448
rect 2128 3435 2130 3448
rect 1823 3433 1827 3434
rect 1863 3434 1867 3435
rect 1480 3428 1482 3433
rect 1478 3427 1484 3428
rect 1478 3423 1479 3427
rect 1483 3423 1484 3427
rect 1478 3422 1484 3423
rect 1824 3418 1826 3433
rect 1863 3429 1867 3430
rect 1903 3434 1907 3435
rect 1903 3429 1907 3430
rect 1911 3434 1915 3435
rect 1911 3429 1915 3430
rect 2007 3434 2011 3435
rect 2007 3429 2011 3430
rect 2071 3434 2075 3435
rect 2071 3429 2075 3430
rect 2127 3434 2131 3435
rect 2127 3429 2131 3430
rect 1822 3417 1828 3418
rect 1822 3413 1823 3417
rect 1827 3413 1828 3417
rect 1864 3414 1866 3429
rect 1912 3424 1914 3429
rect 2072 3424 2074 3429
rect 1910 3423 1916 3424
rect 1910 3419 1911 3423
rect 1915 3419 1916 3423
rect 1910 3418 1916 3419
rect 2070 3423 2076 3424
rect 2070 3419 2071 3423
rect 2075 3419 2076 3423
rect 2070 3418 2076 3419
rect 2144 3416 2146 3498
rect 2264 3494 2266 3505
rect 2350 3503 2356 3504
rect 2350 3499 2351 3503
rect 2355 3499 2356 3503
rect 2350 3498 2356 3499
rect 2262 3493 2268 3494
rect 2262 3489 2263 3493
rect 2267 3489 2268 3493
rect 2262 3488 2268 3489
rect 2352 3476 2354 3498
rect 2392 3494 2394 3505
rect 2458 3503 2464 3504
rect 2458 3499 2459 3503
rect 2463 3499 2464 3503
rect 2458 3498 2464 3499
rect 2390 3493 2396 3494
rect 2390 3489 2391 3493
rect 2395 3489 2396 3493
rect 2390 3488 2396 3489
rect 2460 3476 2462 3498
rect 2528 3494 2530 3505
rect 2572 3504 2574 3546
rect 2598 3535 2604 3536
rect 2598 3531 2599 3535
rect 2603 3531 2604 3535
rect 2598 3530 2604 3531
rect 2686 3535 2692 3536
rect 2686 3531 2687 3535
rect 2691 3531 2692 3535
rect 2686 3530 2692 3531
rect 2774 3535 2780 3536
rect 2774 3531 2775 3535
rect 2779 3531 2780 3535
rect 2774 3530 2780 3531
rect 2862 3535 2868 3536
rect 2862 3531 2863 3535
rect 2867 3531 2868 3535
rect 2862 3530 2868 3531
rect 2950 3535 2956 3536
rect 2950 3531 2951 3535
rect 2955 3531 2956 3535
rect 2950 3530 2956 3531
rect 3038 3535 3044 3536
rect 3038 3531 3039 3535
rect 3043 3531 3044 3535
rect 3038 3530 3044 3531
rect 3126 3535 3132 3536
rect 3126 3531 3127 3535
rect 3131 3531 3132 3535
rect 3126 3530 3132 3531
rect 3214 3535 3220 3536
rect 3214 3531 3215 3535
rect 3219 3531 3220 3535
rect 3214 3530 3220 3531
rect 2600 3511 2602 3530
rect 2630 3523 2636 3524
rect 2630 3519 2631 3523
rect 2635 3519 2636 3523
rect 2630 3518 2636 3519
rect 2599 3510 2603 3511
rect 2599 3505 2603 3506
rect 2570 3503 2576 3504
rect 2570 3499 2571 3503
rect 2575 3499 2576 3503
rect 2570 3498 2576 3499
rect 2526 3493 2532 3494
rect 2526 3489 2527 3493
rect 2531 3489 2532 3493
rect 2526 3488 2532 3489
rect 2632 3476 2634 3518
rect 2688 3511 2690 3530
rect 2776 3511 2778 3530
rect 2864 3511 2866 3530
rect 2952 3511 2954 3530
rect 3040 3511 3042 3530
rect 3128 3511 3130 3530
rect 3216 3511 3218 3530
rect 2663 3510 2667 3511
rect 2663 3505 2667 3506
rect 2687 3510 2691 3511
rect 2687 3505 2691 3506
rect 2775 3510 2779 3511
rect 2775 3505 2779 3506
rect 2799 3510 2803 3511
rect 2799 3505 2803 3506
rect 2863 3510 2867 3511
rect 2863 3505 2867 3506
rect 2943 3510 2947 3511
rect 2943 3505 2947 3506
rect 2951 3510 2955 3511
rect 2951 3505 2955 3506
rect 3039 3510 3043 3511
rect 3039 3505 3043 3506
rect 3087 3510 3091 3511
rect 3087 3505 3091 3506
rect 3127 3510 3131 3511
rect 3127 3505 3131 3506
rect 3215 3510 3219 3511
rect 3215 3505 3219 3506
rect 2664 3494 2666 3505
rect 2702 3503 2708 3504
rect 2702 3499 2703 3503
rect 2707 3499 2708 3503
rect 2702 3498 2708 3499
rect 2662 3493 2668 3494
rect 2662 3489 2663 3493
rect 2667 3489 2668 3493
rect 2662 3488 2668 3489
rect 2350 3475 2356 3476
rect 2350 3471 2351 3475
rect 2355 3471 2356 3475
rect 2350 3470 2356 3471
rect 2458 3475 2464 3476
rect 2458 3471 2459 3475
rect 2463 3471 2464 3475
rect 2458 3470 2464 3471
rect 2630 3475 2636 3476
rect 2630 3471 2631 3475
rect 2635 3471 2636 3475
rect 2630 3470 2636 3471
rect 2390 3463 2396 3464
rect 2390 3459 2391 3463
rect 2395 3459 2396 3463
rect 2390 3458 2396 3459
rect 2254 3453 2260 3454
rect 2254 3449 2255 3453
rect 2259 3449 2260 3453
rect 2254 3448 2260 3449
rect 2382 3453 2388 3454
rect 2382 3449 2383 3453
rect 2387 3449 2388 3453
rect 2382 3448 2388 3449
rect 2256 3435 2258 3448
rect 2384 3435 2386 3448
rect 2223 3434 2227 3435
rect 2223 3429 2227 3430
rect 2255 3434 2259 3435
rect 2255 3429 2259 3430
rect 2367 3434 2371 3435
rect 2367 3429 2371 3430
rect 2383 3434 2387 3435
rect 2383 3429 2387 3430
rect 2224 3424 2226 3429
rect 2368 3424 2370 3429
rect 2222 3423 2228 3424
rect 2222 3419 2223 3423
rect 2227 3419 2228 3423
rect 2222 3418 2228 3419
rect 2366 3423 2372 3424
rect 2366 3419 2367 3423
rect 2371 3419 2372 3423
rect 2366 3418 2372 3419
rect 2142 3415 2148 3416
rect 1822 3412 1828 3413
rect 1862 3413 1868 3414
rect 1862 3409 1863 3413
rect 1867 3409 1868 3413
rect 2142 3411 2143 3415
rect 2147 3411 2148 3415
rect 2142 3410 2148 3411
rect 1862 3408 1868 3409
rect 1586 3403 1592 3404
rect 1586 3399 1587 3403
rect 1591 3399 1592 3403
rect 1586 3398 1592 3399
rect 1822 3400 1828 3401
rect 1486 3387 1492 3388
rect 1486 3383 1487 3387
rect 1491 3383 1492 3387
rect 1486 3382 1492 3383
rect 1334 3375 1340 3376
rect 1334 3371 1335 3375
rect 1339 3371 1340 3375
rect 1334 3370 1340 3371
rect 1488 3363 1490 3382
rect 1143 3362 1147 3363
rect 1143 3357 1147 3358
rect 1279 3362 1283 3363
rect 1279 3357 1283 3358
rect 1303 3362 1307 3363
rect 1303 3357 1307 3358
rect 1415 3362 1419 3363
rect 1415 3357 1419 3358
rect 1487 3362 1491 3363
rect 1487 3357 1491 3358
rect 1559 3362 1563 3363
rect 1559 3357 1563 3358
rect 1144 3346 1146 3357
rect 1280 3346 1282 3357
rect 1416 3346 1418 3357
rect 1560 3346 1562 3357
rect 1588 3356 1590 3398
rect 1822 3396 1823 3400
rect 1827 3396 1828 3400
rect 2214 3399 2220 3400
rect 1822 3395 1828 3396
rect 1862 3396 1868 3397
rect 1824 3363 1826 3395
rect 1862 3392 1863 3396
rect 1867 3392 1868 3396
rect 2214 3395 2215 3399
rect 2219 3395 2220 3399
rect 2214 3394 2220 3395
rect 2290 3399 2296 3400
rect 2290 3395 2291 3399
rect 2295 3395 2296 3399
rect 2290 3394 2296 3395
rect 1862 3391 1868 3392
rect 1864 3363 1866 3391
rect 1918 3383 1924 3384
rect 1918 3379 1919 3383
rect 1923 3379 1924 3383
rect 1918 3378 1924 3379
rect 2078 3383 2084 3384
rect 2078 3379 2079 3383
rect 2083 3379 2084 3383
rect 2078 3378 2084 3379
rect 1920 3363 1922 3378
rect 1950 3371 1956 3372
rect 1950 3367 1951 3371
rect 1955 3367 1956 3371
rect 1950 3366 1956 3367
rect 1823 3362 1827 3363
rect 1823 3357 1827 3358
rect 1863 3362 1867 3363
rect 1863 3357 1867 3358
rect 1895 3362 1899 3363
rect 1895 3357 1899 3358
rect 1919 3362 1923 3363
rect 1919 3357 1923 3358
rect 1586 3355 1592 3356
rect 1586 3351 1587 3355
rect 1591 3351 1592 3355
rect 1586 3350 1592 3351
rect 1142 3345 1148 3346
rect 1142 3341 1143 3345
rect 1147 3341 1148 3345
rect 1142 3340 1148 3341
rect 1278 3345 1284 3346
rect 1278 3341 1279 3345
rect 1283 3341 1284 3345
rect 1278 3340 1284 3341
rect 1414 3345 1420 3346
rect 1414 3341 1415 3345
rect 1419 3341 1420 3345
rect 1414 3340 1420 3341
rect 1558 3345 1564 3346
rect 1558 3341 1559 3345
rect 1563 3341 1564 3345
rect 1558 3340 1564 3341
rect 1824 3333 1826 3357
rect 1864 3333 1866 3357
rect 1896 3346 1898 3357
rect 1894 3345 1900 3346
rect 1894 3341 1895 3345
rect 1899 3341 1900 3345
rect 1894 3340 1900 3341
rect 1952 3340 1954 3366
rect 2080 3363 2082 3378
rect 2047 3362 2051 3363
rect 2047 3357 2051 3358
rect 2079 3362 2083 3363
rect 2079 3357 2083 3358
rect 2207 3362 2211 3363
rect 2207 3357 2211 3358
rect 1990 3355 1996 3356
rect 1990 3351 1991 3355
rect 1995 3351 1996 3355
rect 1990 3350 1996 3351
rect 1950 3339 1956 3340
rect 1950 3335 1951 3339
rect 1955 3335 1956 3339
rect 1950 3334 1956 3335
rect 1822 3332 1828 3333
rect 1822 3328 1823 3332
rect 1827 3328 1828 3332
rect 1134 3327 1140 3328
rect 1822 3327 1828 3328
rect 1862 3332 1868 3333
rect 1862 3328 1863 3332
rect 1867 3328 1868 3332
rect 1992 3328 1994 3350
rect 2048 3346 2050 3357
rect 2070 3355 2076 3356
rect 2070 3351 2071 3355
rect 2075 3351 2076 3355
rect 2070 3350 2076 3351
rect 2046 3345 2052 3346
rect 2046 3341 2047 3345
rect 2051 3341 2052 3345
rect 2046 3340 2052 3341
rect 1862 3327 1868 3328
rect 1990 3327 1996 3328
rect 1134 3323 1135 3327
rect 1139 3323 1140 3327
rect 1134 3322 1140 3323
rect 1990 3323 1991 3327
rect 1995 3323 1996 3327
rect 1990 3322 1996 3323
rect 1378 3315 1384 3316
rect 1378 3311 1379 3315
rect 1383 3311 1384 3315
rect 1378 3310 1384 3311
rect 1822 3315 1828 3316
rect 1822 3311 1823 3315
rect 1827 3311 1828 3315
rect 1822 3310 1828 3311
rect 1862 3315 1868 3316
rect 1862 3311 1863 3315
rect 1867 3311 1868 3315
rect 1862 3310 1868 3311
rect 990 3305 996 3306
rect 990 3301 991 3305
rect 995 3301 996 3305
rect 990 3300 996 3301
rect 1134 3305 1140 3306
rect 1134 3301 1135 3305
rect 1139 3301 1140 3305
rect 1134 3300 1140 3301
rect 1270 3305 1276 3306
rect 1270 3301 1271 3305
rect 1275 3301 1276 3305
rect 1270 3300 1276 3301
rect 992 3291 994 3300
rect 1136 3291 1138 3300
rect 1272 3291 1274 3300
rect 991 3290 995 3291
rect 991 3285 995 3286
rect 1135 3290 1139 3291
rect 1135 3285 1139 3286
rect 1167 3290 1171 3291
rect 1167 3285 1171 3286
rect 1271 3290 1275 3291
rect 1271 3285 1275 3286
rect 1343 3290 1347 3291
rect 1343 3285 1347 3286
rect 992 3280 994 3285
rect 1168 3280 1170 3285
rect 1344 3280 1346 3285
rect 990 3279 996 3280
rect 990 3275 991 3279
rect 995 3275 996 3279
rect 990 3274 996 3275
rect 1166 3279 1172 3280
rect 1166 3275 1167 3279
rect 1171 3275 1172 3279
rect 1166 3274 1172 3275
rect 1342 3279 1348 3280
rect 1342 3275 1343 3279
rect 1347 3275 1348 3279
rect 1342 3274 1348 3275
rect 738 3271 744 3272
rect 110 3265 111 3269
rect 115 3265 116 3269
rect 110 3264 116 3265
rect 295 3268 299 3269
rect 295 3263 299 3264
rect 619 3268 623 3269
rect 738 3267 739 3271
rect 743 3267 744 3271
rect 738 3266 744 3267
rect 950 3271 956 3272
rect 950 3267 951 3271
rect 955 3267 956 3271
rect 950 3266 956 3267
rect 619 3263 623 3264
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 110 3247 116 3248
rect 112 3219 114 3247
rect 262 3239 268 3240
rect 262 3235 263 3239
rect 267 3235 268 3239
rect 262 3234 268 3235
rect 264 3219 266 3234
rect 296 3228 298 3263
rect 382 3239 388 3240
rect 382 3235 383 3239
rect 387 3235 388 3239
rect 518 3239 524 3240
rect 382 3234 388 3235
rect 463 3236 467 3237
rect 294 3227 300 3228
rect 294 3223 295 3227
rect 299 3223 300 3227
rect 294 3222 300 3223
rect 384 3219 386 3234
rect 518 3235 519 3239
rect 523 3235 524 3239
rect 518 3234 524 3235
rect 670 3239 676 3240
rect 670 3235 671 3239
rect 675 3235 676 3239
rect 740 3237 742 3266
rect 1058 3255 1064 3256
rect 1058 3251 1059 3255
rect 1063 3251 1064 3255
rect 1058 3250 1064 3251
rect 830 3239 836 3240
rect 670 3234 676 3235
rect 739 3236 743 3237
rect 463 3231 467 3232
rect 111 3218 115 3219
rect 111 3213 115 3214
rect 263 3218 267 3219
rect 263 3213 267 3214
rect 383 3218 387 3219
rect 383 3213 387 3214
rect 431 3218 435 3219
rect 431 3213 435 3214
rect 112 3189 114 3213
rect 432 3202 434 3213
rect 464 3212 466 3231
rect 520 3219 522 3234
rect 672 3219 674 3234
rect 830 3235 831 3239
rect 835 3235 836 3239
rect 830 3234 836 3235
rect 998 3239 1004 3240
rect 998 3235 999 3239
rect 1003 3235 1004 3239
rect 998 3234 1004 3235
rect 739 3231 743 3232
rect 832 3219 834 3234
rect 1000 3219 1002 3234
rect 1060 3228 1062 3250
rect 1174 3239 1180 3240
rect 1174 3235 1175 3239
rect 1179 3235 1180 3239
rect 1174 3234 1180 3235
rect 1350 3239 1356 3240
rect 1350 3235 1351 3239
rect 1355 3235 1356 3239
rect 1350 3234 1356 3235
rect 1058 3227 1064 3228
rect 1058 3223 1059 3227
rect 1063 3223 1064 3227
rect 1058 3222 1064 3223
rect 1176 3219 1178 3234
rect 1206 3227 1212 3228
rect 1206 3223 1207 3227
rect 1211 3223 1212 3227
rect 1206 3222 1212 3223
rect 519 3218 523 3219
rect 519 3213 523 3214
rect 551 3218 555 3219
rect 551 3213 555 3214
rect 671 3218 675 3219
rect 671 3213 675 3214
rect 799 3218 803 3219
rect 799 3213 803 3214
rect 831 3218 835 3219
rect 831 3213 835 3214
rect 935 3218 939 3219
rect 935 3213 939 3214
rect 999 3218 1003 3219
rect 999 3213 1003 3214
rect 1079 3218 1083 3219
rect 1079 3213 1083 3214
rect 1175 3218 1179 3219
rect 1175 3213 1179 3214
rect 462 3211 468 3212
rect 462 3207 463 3211
rect 467 3207 468 3211
rect 462 3206 468 3207
rect 552 3202 554 3213
rect 672 3202 674 3213
rect 800 3202 802 3213
rect 936 3202 938 3213
rect 1034 3203 1040 3204
rect 430 3201 436 3202
rect 430 3197 431 3201
rect 435 3197 436 3201
rect 430 3196 436 3197
rect 550 3201 556 3202
rect 550 3197 551 3201
rect 555 3197 556 3201
rect 550 3196 556 3197
rect 670 3201 676 3202
rect 670 3197 671 3201
rect 675 3197 676 3201
rect 670 3196 676 3197
rect 798 3201 804 3202
rect 798 3197 799 3201
rect 803 3197 804 3201
rect 798 3196 804 3197
rect 934 3201 940 3202
rect 934 3197 935 3201
rect 939 3197 940 3201
rect 1034 3199 1035 3203
rect 1039 3199 1040 3203
rect 1080 3202 1082 3213
rect 1034 3198 1040 3199
rect 1078 3201 1084 3202
rect 934 3196 940 3197
rect 110 3188 116 3189
rect 110 3184 111 3188
rect 115 3184 116 3188
rect 110 3183 116 3184
rect 110 3171 116 3172
rect 110 3167 111 3171
rect 115 3167 116 3171
rect 110 3166 116 3167
rect 112 3147 114 3166
rect 422 3161 428 3162
rect 422 3157 423 3161
rect 427 3157 428 3161
rect 422 3156 428 3157
rect 542 3161 548 3162
rect 542 3157 543 3161
rect 547 3157 548 3161
rect 542 3156 548 3157
rect 662 3161 668 3162
rect 662 3157 663 3161
rect 667 3157 668 3161
rect 662 3156 668 3157
rect 790 3161 796 3162
rect 790 3157 791 3161
rect 795 3157 796 3161
rect 790 3156 796 3157
rect 926 3161 932 3162
rect 926 3157 927 3161
rect 931 3157 932 3161
rect 926 3156 932 3157
rect 424 3147 426 3156
rect 502 3155 508 3156
rect 502 3151 503 3155
rect 507 3151 508 3155
rect 502 3150 508 3151
rect 111 3146 115 3147
rect 111 3141 115 3142
rect 423 3146 427 3147
rect 423 3141 427 3142
rect 463 3146 467 3147
rect 463 3141 467 3142
rect 112 3126 114 3141
rect 464 3136 466 3141
rect 462 3135 468 3136
rect 462 3131 463 3135
rect 467 3131 468 3135
rect 462 3130 468 3131
rect 110 3125 116 3126
rect 110 3121 111 3125
rect 115 3121 116 3125
rect 110 3120 116 3121
rect 110 3108 116 3109
rect 110 3104 111 3108
rect 115 3104 116 3108
rect 110 3103 116 3104
rect 112 3071 114 3103
rect 470 3095 476 3096
rect 470 3091 471 3095
rect 475 3091 476 3095
rect 470 3090 476 3091
rect 472 3071 474 3090
rect 504 3084 506 3150
rect 544 3147 546 3156
rect 664 3147 666 3156
rect 792 3147 794 3156
rect 928 3147 930 3156
rect 543 3146 547 3147
rect 543 3141 547 3142
rect 551 3146 555 3147
rect 551 3141 555 3142
rect 639 3146 643 3147
rect 639 3141 643 3142
rect 663 3146 667 3147
rect 663 3141 667 3142
rect 735 3146 739 3147
rect 735 3141 739 3142
rect 791 3146 795 3147
rect 791 3141 795 3142
rect 847 3146 851 3147
rect 847 3141 851 3142
rect 927 3146 931 3147
rect 927 3141 931 3142
rect 967 3146 971 3147
rect 967 3141 971 3142
rect 552 3136 554 3141
rect 640 3136 642 3141
rect 736 3136 738 3141
rect 848 3136 850 3141
rect 968 3136 970 3141
rect 550 3135 556 3136
rect 550 3131 551 3135
rect 555 3131 556 3135
rect 550 3130 556 3131
rect 638 3135 644 3136
rect 638 3131 639 3135
rect 643 3131 644 3135
rect 638 3130 644 3131
rect 734 3135 740 3136
rect 734 3131 735 3135
rect 739 3131 740 3135
rect 734 3130 740 3131
rect 846 3135 852 3136
rect 846 3131 847 3135
rect 851 3131 852 3135
rect 846 3130 852 3131
rect 966 3135 972 3136
rect 966 3131 967 3135
rect 971 3131 972 3135
rect 966 3130 972 3131
rect 1036 3128 1038 3198
rect 1078 3197 1079 3201
rect 1083 3197 1084 3201
rect 1078 3196 1084 3197
rect 1208 3184 1210 3222
rect 1352 3219 1354 3234
rect 1380 3228 1382 3310
rect 1406 3305 1412 3306
rect 1406 3301 1407 3305
rect 1411 3301 1412 3305
rect 1406 3300 1412 3301
rect 1550 3305 1556 3306
rect 1550 3301 1551 3305
rect 1555 3301 1556 3305
rect 1550 3300 1556 3301
rect 1408 3291 1410 3300
rect 1552 3291 1554 3300
rect 1824 3291 1826 3310
rect 1864 3291 1866 3310
rect 1886 3305 1892 3306
rect 1886 3301 1887 3305
rect 1891 3301 1892 3305
rect 1886 3300 1892 3301
rect 2038 3305 2044 3306
rect 2038 3301 2039 3305
rect 2043 3301 2044 3305
rect 2038 3300 2044 3301
rect 1888 3291 1890 3300
rect 2040 3291 2042 3300
rect 1407 3290 1411 3291
rect 1407 3285 1411 3286
rect 1519 3290 1523 3291
rect 1519 3285 1523 3286
rect 1551 3290 1555 3291
rect 1551 3285 1555 3286
rect 1823 3290 1827 3291
rect 1823 3285 1827 3286
rect 1863 3290 1867 3291
rect 1863 3285 1867 3286
rect 1887 3290 1891 3291
rect 1887 3285 1891 3286
rect 2039 3290 2043 3291
rect 2039 3285 2043 3286
rect 2063 3290 2067 3291
rect 2063 3285 2067 3286
rect 1520 3280 1522 3285
rect 1518 3279 1524 3280
rect 1518 3275 1519 3279
rect 1523 3275 1524 3279
rect 1518 3274 1524 3275
rect 1824 3270 1826 3285
rect 1864 3270 1866 3285
rect 1888 3280 1890 3285
rect 2064 3280 2066 3285
rect 1886 3279 1892 3280
rect 1886 3275 1887 3279
rect 1891 3275 1892 3279
rect 1886 3274 1892 3275
rect 2062 3279 2068 3280
rect 2062 3275 2063 3279
rect 2067 3275 2068 3279
rect 2062 3274 2068 3275
rect 1822 3269 1828 3270
rect 1822 3265 1823 3269
rect 1827 3265 1828 3269
rect 1822 3264 1828 3265
rect 1862 3269 1868 3270
rect 1862 3265 1863 3269
rect 1867 3265 1868 3269
rect 2072 3268 2074 3350
rect 2208 3346 2210 3357
rect 2216 3356 2218 3394
rect 2230 3383 2236 3384
rect 2230 3379 2231 3383
rect 2235 3379 2236 3383
rect 2230 3378 2236 3379
rect 2232 3363 2234 3378
rect 2292 3372 2294 3394
rect 2374 3383 2380 3384
rect 2374 3379 2375 3383
rect 2379 3379 2380 3383
rect 2374 3378 2380 3379
rect 2290 3371 2296 3372
rect 2290 3367 2291 3371
rect 2295 3367 2296 3371
rect 2290 3366 2296 3367
rect 2376 3363 2378 3378
rect 2392 3372 2394 3458
rect 2518 3453 2524 3454
rect 2518 3449 2519 3453
rect 2523 3449 2524 3453
rect 2518 3448 2524 3449
rect 2654 3453 2660 3454
rect 2654 3449 2655 3453
rect 2659 3449 2660 3453
rect 2654 3448 2660 3449
rect 2520 3435 2522 3448
rect 2656 3435 2658 3448
rect 2503 3434 2507 3435
rect 2503 3429 2507 3430
rect 2519 3434 2523 3435
rect 2519 3429 2523 3430
rect 2631 3434 2635 3435
rect 2631 3429 2635 3430
rect 2655 3434 2659 3435
rect 2655 3429 2659 3430
rect 2504 3424 2506 3429
rect 2632 3424 2634 3429
rect 2502 3423 2508 3424
rect 2502 3419 2503 3423
rect 2507 3419 2508 3423
rect 2502 3418 2508 3419
rect 2630 3423 2636 3424
rect 2630 3419 2631 3423
rect 2635 3419 2636 3423
rect 2630 3418 2636 3419
rect 2704 3416 2706 3498
rect 2800 3494 2802 3505
rect 2890 3503 2896 3504
rect 2890 3499 2891 3503
rect 2895 3499 2896 3503
rect 2890 3498 2896 3499
rect 2798 3493 2804 3494
rect 2798 3489 2799 3493
rect 2803 3489 2804 3493
rect 2798 3488 2804 3489
rect 2892 3476 2894 3498
rect 2944 3494 2946 3505
rect 3088 3494 3090 3505
rect 3276 3504 3278 3562
rect 3574 3561 3575 3565
rect 3579 3561 3580 3565
rect 3574 3560 3580 3561
rect 3574 3548 3580 3549
rect 3574 3544 3575 3548
rect 3579 3544 3580 3548
rect 3574 3543 3580 3544
rect 3302 3535 3308 3536
rect 3302 3531 3303 3535
rect 3307 3531 3308 3535
rect 3302 3530 3308 3531
rect 3304 3511 3306 3530
rect 3576 3511 3578 3543
rect 3303 3510 3307 3511
rect 3303 3505 3307 3506
rect 3575 3510 3579 3511
rect 3575 3505 3579 3506
rect 3274 3503 3280 3504
rect 3274 3499 3275 3503
rect 3279 3499 3280 3503
rect 3274 3498 3280 3499
rect 2942 3493 2948 3494
rect 2942 3489 2943 3493
rect 2947 3489 2948 3493
rect 2942 3488 2948 3489
rect 3086 3493 3092 3494
rect 3086 3489 3087 3493
rect 3091 3489 3092 3493
rect 3086 3488 3092 3489
rect 3576 3481 3578 3505
rect 3574 3480 3580 3481
rect 3574 3476 3575 3480
rect 3579 3476 3580 3480
rect 2890 3475 2896 3476
rect 3574 3475 3580 3476
rect 2890 3471 2891 3475
rect 2895 3471 2896 3475
rect 2890 3470 2896 3471
rect 2798 3463 2804 3464
rect 2798 3459 2799 3463
rect 2803 3459 2804 3463
rect 2798 3458 2804 3459
rect 3574 3463 3580 3464
rect 3574 3459 3575 3463
rect 3579 3459 3580 3463
rect 3574 3458 3580 3459
rect 2790 3453 2796 3454
rect 2790 3449 2791 3453
rect 2795 3449 2796 3453
rect 2790 3448 2796 3449
rect 2792 3435 2794 3448
rect 2759 3434 2763 3435
rect 2759 3429 2763 3430
rect 2791 3434 2795 3435
rect 2791 3429 2795 3430
rect 2760 3424 2762 3429
rect 2758 3423 2764 3424
rect 2758 3419 2759 3423
rect 2763 3419 2764 3423
rect 2758 3418 2764 3419
rect 2702 3415 2708 3416
rect 2702 3411 2703 3415
rect 2707 3411 2708 3415
rect 2702 3410 2708 3411
rect 2510 3383 2516 3384
rect 2510 3379 2511 3383
rect 2515 3379 2516 3383
rect 2510 3378 2516 3379
rect 2638 3383 2644 3384
rect 2638 3379 2639 3383
rect 2643 3379 2644 3383
rect 2638 3378 2644 3379
rect 2766 3383 2772 3384
rect 2766 3379 2767 3383
rect 2771 3379 2772 3383
rect 2766 3378 2772 3379
rect 2390 3371 2396 3372
rect 2390 3367 2391 3371
rect 2395 3367 2396 3371
rect 2390 3366 2396 3367
rect 2512 3363 2514 3378
rect 2602 3371 2608 3372
rect 2602 3367 2603 3371
rect 2607 3367 2608 3371
rect 2602 3366 2608 3367
rect 2231 3362 2235 3363
rect 2231 3357 2235 3358
rect 2367 3362 2371 3363
rect 2367 3357 2371 3358
rect 2375 3362 2379 3363
rect 2375 3357 2379 3358
rect 2511 3362 2515 3363
rect 2511 3357 2515 3358
rect 2535 3362 2539 3363
rect 2535 3357 2539 3358
rect 2214 3355 2220 3356
rect 2214 3351 2215 3355
rect 2219 3351 2220 3355
rect 2214 3350 2220 3351
rect 2368 3346 2370 3357
rect 2536 3346 2538 3357
rect 2206 3345 2212 3346
rect 2206 3341 2207 3345
rect 2211 3341 2212 3345
rect 2206 3340 2212 3341
rect 2366 3345 2372 3346
rect 2366 3341 2367 3345
rect 2371 3341 2372 3345
rect 2366 3340 2372 3341
rect 2534 3345 2540 3346
rect 2534 3341 2535 3345
rect 2539 3341 2540 3345
rect 2534 3340 2540 3341
rect 2604 3328 2606 3366
rect 2640 3363 2642 3378
rect 2768 3363 2770 3378
rect 2800 3372 2802 3458
rect 2934 3453 2940 3454
rect 2934 3449 2935 3453
rect 2939 3449 2940 3453
rect 2934 3448 2940 3449
rect 3078 3453 3084 3454
rect 3078 3449 3079 3453
rect 3083 3449 3084 3453
rect 3078 3448 3084 3449
rect 2936 3435 2938 3448
rect 3080 3435 3082 3448
rect 3576 3435 3578 3458
rect 2887 3434 2891 3435
rect 2887 3429 2891 3430
rect 2935 3434 2939 3435
rect 2935 3429 2939 3430
rect 3023 3434 3027 3435
rect 3023 3429 3027 3430
rect 3079 3434 3083 3435
rect 3079 3429 3083 3430
rect 3575 3434 3579 3435
rect 3575 3429 3579 3430
rect 2888 3424 2890 3429
rect 3024 3424 3026 3429
rect 2886 3423 2892 3424
rect 2886 3419 2887 3423
rect 2891 3419 2892 3423
rect 2886 3418 2892 3419
rect 3022 3423 3028 3424
rect 3022 3419 3023 3423
rect 3027 3419 3028 3423
rect 3022 3418 3028 3419
rect 3576 3414 3578 3429
rect 3574 3413 3580 3414
rect 3574 3409 3575 3413
rect 3579 3409 3580 3413
rect 3574 3408 3580 3409
rect 2842 3399 2848 3400
rect 2842 3395 2843 3399
rect 2847 3395 2848 3399
rect 2842 3394 2848 3395
rect 3090 3399 3096 3400
rect 3090 3395 3091 3399
rect 3095 3395 3096 3399
rect 3090 3394 3096 3395
rect 3574 3396 3580 3397
rect 2844 3372 2846 3394
rect 2894 3383 2900 3384
rect 2894 3379 2895 3383
rect 2899 3379 2900 3383
rect 2894 3378 2900 3379
rect 3030 3383 3036 3384
rect 3030 3379 3031 3383
rect 3035 3379 3036 3383
rect 3030 3378 3036 3379
rect 2798 3371 2804 3372
rect 2798 3367 2799 3371
rect 2803 3367 2804 3371
rect 2798 3366 2804 3367
rect 2842 3371 2848 3372
rect 2842 3367 2843 3371
rect 2847 3367 2848 3371
rect 2842 3366 2848 3367
rect 2896 3363 2898 3378
rect 3032 3363 3034 3378
rect 2639 3362 2643 3363
rect 2639 3357 2643 3358
rect 2703 3362 2707 3363
rect 2703 3357 2707 3358
rect 2767 3362 2771 3363
rect 2767 3357 2771 3358
rect 2879 3362 2883 3363
rect 2879 3357 2883 3358
rect 2895 3362 2899 3363
rect 2895 3357 2899 3358
rect 3031 3362 3035 3363
rect 3031 3357 3035 3358
rect 3055 3362 3059 3363
rect 3055 3357 3059 3358
rect 2704 3346 2706 3357
rect 2710 3355 2716 3356
rect 2710 3351 2711 3355
rect 2715 3351 2716 3355
rect 2710 3350 2716 3351
rect 2702 3345 2708 3346
rect 2702 3341 2703 3345
rect 2707 3341 2708 3345
rect 2702 3340 2708 3341
rect 2602 3327 2608 3328
rect 2602 3323 2603 3327
rect 2607 3323 2608 3327
rect 2602 3322 2608 3323
rect 2494 3315 2500 3316
rect 2494 3311 2495 3315
rect 2499 3311 2500 3315
rect 2494 3310 2500 3311
rect 2198 3305 2204 3306
rect 2198 3301 2199 3305
rect 2203 3301 2204 3305
rect 2198 3300 2204 3301
rect 2358 3305 2364 3306
rect 2358 3301 2359 3305
rect 2363 3301 2364 3305
rect 2358 3300 2364 3301
rect 2200 3291 2202 3300
rect 2360 3291 2362 3300
rect 2199 3290 2203 3291
rect 2199 3285 2203 3286
rect 2263 3290 2267 3291
rect 2263 3285 2267 3286
rect 2359 3290 2363 3291
rect 2359 3285 2363 3286
rect 2455 3290 2459 3291
rect 2455 3285 2459 3286
rect 2264 3280 2266 3285
rect 2456 3280 2458 3285
rect 2262 3279 2268 3280
rect 2262 3275 2263 3279
rect 2267 3275 2268 3279
rect 2262 3274 2268 3275
rect 2454 3279 2460 3280
rect 2454 3275 2455 3279
rect 2459 3275 2460 3279
rect 2454 3274 2460 3275
rect 1862 3264 1868 3265
rect 2070 3267 2076 3268
rect 2070 3263 2071 3267
rect 2075 3263 2076 3267
rect 2070 3262 2076 3263
rect 1586 3255 1592 3256
rect 1586 3251 1587 3255
rect 1591 3251 1592 3255
rect 2330 3255 2336 3256
rect 1586 3250 1592 3251
rect 1822 3252 1828 3253
rect 1526 3239 1532 3240
rect 1526 3235 1527 3239
rect 1531 3235 1532 3239
rect 1526 3234 1532 3235
rect 1378 3227 1384 3228
rect 1378 3223 1379 3227
rect 1383 3223 1384 3227
rect 1378 3222 1384 3223
rect 1528 3219 1530 3234
rect 1231 3218 1235 3219
rect 1231 3213 1235 3214
rect 1351 3218 1355 3219
rect 1351 3213 1355 3214
rect 1383 3218 1387 3219
rect 1383 3213 1387 3214
rect 1527 3218 1531 3219
rect 1527 3213 1531 3214
rect 1535 3218 1539 3219
rect 1535 3213 1539 3214
rect 1232 3202 1234 3213
rect 1384 3202 1386 3213
rect 1536 3202 1538 3213
rect 1588 3212 1590 3250
rect 1822 3248 1823 3252
rect 1827 3248 1828 3252
rect 1822 3247 1828 3248
rect 1862 3252 1868 3253
rect 1862 3248 1863 3252
rect 1867 3248 1868 3252
rect 2330 3251 2331 3255
rect 2335 3251 2336 3255
rect 2330 3250 2336 3251
rect 2338 3255 2344 3256
rect 2338 3251 2339 3255
rect 2343 3251 2344 3255
rect 2338 3250 2344 3251
rect 1862 3247 1868 3248
rect 1824 3219 1826 3247
rect 1864 3223 1866 3247
rect 1894 3239 1900 3240
rect 1894 3235 1895 3239
rect 1899 3235 1900 3239
rect 1894 3234 1900 3235
rect 2070 3239 2076 3240
rect 2070 3235 2071 3239
rect 2075 3235 2076 3239
rect 2070 3234 2076 3235
rect 2270 3239 2276 3240
rect 2270 3235 2271 3239
rect 2275 3235 2276 3239
rect 2270 3234 2276 3235
rect 1896 3223 1898 3234
rect 1954 3227 1960 3228
rect 1954 3223 1955 3227
rect 1959 3223 1960 3227
rect 2072 3223 2074 3234
rect 2272 3223 2274 3234
rect 1863 3222 1867 3223
rect 1823 3218 1827 3219
rect 1863 3217 1867 3218
rect 1895 3222 1899 3223
rect 1954 3222 1960 3223
rect 2071 3222 2075 3223
rect 1895 3217 1899 3218
rect 1823 3213 1827 3214
rect 1586 3211 1592 3212
rect 1586 3207 1587 3211
rect 1591 3207 1592 3211
rect 1586 3206 1592 3207
rect 1230 3201 1236 3202
rect 1230 3197 1231 3201
rect 1235 3197 1236 3201
rect 1230 3196 1236 3197
rect 1382 3201 1388 3202
rect 1382 3197 1383 3201
rect 1387 3197 1388 3201
rect 1382 3196 1388 3197
rect 1534 3201 1540 3202
rect 1534 3197 1535 3201
rect 1539 3197 1540 3201
rect 1534 3196 1540 3197
rect 1824 3189 1826 3213
rect 1864 3193 1866 3217
rect 1896 3206 1898 3217
rect 1894 3205 1900 3206
rect 1894 3201 1895 3205
rect 1899 3201 1900 3205
rect 1894 3200 1900 3201
rect 1862 3192 1868 3193
rect 1956 3192 1958 3222
rect 2071 3217 2075 3218
rect 2087 3222 2091 3223
rect 2087 3217 2091 3218
rect 2271 3222 2275 3223
rect 2271 3217 2275 3218
rect 2303 3222 2307 3223
rect 2303 3217 2307 3218
rect 1962 3215 1968 3216
rect 1962 3211 1963 3215
rect 1967 3211 1968 3215
rect 1962 3210 1968 3211
rect 1822 3188 1828 3189
rect 1822 3184 1823 3188
rect 1827 3184 1828 3188
rect 1862 3188 1863 3192
rect 1867 3188 1868 3192
rect 1862 3187 1868 3188
rect 1954 3191 1960 3192
rect 1954 3187 1955 3191
rect 1959 3187 1960 3191
rect 1964 3188 1966 3210
rect 2088 3206 2090 3217
rect 2146 3215 2152 3216
rect 2146 3211 2147 3215
rect 2151 3211 2152 3215
rect 2146 3210 2152 3211
rect 2086 3205 2092 3206
rect 2086 3201 2087 3205
rect 2091 3201 2092 3205
rect 2086 3200 2092 3201
rect 1954 3186 1960 3187
rect 1962 3187 1968 3188
rect 1206 3183 1212 3184
rect 1822 3183 1828 3184
rect 1962 3183 1963 3187
rect 1967 3183 1968 3187
rect 1206 3179 1207 3183
rect 1211 3179 1212 3183
rect 1962 3182 1968 3183
rect 1206 3178 1212 3179
rect 1862 3175 1868 3176
rect 1822 3171 1828 3172
rect 1822 3167 1823 3171
rect 1827 3167 1828 3171
rect 1862 3171 1863 3175
rect 1867 3171 1868 3175
rect 1862 3170 1868 3171
rect 1822 3166 1828 3167
rect 1070 3161 1076 3162
rect 1070 3157 1071 3161
rect 1075 3157 1076 3161
rect 1070 3156 1076 3157
rect 1222 3161 1228 3162
rect 1222 3157 1223 3161
rect 1227 3157 1228 3161
rect 1222 3156 1228 3157
rect 1374 3161 1380 3162
rect 1374 3157 1375 3161
rect 1379 3157 1380 3161
rect 1374 3156 1380 3157
rect 1526 3161 1532 3162
rect 1526 3157 1527 3161
rect 1531 3157 1532 3161
rect 1526 3156 1532 3157
rect 1072 3147 1074 3156
rect 1224 3147 1226 3156
rect 1376 3147 1378 3156
rect 1414 3155 1420 3156
rect 1414 3151 1415 3155
rect 1419 3151 1420 3155
rect 1414 3150 1420 3151
rect 1071 3146 1075 3147
rect 1071 3141 1075 3142
rect 1095 3146 1099 3147
rect 1095 3141 1099 3142
rect 1223 3146 1227 3147
rect 1223 3141 1227 3142
rect 1231 3146 1235 3147
rect 1231 3141 1235 3142
rect 1375 3146 1379 3147
rect 1375 3141 1379 3142
rect 1096 3136 1098 3141
rect 1232 3136 1234 3141
rect 1376 3136 1378 3141
rect 1094 3135 1100 3136
rect 1094 3131 1095 3135
rect 1099 3131 1100 3135
rect 1094 3130 1100 3131
rect 1230 3135 1236 3136
rect 1230 3131 1231 3135
rect 1235 3131 1236 3135
rect 1230 3130 1236 3131
rect 1374 3135 1380 3136
rect 1374 3131 1375 3135
rect 1379 3131 1380 3135
rect 1374 3130 1380 3131
rect 914 3127 920 3128
rect 914 3123 915 3127
rect 919 3123 920 3127
rect 914 3122 920 3123
rect 1034 3127 1040 3128
rect 1034 3123 1035 3127
rect 1039 3123 1040 3127
rect 1034 3122 1040 3123
rect 558 3095 564 3096
rect 558 3091 559 3095
rect 563 3091 564 3095
rect 558 3090 564 3091
rect 646 3095 652 3096
rect 646 3091 647 3095
rect 651 3091 652 3095
rect 646 3090 652 3091
rect 742 3095 748 3096
rect 742 3091 743 3095
rect 747 3091 748 3095
rect 742 3090 748 3091
rect 854 3095 860 3096
rect 854 3091 855 3095
rect 859 3091 860 3095
rect 854 3090 860 3091
rect 502 3083 508 3084
rect 502 3079 503 3083
rect 507 3079 508 3083
rect 502 3078 508 3079
rect 560 3071 562 3090
rect 648 3071 650 3090
rect 744 3071 746 3090
rect 856 3071 858 3090
rect 111 3070 115 3071
rect 111 3065 115 3066
rect 151 3070 155 3071
rect 151 3065 155 3066
rect 239 3070 243 3071
rect 239 3065 243 3066
rect 327 3070 331 3071
rect 327 3065 331 3066
rect 415 3070 419 3071
rect 415 3065 419 3066
rect 471 3070 475 3071
rect 471 3065 475 3066
rect 503 3070 507 3071
rect 503 3065 507 3066
rect 559 3070 563 3071
rect 559 3065 563 3066
rect 591 3070 595 3071
rect 591 3065 595 3066
rect 647 3070 651 3071
rect 647 3065 651 3066
rect 679 3070 683 3071
rect 679 3065 683 3066
rect 743 3070 747 3071
rect 743 3065 747 3066
rect 767 3070 771 3071
rect 767 3065 771 3066
rect 855 3070 859 3071
rect 855 3065 859 3066
rect 112 3041 114 3065
rect 152 3054 154 3065
rect 222 3063 228 3064
rect 222 3058 223 3063
rect 227 3058 228 3063
rect 230 3063 236 3064
rect 230 3059 231 3063
rect 235 3059 236 3063
rect 230 3058 236 3059
rect 223 3055 227 3056
rect 150 3053 156 3054
rect 150 3049 151 3053
rect 155 3049 156 3053
rect 150 3048 156 3049
rect 110 3040 116 3041
rect 110 3036 111 3040
rect 115 3036 116 3040
rect 232 3036 234 3058
rect 240 3054 242 3065
rect 328 3054 330 3065
rect 416 3054 418 3065
rect 504 3054 506 3065
rect 592 3054 594 3065
rect 680 3054 682 3065
rect 768 3054 770 3065
rect 856 3054 858 3065
rect 916 3061 918 3122
rect 1162 3111 1168 3112
rect 1162 3107 1163 3111
rect 1167 3107 1168 3111
rect 1162 3106 1168 3107
rect 974 3095 980 3096
rect 974 3091 975 3095
rect 979 3091 980 3095
rect 974 3090 980 3091
rect 1102 3095 1108 3096
rect 1102 3091 1103 3095
rect 1107 3091 1108 3095
rect 1102 3090 1108 3091
rect 976 3071 978 3090
rect 1104 3071 1106 3090
rect 1164 3084 1166 3106
rect 1238 3095 1244 3096
rect 1238 3091 1239 3095
rect 1243 3091 1244 3095
rect 1238 3090 1244 3091
rect 1382 3095 1388 3096
rect 1382 3091 1383 3095
rect 1387 3091 1388 3095
rect 1382 3090 1388 3091
rect 1162 3083 1168 3084
rect 1162 3079 1163 3083
rect 1167 3079 1168 3083
rect 1162 3078 1168 3079
rect 1240 3071 1242 3090
rect 1384 3071 1386 3090
rect 1416 3084 1418 3150
rect 1528 3147 1530 3156
rect 1824 3147 1826 3166
rect 1864 3151 1866 3170
rect 1886 3165 1892 3166
rect 1886 3161 1887 3165
rect 1891 3161 1892 3165
rect 1886 3160 1892 3161
rect 2078 3165 2084 3166
rect 2078 3161 2079 3165
rect 2083 3161 2084 3165
rect 2078 3160 2084 3161
rect 1888 3151 1890 3160
rect 2080 3151 2082 3160
rect 1863 3150 1867 3151
rect 1519 3146 1523 3147
rect 1519 3141 1523 3142
rect 1527 3146 1531 3147
rect 1527 3141 1531 3142
rect 1823 3146 1827 3147
rect 1863 3145 1867 3146
rect 1887 3150 1891 3151
rect 1887 3145 1891 3146
rect 2079 3150 2083 3151
rect 2079 3145 2083 3146
rect 1823 3141 1827 3142
rect 1520 3136 1522 3141
rect 1518 3135 1524 3136
rect 1518 3131 1519 3135
rect 1523 3131 1524 3135
rect 1518 3130 1524 3131
rect 1824 3126 1826 3141
rect 1864 3130 1866 3145
rect 1888 3140 1890 3145
rect 2080 3140 2082 3145
rect 1886 3139 1892 3140
rect 1886 3135 1887 3139
rect 1891 3135 1892 3139
rect 1886 3134 1892 3135
rect 2078 3139 2084 3140
rect 2078 3135 2079 3139
rect 2083 3135 2084 3139
rect 2078 3134 2084 3135
rect 2148 3132 2150 3210
rect 2304 3206 2306 3217
rect 2332 3216 2334 3250
rect 2340 3228 2342 3250
rect 2462 3239 2468 3240
rect 2462 3235 2463 3239
rect 2467 3235 2468 3239
rect 2462 3234 2468 3235
rect 2338 3227 2344 3228
rect 2338 3223 2339 3227
rect 2343 3223 2344 3227
rect 2464 3223 2466 3234
rect 2496 3228 2498 3310
rect 2526 3305 2532 3306
rect 2526 3301 2527 3305
rect 2531 3301 2532 3305
rect 2526 3300 2532 3301
rect 2694 3305 2700 3306
rect 2694 3301 2695 3305
rect 2699 3301 2700 3305
rect 2694 3300 2700 3301
rect 2528 3291 2530 3300
rect 2696 3291 2698 3300
rect 2527 3290 2531 3291
rect 2527 3285 2531 3286
rect 2639 3290 2643 3291
rect 2639 3285 2643 3286
rect 2695 3290 2699 3291
rect 2695 3285 2699 3286
rect 2640 3280 2642 3285
rect 2638 3279 2644 3280
rect 2638 3275 2639 3279
rect 2643 3275 2644 3279
rect 2638 3274 2644 3275
rect 2712 3272 2714 3350
rect 2880 3346 2882 3357
rect 2986 3355 2992 3356
rect 2986 3351 2987 3355
rect 2991 3351 2992 3355
rect 2986 3350 2992 3351
rect 2878 3345 2884 3346
rect 2878 3341 2879 3345
rect 2883 3341 2884 3345
rect 2878 3340 2884 3341
rect 2988 3328 2990 3350
rect 3056 3346 3058 3357
rect 3092 3356 3094 3394
rect 3574 3392 3575 3396
rect 3579 3392 3580 3396
rect 3574 3391 3580 3392
rect 3576 3363 3578 3391
rect 3575 3362 3579 3363
rect 3575 3357 3579 3358
rect 3086 3355 3094 3356
rect 3086 3351 3087 3355
rect 3091 3352 3094 3355
rect 3091 3351 3092 3352
rect 3086 3350 3092 3351
rect 3054 3345 3060 3346
rect 3054 3341 3055 3345
rect 3059 3341 3060 3345
rect 3054 3340 3060 3341
rect 3576 3333 3578 3357
rect 3574 3332 3580 3333
rect 3574 3328 3575 3332
rect 3579 3328 3580 3332
rect 2986 3327 2992 3328
rect 3574 3327 3580 3328
rect 2986 3323 2987 3327
rect 2991 3323 2992 3327
rect 2986 3322 2992 3323
rect 2854 3315 2860 3316
rect 2854 3311 2855 3315
rect 2859 3311 2860 3315
rect 2854 3310 2860 3311
rect 3574 3315 3580 3316
rect 3574 3311 3575 3315
rect 3579 3311 3580 3315
rect 3574 3310 3580 3311
rect 2815 3290 2819 3291
rect 2815 3285 2819 3286
rect 2816 3280 2818 3285
rect 2814 3279 2820 3280
rect 2814 3275 2815 3279
rect 2819 3275 2820 3279
rect 2814 3274 2820 3275
rect 2710 3271 2716 3272
rect 2710 3267 2711 3271
rect 2715 3267 2716 3271
rect 2710 3266 2716 3267
rect 2646 3239 2652 3240
rect 2646 3235 2647 3239
rect 2651 3235 2652 3239
rect 2646 3234 2652 3235
rect 2822 3239 2828 3240
rect 2822 3235 2823 3239
rect 2827 3235 2828 3239
rect 2822 3234 2828 3235
rect 2494 3227 2500 3228
rect 2494 3223 2495 3227
rect 2499 3223 2500 3227
rect 2648 3223 2650 3234
rect 2678 3227 2684 3228
rect 2678 3223 2679 3227
rect 2683 3223 2684 3227
rect 2824 3223 2826 3234
rect 2856 3228 2858 3310
rect 2870 3305 2876 3306
rect 2870 3301 2871 3305
rect 2875 3301 2876 3305
rect 2870 3300 2876 3301
rect 3046 3305 3052 3306
rect 3046 3301 3047 3305
rect 3051 3301 3052 3305
rect 3046 3300 3052 3301
rect 2872 3291 2874 3300
rect 3048 3291 3050 3300
rect 3576 3291 3578 3310
rect 2871 3290 2875 3291
rect 2871 3285 2875 3286
rect 2983 3290 2987 3291
rect 2983 3285 2987 3286
rect 3047 3290 3051 3291
rect 3047 3285 3051 3286
rect 3151 3290 3155 3291
rect 3151 3285 3155 3286
rect 3319 3290 3323 3291
rect 3319 3285 3323 3286
rect 3479 3290 3483 3291
rect 3479 3285 3483 3286
rect 3575 3290 3579 3291
rect 3575 3285 3579 3286
rect 2984 3280 2986 3285
rect 3152 3280 3154 3285
rect 3320 3280 3322 3285
rect 3480 3280 3482 3285
rect 2982 3279 2988 3280
rect 2982 3275 2983 3279
rect 2987 3275 2988 3279
rect 2982 3274 2988 3275
rect 3150 3279 3156 3280
rect 3150 3275 3151 3279
rect 3155 3275 3156 3279
rect 3150 3274 3156 3275
rect 3318 3279 3324 3280
rect 3318 3275 3319 3279
rect 3323 3275 3324 3279
rect 3318 3274 3324 3275
rect 3478 3279 3484 3280
rect 3478 3275 3479 3279
rect 3483 3275 3484 3279
rect 3478 3274 3484 3275
rect 3576 3270 3578 3285
rect 3574 3269 3580 3270
rect 3574 3265 3575 3269
rect 3579 3265 3580 3269
rect 3574 3264 3580 3265
rect 3062 3255 3068 3256
rect 3062 3251 3063 3255
rect 3067 3251 3068 3255
rect 3062 3250 3068 3251
rect 3070 3255 3076 3256
rect 3070 3251 3071 3255
rect 3075 3251 3076 3255
rect 3070 3250 3076 3251
rect 3546 3255 3552 3256
rect 3546 3251 3547 3255
rect 3551 3251 3552 3255
rect 3546 3250 3552 3251
rect 3574 3252 3580 3253
rect 2990 3239 2996 3240
rect 2990 3235 2991 3239
rect 2995 3235 2996 3239
rect 2990 3234 2996 3235
rect 2854 3227 2860 3228
rect 2854 3223 2855 3227
rect 2859 3223 2860 3227
rect 2992 3223 2994 3234
rect 3064 3228 3066 3250
rect 3062 3227 3068 3228
rect 3062 3223 3063 3227
rect 3067 3223 3068 3227
rect 2338 3222 2344 3223
rect 2463 3222 2467 3223
rect 2494 3222 2500 3223
rect 2511 3222 2515 3223
rect 2463 3217 2467 3218
rect 2511 3217 2515 3218
rect 2647 3222 2651 3223
rect 2678 3222 2684 3223
rect 2703 3222 2707 3223
rect 2647 3217 2651 3218
rect 2330 3215 2336 3216
rect 2330 3211 2331 3215
rect 2335 3211 2336 3215
rect 2330 3210 2336 3211
rect 2512 3206 2514 3217
rect 2302 3205 2308 3206
rect 2302 3201 2303 3205
rect 2307 3201 2308 3205
rect 2302 3200 2308 3201
rect 2510 3205 2516 3206
rect 2510 3201 2511 3205
rect 2515 3201 2516 3205
rect 2510 3200 2516 3201
rect 2680 3188 2682 3222
rect 2703 3217 2707 3218
rect 2823 3222 2827 3223
rect 2854 3222 2860 3223
rect 2879 3222 2883 3223
rect 2823 3217 2827 3218
rect 2879 3217 2883 3218
rect 2991 3222 2995 3223
rect 2991 3217 2995 3218
rect 3039 3222 3043 3223
rect 3062 3222 3068 3223
rect 3039 3217 3043 3218
rect 2704 3206 2706 3217
rect 2762 3215 2768 3216
rect 2762 3211 2763 3215
rect 2767 3211 2768 3215
rect 2762 3210 2768 3211
rect 2702 3205 2708 3206
rect 2702 3201 2703 3205
rect 2707 3201 2708 3205
rect 2702 3200 2708 3201
rect 2678 3187 2684 3188
rect 2678 3183 2679 3187
rect 2683 3183 2684 3187
rect 2678 3182 2684 3183
rect 2294 3165 2300 3166
rect 2294 3161 2295 3165
rect 2299 3161 2300 3165
rect 2294 3160 2300 3161
rect 2502 3165 2508 3166
rect 2502 3161 2503 3165
rect 2507 3161 2508 3165
rect 2502 3160 2508 3161
rect 2694 3165 2700 3166
rect 2694 3161 2695 3165
rect 2699 3161 2700 3165
rect 2694 3160 2700 3161
rect 2296 3151 2298 3160
rect 2504 3151 2506 3160
rect 2542 3159 2548 3160
rect 2542 3155 2543 3159
rect 2547 3155 2548 3159
rect 2542 3154 2548 3155
rect 2295 3150 2299 3151
rect 2295 3145 2299 3146
rect 2503 3150 2507 3151
rect 2503 3145 2507 3146
rect 2296 3140 2298 3145
rect 2504 3140 2506 3145
rect 2294 3139 2300 3140
rect 2294 3135 2295 3139
rect 2299 3135 2300 3139
rect 2294 3134 2300 3135
rect 2502 3139 2508 3140
rect 2502 3135 2503 3139
rect 2507 3135 2508 3139
rect 2502 3134 2508 3135
rect 2146 3131 2152 3132
rect 1862 3129 1868 3130
rect 1822 3125 1828 3126
rect 1822 3121 1823 3125
rect 1827 3121 1828 3125
rect 1862 3125 1863 3129
rect 1867 3125 1868 3129
rect 2146 3127 2147 3131
rect 2151 3127 2152 3131
rect 2146 3126 2152 3127
rect 1862 3124 1868 3125
rect 1822 3120 1828 3121
rect 2286 3115 2292 3116
rect 1862 3112 1868 3113
rect 1586 3111 1592 3112
rect 1586 3107 1587 3111
rect 1591 3107 1592 3111
rect 1586 3106 1592 3107
rect 1822 3108 1828 3109
rect 1526 3095 1532 3096
rect 1526 3091 1527 3095
rect 1531 3091 1532 3095
rect 1526 3090 1532 3091
rect 1414 3083 1420 3084
rect 1414 3079 1415 3083
rect 1419 3079 1420 3083
rect 1414 3078 1420 3079
rect 1528 3071 1530 3090
rect 943 3070 947 3071
rect 943 3065 947 3066
rect 975 3070 979 3071
rect 975 3065 979 3066
rect 1031 3070 1035 3071
rect 1031 3065 1035 3066
rect 1103 3070 1107 3071
rect 1103 3065 1107 3066
rect 1119 3070 1123 3071
rect 1119 3065 1123 3066
rect 1207 3070 1211 3071
rect 1207 3065 1211 3066
rect 1239 3070 1243 3071
rect 1239 3065 1243 3066
rect 1295 3070 1299 3071
rect 1295 3065 1299 3066
rect 1383 3070 1387 3071
rect 1383 3065 1387 3066
rect 1471 3070 1475 3071
rect 1471 3065 1475 3066
rect 1527 3070 1531 3071
rect 1527 3065 1531 3066
rect 1559 3070 1563 3071
rect 1559 3065 1563 3066
rect 915 3060 919 3061
rect 915 3055 919 3056
rect 944 3054 946 3065
rect 1032 3054 1034 3065
rect 1090 3063 1096 3064
rect 1090 3059 1091 3063
rect 1095 3059 1096 3063
rect 1090 3058 1096 3059
rect 238 3053 244 3054
rect 238 3049 239 3053
rect 243 3049 244 3053
rect 238 3048 244 3049
rect 326 3053 332 3054
rect 326 3049 327 3053
rect 331 3049 332 3053
rect 326 3048 332 3049
rect 414 3053 420 3054
rect 414 3049 415 3053
rect 419 3049 420 3053
rect 414 3048 420 3049
rect 502 3053 508 3054
rect 502 3049 503 3053
rect 507 3049 508 3053
rect 502 3048 508 3049
rect 590 3053 596 3054
rect 590 3049 591 3053
rect 595 3049 596 3053
rect 590 3048 596 3049
rect 678 3053 684 3054
rect 678 3049 679 3053
rect 683 3049 684 3053
rect 678 3048 684 3049
rect 766 3053 772 3054
rect 766 3049 767 3053
rect 771 3049 772 3053
rect 766 3048 772 3049
rect 854 3053 860 3054
rect 854 3049 855 3053
rect 859 3049 860 3053
rect 854 3048 860 3049
rect 942 3053 948 3054
rect 942 3049 943 3053
rect 947 3049 948 3053
rect 942 3048 948 3049
rect 1030 3053 1036 3054
rect 1030 3049 1031 3053
rect 1035 3049 1036 3053
rect 1030 3048 1036 3049
rect 1092 3040 1094 3058
rect 1120 3054 1122 3065
rect 1208 3054 1210 3065
rect 1296 3054 1298 3065
rect 1384 3054 1386 3065
rect 1472 3054 1474 3065
rect 1538 3063 1544 3064
rect 1538 3059 1539 3063
rect 1543 3059 1544 3063
rect 1538 3058 1544 3059
rect 1118 3053 1124 3054
rect 1118 3049 1119 3053
rect 1123 3049 1124 3053
rect 1118 3048 1124 3049
rect 1206 3053 1212 3054
rect 1206 3049 1207 3053
rect 1211 3049 1212 3053
rect 1206 3048 1212 3049
rect 1294 3053 1300 3054
rect 1294 3049 1295 3053
rect 1299 3049 1300 3053
rect 1294 3048 1300 3049
rect 1382 3053 1388 3054
rect 1382 3049 1383 3053
rect 1387 3049 1388 3053
rect 1382 3048 1388 3049
rect 1470 3053 1476 3054
rect 1470 3049 1471 3053
rect 1475 3049 1476 3053
rect 1470 3048 1476 3049
rect 1090 3039 1096 3040
rect 110 3035 116 3036
rect 230 3035 236 3036
rect 230 3031 231 3035
rect 235 3031 236 3035
rect 1090 3035 1091 3039
rect 1095 3035 1096 3039
rect 1540 3036 1542 3058
rect 1560 3054 1562 3065
rect 1588 3064 1590 3106
rect 1822 3104 1823 3108
rect 1827 3104 1828 3108
rect 1862 3108 1863 3112
rect 1867 3108 1868 3112
rect 2286 3111 2287 3115
rect 2291 3111 2292 3115
rect 2286 3110 2292 3111
rect 2362 3115 2368 3116
rect 2362 3111 2363 3115
rect 2367 3111 2368 3115
rect 2362 3110 2368 3111
rect 1862 3107 1868 3108
rect 1822 3103 1828 3104
rect 1824 3071 1826 3103
rect 1864 3071 1866 3107
rect 1894 3099 1900 3100
rect 1894 3095 1895 3099
rect 1899 3095 1900 3099
rect 1894 3094 1900 3095
rect 2086 3099 2092 3100
rect 2086 3095 2087 3099
rect 2091 3095 2092 3099
rect 2086 3094 2092 3095
rect 1896 3071 1898 3094
rect 2088 3071 2090 3094
rect 1647 3070 1651 3071
rect 1647 3065 1651 3066
rect 1735 3070 1739 3071
rect 1735 3065 1739 3066
rect 1823 3070 1827 3071
rect 1823 3065 1827 3066
rect 1863 3070 1867 3071
rect 1863 3065 1867 3066
rect 1895 3070 1899 3071
rect 1895 3065 1899 3066
rect 2087 3070 2091 3071
rect 2087 3065 2091 3066
rect 2255 3070 2259 3071
rect 2255 3065 2259 3066
rect 1586 3063 1592 3064
rect 1586 3059 1587 3063
rect 1591 3059 1592 3063
rect 1586 3058 1592 3059
rect 1648 3054 1650 3065
rect 1698 3063 1704 3064
rect 1698 3059 1699 3063
rect 1703 3059 1704 3063
rect 1698 3058 1704 3059
rect 1558 3053 1564 3054
rect 1558 3049 1559 3053
rect 1563 3049 1564 3053
rect 1558 3048 1564 3049
rect 1646 3053 1652 3054
rect 1646 3049 1647 3053
rect 1651 3049 1652 3053
rect 1646 3048 1652 3049
rect 1090 3034 1096 3035
rect 1538 3035 1544 3036
rect 230 3030 236 3031
rect 1538 3031 1539 3035
rect 1543 3031 1544 3035
rect 1538 3030 1544 3031
rect 110 3023 116 3024
rect 110 3019 111 3023
rect 115 3019 116 3023
rect 110 3018 116 3019
rect 1542 3023 1548 3024
rect 1542 3019 1543 3023
rect 1547 3019 1548 3023
rect 1542 3018 1548 3019
rect 112 2995 114 3018
rect 142 3013 148 3014
rect 142 3009 143 3013
rect 147 3009 148 3013
rect 142 3008 148 3009
rect 230 3013 236 3014
rect 230 3009 231 3013
rect 235 3009 236 3013
rect 230 3008 236 3009
rect 318 3013 324 3014
rect 318 3009 319 3013
rect 323 3009 324 3013
rect 318 3008 324 3009
rect 406 3013 412 3014
rect 406 3009 407 3013
rect 411 3009 412 3013
rect 406 3008 412 3009
rect 494 3013 500 3014
rect 494 3009 495 3013
rect 499 3009 500 3013
rect 494 3008 500 3009
rect 582 3013 588 3014
rect 582 3009 583 3013
rect 587 3009 588 3013
rect 582 3008 588 3009
rect 670 3013 676 3014
rect 670 3009 671 3013
rect 675 3009 676 3013
rect 670 3008 676 3009
rect 758 3013 764 3014
rect 758 3009 759 3013
rect 763 3009 764 3013
rect 758 3008 764 3009
rect 846 3013 852 3014
rect 846 3009 847 3013
rect 851 3009 852 3013
rect 846 3008 852 3009
rect 934 3013 940 3014
rect 934 3009 935 3013
rect 939 3009 940 3013
rect 934 3008 940 3009
rect 1022 3013 1028 3014
rect 1022 3009 1023 3013
rect 1027 3009 1028 3013
rect 1022 3008 1028 3009
rect 1110 3013 1116 3014
rect 1110 3009 1111 3013
rect 1115 3009 1116 3013
rect 1110 3008 1116 3009
rect 1198 3013 1204 3014
rect 1198 3009 1199 3013
rect 1203 3009 1204 3013
rect 1198 3008 1204 3009
rect 1286 3013 1292 3014
rect 1286 3009 1287 3013
rect 1291 3009 1292 3013
rect 1286 3008 1292 3009
rect 1374 3013 1380 3014
rect 1374 3009 1375 3013
rect 1379 3009 1380 3013
rect 1374 3008 1380 3009
rect 1462 3013 1468 3014
rect 1462 3009 1463 3013
rect 1467 3009 1468 3013
rect 1462 3008 1468 3009
rect 144 2995 146 3008
rect 232 2995 234 3008
rect 320 2995 322 3008
rect 408 2995 410 3008
rect 496 2995 498 3008
rect 584 2995 586 3008
rect 672 2995 674 3008
rect 760 2995 762 3008
rect 848 2995 850 3008
rect 936 2995 938 3008
rect 1024 2995 1026 3008
rect 1112 2995 1114 3008
rect 1200 2995 1202 3008
rect 1288 2995 1290 3008
rect 1376 2995 1378 3008
rect 1464 2995 1466 3008
rect 111 2994 115 2995
rect 111 2989 115 2990
rect 143 2994 147 2995
rect 143 2989 147 2990
rect 231 2994 235 2995
rect 231 2989 235 2990
rect 319 2994 323 2995
rect 319 2989 323 2990
rect 407 2994 411 2995
rect 407 2989 411 2990
rect 495 2994 499 2995
rect 495 2989 499 2990
rect 583 2994 587 2995
rect 583 2989 587 2990
rect 671 2994 675 2995
rect 671 2989 675 2990
rect 759 2994 763 2995
rect 759 2989 763 2990
rect 847 2994 851 2995
rect 847 2989 851 2990
rect 935 2994 939 2995
rect 935 2989 939 2990
rect 1023 2994 1027 2995
rect 1023 2989 1027 2990
rect 1111 2994 1115 2995
rect 1111 2989 1115 2990
rect 1199 2994 1203 2995
rect 1199 2989 1203 2990
rect 1287 2994 1291 2995
rect 1287 2989 1291 2990
rect 1375 2994 1379 2995
rect 1375 2989 1379 2990
rect 1407 2994 1411 2995
rect 1407 2989 1411 2990
rect 1463 2994 1467 2995
rect 1463 2989 1467 2990
rect 1519 2994 1523 2995
rect 1519 2989 1523 2990
rect 112 2974 114 2989
rect 1408 2984 1410 2989
rect 1520 2984 1522 2989
rect 1406 2983 1412 2984
rect 1406 2979 1407 2983
rect 1411 2979 1412 2983
rect 1406 2978 1412 2979
rect 1518 2983 1524 2984
rect 1518 2979 1519 2983
rect 1523 2979 1524 2983
rect 1518 2978 1524 2979
rect 110 2973 116 2974
rect 110 2969 111 2973
rect 115 2969 116 2973
rect 110 2968 116 2969
rect 1478 2959 1484 2960
rect 110 2956 116 2957
rect 110 2952 111 2956
rect 115 2952 116 2956
rect 1478 2955 1479 2959
rect 1483 2955 1484 2959
rect 1478 2954 1484 2955
rect 110 2951 116 2952
rect 112 2927 114 2951
rect 1414 2943 1420 2944
rect 1414 2939 1415 2943
rect 1419 2939 1420 2943
rect 1414 2938 1420 2939
rect 1416 2927 1418 2938
rect 1480 2932 1482 2954
rect 1498 2951 1504 2952
rect 1498 2947 1499 2951
rect 1503 2947 1504 2951
rect 1498 2946 1504 2947
rect 1478 2931 1484 2932
rect 1478 2927 1479 2931
rect 1483 2927 1484 2931
rect 111 2926 115 2927
rect 111 2921 115 2922
rect 1359 2926 1363 2927
rect 1359 2921 1363 2922
rect 1415 2926 1419 2927
rect 1415 2921 1419 2922
rect 1471 2926 1475 2927
rect 1478 2926 1484 2927
rect 1471 2921 1475 2922
rect 112 2897 114 2921
rect 1360 2910 1362 2921
rect 1472 2910 1474 2921
rect 1500 2920 1502 2946
rect 1526 2943 1532 2944
rect 1526 2939 1527 2943
rect 1531 2939 1532 2943
rect 1526 2938 1532 2939
rect 1528 2927 1530 2938
rect 1544 2932 1546 3018
rect 1550 3013 1556 3014
rect 1550 3009 1551 3013
rect 1555 3009 1556 3013
rect 1550 3008 1556 3009
rect 1638 3013 1644 3014
rect 1638 3009 1639 3013
rect 1643 3009 1644 3013
rect 1638 3008 1644 3009
rect 1552 2995 1554 3008
rect 1640 2995 1642 3008
rect 1551 2994 1555 2995
rect 1551 2989 1555 2990
rect 1631 2994 1635 2995
rect 1631 2989 1635 2990
rect 1639 2994 1643 2995
rect 1639 2989 1643 2990
rect 1632 2984 1634 2989
rect 1630 2983 1636 2984
rect 1630 2979 1631 2983
rect 1635 2979 1636 2983
rect 1630 2978 1636 2979
rect 1700 2976 1702 3058
rect 1736 3054 1738 3065
rect 1734 3053 1740 3054
rect 1734 3049 1735 3053
rect 1739 3049 1740 3053
rect 1734 3048 1740 3049
rect 1824 3041 1826 3065
rect 1864 3041 1866 3065
rect 2256 3054 2258 3065
rect 2288 3064 2290 3110
rect 2302 3099 2308 3100
rect 2302 3095 2303 3099
rect 2307 3095 2308 3099
rect 2302 3094 2308 3095
rect 2304 3071 2306 3094
rect 2364 3088 2366 3110
rect 2510 3099 2516 3100
rect 2510 3095 2511 3099
rect 2515 3095 2516 3099
rect 2510 3094 2516 3095
rect 2362 3087 2368 3088
rect 2362 3083 2363 3087
rect 2367 3083 2368 3087
rect 2362 3082 2368 3083
rect 2512 3071 2514 3094
rect 2544 3088 2546 3154
rect 2696 3151 2698 3160
rect 2695 3150 2699 3151
rect 2695 3145 2699 3146
rect 2696 3140 2698 3145
rect 2694 3139 2700 3140
rect 2694 3135 2695 3139
rect 2699 3135 2700 3139
rect 2694 3134 2700 3135
rect 2764 3132 2766 3210
rect 2880 3206 2882 3217
rect 2978 3215 2984 3216
rect 2978 3211 2979 3215
rect 2983 3211 2984 3215
rect 2978 3210 2984 3211
rect 2878 3205 2884 3206
rect 2878 3201 2879 3205
rect 2883 3201 2884 3205
rect 2878 3200 2884 3201
rect 2980 3188 2982 3210
rect 3040 3206 3042 3217
rect 3072 3216 3074 3250
rect 3158 3239 3164 3240
rect 3158 3235 3159 3239
rect 3163 3235 3164 3239
rect 3158 3234 3164 3235
rect 3326 3239 3332 3240
rect 3326 3235 3327 3239
rect 3331 3235 3332 3239
rect 3326 3234 3332 3235
rect 3486 3239 3492 3240
rect 3486 3235 3487 3239
rect 3491 3235 3492 3239
rect 3486 3234 3492 3235
rect 3160 3223 3162 3234
rect 3328 3223 3330 3234
rect 3488 3223 3490 3234
rect 3159 3222 3163 3223
rect 3159 3217 3163 3218
rect 3199 3222 3203 3223
rect 3199 3217 3203 3218
rect 3327 3222 3331 3223
rect 3327 3217 3331 3218
rect 3351 3222 3355 3223
rect 3351 3217 3355 3218
rect 3487 3222 3491 3223
rect 3487 3217 3491 3218
rect 3070 3215 3076 3216
rect 3070 3211 3071 3215
rect 3075 3211 3076 3215
rect 3070 3210 3076 3211
rect 3200 3206 3202 3217
rect 3352 3206 3354 3217
rect 3410 3215 3416 3216
rect 3410 3211 3411 3215
rect 3415 3211 3416 3215
rect 3410 3210 3416 3211
rect 3038 3205 3044 3206
rect 3038 3201 3039 3205
rect 3043 3201 3044 3205
rect 3038 3200 3044 3201
rect 3198 3205 3204 3206
rect 3198 3201 3199 3205
rect 3203 3201 3204 3205
rect 3198 3200 3204 3201
rect 3350 3205 3356 3206
rect 3350 3201 3351 3205
rect 3355 3201 3356 3205
rect 3350 3200 3356 3201
rect 2978 3187 2984 3188
rect 2978 3183 2979 3187
rect 2983 3183 2984 3187
rect 2978 3182 2984 3183
rect 2870 3165 2876 3166
rect 2870 3161 2871 3165
rect 2875 3161 2876 3165
rect 2870 3160 2876 3161
rect 3030 3165 3036 3166
rect 3030 3161 3031 3165
rect 3035 3161 3036 3165
rect 3030 3160 3036 3161
rect 3190 3165 3196 3166
rect 3190 3161 3191 3165
rect 3195 3161 3196 3165
rect 3190 3160 3196 3161
rect 3342 3165 3348 3166
rect 3342 3161 3343 3165
rect 3347 3161 3348 3165
rect 3342 3160 3348 3161
rect 2872 3151 2874 3160
rect 2910 3159 2916 3160
rect 2910 3155 2911 3159
rect 2915 3155 2916 3159
rect 2910 3154 2916 3155
rect 2871 3150 2875 3151
rect 2871 3145 2875 3146
rect 2872 3140 2874 3145
rect 2870 3139 2876 3140
rect 2870 3135 2871 3139
rect 2875 3135 2876 3139
rect 2870 3134 2876 3135
rect 2762 3131 2768 3132
rect 2762 3127 2763 3131
rect 2767 3127 2768 3131
rect 2762 3126 2768 3127
rect 2702 3099 2708 3100
rect 2702 3095 2703 3099
rect 2707 3095 2708 3099
rect 2702 3094 2708 3095
rect 2878 3099 2884 3100
rect 2878 3095 2879 3099
rect 2883 3095 2884 3099
rect 2878 3094 2884 3095
rect 2542 3087 2548 3088
rect 2542 3083 2543 3087
rect 2547 3083 2548 3087
rect 2542 3082 2548 3083
rect 2704 3071 2706 3094
rect 2880 3071 2882 3094
rect 2912 3088 2914 3154
rect 3032 3151 3034 3160
rect 3192 3151 3194 3160
rect 3344 3151 3346 3160
rect 3031 3150 3035 3151
rect 3031 3145 3035 3146
rect 3039 3150 3043 3151
rect 3039 3145 3043 3146
rect 3191 3150 3195 3151
rect 3191 3145 3195 3146
rect 3343 3150 3347 3151
rect 3343 3145 3347 3146
rect 3040 3140 3042 3145
rect 3192 3140 3194 3145
rect 3344 3140 3346 3145
rect 3038 3139 3044 3140
rect 3038 3135 3039 3139
rect 3043 3135 3044 3139
rect 3038 3134 3044 3135
rect 3190 3139 3196 3140
rect 3190 3135 3191 3139
rect 3195 3135 3196 3139
rect 3190 3134 3196 3135
rect 3342 3139 3348 3140
rect 3342 3135 3343 3139
rect 3347 3135 3348 3139
rect 3342 3134 3348 3135
rect 3412 3132 3414 3210
rect 3488 3206 3490 3217
rect 3548 3216 3550 3250
rect 3574 3248 3575 3252
rect 3579 3248 3580 3252
rect 3574 3247 3580 3248
rect 3576 3223 3578 3247
rect 3575 3222 3579 3223
rect 3575 3217 3579 3218
rect 3546 3215 3552 3216
rect 3546 3211 3547 3215
rect 3551 3211 3552 3215
rect 3546 3210 3552 3211
rect 3486 3205 3492 3206
rect 3486 3201 3487 3205
rect 3491 3201 3492 3205
rect 3486 3200 3492 3201
rect 3576 3193 3578 3217
rect 3574 3192 3580 3193
rect 3574 3188 3575 3192
rect 3579 3188 3580 3192
rect 3574 3187 3580 3188
rect 3574 3175 3580 3176
rect 3574 3171 3575 3175
rect 3579 3171 3580 3175
rect 3574 3170 3580 3171
rect 3478 3165 3484 3166
rect 3478 3161 3479 3165
rect 3483 3161 3484 3165
rect 3478 3160 3484 3161
rect 3480 3151 3482 3160
rect 3518 3159 3524 3160
rect 3518 3155 3519 3159
rect 3523 3155 3524 3159
rect 3518 3154 3524 3155
rect 3479 3150 3483 3151
rect 3479 3145 3483 3146
rect 3480 3140 3482 3145
rect 3478 3139 3484 3140
rect 3478 3135 3479 3139
rect 3483 3135 3484 3139
rect 3478 3134 3484 3135
rect 3410 3131 3416 3132
rect 3410 3127 3411 3131
rect 3415 3127 3416 3131
rect 3410 3126 3416 3127
rect 3046 3099 3052 3100
rect 3046 3095 3047 3099
rect 3051 3095 3052 3099
rect 3046 3094 3052 3095
rect 3198 3099 3204 3100
rect 3198 3095 3199 3099
rect 3203 3095 3204 3099
rect 3198 3094 3204 3095
rect 3350 3099 3356 3100
rect 3350 3095 3351 3099
rect 3355 3095 3356 3099
rect 3350 3094 3356 3095
rect 3486 3099 3492 3100
rect 3486 3095 3487 3099
rect 3491 3095 3492 3099
rect 3486 3094 3492 3095
rect 2910 3087 2916 3088
rect 2910 3083 2911 3087
rect 2915 3083 2916 3087
rect 2910 3082 2916 3083
rect 3048 3071 3050 3094
rect 3200 3071 3202 3094
rect 3352 3071 3354 3094
rect 3488 3071 3490 3094
rect 3520 3088 3522 3154
rect 3576 3151 3578 3170
rect 3575 3150 3579 3151
rect 3575 3145 3579 3146
rect 3576 3130 3578 3145
rect 3574 3129 3580 3130
rect 3574 3125 3575 3129
rect 3579 3125 3580 3129
rect 3574 3124 3580 3125
rect 3554 3115 3560 3116
rect 3554 3111 3555 3115
rect 3559 3111 3560 3115
rect 3554 3110 3560 3111
rect 3574 3112 3580 3113
rect 3518 3087 3524 3088
rect 3518 3083 3519 3087
rect 3523 3083 3524 3087
rect 3518 3082 3524 3083
rect 2303 3070 2307 3071
rect 2303 3065 2307 3066
rect 2423 3070 2427 3071
rect 2423 3065 2427 3066
rect 2511 3070 2515 3071
rect 2511 3065 2515 3066
rect 2591 3070 2595 3071
rect 2591 3065 2595 3066
rect 2703 3070 2707 3071
rect 2703 3065 2707 3066
rect 2751 3070 2755 3071
rect 2751 3065 2755 3066
rect 2879 3070 2883 3071
rect 2879 3065 2883 3066
rect 2919 3070 2923 3071
rect 2919 3065 2923 3066
rect 3047 3070 3051 3071
rect 3047 3065 3051 3066
rect 3087 3070 3091 3071
rect 3087 3065 3091 3066
rect 3199 3070 3203 3071
rect 3199 3065 3203 3066
rect 3351 3070 3355 3071
rect 3351 3065 3355 3066
rect 3487 3070 3491 3071
rect 3487 3065 3491 3066
rect 2286 3063 2292 3064
rect 2286 3059 2287 3063
rect 2291 3059 2292 3063
rect 2286 3058 2292 3059
rect 2424 3054 2426 3065
rect 2592 3054 2594 3065
rect 2752 3054 2754 3065
rect 2782 3063 2788 3064
rect 2782 3058 2783 3063
rect 2787 3058 2788 3063
rect 2783 3055 2787 3056
rect 2920 3054 2922 3065
rect 2930 3063 2936 3064
rect 2930 3059 2931 3063
rect 2935 3059 2936 3063
rect 2930 3058 2936 3059
rect 3035 3060 3039 3061
rect 2254 3053 2260 3054
rect 2254 3049 2255 3053
rect 2259 3049 2260 3053
rect 2254 3048 2260 3049
rect 2422 3053 2428 3054
rect 2422 3049 2423 3053
rect 2427 3049 2428 3053
rect 2422 3048 2428 3049
rect 2590 3053 2596 3054
rect 2590 3049 2591 3053
rect 2595 3049 2596 3053
rect 2590 3048 2596 3049
rect 2750 3053 2756 3054
rect 2750 3049 2751 3053
rect 2755 3049 2756 3053
rect 2750 3048 2756 3049
rect 2918 3053 2924 3054
rect 2918 3049 2919 3053
rect 2923 3049 2924 3053
rect 2918 3048 2924 3049
rect 1822 3040 1828 3041
rect 1822 3036 1823 3040
rect 1827 3036 1828 3040
rect 1822 3035 1828 3036
rect 1862 3040 1868 3041
rect 1862 3036 1863 3040
rect 1867 3036 1868 3040
rect 1862 3035 1868 3036
rect 1822 3023 1828 3024
rect 1822 3019 1823 3023
rect 1827 3019 1828 3023
rect 1822 3018 1828 3019
rect 1862 3023 1868 3024
rect 1862 3019 1863 3023
rect 1867 3019 1868 3023
rect 1862 3018 1868 3019
rect 2498 3023 2504 3024
rect 2498 3019 2499 3023
rect 2503 3019 2504 3023
rect 2498 3018 2504 3019
rect 1726 3013 1732 3014
rect 1726 3009 1727 3013
rect 1731 3009 1732 3013
rect 1726 3008 1732 3009
rect 1728 2995 1730 3008
rect 1824 2995 1826 3018
rect 1864 2999 1866 3018
rect 2246 3013 2252 3014
rect 2246 3009 2247 3013
rect 2251 3009 2252 3013
rect 2246 3008 2252 3009
rect 2414 3013 2420 3014
rect 2414 3009 2415 3013
rect 2419 3009 2420 3013
rect 2414 3008 2420 3009
rect 2248 2999 2250 3008
rect 2416 2999 2418 3008
rect 1863 2998 1867 2999
rect 1727 2994 1731 2995
rect 1727 2989 1731 2990
rect 1823 2994 1827 2995
rect 1863 2993 1867 2994
rect 2239 2998 2243 2999
rect 2239 2993 2243 2994
rect 2247 2998 2251 2999
rect 2247 2993 2251 2994
rect 2415 2998 2419 2999
rect 2415 2993 2419 2994
rect 2463 2998 2467 2999
rect 2463 2993 2467 2994
rect 1823 2989 1827 2990
rect 1728 2984 1730 2989
rect 1726 2983 1732 2984
rect 1726 2979 1727 2983
rect 1731 2979 1732 2983
rect 1726 2978 1732 2979
rect 1698 2975 1704 2976
rect 1698 2971 1699 2975
rect 1703 2971 1704 2975
rect 1824 2974 1826 2989
rect 1864 2978 1866 2993
rect 2240 2988 2242 2993
rect 2464 2988 2466 2993
rect 2238 2987 2244 2988
rect 2238 2983 2239 2987
rect 2243 2983 2244 2987
rect 2238 2982 2244 2983
rect 2462 2987 2468 2988
rect 2462 2983 2463 2987
rect 2467 2983 2468 2987
rect 2462 2982 2468 2983
rect 1862 2977 1868 2978
rect 1698 2970 1704 2971
rect 1822 2973 1828 2974
rect 1822 2969 1823 2973
rect 1827 2969 1828 2973
rect 1862 2973 1863 2977
rect 1867 2973 1868 2977
rect 1862 2972 1868 2973
rect 1822 2968 1828 2969
rect 2306 2963 2312 2964
rect 1862 2960 1868 2961
rect 1822 2956 1828 2957
rect 1822 2952 1823 2956
rect 1827 2952 1828 2956
rect 1862 2956 1863 2960
rect 1867 2956 1868 2960
rect 2306 2959 2307 2963
rect 2311 2959 2312 2963
rect 2306 2958 2312 2959
rect 2350 2963 2356 2964
rect 2350 2959 2351 2963
rect 2355 2959 2356 2963
rect 2350 2958 2356 2959
rect 1862 2955 1868 2956
rect 1822 2951 1828 2952
rect 1638 2943 1644 2944
rect 1638 2939 1639 2943
rect 1643 2939 1644 2943
rect 1638 2938 1644 2939
rect 1734 2943 1740 2944
rect 1734 2939 1735 2943
rect 1739 2939 1740 2943
rect 1734 2938 1740 2939
rect 1542 2931 1548 2932
rect 1534 2927 1540 2928
rect 1527 2926 1531 2927
rect 1534 2923 1535 2927
rect 1539 2923 1540 2927
rect 1542 2927 1543 2931
rect 1547 2927 1548 2931
rect 1640 2927 1642 2938
rect 1736 2927 1738 2938
rect 1762 2931 1768 2932
rect 1762 2927 1763 2931
rect 1767 2927 1768 2931
rect 1824 2927 1826 2951
rect 1542 2926 1548 2927
rect 1583 2926 1587 2927
rect 1534 2922 1540 2923
rect 1527 2921 1531 2922
rect 1498 2919 1504 2920
rect 1498 2915 1499 2919
rect 1503 2915 1504 2919
rect 1498 2914 1504 2915
rect 1536 2915 1538 2922
rect 1583 2921 1587 2922
rect 1639 2926 1643 2927
rect 1639 2921 1643 2922
rect 1703 2926 1707 2927
rect 1703 2921 1707 2922
rect 1735 2926 1739 2927
rect 1762 2926 1768 2927
rect 1823 2926 1827 2927
rect 1735 2921 1739 2922
rect 1536 2913 1542 2915
rect 1358 2909 1364 2910
rect 1358 2905 1359 2909
rect 1363 2905 1364 2909
rect 1358 2904 1364 2905
rect 1470 2909 1476 2910
rect 1470 2905 1471 2909
rect 1475 2905 1476 2909
rect 1470 2904 1476 2905
rect 110 2896 116 2897
rect 110 2892 111 2896
rect 115 2892 116 2896
rect 110 2891 116 2892
rect 1540 2880 1542 2913
rect 1584 2910 1586 2921
rect 1704 2910 1706 2921
rect 1710 2919 1716 2920
rect 1710 2915 1711 2919
rect 1715 2915 1716 2919
rect 1710 2914 1716 2915
rect 1582 2909 1588 2910
rect 1582 2905 1583 2909
rect 1587 2905 1588 2909
rect 1582 2904 1588 2905
rect 1702 2909 1708 2910
rect 1702 2905 1703 2909
rect 1707 2905 1708 2909
rect 1702 2904 1708 2905
rect 110 2879 116 2880
rect 110 2875 111 2879
rect 115 2875 116 2879
rect 110 2874 116 2875
rect 1538 2879 1544 2880
rect 1538 2875 1539 2879
rect 1543 2875 1544 2879
rect 1538 2874 1544 2875
rect 112 2855 114 2874
rect 1350 2869 1356 2870
rect 1350 2865 1351 2869
rect 1355 2865 1356 2869
rect 1350 2864 1356 2865
rect 1462 2869 1468 2870
rect 1462 2865 1463 2869
rect 1467 2865 1468 2869
rect 1462 2864 1468 2865
rect 1574 2869 1580 2870
rect 1574 2865 1575 2869
rect 1579 2865 1580 2869
rect 1574 2864 1580 2865
rect 1694 2869 1700 2870
rect 1694 2865 1695 2869
rect 1699 2865 1700 2869
rect 1694 2864 1700 2865
rect 1352 2855 1354 2864
rect 1418 2863 1424 2864
rect 1418 2859 1419 2863
rect 1423 2859 1424 2863
rect 1418 2858 1424 2859
rect 111 2854 115 2855
rect 111 2849 115 2850
rect 135 2854 139 2855
rect 135 2849 139 2850
rect 223 2854 227 2855
rect 223 2849 227 2850
rect 311 2854 315 2855
rect 311 2849 315 2850
rect 399 2854 403 2855
rect 399 2849 403 2850
rect 487 2854 491 2855
rect 487 2849 491 2850
rect 599 2854 603 2855
rect 599 2849 603 2850
rect 727 2854 731 2855
rect 727 2849 731 2850
rect 863 2854 867 2855
rect 863 2849 867 2850
rect 999 2854 1003 2855
rect 999 2849 1003 2850
rect 1135 2854 1139 2855
rect 1135 2849 1139 2850
rect 1263 2854 1267 2855
rect 1263 2849 1267 2850
rect 1351 2854 1355 2855
rect 1351 2849 1355 2850
rect 1383 2854 1387 2855
rect 1383 2849 1387 2850
rect 112 2834 114 2849
rect 136 2844 138 2849
rect 224 2844 226 2849
rect 312 2844 314 2849
rect 400 2844 402 2849
rect 488 2844 490 2849
rect 600 2844 602 2849
rect 728 2844 730 2849
rect 864 2844 866 2849
rect 1000 2844 1002 2849
rect 1136 2844 1138 2849
rect 1264 2844 1266 2849
rect 1384 2844 1386 2849
rect 134 2843 140 2844
rect 134 2839 135 2843
rect 139 2839 140 2843
rect 134 2838 140 2839
rect 222 2843 228 2844
rect 222 2839 223 2843
rect 227 2839 228 2843
rect 222 2838 228 2839
rect 310 2843 316 2844
rect 310 2839 311 2843
rect 315 2839 316 2843
rect 310 2838 316 2839
rect 398 2843 404 2844
rect 398 2839 399 2843
rect 403 2839 404 2843
rect 398 2838 404 2839
rect 486 2843 492 2844
rect 486 2839 487 2843
rect 491 2839 492 2843
rect 486 2838 492 2839
rect 598 2843 604 2844
rect 598 2839 599 2843
rect 603 2839 604 2843
rect 598 2838 604 2839
rect 726 2843 732 2844
rect 726 2839 727 2843
rect 731 2839 732 2843
rect 726 2838 732 2839
rect 862 2843 868 2844
rect 862 2839 863 2843
rect 867 2839 868 2843
rect 862 2838 868 2839
rect 998 2843 1004 2844
rect 998 2839 999 2843
rect 1003 2839 1004 2843
rect 998 2838 1004 2839
rect 1134 2843 1140 2844
rect 1134 2839 1135 2843
rect 1139 2839 1140 2843
rect 1134 2838 1140 2839
rect 1262 2843 1268 2844
rect 1262 2839 1263 2843
rect 1267 2839 1268 2843
rect 1262 2838 1268 2839
rect 1382 2843 1388 2844
rect 1382 2839 1383 2843
rect 1387 2839 1388 2843
rect 1382 2838 1388 2839
rect 930 2835 936 2836
rect 110 2833 116 2834
rect 110 2829 111 2833
rect 115 2829 116 2833
rect 930 2831 931 2835
rect 935 2831 936 2835
rect 930 2830 936 2831
rect 110 2828 116 2829
rect 202 2819 208 2820
rect 110 2816 116 2817
rect 110 2812 111 2816
rect 115 2812 116 2816
rect 202 2815 203 2819
rect 207 2815 208 2819
rect 202 2814 208 2815
rect 378 2819 384 2820
rect 378 2815 379 2819
rect 383 2815 384 2819
rect 378 2814 384 2815
rect 466 2819 472 2820
rect 466 2815 467 2819
rect 471 2815 472 2819
rect 466 2814 472 2815
rect 558 2819 564 2820
rect 558 2815 559 2819
rect 563 2815 564 2819
rect 558 2814 564 2815
rect 666 2819 672 2820
rect 666 2815 667 2819
rect 671 2815 672 2819
rect 666 2814 672 2815
rect 110 2811 116 2812
rect 112 2787 114 2811
rect 142 2803 148 2804
rect 142 2799 143 2803
rect 147 2799 148 2803
rect 142 2798 148 2799
rect 144 2787 146 2798
rect 204 2792 206 2814
rect 230 2803 236 2804
rect 230 2799 231 2803
rect 235 2799 236 2803
rect 230 2798 236 2799
rect 318 2803 324 2804
rect 318 2799 319 2803
rect 323 2799 324 2803
rect 318 2798 324 2799
rect 202 2791 208 2792
rect 202 2787 203 2791
rect 207 2787 208 2791
rect 232 2787 234 2798
rect 320 2787 322 2798
rect 380 2792 382 2814
rect 406 2803 412 2804
rect 406 2799 407 2803
rect 411 2799 412 2803
rect 406 2798 412 2799
rect 378 2791 384 2792
rect 378 2787 379 2791
rect 383 2787 384 2791
rect 408 2787 410 2798
rect 468 2792 470 2814
rect 494 2803 500 2804
rect 494 2799 495 2803
rect 499 2799 500 2803
rect 494 2798 500 2799
rect 466 2791 472 2792
rect 466 2787 467 2791
rect 471 2787 472 2791
rect 496 2787 498 2798
rect 560 2792 562 2814
rect 606 2803 612 2804
rect 606 2799 607 2803
rect 611 2799 612 2803
rect 606 2798 612 2799
rect 558 2791 564 2792
rect 558 2787 559 2791
rect 563 2787 564 2791
rect 608 2787 610 2798
rect 668 2792 670 2814
rect 734 2803 740 2804
rect 734 2799 735 2803
rect 739 2799 740 2803
rect 734 2798 740 2799
rect 870 2803 876 2804
rect 870 2799 871 2803
rect 875 2799 876 2803
rect 932 2800 934 2830
rect 1066 2819 1072 2820
rect 1066 2815 1067 2819
rect 1071 2815 1072 2819
rect 1066 2814 1072 2815
rect 1330 2819 1336 2820
rect 1330 2815 1331 2819
rect 1335 2815 1336 2819
rect 1330 2814 1336 2815
rect 1006 2803 1012 2804
rect 870 2798 876 2799
rect 930 2799 936 2800
rect 666 2791 672 2792
rect 666 2787 667 2791
rect 671 2787 672 2791
rect 736 2787 738 2798
rect 872 2787 874 2798
rect 930 2795 931 2799
rect 935 2795 936 2799
rect 1006 2799 1007 2803
rect 1011 2799 1012 2803
rect 1006 2798 1012 2799
rect 930 2794 936 2795
rect 1008 2787 1010 2798
rect 111 2786 115 2787
rect 111 2781 115 2782
rect 143 2786 147 2787
rect 143 2781 147 2782
rect 191 2786 195 2787
rect 202 2786 208 2787
rect 231 2786 235 2787
rect 191 2781 195 2782
rect 231 2781 235 2782
rect 295 2786 299 2787
rect 295 2781 299 2782
rect 319 2786 323 2787
rect 378 2786 384 2787
rect 407 2786 411 2787
rect 319 2781 323 2782
rect 407 2781 411 2782
rect 415 2786 419 2787
rect 466 2786 472 2787
rect 495 2786 499 2787
rect 415 2781 419 2782
rect 495 2781 499 2782
rect 551 2786 555 2787
rect 558 2786 564 2787
rect 607 2786 611 2787
rect 666 2786 672 2787
rect 687 2786 691 2787
rect 551 2781 555 2782
rect 607 2781 611 2782
rect 687 2781 691 2782
rect 735 2786 739 2787
rect 735 2781 739 2782
rect 823 2786 827 2787
rect 823 2781 827 2782
rect 871 2786 875 2787
rect 871 2781 875 2782
rect 959 2786 963 2787
rect 959 2781 963 2782
rect 1007 2786 1011 2787
rect 1007 2781 1011 2782
rect 112 2757 114 2781
rect 192 2770 194 2781
rect 296 2770 298 2781
rect 416 2770 418 2781
rect 552 2770 554 2781
rect 570 2779 576 2780
rect 570 2775 571 2779
rect 575 2775 576 2779
rect 570 2774 576 2775
rect 190 2769 196 2770
rect 190 2765 191 2769
rect 195 2765 196 2769
rect 190 2764 196 2765
rect 294 2769 300 2770
rect 294 2765 295 2769
rect 299 2765 300 2769
rect 294 2764 300 2765
rect 414 2769 420 2770
rect 414 2765 415 2769
rect 419 2765 420 2769
rect 414 2764 420 2765
rect 550 2769 556 2770
rect 550 2765 551 2769
rect 555 2765 556 2769
rect 550 2764 556 2765
rect 110 2756 116 2757
rect 110 2752 111 2756
rect 115 2752 116 2756
rect 110 2751 116 2752
rect 110 2739 116 2740
rect 110 2735 111 2739
rect 115 2735 116 2739
rect 110 2734 116 2735
rect 414 2739 420 2740
rect 414 2735 415 2739
rect 419 2735 420 2739
rect 414 2734 420 2735
rect 112 2711 114 2734
rect 182 2729 188 2730
rect 182 2725 183 2729
rect 187 2725 188 2729
rect 182 2724 188 2725
rect 286 2729 292 2730
rect 286 2725 287 2729
rect 291 2725 292 2729
rect 286 2724 292 2725
rect 406 2729 412 2730
rect 406 2725 407 2729
rect 411 2725 412 2729
rect 406 2724 412 2725
rect 184 2711 186 2724
rect 288 2711 290 2724
rect 408 2711 410 2724
rect 111 2710 115 2711
rect 111 2705 115 2706
rect 167 2710 171 2711
rect 167 2705 171 2706
rect 183 2710 187 2711
rect 183 2705 187 2706
rect 279 2710 283 2711
rect 279 2705 283 2706
rect 287 2710 291 2711
rect 287 2705 291 2706
rect 391 2710 395 2711
rect 391 2705 395 2706
rect 407 2710 411 2711
rect 407 2705 411 2706
rect 112 2690 114 2705
rect 168 2700 170 2705
rect 280 2700 282 2705
rect 392 2700 394 2705
rect 166 2699 172 2700
rect 166 2695 167 2699
rect 171 2695 172 2699
rect 166 2694 172 2695
rect 278 2699 284 2700
rect 278 2695 279 2699
rect 283 2695 284 2699
rect 278 2694 284 2695
rect 390 2699 396 2700
rect 390 2695 391 2699
rect 395 2695 396 2699
rect 390 2694 396 2695
rect 110 2689 116 2690
rect 110 2685 111 2689
rect 115 2685 116 2689
rect 110 2684 116 2685
rect 234 2675 240 2676
rect 110 2672 116 2673
rect 110 2668 111 2672
rect 115 2668 116 2672
rect 234 2671 235 2675
rect 239 2671 240 2675
rect 234 2670 240 2671
rect 346 2675 352 2676
rect 346 2671 347 2675
rect 351 2671 352 2675
rect 346 2670 352 2671
rect 110 2667 116 2668
rect 112 2627 114 2667
rect 174 2659 180 2660
rect 174 2655 175 2659
rect 179 2655 180 2659
rect 174 2654 180 2655
rect 176 2627 178 2654
rect 236 2648 238 2670
rect 250 2667 256 2668
rect 250 2663 251 2667
rect 255 2663 256 2667
rect 250 2662 256 2663
rect 234 2647 240 2648
rect 234 2643 235 2647
rect 239 2643 240 2647
rect 234 2642 240 2643
rect 111 2626 115 2627
rect 111 2621 115 2622
rect 175 2626 179 2627
rect 175 2621 179 2622
rect 223 2626 227 2627
rect 223 2621 227 2622
rect 112 2597 114 2621
rect 224 2610 226 2621
rect 252 2620 254 2662
rect 286 2659 292 2660
rect 286 2655 287 2659
rect 291 2655 292 2659
rect 286 2654 292 2655
rect 288 2627 290 2654
rect 348 2648 350 2670
rect 398 2659 404 2660
rect 398 2655 399 2659
rect 403 2655 404 2659
rect 398 2654 404 2655
rect 346 2647 352 2648
rect 346 2643 347 2647
rect 351 2643 352 2647
rect 346 2642 352 2643
rect 400 2627 402 2654
rect 416 2648 418 2734
rect 542 2729 548 2730
rect 542 2725 543 2729
rect 547 2725 548 2729
rect 542 2724 548 2725
rect 544 2711 546 2724
rect 503 2710 507 2711
rect 503 2705 507 2706
rect 543 2710 547 2711
rect 543 2705 547 2706
rect 504 2700 506 2705
rect 502 2699 508 2700
rect 502 2695 503 2699
rect 507 2695 508 2699
rect 502 2694 508 2695
rect 572 2692 574 2774
rect 688 2770 690 2781
rect 824 2770 826 2781
rect 960 2770 962 2781
rect 1068 2772 1070 2814
rect 1142 2803 1148 2804
rect 1142 2799 1143 2803
rect 1147 2799 1148 2803
rect 1142 2798 1148 2799
rect 1270 2803 1276 2804
rect 1270 2799 1271 2803
rect 1275 2799 1276 2803
rect 1270 2798 1276 2799
rect 1144 2787 1146 2798
rect 1272 2787 1274 2798
rect 1332 2792 1334 2814
rect 1390 2803 1396 2804
rect 1390 2799 1391 2803
rect 1395 2799 1396 2803
rect 1390 2798 1396 2799
rect 1330 2791 1336 2792
rect 1330 2787 1331 2791
rect 1335 2787 1336 2791
rect 1392 2787 1394 2798
rect 1420 2792 1422 2858
rect 1464 2855 1466 2864
rect 1576 2855 1578 2864
rect 1696 2855 1698 2864
rect 1463 2854 1467 2855
rect 1463 2849 1467 2850
rect 1503 2854 1507 2855
rect 1503 2849 1507 2850
rect 1575 2854 1579 2855
rect 1575 2849 1579 2850
rect 1623 2854 1627 2855
rect 1623 2849 1627 2850
rect 1695 2854 1699 2855
rect 1695 2849 1699 2850
rect 1504 2844 1506 2849
rect 1624 2844 1626 2849
rect 1502 2843 1508 2844
rect 1502 2839 1503 2843
rect 1507 2839 1508 2843
rect 1502 2838 1508 2839
rect 1622 2843 1628 2844
rect 1622 2839 1623 2843
rect 1627 2839 1628 2843
rect 1622 2838 1628 2839
rect 1712 2836 1714 2914
rect 1764 2896 1766 2926
rect 1823 2921 1827 2922
rect 1824 2897 1826 2921
rect 1864 2915 1866 2955
rect 2246 2947 2252 2948
rect 2246 2943 2247 2947
rect 2251 2943 2252 2947
rect 2246 2942 2252 2943
rect 2248 2915 2250 2942
rect 1863 2914 1867 2915
rect 1863 2909 1867 2910
rect 2239 2914 2243 2915
rect 2239 2909 2243 2910
rect 2247 2914 2251 2915
rect 2247 2909 2251 2910
rect 1822 2896 1828 2897
rect 1762 2895 1768 2896
rect 1762 2891 1763 2895
rect 1767 2891 1768 2895
rect 1822 2892 1823 2896
rect 1827 2892 1828 2896
rect 1822 2891 1828 2892
rect 1762 2890 1768 2891
rect 1864 2885 1866 2909
rect 2240 2898 2242 2909
rect 2308 2908 2310 2958
rect 2352 2936 2354 2958
rect 2470 2947 2476 2948
rect 2470 2943 2471 2947
rect 2475 2943 2476 2947
rect 2470 2942 2476 2943
rect 2350 2935 2356 2936
rect 2350 2931 2351 2935
rect 2355 2931 2356 2935
rect 2350 2930 2356 2931
rect 2472 2915 2474 2942
rect 2500 2936 2502 3018
rect 2582 3013 2588 3014
rect 2582 3009 2583 3013
rect 2587 3009 2588 3013
rect 2582 3008 2588 3009
rect 2742 3013 2748 3014
rect 2742 3009 2743 3013
rect 2747 3009 2748 3013
rect 2742 3008 2748 3009
rect 2910 3013 2916 3014
rect 2910 3009 2911 3013
rect 2915 3009 2916 3013
rect 2910 3008 2916 3009
rect 2584 2999 2586 3008
rect 2744 2999 2746 3008
rect 2912 2999 2914 3008
rect 2583 2998 2587 2999
rect 2583 2993 2587 2994
rect 2671 2998 2675 2999
rect 2671 2993 2675 2994
rect 2743 2998 2747 2999
rect 2743 2993 2747 2994
rect 2863 2998 2867 2999
rect 2863 2993 2867 2994
rect 2911 2998 2915 2999
rect 2911 2993 2915 2994
rect 2672 2988 2674 2993
rect 2864 2988 2866 2993
rect 2670 2987 2676 2988
rect 2670 2983 2671 2987
rect 2675 2983 2676 2987
rect 2670 2982 2676 2983
rect 2862 2987 2868 2988
rect 2862 2983 2863 2987
rect 2867 2983 2868 2987
rect 2862 2982 2868 2983
rect 2932 2980 2934 3058
rect 3035 3055 3039 3056
rect 3036 3036 3038 3055
rect 3088 3054 3090 3065
rect 3086 3053 3092 3054
rect 3086 3049 3087 3053
rect 3091 3049 3092 3053
rect 3086 3048 3092 3049
rect 3034 3035 3040 3036
rect 3034 3031 3035 3035
rect 3039 3031 3040 3035
rect 3034 3030 3040 3031
rect 3078 3013 3084 3014
rect 3078 3009 3079 3013
rect 3083 3009 3084 3013
rect 3078 3008 3084 3009
rect 3080 2999 3082 3008
rect 3031 2998 3035 2999
rect 3031 2993 3035 2994
rect 3079 2998 3083 2999
rect 3079 2993 3083 2994
rect 3191 2998 3195 2999
rect 3191 2993 3195 2994
rect 3343 2998 3347 2999
rect 3343 2993 3347 2994
rect 3479 2998 3483 2999
rect 3479 2993 3483 2994
rect 3032 2988 3034 2993
rect 3192 2988 3194 2993
rect 3344 2988 3346 2993
rect 3480 2988 3482 2993
rect 3030 2987 3036 2988
rect 3030 2983 3031 2987
rect 3035 2983 3036 2987
rect 3030 2982 3036 2983
rect 3190 2987 3196 2988
rect 3190 2983 3191 2987
rect 3195 2983 3196 2987
rect 3190 2982 3196 2983
rect 3342 2987 3348 2988
rect 3342 2983 3343 2987
rect 3347 2983 3348 2987
rect 3342 2982 3348 2983
rect 3478 2987 3484 2988
rect 3478 2983 3479 2987
rect 3483 2983 3484 2987
rect 3478 2982 3484 2983
rect 2930 2979 2936 2980
rect 2930 2975 2931 2979
rect 2935 2975 2936 2979
rect 2930 2974 2936 2975
rect 2958 2963 2964 2964
rect 2958 2959 2959 2963
rect 2963 2959 2964 2963
rect 2958 2958 2964 2959
rect 3098 2963 3104 2964
rect 3098 2959 3099 2963
rect 3103 2959 3104 2963
rect 3098 2958 3104 2959
rect 3258 2963 3264 2964
rect 3258 2959 3259 2963
rect 3263 2959 3264 2963
rect 3258 2958 3264 2959
rect 3546 2963 3552 2964
rect 3546 2959 3547 2963
rect 3551 2959 3552 2963
rect 3546 2958 3552 2959
rect 2678 2947 2684 2948
rect 2678 2943 2679 2947
rect 2683 2943 2684 2947
rect 2678 2942 2684 2943
rect 2870 2947 2876 2948
rect 2870 2943 2871 2947
rect 2875 2943 2876 2947
rect 2870 2942 2876 2943
rect 2498 2935 2504 2936
rect 2498 2931 2499 2935
rect 2503 2931 2504 2935
rect 2498 2930 2504 2931
rect 2680 2915 2682 2942
rect 2711 2940 2715 2941
rect 2710 2935 2716 2936
rect 2710 2931 2711 2935
rect 2715 2931 2716 2935
rect 2710 2930 2716 2931
rect 2872 2915 2874 2942
rect 2960 2941 2962 2958
rect 3038 2947 3044 2948
rect 3038 2943 3039 2947
rect 3043 2943 3044 2947
rect 3038 2942 3044 2943
rect 2959 2940 2963 2941
rect 2959 2935 2963 2936
rect 3040 2915 3042 2942
rect 3100 2936 3102 2958
rect 3198 2947 3204 2948
rect 3198 2943 3199 2947
rect 3203 2943 3204 2947
rect 3198 2942 3204 2943
rect 3098 2935 3104 2936
rect 3098 2931 3099 2935
rect 3103 2931 3104 2935
rect 3098 2930 3104 2931
rect 3200 2915 3202 2942
rect 3260 2936 3262 2958
rect 3350 2947 3356 2948
rect 3350 2943 3351 2947
rect 3355 2943 3356 2947
rect 3350 2942 3356 2943
rect 3486 2947 3492 2948
rect 3486 2943 3487 2947
rect 3491 2943 3492 2947
rect 3486 2942 3492 2943
rect 3258 2935 3264 2936
rect 3258 2931 3259 2935
rect 3263 2931 3264 2935
rect 3258 2930 3264 2931
rect 3352 2915 3354 2942
rect 3394 2935 3400 2936
rect 3394 2931 3395 2935
rect 3399 2931 3400 2935
rect 3394 2930 3400 2931
rect 2463 2914 2467 2915
rect 2463 2909 2467 2910
rect 2471 2914 2475 2915
rect 2471 2909 2475 2910
rect 2671 2914 2675 2915
rect 2671 2909 2675 2910
rect 2679 2914 2683 2915
rect 2679 2909 2683 2910
rect 2855 2914 2859 2915
rect 2855 2909 2859 2910
rect 2871 2914 2875 2915
rect 2871 2909 2875 2910
rect 3023 2914 3027 2915
rect 3023 2909 3027 2910
rect 3039 2914 3043 2915
rect 3039 2909 3043 2910
rect 3183 2914 3187 2915
rect 3183 2909 3187 2910
rect 3199 2914 3203 2915
rect 3199 2909 3203 2910
rect 3335 2914 3339 2915
rect 3335 2909 3339 2910
rect 3351 2914 3355 2915
rect 3351 2909 3355 2910
rect 2306 2907 2312 2908
rect 2306 2903 2307 2907
rect 2311 2903 2312 2907
rect 2306 2902 2312 2903
rect 2394 2907 2400 2908
rect 2394 2903 2395 2907
rect 2399 2903 2400 2907
rect 2394 2902 2400 2903
rect 2238 2897 2244 2898
rect 2238 2893 2239 2897
rect 2243 2893 2244 2897
rect 2238 2892 2244 2893
rect 1862 2884 1868 2885
rect 2396 2884 2398 2902
rect 2464 2898 2466 2909
rect 2672 2898 2674 2909
rect 2750 2907 2756 2908
rect 2750 2903 2751 2907
rect 2755 2903 2756 2907
rect 2750 2902 2756 2903
rect 2462 2897 2468 2898
rect 2462 2893 2463 2897
rect 2467 2893 2468 2897
rect 2462 2892 2468 2893
rect 2670 2897 2676 2898
rect 2670 2893 2671 2897
rect 2675 2893 2676 2897
rect 2670 2892 2676 2893
rect 1862 2880 1863 2884
rect 1867 2880 1868 2884
rect 1822 2879 1828 2880
rect 1862 2879 1868 2880
rect 2394 2883 2400 2884
rect 2394 2879 2395 2883
rect 2399 2879 2400 2883
rect 1822 2875 1823 2879
rect 1827 2875 1828 2879
rect 2394 2878 2400 2879
rect 1822 2874 1828 2875
rect 1824 2855 1826 2874
rect 2752 2869 2754 2902
rect 2856 2898 2858 2909
rect 3024 2898 3026 2909
rect 3184 2898 3186 2909
rect 3336 2898 3338 2909
rect 2854 2897 2860 2898
rect 2854 2893 2855 2897
rect 2859 2893 2860 2897
rect 2854 2892 2860 2893
rect 3022 2897 3028 2898
rect 3022 2893 3023 2897
rect 3027 2893 3028 2897
rect 3022 2892 3028 2893
rect 3182 2897 3188 2898
rect 3182 2893 3183 2897
rect 3187 2893 3188 2897
rect 3182 2892 3188 2893
rect 3334 2897 3340 2898
rect 3334 2893 3335 2897
rect 3339 2893 3340 2897
rect 3334 2892 3340 2893
rect 3396 2884 3398 2930
rect 3488 2915 3490 2942
rect 3487 2914 3491 2915
rect 3487 2909 3491 2910
rect 3488 2898 3490 2909
rect 3548 2908 3550 2958
rect 3556 2936 3558 3110
rect 3574 3108 3575 3112
rect 3579 3108 3580 3112
rect 3574 3107 3580 3108
rect 3576 3071 3578 3107
rect 3575 3070 3579 3071
rect 3575 3065 3579 3066
rect 3576 3041 3578 3065
rect 3574 3040 3580 3041
rect 3574 3036 3575 3040
rect 3579 3036 3580 3040
rect 3574 3035 3580 3036
rect 3574 3023 3580 3024
rect 3574 3019 3575 3023
rect 3579 3019 3580 3023
rect 3574 3018 3580 3019
rect 3576 2999 3578 3018
rect 3575 2998 3579 2999
rect 3575 2993 3579 2994
rect 3576 2978 3578 2993
rect 3574 2977 3580 2978
rect 3574 2973 3575 2977
rect 3579 2973 3580 2977
rect 3574 2972 3580 2973
rect 3574 2960 3580 2961
rect 3574 2956 3575 2960
rect 3579 2956 3580 2960
rect 3574 2955 3580 2956
rect 3554 2935 3560 2936
rect 3554 2931 3555 2935
rect 3559 2931 3560 2935
rect 3554 2930 3560 2931
rect 3576 2915 3578 2955
rect 3575 2914 3579 2915
rect 3575 2909 3579 2910
rect 3546 2907 3552 2908
rect 3546 2903 3547 2907
rect 3551 2903 3552 2907
rect 3546 2902 3552 2903
rect 3486 2897 3492 2898
rect 3486 2893 3487 2897
rect 3491 2893 3492 2897
rect 3486 2892 3492 2893
rect 3576 2885 3578 2909
rect 3574 2884 3580 2885
rect 3394 2883 3400 2884
rect 3394 2879 3395 2883
rect 3399 2879 3400 2883
rect 3574 2880 3575 2884
rect 3579 2880 3580 2884
rect 3574 2879 3580 2880
rect 3394 2878 3400 2879
rect 2751 2868 2755 2869
rect 1862 2867 1868 2868
rect 1862 2863 1863 2867
rect 1867 2863 1868 2867
rect 1862 2862 1868 2863
rect 2546 2867 2552 2868
rect 2546 2863 2547 2867
rect 2551 2863 2552 2867
rect 2751 2863 2755 2864
rect 3099 2868 3103 2869
rect 3099 2863 3103 2864
rect 3574 2867 3580 2868
rect 3574 2863 3575 2867
rect 3579 2863 3580 2867
rect 2546 2862 2552 2863
rect 1727 2854 1731 2855
rect 1727 2849 1731 2850
rect 1823 2854 1827 2855
rect 1823 2849 1827 2850
rect 1728 2844 1730 2849
rect 1726 2843 1732 2844
rect 1726 2839 1727 2843
rect 1731 2839 1732 2843
rect 1726 2838 1732 2839
rect 1710 2835 1716 2836
rect 1710 2831 1711 2835
rect 1715 2831 1716 2835
rect 1824 2834 1826 2849
rect 1864 2843 1866 2862
rect 2230 2857 2236 2858
rect 2230 2853 2231 2857
rect 2235 2853 2236 2857
rect 2230 2852 2236 2853
rect 2454 2857 2460 2858
rect 2454 2853 2455 2857
rect 2459 2853 2460 2857
rect 2454 2852 2460 2853
rect 2232 2843 2234 2852
rect 2456 2843 2458 2852
rect 1863 2842 1867 2843
rect 1863 2837 1867 2838
rect 1895 2842 1899 2843
rect 1895 2837 1899 2838
rect 1983 2842 1987 2843
rect 1983 2837 1987 2838
rect 2071 2842 2075 2843
rect 2071 2837 2075 2838
rect 2159 2842 2163 2843
rect 2159 2837 2163 2838
rect 2231 2842 2235 2843
rect 2231 2837 2235 2838
rect 2247 2842 2251 2843
rect 2247 2837 2251 2838
rect 2335 2842 2339 2843
rect 2335 2837 2339 2838
rect 2423 2842 2427 2843
rect 2423 2837 2427 2838
rect 2455 2842 2459 2843
rect 2455 2837 2459 2838
rect 2511 2842 2515 2843
rect 2511 2837 2515 2838
rect 1710 2830 1716 2831
rect 1822 2833 1828 2834
rect 1822 2829 1823 2833
rect 1827 2829 1828 2833
rect 1822 2828 1828 2829
rect 1864 2822 1866 2837
rect 1896 2832 1898 2837
rect 1984 2832 1986 2837
rect 2072 2832 2074 2837
rect 2160 2832 2162 2837
rect 2248 2832 2250 2837
rect 2336 2832 2338 2837
rect 2424 2832 2426 2837
rect 2512 2832 2514 2837
rect 1894 2831 1900 2832
rect 1894 2827 1895 2831
rect 1899 2827 1900 2831
rect 1894 2826 1900 2827
rect 1982 2831 1988 2832
rect 1982 2827 1983 2831
rect 1987 2827 1988 2831
rect 1982 2826 1988 2827
rect 2070 2831 2076 2832
rect 2070 2827 2071 2831
rect 2075 2827 2076 2831
rect 2070 2826 2076 2827
rect 2158 2831 2164 2832
rect 2158 2827 2159 2831
rect 2163 2827 2164 2831
rect 2158 2826 2164 2827
rect 2246 2831 2252 2832
rect 2246 2827 2247 2831
rect 2251 2827 2252 2831
rect 2246 2826 2252 2827
rect 2334 2831 2340 2832
rect 2334 2827 2335 2831
rect 2339 2827 2340 2831
rect 2334 2826 2340 2827
rect 2422 2831 2428 2832
rect 2422 2827 2423 2831
rect 2427 2827 2428 2831
rect 2422 2826 2428 2827
rect 2510 2831 2516 2832
rect 2510 2827 2511 2831
rect 2515 2827 2516 2831
rect 2510 2826 2516 2827
rect 2498 2823 2504 2824
rect 1862 2821 1868 2822
rect 1578 2819 1584 2820
rect 1578 2815 1579 2819
rect 1583 2815 1584 2819
rect 1578 2814 1584 2815
rect 1690 2819 1696 2820
rect 1690 2815 1691 2819
rect 1695 2815 1696 2819
rect 1862 2817 1863 2821
rect 1867 2817 1868 2821
rect 2498 2819 2499 2823
rect 2503 2819 2504 2823
rect 2498 2818 2504 2819
rect 1690 2814 1696 2815
rect 1822 2816 1828 2817
rect 1862 2816 1868 2817
rect 1510 2803 1516 2804
rect 1510 2799 1511 2803
rect 1515 2799 1516 2803
rect 1510 2798 1516 2799
rect 1418 2791 1424 2792
rect 1418 2787 1419 2791
rect 1423 2787 1424 2791
rect 1512 2787 1514 2798
rect 1580 2792 1582 2814
rect 1630 2803 1636 2804
rect 1630 2799 1631 2803
rect 1635 2799 1636 2803
rect 1692 2800 1694 2814
rect 1822 2812 1823 2816
rect 1827 2812 1828 2816
rect 1822 2811 1828 2812
rect 1734 2803 1740 2804
rect 1630 2798 1636 2799
rect 1690 2799 1696 2800
rect 1578 2791 1584 2792
rect 1578 2787 1579 2791
rect 1583 2787 1584 2791
rect 1632 2787 1634 2798
rect 1690 2795 1691 2799
rect 1695 2795 1696 2799
rect 1734 2799 1735 2803
rect 1739 2799 1740 2803
rect 1734 2798 1740 2799
rect 1690 2794 1696 2795
rect 1736 2787 1738 2798
rect 1794 2791 1800 2792
rect 1794 2787 1795 2791
rect 1799 2787 1800 2791
rect 1824 2787 1826 2811
rect 2490 2807 2496 2808
rect 1862 2804 1868 2805
rect 1862 2800 1863 2804
rect 1867 2800 1868 2804
rect 2490 2803 2491 2807
rect 2495 2803 2496 2807
rect 2490 2802 2496 2803
rect 1862 2799 1868 2800
rect 1087 2786 1091 2787
rect 1087 2781 1091 2782
rect 1143 2786 1147 2787
rect 1143 2781 1147 2782
rect 1207 2786 1211 2787
rect 1207 2781 1211 2782
rect 1271 2786 1275 2787
rect 1271 2781 1275 2782
rect 1319 2786 1323 2787
rect 1330 2786 1336 2787
rect 1391 2786 1395 2787
rect 1418 2786 1424 2787
rect 1431 2786 1435 2787
rect 1319 2781 1323 2782
rect 1391 2781 1395 2782
rect 1431 2781 1435 2782
rect 1511 2786 1515 2787
rect 1511 2781 1515 2782
rect 1535 2786 1539 2787
rect 1578 2786 1584 2787
rect 1631 2786 1635 2787
rect 1535 2781 1539 2782
rect 1631 2781 1635 2782
rect 1647 2786 1651 2787
rect 1647 2781 1651 2782
rect 1735 2786 1739 2787
rect 1794 2786 1800 2787
rect 1823 2786 1827 2787
rect 1735 2781 1739 2782
rect 1066 2771 1072 2772
rect 686 2769 692 2770
rect 686 2765 687 2769
rect 691 2765 692 2769
rect 686 2764 692 2765
rect 822 2769 828 2770
rect 822 2765 823 2769
rect 827 2765 828 2769
rect 822 2764 828 2765
rect 958 2769 964 2770
rect 958 2765 959 2769
rect 963 2765 964 2769
rect 1066 2767 1067 2771
rect 1071 2767 1072 2771
rect 1088 2770 1090 2781
rect 1190 2779 1196 2780
rect 1190 2775 1191 2779
rect 1195 2775 1196 2779
rect 1190 2774 1196 2775
rect 1066 2766 1072 2767
rect 1086 2769 1092 2770
rect 958 2764 964 2765
rect 1086 2765 1087 2769
rect 1091 2765 1092 2769
rect 1086 2764 1092 2765
rect 1192 2756 1194 2774
rect 1208 2770 1210 2781
rect 1320 2770 1322 2781
rect 1432 2770 1434 2781
rect 1536 2770 1538 2781
rect 1648 2770 1650 2781
rect 1736 2770 1738 2781
rect 1206 2769 1212 2770
rect 1206 2765 1207 2769
rect 1211 2765 1212 2769
rect 1206 2764 1212 2765
rect 1318 2769 1324 2770
rect 1318 2765 1319 2769
rect 1323 2765 1324 2769
rect 1318 2764 1324 2765
rect 1430 2769 1436 2770
rect 1430 2765 1431 2769
rect 1435 2765 1436 2769
rect 1430 2764 1436 2765
rect 1534 2769 1540 2770
rect 1534 2765 1535 2769
rect 1539 2765 1540 2769
rect 1534 2764 1540 2765
rect 1646 2769 1652 2770
rect 1646 2765 1647 2769
rect 1651 2765 1652 2769
rect 1646 2764 1652 2765
rect 1734 2769 1740 2770
rect 1734 2765 1735 2769
rect 1739 2765 1740 2769
rect 1734 2764 1740 2765
rect 1796 2756 1798 2786
rect 1823 2781 1827 2782
rect 1824 2757 1826 2781
rect 1864 2763 1866 2799
rect 1902 2791 1908 2792
rect 1902 2787 1903 2791
rect 1907 2787 1908 2791
rect 1902 2786 1908 2787
rect 1990 2791 1996 2792
rect 1990 2787 1991 2791
rect 1995 2787 1996 2791
rect 1990 2786 1996 2787
rect 2078 2791 2084 2792
rect 2078 2787 2079 2791
rect 2083 2787 2084 2791
rect 2078 2786 2084 2787
rect 2166 2791 2172 2792
rect 2166 2787 2167 2791
rect 2171 2787 2172 2791
rect 2166 2786 2172 2787
rect 2254 2791 2260 2792
rect 2254 2787 2255 2791
rect 2259 2787 2260 2791
rect 2254 2786 2260 2787
rect 2342 2791 2348 2792
rect 2342 2787 2343 2791
rect 2347 2787 2348 2791
rect 2342 2786 2348 2787
rect 2430 2791 2436 2792
rect 2430 2787 2431 2791
rect 2435 2787 2436 2791
rect 2430 2786 2436 2787
rect 1904 2763 1906 2786
rect 1992 2763 1994 2786
rect 2080 2763 2082 2786
rect 2168 2763 2170 2786
rect 2256 2763 2258 2786
rect 2344 2763 2346 2786
rect 2432 2763 2434 2786
rect 2492 2780 2494 2802
rect 2490 2779 2496 2780
rect 2490 2775 2491 2779
rect 2495 2775 2496 2779
rect 2490 2774 2496 2775
rect 1863 2762 1867 2763
rect 1863 2757 1867 2758
rect 1903 2762 1907 2763
rect 1903 2757 1907 2758
rect 1991 2762 1995 2763
rect 1991 2757 1995 2758
rect 2047 2762 2051 2763
rect 2047 2757 2051 2758
rect 2079 2762 2083 2763
rect 2079 2757 2083 2758
rect 2167 2762 2171 2763
rect 2167 2757 2171 2758
rect 2255 2762 2259 2763
rect 2255 2757 2259 2758
rect 2295 2762 2299 2763
rect 2295 2757 2299 2758
rect 2343 2762 2347 2763
rect 2343 2757 2347 2758
rect 2431 2762 2435 2763
rect 2431 2757 2435 2758
rect 2447 2762 2451 2763
rect 2447 2757 2451 2758
rect 1822 2756 1828 2757
rect 1190 2755 1196 2756
rect 1190 2751 1191 2755
rect 1195 2751 1196 2755
rect 1190 2750 1196 2751
rect 1794 2755 1800 2756
rect 1794 2751 1795 2755
rect 1799 2751 1800 2755
rect 1822 2752 1823 2756
rect 1827 2752 1828 2756
rect 1822 2751 1828 2752
rect 1794 2750 1800 2751
rect 1822 2739 1828 2740
rect 1822 2735 1823 2739
rect 1827 2735 1828 2739
rect 1822 2734 1828 2735
rect 678 2729 684 2730
rect 678 2725 679 2729
rect 683 2725 684 2729
rect 678 2724 684 2725
rect 814 2729 820 2730
rect 814 2725 815 2729
rect 819 2725 820 2729
rect 814 2724 820 2725
rect 950 2729 956 2730
rect 950 2725 951 2729
rect 955 2725 956 2729
rect 950 2724 956 2725
rect 1078 2729 1084 2730
rect 1078 2725 1079 2729
rect 1083 2725 1084 2729
rect 1078 2724 1084 2725
rect 1198 2729 1204 2730
rect 1198 2725 1199 2729
rect 1203 2725 1204 2729
rect 1198 2724 1204 2725
rect 1310 2729 1316 2730
rect 1310 2725 1311 2729
rect 1315 2725 1316 2729
rect 1310 2724 1316 2725
rect 1422 2729 1428 2730
rect 1422 2725 1423 2729
rect 1427 2725 1428 2729
rect 1422 2724 1428 2725
rect 1526 2729 1532 2730
rect 1526 2725 1527 2729
rect 1531 2725 1532 2729
rect 1526 2724 1532 2725
rect 1638 2729 1644 2730
rect 1638 2725 1639 2729
rect 1643 2725 1644 2729
rect 1638 2724 1644 2725
rect 1726 2729 1732 2730
rect 1726 2725 1727 2729
rect 1731 2725 1732 2729
rect 1726 2724 1732 2725
rect 680 2711 682 2724
rect 816 2711 818 2724
rect 952 2711 954 2724
rect 1080 2711 1082 2724
rect 1200 2711 1202 2724
rect 1312 2711 1314 2724
rect 1424 2711 1426 2724
rect 1528 2711 1530 2724
rect 1640 2711 1642 2724
rect 1728 2711 1730 2724
rect 1824 2711 1826 2734
rect 1864 2733 1866 2757
rect 2022 2755 2028 2756
rect 2022 2751 2023 2755
rect 2027 2751 2028 2755
rect 2022 2750 2028 2751
rect 1862 2732 1868 2733
rect 1862 2728 1863 2732
rect 1867 2728 1868 2732
rect 1862 2727 1868 2728
rect 1862 2715 1868 2716
rect 1862 2711 1863 2715
rect 1867 2711 1868 2715
rect 615 2710 619 2711
rect 615 2705 619 2706
rect 679 2710 683 2711
rect 679 2705 683 2706
rect 815 2710 819 2711
rect 815 2705 819 2706
rect 951 2710 955 2711
rect 951 2705 955 2706
rect 1079 2710 1083 2711
rect 1079 2705 1083 2706
rect 1199 2710 1203 2711
rect 1199 2705 1203 2706
rect 1311 2710 1315 2711
rect 1311 2705 1315 2706
rect 1423 2710 1427 2711
rect 1423 2705 1427 2706
rect 1527 2710 1531 2711
rect 1527 2705 1531 2706
rect 1639 2710 1643 2711
rect 1639 2705 1643 2706
rect 1727 2710 1731 2711
rect 1727 2705 1731 2706
rect 1823 2710 1827 2711
rect 1862 2710 1868 2711
rect 1823 2705 1827 2706
rect 616 2700 618 2705
rect 614 2699 620 2700
rect 614 2695 615 2699
rect 619 2695 620 2699
rect 614 2694 620 2695
rect 570 2691 576 2692
rect 570 2687 571 2691
rect 575 2687 576 2691
rect 1824 2690 1826 2705
rect 1864 2695 1866 2710
rect 1863 2694 1867 2695
rect 570 2686 576 2687
rect 1822 2689 1828 2690
rect 1863 2689 1867 2690
rect 1943 2694 1947 2695
rect 1943 2689 1947 2690
rect 1822 2685 1823 2689
rect 1827 2685 1828 2689
rect 1822 2684 1828 2685
rect 570 2675 576 2676
rect 570 2671 571 2675
rect 575 2671 576 2675
rect 1864 2674 1866 2689
rect 1944 2684 1946 2689
rect 1942 2683 1948 2684
rect 1942 2679 1943 2683
rect 1947 2679 1948 2683
rect 1942 2678 1948 2679
rect 2024 2676 2026 2750
rect 2048 2746 2050 2757
rect 2168 2746 2170 2757
rect 2296 2746 2298 2757
rect 2448 2746 2450 2757
rect 2500 2756 2502 2818
rect 2518 2791 2524 2792
rect 2518 2787 2519 2791
rect 2523 2787 2524 2791
rect 2518 2786 2524 2787
rect 2520 2763 2522 2786
rect 2548 2780 2550 2862
rect 2662 2857 2668 2858
rect 2662 2853 2663 2857
rect 2667 2853 2668 2857
rect 2662 2852 2668 2853
rect 2846 2857 2852 2858
rect 2846 2853 2847 2857
rect 2851 2853 2852 2857
rect 2846 2852 2852 2853
rect 3014 2857 3020 2858
rect 3014 2853 3015 2857
rect 3019 2853 3020 2857
rect 3014 2852 3020 2853
rect 2664 2843 2666 2852
rect 2848 2843 2850 2852
rect 3016 2843 3018 2852
rect 2599 2842 2603 2843
rect 2599 2837 2603 2838
rect 2663 2842 2667 2843
rect 2663 2837 2667 2838
rect 2687 2842 2691 2843
rect 2687 2837 2691 2838
rect 2791 2842 2795 2843
rect 2791 2837 2795 2838
rect 2847 2842 2851 2843
rect 2847 2837 2851 2838
rect 2903 2842 2907 2843
rect 2903 2837 2907 2838
rect 3015 2842 3019 2843
rect 3015 2837 3019 2838
rect 3031 2842 3035 2843
rect 3031 2837 3035 2838
rect 2600 2832 2602 2837
rect 2688 2832 2690 2837
rect 2792 2832 2794 2837
rect 2904 2832 2906 2837
rect 3032 2832 3034 2837
rect 2598 2831 2604 2832
rect 2598 2827 2599 2831
rect 2603 2827 2604 2831
rect 2598 2826 2604 2827
rect 2686 2831 2692 2832
rect 2686 2827 2687 2831
rect 2691 2827 2692 2831
rect 2686 2826 2692 2827
rect 2790 2831 2796 2832
rect 2790 2827 2791 2831
rect 2795 2827 2796 2831
rect 2790 2826 2796 2827
rect 2902 2831 2908 2832
rect 2902 2827 2903 2831
rect 2907 2827 2908 2831
rect 2902 2826 2908 2827
rect 3030 2831 3036 2832
rect 3030 2827 3031 2831
rect 3035 2827 3036 2831
rect 3030 2826 3036 2827
rect 3100 2824 3102 2863
rect 3574 2862 3580 2863
rect 3174 2857 3180 2858
rect 3174 2853 3175 2857
rect 3179 2853 3180 2857
rect 3174 2852 3180 2853
rect 3326 2857 3332 2858
rect 3326 2853 3327 2857
rect 3331 2853 3332 2857
rect 3326 2852 3332 2853
rect 3478 2857 3484 2858
rect 3478 2853 3479 2857
rect 3483 2853 3484 2857
rect 3478 2852 3484 2853
rect 3176 2843 3178 2852
rect 3328 2843 3330 2852
rect 3480 2843 3482 2852
rect 3518 2851 3524 2852
rect 3518 2847 3519 2851
rect 3523 2847 3524 2851
rect 3518 2846 3524 2847
rect 3175 2842 3179 2843
rect 3175 2837 3179 2838
rect 3327 2842 3331 2843
rect 3327 2837 3331 2838
rect 3479 2842 3483 2843
rect 3479 2837 3483 2838
rect 3176 2832 3178 2837
rect 3328 2832 3330 2837
rect 3480 2832 3482 2837
rect 3174 2831 3180 2832
rect 3174 2827 3175 2831
rect 3179 2827 3180 2831
rect 3174 2826 3180 2827
rect 3326 2831 3332 2832
rect 3326 2827 3327 2831
rect 3331 2827 3332 2831
rect 3326 2826 3332 2827
rect 3478 2831 3484 2832
rect 3478 2827 3479 2831
rect 3483 2827 3484 2831
rect 3478 2826 3484 2827
rect 3098 2823 3104 2824
rect 3098 2819 3099 2823
rect 3103 2819 3104 2823
rect 3098 2818 3104 2819
rect 3098 2807 3104 2808
rect 3098 2803 3099 2807
rect 3103 2803 3104 2807
rect 3098 2802 3104 2803
rect 3242 2807 3248 2808
rect 3242 2803 3243 2807
rect 3247 2803 3248 2807
rect 3242 2802 3248 2803
rect 2606 2791 2612 2792
rect 2606 2787 2607 2791
rect 2611 2787 2612 2791
rect 2606 2786 2612 2787
rect 2694 2791 2700 2792
rect 2694 2787 2695 2791
rect 2699 2787 2700 2791
rect 2694 2786 2700 2787
rect 2798 2791 2804 2792
rect 2798 2787 2799 2791
rect 2803 2787 2804 2791
rect 2798 2786 2804 2787
rect 2910 2791 2916 2792
rect 2910 2787 2911 2791
rect 2915 2787 2916 2791
rect 2910 2786 2916 2787
rect 3038 2791 3044 2792
rect 3038 2787 3039 2791
rect 3043 2787 3044 2791
rect 3038 2786 3044 2787
rect 2546 2779 2552 2780
rect 2546 2775 2547 2779
rect 2551 2775 2552 2779
rect 2546 2774 2552 2775
rect 2608 2763 2610 2786
rect 2696 2763 2698 2786
rect 2800 2763 2802 2786
rect 2912 2763 2914 2786
rect 3040 2763 3042 2786
rect 2519 2762 2523 2763
rect 2519 2757 2523 2758
rect 2607 2762 2611 2763
rect 2607 2757 2611 2758
rect 2623 2762 2627 2763
rect 2623 2757 2627 2758
rect 2695 2762 2699 2763
rect 2695 2757 2699 2758
rect 2799 2762 2803 2763
rect 2799 2757 2803 2758
rect 2823 2762 2827 2763
rect 2823 2757 2827 2758
rect 2911 2762 2915 2763
rect 2911 2757 2915 2758
rect 3039 2762 3043 2763
rect 3039 2757 3043 2758
rect 2498 2755 2504 2756
rect 2498 2751 2499 2755
rect 2503 2751 2504 2755
rect 2498 2750 2504 2751
rect 2624 2746 2626 2757
rect 2706 2755 2712 2756
rect 2706 2751 2707 2755
rect 2711 2751 2712 2755
rect 2706 2750 2712 2751
rect 2046 2745 2052 2746
rect 2046 2741 2047 2745
rect 2051 2741 2052 2745
rect 2046 2740 2052 2741
rect 2166 2745 2172 2746
rect 2166 2741 2167 2745
rect 2171 2741 2172 2745
rect 2166 2740 2172 2741
rect 2294 2745 2300 2746
rect 2294 2741 2295 2745
rect 2299 2741 2300 2745
rect 2294 2740 2300 2741
rect 2446 2745 2452 2746
rect 2446 2741 2447 2745
rect 2451 2741 2452 2745
rect 2446 2740 2452 2741
rect 2622 2745 2628 2746
rect 2622 2741 2623 2745
rect 2627 2741 2628 2745
rect 2622 2740 2628 2741
rect 2708 2728 2710 2750
rect 2824 2746 2826 2757
rect 3040 2746 3042 2757
rect 3100 2756 3102 2802
rect 3182 2791 3188 2792
rect 3182 2787 3183 2791
rect 3187 2787 3188 2791
rect 3182 2786 3188 2787
rect 3184 2763 3186 2786
rect 3244 2780 3246 2802
rect 3334 2791 3340 2792
rect 3334 2787 3335 2791
rect 3339 2787 3340 2791
rect 3334 2786 3340 2787
rect 3486 2791 3492 2792
rect 3486 2787 3487 2791
rect 3491 2787 3492 2791
rect 3486 2786 3492 2787
rect 3242 2779 3248 2780
rect 3242 2775 3243 2779
rect 3247 2775 3248 2779
rect 3242 2774 3248 2775
rect 3336 2763 3338 2786
rect 3488 2763 3490 2786
rect 3520 2780 3522 2846
rect 3576 2843 3578 2862
rect 3575 2842 3579 2843
rect 3575 2837 3579 2838
rect 3576 2822 3578 2837
rect 3574 2821 3580 2822
rect 3574 2817 3575 2821
rect 3579 2817 3580 2821
rect 3574 2816 3580 2817
rect 3546 2807 3552 2808
rect 3546 2803 3547 2807
rect 3551 2803 3552 2807
rect 3546 2802 3552 2803
rect 3574 2804 3580 2805
rect 3518 2779 3524 2780
rect 3518 2775 3519 2779
rect 3523 2775 3524 2779
rect 3518 2774 3524 2775
rect 3183 2762 3187 2763
rect 3183 2757 3187 2758
rect 3271 2762 3275 2763
rect 3271 2757 3275 2758
rect 3335 2762 3339 2763
rect 3335 2757 3339 2758
rect 3487 2762 3491 2763
rect 3487 2757 3491 2758
rect 3098 2755 3104 2756
rect 3098 2751 3099 2755
rect 3103 2751 3104 2755
rect 3098 2750 3104 2751
rect 3198 2755 3204 2756
rect 3198 2751 3199 2755
rect 3203 2751 3204 2755
rect 3198 2750 3204 2751
rect 2822 2745 2828 2746
rect 2822 2741 2823 2745
rect 2827 2741 2828 2745
rect 2822 2740 2828 2741
rect 3038 2745 3044 2746
rect 3038 2741 3039 2745
rect 3043 2741 3044 2745
rect 3038 2740 3044 2741
rect 2706 2727 2712 2728
rect 2706 2723 2707 2727
rect 2711 2723 2712 2727
rect 2706 2722 2712 2723
rect 2370 2715 2376 2716
rect 2370 2711 2371 2715
rect 2375 2711 2376 2715
rect 2370 2710 2376 2711
rect 2558 2715 2564 2716
rect 2558 2711 2559 2715
rect 2563 2711 2564 2715
rect 2558 2710 2564 2711
rect 2038 2705 2044 2706
rect 2038 2701 2039 2705
rect 2043 2701 2044 2705
rect 2038 2700 2044 2701
rect 2158 2705 2164 2706
rect 2158 2701 2159 2705
rect 2163 2701 2164 2705
rect 2158 2700 2164 2701
rect 2286 2705 2292 2706
rect 2286 2701 2287 2705
rect 2291 2701 2292 2705
rect 2286 2700 2292 2701
rect 2040 2695 2042 2700
rect 2160 2695 2162 2700
rect 2288 2695 2290 2700
rect 2039 2694 2043 2695
rect 2039 2689 2043 2690
rect 2055 2694 2059 2695
rect 2055 2689 2059 2690
rect 2159 2694 2163 2695
rect 2159 2689 2163 2690
rect 2167 2694 2171 2695
rect 2167 2689 2171 2690
rect 2287 2694 2291 2695
rect 2287 2689 2291 2690
rect 2056 2684 2058 2689
rect 2168 2684 2170 2689
rect 2288 2684 2290 2689
rect 2054 2683 2060 2684
rect 2054 2679 2055 2683
rect 2059 2679 2060 2683
rect 2054 2678 2060 2679
rect 2166 2683 2172 2684
rect 2166 2679 2167 2683
rect 2171 2679 2172 2683
rect 2166 2678 2172 2679
rect 2286 2683 2292 2684
rect 2286 2679 2287 2683
rect 2291 2679 2292 2683
rect 2286 2678 2292 2679
rect 2022 2675 2028 2676
rect 1862 2673 1868 2674
rect 570 2670 576 2671
rect 1822 2672 1828 2673
rect 510 2659 516 2660
rect 510 2655 511 2659
rect 515 2655 516 2659
rect 510 2654 516 2655
rect 414 2647 420 2648
rect 414 2643 415 2647
rect 419 2643 420 2647
rect 414 2642 420 2643
rect 512 2627 514 2654
rect 572 2648 574 2670
rect 1822 2668 1823 2672
rect 1827 2668 1828 2672
rect 1862 2669 1863 2673
rect 1867 2669 1868 2673
rect 2022 2671 2023 2675
rect 2027 2671 2028 2675
rect 2022 2670 2028 2671
rect 1862 2668 1868 2669
rect 1822 2667 1828 2668
rect 622 2659 628 2660
rect 622 2655 623 2659
rect 627 2655 628 2659
rect 622 2654 628 2655
rect 570 2647 576 2648
rect 570 2643 571 2647
rect 575 2643 576 2647
rect 570 2642 576 2643
rect 624 2627 626 2654
rect 654 2647 660 2648
rect 654 2643 655 2647
rect 659 2643 660 2647
rect 654 2642 660 2643
rect 287 2626 291 2627
rect 287 2621 291 2622
rect 351 2626 355 2627
rect 351 2621 355 2622
rect 399 2626 403 2627
rect 399 2621 403 2622
rect 495 2626 499 2627
rect 495 2621 499 2622
rect 511 2626 515 2627
rect 511 2621 515 2622
rect 623 2626 627 2627
rect 623 2621 627 2622
rect 250 2619 256 2620
rect 250 2615 251 2619
rect 255 2615 256 2619
rect 250 2614 256 2615
rect 352 2610 354 2621
rect 496 2610 498 2621
rect 222 2609 228 2610
rect 222 2605 223 2609
rect 227 2605 228 2609
rect 222 2604 228 2605
rect 350 2609 356 2610
rect 350 2605 351 2609
rect 355 2605 356 2609
rect 350 2604 356 2605
rect 494 2609 500 2610
rect 494 2605 495 2609
rect 499 2605 500 2609
rect 494 2604 500 2605
rect 110 2596 116 2597
rect 110 2592 111 2596
rect 115 2592 116 2596
rect 656 2592 658 2642
rect 1824 2627 1826 2667
rect 2010 2659 2016 2660
rect 1862 2656 1868 2657
rect 1862 2652 1863 2656
rect 1867 2652 1868 2656
rect 2010 2655 2011 2659
rect 2015 2655 2016 2659
rect 2010 2654 2016 2655
rect 2122 2659 2128 2660
rect 2122 2655 2123 2659
rect 2127 2655 2128 2659
rect 2122 2654 2128 2655
rect 1862 2651 1868 2652
rect 663 2626 667 2627
rect 663 2621 667 2622
rect 839 2626 843 2627
rect 839 2621 843 2622
rect 1023 2626 1027 2627
rect 1023 2621 1027 2622
rect 1215 2626 1219 2627
rect 1215 2621 1219 2622
rect 1407 2626 1411 2627
rect 1407 2621 1411 2622
rect 1607 2626 1611 2627
rect 1607 2621 1611 2622
rect 1823 2626 1827 2627
rect 1864 2623 1866 2651
rect 1950 2643 1956 2644
rect 1950 2639 1951 2643
rect 1955 2639 1956 2643
rect 1950 2638 1956 2639
rect 1952 2623 1954 2638
rect 2012 2632 2014 2654
rect 2062 2643 2068 2644
rect 2062 2639 2063 2643
rect 2067 2639 2068 2643
rect 2062 2638 2068 2639
rect 2010 2631 2016 2632
rect 2010 2627 2011 2631
rect 2015 2627 2016 2631
rect 2010 2626 2016 2627
rect 2064 2623 2066 2638
rect 2124 2632 2126 2654
rect 2174 2643 2180 2644
rect 2174 2639 2175 2643
rect 2179 2639 2180 2643
rect 2174 2638 2180 2639
rect 2294 2643 2300 2644
rect 2294 2639 2295 2643
rect 2299 2639 2300 2643
rect 2294 2638 2300 2639
rect 2122 2631 2128 2632
rect 2122 2627 2123 2631
rect 2127 2627 2128 2631
rect 2122 2626 2128 2627
rect 2176 2623 2178 2638
rect 2238 2631 2244 2632
rect 2238 2627 2239 2631
rect 2243 2627 2244 2631
rect 2238 2626 2244 2627
rect 1823 2621 1827 2622
rect 1863 2622 1867 2623
rect 664 2610 666 2621
rect 758 2619 764 2620
rect 758 2615 759 2619
rect 763 2615 764 2619
rect 758 2614 764 2615
rect 662 2609 668 2610
rect 662 2605 663 2609
rect 667 2605 668 2609
rect 662 2604 668 2605
rect 760 2592 762 2614
rect 840 2610 842 2621
rect 906 2619 912 2620
rect 906 2615 907 2619
rect 911 2615 912 2619
rect 906 2614 912 2615
rect 966 2619 972 2620
rect 966 2615 967 2619
rect 971 2615 972 2619
rect 966 2614 972 2615
rect 838 2609 844 2610
rect 838 2605 839 2609
rect 843 2605 844 2609
rect 838 2604 844 2605
rect 908 2592 910 2614
rect 110 2591 116 2592
rect 654 2591 660 2592
rect 654 2587 655 2591
rect 659 2587 660 2591
rect 654 2586 660 2587
rect 758 2591 764 2592
rect 758 2587 759 2591
rect 763 2587 764 2591
rect 758 2586 764 2587
rect 906 2591 912 2592
rect 906 2587 907 2591
rect 911 2587 912 2591
rect 906 2586 912 2587
rect 110 2579 116 2580
rect 110 2575 111 2579
rect 115 2575 116 2579
rect 110 2574 116 2575
rect 494 2579 500 2580
rect 494 2575 495 2579
rect 499 2575 500 2579
rect 494 2574 500 2575
rect 112 2559 114 2574
rect 214 2569 220 2570
rect 214 2565 215 2569
rect 219 2565 220 2569
rect 214 2564 220 2565
rect 342 2569 348 2570
rect 342 2565 343 2569
rect 347 2565 348 2569
rect 342 2564 348 2565
rect 486 2569 492 2570
rect 486 2565 487 2569
rect 491 2565 492 2569
rect 486 2564 492 2565
rect 216 2559 218 2564
rect 344 2559 346 2564
rect 488 2559 490 2564
rect 111 2558 115 2559
rect 111 2553 115 2554
rect 215 2558 219 2559
rect 215 2553 219 2554
rect 271 2558 275 2559
rect 271 2553 275 2554
rect 343 2558 347 2559
rect 343 2553 347 2554
rect 471 2558 475 2559
rect 471 2553 475 2554
rect 487 2558 491 2559
rect 487 2553 491 2554
rect 112 2538 114 2553
rect 272 2548 274 2553
rect 472 2548 474 2553
rect 270 2547 276 2548
rect 270 2543 271 2547
rect 275 2543 276 2547
rect 270 2542 276 2543
rect 470 2547 476 2548
rect 470 2543 471 2547
rect 475 2543 476 2547
rect 470 2542 476 2543
rect 110 2537 116 2538
rect 110 2533 111 2537
rect 115 2533 116 2537
rect 110 2532 116 2533
rect 214 2523 220 2524
rect 110 2520 116 2521
rect 110 2516 111 2520
rect 115 2516 116 2520
rect 214 2519 215 2523
rect 219 2519 220 2523
rect 214 2518 220 2519
rect 338 2523 344 2524
rect 338 2519 339 2523
rect 343 2519 344 2523
rect 338 2518 344 2519
rect 110 2515 116 2516
rect 112 2487 114 2515
rect 111 2486 115 2487
rect 111 2481 115 2482
rect 183 2486 187 2487
rect 183 2481 187 2482
rect 112 2457 114 2481
rect 184 2470 186 2481
rect 216 2480 218 2518
rect 278 2507 284 2508
rect 278 2503 279 2507
rect 283 2503 284 2507
rect 278 2502 284 2503
rect 280 2487 282 2502
rect 340 2496 342 2518
rect 478 2507 484 2508
rect 478 2503 479 2507
rect 483 2503 484 2507
rect 478 2502 484 2503
rect 338 2495 344 2496
rect 338 2491 339 2495
rect 343 2491 344 2495
rect 338 2490 344 2491
rect 480 2487 482 2502
rect 496 2496 498 2574
rect 654 2569 660 2570
rect 654 2565 655 2569
rect 659 2565 660 2569
rect 654 2564 660 2565
rect 830 2569 836 2570
rect 830 2565 831 2569
rect 835 2565 836 2569
rect 830 2564 836 2565
rect 656 2559 658 2564
rect 832 2559 834 2564
rect 655 2558 659 2559
rect 655 2553 659 2554
rect 671 2558 675 2559
rect 671 2553 675 2554
rect 831 2558 835 2559
rect 831 2553 835 2554
rect 855 2558 859 2559
rect 855 2553 859 2554
rect 672 2548 674 2553
rect 856 2548 858 2553
rect 670 2547 676 2548
rect 670 2543 671 2547
rect 675 2543 676 2547
rect 670 2542 676 2543
rect 854 2547 860 2548
rect 854 2543 855 2547
rect 859 2543 860 2547
rect 854 2542 860 2543
rect 968 2540 970 2614
rect 1024 2610 1026 2621
rect 1216 2610 1218 2621
rect 1246 2619 1252 2620
rect 1246 2615 1247 2619
rect 1251 2615 1252 2619
rect 1246 2614 1252 2615
rect 1022 2609 1028 2610
rect 1022 2605 1023 2609
rect 1027 2605 1028 2609
rect 1022 2604 1028 2605
rect 1214 2609 1220 2610
rect 1214 2605 1215 2609
rect 1219 2605 1220 2609
rect 1214 2604 1220 2605
rect 1014 2569 1020 2570
rect 1014 2565 1015 2569
rect 1019 2565 1020 2569
rect 1014 2564 1020 2565
rect 1206 2569 1212 2570
rect 1206 2565 1207 2569
rect 1211 2565 1212 2569
rect 1206 2564 1212 2565
rect 1016 2559 1018 2564
rect 1208 2559 1210 2564
rect 1015 2558 1019 2559
rect 1015 2553 1019 2554
rect 1023 2558 1027 2559
rect 1023 2553 1027 2554
rect 1175 2558 1179 2559
rect 1175 2553 1179 2554
rect 1207 2558 1211 2559
rect 1207 2553 1211 2554
rect 1024 2548 1026 2553
rect 1176 2548 1178 2553
rect 1022 2547 1028 2548
rect 1022 2543 1023 2547
rect 1027 2543 1028 2547
rect 1022 2542 1028 2543
rect 1174 2547 1180 2548
rect 1174 2543 1175 2547
rect 1179 2543 1180 2547
rect 1174 2542 1180 2543
rect 1248 2540 1250 2614
rect 1408 2610 1410 2621
rect 1608 2610 1610 2621
rect 1406 2609 1412 2610
rect 1406 2605 1407 2609
rect 1411 2605 1412 2609
rect 1406 2604 1412 2605
rect 1606 2609 1612 2610
rect 1606 2605 1607 2609
rect 1611 2605 1612 2609
rect 1606 2604 1612 2605
rect 1824 2597 1826 2621
rect 1863 2617 1867 2618
rect 1895 2622 1899 2623
rect 1895 2617 1899 2618
rect 1951 2622 1955 2623
rect 1951 2617 1955 2618
rect 2063 2622 2067 2623
rect 2063 2617 2067 2618
rect 2071 2622 2075 2623
rect 2071 2617 2075 2618
rect 2175 2622 2179 2623
rect 2175 2617 2179 2618
rect 1822 2596 1828 2597
rect 1822 2592 1823 2596
rect 1827 2592 1828 2596
rect 1864 2593 1866 2617
rect 1896 2606 1898 2617
rect 1958 2615 1964 2616
rect 1958 2611 1959 2615
rect 1963 2611 1964 2615
rect 1958 2610 1964 2611
rect 1894 2605 1900 2606
rect 1894 2601 1895 2605
rect 1899 2601 1900 2605
rect 1894 2600 1900 2601
rect 1822 2591 1828 2592
rect 1862 2592 1868 2593
rect 1862 2588 1863 2592
rect 1867 2588 1868 2592
rect 1862 2587 1868 2588
rect 1762 2579 1768 2580
rect 1762 2575 1763 2579
rect 1767 2575 1768 2579
rect 1762 2574 1768 2575
rect 1822 2579 1828 2580
rect 1822 2575 1823 2579
rect 1827 2575 1828 2579
rect 1822 2574 1828 2575
rect 1862 2575 1868 2576
rect 1398 2569 1404 2570
rect 1398 2565 1399 2569
rect 1403 2565 1404 2569
rect 1398 2564 1404 2565
rect 1598 2569 1604 2570
rect 1598 2565 1599 2569
rect 1603 2565 1604 2569
rect 1598 2564 1604 2565
rect 1400 2559 1402 2564
rect 1600 2559 1602 2564
rect 1319 2558 1323 2559
rect 1319 2553 1323 2554
rect 1399 2558 1403 2559
rect 1399 2553 1403 2554
rect 1455 2558 1459 2559
rect 1455 2553 1459 2554
rect 1591 2558 1595 2559
rect 1591 2553 1595 2554
rect 1599 2558 1603 2559
rect 1599 2553 1603 2554
rect 1727 2558 1731 2559
rect 1727 2553 1731 2554
rect 1320 2548 1322 2553
rect 1456 2548 1458 2553
rect 1592 2548 1594 2553
rect 1728 2548 1730 2553
rect 1318 2547 1324 2548
rect 1318 2543 1319 2547
rect 1323 2543 1324 2547
rect 1318 2542 1324 2543
rect 1454 2547 1460 2548
rect 1454 2543 1455 2547
rect 1459 2543 1460 2547
rect 1454 2542 1460 2543
rect 1590 2547 1596 2548
rect 1590 2543 1591 2547
rect 1595 2543 1596 2547
rect 1590 2542 1596 2543
rect 1726 2547 1732 2548
rect 1726 2543 1727 2547
rect 1731 2543 1732 2547
rect 1726 2542 1732 2543
rect 966 2539 972 2540
rect 966 2535 967 2539
rect 971 2535 972 2539
rect 966 2534 972 2535
rect 1246 2539 1252 2540
rect 1246 2535 1247 2539
rect 1251 2535 1252 2539
rect 1246 2534 1252 2535
rect 1158 2523 1164 2524
rect 1158 2519 1159 2523
rect 1163 2519 1164 2523
rect 1158 2518 1164 2519
rect 1386 2523 1392 2524
rect 1386 2519 1387 2523
rect 1391 2519 1392 2523
rect 1386 2518 1392 2519
rect 1522 2523 1528 2524
rect 1522 2519 1523 2523
rect 1527 2519 1528 2523
rect 1522 2518 1528 2519
rect 1658 2523 1664 2524
rect 1658 2519 1659 2523
rect 1663 2519 1664 2523
rect 1658 2518 1664 2519
rect 678 2507 684 2508
rect 678 2503 679 2507
rect 683 2503 684 2507
rect 678 2502 684 2503
rect 862 2507 868 2508
rect 862 2503 863 2507
rect 867 2503 868 2507
rect 862 2502 868 2503
rect 1030 2507 1036 2508
rect 1030 2503 1031 2507
rect 1035 2503 1036 2507
rect 1030 2502 1036 2503
rect 494 2495 500 2496
rect 494 2491 495 2495
rect 499 2491 500 2495
rect 494 2490 500 2491
rect 680 2487 682 2502
rect 864 2487 866 2502
rect 1032 2487 1034 2502
rect 1160 2496 1162 2518
rect 1182 2507 1188 2508
rect 1182 2503 1183 2507
rect 1187 2503 1188 2507
rect 1182 2502 1188 2503
rect 1326 2507 1332 2508
rect 1326 2503 1327 2507
rect 1331 2503 1332 2507
rect 1326 2502 1332 2503
rect 1062 2495 1068 2496
rect 1062 2491 1063 2495
rect 1067 2491 1068 2495
rect 1062 2490 1068 2491
rect 1158 2495 1164 2496
rect 1158 2491 1159 2495
rect 1163 2491 1164 2495
rect 1158 2490 1164 2491
rect 279 2486 283 2487
rect 279 2481 283 2482
rect 319 2486 323 2487
rect 319 2481 323 2482
rect 463 2486 467 2487
rect 463 2481 467 2482
rect 479 2486 483 2487
rect 479 2481 483 2482
rect 607 2486 611 2487
rect 607 2481 611 2482
rect 679 2486 683 2487
rect 679 2481 683 2482
rect 743 2486 747 2487
rect 743 2481 747 2482
rect 863 2486 867 2487
rect 863 2481 867 2482
rect 879 2486 883 2487
rect 879 2481 883 2482
rect 1007 2486 1011 2487
rect 1007 2481 1011 2482
rect 1031 2486 1035 2487
rect 1031 2481 1035 2482
rect 214 2479 220 2480
rect 214 2475 215 2479
rect 219 2475 220 2479
rect 214 2474 220 2475
rect 302 2479 308 2480
rect 302 2475 303 2479
rect 307 2475 308 2479
rect 302 2474 308 2475
rect 182 2469 188 2470
rect 182 2465 183 2469
rect 187 2465 188 2469
rect 182 2464 188 2465
rect 110 2456 116 2457
rect 304 2456 306 2474
rect 320 2470 322 2481
rect 464 2470 466 2481
rect 608 2470 610 2481
rect 744 2470 746 2481
rect 880 2470 882 2481
rect 1008 2470 1010 2481
rect 318 2469 324 2470
rect 318 2465 319 2469
rect 323 2465 324 2469
rect 318 2464 324 2465
rect 462 2469 468 2470
rect 462 2465 463 2469
rect 467 2465 468 2469
rect 462 2464 468 2465
rect 606 2469 612 2470
rect 606 2465 607 2469
rect 611 2465 612 2469
rect 606 2464 612 2465
rect 742 2469 748 2470
rect 742 2465 743 2469
rect 747 2465 748 2469
rect 742 2464 748 2465
rect 878 2469 884 2470
rect 878 2465 879 2469
rect 883 2465 884 2469
rect 878 2464 884 2465
rect 1006 2469 1012 2470
rect 1006 2465 1007 2469
rect 1011 2465 1012 2469
rect 1006 2464 1012 2465
rect 1064 2464 1066 2490
rect 1184 2487 1186 2502
rect 1328 2487 1330 2502
rect 1388 2488 1390 2518
rect 1462 2507 1468 2508
rect 1462 2503 1463 2507
rect 1467 2503 1468 2507
rect 1462 2502 1468 2503
rect 1386 2487 1392 2488
rect 1464 2487 1466 2502
rect 1524 2496 1526 2518
rect 1598 2507 1604 2508
rect 1598 2503 1599 2507
rect 1603 2503 1604 2507
rect 1598 2502 1604 2503
rect 1522 2495 1528 2496
rect 1522 2491 1523 2495
rect 1527 2491 1528 2495
rect 1522 2490 1528 2491
rect 1600 2487 1602 2502
rect 1660 2496 1662 2518
rect 1734 2507 1740 2508
rect 1734 2503 1735 2507
rect 1739 2503 1740 2507
rect 1734 2502 1740 2503
rect 1658 2495 1664 2496
rect 1658 2491 1659 2495
rect 1663 2491 1664 2495
rect 1658 2490 1664 2491
rect 1736 2487 1738 2502
rect 1764 2496 1766 2574
rect 1824 2559 1826 2574
rect 1862 2571 1863 2575
rect 1867 2571 1868 2575
rect 1862 2570 1868 2571
rect 1823 2558 1827 2559
rect 1864 2555 1866 2570
rect 1886 2565 1892 2566
rect 1886 2561 1887 2565
rect 1891 2561 1892 2565
rect 1886 2560 1892 2561
rect 1888 2555 1890 2560
rect 1823 2553 1827 2554
rect 1863 2554 1867 2555
rect 1824 2538 1826 2553
rect 1863 2549 1867 2550
rect 1887 2554 1891 2555
rect 1887 2549 1891 2550
rect 1822 2537 1828 2538
rect 1822 2533 1823 2537
rect 1827 2533 1828 2537
rect 1864 2534 1866 2549
rect 1888 2544 1890 2549
rect 1886 2543 1892 2544
rect 1886 2539 1887 2543
rect 1891 2539 1892 2543
rect 1886 2538 1892 2539
rect 1960 2536 1962 2610
rect 2072 2606 2074 2617
rect 2070 2605 2076 2606
rect 2070 2601 2071 2605
rect 2075 2601 2076 2605
rect 2070 2600 2076 2601
rect 2240 2588 2242 2626
rect 2296 2623 2298 2638
rect 2372 2632 2374 2710
rect 2438 2705 2444 2706
rect 2438 2701 2439 2705
rect 2443 2701 2444 2705
rect 2438 2700 2444 2701
rect 2440 2695 2442 2700
rect 2407 2694 2411 2695
rect 2407 2689 2411 2690
rect 2439 2694 2443 2695
rect 2439 2689 2443 2690
rect 2519 2694 2523 2695
rect 2519 2689 2523 2690
rect 2408 2684 2410 2689
rect 2520 2684 2522 2689
rect 2406 2683 2412 2684
rect 2406 2679 2407 2683
rect 2411 2679 2412 2683
rect 2406 2678 2412 2679
rect 2518 2683 2524 2684
rect 2518 2679 2519 2683
rect 2523 2679 2524 2683
rect 2518 2678 2524 2679
rect 2490 2659 2496 2660
rect 2490 2655 2491 2659
rect 2495 2655 2496 2659
rect 2490 2654 2496 2655
rect 2414 2643 2420 2644
rect 2414 2639 2415 2643
rect 2419 2639 2420 2643
rect 2414 2638 2420 2639
rect 2370 2631 2376 2632
rect 2370 2627 2371 2631
rect 2375 2627 2376 2631
rect 2370 2626 2376 2627
rect 2416 2623 2418 2638
rect 2263 2622 2267 2623
rect 2263 2617 2267 2618
rect 2295 2622 2299 2623
rect 2295 2617 2299 2618
rect 2415 2622 2419 2623
rect 2415 2617 2419 2618
rect 2463 2622 2467 2623
rect 2463 2617 2467 2618
rect 2264 2606 2266 2617
rect 2464 2606 2466 2617
rect 2492 2616 2494 2654
rect 2526 2643 2532 2644
rect 2526 2639 2527 2643
rect 2531 2639 2532 2643
rect 2526 2638 2532 2639
rect 2528 2623 2530 2638
rect 2560 2632 2562 2710
rect 2614 2705 2620 2706
rect 2614 2701 2615 2705
rect 2619 2701 2620 2705
rect 2614 2700 2620 2701
rect 2814 2705 2820 2706
rect 2814 2701 2815 2705
rect 2819 2701 2820 2705
rect 2814 2700 2820 2701
rect 3030 2705 3036 2706
rect 3030 2701 3031 2705
rect 3035 2701 3036 2705
rect 3030 2700 3036 2701
rect 2616 2695 2618 2700
rect 2816 2695 2818 2700
rect 3032 2695 3034 2700
rect 2615 2694 2619 2695
rect 2615 2689 2619 2690
rect 2631 2694 2635 2695
rect 2631 2689 2635 2690
rect 2735 2694 2739 2695
rect 2735 2689 2739 2690
rect 2815 2694 2819 2695
rect 2815 2689 2819 2690
rect 2847 2694 2851 2695
rect 2847 2689 2851 2690
rect 2959 2694 2963 2695
rect 2959 2689 2963 2690
rect 3031 2694 3035 2695
rect 3031 2689 3035 2690
rect 3071 2694 3075 2695
rect 3071 2689 3075 2690
rect 2632 2684 2634 2689
rect 2736 2684 2738 2689
rect 2848 2684 2850 2689
rect 2960 2684 2962 2689
rect 3072 2684 3074 2689
rect 2630 2683 2636 2684
rect 2630 2679 2631 2683
rect 2635 2679 2636 2683
rect 2630 2678 2636 2679
rect 2734 2683 2740 2684
rect 2734 2679 2735 2683
rect 2739 2679 2740 2683
rect 2734 2678 2740 2679
rect 2846 2683 2852 2684
rect 2846 2679 2847 2683
rect 2851 2679 2852 2683
rect 2846 2678 2852 2679
rect 2958 2683 2964 2684
rect 2958 2679 2959 2683
rect 2963 2679 2964 2683
rect 2958 2678 2964 2679
rect 3070 2683 3076 2684
rect 3070 2679 3071 2683
rect 3075 2679 3076 2683
rect 3070 2678 3076 2679
rect 3200 2676 3202 2750
rect 3272 2746 3274 2757
rect 3488 2746 3490 2757
rect 3548 2756 3550 2802
rect 3574 2800 3575 2804
rect 3579 2800 3580 2804
rect 3574 2799 3580 2800
rect 3576 2763 3578 2799
rect 3575 2762 3579 2763
rect 3575 2757 3579 2758
rect 3546 2755 3552 2756
rect 3546 2751 3547 2755
rect 3551 2751 3552 2755
rect 3546 2750 3552 2751
rect 3270 2745 3276 2746
rect 3270 2741 3271 2745
rect 3275 2741 3276 2745
rect 3270 2740 3276 2741
rect 3486 2745 3492 2746
rect 3486 2741 3487 2745
rect 3491 2741 3492 2745
rect 3486 2740 3492 2741
rect 3576 2733 3578 2757
rect 3574 2732 3580 2733
rect 3574 2728 3575 2732
rect 3579 2728 3580 2732
rect 3574 2727 3580 2728
rect 3574 2715 3580 2716
rect 3574 2711 3575 2715
rect 3579 2711 3580 2715
rect 3574 2710 3580 2711
rect 3262 2705 3268 2706
rect 3262 2701 3263 2705
rect 3267 2701 3268 2705
rect 3262 2700 3268 2701
rect 3478 2705 3484 2706
rect 3478 2701 3479 2705
rect 3483 2701 3484 2705
rect 3478 2700 3484 2701
rect 3264 2695 3266 2700
rect 3480 2695 3482 2700
rect 3518 2699 3524 2700
rect 3518 2695 3519 2699
rect 3523 2695 3524 2699
rect 3576 2695 3578 2710
rect 3263 2694 3267 2695
rect 3263 2689 3267 2690
rect 3479 2694 3483 2695
rect 3518 2694 3524 2695
rect 3575 2694 3579 2695
rect 3479 2689 3483 2690
rect 3198 2675 3204 2676
rect 3198 2671 3199 2675
rect 3203 2671 3204 2675
rect 3198 2670 3204 2671
rect 2638 2643 2644 2644
rect 2638 2639 2639 2643
rect 2643 2639 2644 2643
rect 2638 2638 2644 2639
rect 2742 2643 2748 2644
rect 2742 2639 2743 2643
rect 2747 2639 2748 2643
rect 2742 2638 2748 2639
rect 2854 2643 2860 2644
rect 2854 2639 2855 2643
rect 2859 2639 2860 2643
rect 2854 2638 2860 2639
rect 2966 2643 2972 2644
rect 2966 2639 2967 2643
rect 2971 2639 2972 2643
rect 2966 2638 2972 2639
rect 3078 2643 3084 2644
rect 3078 2639 3079 2643
rect 3083 2639 3084 2643
rect 3078 2638 3084 2639
rect 2558 2631 2564 2632
rect 2558 2627 2559 2631
rect 2563 2627 2564 2631
rect 2558 2626 2564 2627
rect 2640 2623 2642 2638
rect 2744 2623 2746 2638
rect 2856 2623 2858 2638
rect 2968 2623 2970 2638
rect 3080 2623 3082 2638
rect 2527 2622 2531 2623
rect 2527 2617 2531 2618
rect 2639 2622 2643 2623
rect 2639 2617 2643 2618
rect 2663 2622 2667 2623
rect 2663 2617 2667 2618
rect 2743 2622 2747 2623
rect 2743 2617 2747 2618
rect 2855 2622 2859 2623
rect 2855 2617 2859 2618
rect 2871 2622 2875 2623
rect 2871 2617 2875 2618
rect 2967 2622 2971 2623
rect 2967 2617 2971 2618
rect 3079 2622 3083 2623
rect 3079 2617 3083 2618
rect 3295 2622 3299 2623
rect 3295 2617 3299 2618
rect 3487 2622 3491 2623
rect 3487 2617 3491 2618
rect 2490 2615 2496 2616
rect 2490 2611 2491 2615
rect 2495 2611 2496 2615
rect 2490 2610 2496 2611
rect 2664 2606 2666 2617
rect 2872 2606 2874 2617
rect 2958 2615 2964 2616
rect 2958 2611 2959 2615
rect 2963 2611 2964 2615
rect 2958 2610 2964 2611
rect 2262 2605 2268 2606
rect 2262 2601 2263 2605
rect 2267 2601 2268 2605
rect 2262 2600 2268 2601
rect 2462 2605 2468 2606
rect 2462 2601 2463 2605
rect 2467 2601 2468 2605
rect 2462 2600 2468 2601
rect 2662 2605 2668 2606
rect 2662 2601 2663 2605
rect 2667 2601 2668 2605
rect 2662 2600 2668 2601
rect 2870 2605 2876 2606
rect 2870 2601 2871 2605
rect 2875 2601 2876 2605
rect 2870 2600 2876 2601
rect 2960 2588 2962 2610
rect 3080 2606 3082 2617
rect 3296 2606 3298 2617
rect 3488 2606 3490 2617
rect 3520 2616 3522 2694
rect 3575 2689 3579 2690
rect 3576 2674 3578 2689
rect 3574 2673 3580 2674
rect 3574 2669 3575 2673
rect 3579 2669 3580 2673
rect 3574 2668 3580 2669
rect 3574 2656 3580 2657
rect 3574 2652 3575 2656
rect 3579 2652 3580 2656
rect 3574 2651 3580 2652
rect 3576 2623 3578 2651
rect 3575 2622 3579 2623
rect 3575 2617 3579 2618
rect 3518 2615 3524 2616
rect 3518 2611 3519 2615
rect 3523 2611 3524 2615
rect 3518 2610 3524 2611
rect 3078 2605 3084 2606
rect 3078 2601 3079 2605
rect 3083 2601 3084 2605
rect 3078 2600 3084 2601
rect 3294 2605 3300 2606
rect 3294 2601 3295 2605
rect 3299 2601 3300 2605
rect 3294 2600 3300 2601
rect 3486 2605 3492 2606
rect 3486 2601 3487 2605
rect 3491 2601 3492 2605
rect 3486 2600 3492 2601
rect 3576 2593 3578 2617
rect 3574 2592 3580 2593
rect 3574 2588 3575 2592
rect 3579 2588 3580 2592
rect 2238 2587 2244 2588
rect 2238 2583 2239 2587
rect 2243 2583 2244 2587
rect 2238 2582 2244 2583
rect 2958 2587 2964 2588
rect 3574 2587 3580 2588
rect 2958 2583 2959 2587
rect 2963 2583 2964 2587
rect 2958 2582 2964 2583
rect 2530 2575 2536 2576
rect 2530 2571 2531 2575
rect 2535 2571 2536 2575
rect 2530 2570 2536 2571
rect 2782 2575 2788 2576
rect 2782 2571 2783 2575
rect 2787 2571 2788 2575
rect 2782 2570 2788 2571
rect 3574 2575 3580 2576
rect 3574 2571 3575 2575
rect 3579 2571 3580 2575
rect 3574 2570 3580 2571
rect 2062 2565 2068 2566
rect 2062 2561 2063 2565
rect 2067 2561 2068 2565
rect 2062 2560 2068 2561
rect 2254 2565 2260 2566
rect 2254 2561 2255 2565
rect 2259 2561 2260 2565
rect 2254 2560 2260 2561
rect 2454 2565 2460 2566
rect 2454 2561 2455 2565
rect 2459 2561 2460 2565
rect 2454 2560 2460 2561
rect 2064 2555 2066 2560
rect 2256 2555 2258 2560
rect 2456 2555 2458 2560
rect 2039 2554 2043 2555
rect 2039 2549 2043 2550
rect 2063 2554 2067 2555
rect 2063 2549 2067 2550
rect 2215 2554 2219 2555
rect 2215 2549 2219 2550
rect 2255 2554 2259 2555
rect 2255 2549 2259 2550
rect 2399 2554 2403 2555
rect 2399 2549 2403 2550
rect 2455 2554 2459 2555
rect 2455 2549 2459 2550
rect 2040 2544 2042 2549
rect 2216 2544 2218 2549
rect 2400 2544 2402 2549
rect 2038 2543 2044 2544
rect 2038 2539 2039 2543
rect 2043 2539 2044 2543
rect 2038 2538 2044 2539
rect 2214 2543 2220 2544
rect 2214 2539 2215 2543
rect 2219 2539 2220 2543
rect 2214 2538 2220 2539
rect 2398 2543 2404 2544
rect 2398 2539 2399 2543
rect 2403 2539 2404 2543
rect 2398 2538 2404 2539
rect 1958 2535 1964 2536
rect 1822 2532 1828 2533
rect 1862 2533 1868 2534
rect 1862 2529 1863 2533
rect 1867 2529 1868 2533
rect 1958 2531 1959 2535
rect 1963 2531 1964 2535
rect 1958 2530 1964 2531
rect 1862 2528 1868 2529
rect 1822 2520 1828 2521
rect 1822 2516 1823 2520
rect 1827 2516 1828 2520
rect 1954 2519 1960 2520
rect 1822 2515 1828 2516
rect 1862 2516 1868 2517
rect 1762 2495 1768 2496
rect 1762 2491 1763 2495
rect 1767 2491 1768 2495
rect 1762 2490 1768 2491
rect 1824 2487 1826 2515
rect 1862 2512 1863 2516
rect 1867 2512 1868 2516
rect 1954 2515 1955 2519
rect 1959 2515 1960 2519
rect 1954 2514 1960 2515
rect 2106 2519 2112 2520
rect 2106 2515 2107 2519
rect 2111 2515 2112 2519
rect 2106 2514 2112 2515
rect 1862 2511 1868 2512
rect 1864 2487 1866 2511
rect 1894 2503 1900 2504
rect 1894 2499 1895 2503
rect 1899 2499 1900 2503
rect 1894 2498 1900 2499
rect 1896 2487 1898 2498
rect 1956 2492 1958 2514
rect 2046 2503 2052 2504
rect 2046 2499 2047 2503
rect 2051 2499 2052 2503
rect 2046 2498 2052 2499
rect 1954 2491 1960 2492
rect 1954 2487 1955 2491
rect 1959 2487 1960 2491
rect 2048 2487 2050 2498
rect 2108 2492 2110 2514
rect 2222 2503 2228 2504
rect 2222 2499 2223 2503
rect 2227 2499 2228 2503
rect 2222 2498 2228 2499
rect 2406 2503 2412 2504
rect 2406 2499 2407 2503
rect 2411 2499 2412 2503
rect 2406 2498 2412 2499
rect 2106 2491 2112 2492
rect 2106 2487 2107 2491
rect 2111 2487 2112 2491
rect 2224 2487 2226 2498
rect 2270 2491 2276 2492
rect 2270 2487 2271 2491
rect 2275 2487 2276 2491
rect 2408 2487 2410 2498
rect 2532 2492 2534 2570
rect 2654 2565 2660 2566
rect 2654 2561 2655 2565
rect 2659 2561 2660 2565
rect 2654 2560 2660 2561
rect 2656 2555 2658 2560
rect 2575 2554 2579 2555
rect 2575 2549 2579 2550
rect 2655 2554 2659 2555
rect 2655 2549 2659 2550
rect 2743 2554 2747 2555
rect 2743 2549 2747 2550
rect 2576 2544 2578 2549
rect 2744 2544 2746 2549
rect 2574 2543 2580 2544
rect 2574 2539 2575 2543
rect 2579 2539 2580 2543
rect 2574 2538 2580 2539
rect 2742 2543 2748 2544
rect 2742 2539 2743 2543
rect 2747 2539 2748 2543
rect 2742 2538 2748 2539
rect 2642 2519 2648 2520
rect 2642 2515 2643 2519
rect 2647 2515 2648 2519
rect 2642 2514 2648 2515
rect 2582 2503 2588 2504
rect 2582 2499 2583 2503
rect 2587 2499 2588 2503
rect 2582 2498 2588 2499
rect 2530 2491 2536 2492
rect 2530 2487 2531 2491
rect 2535 2487 2536 2491
rect 2584 2487 2586 2498
rect 1127 2486 1131 2487
rect 1127 2481 1131 2482
rect 1183 2486 1187 2487
rect 1183 2481 1187 2482
rect 1239 2486 1243 2487
rect 1239 2481 1243 2482
rect 1327 2486 1331 2487
rect 1327 2481 1331 2482
rect 1343 2486 1347 2487
rect 1386 2483 1387 2487
rect 1391 2483 1392 2487
rect 1386 2482 1392 2483
rect 1447 2486 1451 2487
rect 1343 2481 1347 2482
rect 1447 2481 1451 2482
rect 1463 2486 1467 2487
rect 1463 2481 1467 2482
rect 1551 2486 1555 2487
rect 1551 2481 1555 2482
rect 1599 2486 1603 2487
rect 1599 2481 1603 2482
rect 1647 2486 1651 2487
rect 1647 2481 1651 2482
rect 1735 2486 1739 2487
rect 1735 2481 1739 2482
rect 1823 2486 1827 2487
rect 1823 2481 1827 2482
rect 1863 2486 1867 2487
rect 1863 2481 1867 2482
rect 1895 2486 1899 2487
rect 1954 2486 1960 2487
rect 1991 2486 1995 2487
rect 1895 2481 1899 2482
rect 1991 2481 1995 2482
rect 2047 2486 2051 2487
rect 2106 2486 2112 2487
rect 2127 2486 2131 2487
rect 2047 2481 2051 2482
rect 2127 2481 2131 2482
rect 2223 2486 2227 2487
rect 2270 2486 2276 2487
rect 2279 2486 2283 2487
rect 2223 2481 2227 2482
rect 1074 2479 1080 2480
rect 1074 2475 1075 2479
rect 1079 2475 1080 2479
rect 1074 2474 1080 2475
rect 1062 2463 1068 2464
rect 1062 2459 1063 2463
rect 1067 2459 1068 2463
rect 1062 2458 1068 2459
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 110 2451 116 2452
rect 302 2455 308 2456
rect 302 2451 303 2455
rect 307 2451 308 2455
rect 1076 2452 1078 2474
rect 1128 2470 1130 2481
rect 1158 2479 1164 2480
rect 1158 2475 1159 2479
rect 1163 2475 1164 2479
rect 1158 2474 1164 2475
rect 1126 2469 1132 2470
rect 1126 2465 1127 2469
rect 1131 2465 1132 2469
rect 1126 2464 1132 2465
rect 302 2450 308 2451
rect 1074 2451 1080 2452
rect 1074 2447 1075 2451
rect 1079 2447 1080 2451
rect 1074 2446 1080 2447
rect 110 2439 116 2440
rect 110 2435 111 2439
rect 115 2435 116 2439
rect 110 2434 116 2435
rect 386 2439 392 2440
rect 386 2435 387 2439
rect 391 2435 392 2439
rect 386 2434 392 2435
rect 112 2411 114 2434
rect 174 2429 180 2430
rect 174 2425 175 2429
rect 179 2425 180 2429
rect 174 2424 180 2425
rect 310 2429 316 2430
rect 310 2425 311 2429
rect 315 2425 316 2429
rect 310 2424 316 2425
rect 176 2411 178 2424
rect 312 2411 314 2424
rect 111 2410 115 2411
rect 111 2405 115 2406
rect 151 2410 155 2411
rect 151 2405 155 2406
rect 175 2410 179 2411
rect 175 2405 179 2406
rect 311 2410 315 2411
rect 311 2405 315 2406
rect 319 2410 323 2411
rect 319 2405 323 2406
rect 112 2390 114 2405
rect 152 2400 154 2405
rect 320 2400 322 2405
rect 150 2399 156 2400
rect 150 2395 151 2399
rect 155 2395 156 2399
rect 150 2394 156 2395
rect 318 2399 324 2400
rect 318 2395 319 2399
rect 323 2395 324 2399
rect 318 2394 324 2395
rect 110 2389 116 2390
rect 110 2385 111 2389
rect 115 2385 116 2389
rect 110 2384 116 2385
rect 218 2375 224 2376
rect 110 2372 116 2373
rect 110 2368 111 2372
rect 115 2368 116 2372
rect 218 2371 219 2375
rect 223 2371 224 2375
rect 218 2370 224 2371
rect 226 2375 232 2376
rect 226 2371 227 2375
rect 231 2371 232 2375
rect 226 2370 232 2371
rect 110 2367 116 2368
rect 112 2339 114 2367
rect 158 2359 164 2360
rect 158 2355 159 2359
rect 163 2355 164 2359
rect 158 2354 164 2355
rect 160 2339 162 2354
rect 111 2338 115 2339
rect 111 2333 115 2334
rect 143 2338 147 2339
rect 143 2333 147 2334
rect 159 2338 163 2339
rect 159 2333 163 2334
rect 112 2309 114 2333
rect 144 2322 146 2333
rect 220 2332 222 2370
rect 228 2348 230 2370
rect 326 2359 332 2360
rect 326 2355 327 2359
rect 331 2355 332 2359
rect 326 2354 332 2355
rect 226 2347 232 2348
rect 226 2343 227 2347
rect 231 2343 232 2347
rect 226 2342 232 2343
rect 328 2339 330 2354
rect 388 2348 390 2434
rect 454 2429 460 2430
rect 454 2425 455 2429
rect 459 2425 460 2429
rect 454 2424 460 2425
rect 598 2429 604 2430
rect 598 2425 599 2429
rect 603 2425 604 2429
rect 598 2424 604 2425
rect 734 2429 740 2430
rect 734 2425 735 2429
rect 739 2425 740 2429
rect 734 2424 740 2425
rect 870 2429 876 2430
rect 870 2425 871 2429
rect 875 2425 876 2429
rect 870 2424 876 2425
rect 998 2429 1004 2430
rect 998 2425 999 2429
rect 1003 2425 1004 2429
rect 998 2424 1004 2425
rect 1118 2429 1124 2430
rect 1118 2425 1119 2429
rect 1123 2425 1124 2429
rect 1118 2424 1124 2425
rect 456 2411 458 2424
rect 600 2411 602 2424
rect 736 2411 738 2424
rect 872 2411 874 2424
rect 1000 2411 1002 2424
rect 1120 2411 1122 2424
rect 455 2410 459 2411
rect 455 2405 459 2406
rect 479 2410 483 2411
rect 479 2405 483 2406
rect 599 2410 603 2411
rect 599 2405 603 2406
rect 639 2410 643 2411
rect 639 2405 643 2406
rect 735 2410 739 2411
rect 735 2405 739 2406
rect 783 2410 787 2411
rect 783 2405 787 2406
rect 871 2410 875 2411
rect 871 2405 875 2406
rect 919 2410 923 2411
rect 919 2405 923 2406
rect 999 2410 1003 2411
rect 999 2405 1003 2406
rect 1047 2410 1051 2411
rect 1047 2405 1051 2406
rect 1119 2410 1123 2411
rect 1160 2408 1162 2474
rect 1240 2470 1242 2481
rect 1344 2470 1346 2481
rect 1448 2470 1450 2481
rect 1552 2470 1554 2481
rect 1648 2470 1650 2481
rect 1736 2470 1738 2481
rect 1238 2469 1244 2470
rect 1238 2465 1239 2469
rect 1243 2465 1244 2469
rect 1238 2464 1244 2465
rect 1342 2469 1348 2470
rect 1342 2465 1343 2469
rect 1347 2465 1348 2469
rect 1342 2464 1348 2465
rect 1446 2469 1452 2470
rect 1446 2465 1447 2469
rect 1451 2465 1452 2469
rect 1446 2464 1452 2465
rect 1550 2469 1556 2470
rect 1550 2465 1551 2469
rect 1555 2465 1556 2469
rect 1550 2464 1556 2465
rect 1646 2469 1652 2470
rect 1646 2465 1647 2469
rect 1651 2465 1652 2469
rect 1646 2464 1652 2465
rect 1734 2469 1740 2470
rect 1734 2465 1735 2469
rect 1739 2465 1740 2469
rect 1734 2464 1740 2465
rect 1824 2457 1826 2481
rect 1864 2457 1866 2481
rect 1896 2470 1898 2481
rect 1992 2470 1994 2481
rect 2128 2470 2130 2481
rect 1894 2469 1900 2470
rect 1894 2465 1895 2469
rect 1899 2465 1900 2469
rect 1894 2464 1900 2465
rect 1990 2469 1996 2470
rect 1990 2465 1991 2469
rect 1995 2465 1996 2469
rect 1990 2464 1996 2465
rect 2126 2469 2132 2470
rect 2126 2465 2127 2469
rect 2131 2465 2132 2469
rect 2126 2464 2132 2465
rect 1822 2456 1828 2457
rect 1822 2452 1823 2456
rect 1827 2452 1828 2456
rect 1822 2451 1828 2452
rect 1862 2456 1868 2457
rect 1862 2452 1863 2456
rect 1867 2452 1868 2456
rect 2272 2452 2274 2486
rect 2279 2481 2283 2482
rect 2407 2486 2411 2487
rect 2407 2481 2411 2482
rect 2439 2486 2443 2487
rect 2530 2486 2536 2487
rect 2583 2486 2587 2487
rect 2439 2481 2443 2482
rect 2583 2481 2587 2482
rect 2599 2486 2603 2487
rect 2599 2481 2603 2482
rect 2280 2470 2282 2481
rect 2440 2470 2442 2481
rect 2538 2479 2544 2480
rect 2538 2475 2539 2479
rect 2543 2475 2544 2479
rect 2538 2474 2544 2475
rect 2278 2469 2284 2470
rect 2278 2465 2279 2469
rect 2283 2465 2284 2469
rect 2278 2464 2284 2465
rect 2438 2469 2444 2470
rect 2438 2465 2439 2469
rect 2443 2465 2444 2469
rect 2438 2464 2444 2465
rect 2540 2452 2542 2474
rect 2600 2470 2602 2481
rect 2644 2480 2646 2514
rect 2750 2503 2756 2504
rect 2750 2499 2751 2503
rect 2755 2499 2756 2503
rect 2750 2498 2756 2499
rect 2752 2487 2754 2498
rect 2784 2492 2786 2570
rect 2862 2565 2868 2566
rect 2862 2561 2863 2565
rect 2867 2561 2868 2565
rect 2862 2560 2868 2561
rect 3070 2565 3076 2566
rect 3070 2561 3071 2565
rect 3075 2561 3076 2565
rect 3070 2560 3076 2561
rect 3286 2565 3292 2566
rect 3286 2561 3287 2565
rect 3291 2561 3292 2565
rect 3286 2560 3292 2561
rect 3478 2565 3484 2566
rect 3478 2561 3479 2565
rect 3483 2561 3484 2565
rect 3478 2560 3484 2561
rect 2864 2555 2866 2560
rect 3072 2555 3074 2560
rect 3288 2555 3290 2560
rect 3480 2555 3482 2560
rect 3518 2559 3524 2560
rect 3518 2555 3519 2559
rect 3523 2555 3524 2559
rect 3576 2555 3578 2570
rect 2863 2554 2867 2555
rect 2863 2549 2867 2550
rect 2903 2554 2907 2555
rect 2903 2549 2907 2550
rect 3055 2554 3059 2555
rect 3055 2549 3059 2550
rect 3071 2554 3075 2555
rect 3071 2549 3075 2550
rect 3199 2554 3203 2555
rect 3199 2549 3203 2550
rect 3287 2554 3291 2555
rect 3287 2549 3291 2550
rect 3343 2554 3347 2555
rect 3343 2549 3347 2550
rect 3479 2554 3483 2555
rect 3518 2554 3524 2555
rect 3575 2554 3579 2555
rect 3479 2549 3483 2550
rect 2904 2544 2906 2549
rect 3056 2544 3058 2549
rect 3200 2544 3202 2549
rect 3344 2544 3346 2549
rect 3480 2544 3482 2549
rect 2902 2543 2908 2544
rect 2902 2539 2903 2543
rect 2907 2539 2908 2543
rect 2902 2538 2908 2539
rect 3054 2543 3060 2544
rect 3054 2539 3055 2543
rect 3059 2539 3060 2543
rect 3054 2538 3060 2539
rect 3198 2543 3204 2544
rect 3198 2539 3199 2543
rect 3203 2539 3204 2543
rect 3198 2538 3204 2539
rect 3342 2543 3348 2544
rect 3342 2539 3343 2543
rect 3347 2539 3348 2543
rect 3342 2538 3348 2539
rect 3478 2543 3484 2544
rect 3478 2539 3479 2543
rect 3483 2539 3484 2543
rect 3478 2538 3484 2539
rect 3146 2519 3152 2520
rect 3146 2515 3147 2519
rect 3151 2515 3152 2519
rect 3146 2514 3152 2515
rect 3266 2519 3272 2520
rect 3266 2515 3267 2519
rect 3271 2515 3272 2519
rect 3266 2514 3272 2515
rect 2910 2503 2916 2504
rect 2910 2499 2911 2503
rect 2915 2499 2916 2503
rect 2910 2498 2916 2499
rect 3062 2503 3068 2504
rect 3062 2499 3063 2503
rect 3067 2499 3068 2503
rect 3062 2498 3068 2499
rect 2782 2491 2788 2492
rect 2782 2487 2783 2491
rect 2787 2487 2788 2491
rect 2912 2487 2914 2498
rect 3064 2487 3066 2498
rect 2751 2486 2755 2487
rect 2751 2481 2755 2482
rect 2767 2486 2771 2487
rect 2782 2486 2788 2487
rect 2911 2486 2915 2487
rect 2767 2481 2771 2482
rect 2911 2481 2915 2482
rect 2943 2486 2947 2487
rect 2943 2481 2947 2482
rect 3063 2486 3067 2487
rect 3063 2481 3067 2482
rect 3119 2486 3123 2487
rect 3119 2481 3123 2482
rect 2642 2479 2648 2480
rect 2642 2475 2643 2479
rect 2647 2475 2648 2479
rect 2642 2474 2648 2475
rect 2768 2470 2770 2481
rect 2874 2479 2880 2480
rect 2874 2475 2875 2479
rect 2879 2475 2880 2479
rect 2874 2474 2880 2475
rect 2598 2469 2604 2470
rect 2598 2465 2599 2469
rect 2603 2465 2604 2469
rect 2598 2464 2604 2465
rect 2766 2469 2772 2470
rect 2766 2465 2767 2469
rect 2771 2465 2772 2469
rect 2766 2464 2772 2465
rect 2876 2452 2878 2474
rect 2944 2470 2946 2481
rect 3050 2479 3056 2480
rect 3050 2475 3051 2479
rect 3055 2475 3056 2479
rect 3050 2474 3056 2475
rect 2942 2469 2948 2470
rect 2942 2465 2943 2469
rect 2947 2465 2948 2469
rect 2942 2464 2948 2465
rect 3052 2452 3054 2474
rect 3120 2470 3122 2481
rect 3148 2480 3150 2514
rect 3206 2503 3212 2504
rect 3206 2499 3207 2503
rect 3211 2499 3212 2503
rect 3206 2498 3212 2499
rect 3208 2487 3210 2498
rect 3268 2492 3270 2514
rect 3350 2503 3356 2504
rect 3350 2499 3351 2503
rect 3355 2499 3356 2503
rect 3350 2498 3356 2499
rect 3486 2503 3492 2504
rect 3486 2499 3487 2503
rect 3491 2499 3492 2503
rect 3486 2498 3492 2499
rect 3266 2491 3272 2492
rect 3266 2487 3267 2491
rect 3271 2487 3272 2491
rect 3352 2487 3354 2498
rect 3488 2487 3490 2498
rect 3520 2492 3522 2554
rect 3575 2549 3579 2550
rect 3576 2534 3578 2549
rect 3574 2533 3580 2534
rect 3574 2529 3575 2533
rect 3579 2529 3580 2533
rect 3574 2528 3580 2529
rect 3546 2519 3552 2520
rect 3546 2515 3547 2519
rect 3551 2515 3552 2519
rect 3546 2514 3552 2515
rect 3574 2516 3580 2517
rect 3518 2491 3524 2492
rect 3518 2487 3519 2491
rect 3523 2487 3524 2491
rect 3207 2486 3211 2487
rect 3266 2486 3272 2487
rect 3295 2486 3299 2487
rect 3207 2481 3211 2482
rect 3295 2481 3299 2482
rect 3351 2486 3355 2487
rect 3351 2481 3355 2482
rect 3471 2486 3475 2487
rect 3471 2481 3475 2482
rect 3487 2486 3491 2487
rect 3518 2486 3524 2487
rect 3487 2481 3491 2482
rect 3146 2479 3152 2480
rect 3146 2475 3147 2479
rect 3151 2475 3152 2479
rect 3146 2474 3152 2475
rect 3296 2470 3298 2481
rect 3310 2479 3316 2480
rect 3310 2475 3311 2479
rect 3315 2475 3316 2479
rect 3310 2474 3316 2475
rect 3118 2469 3124 2470
rect 3118 2465 3119 2469
rect 3123 2465 3124 2469
rect 3118 2464 3124 2465
rect 3294 2469 3300 2470
rect 3294 2465 3295 2469
rect 3299 2465 3300 2469
rect 3294 2464 3300 2465
rect 1862 2451 1868 2452
rect 2270 2451 2276 2452
rect 2270 2447 2271 2451
rect 2275 2447 2276 2451
rect 2270 2446 2276 2447
rect 2538 2451 2544 2452
rect 2538 2447 2539 2451
rect 2543 2447 2544 2451
rect 2538 2446 2544 2447
rect 2874 2451 2880 2452
rect 2874 2447 2875 2451
rect 2879 2447 2880 2451
rect 2874 2446 2880 2447
rect 3050 2451 3056 2452
rect 3050 2447 3051 2451
rect 3055 2447 3056 2451
rect 3050 2446 3056 2447
rect 1822 2439 1828 2440
rect 1822 2435 1823 2439
rect 1827 2435 1828 2439
rect 1822 2434 1828 2435
rect 1862 2439 1868 2440
rect 1862 2435 1863 2439
rect 1867 2435 1868 2439
rect 1862 2434 1868 2435
rect 2390 2439 2396 2440
rect 2390 2435 2391 2439
rect 2395 2435 2396 2439
rect 2390 2434 2396 2435
rect 2694 2439 2700 2440
rect 2694 2435 2695 2439
rect 2699 2435 2700 2439
rect 2694 2434 2700 2435
rect 1230 2429 1236 2430
rect 1230 2425 1231 2429
rect 1235 2425 1236 2429
rect 1230 2424 1236 2425
rect 1334 2429 1340 2430
rect 1334 2425 1335 2429
rect 1339 2425 1340 2429
rect 1334 2424 1340 2425
rect 1438 2429 1444 2430
rect 1438 2425 1439 2429
rect 1443 2425 1444 2429
rect 1438 2424 1444 2425
rect 1542 2429 1548 2430
rect 1542 2425 1543 2429
rect 1547 2425 1548 2429
rect 1542 2424 1548 2425
rect 1638 2429 1644 2430
rect 1638 2425 1639 2429
rect 1643 2425 1644 2429
rect 1638 2424 1644 2425
rect 1726 2429 1732 2430
rect 1726 2425 1727 2429
rect 1731 2425 1732 2429
rect 1726 2424 1732 2425
rect 1232 2411 1234 2424
rect 1336 2411 1338 2424
rect 1440 2411 1442 2424
rect 1544 2411 1546 2424
rect 1640 2411 1642 2424
rect 1728 2411 1730 2424
rect 1824 2411 1826 2434
rect 1864 2411 1866 2434
rect 1886 2429 1892 2430
rect 1886 2425 1887 2429
rect 1891 2425 1892 2429
rect 1886 2424 1892 2425
rect 1982 2429 1988 2430
rect 1982 2425 1983 2429
rect 1987 2425 1988 2429
rect 1982 2424 1988 2425
rect 2118 2429 2124 2430
rect 2118 2425 2119 2429
rect 2123 2425 2124 2429
rect 2118 2424 2124 2425
rect 2270 2429 2276 2430
rect 2270 2425 2271 2429
rect 2275 2425 2276 2429
rect 2270 2424 2276 2425
rect 1888 2411 1890 2424
rect 1984 2411 1986 2424
rect 2120 2411 2122 2424
rect 2272 2411 2274 2424
rect 1175 2410 1179 2411
rect 1119 2405 1123 2406
rect 1158 2407 1164 2408
rect 480 2400 482 2405
rect 640 2400 642 2405
rect 784 2400 786 2405
rect 920 2400 922 2405
rect 1048 2400 1050 2405
rect 1158 2403 1159 2407
rect 1163 2403 1164 2407
rect 1175 2405 1179 2406
rect 1231 2410 1235 2411
rect 1231 2405 1235 2406
rect 1303 2410 1307 2411
rect 1303 2405 1307 2406
rect 1335 2410 1339 2411
rect 1335 2405 1339 2406
rect 1431 2410 1435 2411
rect 1431 2405 1435 2406
rect 1439 2410 1443 2411
rect 1439 2405 1443 2406
rect 1543 2410 1547 2411
rect 1543 2405 1547 2406
rect 1639 2410 1643 2411
rect 1639 2405 1643 2406
rect 1727 2410 1731 2411
rect 1727 2405 1731 2406
rect 1823 2410 1827 2411
rect 1823 2405 1827 2406
rect 1863 2410 1867 2411
rect 1863 2405 1867 2406
rect 1887 2410 1891 2411
rect 1887 2405 1891 2406
rect 1983 2410 1987 2411
rect 1983 2405 1987 2406
rect 2119 2410 2123 2411
rect 2119 2405 2123 2406
rect 2271 2410 2275 2411
rect 2271 2405 2275 2406
rect 2351 2410 2355 2411
rect 2351 2405 2355 2406
rect 1158 2402 1164 2403
rect 1176 2400 1178 2405
rect 1304 2400 1306 2405
rect 1432 2400 1434 2405
rect 478 2399 484 2400
rect 478 2395 479 2399
rect 483 2395 484 2399
rect 478 2394 484 2395
rect 638 2399 644 2400
rect 638 2395 639 2399
rect 643 2395 644 2399
rect 638 2394 644 2395
rect 782 2399 788 2400
rect 782 2395 783 2399
rect 787 2395 788 2399
rect 782 2394 788 2395
rect 918 2399 924 2400
rect 918 2395 919 2399
rect 923 2395 924 2399
rect 918 2394 924 2395
rect 1046 2399 1052 2400
rect 1046 2395 1047 2399
rect 1051 2395 1052 2399
rect 1046 2394 1052 2395
rect 1174 2399 1180 2400
rect 1174 2395 1175 2399
rect 1179 2395 1180 2399
rect 1174 2394 1180 2395
rect 1302 2399 1308 2400
rect 1302 2395 1303 2399
rect 1307 2395 1308 2399
rect 1302 2394 1308 2395
rect 1430 2399 1436 2400
rect 1430 2395 1431 2399
rect 1435 2395 1436 2399
rect 1430 2394 1436 2395
rect 1824 2390 1826 2405
rect 1864 2390 1866 2405
rect 2352 2400 2354 2405
rect 2350 2399 2356 2400
rect 2350 2395 2351 2399
rect 2355 2395 2356 2399
rect 2350 2394 2356 2395
rect 1822 2389 1828 2390
rect 1822 2385 1823 2389
rect 1827 2385 1828 2389
rect 1822 2384 1828 2385
rect 1862 2389 1868 2390
rect 1862 2385 1863 2389
rect 1867 2385 1868 2389
rect 1862 2384 1868 2385
rect 546 2375 552 2376
rect 546 2371 547 2375
rect 551 2371 552 2375
rect 546 2370 552 2371
rect 706 2375 712 2376
rect 706 2371 707 2375
rect 711 2371 712 2375
rect 706 2370 712 2371
rect 1166 2375 1172 2376
rect 1166 2371 1167 2375
rect 1171 2371 1172 2375
rect 1166 2370 1172 2371
rect 1822 2372 1828 2373
rect 486 2359 492 2360
rect 486 2355 487 2359
rect 491 2355 492 2359
rect 486 2354 492 2355
rect 386 2347 392 2348
rect 386 2343 387 2347
rect 391 2343 392 2347
rect 386 2342 392 2343
rect 488 2339 490 2354
rect 548 2348 550 2370
rect 646 2359 652 2360
rect 646 2355 647 2359
rect 651 2355 652 2359
rect 646 2354 652 2355
rect 546 2347 552 2348
rect 546 2343 547 2347
rect 551 2343 552 2347
rect 546 2342 552 2343
rect 648 2339 650 2354
rect 708 2348 710 2370
rect 790 2359 796 2360
rect 790 2355 791 2359
rect 795 2355 796 2359
rect 790 2354 796 2355
rect 926 2359 932 2360
rect 926 2355 927 2359
rect 931 2355 932 2359
rect 926 2354 932 2355
rect 1054 2359 1060 2360
rect 1054 2355 1055 2359
rect 1059 2355 1060 2359
rect 1054 2354 1060 2355
rect 706 2347 712 2348
rect 706 2343 707 2347
rect 711 2343 712 2347
rect 706 2342 712 2343
rect 792 2339 794 2354
rect 928 2339 930 2354
rect 1026 2347 1032 2348
rect 1026 2343 1027 2347
rect 1031 2343 1032 2347
rect 1026 2342 1032 2343
rect 263 2338 267 2339
rect 263 2333 267 2334
rect 327 2338 331 2339
rect 327 2333 331 2334
rect 407 2338 411 2339
rect 407 2333 411 2334
rect 487 2338 491 2339
rect 487 2333 491 2334
rect 543 2338 547 2339
rect 543 2333 547 2334
rect 647 2338 651 2339
rect 647 2333 651 2334
rect 679 2338 683 2339
rect 679 2333 683 2334
rect 791 2338 795 2339
rect 791 2333 795 2334
rect 807 2338 811 2339
rect 807 2333 811 2334
rect 927 2338 931 2339
rect 927 2333 931 2334
rect 218 2331 224 2332
rect 218 2327 219 2331
rect 223 2327 224 2331
rect 218 2326 224 2327
rect 264 2322 266 2333
rect 408 2322 410 2333
rect 438 2331 444 2332
rect 438 2327 439 2331
rect 443 2327 444 2331
rect 438 2326 444 2327
rect 142 2321 148 2322
rect 142 2317 143 2321
rect 147 2317 148 2321
rect 142 2316 148 2317
rect 262 2321 268 2322
rect 262 2317 263 2321
rect 267 2317 268 2321
rect 262 2316 268 2317
rect 406 2321 412 2322
rect 406 2317 407 2321
rect 411 2317 412 2321
rect 406 2316 412 2317
rect 110 2308 116 2309
rect 110 2304 111 2308
rect 115 2304 116 2308
rect 110 2303 116 2304
rect 110 2291 116 2292
rect 110 2287 111 2291
rect 115 2287 116 2291
rect 110 2286 116 2287
rect 386 2291 392 2292
rect 386 2287 387 2291
rect 391 2287 392 2291
rect 386 2286 392 2287
rect 112 2271 114 2286
rect 134 2281 140 2282
rect 134 2277 135 2281
rect 139 2277 140 2281
rect 134 2276 140 2277
rect 254 2281 260 2282
rect 254 2277 255 2281
rect 259 2277 260 2281
rect 254 2276 260 2277
rect 136 2271 138 2276
rect 256 2271 258 2276
rect 111 2270 115 2271
rect 111 2265 115 2266
rect 135 2270 139 2271
rect 135 2265 139 2266
rect 231 2270 235 2271
rect 231 2265 235 2266
rect 255 2270 259 2271
rect 255 2265 259 2266
rect 351 2270 355 2271
rect 351 2265 355 2266
rect 112 2250 114 2265
rect 136 2260 138 2265
rect 232 2260 234 2265
rect 352 2260 354 2265
rect 134 2259 140 2260
rect 134 2255 135 2259
rect 139 2255 140 2259
rect 134 2254 140 2255
rect 230 2259 236 2260
rect 230 2255 231 2259
rect 235 2255 236 2259
rect 230 2254 236 2255
rect 350 2259 356 2260
rect 350 2255 351 2259
rect 355 2255 356 2259
rect 350 2254 356 2255
rect 110 2249 116 2250
rect 110 2245 111 2249
rect 115 2245 116 2249
rect 110 2244 116 2245
rect 202 2235 208 2236
rect 110 2232 116 2233
rect 110 2228 111 2232
rect 115 2228 116 2232
rect 202 2231 203 2235
rect 207 2231 208 2235
rect 202 2230 208 2231
rect 298 2235 304 2236
rect 298 2231 299 2235
rect 303 2231 304 2235
rect 298 2230 304 2231
rect 110 2227 116 2228
rect 112 2199 114 2227
rect 142 2219 148 2220
rect 142 2215 143 2219
rect 147 2215 148 2219
rect 142 2214 148 2215
rect 144 2199 146 2214
rect 204 2208 206 2230
rect 238 2219 244 2220
rect 238 2215 239 2219
rect 243 2215 244 2219
rect 238 2214 244 2215
rect 202 2207 208 2208
rect 202 2203 203 2207
rect 207 2203 208 2207
rect 202 2202 208 2203
rect 240 2199 242 2214
rect 300 2208 302 2230
rect 358 2219 364 2220
rect 358 2215 359 2219
rect 363 2215 364 2219
rect 358 2214 364 2215
rect 298 2207 304 2208
rect 298 2203 299 2207
rect 303 2203 304 2207
rect 298 2202 304 2203
rect 360 2199 362 2214
rect 388 2208 390 2286
rect 398 2281 404 2282
rect 398 2277 399 2281
rect 403 2277 404 2281
rect 398 2276 404 2277
rect 400 2271 402 2276
rect 399 2270 403 2271
rect 399 2265 403 2266
rect 440 2252 442 2326
rect 544 2322 546 2333
rect 680 2322 682 2333
rect 808 2322 810 2333
rect 928 2322 930 2333
rect 542 2321 548 2322
rect 542 2317 543 2321
rect 547 2317 548 2321
rect 542 2316 548 2317
rect 678 2321 684 2322
rect 678 2317 679 2321
rect 683 2317 684 2321
rect 678 2316 684 2317
rect 806 2321 812 2322
rect 806 2317 807 2321
rect 811 2317 812 2321
rect 806 2316 812 2317
rect 926 2321 932 2322
rect 926 2317 927 2321
rect 931 2317 932 2321
rect 1028 2317 1030 2342
rect 1056 2339 1058 2354
rect 1168 2348 1170 2370
rect 1822 2368 1823 2372
rect 1827 2368 1828 2372
rect 1822 2367 1828 2368
rect 1862 2372 1868 2373
rect 1862 2368 1863 2372
rect 1867 2368 1868 2372
rect 1862 2367 1868 2368
rect 1182 2359 1188 2360
rect 1182 2355 1183 2359
rect 1187 2355 1188 2359
rect 1182 2354 1188 2355
rect 1310 2359 1316 2360
rect 1310 2355 1311 2359
rect 1315 2355 1316 2359
rect 1310 2354 1316 2355
rect 1438 2359 1444 2360
rect 1438 2355 1439 2359
rect 1443 2355 1444 2359
rect 1438 2354 1444 2355
rect 1166 2347 1172 2348
rect 1166 2343 1167 2347
rect 1171 2343 1172 2347
rect 1166 2342 1172 2343
rect 1184 2339 1186 2354
rect 1312 2339 1314 2354
rect 1440 2339 1442 2354
rect 1824 2339 1826 2367
rect 1864 2339 1866 2367
rect 2358 2359 2364 2360
rect 2358 2355 2359 2359
rect 2363 2355 2364 2359
rect 2358 2354 2364 2355
rect 2360 2339 2362 2354
rect 2392 2348 2394 2434
rect 2430 2429 2436 2430
rect 2430 2425 2431 2429
rect 2435 2425 2436 2429
rect 2430 2424 2436 2425
rect 2590 2429 2596 2430
rect 2590 2425 2591 2429
rect 2595 2425 2596 2429
rect 2590 2424 2596 2425
rect 2432 2411 2434 2424
rect 2592 2411 2594 2424
rect 2431 2410 2435 2411
rect 2431 2405 2435 2406
rect 2503 2410 2507 2411
rect 2503 2405 2507 2406
rect 2591 2410 2595 2411
rect 2591 2405 2595 2406
rect 2655 2410 2659 2411
rect 2655 2405 2659 2406
rect 2504 2400 2506 2405
rect 2656 2400 2658 2405
rect 2502 2399 2508 2400
rect 2502 2395 2503 2399
rect 2507 2395 2508 2399
rect 2502 2394 2508 2395
rect 2654 2399 2660 2400
rect 2654 2395 2655 2399
rect 2659 2395 2660 2399
rect 2654 2394 2660 2395
rect 2510 2379 2516 2380
rect 2510 2375 2511 2379
rect 2515 2375 2516 2379
rect 2510 2374 2516 2375
rect 2586 2375 2592 2376
rect 2512 2371 2514 2374
rect 2586 2371 2587 2375
rect 2591 2371 2592 2375
rect 2512 2369 2542 2371
rect 2586 2370 2592 2371
rect 2510 2359 2516 2360
rect 2510 2355 2511 2359
rect 2515 2355 2516 2359
rect 2510 2354 2516 2355
rect 2390 2347 2396 2348
rect 2390 2343 2391 2347
rect 2395 2343 2396 2347
rect 2390 2342 2396 2343
rect 2512 2339 2514 2354
rect 2540 2348 2542 2369
rect 2538 2347 2544 2348
rect 2538 2343 2539 2347
rect 2543 2343 2544 2347
rect 2538 2342 2544 2343
rect 1039 2338 1043 2339
rect 1039 2333 1043 2334
rect 1055 2338 1059 2339
rect 1055 2333 1059 2334
rect 1159 2338 1163 2339
rect 1159 2333 1163 2334
rect 1183 2338 1187 2339
rect 1183 2333 1187 2334
rect 1279 2338 1283 2339
rect 1279 2333 1283 2334
rect 1311 2338 1315 2339
rect 1311 2333 1315 2334
rect 1439 2338 1443 2339
rect 1439 2333 1443 2334
rect 1823 2338 1827 2339
rect 1823 2333 1827 2334
rect 1863 2338 1867 2339
rect 1863 2333 1867 2334
rect 2351 2338 2355 2339
rect 2351 2333 2355 2334
rect 2359 2338 2363 2339
rect 2359 2333 2363 2334
rect 2447 2338 2451 2339
rect 2447 2333 2451 2334
rect 2511 2338 2515 2339
rect 2511 2333 2515 2334
rect 2559 2338 2563 2339
rect 2559 2333 2563 2334
rect 1040 2322 1042 2333
rect 1102 2331 1108 2332
rect 1102 2327 1103 2331
rect 1107 2327 1108 2331
rect 1102 2326 1108 2327
rect 1038 2321 1044 2322
rect 1038 2317 1039 2321
rect 1043 2317 1044 2321
rect 926 2316 932 2317
rect 1027 2316 1031 2317
rect 1038 2316 1044 2317
rect 1027 2311 1031 2312
rect 1104 2308 1106 2326
rect 1160 2322 1162 2333
rect 1218 2331 1224 2332
rect 1218 2327 1219 2331
rect 1223 2327 1224 2331
rect 1218 2326 1224 2327
rect 1158 2321 1164 2322
rect 1158 2317 1159 2321
rect 1163 2317 1164 2321
rect 1158 2316 1164 2317
rect 1220 2308 1222 2326
rect 1280 2322 1282 2333
rect 1278 2321 1284 2322
rect 1278 2317 1279 2321
rect 1283 2317 1284 2321
rect 1227 2316 1231 2317
rect 1278 2316 1284 2317
rect 1227 2311 1231 2312
rect 1102 2307 1108 2308
rect 1102 2303 1103 2307
rect 1107 2303 1108 2307
rect 1102 2302 1108 2303
rect 1218 2307 1224 2308
rect 1218 2303 1219 2307
rect 1223 2303 1224 2307
rect 1228 2304 1230 2311
rect 1824 2309 1826 2333
rect 1864 2309 1866 2333
rect 2352 2322 2354 2333
rect 2418 2331 2424 2332
rect 2418 2327 2419 2331
rect 2423 2327 2424 2331
rect 2418 2326 2424 2327
rect 2350 2321 2356 2322
rect 2350 2317 2351 2321
rect 2355 2317 2356 2321
rect 2350 2316 2356 2317
rect 1822 2308 1828 2309
rect 1822 2304 1823 2308
rect 1827 2304 1828 2308
rect 1218 2302 1224 2303
rect 1226 2303 1232 2304
rect 1822 2303 1828 2304
rect 1862 2308 1868 2309
rect 1862 2304 1863 2308
rect 1867 2304 1868 2308
rect 2420 2304 2422 2326
rect 2448 2322 2450 2333
rect 2522 2331 2528 2332
rect 2522 2327 2523 2331
rect 2527 2327 2528 2331
rect 2522 2326 2528 2327
rect 2446 2321 2452 2322
rect 2446 2317 2447 2321
rect 2451 2317 2452 2321
rect 2446 2316 2452 2317
rect 2524 2304 2526 2326
rect 2560 2322 2562 2333
rect 2588 2332 2590 2370
rect 2662 2359 2668 2360
rect 2662 2355 2663 2359
rect 2667 2355 2668 2359
rect 2662 2354 2668 2355
rect 2664 2339 2666 2354
rect 2696 2348 2698 2434
rect 2758 2429 2764 2430
rect 2758 2425 2759 2429
rect 2763 2425 2764 2429
rect 2758 2424 2764 2425
rect 2934 2429 2940 2430
rect 2934 2425 2935 2429
rect 2939 2425 2940 2429
rect 2934 2424 2940 2425
rect 3110 2429 3116 2430
rect 3110 2425 3111 2429
rect 3115 2425 3116 2429
rect 3110 2424 3116 2425
rect 3286 2429 3292 2430
rect 3286 2425 3287 2429
rect 3291 2425 3292 2429
rect 3286 2424 3292 2425
rect 2760 2411 2762 2424
rect 2936 2411 2938 2424
rect 3112 2411 3114 2424
rect 3288 2411 3290 2424
rect 2759 2410 2763 2411
rect 2759 2405 2763 2406
rect 2807 2410 2811 2411
rect 2807 2405 2811 2406
rect 2935 2410 2939 2411
rect 2935 2405 2939 2406
rect 2967 2410 2971 2411
rect 2967 2405 2971 2406
rect 3111 2410 3115 2411
rect 3111 2405 3115 2406
rect 3135 2410 3139 2411
rect 3135 2405 3139 2406
rect 3287 2410 3291 2411
rect 3287 2405 3291 2406
rect 3303 2410 3307 2411
rect 3303 2405 3307 2406
rect 2808 2400 2810 2405
rect 2968 2400 2970 2405
rect 3136 2400 3138 2405
rect 3304 2400 3306 2405
rect 2806 2399 2812 2400
rect 2806 2395 2807 2399
rect 2811 2395 2812 2399
rect 2806 2394 2812 2395
rect 2966 2399 2972 2400
rect 2966 2395 2967 2399
rect 2971 2395 2972 2399
rect 2966 2394 2972 2395
rect 3134 2399 3140 2400
rect 3134 2395 3135 2399
rect 3139 2395 3140 2399
rect 3134 2394 3140 2395
rect 3302 2399 3308 2400
rect 3302 2395 3303 2399
rect 3307 2395 3308 2399
rect 3302 2394 3308 2395
rect 3312 2388 3314 2474
rect 3472 2470 3474 2481
rect 3548 2480 3550 2514
rect 3574 2512 3575 2516
rect 3579 2512 3580 2516
rect 3574 2511 3580 2512
rect 3576 2487 3578 2511
rect 3575 2486 3579 2487
rect 3575 2481 3579 2482
rect 3546 2479 3552 2480
rect 3546 2475 3547 2479
rect 3551 2475 3552 2479
rect 3546 2474 3552 2475
rect 3470 2469 3476 2470
rect 3470 2465 3471 2469
rect 3475 2465 3476 2469
rect 3470 2464 3476 2465
rect 3576 2457 3578 2481
rect 3574 2456 3580 2457
rect 3574 2452 3575 2456
rect 3579 2452 3580 2456
rect 3574 2451 3580 2452
rect 3574 2439 3580 2440
rect 3574 2435 3575 2439
rect 3579 2435 3580 2439
rect 3574 2434 3580 2435
rect 3462 2429 3468 2430
rect 3462 2425 3463 2429
rect 3467 2425 3468 2429
rect 3462 2424 3468 2425
rect 3464 2411 3466 2424
rect 3510 2423 3516 2424
rect 3510 2419 3511 2423
rect 3515 2419 3516 2423
rect 3510 2418 3516 2419
rect 3463 2410 3467 2411
rect 3463 2405 3467 2406
rect 3471 2410 3475 2411
rect 3471 2405 3475 2406
rect 3472 2400 3474 2405
rect 3470 2399 3476 2400
rect 3470 2395 3471 2399
rect 3475 2395 3476 2399
rect 3470 2394 3476 2395
rect 3310 2387 3316 2388
rect 3310 2383 3311 2387
rect 3315 2383 3316 2387
rect 3310 2382 3316 2383
rect 3294 2375 3300 2376
rect 3294 2371 3295 2375
rect 3299 2371 3300 2375
rect 3294 2370 3300 2371
rect 2814 2359 2820 2360
rect 2814 2355 2815 2359
rect 2819 2355 2820 2359
rect 2814 2354 2820 2355
rect 2974 2359 2980 2360
rect 2974 2355 2975 2359
rect 2979 2355 2980 2359
rect 2974 2354 2980 2355
rect 3142 2359 3148 2360
rect 3142 2355 3143 2359
rect 3147 2355 3148 2359
rect 3142 2354 3148 2355
rect 2694 2347 2700 2348
rect 2694 2343 2695 2347
rect 2699 2343 2700 2347
rect 2694 2342 2700 2343
rect 2816 2339 2818 2354
rect 2958 2339 2964 2340
rect 2976 2339 2978 2354
rect 3144 2339 3146 2354
rect 2663 2338 2667 2339
rect 2663 2333 2667 2334
rect 2703 2338 2707 2339
rect 2703 2333 2707 2334
rect 2815 2338 2819 2339
rect 2815 2333 2819 2334
rect 2879 2338 2883 2339
rect 2958 2335 2959 2339
rect 2963 2335 2964 2339
rect 2958 2334 2964 2335
rect 2975 2338 2979 2339
rect 2879 2333 2883 2334
rect 2586 2331 2592 2332
rect 2586 2327 2587 2331
rect 2591 2327 2592 2331
rect 2586 2326 2592 2327
rect 2704 2322 2706 2333
rect 2880 2322 2882 2333
rect 2558 2321 2564 2322
rect 2558 2317 2559 2321
rect 2563 2317 2564 2321
rect 2558 2316 2564 2317
rect 2702 2321 2708 2322
rect 2702 2317 2703 2321
rect 2707 2317 2708 2321
rect 2702 2316 2708 2317
rect 2878 2321 2884 2322
rect 2878 2317 2879 2321
rect 2883 2317 2884 2321
rect 2878 2316 2884 2317
rect 2960 2304 2962 2334
rect 2975 2333 2979 2334
rect 3079 2338 3083 2339
rect 3079 2333 3083 2334
rect 3143 2338 3147 2339
rect 3143 2333 3147 2334
rect 3287 2338 3291 2339
rect 3287 2333 3291 2334
rect 3080 2322 3082 2333
rect 3150 2331 3156 2332
rect 3150 2327 3151 2331
rect 3155 2327 3156 2331
rect 3150 2326 3156 2327
rect 3078 2321 3084 2322
rect 3078 2317 3079 2321
rect 3083 2317 3084 2321
rect 3078 2316 3084 2317
rect 3152 2304 3154 2326
rect 3288 2322 3290 2333
rect 3296 2332 3298 2370
rect 3310 2359 3316 2360
rect 3310 2355 3311 2359
rect 3315 2355 3316 2359
rect 3310 2354 3316 2355
rect 3478 2359 3484 2360
rect 3478 2355 3479 2359
rect 3483 2355 3484 2359
rect 3478 2354 3484 2355
rect 3312 2339 3314 2354
rect 3370 2347 3376 2348
rect 3370 2343 3371 2347
rect 3375 2343 3376 2347
rect 3370 2342 3376 2343
rect 3311 2338 3315 2339
rect 3311 2333 3315 2334
rect 3294 2331 3300 2332
rect 3294 2327 3295 2331
rect 3299 2327 3300 2331
rect 3294 2326 3300 2327
rect 3286 2321 3292 2322
rect 3286 2317 3287 2321
rect 3291 2317 3292 2321
rect 3286 2316 3292 2317
rect 1862 2303 1868 2304
rect 2418 2303 2424 2304
rect 1226 2299 1227 2303
rect 1231 2299 1232 2303
rect 1226 2298 1232 2299
rect 2418 2299 2419 2303
rect 2423 2299 2424 2303
rect 2418 2298 2424 2299
rect 2522 2303 2528 2304
rect 2522 2299 2523 2303
rect 2527 2299 2528 2303
rect 2522 2298 2528 2299
rect 2958 2303 2964 2304
rect 2958 2299 2959 2303
rect 2963 2299 2964 2303
rect 2958 2298 2964 2299
rect 3150 2303 3156 2304
rect 3150 2299 3151 2303
rect 3155 2299 3156 2303
rect 3150 2298 3156 2299
rect 1822 2291 1828 2292
rect 1822 2287 1823 2291
rect 1827 2287 1828 2291
rect 1822 2286 1828 2287
rect 1862 2291 1868 2292
rect 1862 2287 1863 2291
rect 1867 2287 1868 2291
rect 1862 2286 1868 2287
rect 2946 2291 2952 2292
rect 2946 2287 2947 2291
rect 2951 2287 2952 2291
rect 2946 2286 2952 2287
rect 534 2281 540 2282
rect 534 2277 535 2281
rect 539 2277 540 2281
rect 534 2276 540 2277
rect 670 2281 676 2282
rect 670 2277 671 2281
rect 675 2277 676 2281
rect 670 2276 676 2277
rect 798 2281 804 2282
rect 798 2277 799 2281
rect 803 2277 804 2281
rect 798 2276 804 2277
rect 918 2281 924 2282
rect 918 2277 919 2281
rect 923 2277 924 2281
rect 918 2276 924 2277
rect 1030 2281 1036 2282
rect 1030 2277 1031 2281
rect 1035 2277 1036 2281
rect 1030 2276 1036 2277
rect 1150 2281 1156 2282
rect 1150 2277 1151 2281
rect 1155 2277 1156 2281
rect 1150 2276 1156 2277
rect 1270 2281 1276 2282
rect 1270 2277 1271 2281
rect 1275 2277 1276 2281
rect 1270 2276 1276 2277
rect 536 2271 538 2276
rect 672 2271 674 2276
rect 800 2271 802 2276
rect 920 2271 922 2276
rect 1032 2271 1034 2276
rect 1152 2271 1154 2276
rect 1272 2271 1274 2276
rect 1824 2271 1826 2286
rect 1864 2271 1866 2286
rect 2342 2281 2348 2282
rect 2342 2277 2343 2281
rect 2347 2277 2348 2281
rect 2342 2276 2348 2277
rect 2438 2281 2444 2282
rect 2438 2277 2439 2281
rect 2443 2277 2444 2281
rect 2438 2276 2444 2277
rect 2550 2281 2556 2282
rect 2550 2277 2551 2281
rect 2555 2277 2556 2281
rect 2550 2276 2556 2277
rect 2694 2281 2700 2282
rect 2694 2277 2695 2281
rect 2699 2277 2700 2281
rect 2694 2276 2700 2277
rect 2870 2281 2876 2282
rect 2870 2277 2871 2281
rect 2875 2277 2876 2281
rect 2870 2276 2876 2277
rect 2344 2271 2346 2276
rect 2374 2275 2380 2276
rect 2374 2271 2375 2275
rect 2379 2271 2380 2275
rect 2440 2271 2442 2276
rect 2552 2271 2554 2276
rect 2696 2271 2698 2276
rect 2872 2271 2874 2276
rect 471 2270 475 2271
rect 471 2265 475 2266
rect 535 2270 539 2271
rect 535 2265 539 2266
rect 591 2270 595 2271
rect 591 2265 595 2266
rect 671 2270 675 2271
rect 671 2265 675 2266
rect 711 2270 715 2271
rect 711 2265 715 2266
rect 799 2270 803 2271
rect 799 2265 803 2266
rect 823 2270 827 2271
rect 823 2265 827 2266
rect 919 2270 923 2271
rect 919 2265 923 2266
rect 935 2270 939 2271
rect 935 2265 939 2266
rect 1031 2270 1035 2271
rect 1031 2265 1035 2266
rect 1055 2270 1059 2271
rect 1055 2265 1059 2266
rect 1151 2270 1155 2271
rect 1151 2265 1155 2266
rect 1175 2270 1179 2271
rect 1175 2265 1179 2266
rect 1271 2270 1275 2271
rect 1271 2265 1275 2266
rect 1823 2270 1827 2271
rect 1823 2265 1827 2266
rect 1863 2270 1867 2271
rect 1863 2265 1867 2266
rect 2335 2270 2339 2271
rect 2335 2265 2339 2266
rect 2343 2270 2347 2271
rect 2374 2270 2380 2271
rect 2439 2270 2443 2271
rect 2343 2265 2347 2266
rect 472 2260 474 2265
rect 592 2260 594 2265
rect 712 2260 714 2265
rect 824 2260 826 2265
rect 936 2260 938 2265
rect 1056 2260 1058 2265
rect 1176 2260 1178 2265
rect 470 2259 476 2260
rect 470 2255 471 2259
rect 475 2255 476 2259
rect 470 2254 476 2255
rect 590 2259 596 2260
rect 590 2255 591 2259
rect 595 2255 596 2259
rect 590 2254 596 2255
rect 710 2259 716 2260
rect 710 2255 711 2259
rect 715 2255 716 2259
rect 710 2254 716 2255
rect 822 2259 828 2260
rect 822 2255 823 2259
rect 827 2255 828 2259
rect 822 2254 828 2255
rect 934 2259 940 2260
rect 934 2255 935 2259
rect 939 2255 940 2259
rect 934 2254 940 2255
rect 1054 2259 1060 2260
rect 1054 2255 1055 2259
rect 1059 2255 1060 2259
rect 1054 2254 1060 2255
rect 1174 2259 1180 2260
rect 1174 2255 1175 2259
rect 1179 2255 1180 2259
rect 1174 2254 1180 2255
rect 438 2251 444 2252
rect 438 2247 439 2251
rect 443 2247 444 2251
rect 1824 2250 1826 2265
rect 1864 2250 1866 2265
rect 2336 2260 2338 2265
rect 2334 2259 2340 2260
rect 2334 2255 2335 2259
rect 2339 2255 2340 2259
rect 2334 2254 2340 2255
rect 438 2246 444 2247
rect 1822 2249 1828 2250
rect 1822 2245 1823 2249
rect 1827 2245 1828 2249
rect 1822 2244 1828 2245
rect 1862 2249 1868 2250
rect 1862 2245 1863 2249
rect 1867 2245 1868 2249
rect 1862 2244 1868 2245
rect 538 2235 544 2236
rect 538 2231 539 2235
rect 543 2231 544 2235
rect 538 2230 544 2231
rect 778 2235 784 2236
rect 778 2231 779 2235
rect 783 2231 784 2235
rect 778 2230 784 2231
rect 1138 2235 1144 2236
rect 1138 2231 1139 2235
rect 1143 2231 1144 2235
rect 1138 2230 1144 2231
rect 1146 2235 1152 2236
rect 1146 2231 1147 2235
rect 1151 2231 1152 2235
rect 1146 2230 1152 2231
rect 1822 2232 1828 2233
rect 478 2219 484 2220
rect 478 2215 479 2219
rect 483 2215 484 2219
rect 478 2214 484 2215
rect 386 2207 392 2208
rect 386 2203 387 2207
rect 391 2203 392 2207
rect 386 2202 392 2203
rect 480 2199 482 2214
rect 540 2208 542 2230
rect 598 2219 604 2220
rect 598 2215 599 2219
rect 603 2215 604 2219
rect 598 2214 604 2215
rect 718 2219 724 2220
rect 718 2215 719 2219
rect 723 2215 724 2219
rect 718 2214 724 2215
rect 538 2207 544 2208
rect 538 2203 539 2207
rect 543 2203 544 2207
rect 538 2202 544 2203
rect 600 2199 602 2214
rect 630 2207 636 2208
rect 630 2203 631 2207
rect 635 2203 636 2207
rect 630 2202 636 2203
rect 111 2198 115 2199
rect 111 2193 115 2194
rect 143 2198 147 2199
rect 143 2193 147 2194
rect 239 2198 243 2199
rect 239 2193 243 2194
rect 247 2198 251 2199
rect 247 2193 251 2194
rect 359 2198 363 2199
rect 359 2193 363 2194
rect 383 2198 387 2199
rect 383 2193 387 2194
rect 479 2198 483 2199
rect 479 2193 483 2194
rect 519 2198 523 2199
rect 519 2193 523 2194
rect 599 2198 603 2199
rect 599 2193 603 2194
rect 112 2169 114 2193
rect 144 2182 146 2193
rect 248 2182 250 2193
rect 384 2182 386 2193
rect 426 2191 432 2192
rect 426 2187 427 2191
rect 431 2187 432 2191
rect 426 2186 432 2187
rect 142 2181 148 2182
rect 142 2177 143 2181
rect 147 2177 148 2181
rect 142 2176 148 2177
rect 246 2181 252 2182
rect 246 2177 247 2181
rect 251 2177 252 2181
rect 246 2176 252 2177
rect 382 2181 388 2182
rect 382 2177 383 2181
rect 387 2177 388 2181
rect 382 2176 388 2177
rect 110 2168 116 2169
rect 110 2164 111 2168
rect 115 2164 116 2168
rect 110 2163 116 2164
rect 110 2151 116 2152
rect 110 2147 111 2151
rect 115 2147 116 2151
rect 110 2146 116 2147
rect 112 2123 114 2146
rect 134 2141 140 2142
rect 134 2137 135 2141
rect 139 2137 140 2141
rect 134 2136 140 2137
rect 238 2141 244 2142
rect 238 2137 239 2141
rect 243 2137 244 2141
rect 238 2136 244 2137
rect 374 2141 380 2142
rect 374 2137 375 2141
rect 379 2137 380 2141
rect 374 2136 380 2137
rect 136 2123 138 2136
rect 240 2123 242 2136
rect 270 2135 276 2136
rect 270 2131 271 2135
rect 275 2131 276 2135
rect 270 2130 276 2131
rect 111 2122 115 2123
rect 111 2117 115 2118
rect 135 2122 139 2123
rect 135 2117 139 2118
rect 231 2122 235 2123
rect 231 2117 235 2118
rect 239 2122 243 2123
rect 239 2117 243 2118
rect 112 2102 114 2117
rect 136 2112 138 2117
rect 232 2112 234 2117
rect 134 2111 140 2112
rect 134 2107 135 2111
rect 139 2107 140 2111
rect 134 2106 140 2107
rect 230 2111 236 2112
rect 230 2107 231 2111
rect 235 2107 236 2111
rect 230 2106 236 2107
rect 110 2101 116 2102
rect 110 2097 111 2101
rect 115 2097 116 2101
rect 110 2096 116 2097
rect 202 2087 208 2088
rect 110 2084 116 2085
rect 110 2080 111 2084
rect 115 2080 116 2084
rect 202 2083 203 2087
rect 207 2083 208 2087
rect 202 2082 208 2083
rect 110 2079 116 2080
rect 112 2043 114 2079
rect 142 2071 148 2072
rect 142 2067 143 2071
rect 147 2067 148 2071
rect 142 2066 148 2067
rect 144 2043 146 2066
rect 204 2060 206 2082
rect 238 2071 244 2072
rect 238 2067 239 2071
rect 243 2067 244 2071
rect 238 2066 244 2067
rect 202 2059 208 2060
rect 202 2055 203 2059
rect 207 2055 208 2059
rect 202 2054 208 2055
rect 240 2043 242 2066
rect 272 2060 274 2130
rect 376 2123 378 2136
rect 359 2122 363 2123
rect 359 2117 363 2118
rect 375 2122 379 2123
rect 375 2117 379 2118
rect 360 2112 362 2117
rect 358 2111 364 2112
rect 358 2107 359 2111
rect 363 2107 364 2111
rect 358 2106 364 2107
rect 428 2104 430 2186
rect 520 2182 522 2193
rect 518 2181 524 2182
rect 518 2177 519 2181
rect 523 2177 524 2181
rect 518 2176 524 2177
rect 632 2164 634 2202
rect 720 2199 722 2214
rect 780 2208 782 2230
rect 830 2219 836 2220
rect 830 2215 831 2219
rect 835 2215 836 2219
rect 830 2214 836 2215
rect 942 2219 948 2220
rect 942 2215 943 2219
rect 947 2215 948 2219
rect 942 2214 948 2215
rect 1062 2219 1068 2220
rect 1062 2215 1063 2219
rect 1067 2215 1068 2219
rect 1062 2214 1068 2215
rect 778 2207 784 2208
rect 778 2203 779 2207
rect 783 2203 784 2207
rect 778 2202 784 2203
rect 832 2199 834 2214
rect 944 2199 946 2214
rect 970 2207 976 2208
rect 970 2203 971 2207
rect 975 2203 976 2207
rect 970 2202 976 2203
rect 655 2198 659 2199
rect 655 2193 659 2194
rect 719 2198 723 2199
rect 719 2193 723 2194
rect 783 2198 787 2199
rect 783 2193 787 2194
rect 831 2198 835 2199
rect 831 2193 835 2194
rect 911 2198 915 2199
rect 911 2193 915 2194
rect 943 2198 947 2199
rect 943 2193 947 2194
rect 656 2182 658 2193
rect 784 2182 786 2193
rect 912 2182 914 2193
rect 654 2181 660 2182
rect 654 2177 655 2181
rect 659 2177 660 2181
rect 654 2176 660 2177
rect 782 2181 788 2182
rect 782 2177 783 2181
rect 787 2177 788 2181
rect 782 2176 788 2177
rect 910 2181 916 2182
rect 910 2177 911 2181
rect 915 2177 916 2181
rect 910 2176 916 2177
rect 972 2168 974 2202
rect 978 2199 984 2200
rect 1064 2199 1066 2214
rect 1140 2208 1142 2230
rect 1148 2216 1150 2230
rect 1822 2228 1823 2232
rect 1827 2228 1828 2232
rect 1822 2227 1828 2228
rect 1862 2232 1868 2233
rect 1862 2228 1863 2232
rect 1867 2228 1868 2232
rect 1862 2227 1868 2228
rect 1182 2219 1188 2220
rect 1146 2215 1152 2216
rect 1146 2211 1147 2215
rect 1151 2211 1152 2215
rect 1182 2215 1183 2219
rect 1187 2215 1188 2219
rect 1182 2214 1188 2215
rect 1146 2210 1152 2211
rect 1138 2207 1144 2208
rect 1138 2203 1139 2207
rect 1143 2203 1144 2207
rect 1138 2202 1144 2203
rect 1184 2199 1186 2214
rect 1824 2199 1826 2227
rect 1864 2203 1866 2227
rect 2342 2219 2348 2220
rect 2342 2215 2343 2219
rect 2347 2215 2348 2219
rect 2342 2214 2348 2215
rect 2344 2203 2346 2214
rect 2376 2208 2378 2270
rect 2439 2265 2443 2266
rect 2447 2270 2451 2271
rect 2447 2265 2451 2266
rect 2551 2270 2555 2271
rect 2551 2265 2555 2266
rect 2583 2270 2587 2271
rect 2583 2265 2587 2266
rect 2695 2270 2699 2271
rect 2695 2265 2699 2266
rect 2735 2270 2739 2271
rect 2735 2265 2739 2266
rect 2871 2270 2875 2271
rect 2871 2265 2875 2266
rect 2911 2270 2915 2271
rect 2911 2265 2915 2266
rect 2448 2260 2450 2265
rect 2584 2260 2586 2265
rect 2736 2260 2738 2265
rect 2912 2260 2914 2265
rect 2446 2259 2452 2260
rect 2446 2255 2447 2259
rect 2451 2255 2452 2259
rect 2446 2254 2452 2255
rect 2582 2259 2588 2260
rect 2582 2255 2583 2259
rect 2587 2255 2588 2259
rect 2582 2254 2588 2255
rect 2734 2259 2740 2260
rect 2734 2255 2735 2259
rect 2739 2255 2740 2259
rect 2734 2254 2740 2255
rect 2910 2259 2916 2260
rect 2910 2255 2911 2259
rect 2915 2255 2916 2259
rect 2910 2254 2916 2255
rect 2566 2235 2572 2236
rect 2566 2231 2567 2235
rect 2571 2231 2572 2235
rect 2566 2230 2572 2231
rect 2574 2235 2580 2236
rect 2574 2231 2575 2235
rect 2579 2231 2580 2235
rect 2574 2230 2580 2231
rect 2726 2235 2732 2236
rect 2726 2231 2727 2235
rect 2731 2231 2732 2235
rect 2726 2230 2732 2231
rect 2454 2219 2460 2220
rect 2454 2215 2455 2219
rect 2459 2215 2460 2219
rect 2454 2214 2460 2215
rect 2374 2207 2380 2208
rect 2374 2203 2375 2207
rect 2379 2203 2380 2207
rect 2456 2203 2458 2214
rect 2568 2208 2570 2230
rect 2566 2207 2572 2208
rect 2566 2203 2567 2207
rect 2571 2203 2572 2207
rect 1863 2202 1867 2203
rect 978 2195 979 2199
rect 983 2195 984 2199
rect 978 2194 984 2195
rect 1031 2198 1035 2199
rect 970 2167 976 2168
rect 630 2163 636 2164
rect 630 2159 631 2163
rect 635 2159 636 2163
rect 970 2163 971 2167
rect 975 2163 976 2167
rect 980 2164 982 2194
rect 1031 2193 1035 2194
rect 1063 2198 1067 2199
rect 1063 2193 1067 2194
rect 1159 2198 1163 2199
rect 1159 2193 1163 2194
rect 1183 2198 1187 2199
rect 1183 2193 1187 2194
rect 1287 2198 1291 2199
rect 1287 2193 1291 2194
rect 1823 2198 1827 2199
rect 1863 2197 1867 2198
rect 2255 2202 2259 2203
rect 2255 2197 2259 2198
rect 2343 2202 2347 2203
rect 2374 2202 2380 2203
rect 2439 2202 2443 2203
rect 2343 2197 2347 2198
rect 2439 2197 2443 2198
rect 2455 2202 2459 2203
rect 2455 2197 2459 2198
rect 2551 2202 2555 2203
rect 2566 2202 2572 2203
rect 2551 2197 2555 2198
rect 1823 2193 1827 2194
rect 1032 2182 1034 2193
rect 1160 2182 1162 2193
rect 1230 2191 1236 2192
rect 1230 2187 1231 2191
rect 1235 2187 1236 2191
rect 1230 2186 1236 2187
rect 1030 2181 1036 2182
rect 1030 2177 1031 2181
rect 1035 2177 1036 2181
rect 1030 2176 1036 2177
rect 1158 2181 1164 2182
rect 1158 2177 1159 2181
rect 1163 2177 1164 2181
rect 1158 2176 1164 2177
rect 1232 2164 1234 2186
rect 1288 2182 1290 2193
rect 1286 2181 1292 2182
rect 1286 2177 1287 2181
rect 1291 2177 1292 2181
rect 1286 2176 1292 2177
rect 1824 2169 1826 2193
rect 1864 2173 1866 2197
rect 2256 2186 2258 2197
rect 2322 2195 2328 2196
rect 2322 2191 2323 2195
rect 2327 2191 2328 2195
rect 2322 2190 2328 2191
rect 2254 2185 2260 2186
rect 2254 2181 2255 2185
rect 2259 2181 2260 2185
rect 2254 2180 2260 2181
rect 1862 2172 1868 2173
rect 1822 2168 1828 2169
rect 1822 2164 1823 2168
rect 1827 2164 1828 2168
rect 1862 2168 1863 2172
rect 1867 2168 1868 2172
rect 2324 2168 2326 2190
rect 2344 2186 2346 2197
rect 2410 2195 2416 2196
rect 2410 2191 2411 2195
rect 2415 2191 2416 2195
rect 2410 2190 2416 2191
rect 2342 2185 2348 2186
rect 2342 2181 2343 2185
rect 2347 2181 2348 2185
rect 2342 2180 2348 2181
rect 2412 2168 2414 2190
rect 2440 2186 2442 2197
rect 2514 2195 2520 2196
rect 2514 2191 2515 2195
rect 2519 2191 2520 2195
rect 2514 2190 2520 2191
rect 2438 2185 2444 2186
rect 2438 2181 2439 2185
rect 2443 2181 2444 2185
rect 2438 2180 2444 2181
rect 2516 2168 2518 2190
rect 2552 2186 2554 2197
rect 2576 2196 2578 2230
rect 2590 2219 2596 2220
rect 2590 2215 2591 2219
rect 2595 2215 2596 2219
rect 2590 2214 2596 2215
rect 2592 2203 2594 2214
rect 2591 2202 2595 2203
rect 2591 2197 2595 2198
rect 2695 2202 2699 2203
rect 2695 2197 2699 2198
rect 2574 2195 2580 2196
rect 2574 2191 2575 2195
rect 2579 2191 2580 2195
rect 2574 2190 2580 2191
rect 2696 2186 2698 2197
rect 2728 2196 2730 2230
rect 2742 2219 2748 2220
rect 2742 2215 2743 2219
rect 2747 2215 2748 2219
rect 2742 2214 2748 2215
rect 2918 2219 2924 2220
rect 2918 2215 2919 2219
rect 2923 2215 2924 2219
rect 2918 2214 2924 2215
rect 2744 2203 2746 2214
rect 2920 2203 2922 2214
rect 2948 2208 2950 2286
rect 3070 2281 3076 2282
rect 3070 2277 3071 2281
rect 3075 2277 3076 2281
rect 3070 2276 3076 2277
rect 3278 2281 3284 2282
rect 3278 2277 3279 2281
rect 3283 2277 3284 2281
rect 3278 2276 3284 2277
rect 3072 2271 3074 2276
rect 3280 2271 3282 2276
rect 3071 2270 3075 2271
rect 3071 2265 3075 2266
rect 3103 2270 3107 2271
rect 3103 2265 3107 2266
rect 3279 2270 3283 2271
rect 3279 2265 3283 2266
rect 3303 2270 3307 2271
rect 3303 2265 3307 2266
rect 3104 2260 3106 2265
rect 3304 2260 3306 2265
rect 3102 2259 3108 2260
rect 3102 2255 3103 2259
rect 3107 2255 3108 2259
rect 3102 2254 3108 2255
rect 3302 2259 3308 2260
rect 3302 2255 3303 2259
rect 3307 2255 3308 2259
rect 3302 2254 3308 2255
rect 3372 2252 3374 2342
rect 3480 2339 3482 2354
rect 3512 2348 3514 2418
rect 3576 2411 3578 2434
rect 3575 2410 3579 2411
rect 3575 2405 3579 2406
rect 3576 2390 3578 2405
rect 3574 2389 3580 2390
rect 3574 2385 3575 2389
rect 3579 2385 3580 2389
rect 3574 2384 3580 2385
rect 3538 2375 3544 2376
rect 3538 2371 3539 2375
rect 3543 2371 3544 2375
rect 3538 2370 3544 2371
rect 3574 2372 3580 2373
rect 3510 2347 3516 2348
rect 3510 2343 3511 2347
rect 3515 2343 3516 2347
rect 3510 2342 3516 2343
rect 3479 2338 3483 2339
rect 3479 2333 3483 2334
rect 3487 2338 3491 2339
rect 3487 2333 3491 2334
rect 3488 2322 3490 2333
rect 3540 2332 3542 2370
rect 3574 2368 3575 2372
rect 3579 2368 3580 2372
rect 3574 2367 3580 2368
rect 3576 2339 3578 2367
rect 3575 2338 3579 2339
rect 3575 2333 3579 2334
rect 3538 2331 3544 2332
rect 3538 2327 3539 2331
rect 3543 2327 3544 2331
rect 3538 2326 3544 2327
rect 3486 2321 3492 2322
rect 3486 2317 3487 2321
rect 3491 2317 3492 2321
rect 3486 2316 3492 2317
rect 3576 2309 3578 2333
rect 3574 2308 3580 2309
rect 3574 2304 3575 2308
rect 3579 2304 3580 2308
rect 3574 2303 3580 2304
rect 3574 2291 3580 2292
rect 3574 2287 3575 2291
rect 3579 2287 3580 2291
rect 3574 2286 3580 2287
rect 3478 2281 3484 2282
rect 3478 2277 3479 2281
rect 3483 2277 3484 2281
rect 3478 2276 3484 2277
rect 3480 2271 3482 2276
rect 3518 2275 3524 2276
rect 3518 2271 3519 2275
rect 3523 2271 3524 2275
rect 3576 2271 3578 2286
rect 3479 2270 3483 2271
rect 3518 2270 3524 2271
rect 3575 2270 3579 2271
rect 3479 2265 3483 2266
rect 3480 2260 3482 2265
rect 3478 2259 3484 2260
rect 3478 2255 3479 2259
rect 3483 2255 3484 2259
rect 3478 2254 3484 2255
rect 3370 2251 3376 2252
rect 3370 2247 3371 2251
rect 3375 2247 3376 2251
rect 3370 2246 3376 2247
rect 3014 2235 3020 2236
rect 3014 2231 3015 2235
rect 3019 2231 3020 2235
rect 3014 2230 3020 2231
rect 3022 2235 3028 2236
rect 3022 2231 3023 2235
rect 3027 2231 3028 2235
rect 3022 2230 3028 2231
rect 3016 2208 3018 2230
rect 3024 2216 3026 2230
rect 3110 2219 3116 2220
rect 3022 2215 3028 2216
rect 3022 2211 3023 2215
rect 3027 2211 3028 2215
rect 3110 2215 3111 2219
rect 3115 2215 3116 2219
rect 3110 2214 3116 2215
rect 3310 2219 3316 2220
rect 3310 2215 3311 2219
rect 3315 2215 3316 2219
rect 3310 2214 3316 2215
rect 3486 2219 3492 2220
rect 3486 2215 3487 2219
rect 3491 2215 3492 2219
rect 3486 2214 3492 2215
rect 3022 2210 3028 2211
rect 2946 2207 2952 2208
rect 2946 2203 2947 2207
rect 2951 2203 2952 2207
rect 2743 2202 2747 2203
rect 2743 2197 2747 2198
rect 2871 2202 2875 2203
rect 2871 2197 2875 2198
rect 2919 2202 2923 2203
rect 2946 2202 2952 2203
rect 3014 2207 3020 2208
rect 3014 2203 3015 2207
rect 3019 2203 3020 2207
rect 3112 2203 3114 2214
rect 3312 2203 3314 2214
rect 3342 2207 3348 2208
rect 3342 2203 3343 2207
rect 3347 2203 3348 2207
rect 3488 2203 3490 2214
rect 3520 2208 3522 2270
rect 3575 2265 3579 2266
rect 3576 2250 3578 2265
rect 3574 2249 3580 2250
rect 3574 2245 3575 2249
rect 3579 2245 3580 2249
rect 3574 2244 3580 2245
rect 3546 2235 3552 2236
rect 3546 2231 3547 2235
rect 3551 2231 3552 2235
rect 3546 2230 3552 2231
rect 3574 2232 3580 2233
rect 3518 2207 3524 2208
rect 3518 2203 3519 2207
rect 3523 2203 3524 2207
rect 3014 2202 3020 2203
rect 3071 2202 3075 2203
rect 2919 2197 2923 2198
rect 3071 2197 3075 2198
rect 3111 2202 3115 2203
rect 3111 2197 3115 2198
rect 3287 2202 3291 2203
rect 3287 2197 3291 2198
rect 3311 2202 3315 2203
rect 3342 2202 3348 2203
rect 3487 2202 3491 2203
rect 3518 2202 3524 2203
rect 3311 2197 3315 2198
rect 2726 2195 2732 2196
rect 2726 2191 2727 2195
rect 2731 2191 2732 2195
rect 2726 2190 2732 2191
rect 2822 2195 2828 2196
rect 2822 2191 2823 2195
rect 2827 2191 2828 2195
rect 2822 2190 2828 2191
rect 2550 2185 2556 2186
rect 2550 2181 2551 2185
rect 2555 2181 2556 2185
rect 2550 2180 2556 2181
rect 2694 2185 2700 2186
rect 2694 2181 2695 2185
rect 2699 2181 2700 2185
rect 2694 2180 2700 2181
rect 2824 2172 2826 2190
rect 2872 2186 2874 2197
rect 3072 2186 3074 2197
rect 3288 2186 3290 2197
rect 2870 2185 2876 2186
rect 2870 2181 2871 2185
rect 2875 2181 2876 2185
rect 2870 2180 2876 2181
rect 3070 2185 3076 2186
rect 3070 2181 3071 2185
rect 3075 2181 3076 2185
rect 3070 2180 3076 2181
rect 3286 2185 3292 2186
rect 3286 2181 3287 2185
rect 3291 2181 3292 2185
rect 3286 2180 3292 2181
rect 2822 2171 2828 2172
rect 1862 2167 1868 2168
rect 2322 2167 2328 2168
rect 970 2162 976 2163
rect 978 2163 984 2164
rect 630 2158 636 2159
rect 978 2159 979 2163
rect 983 2159 984 2163
rect 978 2158 984 2159
rect 1230 2163 1236 2164
rect 1822 2163 1828 2164
rect 2322 2163 2323 2167
rect 2327 2163 2328 2167
rect 1230 2159 1231 2163
rect 1235 2159 1236 2163
rect 2322 2162 2328 2163
rect 2410 2167 2416 2168
rect 2410 2163 2411 2167
rect 2415 2163 2416 2167
rect 2410 2162 2416 2163
rect 2514 2167 2520 2168
rect 2514 2163 2515 2167
rect 2519 2163 2520 2167
rect 2822 2167 2823 2171
rect 2827 2167 2828 2171
rect 2822 2166 2828 2167
rect 2514 2162 2520 2163
rect 1230 2158 1236 2159
rect 1862 2155 1868 2156
rect 1822 2151 1828 2152
rect 1822 2147 1823 2151
rect 1827 2147 1828 2151
rect 1862 2151 1863 2155
rect 1867 2151 1868 2155
rect 1862 2150 1868 2151
rect 2342 2155 2348 2156
rect 2342 2151 2343 2155
rect 2347 2151 2348 2155
rect 2342 2150 2348 2151
rect 3198 2155 3204 2156
rect 3198 2151 3199 2155
rect 3203 2151 3204 2155
rect 3198 2150 3204 2151
rect 1822 2146 1828 2147
rect 510 2141 516 2142
rect 510 2137 511 2141
rect 515 2137 516 2141
rect 510 2136 516 2137
rect 646 2141 652 2142
rect 646 2137 647 2141
rect 651 2137 652 2141
rect 646 2136 652 2137
rect 774 2141 780 2142
rect 774 2137 775 2141
rect 779 2137 780 2141
rect 774 2136 780 2137
rect 902 2141 908 2142
rect 902 2137 903 2141
rect 907 2137 908 2141
rect 902 2136 908 2137
rect 1022 2141 1028 2142
rect 1022 2137 1023 2141
rect 1027 2137 1028 2141
rect 1022 2136 1028 2137
rect 1150 2141 1156 2142
rect 1150 2137 1151 2141
rect 1155 2137 1156 2141
rect 1150 2136 1156 2137
rect 1278 2141 1284 2142
rect 1278 2137 1279 2141
rect 1283 2137 1284 2141
rect 1278 2136 1284 2137
rect 512 2123 514 2136
rect 648 2123 650 2136
rect 776 2123 778 2136
rect 904 2123 906 2136
rect 1024 2123 1026 2136
rect 1152 2123 1154 2136
rect 1280 2123 1282 2136
rect 1824 2123 1826 2146
rect 1864 2127 1866 2150
rect 2246 2145 2252 2146
rect 2246 2141 2247 2145
rect 2251 2141 2252 2145
rect 2246 2140 2252 2141
rect 2334 2145 2340 2146
rect 2334 2141 2335 2145
rect 2339 2141 2340 2145
rect 2334 2140 2340 2141
rect 2248 2127 2250 2140
rect 2336 2127 2338 2140
rect 1863 2126 1867 2127
rect 479 2122 483 2123
rect 479 2117 483 2118
rect 511 2122 515 2123
rect 511 2117 515 2118
rect 599 2122 603 2123
rect 599 2117 603 2118
rect 647 2122 651 2123
rect 647 2117 651 2118
rect 719 2122 723 2123
rect 719 2117 723 2118
rect 775 2122 779 2123
rect 775 2117 779 2118
rect 831 2122 835 2123
rect 831 2117 835 2118
rect 903 2122 907 2123
rect 903 2117 907 2118
rect 943 2122 947 2123
rect 943 2117 947 2118
rect 1023 2122 1027 2123
rect 1023 2117 1027 2118
rect 1055 2122 1059 2123
rect 1055 2117 1059 2118
rect 1151 2122 1155 2123
rect 1151 2117 1155 2118
rect 1175 2122 1179 2123
rect 1175 2117 1179 2118
rect 1279 2122 1283 2123
rect 1279 2117 1283 2118
rect 1823 2122 1827 2123
rect 1863 2121 1867 2122
rect 2151 2126 2155 2127
rect 2151 2121 2155 2122
rect 2239 2126 2243 2127
rect 2239 2121 2243 2122
rect 2247 2126 2251 2127
rect 2247 2121 2251 2122
rect 2327 2126 2331 2127
rect 2327 2121 2331 2122
rect 2335 2126 2339 2127
rect 2335 2121 2339 2122
rect 1823 2117 1827 2118
rect 480 2112 482 2117
rect 600 2112 602 2117
rect 720 2112 722 2117
rect 832 2112 834 2117
rect 944 2112 946 2117
rect 1056 2112 1058 2117
rect 1176 2112 1178 2117
rect 478 2111 484 2112
rect 478 2107 479 2111
rect 483 2107 484 2111
rect 478 2106 484 2107
rect 598 2111 604 2112
rect 598 2107 599 2111
rect 603 2107 604 2111
rect 598 2106 604 2107
rect 718 2111 724 2112
rect 718 2107 719 2111
rect 723 2107 724 2111
rect 718 2106 724 2107
rect 830 2111 836 2112
rect 830 2107 831 2111
rect 835 2107 836 2111
rect 830 2106 836 2107
rect 942 2111 948 2112
rect 942 2107 943 2111
rect 947 2107 948 2111
rect 942 2106 948 2107
rect 1054 2111 1060 2112
rect 1054 2107 1055 2111
rect 1059 2107 1060 2111
rect 1054 2106 1060 2107
rect 1174 2111 1180 2112
rect 1174 2107 1175 2111
rect 1179 2107 1180 2111
rect 1174 2106 1180 2107
rect 426 2103 432 2104
rect 426 2099 427 2103
rect 431 2099 432 2103
rect 1824 2102 1826 2117
rect 1864 2106 1866 2121
rect 2152 2116 2154 2121
rect 2240 2116 2242 2121
rect 2328 2116 2330 2121
rect 2150 2115 2156 2116
rect 2150 2111 2151 2115
rect 2155 2111 2156 2115
rect 2150 2110 2156 2111
rect 2238 2115 2244 2116
rect 2238 2111 2239 2115
rect 2243 2111 2244 2115
rect 2238 2110 2244 2111
rect 2326 2115 2332 2116
rect 2326 2111 2327 2115
rect 2331 2111 2332 2115
rect 2326 2110 2332 2111
rect 1862 2105 1868 2106
rect 426 2098 432 2099
rect 1822 2101 1828 2102
rect 1822 2097 1823 2101
rect 1827 2097 1828 2101
rect 1862 2101 1863 2105
rect 1867 2101 1868 2105
rect 1862 2100 1868 2101
rect 1822 2096 1828 2097
rect 2306 2091 2312 2092
rect 1862 2088 1868 2089
rect 426 2087 432 2088
rect 426 2083 427 2087
rect 431 2083 432 2087
rect 426 2082 432 2083
rect 546 2087 552 2088
rect 546 2083 547 2087
rect 551 2083 552 2087
rect 546 2082 552 2083
rect 1822 2084 1828 2085
rect 366 2071 372 2072
rect 366 2067 367 2071
rect 371 2067 372 2071
rect 366 2066 372 2067
rect 270 2059 276 2060
rect 270 2055 271 2059
rect 275 2055 276 2059
rect 270 2054 276 2055
rect 368 2043 370 2066
rect 428 2060 430 2082
rect 486 2071 492 2072
rect 486 2067 487 2071
rect 491 2067 492 2071
rect 486 2066 492 2067
rect 426 2059 432 2060
rect 426 2055 427 2059
rect 431 2055 432 2059
rect 426 2054 432 2055
rect 488 2043 490 2066
rect 548 2060 550 2082
rect 1822 2080 1823 2084
rect 1827 2080 1828 2084
rect 1862 2084 1863 2088
rect 1867 2084 1868 2088
rect 2306 2087 2307 2091
rect 2311 2087 2312 2091
rect 2306 2086 2312 2087
rect 1862 2083 1868 2084
rect 1822 2079 1828 2080
rect 606 2071 612 2072
rect 606 2067 607 2071
rect 611 2067 612 2071
rect 606 2066 612 2067
rect 726 2071 732 2072
rect 726 2067 727 2071
rect 731 2067 732 2071
rect 726 2066 732 2067
rect 838 2071 844 2072
rect 838 2067 839 2071
rect 843 2067 844 2071
rect 838 2066 844 2067
rect 950 2071 956 2072
rect 950 2067 951 2071
rect 955 2067 956 2071
rect 950 2066 956 2067
rect 1062 2071 1068 2072
rect 1062 2067 1063 2071
rect 1067 2067 1068 2071
rect 1062 2066 1068 2067
rect 1182 2071 1188 2072
rect 1182 2067 1183 2071
rect 1187 2067 1188 2071
rect 1182 2066 1188 2067
rect 546 2059 552 2060
rect 546 2055 547 2059
rect 551 2055 552 2059
rect 546 2054 552 2055
rect 608 2043 610 2066
rect 634 2059 640 2060
rect 634 2055 635 2059
rect 639 2055 640 2059
rect 634 2054 640 2055
rect 111 2042 115 2043
rect 111 2037 115 2038
rect 143 2042 147 2043
rect 143 2037 147 2038
rect 167 2042 171 2043
rect 167 2037 171 2038
rect 239 2042 243 2043
rect 239 2037 243 2038
rect 311 2042 315 2043
rect 311 2037 315 2038
rect 367 2042 371 2043
rect 367 2037 371 2038
rect 447 2042 451 2043
rect 447 2037 451 2038
rect 487 2042 491 2043
rect 487 2037 491 2038
rect 575 2042 579 2043
rect 575 2037 579 2038
rect 607 2042 611 2043
rect 607 2037 611 2038
rect 112 2013 114 2037
rect 168 2026 170 2037
rect 312 2026 314 2037
rect 386 2035 392 2036
rect 386 2031 387 2035
rect 391 2031 392 2035
rect 386 2030 392 2031
rect 398 2035 404 2036
rect 398 2031 399 2035
rect 403 2031 404 2035
rect 398 2030 404 2031
rect 166 2025 172 2026
rect 166 2021 167 2025
rect 171 2021 172 2025
rect 166 2020 172 2021
rect 310 2025 316 2026
rect 310 2021 311 2025
rect 315 2021 316 2025
rect 310 2020 316 2021
rect 110 2012 116 2013
rect 110 2008 111 2012
rect 115 2008 116 2012
rect 110 2007 116 2008
rect 110 1995 116 1996
rect 110 1991 111 1995
rect 115 1991 116 1995
rect 110 1990 116 1991
rect 112 1975 114 1990
rect 158 1985 164 1986
rect 158 1981 159 1985
rect 163 1981 164 1985
rect 158 1980 164 1981
rect 302 1985 308 1986
rect 302 1981 303 1985
rect 307 1981 308 1985
rect 302 1980 308 1981
rect 160 1975 162 1980
rect 206 1979 212 1980
rect 206 1975 207 1979
rect 211 1975 212 1979
rect 304 1975 306 1980
rect 111 1974 115 1975
rect 111 1969 115 1970
rect 159 1974 163 1975
rect 206 1974 212 1975
rect 295 1974 299 1975
rect 159 1969 163 1970
rect 112 1954 114 1969
rect 160 1964 162 1969
rect 158 1963 164 1964
rect 158 1959 159 1963
rect 163 1959 164 1963
rect 158 1958 164 1959
rect 110 1953 116 1954
rect 110 1949 111 1953
rect 115 1949 116 1953
rect 110 1948 116 1949
rect 110 1936 116 1937
rect 110 1932 111 1936
rect 115 1932 116 1936
rect 110 1931 116 1932
rect 112 1899 114 1931
rect 166 1923 172 1924
rect 166 1919 167 1923
rect 171 1919 172 1923
rect 166 1918 172 1919
rect 168 1899 170 1918
rect 208 1912 210 1974
rect 295 1969 299 1970
rect 303 1974 307 1975
rect 303 1969 307 1970
rect 296 1964 298 1969
rect 294 1963 300 1964
rect 294 1959 295 1963
rect 299 1959 300 1963
rect 294 1958 300 1959
rect 388 1956 390 2030
rect 400 2012 402 2030
rect 448 2026 450 2037
rect 576 2026 578 2037
rect 446 2025 452 2026
rect 446 2021 447 2025
rect 451 2021 452 2025
rect 446 2020 452 2021
rect 574 2025 580 2026
rect 574 2021 575 2025
rect 579 2021 580 2025
rect 574 2020 580 2021
rect 636 2012 638 2054
rect 728 2043 730 2066
rect 758 2059 764 2060
rect 758 2055 759 2059
rect 763 2055 764 2059
rect 758 2054 764 2055
rect 760 2051 762 2054
rect 760 2049 766 2051
rect 695 2042 699 2043
rect 695 2037 699 2038
rect 727 2042 731 2043
rect 727 2037 731 2038
rect 696 2026 698 2037
rect 754 2035 760 2036
rect 726 2031 732 2032
rect 726 2027 727 2031
rect 731 2027 732 2031
rect 754 2031 755 2035
rect 759 2031 760 2035
rect 754 2030 760 2031
rect 726 2026 732 2027
rect 694 2025 700 2026
rect 694 2021 695 2025
rect 699 2021 700 2025
rect 694 2020 700 2021
rect 398 2011 404 2012
rect 398 2007 399 2011
rect 403 2007 404 2011
rect 398 2006 404 2007
rect 634 2011 640 2012
rect 634 2007 635 2011
rect 639 2007 640 2011
rect 634 2006 640 2007
rect 438 1985 444 1986
rect 438 1981 439 1985
rect 443 1981 444 1985
rect 438 1980 444 1981
rect 566 1985 572 1986
rect 566 1981 567 1985
rect 571 1981 572 1985
rect 566 1980 572 1981
rect 686 1985 692 1986
rect 686 1981 687 1985
rect 691 1981 692 1985
rect 686 1980 692 1981
rect 440 1975 442 1980
rect 568 1975 570 1980
rect 688 1975 690 1980
rect 439 1974 443 1975
rect 439 1969 443 1970
rect 567 1974 571 1975
rect 567 1969 571 1970
rect 583 1974 587 1975
rect 583 1969 587 1970
rect 687 1974 691 1975
rect 687 1969 691 1970
rect 719 1974 723 1975
rect 719 1969 723 1970
rect 440 1964 442 1969
rect 584 1964 586 1969
rect 720 1964 722 1969
rect 438 1963 444 1964
rect 438 1959 439 1963
rect 443 1959 444 1963
rect 438 1958 444 1959
rect 582 1963 588 1964
rect 582 1959 583 1963
rect 587 1959 588 1963
rect 582 1958 588 1959
rect 718 1963 724 1964
rect 718 1959 719 1963
rect 723 1959 724 1963
rect 718 1958 724 1959
rect 386 1955 392 1956
rect 386 1951 387 1955
rect 391 1951 392 1955
rect 728 1952 730 2026
rect 756 2012 758 2030
rect 754 2011 760 2012
rect 754 2007 755 2011
rect 759 2007 760 2011
rect 764 2008 766 2049
rect 840 2043 842 2066
rect 952 2043 954 2066
rect 1064 2043 1066 2066
rect 1184 2043 1186 2066
rect 1824 2043 1826 2079
rect 1864 2055 1866 2083
rect 2158 2075 2164 2076
rect 2158 2071 2159 2075
rect 2163 2071 2164 2075
rect 2158 2070 2164 2071
rect 2246 2075 2252 2076
rect 2246 2071 2247 2075
rect 2251 2071 2252 2075
rect 2246 2070 2252 2071
rect 2160 2055 2162 2070
rect 2191 2068 2195 2069
rect 2190 2063 2196 2064
rect 2190 2059 2191 2063
rect 2195 2059 2196 2063
rect 2190 2058 2196 2059
rect 2248 2055 2250 2070
rect 1863 2054 1867 2055
rect 1863 2049 1867 2050
rect 1999 2054 2003 2055
rect 1999 2049 2003 2050
rect 2127 2054 2131 2055
rect 2127 2049 2131 2050
rect 2159 2054 2163 2055
rect 2159 2049 2163 2050
rect 2247 2054 2251 2055
rect 2247 2049 2251 2050
rect 2255 2054 2259 2055
rect 2255 2049 2259 2050
rect 807 2042 811 2043
rect 807 2037 811 2038
rect 839 2042 843 2043
rect 839 2037 843 2038
rect 911 2042 915 2043
rect 911 2037 915 2038
rect 951 2042 955 2043
rect 951 2037 955 2038
rect 1015 2042 1019 2043
rect 1015 2037 1019 2038
rect 1063 2042 1067 2043
rect 1063 2037 1067 2038
rect 1119 2042 1123 2043
rect 1119 2037 1123 2038
rect 1183 2042 1187 2043
rect 1183 2037 1187 2038
rect 1223 2042 1227 2043
rect 1223 2037 1227 2038
rect 1327 2042 1331 2043
rect 1327 2037 1331 2038
rect 1823 2042 1827 2043
rect 1823 2037 1827 2038
rect 808 2026 810 2037
rect 912 2026 914 2037
rect 982 2035 988 2036
rect 982 2031 983 2035
rect 987 2031 988 2035
rect 982 2030 988 2031
rect 806 2025 812 2026
rect 806 2021 807 2025
rect 811 2021 812 2025
rect 806 2020 812 2021
rect 910 2025 916 2026
rect 910 2021 911 2025
rect 915 2021 916 2025
rect 910 2020 916 2021
rect 984 2008 986 2030
rect 1016 2026 1018 2037
rect 1082 2035 1088 2036
rect 1082 2031 1083 2035
rect 1087 2031 1088 2035
rect 1082 2030 1088 2031
rect 1014 2025 1020 2026
rect 1014 2021 1015 2025
rect 1019 2021 1020 2025
rect 1014 2020 1020 2021
rect 1084 2008 1086 2030
rect 1120 2026 1122 2037
rect 1190 2035 1196 2036
rect 1190 2031 1191 2035
rect 1195 2031 1196 2035
rect 1190 2030 1196 2031
rect 1118 2025 1124 2026
rect 1118 2021 1119 2025
rect 1123 2021 1124 2025
rect 1118 2020 1124 2021
rect 1192 2008 1194 2030
rect 1224 2026 1226 2037
rect 1310 2035 1316 2036
rect 1310 2031 1311 2035
rect 1315 2031 1316 2035
rect 1310 2030 1316 2031
rect 1222 2025 1228 2026
rect 1222 2021 1223 2025
rect 1227 2021 1228 2025
rect 1222 2020 1228 2021
rect 754 2006 760 2007
rect 762 2007 768 2008
rect 762 2003 763 2007
rect 767 2003 768 2007
rect 762 2002 768 2003
rect 982 2007 988 2008
rect 982 2003 983 2007
rect 987 2003 988 2007
rect 982 2002 988 2003
rect 1082 2007 1088 2008
rect 1082 2003 1083 2007
rect 1087 2003 1088 2007
rect 1082 2002 1088 2003
rect 1190 2007 1196 2008
rect 1190 2003 1191 2007
rect 1195 2003 1196 2007
rect 1190 2002 1196 2003
rect 1014 1995 1020 1996
rect 1014 1991 1015 1995
rect 1019 1991 1020 1995
rect 1014 1990 1020 1991
rect 798 1985 804 1986
rect 798 1981 799 1985
rect 803 1981 804 1985
rect 798 1980 804 1981
rect 902 1985 908 1986
rect 902 1981 903 1985
rect 907 1981 908 1985
rect 902 1980 908 1981
rect 1006 1985 1012 1986
rect 1006 1981 1007 1985
rect 1011 1981 1012 1985
rect 1006 1980 1012 1981
rect 800 1975 802 1980
rect 904 1975 906 1980
rect 1008 1975 1010 1980
rect 799 1974 803 1975
rect 799 1969 803 1970
rect 855 1974 859 1975
rect 855 1969 859 1970
rect 903 1974 907 1975
rect 903 1969 907 1970
rect 991 1974 995 1975
rect 991 1969 995 1970
rect 1007 1974 1011 1975
rect 1007 1969 1011 1970
rect 856 1964 858 1969
rect 992 1964 994 1969
rect 854 1963 860 1964
rect 854 1959 855 1963
rect 859 1959 860 1963
rect 854 1958 860 1959
rect 990 1963 996 1964
rect 990 1959 991 1963
rect 995 1959 996 1963
rect 990 1958 996 1959
rect 386 1950 392 1951
rect 726 1951 732 1952
rect 726 1947 727 1951
rect 731 1947 732 1951
rect 726 1946 732 1947
rect 506 1939 512 1940
rect 506 1935 507 1939
rect 511 1935 512 1939
rect 506 1934 512 1935
rect 786 1939 792 1940
rect 786 1935 787 1939
rect 791 1935 792 1939
rect 786 1934 792 1935
rect 922 1939 928 1940
rect 922 1935 923 1939
rect 927 1935 928 1939
rect 922 1934 928 1935
rect 302 1923 308 1924
rect 302 1919 303 1923
rect 307 1919 308 1923
rect 302 1918 308 1919
rect 446 1923 452 1924
rect 446 1919 447 1923
rect 451 1919 452 1923
rect 446 1918 452 1919
rect 206 1911 212 1912
rect 206 1907 207 1911
rect 211 1907 212 1911
rect 206 1906 212 1907
rect 304 1899 306 1918
rect 448 1899 450 1918
rect 508 1912 510 1934
rect 590 1923 596 1924
rect 590 1919 591 1923
rect 595 1919 596 1923
rect 590 1918 596 1919
rect 726 1923 732 1924
rect 726 1919 727 1923
rect 731 1919 732 1923
rect 788 1920 790 1934
rect 862 1923 868 1924
rect 726 1918 732 1919
rect 786 1919 792 1920
rect 506 1911 512 1912
rect 506 1907 507 1911
rect 511 1907 512 1911
rect 506 1906 512 1907
rect 592 1899 594 1918
rect 728 1899 730 1918
rect 786 1915 787 1919
rect 791 1915 792 1919
rect 862 1919 863 1923
rect 867 1919 868 1923
rect 862 1918 868 1919
rect 786 1914 792 1915
rect 778 1911 784 1912
rect 778 1907 779 1911
rect 783 1907 784 1911
rect 778 1906 784 1907
rect 111 1898 115 1899
rect 111 1893 115 1894
rect 167 1898 171 1899
rect 167 1893 171 1894
rect 223 1898 227 1899
rect 223 1893 227 1894
rect 303 1898 307 1899
rect 303 1893 307 1894
rect 447 1898 451 1899
rect 447 1893 451 1894
rect 479 1898 483 1899
rect 479 1893 483 1894
rect 591 1898 595 1899
rect 591 1893 595 1894
rect 719 1898 723 1899
rect 719 1893 723 1894
rect 727 1898 731 1899
rect 727 1893 731 1894
rect 112 1869 114 1893
rect 224 1882 226 1893
rect 480 1882 482 1893
rect 720 1882 722 1893
rect 750 1891 756 1892
rect 750 1887 751 1891
rect 755 1887 756 1891
rect 750 1886 756 1887
rect 222 1881 228 1882
rect 222 1877 223 1881
rect 227 1877 228 1881
rect 222 1876 228 1877
rect 478 1881 484 1882
rect 478 1877 479 1881
rect 483 1877 484 1881
rect 478 1876 484 1877
rect 718 1881 724 1882
rect 718 1877 719 1881
rect 723 1877 724 1881
rect 718 1876 724 1877
rect 110 1868 116 1869
rect 110 1864 111 1868
rect 115 1864 116 1868
rect 110 1863 116 1864
rect 110 1851 116 1852
rect 110 1847 111 1851
rect 115 1847 116 1851
rect 110 1846 116 1847
rect 112 1831 114 1846
rect 214 1841 220 1842
rect 214 1837 215 1841
rect 219 1837 220 1841
rect 214 1836 220 1837
rect 470 1841 476 1842
rect 470 1837 471 1841
rect 475 1837 476 1841
rect 470 1836 476 1837
rect 710 1841 716 1842
rect 710 1837 711 1841
rect 715 1837 716 1841
rect 710 1836 716 1837
rect 216 1831 218 1836
rect 282 1835 288 1836
rect 282 1831 283 1835
rect 287 1831 288 1835
rect 472 1831 474 1836
rect 712 1831 714 1836
rect 111 1830 115 1831
rect 111 1825 115 1826
rect 215 1830 219 1831
rect 215 1825 219 1826
rect 247 1830 251 1831
rect 282 1830 288 1831
rect 415 1830 419 1831
rect 247 1825 251 1826
rect 112 1810 114 1825
rect 248 1820 250 1825
rect 246 1819 252 1820
rect 246 1815 247 1819
rect 251 1815 252 1819
rect 246 1814 252 1815
rect 110 1809 116 1810
rect 110 1805 111 1809
rect 115 1805 116 1809
rect 110 1804 116 1805
rect 110 1792 116 1793
rect 110 1788 111 1792
rect 115 1788 116 1792
rect 110 1787 116 1788
rect 112 1759 114 1787
rect 254 1779 260 1780
rect 254 1775 255 1779
rect 259 1775 260 1779
rect 254 1774 260 1775
rect 256 1759 258 1774
rect 284 1768 286 1830
rect 415 1825 419 1826
rect 471 1830 475 1831
rect 471 1825 475 1826
rect 591 1830 595 1831
rect 591 1825 595 1826
rect 711 1830 715 1831
rect 711 1825 715 1826
rect 416 1820 418 1825
rect 592 1820 594 1825
rect 414 1819 420 1820
rect 414 1815 415 1819
rect 419 1815 420 1819
rect 414 1814 420 1815
rect 590 1819 596 1820
rect 590 1815 591 1819
rect 595 1815 596 1819
rect 590 1814 596 1815
rect 752 1812 754 1886
rect 780 1868 782 1906
rect 864 1899 866 1918
rect 924 1912 926 1934
rect 998 1923 1004 1924
rect 998 1919 999 1923
rect 1003 1919 1004 1923
rect 998 1918 1004 1919
rect 922 1911 928 1912
rect 922 1907 923 1911
rect 927 1907 928 1911
rect 922 1906 928 1907
rect 1000 1899 1002 1918
rect 1016 1912 1018 1990
rect 1110 1985 1116 1986
rect 1110 1981 1111 1985
rect 1115 1981 1116 1985
rect 1110 1980 1116 1981
rect 1214 1985 1220 1986
rect 1214 1981 1215 1985
rect 1219 1981 1220 1985
rect 1214 1980 1220 1981
rect 1112 1975 1114 1980
rect 1216 1975 1218 1980
rect 1111 1974 1115 1975
rect 1111 1969 1115 1970
rect 1119 1974 1123 1975
rect 1119 1969 1123 1970
rect 1215 1974 1219 1975
rect 1215 1969 1219 1970
rect 1239 1974 1243 1975
rect 1239 1969 1243 1970
rect 1120 1964 1122 1969
rect 1240 1964 1242 1969
rect 1118 1963 1124 1964
rect 1118 1959 1119 1963
rect 1123 1959 1124 1963
rect 1118 1958 1124 1959
rect 1238 1963 1244 1964
rect 1238 1959 1239 1963
rect 1243 1959 1244 1963
rect 1238 1958 1244 1959
rect 1312 1956 1314 2030
rect 1328 2026 1330 2037
rect 1326 2025 1332 2026
rect 1326 2021 1327 2025
rect 1331 2021 1332 2025
rect 1326 2020 1332 2021
rect 1824 2013 1826 2037
rect 1864 2025 1866 2049
rect 2000 2038 2002 2049
rect 2070 2047 2076 2048
rect 2070 2043 2071 2047
rect 2075 2043 2076 2047
rect 2070 2042 2076 2043
rect 1998 2037 2004 2038
rect 1998 2033 1999 2037
rect 2003 2033 2004 2037
rect 1998 2032 2004 2033
rect 1862 2024 1868 2025
rect 1862 2020 1863 2024
rect 1867 2020 1868 2024
rect 2072 2021 2074 2042
rect 2128 2038 2130 2049
rect 2256 2038 2258 2049
rect 2308 2048 2310 2086
rect 2334 2075 2340 2076
rect 2334 2071 2335 2075
rect 2339 2071 2340 2075
rect 2334 2070 2340 2071
rect 2336 2055 2338 2070
rect 2344 2064 2346 2150
rect 2430 2145 2436 2146
rect 2430 2141 2431 2145
rect 2435 2141 2436 2145
rect 2430 2140 2436 2141
rect 2542 2145 2548 2146
rect 2542 2141 2543 2145
rect 2547 2141 2548 2145
rect 2542 2140 2548 2141
rect 2686 2145 2692 2146
rect 2686 2141 2687 2145
rect 2691 2141 2692 2145
rect 2686 2140 2692 2141
rect 2862 2145 2868 2146
rect 2862 2141 2863 2145
rect 2867 2141 2868 2145
rect 2862 2140 2868 2141
rect 3062 2145 3068 2146
rect 3062 2141 3063 2145
rect 3067 2141 3068 2145
rect 3062 2140 3068 2141
rect 2432 2127 2434 2140
rect 2544 2127 2546 2140
rect 2688 2127 2690 2140
rect 2864 2127 2866 2140
rect 3064 2127 3066 2140
rect 2415 2126 2419 2127
rect 2415 2121 2419 2122
rect 2431 2126 2435 2127
rect 2431 2121 2435 2122
rect 2503 2126 2507 2127
rect 2503 2121 2507 2122
rect 2543 2126 2547 2127
rect 2543 2121 2547 2122
rect 2615 2126 2619 2127
rect 2615 2121 2619 2122
rect 2687 2126 2691 2127
rect 2687 2121 2691 2122
rect 2751 2126 2755 2127
rect 2751 2121 2755 2122
rect 2863 2126 2867 2127
rect 2863 2121 2867 2122
rect 2919 2126 2923 2127
rect 2919 2121 2923 2122
rect 3063 2126 3067 2127
rect 3063 2121 3067 2122
rect 3103 2126 3107 2127
rect 3103 2121 3107 2122
rect 2416 2116 2418 2121
rect 2504 2116 2506 2121
rect 2616 2116 2618 2121
rect 2752 2116 2754 2121
rect 2920 2116 2922 2121
rect 3104 2116 3106 2121
rect 2414 2115 2420 2116
rect 2414 2111 2415 2115
rect 2419 2111 2420 2115
rect 2414 2110 2420 2111
rect 2502 2115 2508 2116
rect 2502 2111 2503 2115
rect 2507 2111 2508 2115
rect 2502 2110 2508 2111
rect 2614 2115 2620 2116
rect 2614 2111 2615 2115
rect 2619 2111 2620 2115
rect 2614 2110 2620 2111
rect 2750 2115 2756 2116
rect 2750 2111 2751 2115
rect 2755 2111 2756 2115
rect 2750 2110 2756 2111
rect 2918 2115 2924 2116
rect 2918 2111 2919 2115
rect 2923 2111 2924 2115
rect 2918 2110 2924 2111
rect 3102 2115 3108 2116
rect 3102 2111 3103 2115
rect 3107 2111 3108 2115
rect 3102 2110 3108 2111
rect 3200 2109 3202 2150
rect 3278 2145 3284 2146
rect 3278 2141 3279 2145
rect 3283 2141 3284 2145
rect 3278 2140 3284 2141
rect 3280 2127 3282 2140
rect 3279 2126 3283 2127
rect 3279 2121 3283 2122
rect 3303 2126 3307 2127
rect 3303 2121 3307 2122
rect 3304 2116 3306 2121
rect 3302 2115 3308 2116
rect 3302 2111 3303 2115
rect 3307 2111 3308 2115
rect 3302 2110 3308 2111
rect 2663 2108 2667 2109
rect 2482 2107 2488 2108
rect 2482 2103 2483 2107
rect 2487 2103 2488 2107
rect 2663 2103 2667 2104
rect 3199 2108 3203 2109
rect 3199 2103 3203 2104
rect 2482 2102 2488 2103
rect 2422 2075 2428 2076
rect 2422 2071 2423 2075
rect 2427 2071 2428 2075
rect 2422 2070 2428 2071
rect 2342 2063 2348 2064
rect 2342 2059 2343 2063
rect 2347 2059 2348 2063
rect 2342 2058 2348 2059
rect 2424 2055 2426 2070
rect 2484 2069 2486 2102
rect 2510 2075 2516 2076
rect 2510 2071 2511 2075
rect 2515 2071 2516 2075
rect 2510 2070 2516 2071
rect 2622 2075 2628 2076
rect 2622 2071 2623 2075
rect 2627 2071 2628 2075
rect 2622 2070 2628 2071
rect 2483 2068 2487 2069
rect 2483 2063 2487 2064
rect 2512 2055 2514 2070
rect 2624 2055 2626 2070
rect 2664 2064 2666 2103
rect 3094 2091 3100 2092
rect 3094 2087 3095 2091
rect 3099 2087 3100 2091
rect 3094 2086 3100 2087
rect 2758 2075 2764 2076
rect 2758 2071 2759 2075
rect 2763 2071 2764 2075
rect 2758 2070 2764 2071
rect 2926 2075 2932 2076
rect 2926 2071 2927 2075
rect 2931 2071 2932 2075
rect 2926 2070 2932 2071
rect 2662 2063 2668 2064
rect 2662 2059 2663 2063
rect 2667 2059 2668 2063
rect 2662 2058 2668 2059
rect 2760 2055 2762 2070
rect 2928 2055 2930 2070
rect 3096 2064 3098 2086
rect 3110 2075 3116 2076
rect 3110 2071 3111 2075
rect 3115 2071 3116 2075
rect 3110 2070 3116 2071
rect 3310 2075 3316 2076
rect 3310 2071 3311 2075
rect 3315 2071 3316 2075
rect 3310 2070 3316 2071
rect 3094 2063 3100 2064
rect 3094 2059 3095 2063
rect 3099 2059 3100 2063
rect 3094 2058 3100 2059
rect 3112 2055 3114 2070
rect 3312 2055 3314 2070
rect 2335 2054 2339 2055
rect 2335 2049 2339 2050
rect 2399 2054 2403 2055
rect 2399 2049 2403 2050
rect 2423 2054 2427 2055
rect 2423 2049 2427 2050
rect 2511 2054 2515 2055
rect 2511 2049 2515 2050
rect 2551 2054 2555 2055
rect 2551 2049 2555 2050
rect 2623 2054 2627 2055
rect 2623 2049 2627 2050
rect 2711 2054 2715 2055
rect 2711 2049 2715 2050
rect 2759 2054 2763 2055
rect 2759 2049 2763 2050
rect 2879 2054 2883 2055
rect 2879 2049 2883 2050
rect 2927 2054 2931 2055
rect 2927 2049 2931 2050
rect 3063 2054 3067 2055
rect 3063 2049 3067 2050
rect 3111 2054 3115 2055
rect 3111 2049 3115 2050
rect 3247 2054 3251 2055
rect 3247 2049 3251 2050
rect 3311 2054 3315 2055
rect 3311 2049 3315 2050
rect 2306 2047 2312 2048
rect 2306 2043 2307 2047
rect 2311 2043 2312 2047
rect 2306 2042 2312 2043
rect 2366 2047 2372 2048
rect 2366 2043 2367 2047
rect 2371 2043 2372 2047
rect 2366 2042 2372 2043
rect 2126 2037 2132 2038
rect 2126 2033 2127 2037
rect 2131 2033 2132 2037
rect 2126 2032 2132 2033
rect 2254 2037 2260 2038
rect 2254 2033 2255 2037
rect 2259 2033 2260 2037
rect 2254 2032 2260 2033
rect 2368 2024 2370 2042
rect 2400 2038 2402 2049
rect 2552 2038 2554 2049
rect 2712 2038 2714 2049
rect 2830 2047 2836 2048
rect 2830 2043 2831 2047
rect 2835 2043 2836 2047
rect 2830 2042 2836 2043
rect 2398 2037 2404 2038
rect 2398 2033 2399 2037
rect 2403 2033 2404 2037
rect 2398 2032 2404 2033
rect 2550 2037 2556 2038
rect 2550 2033 2551 2037
rect 2555 2033 2556 2037
rect 2550 2032 2556 2033
rect 2710 2037 2716 2038
rect 2710 2033 2711 2037
rect 2715 2033 2716 2037
rect 2710 2032 2716 2033
rect 2832 2024 2834 2042
rect 2880 2038 2882 2049
rect 2990 2047 2996 2048
rect 2990 2043 2991 2047
rect 2995 2043 2996 2047
rect 2990 2042 2996 2043
rect 2878 2037 2884 2038
rect 2878 2033 2879 2037
rect 2883 2033 2884 2037
rect 2878 2032 2884 2033
rect 2992 2024 2994 2042
rect 3064 2038 3066 2049
rect 3174 2047 3180 2048
rect 3174 2043 3175 2047
rect 3179 2043 3180 2047
rect 3174 2042 3180 2043
rect 3062 2037 3068 2038
rect 3062 2033 3063 2037
rect 3067 2033 3068 2037
rect 3062 2032 3068 2033
rect 3176 2024 3178 2042
rect 3248 2038 3250 2049
rect 3246 2037 3252 2038
rect 3246 2033 3247 2037
rect 3251 2033 3252 2037
rect 3246 2032 3252 2033
rect 2366 2023 2372 2024
rect 1862 2019 1868 2020
rect 2071 2020 2075 2021
rect 2366 2019 2367 2023
rect 2371 2019 2372 2023
rect 2830 2023 2836 2024
rect 2479 2020 2483 2021
rect 2366 2018 2372 2019
rect 2071 2015 2075 2016
rect 2478 2015 2479 2020
rect 2483 2015 2484 2020
rect 2830 2019 2831 2023
rect 2835 2019 2836 2023
rect 2830 2018 2836 2019
rect 2990 2023 2996 2024
rect 2990 2019 2991 2023
rect 2995 2019 2996 2023
rect 2990 2018 2996 2019
rect 3174 2023 3180 2024
rect 3174 2019 3175 2023
rect 3179 2019 3180 2023
rect 3344 2020 3346 2202
rect 3487 2197 3491 2198
rect 3488 2186 3490 2197
rect 3548 2196 3550 2230
rect 3574 2228 3575 2232
rect 3579 2228 3580 2232
rect 3574 2227 3580 2228
rect 3576 2203 3578 2227
rect 3575 2202 3579 2203
rect 3575 2197 3579 2198
rect 3546 2195 3552 2196
rect 3546 2191 3547 2195
rect 3551 2191 3552 2195
rect 3546 2190 3552 2191
rect 3486 2185 3492 2186
rect 3486 2181 3487 2185
rect 3491 2181 3492 2185
rect 3486 2180 3492 2181
rect 3576 2173 3578 2197
rect 3574 2172 3580 2173
rect 3574 2168 3575 2172
rect 3579 2168 3580 2172
rect 3574 2167 3580 2168
rect 3574 2155 3580 2156
rect 3574 2151 3575 2155
rect 3579 2151 3580 2155
rect 3574 2150 3580 2151
rect 3478 2145 3484 2146
rect 3478 2141 3479 2145
rect 3483 2141 3484 2145
rect 3478 2140 3484 2141
rect 3480 2127 3482 2140
rect 3518 2139 3524 2140
rect 3518 2135 3519 2139
rect 3523 2135 3524 2139
rect 3518 2134 3524 2135
rect 3479 2126 3483 2127
rect 3479 2121 3483 2122
rect 3480 2116 3482 2121
rect 3478 2115 3484 2116
rect 3478 2111 3479 2115
rect 3483 2111 3484 2115
rect 3478 2110 3484 2111
rect 3486 2075 3492 2076
rect 3486 2071 3487 2075
rect 3491 2071 3492 2075
rect 3486 2070 3492 2071
rect 3488 2055 3490 2070
rect 3520 2064 3522 2134
rect 3576 2127 3578 2150
rect 3575 2126 3579 2127
rect 3575 2121 3579 2122
rect 3576 2106 3578 2121
rect 3574 2105 3580 2106
rect 3574 2101 3575 2105
rect 3579 2101 3580 2105
rect 3574 2100 3580 2101
rect 3554 2091 3560 2092
rect 3554 2087 3555 2091
rect 3559 2087 3560 2091
rect 3554 2086 3560 2087
rect 3574 2088 3580 2089
rect 3518 2063 3524 2064
rect 3518 2059 3519 2063
rect 3523 2059 3524 2063
rect 3518 2058 3524 2059
rect 3439 2054 3443 2055
rect 3439 2049 3443 2050
rect 3487 2054 3491 2055
rect 3487 2049 3491 2050
rect 3418 2047 3424 2048
rect 3418 2043 3419 2047
rect 3423 2043 3424 2047
rect 3418 2042 3424 2043
rect 3174 2018 3180 2019
rect 3342 2019 3348 2020
rect 2478 2014 2484 2015
rect 3342 2015 3343 2019
rect 3347 2015 3348 2019
rect 3342 2014 3348 2015
rect 1822 2012 1828 2013
rect 1822 2008 1823 2012
rect 1827 2008 1828 2012
rect 1822 2007 1828 2008
rect 1862 2007 1868 2008
rect 1862 2003 1863 2007
rect 1867 2003 1868 2007
rect 1862 2002 1868 2003
rect 2194 2007 2200 2008
rect 2194 2003 2195 2007
rect 2199 2003 2200 2007
rect 2194 2002 2200 2003
rect 3150 2007 3156 2008
rect 3150 2003 3151 2007
rect 3155 2003 3156 2007
rect 3150 2002 3156 2003
rect 1822 1995 1828 1996
rect 1822 1991 1823 1995
rect 1827 1991 1828 1995
rect 1822 1990 1828 1991
rect 1318 1985 1324 1986
rect 1318 1981 1319 1985
rect 1323 1981 1324 1985
rect 1318 1980 1324 1981
rect 1320 1975 1322 1980
rect 1824 1975 1826 1990
rect 1864 1979 1866 2002
rect 1990 1997 1996 1998
rect 1990 1993 1991 1997
rect 1995 1993 1996 1997
rect 1990 1992 1996 1993
rect 2118 1997 2124 1998
rect 2118 1993 2119 1997
rect 2123 1993 2124 1997
rect 2118 1992 2124 1993
rect 1992 1979 1994 1992
rect 2120 1979 2122 1992
rect 1863 1978 1867 1979
rect 1319 1974 1323 1975
rect 1319 1969 1323 1970
rect 1359 1974 1363 1975
rect 1359 1969 1363 1970
rect 1479 1974 1483 1975
rect 1479 1969 1483 1970
rect 1599 1974 1603 1975
rect 1599 1969 1603 1970
rect 1823 1974 1827 1975
rect 1863 1973 1867 1974
rect 1903 1978 1907 1979
rect 1903 1973 1907 1974
rect 1991 1978 1995 1979
rect 1991 1973 1995 1974
rect 2119 1978 2123 1979
rect 2119 1973 2123 1974
rect 2159 1978 2163 1979
rect 2159 1973 2163 1974
rect 1823 1969 1827 1970
rect 1360 1964 1362 1969
rect 1480 1964 1482 1969
rect 1600 1964 1602 1969
rect 1358 1963 1364 1964
rect 1358 1959 1359 1963
rect 1363 1959 1364 1963
rect 1358 1958 1364 1959
rect 1478 1963 1484 1964
rect 1478 1959 1479 1963
rect 1483 1959 1484 1963
rect 1478 1958 1484 1959
rect 1598 1963 1604 1964
rect 1598 1959 1599 1963
rect 1603 1959 1604 1963
rect 1598 1958 1604 1959
rect 1310 1955 1316 1956
rect 1310 1951 1311 1955
rect 1315 1951 1316 1955
rect 1824 1954 1826 1969
rect 1864 1958 1866 1973
rect 1904 1968 1906 1973
rect 2160 1968 2162 1973
rect 1902 1967 1908 1968
rect 1902 1963 1903 1967
rect 1907 1963 1908 1967
rect 1902 1962 1908 1963
rect 2158 1967 2164 1968
rect 2158 1963 2159 1967
rect 2163 1963 2164 1967
rect 2158 1962 2164 1963
rect 1862 1957 1868 1958
rect 1310 1950 1316 1951
rect 1822 1953 1828 1954
rect 1822 1949 1823 1953
rect 1827 1949 1828 1953
rect 1862 1953 1863 1957
rect 1867 1953 1868 1957
rect 1862 1952 1868 1953
rect 1822 1948 1828 1949
rect 2010 1943 2016 1944
rect 1862 1940 1868 1941
rect 1306 1939 1312 1940
rect 1306 1935 1307 1939
rect 1311 1935 1312 1939
rect 1306 1934 1312 1935
rect 1426 1939 1432 1940
rect 1426 1935 1427 1939
rect 1431 1935 1432 1939
rect 1426 1934 1432 1935
rect 1546 1939 1552 1940
rect 1546 1935 1547 1939
rect 1551 1935 1552 1939
rect 1546 1934 1552 1935
rect 1822 1936 1828 1937
rect 1126 1923 1132 1924
rect 1126 1919 1127 1923
rect 1131 1919 1132 1923
rect 1126 1918 1132 1919
rect 1246 1923 1252 1924
rect 1246 1919 1247 1923
rect 1251 1919 1252 1923
rect 1246 1918 1252 1919
rect 1014 1911 1020 1912
rect 1014 1907 1015 1911
rect 1019 1907 1020 1911
rect 1014 1906 1020 1907
rect 1128 1899 1130 1918
rect 1248 1899 1250 1918
rect 1308 1904 1310 1934
rect 1366 1923 1372 1924
rect 1366 1919 1367 1923
rect 1371 1919 1372 1923
rect 1366 1918 1372 1919
rect 1306 1903 1312 1904
rect 1306 1899 1307 1903
rect 1311 1899 1312 1903
rect 1368 1899 1370 1918
rect 1428 1912 1430 1934
rect 1486 1923 1492 1924
rect 1486 1919 1487 1923
rect 1491 1919 1492 1923
rect 1486 1918 1492 1919
rect 1426 1911 1432 1912
rect 1426 1907 1427 1911
rect 1431 1907 1432 1911
rect 1426 1906 1432 1907
rect 1488 1899 1490 1918
rect 1548 1912 1550 1934
rect 1822 1932 1823 1936
rect 1827 1932 1828 1936
rect 1862 1936 1863 1940
rect 1867 1936 1868 1940
rect 2010 1939 2011 1943
rect 2015 1939 2016 1943
rect 2010 1938 2016 1939
rect 1862 1935 1868 1936
rect 1822 1931 1828 1932
rect 1606 1923 1612 1924
rect 1606 1919 1607 1923
rect 1611 1919 1612 1923
rect 1606 1918 1612 1919
rect 1546 1911 1552 1912
rect 1546 1907 1547 1911
rect 1551 1907 1552 1911
rect 1546 1906 1552 1907
rect 1608 1899 1610 1918
rect 1666 1911 1672 1912
rect 1666 1907 1667 1911
rect 1671 1907 1672 1911
rect 1666 1906 1672 1907
rect 863 1898 867 1899
rect 863 1893 867 1894
rect 935 1898 939 1899
rect 935 1893 939 1894
rect 999 1898 1003 1899
rect 999 1893 1003 1894
rect 1127 1898 1131 1899
rect 1127 1893 1131 1894
rect 1247 1898 1251 1899
rect 1247 1893 1251 1894
rect 1295 1898 1299 1899
rect 1306 1898 1312 1899
rect 1367 1898 1371 1899
rect 1295 1893 1299 1894
rect 1367 1893 1371 1894
rect 1455 1898 1459 1899
rect 1455 1893 1459 1894
rect 1487 1898 1491 1899
rect 1487 1893 1491 1894
rect 1607 1898 1611 1899
rect 1607 1893 1611 1894
rect 936 1882 938 1893
rect 1030 1891 1036 1892
rect 1030 1887 1031 1891
rect 1035 1887 1036 1891
rect 1030 1886 1036 1887
rect 934 1881 940 1882
rect 934 1877 935 1881
rect 939 1877 940 1881
rect 934 1876 940 1877
rect 778 1867 784 1868
rect 778 1863 779 1867
rect 783 1863 784 1867
rect 778 1862 784 1863
rect 926 1841 932 1842
rect 926 1837 927 1841
rect 931 1837 932 1841
rect 926 1836 932 1837
rect 928 1831 930 1836
rect 759 1830 763 1831
rect 759 1825 763 1826
rect 927 1830 931 1831
rect 927 1825 931 1826
rect 760 1820 762 1825
rect 928 1820 930 1825
rect 758 1819 764 1820
rect 758 1815 759 1819
rect 763 1815 764 1819
rect 758 1814 764 1815
rect 926 1819 932 1820
rect 926 1815 927 1819
rect 931 1815 932 1819
rect 926 1814 932 1815
rect 1032 1812 1034 1886
rect 1128 1882 1130 1893
rect 1296 1882 1298 1893
rect 1456 1882 1458 1893
rect 1608 1882 1610 1893
rect 1126 1881 1132 1882
rect 1126 1877 1127 1881
rect 1131 1877 1132 1881
rect 1126 1876 1132 1877
rect 1294 1881 1300 1882
rect 1294 1877 1295 1881
rect 1299 1877 1300 1881
rect 1294 1876 1300 1877
rect 1454 1881 1460 1882
rect 1454 1877 1455 1881
rect 1459 1877 1460 1881
rect 1454 1876 1460 1877
rect 1606 1881 1612 1882
rect 1606 1877 1607 1881
rect 1611 1877 1612 1881
rect 1606 1876 1612 1877
rect 1668 1868 1670 1906
rect 1824 1899 1826 1931
rect 1864 1911 1866 1935
rect 1910 1927 1916 1928
rect 1910 1923 1911 1927
rect 1915 1923 1916 1927
rect 1910 1922 1916 1923
rect 1912 1911 1914 1922
rect 1942 1915 1948 1916
rect 1942 1911 1943 1915
rect 1947 1911 1948 1915
rect 1863 1910 1867 1911
rect 1863 1905 1867 1906
rect 1895 1910 1899 1911
rect 1895 1905 1899 1906
rect 1911 1910 1915 1911
rect 1942 1910 1948 1911
rect 1983 1910 1987 1911
rect 1911 1905 1915 1906
rect 1735 1898 1739 1899
rect 1735 1893 1739 1894
rect 1823 1898 1827 1899
rect 1823 1893 1827 1894
rect 1736 1882 1738 1893
rect 1734 1881 1740 1882
rect 1734 1877 1735 1881
rect 1739 1877 1740 1881
rect 1734 1876 1740 1877
rect 1824 1869 1826 1893
rect 1864 1881 1866 1905
rect 1896 1894 1898 1905
rect 1894 1893 1900 1894
rect 1894 1889 1895 1893
rect 1899 1889 1900 1893
rect 1894 1888 1900 1889
rect 1944 1885 1946 1910
rect 1983 1905 1987 1906
rect 1984 1894 1986 1905
rect 2012 1904 2014 1938
rect 2166 1927 2172 1928
rect 2166 1923 2167 1927
rect 2171 1923 2172 1927
rect 2166 1922 2172 1923
rect 2168 1911 2170 1922
rect 2196 1916 2198 2002
rect 2246 1997 2252 1998
rect 2246 1993 2247 1997
rect 2251 1993 2252 1997
rect 2246 1992 2252 1993
rect 2390 1997 2396 1998
rect 2390 1993 2391 1997
rect 2395 1993 2396 1997
rect 2390 1992 2396 1993
rect 2542 1997 2548 1998
rect 2542 1993 2543 1997
rect 2547 1993 2548 1997
rect 2542 1992 2548 1993
rect 2702 1997 2708 1998
rect 2702 1993 2703 1997
rect 2707 1993 2708 1997
rect 2702 1992 2708 1993
rect 2870 1997 2876 1998
rect 2870 1993 2871 1997
rect 2875 1993 2876 1997
rect 2870 1992 2876 1993
rect 3054 1997 3060 1998
rect 3054 1993 3055 1997
rect 3059 1993 3060 1997
rect 3054 1992 3060 1993
rect 2248 1979 2250 1992
rect 2392 1979 2394 1992
rect 2544 1979 2546 1992
rect 2704 1979 2706 1992
rect 2872 1979 2874 1992
rect 3056 1979 3058 1992
rect 2247 1978 2251 1979
rect 2247 1973 2251 1974
rect 2391 1978 2395 1979
rect 2391 1973 2395 1974
rect 2399 1978 2403 1979
rect 2399 1973 2403 1974
rect 2543 1978 2547 1979
rect 2543 1973 2547 1974
rect 2615 1978 2619 1979
rect 2615 1973 2619 1974
rect 2703 1978 2707 1979
rect 2703 1973 2707 1974
rect 2815 1978 2819 1979
rect 2815 1973 2819 1974
rect 2871 1978 2875 1979
rect 2871 1973 2875 1974
rect 2999 1978 3003 1979
rect 2999 1973 3003 1974
rect 3055 1978 3059 1979
rect 3055 1973 3059 1974
rect 2400 1968 2402 1973
rect 2616 1968 2618 1973
rect 2816 1968 2818 1973
rect 3000 1968 3002 1973
rect 2398 1967 2404 1968
rect 2398 1963 2399 1967
rect 2403 1963 2404 1967
rect 2398 1962 2404 1963
rect 2614 1967 2620 1968
rect 2614 1963 2615 1967
rect 2619 1963 2620 1967
rect 2614 1962 2620 1963
rect 2814 1967 2820 1968
rect 2814 1963 2815 1967
rect 2819 1963 2820 1967
rect 2814 1962 2820 1963
rect 2998 1967 3004 1968
rect 2998 1963 2999 1967
rect 3003 1963 3004 1967
rect 2998 1962 3004 1963
rect 3152 1941 3154 2002
rect 3238 1997 3244 1998
rect 3238 1993 3239 1997
rect 3243 1993 3244 1997
rect 3238 1992 3244 1993
rect 3240 1979 3242 1992
rect 3167 1978 3171 1979
rect 3167 1973 3171 1974
rect 3239 1978 3243 1979
rect 3239 1973 3243 1974
rect 3335 1978 3339 1979
rect 3335 1973 3339 1974
rect 3168 1968 3170 1973
rect 3336 1968 3338 1973
rect 3166 1967 3172 1968
rect 3166 1963 3167 1967
rect 3171 1963 3172 1967
rect 3166 1962 3172 1963
rect 3334 1967 3340 1968
rect 3334 1963 3335 1967
rect 3339 1963 3340 1967
rect 3334 1962 3340 1963
rect 3258 1959 3264 1960
rect 3258 1955 3259 1959
rect 3263 1955 3264 1959
rect 3258 1954 3264 1955
rect 2655 1940 2659 1941
rect 2655 1935 2659 1936
rect 3151 1940 3155 1941
rect 3151 1935 3155 1936
rect 2406 1927 2412 1928
rect 2406 1923 2407 1927
rect 2411 1923 2412 1927
rect 2406 1922 2412 1923
rect 2622 1927 2628 1928
rect 2622 1923 2623 1927
rect 2627 1923 2628 1927
rect 2622 1922 2628 1923
rect 2194 1915 2200 1916
rect 2194 1911 2195 1915
rect 2199 1911 2200 1915
rect 2408 1911 2410 1922
rect 2624 1911 2626 1922
rect 2656 1916 2658 1935
rect 2822 1927 2828 1928
rect 2822 1923 2823 1927
rect 2827 1923 2828 1927
rect 3006 1927 3012 1928
rect 2822 1922 2828 1923
rect 2951 1924 2955 1925
rect 2654 1915 2660 1916
rect 2654 1911 2655 1915
rect 2659 1911 2660 1915
rect 2824 1911 2826 1922
rect 3006 1923 3007 1927
rect 3011 1923 3012 1927
rect 3006 1922 3012 1923
rect 3174 1927 3180 1928
rect 3174 1923 3175 1927
rect 3179 1923 3180 1927
rect 3260 1925 3262 1954
rect 3342 1927 3348 1928
rect 3174 1922 3180 1923
rect 3259 1924 3263 1925
rect 2951 1919 2955 1920
rect 2071 1910 2075 1911
rect 2071 1905 2075 1906
rect 2167 1910 2171 1911
rect 2194 1910 2200 1911
rect 2295 1910 2299 1911
rect 2167 1905 2171 1906
rect 2295 1905 2299 1906
rect 2407 1910 2411 1911
rect 2407 1905 2411 1906
rect 2447 1910 2451 1911
rect 2447 1905 2451 1906
rect 2607 1910 2611 1911
rect 2607 1905 2611 1906
rect 2623 1910 2627 1911
rect 2654 1910 2660 1911
rect 2767 1910 2771 1911
rect 2623 1905 2627 1906
rect 2767 1905 2771 1906
rect 2823 1910 2827 1911
rect 2823 1905 2827 1906
rect 2919 1910 2923 1911
rect 2919 1905 2923 1906
rect 2010 1903 2016 1904
rect 2010 1899 2011 1903
rect 2015 1899 2016 1903
rect 2010 1898 2016 1899
rect 2072 1894 2074 1905
rect 2110 1903 2116 1904
rect 2110 1899 2111 1903
rect 2115 1899 2116 1903
rect 2110 1898 2116 1899
rect 1982 1893 1988 1894
rect 1982 1889 1983 1893
rect 1987 1889 1988 1893
rect 1982 1888 1988 1889
rect 2070 1893 2076 1894
rect 2070 1889 2071 1893
rect 2075 1889 2076 1893
rect 2070 1888 2076 1889
rect 1943 1884 1947 1885
rect 1862 1880 1868 1881
rect 1862 1876 1863 1880
rect 1867 1876 1868 1880
rect 1943 1879 1947 1880
rect 1862 1875 1868 1876
rect 1822 1868 1828 1869
rect 1666 1867 1672 1868
rect 1666 1863 1667 1867
rect 1671 1863 1672 1867
rect 1822 1864 1823 1868
rect 1827 1864 1828 1868
rect 1822 1863 1828 1864
rect 1862 1863 1868 1864
rect 1666 1862 1672 1863
rect 1862 1859 1863 1863
rect 1867 1859 1868 1863
rect 1862 1858 1868 1859
rect 1822 1851 1828 1852
rect 1822 1847 1823 1851
rect 1827 1847 1828 1851
rect 1822 1846 1828 1847
rect 1118 1841 1124 1842
rect 1118 1837 1119 1841
rect 1123 1837 1124 1841
rect 1118 1836 1124 1837
rect 1286 1841 1292 1842
rect 1286 1837 1287 1841
rect 1291 1837 1292 1841
rect 1286 1836 1292 1837
rect 1446 1841 1452 1842
rect 1446 1837 1447 1841
rect 1451 1837 1452 1841
rect 1446 1836 1452 1837
rect 1598 1841 1604 1842
rect 1598 1837 1599 1841
rect 1603 1837 1604 1841
rect 1598 1836 1604 1837
rect 1726 1841 1732 1842
rect 1726 1837 1727 1841
rect 1731 1837 1732 1841
rect 1726 1836 1732 1837
rect 1120 1831 1122 1836
rect 1288 1831 1290 1836
rect 1448 1831 1450 1836
rect 1600 1831 1602 1836
rect 1728 1831 1730 1836
rect 1766 1835 1772 1836
rect 1766 1831 1767 1835
rect 1771 1831 1772 1835
rect 1824 1831 1826 1846
rect 1864 1839 1866 1858
rect 1886 1853 1892 1854
rect 1886 1849 1887 1853
rect 1891 1849 1892 1853
rect 1886 1848 1892 1849
rect 1974 1853 1980 1854
rect 1974 1849 1975 1853
rect 1979 1849 1980 1853
rect 1974 1848 1980 1849
rect 2062 1853 2068 1854
rect 2062 1849 2063 1853
rect 2067 1849 2068 1853
rect 2062 1848 2068 1849
rect 1888 1839 1890 1848
rect 1976 1839 1978 1848
rect 2064 1839 2066 1848
rect 1863 1838 1867 1839
rect 1863 1833 1867 1834
rect 1887 1838 1891 1839
rect 1887 1833 1891 1834
rect 1975 1838 1979 1839
rect 1975 1833 1979 1834
rect 1999 1838 2003 1839
rect 1999 1833 2003 1834
rect 2063 1838 2067 1839
rect 2063 1833 2067 1834
rect 1079 1830 1083 1831
rect 1079 1825 1083 1826
rect 1119 1830 1123 1831
rect 1119 1825 1123 1826
rect 1223 1830 1227 1831
rect 1223 1825 1227 1826
rect 1287 1830 1291 1831
rect 1287 1825 1291 1826
rect 1359 1830 1363 1831
rect 1359 1825 1363 1826
rect 1447 1830 1451 1831
rect 1447 1825 1451 1826
rect 1487 1830 1491 1831
rect 1487 1825 1491 1826
rect 1599 1830 1603 1831
rect 1599 1825 1603 1826
rect 1615 1830 1619 1831
rect 1615 1825 1619 1826
rect 1727 1830 1731 1831
rect 1766 1830 1772 1831
rect 1823 1830 1827 1831
rect 1727 1825 1731 1826
rect 1080 1820 1082 1825
rect 1224 1820 1226 1825
rect 1360 1820 1362 1825
rect 1488 1820 1490 1825
rect 1616 1820 1618 1825
rect 1728 1820 1730 1825
rect 1078 1819 1084 1820
rect 1078 1815 1079 1819
rect 1083 1815 1084 1819
rect 1078 1814 1084 1815
rect 1222 1819 1228 1820
rect 1222 1815 1223 1819
rect 1227 1815 1228 1819
rect 1222 1814 1228 1815
rect 1358 1819 1364 1820
rect 1358 1815 1359 1819
rect 1363 1815 1364 1819
rect 1358 1814 1364 1815
rect 1486 1819 1492 1820
rect 1486 1815 1487 1819
rect 1491 1815 1492 1819
rect 1486 1814 1492 1815
rect 1614 1819 1620 1820
rect 1614 1815 1615 1819
rect 1619 1815 1620 1819
rect 1614 1814 1620 1815
rect 1726 1819 1732 1820
rect 1726 1815 1727 1819
rect 1731 1815 1732 1819
rect 1726 1814 1732 1815
rect 750 1811 756 1812
rect 750 1807 751 1811
rect 755 1807 756 1811
rect 750 1806 756 1807
rect 1030 1811 1036 1812
rect 1030 1807 1031 1811
rect 1035 1807 1036 1811
rect 1030 1806 1036 1807
rect 574 1795 580 1796
rect 574 1791 575 1795
rect 579 1791 580 1795
rect 574 1790 580 1791
rect 658 1795 664 1796
rect 658 1791 659 1795
rect 663 1791 664 1795
rect 658 1790 664 1791
rect 826 1795 832 1796
rect 826 1791 827 1795
rect 831 1791 832 1795
rect 826 1790 832 1791
rect 1146 1795 1152 1796
rect 1146 1791 1147 1795
rect 1151 1791 1152 1795
rect 1146 1790 1152 1791
rect 1290 1795 1296 1796
rect 1290 1791 1291 1795
rect 1295 1791 1296 1795
rect 1290 1790 1296 1791
rect 1554 1795 1560 1796
rect 1554 1791 1555 1795
rect 1559 1791 1560 1795
rect 1554 1790 1560 1791
rect 1682 1795 1688 1796
rect 1682 1791 1683 1795
rect 1687 1791 1688 1795
rect 1682 1790 1688 1791
rect 422 1779 428 1780
rect 422 1775 423 1779
rect 427 1775 428 1779
rect 422 1774 428 1775
rect 282 1767 288 1768
rect 282 1763 283 1767
rect 287 1763 288 1767
rect 282 1762 288 1763
rect 424 1759 426 1774
rect 576 1768 578 1790
rect 598 1779 604 1780
rect 598 1775 599 1779
rect 603 1775 604 1779
rect 598 1774 604 1775
rect 574 1767 580 1768
rect 574 1763 575 1767
rect 579 1763 580 1767
rect 574 1762 580 1763
rect 538 1759 544 1760
rect 600 1759 602 1774
rect 111 1758 115 1759
rect 111 1753 115 1754
rect 255 1758 259 1759
rect 255 1753 259 1754
rect 327 1758 331 1759
rect 327 1753 331 1754
rect 423 1758 427 1759
rect 423 1753 427 1754
rect 471 1758 475 1759
rect 538 1755 539 1759
rect 543 1755 544 1759
rect 538 1754 544 1755
rect 599 1758 603 1759
rect 471 1753 475 1754
rect 112 1729 114 1753
rect 328 1742 330 1753
rect 472 1742 474 1753
rect 326 1741 332 1742
rect 326 1737 327 1741
rect 331 1737 332 1741
rect 326 1736 332 1737
rect 470 1741 476 1742
rect 470 1737 471 1741
rect 475 1737 476 1741
rect 470 1736 476 1737
rect 110 1728 116 1729
rect 110 1724 111 1728
rect 115 1724 116 1728
rect 540 1724 542 1754
rect 599 1753 603 1754
rect 615 1758 619 1759
rect 615 1753 619 1754
rect 616 1742 618 1753
rect 660 1752 662 1790
rect 766 1779 772 1780
rect 766 1775 767 1779
rect 771 1775 772 1779
rect 766 1774 772 1775
rect 768 1759 770 1774
rect 828 1768 830 1790
rect 934 1779 940 1780
rect 934 1775 935 1779
rect 939 1775 940 1779
rect 934 1774 940 1775
rect 1086 1779 1092 1780
rect 1086 1775 1087 1779
rect 1091 1775 1092 1779
rect 1086 1774 1092 1775
rect 826 1767 832 1768
rect 826 1763 827 1767
rect 831 1763 832 1767
rect 826 1762 832 1763
rect 936 1759 938 1774
rect 978 1767 984 1768
rect 978 1763 979 1767
rect 983 1763 984 1767
rect 978 1762 984 1763
rect 767 1758 771 1759
rect 767 1753 771 1754
rect 919 1758 923 1759
rect 919 1753 923 1754
rect 935 1758 939 1759
rect 935 1753 939 1754
rect 658 1751 664 1752
rect 658 1747 659 1751
rect 663 1747 664 1751
rect 658 1746 664 1747
rect 768 1742 770 1753
rect 838 1751 844 1752
rect 838 1747 839 1751
rect 843 1747 844 1751
rect 838 1746 844 1747
rect 614 1741 620 1742
rect 614 1737 615 1741
rect 619 1737 620 1741
rect 614 1736 620 1737
rect 766 1741 772 1742
rect 766 1737 767 1741
rect 771 1737 772 1741
rect 766 1736 772 1737
rect 110 1723 116 1724
rect 538 1723 544 1724
rect 538 1719 539 1723
rect 543 1719 544 1723
rect 538 1718 544 1719
rect 110 1711 116 1712
rect 110 1707 111 1711
rect 115 1707 116 1711
rect 110 1706 116 1707
rect 614 1711 620 1712
rect 614 1707 615 1711
rect 619 1707 620 1711
rect 614 1706 620 1707
rect 112 1687 114 1706
rect 318 1701 324 1702
rect 318 1697 319 1701
rect 323 1697 324 1701
rect 318 1696 324 1697
rect 462 1701 468 1702
rect 462 1697 463 1701
rect 467 1697 468 1701
rect 462 1696 468 1697
rect 606 1701 612 1702
rect 606 1697 607 1701
rect 611 1697 612 1701
rect 606 1696 612 1697
rect 320 1687 322 1696
rect 464 1687 466 1696
rect 608 1687 610 1696
rect 111 1686 115 1687
rect 111 1681 115 1682
rect 311 1686 315 1687
rect 311 1681 315 1682
rect 319 1686 323 1687
rect 319 1681 323 1682
rect 447 1686 451 1687
rect 447 1681 451 1682
rect 463 1686 467 1687
rect 463 1681 467 1682
rect 591 1686 595 1687
rect 591 1681 595 1682
rect 607 1686 611 1687
rect 607 1681 611 1682
rect 112 1666 114 1681
rect 312 1676 314 1681
rect 448 1676 450 1681
rect 592 1676 594 1681
rect 310 1675 316 1676
rect 310 1671 311 1675
rect 315 1671 316 1675
rect 310 1670 316 1671
rect 446 1675 452 1676
rect 446 1671 447 1675
rect 451 1671 452 1675
rect 446 1670 452 1671
rect 590 1675 596 1676
rect 590 1671 591 1675
rect 595 1671 596 1675
rect 590 1670 596 1671
rect 110 1665 116 1666
rect 110 1661 111 1665
rect 115 1661 116 1665
rect 110 1660 116 1661
rect 254 1651 260 1652
rect 110 1648 116 1649
rect 110 1644 111 1648
rect 115 1644 116 1648
rect 254 1647 255 1651
rect 259 1647 260 1651
rect 254 1646 260 1647
rect 378 1651 384 1652
rect 378 1647 379 1651
rect 383 1647 384 1651
rect 378 1646 384 1647
rect 514 1651 520 1652
rect 514 1647 515 1651
rect 519 1647 520 1651
rect 514 1646 520 1647
rect 110 1643 116 1644
rect 112 1611 114 1643
rect 111 1610 115 1611
rect 111 1605 115 1606
rect 223 1610 227 1611
rect 223 1605 227 1606
rect 112 1581 114 1605
rect 224 1594 226 1605
rect 256 1604 258 1646
rect 318 1635 324 1636
rect 318 1631 319 1635
rect 323 1631 324 1635
rect 318 1630 324 1631
rect 320 1611 322 1630
rect 380 1624 382 1646
rect 454 1635 460 1636
rect 454 1631 455 1635
rect 459 1631 460 1635
rect 454 1630 460 1631
rect 378 1623 384 1624
rect 378 1619 379 1623
rect 383 1619 384 1623
rect 378 1618 384 1619
rect 456 1611 458 1630
rect 516 1624 518 1646
rect 598 1635 604 1636
rect 598 1631 599 1635
rect 603 1631 604 1635
rect 598 1630 604 1631
rect 514 1623 520 1624
rect 514 1619 515 1623
rect 519 1619 520 1623
rect 514 1618 520 1619
rect 600 1611 602 1630
rect 616 1624 618 1706
rect 758 1701 764 1702
rect 758 1697 759 1701
rect 763 1697 764 1701
rect 758 1696 764 1697
rect 760 1687 762 1696
rect 735 1686 739 1687
rect 735 1681 739 1682
rect 759 1686 763 1687
rect 759 1681 763 1682
rect 736 1676 738 1681
rect 734 1675 740 1676
rect 734 1671 735 1675
rect 739 1671 740 1675
rect 734 1670 740 1671
rect 840 1668 842 1746
rect 920 1742 922 1753
rect 918 1741 924 1742
rect 918 1737 919 1741
rect 923 1737 924 1741
rect 918 1736 924 1737
rect 980 1728 982 1762
rect 1088 1759 1090 1774
rect 1148 1768 1150 1790
rect 1230 1779 1236 1780
rect 1230 1775 1231 1779
rect 1235 1775 1236 1779
rect 1230 1774 1236 1775
rect 1146 1767 1152 1768
rect 1146 1763 1147 1767
rect 1151 1763 1152 1767
rect 1146 1762 1152 1763
rect 1232 1759 1234 1774
rect 1292 1768 1294 1790
rect 1366 1779 1372 1780
rect 1366 1775 1367 1779
rect 1371 1775 1372 1779
rect 1366 1774 1372 1775
rect 1494 1779 1500 1780
rect 1494 1775 1495 1779
rect 1499 1775 1500 1779
rect 1494 1774 1500 1775
rect 1290 1767 1296 1768
rect 1290 1763 1291 1767
rect 1295 1763 1296 1767
rect 1290 1762 1296 1763
rect 1368 1759 1370 1774
rect 1434 1767 1440 1768
rect 1434 1763 1435 1767
rect 1439 1763 1440 1767
rect 1434 1762 1440 1763
rect 1071 1758 1075 1759
rect 1071 1753 1075 1754
rect 1087 1758 1091 1759
rect 1087 1753 1091 1754
rect 1223 1758 1227 1759
rect 1223 1753 1227 1754
rect 1231 1758 1235 1759
rect 1231 1753 1235 1754
rect 1367 1758 1371 1759
rect 1367 1753 1371 1754
rect 1375 1758 1379 1759
rect 1375 1753 1379 1754
rect 1072 1742 1074 1753
rect 1110 1751 1116 1752
rect 1110 1747 1111 1751
rect 1115 1747 1116 1751
rect 1110 1746 1116 1747
rect 1070 1741 1076 1742
rect 1070 1737 1071 1741
rect 1075 1737 1076 1741
rect 1070 1736 1076 1737
rect 978 1727 984 1728
rect 978 1723 979 1727
rect 983 1723 984 1727
rect 978 1722 984 1723
rect 910 1701 916 1702
rect 910 1697 911 1701
rect 915 1697 916 1701
rect 910 1696 916 1697
rect 1062 1701 1068 1702
rect 1062 1697 1063 1701
rect 1067 1697 1068 1701
rect 1062 1696 1068 1697
rect 912 1687 914 1696
rect 1064 1687 1066 1696
rect 887 1686 891 1687
rect 887 1681 891 1682
rect 911 1686 915 1687
rect 911 1681 915 1682
rect 1039 1686 1043 1687
rect 1039 1681 1043 1682
rect 1063 1686 1067 1687
rect 1063 1681 1067 1682
rect 888 1676 890 1681
rect 1040 1676 1042 1681
rect 886 1675 892 1676
rect 886 1671 887 1675
rect 891 1671 892 1675
rect 886 1670 892 1671
rect 1038 1675 1044 1676
rect 1038 1671 1039 1675
rect 1043 1671 1044 1675
rect 1038 1670 1044 1671
rect 1112 1668 1114 1746
rect 1224 1742 1226 1753
rect 1376 1742 1378 1753
rect 1222 1741 1228 1742
rect 1222 1737 1223 1741
rect 1227 1737 1228 1741
rect 1222 1736 1228 1737
rect 1374 1741 1380 1742
rect 1374 1737 1375 1741
rect 1379 1737 1380 1741
rect 1374 1736 1380 1737
rect 1436 1728 1438 1762
rect 1496 1759 1498 1774
rect 1556 1768 1558 1790
rect 1562 1787 1568 1788
rect 1562 1783 1563 1787
rect 1567 1783 1568 1787
rect 1562 1782 1568 1783
rect 1554 1767 1560 1768
rect 1554 1763 1555 1767
rect 1559 1763 1560 1767
rect 1554 1762 1560 1763
rect 1495 1758 1499 1759
rect 1495 1753 1499 1754
rect 1527 1758 1531 1759
rect 1564 1756 1566 1782
rect 1622 1779 1628 1780
rect 1622 1775 1623 1779
rect 1627 1775 1628 1779
rect 1622 1774 1628 1775
rect 1624 1759 1626 1774
rect 1684 1768 1686 1790
rect 1734 1779 1740 1780
rect 1734 1775 1735 1779
rect 1739 1775 1740 1779
rect 1734 1774 1740 1775
rect 1682 1767 1688 1768
rect 1682 1763 1683 1767
rect 1687 1763 1688 1767
rect 1682 1762 1688 1763
rect 1736 1759 1738 1774
rect 1768 1768 1770 1830
rect 1823 1825 1827 1826
rect 1824 1810 1826 1825
rect 1864 1818 1866 1833
rect 2000 1828 2002 1833
rect 1998 1827 2004 1828
rect 1998 1823 1999 1827
rect 2003 1823 2004 1827
rect 1998 1822 2004 1823
rect 2112 1820 2114 1898
rect 2168 1894 2170 1905
rect 2296 1894 2298 1905
rect 2448 1894 2450 1905
rect 2608 1894 2610 1905
rect 2768 1894 2770 1905
rect 2920 1894 2922 1905
rect 2952 1904 2954 1919
rect 3008 1911 3010 1922
rect 3176 1911 3178 1922
rect 3342 1923 3343 1927
rect 3347 1923 3348 1927
rect 3342 1922 3348 1923
rect 3259 1919 3263 1920
rect 3344 1911 3346 1922
rect 3007 1910 3011 1911
rect 3007 1905 3011 1906
rect 3071 1910 3075 1911
rect 3071 1905 3075 1906
rect 3175 1910 3179 1911
rect 3175 1905 3179 1906
rect 3215 1910 3219 1911
rect 3215 1905 3219 1906
rect 3343 1910 3347 1911
rect 3343 1905 3347 1906
rect 3359 1910 3363 1911
rect 3359 1905 3363 1906
rect 2950 1903 2956 1904
rect 2950 1899 2951 1903
rect 2955 1899 2956 1903
rect 2950 1898 2956 1899
rect 3072 1894 3074 1905
rect 3216 1894 3218 1905
rect 3360 1894 3362 1905
rect 2166 1893 2172 1894
rect 2166 1889 2167 1893
rect 2171 1889 2172 1893
rect 2166 1888 2172 1889
rect 2294 1893 2300 1894
rect 2294 1889 2295 1893
rect 2299 1889 2300 1893
rect 2294 1888 2300 1889
rect 2446 1893 2452 1894
rect 2446 1889 2447 1893
rect 2451 1889 2452 1893
rect 2446 1888 2452 1889
rect 2606 1893 2612 1894
rect 2606 1889 2607 1893
rect 2611 1889 2612 1893
rect 2606 1888 2612 1889
rect 2766 1893 2772 1894
rect 2766 1889 2767 1893
rect 2771 1889 2772 1893
rect 2766 1888 2772 1889
rect 2918 1893 2924 1894
rect 2918 1889 2919 1893
rect 2923 1889 2924 1893
rect 2918 1888 2924 1889
rect 3070 1893 3076 1894
rect 3070 1889 3071 1893
rect 3075 1889 3076 1893
rect 3070 1888 3076 1889
rect 3214 1893 3220 1894
rect 3214 1889 3215 1893
rect 3219 1889 3220 1893
rect 3214 1888 3220 1889
rect 3358 1893 3364 1894
rect 3358 1889 3359 1893
rect 3363 1889 3364 1893
rect 3358 1888 3364 1889
rect 2403 1884 2407 1885
rect 3420 1880 3422 2042
rect 3440 2038 3442 2049
rect 3438 2037 3444 2038
rect 3438 2033 3439 2037
rect 3443 2033 3444 2037
rect 3438 2032 3444 2033
rect 3430 1997 3436 1998
rect 3430 1993 3431 1997
rect 3435 1993 3436 1997
rect 3430 1992 3436 1993
rect 3432 1979 3434 1992
rect 3431 1978 3435 1979
rect 3431 1973 3435 1974
rect 3479 1978 3483 1979
rect 3479 1973 3483 1974
rect 3480 1968 3482 1973
rect 3478 1967 3484 1968
rect 3478 1963 3479 1967
rect 3483 1963 3484 1967
rect 3478 1962 3484 1963
rect 3546 1943 3552 1944
rect 3546 1939 3547 1943
rect 3551 1939 3552 1943
rect 3546 1938 3552 1939
rect 3486 1927 3492 1928
rect 3486 1923 3487 1927
rect 3491 1923 3492 1927
rect 3486 1922 3492 1923
rect 3488 1911 3490 1922
rect 3487 1910 3491 1911
rect 3487 1905 3491 1906
rect 3426 1903 3432 1904
rect 3426 1899 3427 1903
rect 3431 1899 3432 1903
rect 3426 1898 3432 1899
rect 2403 1879 2407 1880
rect 3418 1879 3424 1880
rect 2404 1876 2406 1879
rect 2402 1875 2408 1876
rect 2402 1871 2403 1875
rect 2407 1871 2408 1875
rect 3418 1875 3419 1879
rect 3423 1875 3424 1879
rect 3428 1876 3430 1898
rect 3488 1894 3490 1905
rect 3548 1904 3550 1938
rect 3556 1916 3558 2086
rect 3574 2084 3575 2088
rect 3579 2084 3580 2088
rect 3574 2083 3580 2084
rect 3576 2055 3578 2083
rect 3575 2054 3579 2055
rect 3575 2049 3579 2050
rect 3576 2025 3578 2049
rect 3574 2024 3580 2025
rect 3574 2020 3575 2024
rect 3579 2020 3580 2024
rect 3574 2019 3580 2020
rect 3574 2007 3580 2008
rect 3574 2003 3575 2007
rect 3579 2003 3580 2007
rect 3574 2002 3580 2003
rect 3576 1979 3578 2002
rect 3575 1978 3579 1979
rect 3575 1973 3579 1974
rect 3576 1958 3578 1973
rect 3574 1957 3580 1958
rect 3574 1953 3575 1957
rect 3579 1953 3580 1957
rect 3574 1952 3580 1953
rect 3574 1940 3580 1941
rect 3574 1936 3575 1940
rect 3579 1936 3580 1940
rect 3574 1935 3580 1936
rect 3554 1915 3560 1916
rect 3554 1911 3555 1915
rect 3559 1911 3560 1915
rect 3576 1911 3578 1935
rect 3554 1910 3560 1911
rect 3575 1910 3579 1911
rect 3575 1905 3579 1906
rect 3546 1903 3552 1904
rect 3546 1899 3547 1903
rect 3551 1899 3552 1903
rect 3546 1898 3552 1899
rect 3486 1893 3492 1894
rect 3486 1889 3487 1893
rect 3491 1889 3492 1893
rect 3486 1888 3492 1889
rect 3576 1881 3578 1905
rect 3574 1880 3580 1881
rect 3574 1876 3575 1880
rect 3579 1876 3580 1880
rect 3418 1874 3424 1875
rect 3426 1875 3432 1876
rect 3574 1875 3580 1876
rect 2402 1870 2408 1871
rect 3426 1871 3427 1875
rect 3431 1871 3432 1875
rect 3426 1870 3432 1871
rect 2674 1863 2680 1864
rect 2674 1859 2675 1863
rect 2679 1859 2680 1863
rect 2674 1858 2680 1859
rect 3574 1863 3580 1864
rect 3574 1859 3575 1863
rect 3579 1859 3580 1863
rect 3574 1858 3580 1859
rect 2158 1853 2164 1854
rect 2158 1849 2159 1853
rect 2163 1849 2164 1853
rect 2158 1848 2164 1849
rect 2286 1853 2292 1854
rect 2286 1849 2287 1853
rect 2291 1849 2292 1853
rect 2286 1848 2292 1849
rect 2438 1853 2444 1854
rect 2438 1849 2439 1853
rect 2443 1849 2444 1853
rect 2438 1848 2444 1849
rect 2598 1853 2604 1854
rect 2598 1849 2599 1853
rect 2603 1849 2604 1853
rect 2598 1848 2604 1849
rect 2160 1839 2162 1848
rect 2288 1839 2290 1848
rect 2440 1839 2442 1848
rect 2600 1839 2602 1848
rect 2159 1838 2163 1839
rect 2159 1833 2163 1834
rect 2223 1838 2227 1839
rect 2223 1833 2227 1834
rect 2287 1838 2291 1839
rect 2287 1833 2291 1834
rect 2439 1838 2443 1839
rect 2439 1833 2443 1834
rect 2599 1838 2603 1839
rect 2599 1833 2603 1834
rect 2639 1838 2643 1839
rect 2639 1833 2643 1834
rect 2224 1828 2226 1833
rect 2440 1828 2442 1833
rect 2640 1828 2642 1833
rect 2222 1827 2228 1828
rect 2222 1823 2223 1827
rect 2227 1823 2228 1827
rect 2222 1822 2228 1823
rect 2438 1827 2444 1828
rect 2438 1823 2439 1827
rect 2443 1823 2444 1827
rect 2438 1822 2444 1823
rect 2638 1827 2644 1828
rect 2638 1823 2639 1827
rect 2643 1823 2644 1827
rect 2638 1822 2644 1823
rect 2110 1819 2116 1820
rect 1862 1817 1868 1818
rect 1862 1813 1863 1817
rect 1867 1813 1868 1817
rect 2110 1815 2111 1819
rect 2115 1815 2116 1819
rect 2110 1814 2116 1815
rect 1862 1812 1868 1813
rect 1822 1809 1828 1810
rect 1822 1805 1823 1809
rect 1827 1805 1828 1809
rect 1822 1804 1828 1805
rect 1862 1800 1868 1801
rect 1862 1796 1863 1800
rect 1867 1796 1868 1800
rect 2676 1797 2678 1858
rect 2758 1853 2764 1854
rect 2758 1849 2759 1853
rect 2763 1849 2764 1853
rect 2758 1848 2764 1849
rect 2910 1853 2916 1854
rect 2910 1849 2911 1853
rect 2915 1849 2916 1853
rect 2910 1848 2916 1849
rect 3062 1853 3068 1854
rect 3062 1849 3063 1853
rect 3067 1849 3068 1853
rect 3062 1848 3068 1849
rect 3206 1853 3212 1854
rect 3206 1849 3207 1853
rect 3211 1849 3212 1853
rect 3206 1848 3212 1849
rect 3350 1853 3356 1854
rect 3350 1849 3351 1853
rect 3355 1849 3356 1853
rect 3350 1848 3356 1849
rect 3478 1853 3484 1854
rect 3478 1849 3479 1853
rect 3483 1849 3484 1853
rect 3478 1848 3484 1849
rect 2760 1839 2762 1848
rect 2912 1839 2914 1848
rect 3064 1839 3066 1848
rect 3208 1839 3210 1848
rect 3352 1839 3354 1848
rect 3480 1839 3482 1848
rect 3576 1839 3578 1858
rect 2759 1838 2763 1839
rect 2759 1833 2763 1834
rect 2831 1838 2835 1839
rect 2831 1833 2835 1834
rect 2911 1838 2915 1839
rect 2911 1833 2915 1834
rect 3015 1838 3019 1839
rect 3015 1833 3019 1834
rect 3063 1838 3067 1839
rect 3063 1833 3067 1834
rect 3199 1838 3203 1839
rect 3199 1833 3203 1834
rect 3207 1838 3211 1839
rect 3207 1833 3211 1834
rect 3351 1838 3355 1839
rect 3351 1833 3355 1834
rect 3391 1838 3395 1839
rect 3391 1833 3395 1834
rect 3479 1838 3483 1839
rect 3479 1833 3483 1834
rect 3575 1838 3579 1839
rect 3575 1833 3579 1834
rect 2832 1828 2834 1833
rect 3016 1828 3018 1833
rect 3200 1828 3202 1833
rect 3392 1828 3394 1833
rect 2830 1827 2836 1828
rect 2830 1823 2831 1827
rect 2835 1823 2836 1827
rect 2830 1822 2836 1823
rect 3014 1827 3020 1828
rect 3014 1823 3015 1827
rect 3019 1823 3020 1827
rect 3014 1822 3020 1823
rect 3198 1827 3204 1828
rect 3198 1823 3199 1827
rect 3203 1823 3204 1827
rect 3198 1822 3204 1823
rect 3390 1827 3396 1828
rect 3390 1823 3391 1827
rect 3395 1823 3396 1827
rect 3390 1822 3396 1823
rect 2718 1819 2724 1820
rect 2718 1815 2719 1819
rect 2723 1815 2724 1819
rect 3576 1818 3578 1833
rect 2718 1814 2724 1815
rect 3574 1817 3580 1818
rect 1862 1795 1868 1796
rect 2263 1796 2267 1797
rect 1822 1792 1828 1793
rect 1822 1788 1823 1792
rect 1827 1788 1828 1792
rect 1822 1787 1828 1788
rect 1766 1767 1772 1768
rect 1766 1763 1767 1767
rect 1771 1763 1772 1767
rect 1766 1762 1772 1763
rect 1824 1759 1826 1787
rect 1864 1767 1866 1795
rect 2263 1791 2267 1792
rect 2675 1796 2679 1797
rect 2675 1791 2679 1792
rect 2006 1787 2012 1788
rect 2006 1783 2007 1787
rect 2011 1783 2012 1787
rect 2006 1782 2012 1783
rect 2230 1787 2236 1788
rect 2230 1783 2231 1787
rect 2235 1783 2236 1787
rect 2230 1782 2236 1783
rect 2008 1767 2010 1782
rect 2232 1767 2234 1782
rect 2264 1776 2266 1791
rect 2446 1787 2452 1788
rect 2446 1783 2447 1787
rect 2451 1783 2452 1787
rect 2446 1782 2452 1783
rect 2646 1787 2652 1788
rect 2646 1783 2647 1787
rect 2651 1783 2652 1787
rect 2646 1782 2652 1783
rect 2262 1775 2268 1776
rect 2262 1771 2263 1775
rect 2267 1771 2268 1775
rect 2262 1770 2268 1771
rect 2448 1767 2450 1782
rect 2479 1780 2483 1781
rect 2478 1775 2484 1776
rect 2478 1771 2479 1775
rect 2483 1771 2484 1775
rect 2478 1770 2484 1771
rect 2648 1767 2650 1782
rect 2720 1781 2722 1814
rect 3574 1813 3575 1817
rect 3579 1813 3580 1817
rect 3574 1812 3580 1813
rect 2818 1803 2824 1804
rect 2818 1799 2819 1803
rect 2823 1799 2824 1803
rect 2818 1798 2824 1799
rect 2898 1803 2904 1804
rect 2898 1799 2899 1803
rect 2903 1799 2904 1803
rect 2898 1798 2904 1799
rect 3082 1803 3088 1804
rect 3082 1799 3083 1803
rect 3087 1799 3088 1803
rect 3082 1798 3088 1799
rect 3458 1803 3464 1804
rect 3458 1799 3459 1803
rect 3463 1799 3464 1803
rect 3458 1798 3464 1799
rect 3574 1800 3580 1801
rect 2719 1780 2723 1781
rect 2719 1775 2723 1776
rect 1863 1766 1867 1767
rect 1863 1761 1867 1762
rect 1943 1766 1947 1767
rect 1943 1761 1947 1762
rect 2007 1766 2011 1767
rect 2007 1761 2011 1762
rect 2087 1766 2091 1767
rect 2087 1761 2091 1762
rect 2231 1766 2235 1767
rect 2231 1761 2235 1762
rect 2247 1766 2251 1767
rect 2247 1761 2251 1762
rect 2415 1766 2419 1767
rect 2415 1761 2419 1762
rect 2447 1766 2451 1767
rect 2447 1761 2451 1762
rect 2599 1766 2603 1767
rect 2599 1761 2603 1762
rect 2647 1766 2651 1767
rect 2647 1761 2651 1762
rect 2791 1766 2795 1767
rect 2791 1761 2795 1762
rect 1623 1758 1627 1759
rect 1527 1753 1531 1754
rect 1562 1755 1568 1756
rect 1528 1742 1530 1753
rect 1562 1751 1563 1755
rect 1567 1751 1568 1755
rect 1623 1753 1627 1754
rect 1687 1758 1691 1759
rect 1687 1753 1691 1754
rect 1735 1758 1739 1759
rect 1735 1753 1739 1754
rect 1823 1758 1827 1759
rect 1823 1753 1827 1754
rect 1562 1750 1568 1751
rect 1688 1742 1690 1753
rect 1526 1741 1532 1742
rect 1526 1737 1527 1741
rect 1531 1737 1532 1741
rect 1526 1736 1532 1737
rect 1686 1741 1692 1742
rect 1686 1737 1687 1741
rect 1691 1737 1692 1741
rect 1686 1736 1692 1737
rect 1824 1729 1826 1753
rect 1864 1737 1866 1761
rect 1944 1750 1946 1761
rect 2034 1759 2040 1760
rect 2034 1755 2035 1759
rect 2039 1755 2040 1759
rect 2034 1754 2040 1755
rect 1942 1749 1948 1750
rect 1942 1745 1943 1749
rect 1947 1745 1948 1749
rect 1942 1744 1948 1745
rect 1862 1736 1868 1737
rect 1862 1732 1863 1736
rect 1867 1732 1868 1736
rect 2036 1732 2038 1754
rect 2088 1750 2090 1761
rect 2186 1759 2192 1760
rect 2186 1755 2187 1759
rect 2191 1755 2192 1759
rect 2186 1754 2192 1755
rect 2086 1749 2092 1750
rect 2086 1745 2087 1749
rect 2091 1745 2092 1749
rect 2086 1744 2092 1745
rect 2188 1732 2190 1754
rect 2248 1750 2250 1761
rect 2416 1750 2418 1761
rect 2600 1750 2602 1761
rect 2792 1750 2794 1761
rect 2820 1760 2822 1798
rect 2838 1787 2844 1788
rect 2838 1783 2839 1787
rect 2843 1783 2844 1787
rect 2838 1782 2844 1783
rect 2840 1767 2842 1782
rect 2900 1776 2902 1798
rect 3022 1787 3028 1788
rect 3022 1783 3023 1787
rect 3027 1783 3028 1787
rect 3022 1782 3028 1783
rect 2898 1775 2904 1776
rect 2898 1771 2899 1775
rect 2903 1771 2904 1775
rect 2898 1770 2904 1771
rect 3024 1767 3026 1782
rect 3084 1776 3086 1798
rect 3206 1787 3212 1788
rect 3206 1783 3207 1787
rect 3211 1783 3212 1787
rect 3206 1782 3212 1783
rect 3398 1787 3404 1788
rect 3398 1783 3399 1787
rect 3403 1783 3404 1787
rect 3398 1782 3404 1783
rect 3082 1775 3088 1776
rect 3082 1771 3083 1775
rect 3087 1771 3088 1775
rect 3082 1770 3088 1771
rect 3208 1767 3210 1782
rect 3258 1775 3264 1776
rect 3258 1771 3259 1775
rect 3263 1771 3264 1775
rect 3258 1770 3264 1771
rect 2839 1766 2843 1767
rect 2839 1761 2843 1762
rect 2991 1766 2995 1767
rect 2991 1761 2995 1762
rect 3023 1766 3027 1767
rect 3023 1761 3027 1762
rect 3199 1766 3203 1767
rect 3199 1761 3203 1762
rect 3207 1766 3211 1767
rect 3207 1761 3211 1762
rect 2818 1759 2824 1760
rect 2818 1755 2819 1759
rect 2823 1755 2824 1759
rect 2818 1754 2824 1755
rect 2992 1750 2994 1761
rect 3200 1750 3202 1761
rect 3230 1759 3236 1760
rect 3230 1755 3231 1759
rect 3235 1755 3236 1759
rect 3230 1754 3236 1755
rect 2246 1749 2252 1750
rect 2246 1745 2247 1749
rect 2251 1745 2252 1749
rect 2246 1744 2252 1745
rect 2414 1749 2420 1750
rect 2414 1745 2415 1749
rect 2419 1745 2420 1749
rect 2414 1744 2420 1745
rect 2598 1749 2604 1750
rect 2598 1745 2599 1749
rect 2603 1745 2604 1749
rect 2598 1744 2604 1745
rect 2790 1749 2796 1750
rect 2790 1745 2791 1749
rect 2795 1745 2796 1749
rect 2790 1744 2796 1745
rect 2990 1749 2996 1750
rect 2990 1745 2991 1749
rect 2995 1745 2996 1749
rect 2990 1744 2996 1745
rect 3198 1749 3204 1750
rect 3198 1745 3199 1749
rect 3203 1745 3204 1749
rect 3198 1744 3204 1745
rect 1862 1731 1868 1732
rect 2034 1731 2040 1732
rect 1822 1728 1828 1729
rect 1434 1727 1440 1728
rect 1434 1723 1435 1727
rect 1439 1723 1440 1727
rect 1822 1724 1823 1728
rect 1827 1724 1828 1728
rect 2034 1727 2035 1731
rect 2039 1727 2040 1731
rect 2034 1726 2040 1727
rect 2186 1731 2192 1732
rect 2186 1727 2187 1731
rect 2191 1727 2192 1731
rect 2186 1726 2192 1727
rect 1822 1723 1828 1724
rect 1434 1722 1440 1723
rect 1862 1719 1868 1720
rect 1862 1715 1863 1719
rect 1867 1715 1868 1719
rect 1862 1714 1868 1715
rect 3082 1719 3088 1720
rect 3082 1715 3083 1719
rect 3087 1715 3088 1719
rect 3082 1714 3088 1715
rect 1686 1711 1692 1712
rect 1686 1707 1687 1711
rect 1691 1707 1692 1711
rect 1686 1706 1692 1707
rect 1822 1711 1828 1712
rect 1822 1707 1823 1711
rect 1827 1707 1828 1711
rect 1822 1706 1828 1707
rect 1214 1701 1220 1702
rect 1214 1697 1215 1701
rect 1219 1697 1220 1701
rect 1214 1696 1220 1697
rect 1366 1701 1372 1702
rect 1366 1697 1367 1701
rect 1371 1697 1372 1701
rect 1366 1696 1372 1697
rect 1518 1701 1524 1702
rect 1518 1697 1519 1701
rect 1523 1697 1524 1701
rect 1518 1696 1524 1697
rect 1678 1701 1684 1702
rect 1678 1697 1679 1701
rect 1683 1697 1684 1701
rect 1678 1696 1684 1697
rect 1216 1687 1218 1696
rect 1368 1687 1370 1696
rect 1520 1687 1522 1696
rect 1680 1687 1682 1696
rect 1191 1686 1195 1687
rect 1191 1681 1195 1682
rect 1215 1686 1219 1687
rect 1215 1681 1219 1682
rect 1343 1686 1347 1687
rect 1343 1681 1347 1682
rect 1367 1686 1371 1687
rect 1367 1681 1371 1682
rect 1495 1686 1499 1687
rect 1495 1681 1499 1682
rect 1519 1686 1523 1687
rect 1519 1681 1523 1682
rect 1647 1686 1651 1687
rect 1647 1681 1651 1682
rect 1679 1686 1683 1687
rect 1679 1681 1683 1682
rect 1192 1676 1194 1681
rect 1344 1676 1346 1681
rect 1496 1676 1498 1681
rect 1648 1676 1650 1681
rect 1190 1675 1196 1676
rect 1190 1671 1191 1675
rect 1195 1671 1196 1675
rect 1190 1670 1196 1671
rect 1342 1675 1348 1676
rect 1342 1671 1343 1675
rect 1347 1671 1348 1675
rect 1342 1670 1348 1671
rect 1494 1675 1500 1676
rect 1494 1671 1495 1675
rect 1499 1671 1500 1675
rect 1494 1670 1500 1671
rect 1646 1675 1652 1676
rect 1646 1671 1647 1675
rect 1651 1671 1652 1675
rect 1646 1670 1652 1671
rect 838 1667 844 1668
rect 838 1663 839 1667
rect 843 1663 844 1667
rect 838 1662 844 1663
rect 1110 1667 1116 1668
rect 1110 1663 1111 1667
rect 1115 1663 1116 1667
rect 1110 1662 1116 1663
rect 1142 1651 1148 1652
rect 1142 1647 1143 1651
rect 1147 1647 1148 1651
rect 1142 1646 1148 1647
rect 1410 1651 1416 1652
rect 1410 1647 1411 1651
rect 1415 1647 1416 1651
rect 1410 1646 1416 1647
rect 1562 1651 1568 1652
rect 1562 1647 1563 1651
rect 1567 1647 1568 1651
rect 1562 1646 1568 1647
rect 742 1635 748 1636
rect 742 1631 743 1635
rect 747 1631 748 1635
rect 742 1630 748 1631
rect 894 1635 900 1636
rect 894 1631 895 1635
rect 899 1631 900 1635
rect 894 1630 900 1631
rect 1046 1635 1052 1636
rect 1046 1631 1047 1635
rect 1051 1631 1052 1635
rect 1046 1630 1052 1631
rect 614 1623 620 1624
rect 614 1619 615 1623
rect 619 1619 620 1623
rect 614 1618 620 1619
rect 744 1611 746 1630
rect 750 1623 756 1624
rect 750 1619 751 1623
rect 755 1619 756 1623
rect 750 1618 756 1619
rect 319 1610 323 1611
rect 319 1605 323 1606
rect 351 1610 355 1611
rect 351 1605 355 1606
rect 455 1610 459 1611
rect 455 1605 459 1606
rect 487 1610 491 1611
rect 487 1605 491 1606
rect 599 1610 603 1611
rect 599 1605 603 1606
rect 623 1610 627 1611
rect 623 1605 627 1606
rect 743 1610 747 1611
rect 743 1605 747 1606
rect 254 1603 260 1604
rect 254 1599 255 1603
rect 259 1599 260 1603
rect 254 1598 260 1599
rect 352 1594 354 1605
rect 488 1594 490 1605
rect 624 1594 626 1605
rect 650 1603 656 1604
rect 650 1599 651 1603
rect 655 1599 656 1603
rect 650 1598 656 1599
rect 222 1593 228 1594
rect 222 1589 223 1593
rect 227 1589 228 1593
rect 222 1588 228 1589
rect 350 1593 356 1594
rect 350 1589 351 1593
rect 355 1589 356 1593
rect 350 1588 356 1589
rect 486 1593 492 1594
rect 486 1589 487 1593
rect 491 1589 492 1593
rect 486 1588 492 1589
rect 622 1593 628 1594
rect 622 1589 623 1593
rect 627 1589 628 1593
rect 622 1588 628 1589
rect 110 1580 116 1581
rect 110 1576 111 1580
rect 115 1576 116 1580
rect 110 1575 116 1576
rect 110 1563 116 1564
rect 110 1559 111 1563
rect 115 1559 116 1563
rect 110 1558 116 1559
rect 462 1563 468 1564
rect 462 1559 463 1563
rect 467 1559 468 1563
rect 462 1558 468 1559
rect 112 1539 114 1558
rect 214 1553 220 1554
rect 214 1549 215 1553
rect 219 1549 220 1553
rect 214 1548 220 1549
rect 342 1553 348 1554
rect 342 1549 343 1553
rect 347 1549 348 1553
rect 342 1548 348 1549
rect 216 1539 218 1548
rect 344 1539 346 1548
rect 111 1538 115 1539
rect 111 1533 115 1534
rect 135 1538 139 1539
rect 135 1533 139 1534
rect 215 1538 219 1539
rect 215 1533 219 1534
rect 271 1538 275 1539
rect 271 1533 275 1534
rect 343 1538 347 1539
rect 343 1533 347 1534
rect 423 1538 427 1539
rect 423 1533 427 1534
rect 112 1518 114 1533
rect 136 1528 138 1533
rect 272 1528 274 1533
rect 424 1528 426 1533
rect 134 1527 140 1528
rect 134 1523 135 1527
rect 139 1523 140 1527
rect 134 1522 140 1523
rect 270 1527 276 1528
rect 270 1523 271 1527
rect 275 1523 276 1527
rect 270 1522 276 1523
rect 422 1527 428 1528
rect 422 1523 423 1527
rect 427 1523 428 1527
rect 422 1522 428 1523
rect 110 1517 116 1518
rect 110 1513 111 1517
rect 115 1513 116 1517
rect 110 1512 116 1513
rect 338 1503 344 1504
rect 110 1500 116 1501
rect 110 1496 111 1500
rect 115 1496 116 1500
rect 338 1499 339 1503
rect 343 1499 344 1503
rect 338 1498 344 1499
rect 110 1495 116 1496
rect 198 1495 204 1496
rect 112 1463 114 1495
rect 198 1491 199 1495
rect 203 1491 204 1495
rect 198 1490 204 1491
rect 142 1487 148 1488
rect 142 1483 143 1487
rect 147 1483 148 1487
rect 142 1482 148 1483
rect 144 1463 146 1482
rect 111 1462 115 1463
rect 111 1457 115 1458
rect 143 1462 147 1463
rect 143 1457 147 1458
rect 112 1433 114 1457
rect 144 1446 146 1457
rect 200 1456 202 1490
rect 278 1487 284 1488
rect 278 1483 279 1487
rect 283 1483 284 1487
rect 278 1482 284 1483
rect 280 1463 282 1482
rect 340 1476 342 1498
rect 430 1487 436 1488
rect 430 1483 431 1487
rect 435 1483 436 1487
rect 430 1482 436 1483
rect 338 1475 344 1476
rect 338 1471 339 1475
rect 343 1471 344 1475
rect 338 1470 344 1471
rect 432 1463 434 1482
rect 464 1476 466 1558
rect 478 1553 484 1554
rect 478 1549 479 1553
rect 483 1549 484 1553
rect 478 1548 484 1549
rect 614 1553 620 1554
rect 614 1549 615 1553
rect 619 1549 620 1553
rect 614 1548 620 1549
rect 480 1539 482 1548
rect 616 1539 618 1548
rect 479 1538 483 1539
rect 479 1533 483 1534
rect 583 1538 587 1539
rect 583 1533 587 1534
rect 615 1538 619 1539
rect 615 1533 619 1534
rect 584 1528 586 1533
rect 582 1527 588 1528
rect 582 1523 583 1527
rect 587 1523 588 1527
rect 582 1522 588 1523
rect 652 1520 654 1598
rect 752 1576 754 1618
rect 896 1611 898 1630
rect 1048 1611 1050 1630
rect 1144 1624 1146 1646
rect 1198 1635 1204 1636
rect 1198 1631 1199 1635
rect 1203 1631 1204 1635
rect 1198 1630 1204 1631
rect 1350 1635 1356 1636
rect 1350 1631 1351 1635
rect 1355 1631 1356 1635
rect 1350 1630 1356 1631
rect 1142 1623 1148 1624
rect 1142 1619 1143 1623
rect 1147 1619 1148 1623
rect 1142 1618 1148 1619
rect 1200 1611 1202 1630
rect 1206 1623 1212 1624
rect 1206 1619 1207 1623
rect 1211 1619 1212 1623
rect 1206 1618 1212 1619
rect 759 1610 763 1611
rect 759 1605 763 1606
rect 895 1610 899 1611
rect 895 1605 899 1606
rect 903 1610 907 1611
rect 903 1605 907 1606
rect 1047 1610 1051 1611
rect 1047 1605 1051 1606
rect 1055 1610 1059 1611
rect 1055 1605 1059 1606
rect 1199 1610 1203 1611
rect 1199 1605 1203 1606
rect 760 1594 762 1605
rect 904 1594 906 1605
rect 954 1603 960 1604
rect 954 1599 955 1603
rect 959 1599 960 1603
rect 954 1598 960 1599
rect 758 1593 764 1594
rect 758 1589 759 1593
rect 763 1589 764 1593
rect 758 1588 764 1589
rect 902 1593 908 1594
rect 902 1589 903 1593
rect 907 1589 908 1593
rect 902 1588 908 1589
rect 750 1575 756 1576
rect 750 1571 751 1575
rect 755 1571 756 1575
rect 750 1570 756 1571
rect 750 1553 756 1554
rect 750 1549 751 1553
rect 755 1549 756 1553
rect 750 1548 756 1549
rect 894 1553 900 1554
rect 894 1549 895 1553
rect 899 1549 900 1553
rect 894 1548 900 1549
rect 752 1539 754 1548
rect 896 1539 898 1548
rect 735 1538 739 1539
rect 735 1533 739 1534
rect 751 1538 755 1539
rect 751 1533 755 1534
rect 887 1538 891 1539
rect 887 1533 891 1534
rect 895 1538 899 1539
rect 895 1533 899 1534
rect 736 1528 738 1533
rect 888 1528 890 1533
rect 734 1527 740 1528
rect 734 1523 735 1527
rect 739 1523 740 1527
rect 734 1522 740 1523
rect 886 1527 892 1528
rect 886 1523 887 1527
rect 891 1523 892 1527
rect 886 1522 892 1523
rect 956 1520 958 1598
rect 1056 1594 1058 1605
rect 1174 1603 1180 1604
rect 1174 1599 1175 1603
rect 1179 1599 1180 1603
rect 1174 1598 1180 1599
rect 1054 1593 1060 1594
rect 1054 1589 1055 1593
rect 1059 1589 1060 1593
rect 1054 1588 1060 1589
rect 1176 1580 1178 1598
rect 1174 1579 1180 1580
rect 1174 1575 1175 1579
rect 1179 1575 1180 1579
rect 1208 1576 1210 1618
rect 1352 1611 1354 1630
rect 1412 1624 1414 1646
rect 1502 1635 1508 1636
rect 1502 1631 1503 1635
rect 1507 1631 1508 1635
rect 1502 1630 1508 1631
rect 1410 1623 1416 1624
rect 1410 1619 1411 1623
rect 1415 1619 1416 1623
rect 1410 1618 1416 1619
rect 1504 1611 1506 1630
rect 1564 1624 1566 1646
rect 1654 1635 1660 1636
rect 1654 1631 1655 1635
rect 1659 1631 1660 1635
rect 1654 1630 1660 1631
rect 1562 1623 1568 1624
rect 1562 1619 1563 1623
rect 1567 1619 1568 1623
rect 1562 1618 1568 1619
rect 1656 1611 1658 1630
rect 1688 1624 1690 1706
rect 1824 1687 1826 1706
rect 1864 1695 1866 1714
rect 1934 1709 1940 1710
rect 1934 1705 1935 1709
rect 1939 1705 1940 1709
rect 1934 1704 1940 1705
rect 2078 1709 2084 1710
rect 2078 1705 2079 1709
rect 2083 1705 2084 1709
rect 2078 1704 2084 1705
rect 2238 1709 2244 1710
rect 2238 1705 2239 1709
rect 2243 1705 2244 1709
rect 2238 1704 2244 1705
rect 2406 1709 2412 1710
rect 2406 1705 2407 1709
rect 2411 1705 2412 1709
rect 2406 1704 2412 1705
rect 2590 1709 2596 1710
rect 2590 1705 2591 1709
rect 2595 1705 2596 1709
rect 2590 1704 2596 1705
rect 2782 1709 2788 1710
rect 2782 1705 2783 1709
rect 2787 1705 2788 1709
rect 2782 1704 2788 1705
rect 2982 1709 2988 1710
rect 2982 1705 2983 1709
rect 2987 1705 2988 1709
rect 2982 1704 2988 1705
rect 1936 1695 1938 1704
rect 2080 1695 2082 1704
rect 2240 1695 2242 1704
rect 2310 1703 2316 1704
rect 2310 1699 2311 1703
rect 2315 1699 2316 1703
rect 2310 1698 2316 1699
rect 1863 1694 1867 1695
rect 1863 1689 1867 1690
rect 1911 1694 1915 1695
rect 1911 1689 1915 1690
rect 1935 1694 1939 1695
rect 1935 1689 1939 1690
rect 2031 1694 2035 1695
rect 2031 1689 2035 1690
rect 2079 1694 2083 1695
rect 2079 1689 2083 1690
rect 2151 1694 2155 1695
rect 2151 1689 2155 1690
rect 2239 1694 2243 1695
rect 2239 1689 2243 1690
rect 2271 1694 2275 1695
rect 2271 1689 2275 1690
rect 1823 1686 1827 1687
rect 1823 1681 1827 1682
rect 1824 1666 1826 1681
rect 1864 1674 1866 1689
rect 1912 1684 1914 1689
rect 2032 1684 2034 1689
rect 2152 1684 2154 1689
rect 2272 1684 2274 1689
rect 1910 1683 1916 1684
rect 1910 1679 1911 1683
rect 1915 1679 1916 1683
rect 1910 1678 1916 1679
rect 2030 1683 2036 1684
rect 2030 1679 2031 1683
rect 2035 1679 2036 1683
rect 2030 1678 2036 1679
rect 2150 1683 2156 1684
rect 2150 1679 2151 1683
rect 2155 1679 2156 1683
rect 2150 1678 2156 1679
rect 2270 1683 2276 1684
rect 2270 1679 2271 1683
rect 2275 1679 2276 1683
rect 2270 1678 2276 1679
rect 1862 1673 1868 1674
rect 1862 1669 1863 1673
rect 1867 1669 1868 1673
rect 1862 1668 1868 1669
rect 1822 1665 1828 1666
rect 1822 1661 1823 1665
rect 1827 1661 1828 1665
rect 1822 1660 1828 1661
rect 1862 1656 1868 1657
rect 1862 1652 1863 1656
rect 1867 1652 1868 1656
rect 1862 1651 1868 1652
rect 1822 1648 1828 1649
rect 1822 1644 1823 1648
rect 1827 1644 1828 1648
rect 1822 1643 1828 1644
rect 1686 1623 1692 1624
rect 1686 1619 1687 1623
rect 1691 1619 1692 1623
rect 1686 1618 1692 1619
rect 1824 1611 1826 1643
rect 1864 1619 1866 1651
rect 1918 1643 1924 1644
rect 1918 1639 1919 1643
rect 1923 1639 1924 1643
rect 1918 1638 1924 1639
rect 2038 1643 2044 1644
rect 2038 1639 2039 1643
rect 2043 1639 2044 1643
rect 2038 1638 2044 1639
rect 2158 1643 2164 1644
rect 2158 1639 2159 1643
rect 2163 1639 2164 1643
rect 2158 1638 2164 1639
rect 2278 1643 2284 1644
rect 2278 1639 2279 1643
rect 2283 1639 2284 1643
rect 2278 1638 2284 1639
rect 1920 1619 1922 1638
rect 1958 1631 1964 1632
rect 1958 1627 1959 1631
rect 1963 1627 1964 1631
rect 1958 1626 1964 1627
rect 1863 1618 1867 1619
rect 1863 1613 1867 1614
rect 1895 1618 1899 1619
rect 1895 1613 1899 1614
rect 1919 1618 1923 1619
rect 1919 1613 1923 1614
rect 1215 1610 1219 1611
rect 1215 1605 1219 1606
rect 1351 1610 1355 1611
rect 1351 1605 1355 1606
rect 1375 1610 1379 1611
rect 1375 1605 1379 1606
rect 1503 1610 1507 1611
rect 1503 1605 1507 1606
rect 1543 1610 1547 1611
rect 1543 1605 1547 1606
rect 1655 1610 1659 1611
rect 1655 1605 1659 1606
rect 1823 1610 1827 1611
rect 1823 1605 1827 1606
rect 1216 1594 1218 1605
rect 1376 1594 1378 1605
rect 1544 1594 1546 1605
rect 1214 1593 1220 1594
rect 1214 1589 1215 1593
rect 1219 1589 1220 1593
rect 1214 1588 1220 1589
rect 1374 1593 1380 1594
rect 1374 1589 1375 1593
rect 1379 1589 1380 1593
rect 1374 1588 1380 1589
rect 1542 1593 1548 1594
rect 1542 1589 1543 1593
rect 1547 1589 1548 1593
rect 1542 1588 1548 1589
rect 1824 1581 1826 1605
rect 1864 1589 1866 1613
rect 1896 1602 1898 1613
rect 1894 1601 1900 1602
rect 1894 1597 1895 1601
rect 1899 1597 1900 1601
rect 1894 1596 1900 1597
rect 1862 1588 1868 1589
rect 1960 1588 1962 1626
rect 2040 1619 2042 1638
rect 2160 1619 2162 1638
rect 2280 1619 2282 1638
rect 2312 1632 2314 1698
rect 2408 1695 2410 1704
rect 2592 1695 2594 1704
rect 2784 1695 2786 1704
rect 2984 1695 2986 1704
rect 2399 1694 2403 1695
rect 2399 1689 2403 1690
rect 2407 1694 2411 1695
rect 2407 1689 2411 1690
rect 2543 1694 2547 1695
rect 2543 1689 2547 1690
rect 2591 1694 2595 1695
rect 2591 1689 2595 1690
rect 2695 1694 2699 1695
rect 2695 1689 2699 1690
rect 2783 1694 2787 1695
rect 2783 1689 2787 1690
rect 2863 1694 2867 1695
rect 2863 1689 2867 1690
rect 2983 1694 2987 1695
rect 2983 1689 2987 1690
rect 3047 1694 3051 1695
rect 3047 1689 3051 1690
rect 2400 1684 2402 1689
rect 2544 1684 2546 1689
rect 2696 1684 2698 1689
rect 2864 1684 2866 1689
rect 3048 1684 3050 1689
rect 2398 1683 2404 1684
rect 2398 1679 2399 1683
rect 2403 1679 2404 1683
rect 2398 1678 2404 1679
rect 2542 1683 2548 1684
rect 2542 1679 2543 1683
rect 2547 1679 2548 1683
rect 2542 1678 2548 1679
rect 2694 1683 2700 1684
rect 2694 1679 2695 1683
rect 2699 1679 2700 1683
rect 2694 1678 2700 1679
rect 2862 1683 2868 1684
rect 2862 1679 2863 1683
rect 2867 1679 2868 1683
rect 2862 1678 2868 1679
rect 3046 1683 3052 1684
rect 3046 1679 3047 1683
rect 3051 1679 3052 1683
rect 3046 1678 3052 1679
rect 2466 1659 2472 1660
rect 2466 1655 2467 1659
rect 2471 1655 2472 1659
rect 2466 1654 2472 1655
rect 2610 1659 2616 1660
rect 2610 1655 2611 1659
rect 2615 1655 2616 1659
rect 2610 1654 2616 1655
rect 2762 1659 2768 1660
rect 2762 1655 2763 1659
rect 2767 1655 2768 1659
rect 2762 1654 2768 1655
rect 2930 1659 2936 1660
rect 2930 1655 2931 1659
rect 2935 1655 2936 1659
rect 2930 1654 2936 1655
rect 2406 1643 2412 1644
rect 2406 1639 2407 1643
rect 2411 1639 2412 1643
rect 2406 1638 2412 1639
rect 2310 1631 2316 1632
rect 2310 1627 2311 1631
rect 2315 1627 2316 1631
rect 2310 1626 2316 1627
rect 2408 1619 2410 1638
rect 2015 1618 2019 1619
rect 2015 1613 2019 1614
rect 2039 1618 2043 1619
rect 2039 1613 2043 1614
rect 2151 1618 2155 1619
rect 2151 1613 2155 1614
rect 2159 1618 2163 1619
rect 2159 1613 2163 1614
rect 2279 1618 2283 1619
rect 2279 1613 2283 1614
rect 2287 1618 2291 1619
rect 2287 1613 2291 1614
rect 2407 1618 2411 1619
rect 2407 1613 2411 1614
rect 2431 1618 2435 1619
rect 2431 1613 2435 1614
rect 1974 1611 1980 1612
rect 1974 1607 1975 1611
rect 1979 1607 1980 1611
rect 1974 1606 1980 1607
rect 1862 1584 1863 1588
rect 1867 1584 1868 1588
rect 1862 1583 1868 1584
rect 1958 1587 1964 1588
rect 1958 1583 1959 1587
rect 1963 1583 1964 1587
rect 1976 1584 1978 1606
rect 2016 1602 2018 1613
rect 2082 1611 2088 1612
rect 2082 1607 2083 1611
rect 2087 1607 2088 1611
rect 2082 1606 2088 1607
rect 2014 1601 2020 1602
rect 2014 1597 2015 1601
rect 2019 1597 2020 1601
rect 2014 1596 2020 1597
rect 2084 1584 2086 1606
rect 2152 1602 2154 1613
rect 2288 1602 2290 1613
rect 2432 1602 2434 1613
rect 2468 1612 2470 1654
rect 2550 1643 2556 1644
rect 2550 1639 2551 1643
rect 2555 1639 2556 1643
rect 2550 1638 2556 1639
rect 2552 1619 2554 1638
rect 2612 1632 2614 1654
rect 2618 1651 2624 1652
rect 2618 1647 2619 1651
rect 2623 1647 2624 1651
rect 2618 1646 2624 1647
rect 2610 1631 2616 1632
rect 2610 1627 2611 1631
rect 2615 1627 2616 1631
rect 2610 1626 2616 1627
rect 2551 1618 2555 1619
rect 2551 1613 2555 1614
rect 2583 1618 2587 1619
rect 2620 1616 2622 1646
rect 2702 1643 2708 1644
rect 2702 1639 2703 1643
rect 2707 1639 2708 1643
rect 2702 1638 2708 1639
rect 2704 1619 2706 1638
rect 2764 1632 2766 1654
rect 2870 1643 2876 1644
rect 2870 1639 2871 1643
rect 2875 1639 2876 1643
rect 2870 1638 2876 1639
rect 2762 1631 2768 1632
rect 2762 1627 2763 1631
rect 2767 1627 2768 1631
rect 2762 1626 2768 1627
rect 2872 1619 2874 1638
rect 2932 1632 2934 1654
rect 3054 1643 3060 1644
rect 3054 1639 3055 1643
rect 3059 1639 3060 1643
rect 3054 1638 3060 1639
rect 2930 1631 2936 1632
rect 2930 1627 2931 1631
rect 2935 1627 2936 1631
rect 2930 1626 2936 1627
rect 3056 1619 3058 1638
rect 3084 1632 3086 1714
rect 3190 1709 3196 1710
rect 3190 1705 3191 1709
rect 3195 1705 3196 1709
rect 3190 1704 3196 1705
rect 3192 1695 3194 1704
rect 3191 1694 3195 1695
rect 3191 1689 3195 1690
rect 3232 1676 3234 1754
rect 3260 1736 3262 1770
rect 3400 1767 3402 1782
rect 3399 1766 3403 1767
rect 3399 1761 3403 1762
rect 3415 1766 3419 1767
rect 3415 1761 3419 1762
rect 3416 1750 3418 1761
rect 3460 1760 3462 1798
rect 3574 1796 3575 1800
rect 3579 1796 3580 1800
rect 3574 1795 3580 1796
rect 3576 1767 3578 1795
rect 3575 1766 3579 1767
rect 3575 1761 3579 1762
rect 3458 1759 3464 1760
rect 3458 1755 3459 1759
rect 3463 1755 3464 1759
rect 3458 1754 3464 1755
rect 3414 1749 3420 1750
rect 3414 1745 3415 1749
rect 3419 1745 3420 1749
rect 3414 1744 3420 1745
rect 3576 1737 3578 1761
rect 3574 1736 3580 1737
rect 3258 1735 3264 1736
rect 3258 1731 3259 1735
rect 3263 1731 3264 1735
rect 3574 1732 3575 1736
rect 3579 1732 3580 1736
rect 3574 1731 3580 1732
rect 3258 1730 3264 1731
rect 3574 1719 3580 1720
rect 3574 1715 3575 1719
rect 3579 1715 3580 1719
rect 3574 1714 3580 1715
rect 3406 1709 3412 1710
rect 3406 1705 3407 1709
rect 3411 1705 3412 1709
rect 3406 1704 3412 1705
rect 3408 1695 3410 1704
rect 3466 1703 3472 1704
rect 3466 1699 3467 1703
rect 3471 1699 3472 1703
rect 3466 1698 3472 1699
rect 3239 1694 3243 1695
rect 3239 1689 3243 1690
rect 3407 1694 3411 1695
rect 3407 1689 3411 1690
rect 3431 1694 3435 1695
rect 3431 1689 3435 1690
rect 3240 1684 3242 1689
rect 3432 1684 3434 1689
rect 3238 1683 3244 1684
rect 3238 1679 3239 1683
rect 3243 1679 3244 1683
rect 3238 1678 3244 1679
rect 3430 1683 3436 1684
rect 3430 1679 3431 1683
rect 3435 1679 3436 1683
rect 3430 1678 3436 1679
rect 3230 1675 3236 1676
rect 3230 1671 3231 1675
rect 3235 1671 3236 1675
rect 3230 1670 3236 1671
rect 3246 1643 3252 1644
rect 3246 1639 3247 1643
rect 3251 1639 3252 1643
rect 3246 1638 3252 1639
rect 3438 1643 3444 1644
rect 3438 1639 3439 1643
rect 3443 1639 3444 1643
rect 3438 1638 3444 1639
rect 3082 1631 3088 1632
rect 3082 1627 3083 1631
rect 3087 1627 3088 1631
rect 3082 1626 3088 1627
rect 3248 1619 3250 1638
rect 3270 1631 3276 1632
rect 3270 1627 3271 1631
rect 3275 1627 3276 1631
rect 3270 1626 3276 1627
rect 2703 1618 2707 1619
rect 2583 1613 2587 1614
rect 2618 1615 2624 1616
rect 2462 1611 2470 1612
rect 2462 1607 2463 1611
rect 2467 1608 2470 1611
rect 2467 1607 2468 1608
rect 2462 1606 2468 1607
rect 2584 1602 2586 1613
rect 2618 1611 2619 1615
rect 2623 1611 2624 1615
rect 2703 1613 2707 1614
rect 2743 1618 2747 1619
rect 2743 1613 2747 1614
rect 2871 1618 2875 1619
rect 2871 1613 2875 1614
rect 2911 1618 2915 1619
rect 2911 1613 2915 1614
rect 3055 1618 3059 1619
rect 3055 1613 3059 1614
rect 3095 1618 3099 1619
rect 3095 1613 3099 1614
rect 3247 1618 3251 1619
rect 3247 1613 3251 1614
rect 2618 1610 2624 1611
rect 2744 1602 2746 1613
rect 2912 1602 2914 1613
rect 3096 1602 3098 1613
rect 2150 1601 2156 1602
rect 2150 1597 2151 1601
rect 2155 1597 2156 1601
rect 2150 1596 2156 1597
rect 2286 1601 2292 1602
rect 2286 1597 2287 1601
rect 2291 1597 2292 1601
rect 2286 1596 2292 1597
rect 2430 1601 2436 1602
rect 2430 1597 2431 1601
rect 2435 1597 2436 1601
rect 2430 1596 2436 1597
rect 2582 1601 2588 1602
rect 2582 1597 2583 1601
rect 2587 1597 2588 1601
rect 2582 1596 2588 1597
rect 2742 1601 2748 1602
rect 2742 1597 2743 1601
rect 2747 1597 2748 1601
rect 2742 1596 2748 1597
rect 2910 1601 2916 1602
rect 2910 1597 2911 1601
rect 2915 1597 2916 1601
rect 2910 1596 2916 1597
rect 3094 1601 3100 1602
rect 3094 1597 3095 1601
rect 3099 1597 3100 1601
rect 3094 1596 3100 1597
rect 3272 1584 3274 1626
rect 3440 1619 3442 1638
rect 3468 1632 3470 1698
rect 3576 1695 3578 1714
rect 3575 1694 3579 1695
rect 3575 1689 3579 1690
rect 3576 1674 3578 1689
rect 3574 1673 3580 1674
rect 3574 1669 3575 1673
rect 3579 1669 3580 1673
rect 3574 1668 3580 1669
rect 3498 1659 3504 1660
rect 3498 1655 3499 1659
rect 3503 1655 3504 1659
rect 3498 1654 3504 1655
rect 3574 1656 3580 1657
rect 3466 1631 3472 1632
rect 3466 1627 3467 1631
rect 3471 1627 3472 1631
rect 3466 1626 3472 1627
rect 3279 1618 3283 1619
rect 3279 1613 3283 1614
rect 3439 1618 3443 1619
rect 3439 1613 3443 1614
rect 3471 1618 3475 1619
rect 3471 1613 3475 1614
rect 3280 1602 3282 1613
rect 3310 1611 3316 1612
rect 3310 1607 3311 1611
rect 3315 1607 3316 1611
rect 3310 1606 3316 1607
rect 3278 1601 3284 1602
rect 3278 1597 3279 1601
rect 3283 1597 3284 1601
rect 3278 1596 3284 1597
rect 1958 1582 1964 1583
rect 1974 1583 1980 1584
rect 1822 1580 1828 1581
rect 1822 1576 1823 1580
rect 1827 1576 1828 1580
rect 1974 1579 1975 1583
rect 1979 1579 1980 1583
rect 1974 1578 1980 1579
rect 2082 1583 2088 1584
rect 2082 1579 2083 1583
rect 2087 1579 2088 1583
rect 2082 1578 2088 1579
rect 3270 1583 3276 1584
rect 3270 1579 3271 1583
rect 3275 1579 3276 1583
rect 3270 1578 3276 1579
rect 1174 1574 1180 1575
rect 1206 1575 1212 1576
rect 1822 1575 1828 1576
rect 1206 1571 1207 1575
rect 1211 1571 1212 1575
rect 1206 1570 1212 1571
rect 1862 1571 1868 1572
rect 1862 1567 1863 1571
rect 1867 1567 1868 1571
rect 1862 1566 1868 1567
rect 2222 1571 2228 1572
rect 2222 1567 2223 1571
rect 2227 1567 2228 1571
rect 2222 1566 2228 1567
rect 3018 1571 3024 1572
rect 3018 1567 3019 1571
rect 3023 1567 3024 1571
rect 3018 1566 3024 1567
rect 1542 1563 1548 1564
rect 1542 1559 1543 1563
rect 1547 1559 1548 1563
rect 1542 1558 1548 1559
rect 1822 1563 1828 1564
rect 1822 1559 1823 1563
rect 1827 1559 1828 1563
rect 1822 1558 1828 1559
rect 1046 1553 1052 1554
rect 1046 1549 1047 1553
rect 1051 1549 1052 1553
rect 1046 1548 1052 1549
rect 1206 1553 1212 1554
rect 1206 1549 1207 1553
rect 1211 1549 1212 1553
rect 1206 1548 1212 1549
rect 1366 1553 1372 1554
rect 1366 1549 1367 1553
rect 1371 1549 1372 1553
rect 1366 1548 1372 1549
rect 1534 1553 1540 1554
rect 1534 1549 1535 1553
rect 1539 1549 1540 1553
rect 1534 1548 1540 1549
rect 1048 1539 1050 1548
rect 1208 1539 1210 1548
rect 1368 1539 1370 1548
rect 1536 1539 1538 1548
rect 1039 1538 1043 1539
rect 1039 1533 1043 1534
rect 1047 1538 1051 1539
rect 1047 1533 1051 1534
rect 1191 1538 1195 1539
rect 1191 1533 1195 1534
rect 1207 1538 1211 1539
rect 1207 1533 1211 1534
rect 1343 1538 1347 1539
rect 1343 1533 1347 1534
rect 1367 1538 1371 1539
rect 1367 1533 1371 1534
rect 1495 1538 1499 1539
rect 1495 1533 1499 1534
rect 1535 1538 1539 1539
rect 1535 1533 1539 1534
rect 1040 1528 1042 1533
rect 1192 1528 1194 1533
rect 1344 1528 1346 1533
rect 1496 1528 1498 1533
rect 1038 1527 1044 1528
rect 1038 1523 1039 1527
rect 1043 1523 1044 1527
rect 1038 1522 1044 1523
rect 1190 1527 1196 1528
rect 1190 1523 1191 1527
rect 1195 1523 1196 1527
rect 1190 1522 1196 1523
rect 1342 1527 1348 1528
rect 1342 1523 1343 1527
rect 1347 1523 1348 1527
rect 1342 1522 1348 1523
rect 1494 1527 1500 1528
rect 1494 1523 1495 1527
rect 1499 1523 1500 1527
rect 1494 1522 1500 1523
rect 650 1519 656 1520
rect 650 1515 651 1519
rect 655 1515 656 1519
rect 650 1514 656 1515
rect 954 1519 960 1520
rect 954 1515 955 1519
rect 959 1515 960 1519
rect 954 1514 960 1515
rect 650 1503 656 1504
rect 650 1499 651 1503
rect 655 1499 656 1503
rect 650 1498 656 1499
rect 954 1503 960 1504
rect 954 1499 955 1503
rect 959 1499 960 1503
rect 954 1498 960 1499
rect 1410 1503 1416 1504
rect 1410 1499 1411 1503
rect 1415 1499 1416 1503
rect 1410 1498 1416 1499
rect 1418 1503 1424 1504
rect 1418 1499 1419 1503
rect 1423 1499 1424 1503
rect 1418 1498 1424 1499
rect 590 1487 596 1488
rect 590 1483 591 1487
rect 595 1483 596 1487
rect 590 1482 596 1483
rect 462 1475 468 1476
rect 462 1471 463 1475
rect 467 1471 468 1475
rect 462 1470 468 1471
rect 592 1463 594 1482
rect 652 1476 654 1498
rect 742 1487 748 1488
rect 742 1483 743 1487
rect 747 1483 748 1487
rect 742 1482 748 1483
rect 894 1487 900 1488
rect 894 1483 895 1487
rect 899 1483 900 1487
rect 894 1482 900 1483
rect 650 1475 656 1476
rect 650 1471 651 1475
rect 655 1471 656 1475
rect 650 1470 656 1471
rect 744 1463 746 1482
rect 896 1463 898 1482
rect 956 1476 958 1498
rect 1046 1487 1052 1488
rect 1046 1483 1047 1487
rect 1051 1483 1052 1487
rect 1046 1482 1052 1483
rect 1198 1487 1204 1488
rect 1198 1483 1199 1487
rect 1203 1483 1204 1487
rect 1198 1482 1204 1483
rect 1350 1487 1356 1488
rect 1350 1483 1351 1487
rect 1355 1483 1356 1487
rect 1350 1482 1356 1483
rect 954 1475 960 1476
rect 954 1471 955 1475
rect 959 1471 960 1475
rect 954 1470 960 1471
rect 1048 1463 1050 1482
rect 1078 1475 1084 1476
rect 1078 1471 1079 1475
rect 1083 1471 1084 1475
rect 1078 1470 1084 1471
rect 263 1462 267 1463
rect 263 1457 267 1458
rect 279 1462 283 1463
rect 279 1457 283 1458
rect 399 1462 403 1463
rect 399 1457 403 1458
rect 431 1462 435 1463
rect 431 1457 435 1458
rect 535 1462 539 1463
rect 535 1457 539 1458
rect 591 1462 595 1463
rect 591 1457 595 1458
rect 663 1462 667 1463
rect 663 1457 667 1458
rect 743 1462 747 1463
rect 743 1457 747 1458
rect 791 1462 795 1463
rect 791 1457 795 1458
rect 895 1462 899 1463
rect 895 1457 899 1458
rect 911 1462 915 1463
rect 911 1457 915 1458
rect 1023 1462 1027 1463
rect 1023 1457 1027 1458
rect 1047 1462 1051 1463
rect 1047 1457 1051 1458
rect 198 1455 204 1456
rect 198 1451 199 1455
rect 203 1451 204 1455
rect 198 1450 204 1451
rect 264 1446 266 1457
rect 400 1446 402 1457
rect 536 1446 538 1457
rect 622 1447 628 1448
rect 142 1445 148 1446
rect 142 1441 143 1445
rect 147 1441 148 1445
rect 142 1440 148 1441
rect 262 1445 268 1446
rect 262 1441 263 1445
rect 267 1441 268 1445
rect 262 1440 268 1441
rect 398 1445 404 1446
rect 398 1441 399 1445
rect 403 1441 404 1445
rect 398 1440 404 1441
rect 534 1445 540 1446
rect 534 1441 535 1445
rect 539 1441 540 1445
rect 622 1443 623 1447
rect 627 1443 628 1447
rect 664 1446 666 1457
rect 792 1446 794 1457
rect 912 1446 914 1457
rect 1024 1446 1026 1457
rect 622 1442 628 1443
rect 662 1445 668 1446
rect 534 1440 540 1441
rect 110 1432 116 1433
rect 110 1428 111 1432
rect 115 1428 116 1432
rect 110 1427 116 1428
rect 110 1415 116 1416
rect 110 1411 111 1415
rect 115 1411 116 1415
rect 110 1410 116 1411
rect 534 1415 540 1416
rect 534 1411 535 1415
rect 539 1411 540 1415
rect 534 1410 540 1411
rect 112 1395 114 1410
rect 134 1405 140 1406
rect 134 1401 135 1405
rect 139 1401 140 1405
rect 134 1400 140 1401
rect 254 1405 260 1406
rect 254 1401 255 1405
rect 259 1401 260 1405
rect 254 1400 260 1401
rect 390 1405 396 1406
rect 390 1401 391 1405
rect 395 1401 396 1405
rect 390 1400 396 1401
rect 526 1405 532 1406
rect 526 1401 527 1405
rect 531 1401 532 1405
rect 526 1400 532 1401
rect 136 1395 138 1400
rect 256 1395 258 1400
rect 392 1395 394 1400
rect 528 1395 530 1400
rect 111 1394 115 1395
rect 111 1389 115 1390
rect 135 1394 139 1395
rect 135 1389 139 1390
rect 255 1394 259 1395
rect 255 1389 259 1390
rect 327 1394 331 1395
rect 327 1389 331 1390
rect 391 1394 395 1395
rect 391 1389 395 1390
rect 527 1394 531 1395
rect 527 1389 531 1390
rect 112 1374 114 1389
rect 136 1384 138 1389
rect 328 1384 330 1389
rect 134 1383 140 1384
rect 134 1379 135 1383
rect 139 1379 140 1383
rect 134 1378 140 1379
rect 326 1383 332 1384
rect 326 1379 327 1383
rect 331 1379 332 1383
rect 326 1378 332 1379
rect 110 1373 116 1374
rect 110 1369 111 1373
rect 115 1369 116 1373
rect 110 1368 116 1369
rect 394 1359 400 1360
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 394 1355 395 1359
rect 399 1355 400 1359
rect 394 1354 400 1355
rect 110 1351 116 1352
rect 198 1351 204 1352
rect 112 1319 114 1351
rect 198 1347 199 1351
rect 203 1347 204 1351
rect 198 1346 204 1347
rect 142 1343 148 1344
rect 142 1339 143 1343
rect 147 1339 148 1343
rect 142 1338 148 1339
rect 144 1319 146 1338
rect 111 1318 115 1319
rect 111 1313 115 1314
rect 143 1318 147 1319
rect 143 1313 147 1314
rect 112 1289 114 1313
rect 144 1302 146 1313
rect 200 1312 202 1346
rect 334 1343 340 1344
rect 334 1339 335 1343
rect 339 1339 340 1343
rect 334 1338 340 1339
rect 336 1319 338 1338
rect 396 1332 398 1354
rect 536 1332 538 1410
rect 551 1394 555 1395
rect 551 1389 555 1390
rect 552 1384 554 1389
rect 550 1383 556 1384
rect 550 1379 551 1383
rect 555 1379 556 1383
rect 550 1378 556 1379
rect 624 1376 626 1442
rect 662 1441 663 1445
rect 667 1441 668 1445
rect 662 1440 668 1441
rect 790 1445 796 1446
rect 790 1441 791 1445
rect 795 1441 796 1445
rect 790 1440 796 1441
rect 910 1445 916 1446
rect 910 1441 911 1445
rect 915 1441 916 1445
rect 910 1440 916 1441
rect 1022 1445 1028 1446
rect 1022 1441 1023 1445
rect 1027 1441 1028 1445
rect 1022 1440 1028 1441
rect 1080 1440 1082 1470
rect 1090 1463 1096 1464
rect 1200 1463 1202 1482
rect 1352 1463 1354 1482
rect 1090 1459 1091 1463
rect 1095 1459 1096 1463
rect 1090 1458 1096 1459
rect 1143 1462 1147 1463
rect 1078 1439 1084 1440
rect 1078 1435 1079 1439
rect 1083 1435 1084 1439
rect 1078 1434 1084 1435
rect 1092 1428 1094 1458
rect 1143 1457 1147 1458
rect 1199 1462 1203 1463
rect 1199 1457 1203 1458
rect 1263 1462 1267 1463
rect 1263 1457 1267 1458
rect 1351 1462 1355 1463
rect 1351 1457 1355 1458
rect 1383 1462 1387 1463
rect 1383 1457 1387 1458
rect 1144 1446 1146 1457
rect 1210 1455 1216 1456
rect 1210 1451 1211 1455
rect 1215 1451 1216 1455
rect 1210 1450 1216 1451
rect 1142 1445 1148 1446
rect 1142 1441 1143 1445
rect 1147 1441 1148 1445
rect 1142 1440 1148 1441
rect 1212 1428 1214 1450
rect 1264 1446 1266 1457
rect 1384 1446 1386 1457
rect 1412 1456 1414 1498
rect 1420 1468 1422 1498
rect 1502 1487 1508 1488
rect 1502 1483 1503 1487
rect 1507 1483 1508 1487
rect 1502 1482 1508 1483
rect 1418 1467 1424 1468
rect 1418 1463 1419 1467
rect 1423 1463 1424 1467
rect 1504 1463 1506 1482
rect 1544 1476 1546 1558
rect 1824 1539 1826 1558
rect 1864 1543 1866 1566
rect 1886 1561 1892 1562
rect 1886 1557 1887 1561
rect 1891 1557 1892 1561
rect 1886 1556 1892 1557
rect 2006 1561 2012 1562
rect 2006 1557 2007 1561
rect 2011 1557 2012 1561
rect 2006 1556 2012 1557
rect 2142 1561 2148 1562
rect 2142 1557 2143 1561
rect 2147 1557 2148 1561
rect 2142 1556 2148 1557
rect 1888 1543 1890 1556
rect 2008 1543 2010 1556
rect 2144 1543 2146 1556
rect 1863 1542 1867 1543
rect 1823 1538 1827 1539
rect 1863 1537 1867 1538
rect 1887 1542 1891 1543
rect 1887 1537 1891 1538
rect 2007 1542 2011 1543
rect 2007 1537 2011 1538
rect 2023 1542 2027 1543
rect 2023 1537 2027 1538
rect 2143 1542 2147 1543
rect 2143 1537 2147 1538
rect 2183 1542 2187 1543
rect 2183 1537 2187 1538
rect 1823 1533 1827 1534
rect 1824 1518 1826 1533
rect 1864 1522 1866 1537
rect 1888 1532 1890 1537
rect 2024 1532 2026 1537
rect 2184 1532 2186 1537
rect 1886 1531 1892 1532
rect 1886 1527 1887 1531
rect 1891 1527 1892 1531
rect 1886 1526 1892 1527
rect 2022 1531 2028 1532
rect 2022 1527 2023 1531
rect 2027 1527 2028 1531
rect 2022 1526 2028 1527
rect 2182 1531 2188 1532
rect 2182 1527 2183 1531
rect 2187 1527 2188 1531
rect 2182 1526 2188 1527
rect 1862 1521 1868 1522
rect 1822 1517 1828 1518
rect 1822 1513 1823 1517
rect 1827 1513 1828 1517
rect 1862 1517 1863 1521
rect 1867 1517 1868 1521
rect 1862 1516 1868 1517
rect 1822 1512 1828 1513
rect 1862 1504 1868 1505
rect 1822 1500 1828 1501
rect 1822 1496 1823 1500
rect 1827 1496 1828 1500
rect 1862 1500 1863 1504
rect 1867 1500 1868 1504
rect 1862 1499 1868 1500
rect 1822 1495 1828 1496
rect 1542 1475 1548 1476
rect 1542 1471 1543 1475
rect 1547 1471 1548 1475
rect 1542 1470 1548 1471
rect 1824 1463 1826 1495
rect 1864 1467 1866 1499
rect 1894 1491 1900 1492
rect 1894 1487 1895 1491
rect 1899 1487 1900 1491
rect 1894 1486 1900 1487
rect 2030 1491 2036 1492
rect 2030 1487 2031 1491
rect 2035 1487 2036 1491
rect 2030 1486 2036 1487
rect 2190 1491 2196 1492
rect 2190 1487 2191 1491
rect 2195 1487 2196 1491
rect 2190 1486 2196 1487
rect 1896 1467 1898 1486
rect 2032 1467 2034 1486
rect 2192 1467 2194 1486
rect 2224 1480 2226 1566
rect 2278 1561 2284 1562
rect 2278 1557 2279 1561
rect 2283 1557 2284 1561
rect 2278 1556 2284 1557
rect 2422 1561 2428 1562
rect 2422 1557 2423 1561
rect 2427 1557 2428 1561
rect 2422 1556 2428 1557
rect 2574 1561 2580 1562
rect 2574 1557 2575 1561
rect 2579 1557 2580 1561
rect 2574 1556 2580 1557
rect 2734 1561 2740 1562
rect 2734 1557 2735 1561
rect 2739 1557 2740 1561
rect 2734 1556 2740 1557
rect 2902 1561 2908 1562
rect 2902 1557 2903 1561
rect 2907 1557 2908 1561
rect 2902 1556 2908 1557
rect 2280 1543 2282 1556
rect 2424 1543 2426 1556
rect 2576 1543 2578 1556
rect 2736 1543 2738 1556
rect 2904 1543 2906 1556
rect 2279 1542 2283 1543
rect 2279 1537 2283 1538
rect 2343 1542 2347 1543
rect 2343 1537 2347 1538
rect 2423 1542 2427 1543
rect 2423 1537 2427 1538
rect 2503 1542 2507 1543
rect 2503 1537 2507 1538
rect 2575 1542 2579 1543
rect 2575 1537 2579 1538
rect 2663 1542 2667 1543
rect 2663 1537 2667 1538
rect 2735 1542 2739 1543
rect 2735 1537 2739 1538
rect 2823 1542 2827 1543
rect 2823 1537 2827 1538
rect 2903 1542 2907 1543
rect 2903 1537 2907 1538
rect 2983 1542 2987 1543
rect 2983 1537 2987 1538
rect 2344 1532 2346 1537
rect 2504 1532 2506 1537
rect 2664 1532 2666 1537
rect 2703 1532 2707 1533
rect 2824 1532 2826 1537
rect 2984 1532 2986 1537
rect 3020 1533 3022 1566
rect 3086 1561 3092 1562
rect 3086 1557 3087 1561
rect 3091 1557 3092 1561
rect 3086 1556 3092 1557
rect 3270 1561 3276 1562
rect 3270 1557 3271 1561
rect 3275 1557 3276 1561
rect 3270 1556 3276 1557
rect 3088 1543 3090 1556
rect 3272 1543 3274 1556
rect 3087 1542 3091 1543
rect 3087 1537 3091 1538
rect 3151 1542 3155 1543
rect 3151 1537 3155 1538
rect 3271 1542 3275 1543
rect 3271 1537 3275 1538
rect 3019 1532 3023 1533
rect 3152 1532 3154 1537
rect 2342 1531 2348 1532
rect 2342 1527 2343 1531
rect 2347 1527 2348 1531
rect 2342 1526 2348 1527
rect 2502 1531 2508 1532
rect 2502 1527 2503 1531
rect 2507 1527 2508 1531
rect 2502 1526 2508 1527
rect 2662 1531 2668 1532
rect 2662 1527 2663 1531
rect 2667 1527 2668 1531
rect 2703 1527 2707 1528
rect 2822 1531 2828 1532
rect 2822 1527 2823 1531
rect 2827 1527 2828 1531
rect 2662 1526 2668 1527
rect 2566 1499 2572 1500
rect 2566 1495 2567 1499
rect 2571 1495 2572 1499
rect 2566 1494 2572 1495
rect 2350 1491 2356 1492
rect 2350 1487 2351 1491
rect 2355 1487 2356 1491
rect 2350 1486 2356 1487
rect 2510 1491 2516 1492
rect 2510 1487 2511 1491
rect 2515 1487 2516 1491
rect 2510 1486 2516 1487
rect 2222 1479 2228 1480
rect 2222 1475 2223 1479
rect 2227 1475 2228 1479
rect 2222 1474 2228 1475
rect 2352 1467 2354 1486
rect 2512 1467 2514 1486
rect 1863 1466 1867 1467
rect 1418 1462 1424 1463
rect 1503 1462 1507 1463
rect 1503 1457 1507 1458
rect 1631 1462 1635 1463
rect 1631 1457 1635 1458
rect 1735 1462 1739 1463
rect 1735 1457 1739 1458
rect 1823 1462 1827 1463
rect 1863 1461 1867 1462
rect 1895 1466 1899 1467
rect 1895 1461 1899 1462
rect 2031 1466 2035 1467
rect 2031 1461 2035 1462
rect 2183 1466 2187 1467
rect 2183 1461 2187 1462
rect 2191 1466 2195 1467
rect 2191 1461 2195 1462
rect 2351 1466 2355 1467
rect 2351 1461 2355 1462
rect 2359 1466 2363 1467
rect 2359 1461 2363 1462
rect 2511 1466 2515 1467
rect 2511 1461 2515 1462
rect 2527 1466 2531 1467
rect 2527 1461 2531 1462
rect 1823 1457 1827 1458
rect 1402 1455 1408 1456
rect 1402 1451 1403 1455
rect 1407 1451 1408 1455
rect 1402 1450 1408 1451
rect 1410 1455 1416 1456
rect 1410 1451 1411 1455
rect 1415 1451 1416 1455
rect 1410 1450 1416 1451
rect 1262 1445 1268 1446
rect 1262 1441 1263 1445
rect 1267 1441 1268 1445
rect 1262 1440 1268 1441
rect 1382 1445 1388 1446
rect 1382 1441 1383 1445
rect 1387 1441 1388 1445
rect 1382 1440 1388 1441
rect 1090 1427 1096 1428
rect 1090 1423 1091 1427
rect 1095 1423 1096 1427
rect 1090 1422 1096 1423
rect 1210 1427 1216 1428
rect 1210 1423 1211 1427
rect 1215 1423 1216 1427
rect 1210 1422 1216 1423
rect 654 1405 660 1406
rect 654 1401 655 1405
rect 659 1401 660 1405
rect 654 1400 660 1401
rect 782 1405 788 1406
rect 782 1401 783 1405
rect 787 1401 788 1405
rect 782 1400 788 1401
rect 902 1405 908 1406
rect 902 1401 903 1405
rect 907 1401 908 1405
rect 902 1400 908 1401
rect 1014 1405 1020 1406
rect 1014 1401 1015 1405
rect 1019 1401 1020 1405
rect 1014 1400 1020 1401
rect 1134 1405 1140 1406
rect 1134 1401 1135 1405
rect 1139 1401 1140 1405
rect 1134 1400 1140 1401
rect 1254 1405 1260 1406
rect 1254 1401 1255 1405
rect 1259 1401 1260 1405
rect 1254 1400 1260 1401
rect 1374 1405 1380 1406
rect 1374 1401 1375 1405
rect 1379 1401 1380 1405
rect 1374 1400 1380 1401
rect 1404 1400 1406 1450
rect 1504 1446 1506 1457
rect 1632 1446 1634 1457
rect 1736 1446 1738 1457
rect 1502 1445 1508 1446
rect 1502 1441 1503 1445
rect 1507 1441 1508 1445
rect 1502 1440 1508 1441
rect 1630 1445 1636 1446
rect 1630 1441 1631 1445
rect 1635 1441 1636 1445
rect 1630 1440 1636 1441
rect 1734 1445 1740 1446
rect 1734 1441 1735 1445
rect 1739 1441 1740 1445
rect 1734 1440 1740 1441
rect 1824 1433 1826 1457
rect 1864 1437 1866 1461
rect 2184 1450 2186 1461
rect 2222 1459 2228 1460
rect 2222 1455 2223 1459
rect 2227 1455 2228 1459
rect 2222 1454 2228 1455
rect 2182 1449 2188 1450
rect 2182 1445 2183 1449
rect 2187 1445 2188 1449
rect 2182 1444 2188 1445
rect 2224 1437 2226 1454
rect 2360 1450 2362 1461
rect 2528 1450 2530 1461
rect 2568 1460 2570 1494
rect 2670 1491 2676 1492
rect 2670 1487 2671 1491
rect 2675 1487 2676 1491
rect 2670 1486 2676 1487
rect 2672 1467 2674 1486
rect 2704 1480 2706 1527
rect 2822 1526 2828 1527
rect 2982 1531 2988 1532
rect 2982 1527 2983 1531
rect 2987 1527 2988 1531
rect 3019 1527 3023 1528
rect 3150 1531 3156 1532
rect 3150 1527 3151 1531
rect 3155 1527 3156 1531
rect 2982 1526 2988 1527
rect 3150 1526 3156 1527
rect 3312 1524 3314 1606
rect 3472 1602 3474 1613
rect 3500 1612 3502 1654
rect 3574 1652 3575 1656
rect 3579 1652 3580 1656
rect 3574 1651 3580 1652
rect 3576 1619 3578 1651
rect 3575 1618 3579 1619
rect 3575 1613 3579 1614
rect 3498 1611 3504 1612
rect 3498 1607 3499 1611
rect 3503 1607 3504 1611
rect 3498 1606 3504 1607
rect 3470 1601 3476 1602
rect 3470 1597 3471 1601
rect 3475 1597 3476 1601
rect 3470 1596 3476 1597
rect 3576 1589 3578 1613
rect 3574 1588 3580 1589
rect 3574 1584 3575 1588
rect 3579 1584 3580 1588
rect 3574 1583 3580 1584
rect 3574 1571 3580 1572
rect 3574 1567 3575 1571
rect 3579 1567 3580 1571
rect 3574 1566 3580 1567
rect 3462 1561 3468 1562
rect 3462 1557 3463 1561
rect 3467 1557 3468 1561
rect 3462 1556 3468 1557
rect 3464 1543 3466 1556
rect 3514 1555 3520 1556
rect 3514 1551 3515 1555
rect 3519 1551 3520 1555
rect 3514 1550 3520 1551
rect 3319 1542 3323 1543
rect 3319 1537 3323 1538
rect 3463 1542 3467 1543
rect 3463 1537 3467 1538
rect 3479 1542 3483 1543
rect 3479 1537 3483 1538
rect 3320 1532 3322 1537
rect 3480 1532 3482 1537
rect 3318 1531 3324 1532
rect 3318 1527 3319 1531
rect 3323 1527 3324 1531
rect 3318 1526 3324 1527
rect 3478 1531 3484 1532
rect 3478 1527 3479 1531
rect 3483 1527 3484 1531
rect 3478 1526 3484 1527
rect 3078 1523 3084 1524
rect 3078 1519 3079 1523
rect 3083 1519 3084 1523
rect 3078 1518 3084 1519
rect 3310 1523 3316 1524
rect 3310 1519 3311 1523
rect 3315 1519 3316 1523
rect 3310 1518 3316 1519
rect 2730 1507 2736 1508
rect 2730 1503 2731 1507
rect 2735 1503 2736 1507
rect 2730 1502 2736 1503
rect 2719 1484 2723 1485
rect 2732 1480 2734 1502
rect 2830 1491 2836 1492
rect 2830 1487 2831 1491
rect 2835 1487 2836 1491
rect 2830 1486 2836 1487
rect 2990 1491 2996 1492
rect 2990 1487 2991 1491
rect 2995 1487 2996 1491
rect 2990 1486 2996 1487
rect 2702 1479 2708 1480
rect 2719 1479 2723 1480
rect 2730 1479 2736 1480
rect 2702 1475 2703 1479
rect 2707 1475 2708 1479
rect 2702 1474 2708 1475
rect 2671 1466 2675 1467
rect 2671 1461 2675 1462
rect 2687 1466 2691 1467
rect 2687 1461 2691 1462
rect 2566 1459 2572 1460
rect 2566 1455 2567 1459
rect 2571 1455 2572 1459
rect 2566 1454 2572 1455
rect 2688 1450 2690 1461
rect 2720 1460 2722 1479
rect 2730 1475 2731 1479
rect 2735 1475 2736 1479
rect 2730 1474 2736 1475
rect 2832 1467 2834 1486
rect 2992 1467 2994 1486
rect 3080 1485 3082 1518
rect 3158 1491 3164 1492
rect 3158 1487 3159 1491
rect 3163 1487 3164 1491
rect 3158 1486 3164 1487
rect 3326 1491 3332 1492
rect 3326 1487 3327 1491
rect 3331 1487 3332 1491
rect 3326 1486 3332 1487
rect 3486 1491 3492 1492
rect 3486 1487 3487 1491
rect 3491 1487 3492 1491
rect 3486 1486 3492 1487
rect 3079 1484 3083 1485
rect 3079 1479 3083 1480
rect 3160 1467 3162 1486
rect 3328 1467 3330 1486
rect 3350 1479 3356 1480
rect 3350 1475 3351 1479
rect 3355 1475 3356 1479
rect 3350 1474 3356 1475
rect 2831 1466 2835 1467
rect 2831 1461 2835 1462
rect 2847 1466 2851 1467
rect 2847 1461 2851 1462
rect 2991 1466 2995 1467
rect 2991 1461 2995 1462
rect 3007 1466 3011 1467
rect 3007 1461 3011 1462
rect 3159 1466 3163 1467
rect 3159 1461 3163 1462
rect 3175 1466 3179 1467
rect 3175 1461 3179 1462
rect 3327 1466 3331 1467
rect 3327 1461 3331 1462
rect 3343 1466 3347 1467
rect 3343 1461 3347 1462
rect 2718 1459 2724 1460
rect 2718 1455 2719 1459
rect 2723 1455 2724 1459
rect 2718 1454 2724 1455
rect 2848 1450 2850 1461
rect 3008 1450 3010 1461
rect 3176 1450 3178 1461
rect 3344 1450 3346 1461
rect 2358 1449 2364 1450
rect 2358 1445 2359 1449
rect 2363 1445 2364 1449
rect 2358 1444 2364 1445
rect 2526 1449 2532 1450
rect 2526 1445 2527 1449
rect 2531 1445 2532 1449
rect 2526 1444 2532 1445
rect 2686 1449 2692 1450
rect 2686 1445 2687 1449
rect 2691 1445 2692 1449
rect 2686 1444 2692 1445
rect 2846 1449 2852 1450
rect 2846 1445 2847 1449
rect 2851 1445 2852 1449
rect 2846 1444 2852 1445
rect 3006 1449 3012 1450
rect 3006 1445 3007 1449
rect 3011 1445 3012 1449
rect 3006 1444 3012 1445
rect 3174 1449 3180 1450
rect 3174 1445 3175 1449
rect 3179 1445 3180 1449
rect 3174 1444 3180 1445
rect 3342 1449 3348 1450
rect 3342 1445 3343 1449
rect 3347 1445 3348 1449
rect 3342 1444 3348 1445
rect 1862 1436 1868 1437
rect 1822 1432 1828 1433
rect 1822 1428 1823 1432
rect 1827 1428 1828 1432
rect 1862 1432 1863 1436
rect 1867 1432 1868 1436
rect 1862 1431 1868 1432
rect 2223 1436 2227 1437
rect 2427 1436 2431 1437
rect 2223 1431 2227 1432
rect 2426 1431 2432 1432
rect 1822 1427 1828 1428
rect 2426 1427 2427 1431
rect 2431 1427 2432 1431
rect 2426 1426 2432 1427
rect 1862 1419 1868 1420
rect 1822 1415 1828 1416
rect 1822 1411 1823 1415
rect 1827 1411 1828 1415
rect 1862 1415 1863 1419
rect 1867 1415 1868 1419
rect 1862 1414 1868 1415
rect 2474 1419 2480 1420
rect 2474 1415 2475 1419
rect 2479 1415 2480 1419
rect 2474 1414 2480 1415
rect 3258 1419 3264 1420
rect 3258 1415 3259 1419
rect 3263 1415 3264 1419
rect 3258 1414 3264 1415
rect 1822 1410 1828 1411
rect 1494 1405 1500 1406
rect 1494 1401 1495 1405
rect 1499 1401 1500 1405
rect 1494 1400 1500 1401
rect 1622 1405 1628 1406
rect 1622 1401 1623 1405
rect 1627 1401 1628 1405
rect 1622 1400 1628 1401
rect 1726 1405 1732 1406
rect 1726 1401 1727 1405
rect 1731 1401 1732 1405
rect 1726 1400 1732 1401
rect 656 1395 658 1400
rect 784 1395 786 1400
rect 904 1395 906 1400
rect 1016 1395 1018 1400
rect 1136 1395 1138 1400
rect 1256 1395 1258 1400
rect 1376 1395 1378 1400
rect 1402 1399 1408 1400
rect 1402 1395 1403 1399
rect 1407 1395 1408 1399
rect 1496 1395 1498 1400
rect 1624 1395 1626 1400
rect 1728 1395 1730 1400
rect 1824 1395 1826 1410
rect 655 1394 659 1395
rect 655 1389 659 1390
rect 783 1394 787 1395
rect 783 1389 787 1390
rect 903 1394 907 1395
rect 903 1389 907 1390
rect 1015 1394 1019 1395
rect 1015 1389 1019 1390
rect 1023 1394 1027 1395
rect 1023 1389 1027 1390
rect 1135 1394 1139 1395
rect 1135 1389 1139 1390
rect 1255 1394 1259 1395
rect 1255 1389 1259 1390
rect 1263 1394 1267 1395
rect 1263 1389 1267 1390
rect 1375 1394 1379 1395
rect 1402 1394 1408 1395
rect 1495 1394 1499 1395
rect 1375 1389 1379 1390
rect 1495 1389 1499 1390
rect 1503 1394 1507 1395
rect 1503 1389 1507 1390
rect 1623 1394 1627 1395
rect 1623 1389 1627 1390
rect 1727 1394 1731 1395
rect 1727 1389 1731 1390
rect 1823 1394 1827 1395
rect 1864 1391 1866 1414
rect 2174 1409 2180 1410
rect 2174 1405 2175 1409
rect 2179 1405 2180 1409
rect 2174 1404 2180 1405
rect 2350 1409 2356 1410
rect 2350 1405 2351 1409
rect 2355 1405 2356 1409
rect 2350 1404 2356 1405
rect 2176 1391 2178 1404
rect 2352 1391 2354 1404
rect 1823 1389 1827 1390
rect 1863 1390 1867 1391
rect 784 1384 786 1389
rect 1024 1384 1026 1389
rect 1264 1384 1266 1389
rect 1504 1384 1506 1389
rect 1728 1384 1730 1389
rect 782 1383 788 1384
rect 782 1379 783 1383
rect 787 1379 788 1383
rect 782 1378 788 1379
rect 1022 1383 1028 1384
rect 1022 1379 1023 1383
rect 1027 1379 1028 1383
rect 1022 1378 1028 1379
rect 1262 1383 1268 1384
rect 1262 1379 1263 1383
rect 1267 1379 1268 1383
rect 1262 1378 1268 1379
rect 1502 1383 1508 1384
rect 1502 1379 1503 1383
rect 1507 1379 1508 1383
rect 1502 1378 1508 1379
rect 1726 1383 1732 1384
rect 1726 1379 1727 1383
rect 1731 1379 1732 1383
rect 1726 1378 1732 1379
rect 622 1375 628 1376
rect 622 1371 623 1375
rect 627 1371 628 1375
rect 1824 1374 1826 1389
rect 1863 1385 1867 1386
rect 2079 1390 2083 1391
rect 2079 1385 2083 1386
rect 2175 1390 2179 1391
rect 2175 1385 2179 1386
rect 2263 1390 2267 1391
rect 2263 1385 2267 1386
rect 2351 1390 2355 1391
rect 2351 1385 2355 1386
rect 2439 1390 2443 1391
rect 2439 1385 2443 1386
rect 622 1370 628 1371
rect 1822 1373 1828 1374
rect 1822 1369 1823 1373
rect 1827 1369 1828 1373
rect 1864 1370 1866 1385
rect 2080 1380 2082 1385
rect 2264 1380 2266 1385
rect 2440 1380 2442 1385
rect 2078 1379 2084 1380
rect 2078 1375 2079 1379
rect 2083 1375 2084 1379
rect 2078 1374 2084 1375
rect 2262 1379 2268 1380
rect 2262 1375 2263 1379
rect 2267 1375 2268 1379
rect 2262 1374 2268 1375
rect 2438 1379 2444 1380
rect 2438 1375 2439 1379
rect 2443 1375 2444 1379
rect 2438 1374 2444 1375
rect 1822 1368 1828 1369
rect 1862 1369 1868 1370
rect 1862 1365 1863 1369
rect 1867 1365 1868 1369
rect 1862 1364 1868 1365
rect 850 1359 856 1360
rect 850 1355 851 1359
rect 855 1355 856 1359
rect 850 1354 856 1355
rect 1638 1359 1644 1360
rect 1638 1355 1639 1359
rect 1643 1355 1644 1359
rect 1638 1354 1644 1355
rect 1822 1356 1828 1357
rect 558 1343 564 1344
rect 558 1339 559 1343
rect 563 1339 564 1343
rect 558 1338 564 1339
rect 790 1343 796 1344
rect 790 1339 791 1343
rect 795 1339 796 1343
rect 790 1338 796 1339
rect 394 1331 400 1332
rect 394 1327 395 1331
rect 399 1327 400 1331
rect 394 1326 400 1327
rect 534 1331 540 1332
rect 534 1327 535 1331
rect 539 1327 540 1331
rect 534 1326 540 1327
rect 560 1319 562 1338
rect 792 1319 794 1338
rect 852 1332 854 1354
rect 1030 1343 1036 1344
rect 1030 1339 1031 1343
rect 1035 1339 1036 1343
rect 1030 1338 1036 1339
rect 1270 1343 1276 1344
rect 1270 1339 1271 1343
rect 1275 1339 1276 1343
rect 1510 1343 1516 1344
rect 1270 1338 1276 1339
rect 1303 1340 1307 1341
rect 850 1331 856 1332
rect 850 1327 851 1331
rect 855 1327 856 1331
rect 850 1326 856 1327
rect 1032 1319 1034 1338
rect 1272 1319 1274 1338
rect 1510 1339 1511 1343
rect 1515 1339 1516 1343
rect 1640 1341 1642 1354
rect 1822 1352 1823 1356
rect 1827 1352 1828 1356
rect 2338 1355 2344 1356
rect 1822 1351 1828 1352
rect 1862 1352 1868 1353
rect 1734 1343 1740 1344
rect 1510 1338 1516 1339
rect 1639 1340 1643 1341
rect 1303 1335 1307 1336
rect 1304 1332 1306 1335
rect 1302 1331 1308 1332
rect 1302 1327 1303 1331
rect 1307 1327 1308 1331
rect 1302 1326 1308 1327
rect 1458 1319 1464 1320
rect 1512 1319 1514 1338
rect 1734 1339 1735 1343
rect 1739 1339 1740 1343
rect 1734 1338 1740 1339
rect 1639 1335 1643 1336
rect 1736 1319 1738 1338
rect 1824 1319 1826 1351
rect 1862 1348 1863 1352
rect 1867 1348 1868 1352
rect 2338 1351 2339 1355
rect 2343 1351 2344 1355
rect 2338 1350 2344 1351
rect 1862 1347 1868 1348
rect 1864 1323 1866 1347
rect 2086 1339 2092 1340
rect 2086 1335 2087 1339
rect 2091 1335 2092 1339
rect 2086 1334 2092 1335
rect 2270 1339 2276 1340
rect 2270 1335 2271 1339
rect 2275 1335 2276 1339
rect 2270 1334 2276 1335
rect 2088 1323 2090 1334
rect 2119 1332 2123 1333
rect 2118 1327 2124 1328
rect 2118 1323 2119 1327
rect 2123 1323 2124 1327
rect 2272 1323 2274 1334
rect 1863 1322 1867 1323
rect 327 1318 331 1319
rect 327 1313 331 1314
rect 335 1318 339 1319
rect 335 1313 339 1314
rect 527 1318 531 1319
rect 527 1313 531 1314
rect 559 1318 563 1319
rect 559 1313 563 1314
rect 719 1318 723 1319
rect 719 1313 723 1314
rect 791 1318 795 1319
rect 791 1313 795 1314
rect 903 1318 907 1319
rect 903 1313 907 1314
rect 1031 1318 1035 1319
rect 1031 1313 1035 1314
rect 1071 1318 1075 1319
rect 1071 1313 1075 1314
rect 1231 1318 1235 1319
rect 1231 1313 1235 1314
rect 1271 1318 1275 1319
rect 1271 1313 1275 1314
rect 1383 1318 1387 1319
rect 1458 1315 1459 1319
rect 1463 1315 1464 1319
rect 1458 1314 1464 1315
rect 1511 1318 1515 1319
rect 1383 1313 1387 1314
rect 198 1311 204 1312
rect 198 1307 199 1311
rect 203 1307 204 1311
rect 198 1306 204 1307
rect 328 1302 330 1313
rect 528 1302 530 1313
rect 614 1311 620 1312
rect 614 1307 615 1311
rect 619 1307 620 1311
rect 614 1306 620 1307
rect 142 1301 148 1302
rect 142 1297 143 1301
rect 147 1297 148 1301
rect 142 1296 148 1297
rect 326 1301 332 1302
rect 326 1297 327 1301
rect 331 1297 332 1301
rect 326 1296 332 1297
rect 526 1301 532 1302
rect 526 1297 527 1301
rect 531 1297 532 1301
rect 526 1296 532 1297
rect 110 1288 116 1289
rect 110 1284 111 1288
rect 115 1284 116 1288
rect 110 1283 116 1284
rect 110 1271 116 1272
rect 110 1267 111 1271
rect 115 1267 116 1271
rect 110 1266 116 1267
rect 210 1271 216 1272
rect 210 1267 211 1271
rect 215 1267 216 1271
rect 210 1266 216 1267
rect 112 1247 114 1266
rect 134 1261 140 1262
rect 134 1257 135 1261
rect 139 1257 140 1261
rect 134 1256 140 1257
rect 136 1247 138 1256
rect 111 1246 115 1247
rect 111 1241 115 1242
rect 135 1246 139 1247
rect 135 1241 139 1242
rect 112 1226 114 1241
rect 136 1236 138 1241
rect 134 1235 140 1236
rect 134 1231 135 1235
rect 139 1231 140 1235
rect 134 1230 140 1231
rect 110 1225 116 1226
rect 110 1221 111 1225
rect 115 1221 116 1225
rect 110 1220 116 1221
rect 110 1208 116 1209
rect 110 1204 111 1208
rect 115 1204 116 1208
rect 110 1203 116 1204
rect 112 1175 114 1203
rect 142 1195 148 1196
rect 142 1191 143 1195
rect 147 1191 148 1195
rect 142 1190 148 1191
rect 144 1175 146 1190
rect 212 1184 214 1266
rect 318 1261 324 1262
rect 318 1257 319 1261
rect 323 1257 324 1261
rect 318 1256 324 1257
rect 518 1261 524 1262
rect 518 1257 519 1261
rect 523 1257 524 1261
rect 518 1256 524 1257
rect 320 1247 322 1256
rect 520 1247 522 1256
rect 295 1246 299 1247
rect 295 1241 299 1242
rect 319 1246 323 1247
rect 319 1241 323 1242
rect 479 1246 483 1247
rect 479 1241 483 1242
rect 519 1246 523 1247
rect 519 1241 523 1242
rect 296 1236 298 1241
rect 480 1236 482 1241
rect 294 1235 300 1236
rect 294 1231 295 1235
rect 299 1231 300 1235
rect 294 1230 300 1231
rect 478 1235 484 1236
rect 478 1231 479 1235
rect 483 1231 484 1235
rect 478 1230 484 1231
rect 616 1228 618 1306
rect 720 1302 722 1313
rect 904 1302 906 1313
rect 1072 1302 1074 1313
rect 1214 1311 1220 1312
rect 1214 1307 1215 1311
rect 1219 1307 1220 1311
rect 1214 1306 1220 1307
rect 718 1301 724 1302
rect 718 1297 719 1301
rect 723 1297 724 1301
rect 718 1296 724 1297
rect 902 1301 908 1302
rect 902 1297 903 1301
rect 907 1297 908 1301
rect 902 1296 908 1297
rect 1070 1301 1076 1302
rect 1070 1297 1071 1301
rect 1075 1297 1076 1301
rect 1070 1296 1076 1297
rect 1216 1288 1218 1306
rect 1232 1302 1234 1313
rect 1384 1302 1386 1313
rect 1230 1301 1236 1302
rect 1230 1297 1231 1301
rect 1235 1297 1236 1301
rect 1230 1296 1236 1297
rect 1382 1301 1388 1302
rect 1382 1297 1383 1301
rect 1387 1297 1388 1301
rect 1382 1296 1388 1297
rect 1214 1287 1220 1288
rect 1214 1283 1215 1287
rect 1219 1283 1220 1287
rect 1214 1282 1220 1283
rect 710 1261 716 1262
rect 710 1257 711 1261
rect 715 1257 716 1261
rect 710 1256 716 1257
rect 894 1261 900 1262
rect 894 1257 895 1261
rect 899 1257 900 1261
rect 894 1256 900 1257
rect 1062 1261 1068 1262
rect 1062 1257 1063 1261
rect 1067 1257 1068 1261
rect 1062 1256 1068 1257
rect 1222 1261 1228 1262
rect 1222 1257 1223 1261
rect 1227 1257 1228 1261
rect 1222 1256 1228 1257
rect 1374 1261 1380 1262
rect 1374 1257 1375 1261
rect 1379 1257 1380 1261
rect 1374 1256 1380 1257
rect 712 1247 714 1256
rect 896 1247 898 1256
rect 1064 1247 1066 1256
rect 1224 1247 1226 1256
rect 1376 1247 1378 1256
rect 655 1246 659 1247
rect 655 1241 659 1242
rect 711 1246 715 1247
rect 711 1241 715 1242
rect 815 1246 819 1247
rect 815 1241 819 1242
rect 895 1246 899 1247
rect 895 1241 899 1242
rect 967 1246 971 1247
rect 967 1241 971 1242
rect 1063 1246 1067 1247
rect 1063 1241 1067 1242
rect 1111 1246 1115 1247
rect 1111 1241 1115 1242
rect 1223 1246 1227 1247
rect 1223 1241 1227 1242
rect 1247 1246 1251 1247
rect 1247 1241 1251 1242
rect 1375 1246 1379 1247
rect 1375 1241 1379 1242
rect 1383 1246 1387 1247
rect 1383 1241 1387 1242
rect 656 1236 658 1241
rect 816 1236 818 1241
rect 968 1236 970 1241
rect 1112 1236 1114 1241
rect 1248 1236 1250 1241
rect 1384 1236 1386 1241
rect 654 1235 660 1236
rect 654 1231 655 1235
rect 659 1231 660 1235
rect 654 1230 660 1231
rect 814 1235 820 1236
rect 814 1231 815 1235
rect 819 1231 820 1235
rect 814 1230 820 1231
rect 966 1235 972 1236
rect 966 1231 967 1235
rect 971 1231 972 1235
rect 966 1230 972 1231
rect 1110 1235 1116 1236
rect 1110 1231 1111 1235
rect 1115 1231 1116 1235
rect 1110 1230 1116 1231
rect 1246 1235 1252 1236
rect 1246 1231 1247 1235
rect 1251 1231 1252 1235
rect 1246 1230 1252 1231
rect 1382 1235 1388 1236
rect 1382 1231 1383 1235
rect 1387 1231 1388 1235
rect 1382 1230 1388 1231
rect 1460 1228 1462 1314
rect 1511 1313 1515 1314
rect 1535 1318 1539 1319
rect 1535 1313 1539 1314
rect 1687 1318 1691 1319
rect 1687 1313 1691 1314
rect 1735 1318 1739 1319
rect 1735 1313 1739 1314
rect 1823 1318 1827 1319
rect 1863 1317 1867 1318
rect 2087 1322 2091 1323
rect 2118 1322 2124 1323
rect 2271 1322 2275 1323
rect 2087 1317 2091 1318
rect 2271 1317 2275 1318
rect 2311 1322 2315 1323
rect 2311 1317 2315 1318
rect 1823 1313 1827 1314
rect 1536 1302 1538 1313
rect 1688 1302 1690 1313
rect 1534 1301 1540 1302
rect 1534 1297 1535 1301
rect 1539 1297 1540 1301
rect 1534 1296 1540 1297
rect 1686 1301 1692 1302
rect 1686 1297 1687 1301
rect 1691 1297 1692 1301
rect 1686 1296 1692 1297
rect 1824 1289 1826 1313
rect 1864 1293 1866 1317
rect 2088 1306 2090 1317
rect 2294 1315 2300 1316
rect 2294 1311 2295 1315
rect 2299 1311 2300 1315
rect 2294 1310 2300 1311
rect 2086 1305 2092 1306
rect 2086 1301 2087 1305
rect 2091 1301 2092 1305
rect 2086 1300 2092 1301
rect 2296 1293 2298 1310
rect 2312 1306 2314 1317
rect 2340 1316 2342 1350
rect 2446 1339 2452 1340
rect 2446 1335 2447 1339
rect 2451 1335 2452 1339
rect 2446 1334 2452 1335
rect 2448 1323 2450 1334
rect 2476 1328 2478 1414
rect 2518 1409 2524 1410
rect 2518 1405 2519 1409
rect 2523 1405 2524 1409
rect 2518 1404 2524 1405
rect 2678 1409 2684 1410
rect 2678 1405 2679 1409
rect 2683 1405 2684 1409
rect 2678 1404 2684 1405
rect 2838 1409 2844 1410
rect 2838 1405 2839 1409
rect 2843 1405 2844 1409
rect 2838 1404 2844 1405
rect 2998 1409 3004 1410
rect 2998 1405 2999 1409
rect 3003 1405 3004 1409
rect 2998 1404 3004 1405
rect 3166 1409 3172 1410
rect 3166 1405 3167 1409
rect 3171 1405 3172 1409
rect 3166 1404 3172 1405
rect 2520 1391 2522 1404
rect 2680 1391 2682 1404
rect 2840 1391 2842 1404
rect 3000 1391 3002 1404
rect 3168 1391 3170 1404
rect 2519 1390 2523 1391
rect 2519 1385 2523 1386
rect 2615 1390 2619 1391
rect 2615 1385 2619 1386
rect 2679 1390 2683 1391
rect 2679 1385 2683 1386
rect 2783 1390 2787 1391
rect 2783 1385 2787 1386
rect 2839 1390 2843 1391
rect 2839 1385 2843 1386
rect 2935 1390 2939 1391
rect 2935 1385 2939 1386
rect 2999 1390 3003 1391
rect 2999 1385 3003 1386
rect 3079 1390 3083 1391
rect 3079 1385 3083 1386
rect 3167 1390 3171 1391
rect 3167 1385 3171 1386
rect 3223 1390 3227 1391
rect 3223 1385 3227 1386
rect 2616 1380 2618 1385
rect 2784 1380 2786 1385
rect 2936 1380 2938 1385
rect 3080 1380 3082 1385
rect 3224 1380 3226 1385
rect 2614 1379 2620 1380
rect 2614 1375 2615 1379
rect 2619 1375 2620 1379
rect 2614 1374 2620 1375
rect 2782 1379 2788 1380
rect 2782 1375 2783 1379
rect 2787 1375 2788 1379
rect 2782 1374 2788 1375
rect 2934 1379 2940 1380
rect 2934 1375 2935 1379
rect 2939 1375 2940 1379
rect 2934 1374 2940 1375
rect 3078 1379 3084 1380
rect 3078 1375 3079 1379
rect 3083 1375 3084 1379
rect 3078 1374 3084 1375
rect 3222 1379 3228 1380
rect 3222 1375 3223 1379
rect 3227 1375 3228 1379
rect 3222 1374 3228 1375
rect 2538 1371 2544 1372
rect 2538 1367 2539 1371
rect 2543 1367 2544 1371
rect 2538 1366 2544 1367
rect 2540 1333 2542 1366
rect 3260 1341 3262 1414
rect 3334 1409 3340 1410
rect 3334 1405 3335 1409
rect 3339 1405 3340 1409
rect 3334 1404 3340 1405
rect 3336 1391 3338 1404
rect 3335 1390 3339 1391
rect 3335 1385 3339 1386
rect 3352 1372 3354 1474
rect 3488 1467 3490 1486
rect 3516 1480 3518 1550
rect 3576 1543 3578 1566
rect 3575 1542 3579 1543
rect 3575 1537 3579 1538
rect 3576 1522 3578 1537
rect 3574 1521 3580 1522
rect 3574 1517 3575 1521
rect 3579 1517 3580 1521
rect 3574 1516 3580 1517
rect 3546 1507 3552 1508
rect 3546 1503 3547 1507
rect 3551 1503 3552 1507
rect 3546 1502 3552 1503
rect 3574 1504 3580 1505
rect 3514 1479 3520 1480
rect 3514 1475 3515 1479
rect 3519 1475 3520 1479
rect 3514 1474 3520 1475
rect 3487 1466 3491 1467
rect 3487 1461 3491 1462
rect 3488 1450 3490 1461
rect 3548 1460 3550 1502
rect 3574 1500 3575 1504
rect 3579 1500 3580 1504
rect 3574 1499 3580 1500
rect 3576 1467 3578 1499
rect 3575 1466 3579 1467
rect 3575 1461 3579 1462
rect 3546 1459 3552 1460
rect 3546 1455 3547 1459
rect 3551 1455 3552 1459
rect 3546 1454 3552 1455
rect 3486 1449 3492 1450
rect 3486 1445 3487 1449
rect 3491 1445 3492 1449
rect 3486 1444 3492 1445
rect 3576 1437 3578 1461
rect 3574 1436 3580 1437
rect 3574 1432 3575 1436
rect 3579 1432 3580 1436
rect 3574 1431 3580 1432
rect 3574 1419 3580 1420
rect 3574 1415 3575 1419
rect 3579 1415 3580 1419
rect 3574 1414 3580 1415
rect 3478 1409 3484 1410
rect 3478 1405 3479 1409
rect 3483 1405 3484 1409
rect 3478 1404 3484 1405
rect 3480 1391 3482 1404
rect 3518 1403 3524 1404
rect 3518 1399 3519 1403
rect 3523 1399 3524 1403
rect 3518 1398 3524 1399
rect 3359 1390 3363 1391
rect 3359 1385 3363 1386
rect 3479 1390 3483 1391
rect 3479 1385 3483 1386
rect 3360 1380 3362 1385
rect 3480 1380 3482 1385
rect 3358 1379 3364 1380
rect 3358 1375 3359 1379
rect 3363 1375 3364 1379
rect 3358 1374 3364 1375
rect 3478 1379 3484 1380
rect 3478 1375 3479 1379
rect 3483 1375 3484 1379
rect 3478 1374 3484 1375
rect 3350 1371 3356 1372
rect 3350 1367 3351 1371
rect 3355 1367 3356 1371
rect 3350 1366 3356 1367
rect 2823 1340 2827 1341
rect 3259 1340 3263 1341
rect 2622 1339 2628 1340
rect 2622 1335 2623 1339
rect 2627 1335 2628 1339
rect 2622 1334 2628 1335
rect 2790 1339 2796 1340
rect 2790 1335 2791 1339
rect 2795 1335 2796 1339
rect 2823 1335 2827 1336
rect 2942 1339 2948 1340
rect 2942 1335 2943 1339
rect 2947 1335 2948 1339
rect 2790 1334 2796 1335
rect 2539 1332 2543 1333
rect 2474 1327 2480 1328
rect 2539 1327 2543 1328
rect 2474 1323 2475 1327
rect 2479 1323 2480 1327
rect 2624 1323 2626 1334
rect 2792 1323 2794 1334
rect 2824 1328 2826 1335
rect 2942 1334 2948 1335
rect 3086 1339 3092 1340
rect 3086 1335 3087 1339
rect 3091 1335 3092 1339
rect 3086 1334 3092 1335
rect 3230 1339 3236 1340
rect 3230 1335 3231 1339
rect 3235 1335 3236 1339
rect 3259 1335 3263 1336
rect 3366 1339 3372 1340
rect 3366 1335 3367 1339
rect 3371 1335 3372 1339
rect 3230 1334 3236 1335
rect 3366 1334 3372 1335
rect 3486 1339 3492 1340
rect 3486 1335 3487 1339
rect 3491 1335 3492 1339
rect 3486 1334 3492 1335
rect 2822 1327 2828 1328
rect 2822 1323 2823 1327
rect 2827 1323 2828 1327
rect 2944 1323 2946 1334
rect 3088 1323 3090 1334
rect 3232 1323 3234 1334
rect 3368 1323 3370 1334
rect 3418 1327 3424 1328
rect 3418 1323 3419 1327
rect 3423 1323 3424 1327
rect 3488 1323 3490 1334
rect 3520 1328 3522 1398
rect 3576 1391 3578 1414
rect 3575 1390 3579 1391
rect 3575 1385 3579 1386
rect 3576 1370 3578 1385
rect 3574 1369 3580 1370
rect 3574 1365 3575 1369
rect 3579 1365 3580 1369
rect 3574 1364 3580 1365
rect 3546 1355 3552 1356
rect 3546 1351 3547 1355
rect 3551 1351 3552 1355
rect 3546 1350 3552 1351
rect 3574 1352 3580 1353
rect 3518 1327 3524 1328
rect 3518 1323 3519 1327
rect 3523 1323 3524 1327
rect 2447 1322 2451 1323
rect 2474 1322 2480 1323
rect 2519 1322 2523 1323
rect 2447 1317 2451 1318
rect 2519 1317 2523 1318
rect 2623 1322 2627 1323
rect 2623 1317 2627 1318
rect 2711 1322 2715 1323
rect 2711 1317 2715 1318
rect 2791 1322 2795 1323
rect 2822 1322 2828 1323
rect 2887 1322 2891 1323
rect 2791 1317 2795 1318
rect 2887 1317 2891 1318
rect 2943 1322 2947 1323
rect 2943 1317 2947 1318
rect 3047 1322 3051 1323
rect 3047 1317 3051 1318
rect 3087 1322 3091 1323
rect 3087 1317 3091 1318
rect 3199 1322 3203 1323
rect 3199 1317 3203 1318
rect 3231 1322 3235 1323
rect 3231 1317 3235 1318
rect 3351 1322 3355 1323
rect 3351 1317 3355 1318
rect 3367 1322 3371 1323
rect 3418 1322 3424 1323
rect 3487 1322 3491 1323
rect 3518 1322 3524 1323
rect 3367 1317 3371 1318
rect 2338 1315 2344 1316
rect 2338 1311 2339 1315
rect 2343 1311 2344 1315
rect 2338 1310 2344 1311
rect 2520 1306 2522 1317
rect 2712 1306 2714 1317
rect 2762 1315 2768 1316
rect 2762 1311 2763 1315
rect 2767 1311 2768 1315
rect 2762 1310 2768 1311
rect 2310 1305 2316 1306
rect 2310 1301 2311 1305
rect 2315 1301 2316 1305
rect 2310 1300 2316 1301
rect 2518 1305 2524 1306
rect 2518 1301 2519 1305
rect 2523 1301 2524 1305
rect 2518 1300 2524 1301
rect 2710 1305 2716 1306
rect 2710 1301 2711 1305
rect 2715 1301 2716 1305
rect 2710 1300 2716 1301
rect 1862 1292 1868 1293
rect 1822 1288 1828 1289
rect 1822 1284 1823 1288
rect 1827 1284 1828 1288
rect 1862 1288 1863 1292
rect 1867 1288 1868 1292
rect 1862 1287 1868 1288
rect 2295 1292 2299 1293
rect 2443 1292 2447 1293
rect 2295 1287 2299 1288
rect 2442 1287 2448 1288
rect 1822 1283 1828 1284
rect 2442 1283 2443 1287
rect 2447 1283 2448 1287
rect 2442 1282 2448 1283
rect 1862 1275 1868 1276
rect 1822 1271 1828 1272
rect 1822 1267 1823 1271
rect 1827 1267 1828 1271
rect 1862 1271 1863 1275
rect 1867 1271 1868 1275
rect 1862 1270 1868 1271
rect 1822 1266 1828 1267
rect 1526 1261 1532 1262
rect 1526 1257 1527 1261
rect 1531 1257 1532 1261
rect 1526 1256 1532 1257
rect 1678 1261 1684 1262
rect 1678 1257 1679 1261
rect 1683 1257 1684 1261
rect 1678 1256 1684 1257
rect 1528 1247 1530 1256
rect 1680 1247 1682 1256
rect 1824 1247 1826 1266
rect 1864 1251 1866 1270
rect 2078 1265 2084 1266
rect 2078 1261 2079 1265
rect 2083 1261 2084 1265
rect 2078 1260 2084 1261
rect 2302 1265 2308 1266
rect 2302 1261 2303 1265
rect 2307 1261 2308 1265
rect 2302 1260 2308 1261
rect 2510 1265 2516 1266
rect 2510 1261 2511 1265
rect 2515 1261 2516 1265
rect 2510 1260 2516 1261
rect 2702 1265 2708 1266
rect 2702 1261 2703 1265
rect 2707 1261 2708 1265
rect 2702 1260 2708 1261
rect 2080 1251 2082 1260
rect 2130 1259 2136 1260
rect 2130 1255 2131 1259
rect 2135 1255 2136 1259
rect 2130 1254 2136 1255
rect 1863 1250 1867 1251
rect 1527 1246 1531 1247
rect 1527 1241 1531 1242
rect 1679 1246 1683 1247
rect 1679 1241 1683 1242
rect 1823 1246 1827 1247
rect 1863 1245 1867 1246
rect 1903 1250 1907 1251
rect 1903 1245 1907 1246
rect 1991 1250 1995 1251
rect 1991 1245 1995 1246
rect 2079 1250 2083 1251
rect 2079 1245 2083 1246
rect 2095 1250 2099 1251
rect 2095 1245 2099 1246
rect 1823 1241 1827 1242
rect 1528 1236 1530 1241
rect 1526 1235 1532 1236
rect 1526 1231 1527 1235
rect 1531 1231 1532 1235
rect 1526 1230 1532 1231
rect 614 1227 620 1228
rect 614 1223 615 1227
rect 619 1223 620 1227
rect 614 1222 620 1223
rect 1458 1227 1464 1228
rect 1458 1223 1459 1227
rect 1463 1223 1464 1227
rect 1824 1226 1826 1241
rect 1864 1230 1866 1245
rect 1904 1240 1906 1245
rect 1992 1240 1994 1245
rect 2096 1240 2098 1245
rect 1902 1239 1908 1240
rect 1902 1235 1903 1239
rect 1907 1235 1908 1239
rect 1902 1234 1908 1235
rect 1990 1239 1996 1240
rect 1990 1235 1991 1239
rect 1995 1235 1996 1239
rect 1990 1234 1996 1235
rect 2094 1239 2100 1240
rect 2094 1235 2095 1239
rect 2099 1235 2100 1239
rect 2094 1234 2100 1235
rect 1862 1229 1868 1230
rect 1458 1222 1464 1223
rect 1822 1225 1828 1226
rect 1822 1221 1823 1225
rect 1827 1221 1828 1225
rect 1862 1225 1863 1229
rect 1867 1225 1868 1229
rect 1862 1224 1868 1225
rect 1822 1220 1828 1221
rect 1970 1215 1976 1216
rect 1862 1212 1868 1213
rect 546 1211 552 1212
rect 546 1207 547 1211
rect 551 1207 552 1211
rect 546 1206 552 1207
rect 722 1211 728 1212
rect 722 1207 723 1211
rect 727 1207 728 1211
rect 722 1206 728 1207
rect 1822 1208 1828 1209
rect 302 1195 308 1196
rect 302 1191 303 1195
rect 307 1191 308 1195
rect 302 1190 308 1191
rect 486 1195 492 1196
rect 486 1191 487 1195
rect 491 1191 492 1195
rect 486 1190 492 1191
rect 210 1183 216 1184
rect 210 1179 211 1183
rect 215 1179 216 1183
rect 210 1178 216 1179
rect 304 1175 306 1190
rect 488 1175 490 1190
rect 111 1174 115 1175
rect 111 1169 115 1170
rect 143 1174 147 1175
rect 143 1169 147 1170
rect 167 1174 171 1175
rect 167 1169 171 1170
rect 303 1174 307 1175
rect 303 1169 307 1170
rect 319 1174 323 1175
rect 319 1169 323 1170
rect 471 1174 475 1175
rect 471 1169 475 1170
rect 487 1174 491 1175
rect 487 1169 491 1170
rect 112 1145 114 1169
rect 168 1158 170 1169
rect 234 1167 240 1168
rect 234 1163 235 1167
rect 239 1163 240 1167
rect 234 1162 240 1163
rect 166 1157 172 1158
rect 166 1153 167 1157
rect 171 1153 172 1157
rect 166 1152 172 1153
rect 110 1144 116 1145
rect 110 1140 111 1144
rect 115 1140 116 1144
rect 236 1140 238 1162
rect 320 1158 322 1169
rect 390 1167 396 1168
rect 390 1163 391 1167
rect 395 1163 396 1167
rect 390 1162 396 1163
rect 318 1157 324 1158
rect 318 1153 319 1157
rect 323 1153 324 1157
rect 318 1152 324 1153
rect 392 1140 394 1162
rect 472 1158 474 1169
rect 548 1168 550 1206
rect 662 1195 668 1196
rect 662 1191 663 1195
rect 667 1191 668 1195
rect 662 1190 668 1191
rect 664 1175 666 1190
rect 724 1184 726 1206
rect 1822 1204 1823 1208
rect 1827 1204 1828 1208
rect 1862 1208 1863 1212
rect 1867 1208 1868 1212
rect 1970 1211 1971 1215
rect 1975 1211 1976 1215
rect 1970 1210 1976 1211
rect 1978 1215 1984 1216
rect 1978 1211 1979 1215
rect 1983 1211 1984 1215
rect 1978 1210 1984 1211
rect 2086 1215 2092 1216
rect 2086 1211 2087 1215
rect 2091 1211 2092 1215
rect 2086 1210 2092 1211
rect 1862 1207 1868 1208
rect 1822 1203 1828 1204
rect 822 1195 828 1196
rect 822 1191 823 1195
rect 827 1191 828 1195
rect 822 1190 828 1191
rect 974 1195 980 1196
rect 974 1191 975 1195
rect 979 1191 980 1195
rect 974 1190 980 1191
rect 1118 1195 1124 1196
rect 1118 1191 1119 1195
rect 1123 1191 1124 1195
rect 1118 1190 1124 1191
rect 1254 1195 1260 1196
rect 1254 1191 1255 1195
rect 1259 1191 1260 1195
rect 1254 1190 1260 1191
rect 1390 1195 1396 1196
rect 1390 1191 1391 1195
rect 1395 1191 1396 1195
rect 1390 1190 1396 1191
rect 1534 1195 1540 1196
rect 1534 1191 1535 1195
rect 1539 1191 1540 1195
rect 1534 1190 1540 1191
rect 722 1183 728 1184
rect 722 1179 723 1183
rect 727 1179 728 1183
rect 722 1178 728 1179
rect 824 1175 826 1190
rect 976 1175 978 1190
rect 1050 1183 1056 1184
rect 1050 1179 1051 1183
rect 1055 1179 1056 1183
rect 1050 1178 1056 1179
rect 615 1174 619 1175
rect 615 1169 619 1170
rect 663 1174 667 1175
rect 663 1169 667 1170
rect 759 1174 763 1175
rect 759 1169 763 1170
rect 823 1174 827 1175
rect 823 1169 827 1170
rect 911 1174 915 1175
rect 911 1169 915 1170
rect 975 1174 979 1175
rect 975 1169 979 1170
rect 546 1167 552 1168
rect 546 1163 547 1167
rect 551 1163 552 1167
rect 546 1162 552 1163
rect 616 1158 618 1169
rect 646 1167 652 1168
rect 646 1163 647 1167
rect 651 1163 652 1167
rect 646 1162 652 1163
rect 470 1157 476 1158
rect 470 1153 471 1157
rect 475 1153 476 1157
rect 470 1152 476 1153
rect 614 1157 620 1158
rect 614 1153 615 1157
rect 619 1153 620 1157
rect 614 1152 620 1153
rect 110 1139 116 1140
rect 234 1139 240 1140
rect 234 1135 235 1139
rect 239 1135 240 1139
rect 234 1134 240 1135
rect 390 1139 396 1140
rect 390 1135 391 1139
rect 395 1135 396 1139
rect 390 1134 396 1135
rect 110 1127 116 1128
rect 110 1123 111 1127
rect 115 1123 116 1127
rect 110 1122 116 1123
rect 250 1127 256 1128
rect 250 1123 251 1127
rect 255 1123 256 1127
rect 250 1122 256 1123
rect 112 1103 114 1122
rect 158 1117 164 1118
rect 158 1113 159 1117
rect 163 1113 164 1117
rect 158 1112 164 1113
rect 160 1103 162 1112
rect 111 1102 115 1103
rect 111 1097 115 1098
rect 159 1102 163 1103
rect 159 1097 163 1098
rect 215 1102 219 1103
rect 215 1097 219 1098
rect 112 1082 114 1097
rect 216 1092 218 1097
rect 214 1091 220 1092
rect 214 1087 215 1091
rect 219 1087 220 1091
rect 214 1086 220 1087
rect 110 1081 116 1082
rect 110 1077 111 1081
rect 115 1077 116 1081
rect 110 1076 116 1077
rect 110 1064 116 1065
rect 110 1060 111 1064
rect 115 1060 116 1064
rect 110 1059 116 1060
rect 112 1027 114 1059
rect 222 1051 228 1052
rect 222 1047 223 1051
rect 227 1047 228 1051
rect 222 1046 228 1047
rect 224 1027 226 1046
rect 252 1040 254 1122
rect 310 1117 316 1118
rect 310 1113 311 1117
rect 315 1113 316 1117
rect 310 1112 316 1113
rect 462 1117 468 1118
rect 462 1113 463 1117
rect 467 1113 468 1117
rect 462 1112 468 1113
rect 606 1117 612 1118
rect 606 1113 607 1117
rect 611 1113 612 1117
rect 606 1112 612 1113
rect 312 1103 314 1112
rect 464 1103 466 1112
rect 608 1103 610 1112
rect 311 1102 315 1103
rect 311 1097 315 1098
rect 327 1102 331 1103
rect 327 1097 331 1098
rect 439 1102 443 1103
rect 439 1097 443 1098
rect 463 1102 467 1103
rect 463 1097 467 1098
rect 559 1102 563 1103
rect 559 1097 563 1098
rect 607 1102 611 1103
rect 607 1097 611 1098
rect 328 1092 330 1097
rect 440 1092 442 1097
rect 560 1092 562 1097
rect 326 1091 332 1092
rect 326 1087 327 1091
rect 331 1087 332 1091
rect 326 1086 332 1087
rect 438 1091 444 1092
rect 438 1087 439 1091
rect 443 1087 444 1091
rect 438 1086 444 1087
rect 558 1091 564 1092
rect 558 1087 559 1091
rect 563 1087 564 1091
rect 558 1086 564 1087
rect 648 1084 650 1162
rect 760 1158 762 1169
rect 912 1158 914 1169
rect 998 1167 1004 1168
rect 998 1163 999 1167
rect 1003 1163 1004 1167
rect 1052 1165 1054 1178
rect 1120 1175 1122 1190
rect 1256 1175 1258 1190
rect 1392 1175 1394 1190
rect 1536 1175 1538 1190
rect 1824 1175 1826 1203
rect 1864 1179 1866 1207
rect 1910 1199 1916 1200
rect 1910 1195 1911 1199
rect 1915 1195 1916 1199
rect 1910 1194 1916 1195
rect 1912 1179 1914 1194
rect 1863 1178 1867 1179
rect 1063 1174 1067 1175
rect 1063 1169 1067 1170
rect 1119 1174 1123 1175
rect 1119 1169 1123 1170
rect 1231 1174 1235 1175
rect 1231 1169 1235 1170
rect 1255 1174 1259 1175
rect 1255 1169 1259 1170
rect 1391 1174 1395 1175
rect 1391 1169 1395 1170
rect 1399 1174 1403 1175
rect 1399 1169 1403 1170
rect 1535 1174 1539 1175
rect 1535 1169 1539 1170
rect 1575 1174 1579 1175
rect 1575 1169 1579 1170
rect 1735 1174 1739 1175
rect 1735 1169 1739 1170
rect 1823 1174 1827 1175
rect 1863 1173 1867 1174
rect 1895 1178 1899 1179
rect 1895 1173 1899 1174
rect 1911 1178 1915 1179
rect 1911 1173 1915 1174
rect 1823 1169 1827 1170
rect 998 1162 1004 1163
rect 1051 1164 1055 1165
rect 758 1157 764 1158
rect 758 1153 759 1157
rect 763 1153 764 1157
rect 758 1152 764 1153
rect 910 1157 916 1158
rect 910 1153 911 1157
rect 915 1153 916 1157
rect 910 1152 916 1153
rect 750 1117 756 1118
rect 750 1113 751 1117
rect 755 1113 756 1117
rect 750 1112 756 1113
rect 902 1117 908 1118
rect 902 1113 903 1117
rect 907 1113 908 1117
rect 902 1112 908 1113
rect 752 1103 754 1112
rect 904 1103 906 1112
rect 679 1102 683 1103
rect 679 1097 683 1098
rect 751 1102 755 1103
rect 751 1097 755 1098
rect 807 1102 811 1103
rect 807 1097 811 1098
rect 903 1102 907 1103
rect 903 1097 907 1098
rect 943 1102 947 1103
rect 943 1097 947 1098
rect 680 1092 682 1097
rect 808 1092 810 1097
rect 944 1092 946 1097
rect 678 1091 684 1092
rect 678 1087 679 1091
rect 683 1087 684 1091
rect 678 1086 684 1087
rect 806 1091 812 1092
rect 806 1087 807 1091
rect 811 1087 812 1091
rect 806 1086 812 1087
rect 942 1091 948 1092
rect 942 1087 943 1091
rect 947 1087 948 1091
rect 942 1086 948 1087
rect 1000 1085 1002 1162
rect 1051 1159 1055 1160
rect 1064 1158 1066 1169
rect 1232 1158 1234 1169
rect 1400 1158 1402 1169
rect 1539 1164 1543 1165
rect 1539 1159 1543 1160
rect 1062 1157 1068 1158
rect 1062 1153 1063 1157
rect 1067 1153 1068 1157
rect 1062 1152 1068 1153
rect 1230 1157 1236 1158
rect 1230 1153 1231 1157
rect 1235 1153 1236 1157
rect 1230 1152 1236 1153
rect 1398 1157 1404 1158
rect 1398 1153 1399 1157
rect 1403 1153 1404 1157
rect 1398 1152 1404 1153
rect 1540 1140 1542 1159
rect 1576 1158 1578 1169
rect 1736 1158 1738 1169
rect 1574 1157 1580 1158
rect 1574 1153 1575 1157
rect 1579 1153 1580 1157
rect 1574 1152 1580 1153
rect 1734 1157 1740 1158
rect 1734 1153 1735 1157
rect 1739 1153 1740 1157
rect 1734 1152 1740 1153
rect 1824 1145 1826 1169
rect 1864 1149 1866 1173
rect 1870 1167 1876 1168
rect 1870 1163 1871 1167
rect 1875 1163 1876 1167
rect 1870 1162 1876 1163
rect 1896 1162 1898 1173
rect 1972 1172 1974 1210
rect 1980 1188 1982 1210
rect 1998 1199 2004 1200
rect 1998 1195 1999 1199
rect 2003 1195 2004 1199
rect 1998 1194 2004 1195
rect 1978 1187 1984 1188
rect 1978 1183 1979 1187
rect 1983 1183 1984 1187
rect 1978 1182 1984 1183
rect 2000 1179 2002 1194
rect 1999 1178 2003 1179
rect 1999 1173 2003 1174
rect 2063 1178 2067 1179
rect 2063 1173 2067 1174
rect 1970 1171 1976 1172
rect 1970 1167 1971 1171
rect 1975 1167 1976 1171
rect 1970 1166 1976 1167
rect 2064 1162 2066 1173
rect 2088 1172 2090 1210
rect 2102 1199 2108 1200
rect 2102 1195 2103 1199
rect 2107 1195 2108 1199
rect 2102 1194 2108 1195
rect 2104 1179 2106 1194
rect 2132 1188 2134 1254
rect 2304 1251 2306 1260
rect 2512 1251 2514 1260
rect 2704 1251 2706 1260
rect 2764 1252 2766 1310
rect 2888 1306 2890 1317
rect 3048 1306 3050 1317
rect 3114 1315 3120 1316
rect 3114 1311 3115 1315
rect 3119 1311 3120 1315
rect 3114 1310 3120 1311
rect 2886 1305 2892 1306
rect 2886 1301 2887 1305
rect 2891 1301 2892 1305
rect 2886 1300 2892 1301
rect 3046 1305 3052 1306
rect 3046 1301 3047 1305
rect 3051 1301 3052 1305
rect 3046 1300 3052 1301
rect 3116 1288 3118 1310
rect 3200 1306 3202 1317
rect 3352 1306 3354 1317
rect 3198 1305 3204 1306
rect 3198 1301 3199 1305
rect 3203 1301 3204 1305
rect 3198 1300 3204 1301
rect 3350 1305 3356 1306
rect 3350 1301 3351 1305
rect 3355 1301 3356 1305
rect 3350 1300 3356 1301
rect 3114 1287 3120 1288
rect 3114 1283 3115 1287
rect 3119 1283 3120 1287
rect 3114 1282 3120 1283
rect 2958 1275 2964 1276
rect 2958 1271 2959 1275
rect 2963 1271 2964 1275
rect 2958 1270 2964 1271
rect 2878 1265 2884 1266
rect 2878 1261 2879 1265
rect 2883 1261 2884 1265
rect 2878 1260 2884 1261
rect 2762 1251 2768 1252
rect 2880 1251 2882 1260
rect 2950 1259 2956 1260
rect 2950 1255 2951 1259
rect 2955 1255 2956 1259
rect 2950 1254 2956 1255
rect 2215 1250 2219 1251
rect 2215 1245 2219 1246
rect 2303 1250 2307 1251
rect 2303 1245 2307 1246
rect 2351 1250 2355 1251
rect 2351 1245 2355 1246
rect 2487 1250 2491 1251
rect 2487 1245 2491 1246
rect 2511 1250 2515 1251
rect 2511 1245 2515 1246
rect 2631 1250 2635 1251
rect 2631 1245 2635 1246
rect 2703 1250 2707 1251
rect 2762 1247 2763 1251
rect 2767 1247 2768 1251
rect 2762 1246 2768 1247
rect 2775 1250 2779 1251
rect 2703 1245 2707 1246
rect 2775 1245 2779 1246
rect 2879 1250 2883 1251
rect 2879 1245 2883 1246
rect 2919 1250 2923 1251
rect 2919 1245 2923 1246
rect 2216 1240 2218 1245
rect 2352 1240 2354 1245
rect 2488 1240 2490 1245
rect 2632 1240 2634 1245
rect 2776 1240 2778 1245
rect 2920 1240 2922 1245
rect 2214 1239 2220 1240
rect 2214 1235 2215 1239
rect 2219 1235 2220 1239
rect 2214 1234 2220 1235
rect 2350 1239 2356 1240
rect 2350 1235 2351 1239
rect 2355 1235 2356 1239
rect 2350 1234 2356 1235
rect 2486 1239 2492 1240
rect 2486 1235 2487 1239
rect 2491 1235 2492 1239
rect 2486 1234 2492 1235
rect 2630 1239 2636 1240
rect 2630 1235 2631 1239
rect 2635 1235 2636 1239
rect 2630 1234 2636 1235
rect 2774 1239 2780 1240
rect 2774 1235 2775 1239
rect 2779 1235 2780 1239
rect 2774 1234 2780 1235
rect 2918 1239 2924 1240
rect 2918 1235 2919 1239
rect 2923 1235 2924 1239
rect 2918 1234 2924 1235
rect 2554 1231 2560 1232
rect 2554 1227 2555 1231
rect 2559 1227 2560 1231
rect 2554 1226 2560 1227
rect 2162 1215 2168 1216
rect 2162 1211 2163 1215
rect 2167 1211 2168 1215
rect 2162 1210 2168 1211
rect 2282 1215 2288 1216
rect 2282 1211 2283 1215
rect 2287 1211 2288 1215
rect 2282 1210 2288 1211
rect 2164 1196 2166 1210
rect 2222 1199 2228 1200
rect 2162 1195 2168 1196
rect 2162 1191 2163 1195
rect 2167 1191 2168 1195
rect 2222 1195 2223 1199
rect 2227 1195 2228 1199
rect 2222 1194 2228 1195
rect 2162 1190 2168 1191
rect 2130 1187 2136 1188
rect 2130 1183 2131 1187
rect 2135 1183 2136 1187
rect 2130 1182 2136 1183
rect 2224 1179 2226 1194
rect 2284 1188 2286 1210
rect 2358 1199 2364 1200
rect 2358 1195 2359 1199
rect 2363 1195 2364 1199
rect 2358 1194 2364 1195
rect 2494 1199 2500 1200
rect 2494 1195 2495 1199
rect 2499 1195 2500 1199
rect 2556 1196 2558 1226
rect 2698 1215 2704 1216
rect 2698 1211 2699 1215
rect 2703 1211 2704 1215
rect 2698 1210 2704 1211
rect 2638 1199 2644 1200
rect 2494 1194 2500 1195
rect 2554 1195 2560 1196
rect 2282 1187 2288 1188
rect 2282 1183 2283 1187
rect 2287 1183 2288 1187
rect 2282 1182 2288 1183
rect 2360 1179 2362 1194
rect 2496 1179 2498 1194
rect 2554 1191 2555 1195
rect 2559 1191 2560 1195
rect 2638 1195 2639 1199
rect 2643 1195 2644 1199
rect 2638 1194 2644 1195
rect 2554 1190 2560 1191
rect 2640 1179 2642 1194
rect 2103 1178 2107 1179
rect 2103 1173 2107 1174
rect 2223 1178 2227 1179
rect 2223 1173 2227 1174
rect 2255 1178 2259 1179
rect 2255 1173 2259 1174
rect 2359 1178 2363 1179
rect 2359 1173 2363 1174
rect 2439 1178 2443 1179
rect 2439 1173 2443 1174
rect 2495 1178 2499 1179
rect 2495 1173 2499 1174
rect 2615 1178 2619 1179
rect 2615 1173 2619 1174
rect 2639 1178 2643 1179
rect 2639 1173 2643 1174
rect 2086 1171 2092 1172
rect 2086 1167 2087 1171
rect 2091 1167 2092 1171
rect 2086 1166 2092 1167
rect 2256 1162 2258 1173
rect 2440 1162 2442 1173
rect 2478 1171 2484 1172
rect 2478 1167 2479 1171
rect 2483 1167 2484 1171
rect 2478 1166 2484 1167
rect 1862 1148 1868 1149
rect 1822 1144 1828 1145
rect 1822 1140 1823 1144
rect 1827 1140 1828 1144
rect 1862 1144 1863 1148
rect 1867 1144 1868 1148
rect 1872 1144 1874 1162
rect 1894 1161 1900 1162
rect 1894 1157 1895 1161
rect 1899 1157 1900 1161
rect 1894 1156 1900 1157
rect 2062 1161 2068 1162
rect 2062 1157 2063 1161
rect 2067 1157 2068 1161
rect 2062 1156 2068 1157
rect 2254 1161 2260 1162
rect 2254 1157 2255 1161
rect 2259 1157 2260 1161
rect 2254 1156 2260 1157
rect 2438 1161 2444 1162
rect 2438 1157 2439 1161
rect 2443 1157 2444 1161
rect 2438 1156 2444 1157
rect 1862 1143 1868 1144
rect 1870 1143 1876 1144
rect 1538 1139 1544 1140
rect 1822 1139 1828 1140
rect 1870 1139 1871 1143
rect 1875 1139 1876 1143
rect 1538 1135 1539 1139
rect 1543 1135 1544 1139
rect 1870 1138 1876 1139
rect 1538 1134 1544 1135
rect 1862 1131 1868 1132
rect 1822 1127 1828 1128
rect 1822 1123 1823 1127
rect 1827 1123 1828 1127
rect 1862 1127 1863 1131
rect 1867 1127 1868 1131
rect 1862 1126 1868 1127
rect 2134 1131 2140 1132
rect 2134 1127 2135 1131
rect 2139 1127 2140 1131
rect 2134 1126 2140 1127
rect 1822 1122 1828 1123
rect 1054 1117 1060 1118
rect 1054 1113 1055 1117
rect 1059 1113 1060 1117
rect 1054 1112 1060 1113
rect 1222 1117 1228 1118
rect 1222 1113 1223 1117
rect 1227 1113 1228 1117
rect 1222 1112 1228 1113
rect 1390 1117 1396 1118
rect 1390 1113 1391 1117
rect 1395 1113 1396 1117
rect 1390 1112 1396 1113
rect 1566 1117 1572 1118
rect 1566 1113 1567 1117
rect 1571 1113 1572 1117
rect 1566 1112 1572 1113
rect 1726 1117 1732 1118
rect 1726 1113 1727 1117
rect 1731 1113 1732 1117
rect 1726 1112 1732 1113
rect 1056 1103 1058 1112
rect 1224 1103 1226 1112
rect 1392 1103 1394 1112
rect 1568 1103 1570 1112
rect 1728 1103 1730 1112
rect 1766 1111 1772 1112
rect 1766 1107 1767 1111
rect 1771 1107 1772 1111
rect 1766 1106 1772 1107
rect 1055 1102 1059 1103
rect 1055 1097 1059 1098
rect 1087 1102 1091 1103
rect 1087 1097 1091 1098
rect 1223 1102 1227 1103
rect 1223 1097 1227 1098
rect 1247 1102 1251 1103
rect 1247 1097 1251 1098
rect 1391 1102 1395 1103
rect 1391 1097 1395 1098
rect 1407 1102 1411 1103
rect 1407 1097 1411 1098
rect 1567 1102 1571 1103
rect 1567 1097 1571 1098
rect 1575 1102 1579 1103
rect 1575 1097 1579 1098
rect 1727 1102 1731 1103
rect 1727 1097 1731 1098
rect 1088 1092 1090 1097
rect 1248 1092 1250 1097
rect 1408 1092 1410 1097
rect 1576 1092 1578 1097
rect 1728 1092 1730 1097
rect 1086 1091 1092 1092
rect 1086 1087 1087 1091
rect 1091 1087 1092 1091
rect 1086 1086 1092 1087
rect 1246 1091 1252 1092
rect 1246 1087 1247 1091
rect 1251 1087 1252 1091
rect 1246 1086 1252 1087
rect 1406 1091 1412 1092
rect 1406 1087 1407 1091
rect 1411 1087 1412 1091
rect 1406 1086 1412 1087
rect 1574 1091 1580 1092
rect 1574 1087 1575 1091
rect 1579 1087 1580 1091
rect 1574 1086 1580 1087
rect 1726 1091 1732 1092
rect 1726 1087 1727 1091
rect 1731 1087 1732 1091
rect 1726 1086 1732 1087
rect 999 1084 1003 1085
rect 1339 1084 1343 1085
rect 646 1083 652 1084
rect 646 1079 647 1083
rect 651 1079 652 1083
rect 999 1079 1003 1080
rect 1338 1079 1339 1084
rect 1343 1079 1344 1084
rect 646 1078 652 1079
rect 1338 1078 1344 1079
rect 1566 1067 1572 1068
rect 1566 1063 1567 1067
rect 1571 1063 1572 1067
rect 1566 1062 1572 1063
rect 1642 1067 1648 1068
rect 1642 1063 1643 1067
rect 1647 1063 1648 1067
rect 1642 1062 1648 1063
rect 334 1051 340 1052
rect 334 1047 335 1051
rect 339 1047 340 1051
rect 334 1046 340 1047
rect 446 1051 452 1052
rect 446 1047 447 1051
rect 451 1047 452 1051
rect 446 1046 452 1047
rect 566 1051 572 1052
rect 566 1047 567 1051
rect 571 1047 572 1051
rect 566 1046 572 1047
rect 686 1051 692 1052
rect 686 1047 687 1051
rect 691 1047 692 1051
rect 686 1046 692 1047
rect 814 1051 820 1052
rect 814 1047 815 1051
rect 819 1047 820 1051
rect 814 1046 820 1047
rect 950 1051 956 1052
rect 950 1047 951 1051
rect 955 1047 956 1051
rect 950 1046 956 1047
rect 1094 1051 1100 1052
rect 1094 1047 1095 1051
rect 1099 1047 1100 1051
rect 1094 1046 1100 1047
rect 1254 1051 1260 1052
rect 1254 1047 1255 1051
rect 1259 1047 1260 1051
rect 1254 1046 1260 1047
rect 1414 1051 1420 1052
rect 1414 1047 1415 1051
rect 1419 1047 1420 1051
rect 1414 1046 1420 1047
rect 250 1039 256 1040
rect 250 1035 251 1039
rect 255 1035 256 1039
rect 250 1034 256 1035
rect 336 1027 338 1046
rect 448 1027 450 1046
rect 568 1027 570 1046
rect 688 1027 690 1046
rect 714 1039 720 1040
rect 714 1035 715 1039
rect 719 1035 720 1039
rect 714 1034 720 1035
rect 111 1026 115 1027
rect 111 1021 115 1022
rect 223 1026 227 1027
rect 223 1021 227 1022
rect 335 1026 339 1027
rect 335 1021 339 1022
rect 343 1026 347 1027
rect 343 1021 347 1022
rect 431 1026 435 1027
rect 431 1021 435 1022
rect 447 1026 451 1027
rect 447 1021 451 1022
rect 535 1026 539 1027
rect 535 1021 539 1022
rect 567 1026 571 1027
rect 567 1021 571 1022
rect 655 1026 659 1027
rect 655 1021 659 1022
rect 687 1026 691 1027
rect 687 1021 691 1022
rect 112 997 114 1021
rect 344 1010 346 1021
rect 410 1019 416 1020
rect 410 1015 411 1019
rect 415 1015 416 1019
rect 410 1014 416 1015
rect 342 1009 348 1010
rect 342 1005 343 1009
rect 347 1005 348 1009
rect 342 1004 348 1005
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 412 992 414 1014
rect 432 1010 434 1021
rect 502 1019 508 1020
rect 502 1015 503 1019
rect 507 1015 508 1019
rect 502 1014 508 1015
rect 430 1009 436 1010
rect 430 1005 431 1009
rect 435 1005 436 1009
rect 430 1004 436 1005
rect 504 992 506 1014
rect 536 1010 538 1021
rect 656 1010 658 1021
rect 534 1009 540 1010
rect 534 1005 535 1009
rect 539 1005 540 1009
rect 534 1004 540 1005
rect 654 1009 660 1010
rect 654 1005 655 1009
rect 659 1005 660 1009
rect 654 1004 660 1005
rect 716 996 718 1034
rect 816 1027 818 1046
rect 858 1039 864 1040
rect 858 1035 859 1039
rect 863 1035 864 1039
rect 858 1034 864 1035
rect 791 1026 795 1027
rect 791 1021 795 1022
rect 815 1026 819 1027
rect 815 1021 819 1022
rect 722 1019 728 1020
rect 722 1015 723 1019
rect 727 1015 728 1019
rect 722 1014 728 1015
rect 714 995 720 996
rect 110 991 116 992
rect 410 991 416 992
rect 410 987 411 991
rect 415 987 416 991
rect 410 986 416 987
rect 502 991 508 992
rect 502 987 503 991
rect 507 987 508 991
rect 714 991 715 995
rect 719 991 720 995
rect 724 992 726 1014
rect 792 1010 794 1021
rect 822 1019 828 1020
rect 822 1015 823 1019
rect 827 1015 828 1019
rect 822 1014 828 1015
rect 790 1009 796 1010
rect 790 1005 791 1009
rect 795 1005 796 1009
rect 790 1004 796 1005
rect 714 990 720 991
rect 722 991 728 992
rect 502 986 508 987
rect 722 987 723 991
rect 727 987 728 991
rect 722 986 728 987
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 110 974 116 975
rect 112 955 114 974
rect 334 969 340 970
rect 334 965 335 969
rect 339 965 340 969
rect 334 964 340 965
rect 422 969 428 970
rect 422 965 423 969
rect 427 965 428 969
rect 422 964 428 965
rect 526 969 532 970
rect 526 965 527 969
rect 531 965 532 969
rect 526 964 532 965
rect 646 969 652 970
rect 646 965 647 969
rect 651 965 652 969
rect 646 964 652 965
rect 782 969 788 970
rect 782 965 783 969
rect 787 965 788 969
rect 782 964 788 965
rect 336 955 338 964
rect 402 963 408 964
rect 402 959 403 963
rect 407 959 408 963
rect 402 958 408 959
rect 111 954 115 955
rect 111 949 115 950
rect 335 954 339 955
rect 335 949 339 950
rect 367 954 371 955
rect 367 949 371 950
rect 112 934 114 949
rect 368 944 370 949
rect 366 943 372 944
rect 366 939 367 943
rect 371 939 372 943
rect 366 938 372 939
rect 110 933 116 934
rect 110 929 111 933
rect 115 929 116 933
rect 110 928 116 929
rect 110 916 116 917
rect 110 912 111 916
rect 115 912 116 916
rect 110 911 116 912
rect 112 883 114 911
rect 374 903 380 904
rect 374 899 375 903
rect 379 899 380 903
rect 374 898 380 899
rect 376 883 378 898
rect 404 892 406 958
rect 424 955 426 964
rect 528 955 530 964
rect 648 955 650 964
rect 784 955 786 964
rect 423 954 427 955
rect 423 949 427 950
rect 463 954 467 955
rect 463 949 467 950
rect 527 954 531 955
rect 527 949 531 950
rect 575 954 579 955
rect 575 949 579 950
rect 647 954 651 955
rect 647 949 651 950
rect 703 954 707 955
rect 703 949 707 950
rect 783 954 787 955
rect 783 949 787 950
rect 464 944 466 949
rect 576 944 578 949
rect 704 944 706 949
rect 462 943 468 944
rect 462 939 463 943
rect 467 939 468 943
rect 462 938 468 939
rect 574 943 580 944
rect 574 939 575 943
rect 579 939 580 943
rect 574 938 580 939
rect 702 943 708 944
rect 702 939 703 943
rect 707 939 708 943
rect 702 938 708 939
rect 824 936 826 1014
rect 860 992 862 1034
rect 952 1027 954 1046
rect 1096 1027 1098 1046
rect 1256 1027 1258 1046
rect 1416 1027 1418 1046
rect 951 1026 955 1027
rect 951 1021 955 1022
rect 1095 1026 1099 1027
rect 1095 1021 1099 1022
rect 1135 1026 1139 1027
rect 1135 1021 1139 1022
rect 1255 1026 1259 1027
rect 1255 1021 1259 1022
rect 1327 1026 1331 1027
rect 1327 1021 1331 1022
rect 1415 1026 1419 1027
rect 1415 1021 1419 1022
rect 1535 1026 1539 1027
rect 1535 1021 1539 1022
rect 952 1010 954 1021
rect 1038 1019 1044 1020
rect 1038 1015 1039 1019
rect 1043 1015 1044 1019
rect 1038 1014 1044 1015
rect 950 1009 956 1010
rect 950 1005 951 1009
rect 955 1005 956 1009
rect 950 1004 956 1005
rect 1040 992 1042 1014
rect 1136 1010 1138 1021
rect 1202 1019 1208 1020
rect 1202 1015 1203 1019
rect 1207 1015 1208 1019
rect 1202 1014 1208 1015
rect 1278 1019 1284 1020
rect 1278 1015 1279 1019
rect 1283 1015 1284 1019
rect 1278 1014 1284 1015
rect 1134 1009 1140 1010
rect 1134 1005 1135 1009
rect 1139 1005 1140 1009
rect 1134 1004 1140 1005
rect 1204 992 1206 1014
rect 858 991 864 992
rect 858 987 859 991
rect 863 987 864 991
rect 858 986 864 987
rect 1038 991 1044 992
rect 1038 987 1039 991
rect 1043 987 1044 991
rect 1038 986 1044 987
rect 1202 991 1208 992
rect 1202 987 1203 991
rect 1207 987 1208 991
rect 1202 986 1208 987
rect 942 969 948 970
rect 942 965 943 969
rect 947 965 948 969
rect 942 964 948 965
rect 1126 969 1132 970
rect 1126 965 1127 969
rect 1131 965 1132 969
rect 1126 964 1132 965
rect 944 955 946 964
rect 1128 955 1130 964
rect 847 954 851 955
rect 847 949 851 950
rect 943 954 947 955
rect 943 949 947 950
rect 1007 954 1011 955
rect 1007 949 1011 950
rect 1127 954 1131 955
rect 1127 949 1131 950
rect 1175 954 1179 955
rect 1175 949 1179 950
rect 848 944 850 949
rect 1008 944 1010 949
rect 1176 944 1178 949
rect 846 943 852 944
rect 846 939 847 943
rect 851 939 852 943
rect 846 938 852 939
rect 1006 943 1012 944
rect 1006 939 1007 943
rect 1011 939 1012 943
rect 1006 938 1012 939
rect 1174 943 1180 944
rect 1174 939 1175 943
rect 1179 939 1180 943
rect 1174 938 1180 939
rect 1280 936 1282 1014
rect 1328 1010 1330 1021
rect 1536 1010 1538 1021
rect 1568 1020 1570 1062
rect 1582 1051 1588 1052
rect 1582 1047 1583 1051
rect 1587 1047 1588 1051
rect 1582 1046 1588 1047
rect 1584 1027 1586 1046
rect 1644 1040 1646 1062
rect 1734 1051 1740 1052
rect 1734 1047 1735 1051
rect 1739 1047 1740 1051
rect 1734 1046 1740 1047
rect 1642 1039 1648 1040
rect 1642 1035 1643 1039
rect 1647 1035 1648 1039
rect 1642 1034 1648 1035
rect 1736 1027 1738 1046
rect 1768 1040 1770 1106
rect 1824 1103 1826 1122
rect 1823 1102 1827 1103
rect 1864 1099 1866 1126
rect 1886 1121 1892 1122
rect 1886 1117 1887 1121
rect 1891 1117 1892 1121
rect 1886 1116 1892 1117
rect 2054 1121 2060 1122
rect 2054 1117 2055 1121
rect 2059 1117 2060 1121
rect 2054 1116 2060 1117
rect 1888 1099 1890 1116
rect 2056 1099 2058 1116
rect 1823 1097 1827 1098
rect 1863 1098 1867 1099
rect 1824 1082 1826 1097
rect 1863 1093 1867 1094
rect 1887 1098 1891 1099
rect 1887 1093 1891 1094
rect 1935 1098 1939 1099
rect 1935 1093 1939 1094
rect 2055 1098 2059 1099
rect 2055 1093 2059 1094
rect 2095 1098 2099 1099
rect 2095 1093 2099 1094
rect 1822 1081 1828 1082
rect 1822 1077 1823 1081
rect 1827 1077 1828 1081
rect 1864 1078 1866 1093
rect 1936 1088 1938 1093
rect 2096 1088 2098 1093
rect 1934 1087 1940 1088
rect 1934 1083 1935 1087
rect 1939 1083 1940 1087
rect 1934 1082 1940 1083
rect 2094 1087 2100 1088
rect 2094 1083 2095 1087
rect 2099 1083 2100 1087
rect 2094 1082 2100 1083
rect 2010 1079 2016 1080
rect 1822 1076 1828 1077
rect 1862 1077 1868 1078
rect 1862 1073 1863 1077
rect 1867 1073 1868 1077
rect 2010 1075 2011 1079
rect 2015 1075 2016 1079
rect 2010 1074 2016 1075
rect 1862 1072 1868 1073
rect 1822 1064 1828 1065
rect 1822 1060 1823 1064
rect 1827 1060 1828 1064
rect 2002 1063 2008 1064
rect 1822 1059 1828 1060
rect 1862 1060 1868 1061
rect 1766 1039 1772 1040
rect 1766 1035 1767 1039
rect 1771 1035 1772 1039
rect 1766 1034 1772 1035
rect 1824 1027 1826 1059
rect 1862 1056 1863 1060
rect 1867 1056 1868 1060
rect 2002 1059 2003 1063
rect 2007 1059 2008 1063
rect 2002 1058 2008 1059
rect 1862 1055 1868 1056
rect 1864 1027 1866 1055
rect 1942 1047 1948 1048
rect 1942 1043 1943 1047
rect 1947 1043 1948 1047
rect 1942 1042 1948 1043
rect 1944 1027 1946 1042
rect 2004 1036 2006 1058
rect 2002 1035 2008 1036
rect 2002 1031 2003 1035
rect 2007 1031 2008 1035
rect 2002 1030 2008 1031
rect 1583 1026 1587 1027
rect 1583 1021 1587 1022
rect 1735 1026 1739 1027
rect 1735 1021 1739 1022
rect 1823 1026 1827 1027
rect 1823 1021 1827 1022
rect 1863 1026 1867 1027
rect 1863 1021 1867 1022
rect 1943 1026 1947 1027
rect 1943 1021 1947 1022
rect 1566 1019 1572 1020
rect 1566 1015 1567 1019
rect 1571 1015 1572 1019
rect 1566 1014 1572 1015
rect 1736 1010 1738 1021
rect 1326 1009 1332 1010
rect 1326 1005 1327 1009
rect 1331 1005 1332 1009
rect 1326 1004 1332 1005
rect 1534 1009 1540 1010
rect 1534 1005 1535 1009
rect 1539 1005 1540 1009
rect 1534 1004 1540 1005
rect 1734 1009 1740 1010
rect 1734 1005 1735 1009
rect 1739 1005 1740 1009
rect 1734 1004 1740 1005
rect 1824 997 1826 1021
rect 1864 997 1866 1021
rect 1944 1010 1946 1021
rect 2012 1020 2014 1074
rect 2102 1047 2108 1048
rect 2102 1043 2103 1047
rect 2107 1043 2108 1047
rect 2102 1042 2108 1043
rect 2104 1027 2106 1042
rect 2136 1036 2138 1126
rect 2246 1121 2252 1122
rect 2246 1117 2247 1121
rect 2251 1117 2252 1121
rect 2246 1116 2252 1117
rect 2430 1121 2436 1122
rect 2430 1117 2431 1121
rect 2435 1117 2436 1121
rect 2430 1116 2436 1117
rect 2248 1099 2250 1116
rect 2432 1099 2434 1116
rect 2247 1098 2251 1099
rect 2247 1093 2251 1094
rect 2407 1098 2411 1099
rect 2407 1093 2411 1094
rect 2431 1098 2435 1099
rect 2431 1093 2435 1094
rect 2248 1088 2250 1093
rect 2408 1088 2410 1093
rect 2246 1087 2252 1088
rect 2246 1083 2247 1087
rect 2251 1083 2252 1087
rect 2246 1082 2252 1083
rect 2406 1087 2412 1088
rect 2406 1083 2407 1087
rect 2411 1083 2412 1087
rect 2406 1082 2412 1083
rect 2480 1080 2482 1166
rect 2616 1162 2618 1173
rect 2700 1172 2702 1210
rect 2782 1199 2788 1200
rect 2782 1195 2783 1199
rect 2787 1195 2788 1199
rect 2926 1199 2932 1200
rect 2782 1194 2788 1195
rect 2815 1196 2819 1197
rect 2784 1179 2786 1194
rect 2926 1195 2927 1199
rect 2931 1195 2932 1199
rect 2926 1194 2932 1195
rect 2815 1191 2819 1192
rect 2816 1188 2818 1191
rect 2814 1187 2820 1188
rect 2814 1183 2815 1187
rect 2819 1183 2820 1187
rect 2814 1182 2820 1183
rect 2928 1179 2930 1194
rect 2952 1188 2954 1254
rect 2960 1252 2962 1270
rect 3038 1265 3044 1266
rect 3038 1261 3039 1265
rect 3043 1261 3044 1265
rect 3038 1260 3044 1261
rect 3190 1265 3196 1266
rect 3190 1261 3191 1265
rect 3195 1261 3196 1265
rect 3190 1260 3196 1261
rect 3342 1265 3348 1266
rect 3342 1261 3343 1265
rect 3347 1261 3348 1265
rect 3342 1260 3348 1261
rect 2958 1251 2964 1252
rect 3040 1251 3042 1260
rect 3192 1251 3194 1260
rect 3344 1251 3346 1260
rect 2958 1247 2959 1251
rect 2963 1247 2964 1251
rect 2958 1246 2964 1247
rect 3039 1250 3043 1251
rect 3039 1245 3043 1246
rect 3063 1250 3067 1251
rect 3063 1245 3067 1246
rect 3191 1250 3195 1251
rect 3191 1245 3195 1246
rect 3207 1250 3211 1251
rect 3207 1245 3211 1246
rect 3343 1250 3347 1251
rect 3343 1245 3347 1246
rect 3351 1250 3355 1251
rect 3351 1245 3355 1246
rect 3064 1240 3066 1245
rect 3208 1240 3210 1245
rect 3352 1240 3354 1245
rect 3062 1239 3068 1240
rect 3062 1235 3063 1239
rect 3067 1235 3068 1239
rect 3062 1234 3068 1235
rect 3206 1239 3212 1240
rect 3206 1235 3207 1239
rect 3211 1235 3212 1239
rect 3206 1234 3212 1235
rect 3350 1239 3356 1240
rect 3350 1235 3351 1239
rect 3355 1235 3356 1239
rect 3350 1234 3356 1235
rect 3420 1232 3422 1322
rect 3487 1317 3491 1318
rect 3488 1306 3490 1317
rect 3548 1316 3550 1350
rect 3574 1348 3575 1352
rect 3579 1348 3580 1352
rect 3574 1347 3580 1348
rect 3576 1323 3578 1347
rect 3575 1322 3579 1323
rect 3575 1317 3579 1318
rect 3546 1315 3552 1316
rect 3546 1311 3547 1315
rect 3551 1311 3552 1315
rect 3546 1310 3552 1311
rect 3486 1305 3492 1306
rect 3486 1301 3487 1305
rect 3491 1301 3492 1305
rect 3486 1300 3492 1301
rect 3576 1293 3578 1317
rect 3574 1292 3580 1293
rect 3574 1288 3575 1292
rect 3579 1288 3580 1292
rect 3574 1287 3580 1288
rect 3574 1275 3580 1276
rect 3574 1271 3575 1275
rect 3579 1271 3580 1275
rect 3574 1270 3580 1271
rect 3478 1265 3484 1266
rect 3478 1261 3479 1265
rect 3483 1261 3484 1265
rect 3478 1260 3484 1261
rect 3480 1251 3482 1260
rect 3518 1259 3524 1260
rect 3518 1255 3519 1259
rect 3523 1255 3524 1259
rect 3518 1254 3524 1255
rect 3479 1250 3483 1251
rect 3479 1245 3483 1246
rect 3480 1240 3482 1245
rect 3478 1239 3484 1240
rect 3478 1235 3479 1239
rect 3483 1235 3484 1239
rect 3478 1234 3484 1235
rect 3138 1231 3144 1232
rect 3138 1227 3139 1231
rect 3143 1227 3144 1231
rect 3138 1226 3144 1227
rect 3418 1231 3424 1232
rect 3418 1227 3419 1231
rect 3423 1227 3424 1231
rect 3418 1226 3424 1227
rect 3070 1199 3076 1200
rect 3070 1195 3071 1199
rect 3075 1195 3076 1199
rect 3140 1197 3142 1226
rect 3214 1199 3220 1200
rect 3070 1194 3076 1195
rect 3139 1196 3143 1197
rect 2950 1187 2956 1188
rect 2950 1183 2951 1187
rect 2955 1183 2956 1187
rect 2950 1182 2956 1183
rect 3072 1179 3074 1194
rect 3214 1195 3215 1199
rect 3219 1195 3220 1199
rect 3214 1194 3220 1195
rect 3358 1199 3364 1200
rect 3358 1195 3359 1199
rect 3363 1195 3364 1199
rect 3358 1194 3364 1195
rect 3486 1199 3492 1200
rect 3486 1195 3487 1199
rect 3491 1195 3492 1199
rect 3486 1194 3492 1195
rect 3139 1191 3143 1192
rect 3216 1179 3218 1194
rect 3360 1179 3362 1194
rect 3386 1187 3392 1188
rect 3386 1183 3387 1187
rect 3391 1183 3392 1187
rect 3386 1182 3392 1183
rect 2783 1178 2787 1179
rect 2783 1173 2787 1174
rect 2791 1178 2795 1179
rect 2791 1173 2795 1174
rect 2927 1178 2931 1179
rect 2927 1173 2931 1174
rect 2967 1178 2971 1179
rect 2967 1173 2971 1174
rect 3071 1178 3075 1179
rect 3071 1173 3075 1174
rect 3143 1178 3147 1179
rect 3143 1173 3147 1174
rect 3215 1178 3219 1179
rect 3215 1173 3219 1174
rect 3327 1178 3331 1179
rect 3327 1173 3331 1174
rect 3359 1178 3363 1179
rect 3359 1173 3363 1174
rect 2698 1171 2704 1172
rect 2698 1167 2699 1171
rect 2703 1167 2704 1171
rect 2698 1166 2704 1167
rect 2792 1162 2794 1173
rect 2968 1162 2970 1173
rect 3144 1162 3146 1173
rect 3328 1162 3330 1173
rect 3354 1167 3360 1168
rect 3354 1163 3355 1167
rect 3359 1163 3360 1167
rect 3354 1162 3360 1163
rect 2614 1161 2620 1162
rect 2614 1157 2615 1161
rect 2619 1157 2620 1161
rect 2614 1156 2620 1157
rect 2790 1161 2796 1162
rect 2790 1157 2791 1161
rect 2795 1157 2796 1161
rect 2790 1156 2796 1157
rect 2966 1161 2972 1162
rect 2966 1157 2967 1161
rect 2971 1157 2972 1161
rect 2966 1156 2972 1157
rect 3142 1161 3148 1162
rect 3142 1157 3143 1161
rect 3147 1157 3148 1161
rect 3142 1156 3148 1157
rect 3326 1161 3332 1162
rect 3326 1157 3327 1161
rect 3331 1157 3332 1161
rect 3326 1156 3332 1157
rect 3142 1131 3148 1132
rect 3142 1127 3143 1131
rect 3147 1127 3148 1131
rect 3142 1126 3148 1127
rect 2606 1121 2612 1122
rect 2606 1117 2607 1121
rect 2611 1117 2612 1121
rect 2606 1116 2612 1117
rect 2782 1121 2788 1122
rect 2782 1117 2783 1121
rect 2787 1117 2788 1121
rect 2782 1116 2788 1117
rect 2958 1121 2964 1122
rect 2958 1117 2959 1121
rect 2963 1117 2964 1121
rect 2958 1116 2964 1117
rect 3134 1121 3140 1122
rect 3134 1117 3135 1121
rect 3139 1117 3140 1121
rect 3134 1116 3140 1117
rect 2608 1099 2610 1116
rect 2784 1099 2786 1116
rect 2960 1099 2962 1116
rect 3136 1099 3138 1116
rect 2567 1098 2571 1099
rect 2567 1093 2571 1094
rect 2607 1098 2611 1099
rect 2607 1093 2611 1094
rect 2735 1098 2739 1099
rect 2735 1093 2739 1094
rect 2783 1098 2787 1099
rect 2783 1093 2787 1094
rect 2911 1098 2915 1099
rect 2911 1093 2915 1094
rect 2959 1098 2963 1099
rect 2959 1093 2963 1094
rect 3095 1098 3099 1099
rect 3095 1093 3099 1094
rect 3135 1098 3139 1099
rect 3135 1093 3139 1094
rect 2568 1088 2570 1093
rect 2736 1088 2738 1093
rect 2912 1088 2914 1093
rect 3096 1088 3098 1093
rect 2566 1087 2572 1088
rect 2566 1083 2567 1087
rect 2571 1083 2572 1087
rect 2566 1082 2572 1083
rect 2734 1087 2740 1088
rect 2734 1083 2735 1087
rect 2739 1083 2740 1087
rect 2734 1082 2740 1083
rect 2910 1087 2916 1088
rect 2910 1083 2911 1087
rect 2915 1083 2916 1087
rect 2910 1082 2916 1083
rect 3094 1087 3100 1088
rect 3094 1083 3095 1087
rect 3099 1083 3100 1087
rect 3094 1082 3100 1083
rect 2478 1079 2484 1080
rect 2478 1075 2479 1079
rect 2483 1075 2484 1079
rect 2478 1074 2484 1075
rect 2642 1079 2648 1080
rect 2642 1075 2643 1079
rect 2647 1075 2648 1079
rect 2642 1074 2648 1075
rect 2634 1063 2640 1064
rect 2634 1059 2635 1063
rect 2639 1059 2640 1063
rect 2634 1058 2640 1059
rect 2254 1047 2260 1048
rect 2254 1043 2255 1047
rect 2259 1043 2260 1047
rect 2254 1042 2260 1043
rect 2414 1047 2420 1048
rect 2414 1043 2415 1047
rect 2419 1043 2420 1047
rect 2414 1042 2420 1043
rect 2574 1047 2580 1048
rect 2574 1043 2575 1047
rect 2579 1043 2580 1047
rect 2574 1042 2580 1043
rect 2134 1035 2140 1036
rect 2134 1031 2135 1035
rect 2139 1031 2140 1035
rect 2134 1030 2140 1031
rect 2256 1027 2258 1042
rect 2378 1035 2384 1036
rect 2378 1031 2379 1035
rect 2383 1031 2384 1035
rect 2378 1030 2384 1031
rect 2071 1026 2075 1027
rect 2071 1021 2075 1022
rect 2103 1026 2107 1027
rect 2103 1021 2107 1022
rect 2191 1026 2195 1027
rect 2191 1021 2195 1022
rect 2255 1026 2259 1027
rect 2255 1021 2259 1022
rect 2311 1026 2315 1027
rect 2311 1021 2315 1022
rect 2010 1019 2016 1020
rect 2010 1015 2011 1019
rect 2015 1015 2016 1019
rect 2010 1014 2016 1015
rect 2072 1010 2074 1021
rect 2114 1019 2120 1020
rect 2114 1015 2115 1019
rect 2119 1015 2120 1019
rect 2114 1014 2120 1015
rect 1942 1009 1948 1010
rect 1942 1005 1943 1009
rect 1947 1005 1948 1009
rect 1942 1004 1948 1005
rect 2070 1009 2076 1010
rect 2070 1005 2071 1009
rect 2075 1005 2076 1009
rect 2070 1004 2076 1005
rect 1822 996 1828 997
rect 1822 992 1823 996
rect 1827 992 1828 996
rect 1822 991 1828 992
rect 1862 996 1868 997
rect 1862 992 1863 996
rect 1867 992 1868 996
rect 1862 991 1868 992
rect 1734 979 1740 980
rect 1734 975 1735 979
rect 1739 975 1740 979
rect 1734 974 1740 975
rect 1822 979 1828 980
rect 1822 975 1823 979
rect 1827 975 1828 979
rect 1822 974 1828 975
rect 1862 979 1868 980
rect 1862 975 1863 979
rect 1867 975 1868 979
rect 1862 974 1868 975
rect 1942 979 1948 980
rect 1942 975 1943 979
rect 1947 975 1948 979
rect 1942 974 1948 975
rect 1318 969 1324 970
rect 1318 965 1319 969
rect 1323 965 1324 969
rect 1318 964 1324 965
rect 1526 969 1532 970
rect 1526 965 1527 969
rect 1531 965 1532 969
rect 1526 964 1532 965
rect 1726 969 1732 970
rect 1726 965 1727 969
rect 1731 965 1732 969
rect 1726 964 1732 965
rect 1320 955 1322 964
rect 1528 955 1530 964
rect 1728 955 1730 964
rect 1319 954 1323 955
rect 1319 949 1323 950
rect 1351 954 1355 955
rect 1351 949 1355 950
rect 1527 954 1531 955
rect 1527 949 1531 950
rect 1711 954 1715 955
rect 1711 949 1715 950
rect 1727 954 1731 955
rect 1727 949 1731 950
rect 1352 944 1354 949
rect 1528 944 1530 949
rect 1712 944 1714 949
rect 1350 943 1356 944
rect 1350 939 1351 943
rect 1355 939 1356 943
rect 1350 938 1356 939
rect 1526 943 1532 944
rect 1526 939 1527 943
rect 1531 939 1532 943
rect 1526 938 1532 939
rect 1710 943 1716 944
rect 1710 939 1711 943
rect 1715 939 1716 943
rect 1710 938 1716 939
rect 822 935 828 936
rect 822 931 823 935
rect 827 931 828 935
rect 822 930 828 931
rect 1278 935 1284 936
rect 1278 931 1279 935
rect 1283 931 1284 935
rect 1278 930 1284 931
rect 562 919 568 920
rect 562 915 563 919
rect 567 915 568 919
rect 562 914 568 915
rect 1166 919 1172 920
rect 1166 915 1167 919
rect 1171 915 1172 919
rect 1166 914 1172 915
rect 1658 919 1664 920
rect 1658 915 1659 919
rect 1663 915 1664 919
rect 1658 914 1664 915
rect 1666 919 1672 920
rect 1666 915 1667 919
rect 1671 915 1672 919
rect 1666 914 1672 915
rect 470 903 476 904
rect 470 899 471 903
rect 475 899 476 903
rect 470 898 476 899
rect 402 891 408 892
rect 402 887 403 891
rect 407 887 408 891
rect 402 886 408 887
rect 472 883 474 898
rect 111 882 115 883
rect 111 877 115 878
rect 343 882 347 883
rect 343 877 347 878
rect 375 882 379 883
rect 375 877 379 878
rect 431 882 435 883
rect 431 877 435 878
rect 471 882 475 883
rect 471 877 475 878
rect 535 882 539 883
rect 535 877 539 878
rect 112 853 114 877
rect 344 866 346 877
rect 410 875 416 876
rect 410 871 411 875
rect 415 871 416 875
rect 410 870 416 871
rect 342 865 348 866
rect 342 861 343 865
rect 347 861 348 865
rect 342 860 348 861
rect 110 852 116 853
rect 110 848 111 852
rect 115 848 116 852
rect 412 848 414 870
rect 432 866 434 877
rect 502 875 508 876
rect 502 871 503 875
rect 507 871 508 875
rect 502 870 508 871
rect 430 865 436 866
rect 430 861 431 865
rect 435 861 436 865
rect 430 860 436 861
rect 504 848 506 870
rect 536 866 538 877
rect 564 876 566 914
rect 582 903 588 904
rect 582 899 583 903
rect 587 899 588 903
rect 582 898 588 899
rect 710 903 716 904
rect 710 899 711 903
rect 715 899 716 903
rect 710 898 716 899
rect 854 903 860 904
rect 854 899 855 903
rect 859 899 860 903
rect 854 898 860 899
rect 1014 903 1020 904
rect 1014 899 1015 903
rect 1019 899 1020 903
rect 1014 898 1020 899
rect 584 883 586 898
rect 634 891 640 892
rect 634 887 635 891
rect 639 887 640 891
rect 634 886 640 887
rect 583 882 587 883
rect 583 877 587 878
rect 562 875 568 876
rect 562 871 563 875
rect 567 871 568 875
rect 562 870 568 871
rect 534 865 540 866
rect 534 861 535 865
rect 539 861 540 865
rect 534 860 540 861
rect 636 848 638 886
rect 712 883 714 898
rect 856 883 858 898
rect 1016 883 1018 898
rect 1168 892 1170 914
rect 1182 903 1188 904
rect 1182 899 1183 903
rect 1187 899 1188 903
rect 1182 898 1188 899
rect 1358 903 1364 904
rect 1358 899 1359 903
rect 1363 899 1364 903
rect 1534 903 1540 904
rect 1358 898 1364 899
rect 1391 900 1395 901
rect 1166 891 1172 892
rect 1166 887 1167 891
rect 1171 887 1172 891
rect 1166 886 1172 887
rect 1184 883 1186 898
rect 1360 883 1362 898
rect 1534 899 1535 903
rect 1539 899 1540 903
rect 1534 898 1540 899
rect 1391 895 1395 896
rect 1392 892 1394 895
rect 1390 891 1396 892
rect 1390 887 1391 891
rect 1395 887 1396 891
rect 1390 886 1396 887
rect 1536 883 1538 898
rect 647 882 651 883
rect 647 877 651 878
rect 711 882 715 883
rect 711 877 715 878
rect 783 882 787 883
rect 783 877 787 878
rect 855 882 859 883
rect 855 877 859 878
rect 927 882 931 883
rect 927 877 931 878
rect 1015 882 1019 883
rect 1015 877 1019 878
rect 1087 882 1091 883
rect 1087 877 1091 878
rect 1183 882 1187 883
rect 1183 877 1187 878
rect 1263 882 1267 883
rect 1263 877 1267 878
rect 1359 882 1363 883
rect 1359 877 1363 878
rect 1447 882 1451 883
rect 1447 877 1451 878
rect 1535 882 1539 883
rect 1535 877 1539 878
rect 1631 882 1635 883
rect 1631 877 1635 878
rect 648 866 650 877
rect 718 875 724 876
rect 718 871 719 875
rect 723 871 724 875
rect 718 870 724 871
rect 646 865 652 866
rect 646 861 647 865
rect 651 861 652 865
rect 646 860 652 861
rect 720 848 722 870
rect 784 866 786 877
rect 814 875 820 876
rect 814 871 815 875
rect 819 871 820 875
rect 814 870 820 871
rect 782 865 788 866
rect 782 861 783 865
rect 787 861 788 865
rect 782 860 788 861
rect 110 847 116 848
rect 410 847 416 848
rect 410 843 411 847
rect 415 843 416 847
rect 410 842 416 843
rect 502 847 508 848
rect 502 843 503 847
rect 507 843 508 847
rect 502 842 508 843
rect 634 847 640 848
rect 634 843 635 847
rect 639 843 640 847
rect 634 842 640 843
rect 718 847 724 848
rect 718 843 719 847
rect 723 843 724 847
rect 718 842 724 843
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 110 830 116 831
rect 430 835 436 836
rect 430 831 431 835
rect 435 831 436 835
rect 430 830 436 831
rect 112 815 114 830
rect 334 825 340 826
rect 334 821 335 825
rect 339 821 340 825
rect 334 820 340 821
rect 422 825 428 826
rect 422 821 423 825
rect 427 821 428 825
rect 422 820 428 821
rect 336 815 338 820
rect 424 815 426 820
rect 111 814 115 815
rect 111 809 115 810
rect 287 814 291 815
rect 287 809 291 810
rect 335 814 339 815
rect 335 809 339 810
rect 407 814 411 815
rect 407 809 411 810
rect 423 814 427 815
rect 423 809 427 810
rect 112 794 114 809
rect 288 804 290 809
rect 408 804 410 809
rect 286 803 292 804
rect 286 799 287 803
rect 291 799 292 803
rect 286 798 292 799
rect 406 803 412 804
rect 406 799 407 803
rect 411 799 412 803
rect 406 798 412 799
rect 110 793 116 794
rect 110 789 111 793
rect 115 789 116 793
rect 110 788 116 789
rect 246 779 252 780
rect 110 776 116 777
rect 110 772 111 776
rect 115 772 116 776
rect 246 775 247 779
rect 251 775 252 779
rect 246 774 252 775
rect 110 771 116 772
rect 112 743 114 771
rect 111 742 115 743
rect 111 737 115 738
rect 215 742 219 743
rect 215 737 219 738
rect 112 713 114 737
rect 216 726 218 737
rect 248 736 250 774
rect 294 763 300 764
rect 294 759 295 763
rect 299 759 300 763
rect 294 758 300 759
rect 414 763 420 764
rect 414 759 415 763
rect 419 759 420 763
rect 414 758 420 759
rect 296 743 298 758
rect 416 743 418 758
rect 432 752 434 830
rect 526 825 532 826
rect 526 821 527 825
rect 531 821 532 825
rect 526 820 532 821
rect 638 825 644 826
rect 638 821 639 825
rect 643 821 644 825
rect 638 820 644 821
rect 774 825 780 826
rect 774 821 775 825
rect 779 821 780 825
rect 774 820 780 821
rect 528 815 530 820
rect 640 815 642 820
rect 776 815 778 820
rect 527 814 531 815
rect 527 809 531 810
rect 535 814 539 815
rect 535 809 539 810
rect 639 814 643 815
rect 639 809 643 810
rect 679 814 683 815
rect 679 809 683 810
rect 775 814 779 815
rect 775 809 779 810
rect 536 804 538 809
rect 680 804 682 809
rect 534 803 540 804
rect 534 799 535 803
rect 539 799 540 803
rect 534 798 540 799
rect 678 803 684 804
rect 678 799 679 803
rect 683 799 684 803
rect 678 798 684 799
rect 816 796 818 870
rect 928 866 930 877
rect 1026 875 1032 876
rect 1026 871 1027 875
rect 1031 871 1032 875
rect 1026 870 1032 871
rect 926 865 932 866
rect 926 861 927 865
rect 931 861 932 865
rect 926 860 932 861
rect 1028 848 1030 870
rect 1088 866 1090 877
rect 1194 875 1200 876
rect 1194 871 1195 875
rect 1199 871 1200 875
rect 1194 870 1200 871
rect 1222 875 1228 876
rect 1222 871 1223 875
rect 1227 871 1228 875
rect 1222 870 1228 871
rect 1086 865 1092 866
rect 1086 861 1087 865
rect 1091 861 1092 865
rect 1086 860 1092 861
rect 1196 848 1198 870
rect 1026 847 1032 848
rect 1026 843 1027 847
rect 1031 843 1032 847
rect 1026 842 1032 843
rect 1194 847 1200 848
rect 1194 843 1195 847
rect 1199 843 1200 847
rect 1194 842 1200 843
rect 918 825 924 826
rect 918 821 919 825
rect 923 821 924 825
rect 918 820 924 821
rect 1078 825 1084 826
rect 1078 821 1079 825
rect 1083 821 1084 825
rect 1078 820 1084 821
rect 920 815 922 820
rect 1080 815 1082 820
rect 823 814 827 815
rect 823 809 827 810
rect 919 814 923 815
rect 919 809 923 810
rect 975 814 979 815
rect 975 809 979 810
rect 1079 814 1083 815
rect 1079 809 1083 810
rect 1127 814 1131 815
rect 1127 809 1131 810
rect 824 804 826 809
rect 976 804 978 809
rect 1128 804 1130 809
rect 822 803 828 804
rect 822 799 823 803
rect 827 799 828 803
rect 822 798 828 799
rect 974 803 980 804
rect 974 799 975 803
rect 979 799 980 803
rect 974 798 980 799
rect 1126 803 1132 804
rect 1126 799 1127 803
rect 1131 799 1132 803
rect 1126 798 1132 799
rect 1224 796 1226 870
rect 1264 866 1266 877
rect 1448 866 1450 877
rect 1518 875 1524 876
rect 1518 871 1519 875
rect 1523 871 1524 875
rect 1518 870 1524 871
rect 1262 865 1268 866
rect 1262 861 1263 865
rect 1267 861 1268 865
rect 1262 860 1268 861
rect 1446 865 1452 866
rect 1446 861 1447 865
rect 1451 861 1452 865
rect 1446 860 1452 861
rect 1520 848 1522 870
rect 1632 866 1634 877
rect 1660 876 1662 914
rect 1668 901 1670 914
rect 1718 903 1724 904
rect 1667 900 1671 901
rect 1718 899 1719 903
rect 1723 899 1724 903
rect 1718 898 1724 899
rect 1667 895 1671 896
rect 1720 883 1722 898
rect 1736 892 1738 974
rect 1824 955 1826 974
rect 1864 955 1866 974
rect 1934 969 1940 970
rect 1934 965 1935 969
rect 1939 965 1940 969
rect 1934 964 1940 965
rect 1936 955 1938 964
rect 1823 954 1827 955
rect 1823 949 1827 950
rect 1863 954 1867 955
rect 1863 949 1867 950
rect 1887 954 1891 955
rect 1887 949 1891 950
rect 1935 954 1939 955
rect 1935 949 1939 950
rect 1824 934 1826 949
rect 1864 934 1866 949
rect 1888 944 1890 949
rect 1886 943 1892 944
rect 1886 939 1887 943
rect 1891 939 1892 943
rect 1886 938 1892 939
rect 1822 933 1828 934
rect 1822 929 1823 933
rect 1827 929 1828 933
rect 1822 928 1828 929
rect 1862 933 1868 934
rect 1862 929 1863 933
rect 1867 929 1868 933
rect 1862 928 1868 929
rect 1822 916 1828 917
rect 1822 912 1823 916
rect 1827 912 1828 916
rect 1822 911 1828 912
rect 1862 916 1868 917
rect 1862 912 1863 916
rect 1867 912 1868 916
rect 1862 911 1868 912
rect 1734 891 1740 892
rect 1734 887 1735 891
rect 1739 887 1740 891
rect 1734 886 1740 887
rect 1824 883 1826 911
rect 1864 887 1866 911
rect 1894 903 1900 904
rect 1894 899 1895 903
rect 1899 899 1900 903
rect 1894 898 1900 899
rect 1896 887 1898 898
rect 1944 892 1946 974
rect 2062 969 2068 970
rect 2062 965 2063 969
rect 2067 965 2068 969
rect 2062 964 2068 965
rect 2064 955 2066 964
rect 2047 954 2051 955
rect 2047 949 2051 950
rect 2063 954 2067 955
rect 2063 949 2067 950
rect 2048 944 2050 949
rect 2046 943 2052 944
rect 2046 939 2047 943
rect 2051 939 2052 943
rect 2046 938 2052 939
rect 2116 936 2118 1014
rect 2192 1010 2194 1021
rect 2312 1010 2314 1021
rect 2190 1009 2196 1010
rect 2190 1005 2191 1009
rect 2195 1005 2196 1009
rect 2190 1004 2196 1005
rect 2310 1009 2316 1010
rect 2310 1005 2311 1009
rect 2315 1005 2316 1009
rect 2310 1004 2316 1005
rect 2380 980 2382 1030
rect 2416 1027 2418 1042
rect 2576 1027 2578 1042
rect 2636 1036 2638 1058
rect 2634 1035 2640 1036
rect 2634 1031 2635 1035
rect 2639 1031 2640 1035
rect 2634 1030 2640 1031
rect 2415 1026 2419 1027
rect 2415 1021 2419 1022
rect 2439 1026 2443 1027
rect 2439 1021 2443 1022
rect 2575 1026 2579 1027
rect 2575 1021 2579 1022
rect 2440 1010 2442 1021
rect 2576 1010 2578 1021
rect 2644 1020 2646 1074
rect 2978 1063 2984 1064
rect 2978 1059 2979 1063
rect 2983 1059 2984 1063
rect 2978 1058 2984 1059
rect 2742 1047 2748 1048
rect 2742 1043 2743 1047
rect 2747 1043 2748 1047
rect 2742 1042 2748 1043
rect 2918 1047 2924 1048
rect 2918 1043 2919 1047
rect 2923 1043 2924 1047
rect 2918 1042 2924 1043
rect 2744 1027 2746 1042
rect 2920 1027 2922 1042
rect 2980 1036 2982 1058
rect 3102 1047 3108 1048
rect 3102 1043 3103 1047
rect 3107 1043 3108 1047
rect 3102 1042 3108 1043
rect 2978 1035 2984 1036
rect 2978 1031 2979 1035
rect 2983 1031 2984 1035
rect 2978 1030 2984 1031
rect 3104 1027 3106 1042
rect 3144 1036 3146 1126
rect 3318 1121 3324 1122
rect 3318 1117 3319 1121
rect 3323 1117 3324 1121
rect 3318 1116 3324 1117
rect 3320 1099 3322 1116
rect 3287 1098 3291 1099
rect 3287 1093 3291 1094
rect 3319 1098 3323 1099
rect 3319 1093 3323 1094
rect 3288 1088 3290 1093
rect 3286 1087 3292 1088
rect 3286 1083 3287 1087
rect 3291 1083 3292 1087
rect 3286 1082 3292 1083
rect 3356 1080 3358 1162
rect 3388 1148 3390 1182
rect 3488 1179 3490 1194
rect 3520 1188 3522 1254
rect 3576 1251 3578 1270
rect 3575 1250 3579 1251
rect 3575 1245 3579 1246
rect 3576 1230 3578 1245
rect 3574 1229 3580 1230
rect 3574 1225 3575 1229
rect 3579 1225 3580 1229
rect 3574 1224 3580 1225
rect 3546 1215 3552 1216
rect 3546 1211 3547 1215
rect 3551 1211 3552 1215
rect 3546 1210 3552 1211
rect 3574 1212 3580 1213
rect 3518 1187 3524 1188
rect 3518 1183 3519 1187
rect 3523 1183 3524 1187
rect 3518 1182 3524 1183
rect 3487 1178 3491 1179
rect 3487 1173 3491 1174
rect 3488 1162 3490 1173
rect 3548 1172 3550 1210
rect 3574 1208 3575 1212
rect 3579 1208 3580 1212
rect 3574 1207 3580 1208
rect 3576 1179 3578 1207
rect 3575 1178 3579 1179
rect 3575 1173 3579 1174
rect 3546 1171 3552 1172
rect 3546 1167 3547 1171
rect 3551 1167 3552 1171
rect 3546 1166 3552 1167
rect 3486 1161 3492 1162
rect 3486 1157 3487 1161
rect 3491 1157 3492 1161
rect 3486 1156 3492 1157
rect 3576 1149 3578 1173
rect 3574 1148 3580 1149
rect 3386 1147 3392 1148
rect 3386 1143 3387 1147
rect 3391 1143 3392 1147
rect 3574 1144 3575 1148
rect 3579 1144 3580 1148
rect 3574 1143 3580 1144
rect 3386 1142 3392 1143
rect 3574 1131 3580 1132
rect 3574 1127 3575 1131
rect 3579 1127 3580 1131
rect 3574 1126 3580 1127
rect 3478 1121 3484 1122
rect 3478 1117 3479 1121
rect 3483 1117 3484 1121
rect 3478 1116 3484 1117
rect 3480 1099 3482 1116
rect 3518 1115 3524 1116
rect 3518 1111 3519 1115
rect 3523 1111 3524 1115
rect 3518 1110 3524 1111
rect 3479 1098 3483 1099
rect 3479 1093 3483 1094
rect 3480 1088 3482 1093
rect 3478 1087 3484 1088
rect 3478 1083 3479 1087
rect 3483 1083 3484 1087
rect 3478 1082 3484 1083
rect 3354 1079 3360 1080
rect 3354 1075 3355 1079
rect 3359 1075 3360 1079
rect 3354 1074 3360 1075
rect 3294 1047 3300 1048
rect 3294 1043 3295 1047
rect 3299 1043 3300 1047
rect 3294 1042 3300 1043
rect 3486 1047 3492 1048
rect 3486 1043 3487 1047
rect 3491 1043 3492 1047
rect 3486 1042 3492 1043
rect 3142 1035 3148 1036
rect 3142 1031 3143 1035
rect 3147 1031 3148 1035
rect 3142 1030 3148 1031
rect 3296 1027 3298 1042
rect 3488 1027 3490 1042
rect 3520 1036 3522 1110
rect 3576 1099 3578 1126
rect 3575 1098 3579 1099
rect 3575 1093 3579 1094
rect 3576 1078 3578 1093
rect 3574 1077 3580 1078
rect 3574 1073 3575 1077
rect 3579 1073 3580 1077
rect 3574 1072 3580 1073
rect 3546 1063 3552 1064
rect 3546 1059 3547 1063
rect 3551 1059 3552 1063
rect 3546 1058 3552 1059
rect 3574 1060 3580 1061
rect 3518 1035 3524 1036
rect 3518 1031 3519 1035
rect 3523 1031 3524 1035
rect 3518 1030 3524 1031
rect 2719 1026 2723 1027
rect 2719 1021 2723 1022
rect 2743 1026 2747 1027
rect 2743 1021 2747 1022
rect 2871 1026 2875 1027
rect 2871 1021 2875 1022
rect 2919 1026 2923 1027
rect 2919 1021 2923 1022
rect 3031 1026 3035 1027
rect 3031 1021 3035 1022
rect 3103 1026 3107 1027
rect 3103 1021 3107 1022
rect 3191 1026 3195 1027
rect 3191 1021 3195 1022
rect 3295 1026 3299 1027
rect 3295 1021 3299 1022
rect 3351 1026 3355 1027
rect 3351 1021 3355 1022
rect 3487 1026 3491 1027
rect 3487 1021 3491 1022
rect 2642 1019 2648 1020
rect 2642 1015 2643 1019
rect 2647 1015 2648 1019
rect 2642 1014 2648 1015
rect 2720 1010 2722 1021
rect 2872 1010 2874 1021
rect 3032 1010 3034 1021
rect 3192 1010 3194 1021
rect 3352 1010 3354 1021
rect 3418 1019 3424 1020
rect 3418 1015 3419 1019
rect 3423 1015 3424 1019
rect 3418 1014 3424 1015
rect 2438 1009 2444 1010
rect 2438 1005 2439 1009
rect 2443 1005 2444 1009
rect 2438 1004 2444 1005
rect 2574 1009 2580 1010
rect 2574 1005 2575 1009
rect 2579 1005 2580 1009
rect 2574 1004 2580 1005
rect 2718 1009 2724 1010
rect 2718 1005 2719 1009
rect 2723 1005 2724 1009
rect 2718 1004 2724 1005
rect 2870 1009 2876 1010
rect 2870 1005 2871 1009
rect 2875 1005 2876 1009
rect 2870 1004 2876 1005
rect 3030 1009 3036 1010
rect 3030 1005 3031 1009
rect 3035 1005 3036 1009
rect 3030 1004 3036 1005
rect 3190 1009 3196 1010
rect 3190 1005 3191 1009
rect 3195 1005 3196 1009
rect 3190 1004 3196 1005
rect 3350 1009 3356 1010
rect 3350 1005 3351 1009
rect 3355 1005 3356 1009
rect 3350 1004 3356 1005
rect 3420 992 3422 1014
rect 3488 1010 3490 1021
rect 3548 1020 3550 1058
rect 3574 1056 3575 1060
rect 3579 1056 3580 1060
rect 3574 1055 3580 1056
rect 3576 1027 3578 1055
rect 3575 1026 3579 1027
rect 3575 1021 3579 1022
rect 3546 1019 3552 1020
rect 3546 1015 3547 1019
rect 3551 1015 3552 1019
rect 3546 1014 3552 1015
rect 3486 1009 3492 1010
rect 3486 1005 3487 1009
rect 3491 1005 3492 1009
rect 3486 1004 3492 1005
rect 3576 997 3578 1021
rect 3574 996 3580 997
rect 3574 992 3575 996
rect 3579 992 3580 996
rect 3418 991 3424 992
rect 3574 991 3580 992
rect 3418 987 3419 991
rect 3423 987 3424 991
rect 3418 986 3424 987
rect 2378 979 2384 980
rect 2378 975 2379 979
rect 2383 975 2384 979
rect 2378 974 2384 975
rect 2958 979 2964 980
rect 2958 975 2959 979
rect 2963 975 2964 979
rect 2958 974 2964 975
rect 3574 979 3580 980
rect 3574 975 3575 979
rect 3579 975 3580 979
rect 3574 974 3580 975
rect 2182 969 2188 970
rect 2182 965 2183 969
rect 2187 965 2188 969
rect 2182 964 2188 965
rect 2302 969 2308 970
rect 2302 965 2303 969
rect 2307 965 2308 969
rect 2302 964 2308 965
rect 2430 969 2436 970
rect 2430 965 2431 969
rect 2435 965 2436 969
rect 2430 964 2436 965
rect 2566 969 2572 970
rect 2566 965 2567 969
rect 2571 965 2572 969
rect 2566 964 2572 965
rect 2710 969 2716 970
rect 2710 965 2711 969
rect 2715 965 2716 969
rect 2710 964 2716 965
rect 2862 969 2868 970
rect 2862 965 2863 969
rect 2867 965 2868 969
rect 2862 964 2868 965
rect 2184 955 2186 964
rect 2304 955 2306 964
rect 2432 955 2434 964
rect 2534 955 2540 956
rect 2568 955 2570 964
rect 2712 955 2714 964
rect 2864 955 2866 964
rect 2960 956 2962 974
rect 3022 969 3028 970
rect 3022 965 3023 969
rect 3027 965 3028 969
rect 3022 964 3028 965
rect 3182 969 3188 970
rect 3182 965 3183 969
rect 3187 965 3188 969
rect 3182 964 3188 965
rect 3342 969 3348 970
rect 3342 965 3343 969
rect 3347 965 3348 969
rect 3342 964 3348 965
rect 3478 969 3484 970
rect 3478 965 3479 969
rect 3483 965 3484 969
rect 3478 964 3484 965
rect 2958 955 2964 956
rect 3024 955 3026 964
rect 3184 955 3186 964
rect 3344 955 3346 964
rect 3480 955 3482 964
rect 3576 955 3578 974
rect 2183 954 2187 955
rect 2183 949 2187 950
rect 2199 954 2203 955
rect 2199 949 2203 950
rect 2303 954 2307 955
rect 2303 949 2307 950
rect 2351 954 2355 955
rect 2351 949 2355 950
rect 2431 954 2435 955
rect 2431 949 2435 950
rect 2495 954 2499 955
rect 2534 951 2535 955
rect 2539 951 2540 955
rect 2534 950 2540 951
rect 2567 954 2571 955
rect 2495 949 2499 950
rect 2200 944 2202 949
rect 2352 944 2354 949
rect 2496 944 2498 949
rect 2198 943 2204 944
rect 2198 939 2199 943
rect 2203 939 2204 943
rect 2198 938 2204 939
rect 2350 943 2356 944
rect 2350 939 2351 943
rect 2355 939 2356 943
rect 2350 938 2356 939
rect 2494 943 2500 944
rect 2494 939 2495 943
rect 2499 939 2500 943
rect 2494 938 2500 939
rect 2114 935 2120 936
rect 2114 931 2115 935
rect 2119 931 2120 935
rect 2114 930 2120 931
rect 2038 919 2044 920
rect 2038 915 2039 919
rect 2043 915 2044 919
rect 2038 914 2044 915
rect 2266 919 2272 920
rect 2266 915 2267 919
rect 2271 915 2272 919
rect 2266 914 2272 915
rect 1942 891 1948 892
rect 1942 887 1943 891
rect 1947 887 1948 891
rect 1863 886 1867 887
rect 1719 882 1723 883
rect 1719 877 1723 878
rect 1823 882 1827 883
rect 1863 881 1867 882
rect 1895 886 1899 887
rect 1942 886 1948 887
rect 2015 886 2019 887
rect 1895 881 1899 882
rect 2015 881 2019 882
rect 1823 877 1827 878
rect 1658 875 1664 876
rect 1658 871 1659 875
rect 1663 871 1664 875
rect 1658 870 1664 871
rect 1630 865 1636 866
rect 1630 861 1631 865
rect 1635 861 1636 865
rect 1630 860 1636 861
rect 1824 853 1826 877
rect 1864 857 1866 881
rect 1896 870 1898 881
rect 1966 879 1972 880
rect 1966 875 1967 879
rect 1971 875 1972 879
rect 1966 874 1972 875
rect 1894 869 1900 870
rect 1894 865 1895 869
rect 1899 865 1900 869
rect 1894 864 1900 865
rect 1862 856 1868 857
rect 1822 852 1828 853
rect 1822 848 1823 852
rect 1827 848 1828 852
rect 1862 852 1863 856
rect 1867 852 1868 856
rect 1968 852 1970 874
rect 2016 870 2018 881
rect 2040 880 2042 914
rect 2054 903 2060 904
rect 2054 899 2055 903
rect 2059 899 2060 903
rect 2054 898 2060 899
rect 2206 903 2212 904
rect 2206 899 2207 903
rect 2211 899 2212 903
rect 2206 898 2212 899
rect 2056 887 2058 898
rect 2208 887 2210 898
rect 2268 892 2270 914
rect 2358 903 2364 904
rect 2358 899 2359 903
rect 2363 899 2364 903
rect 2358 898 2364 899
rect 2502 903 2508 904
rect 2502 899 2503 903
rect 2507 899 2508 903
rect 2502 898 2508 899
rect 2266 891 2272 892
rect 2266 887 2267 891
rect 2271 887 2272 891
rect 2360 887 2362 898
rect 2390 891 2396 892
rect 2390 887 2391 891
rect 2395 887 2396 891
rect 2504 887 2506 898
rect 2536 892 2538 950
rect 2567 949 2571 950
rect 2631 954 2635 955
rect 2631 949 2635 950
rect 2711 954 2715 955
rect 2711 949 2715 950
rect 2759 954 2763 955
rect 2759 949 2763 950
rect 2863 954 2867 955
rect 2863 949 2867 950
rect 2887 954 2891 955
rect 2958 951 2959 955
rect 2963 951 2964 955
rect 2958 950 2964 951
rect 3023 954 3027 955
rect 2887 949 2891 950
rect 3023 949 3027 950
rect 3183 954 3187 955
rect 3183 949 3187 950
rect 3343 954 3347 955
rect 3343 949 3347 950
rect 3479 954 3483 955
rect 3479 949 3483 950
rect 3575 954 3579 955
rect 3575 949 3579 950
rect 2632 944 2634 949
rect 2760 944 2762 949
rect 2888 944 2890 949
rect 3024 944 3026 949
rect 2630 943 2636 944
rect 2630 939 2631 943
rect 2635 939 2636 943
rect 2630 938 2636 939
rect 2758 943 2764 944
rect 2758 939 2759 943
rect 2763 939 2764 943
rect 2758 938 2764 939
rect 2886 943 2892 944
rect 2886 939 2887 943
rect 2891 939 2892 943
rect 2886 938 2892 939
rect 3022 943 3028 944
rect 3022 939 3023 943
rect 3027 939 3028 943
rect 3022 938 3028 939
rect 3576 934 3578 949
rect 3574 933 3580 934
rect 3574 929 3575 933
rect 3579 929 3580 933
rect 3574 928 3580 929
rect 2714 919 2720 920
rect 2714 915 2715 919
rect 2719 915 2720 919
rect 2714 914 2720 915
rect 2854 919 2860 920
rect 2854 915 2855 919
rect 2859 915 2860 919
rect 2854 914 2860 915
rect 3090 919 3096 920
rect 3090 915 3091 919
rect 3095 915 3096 919
rect 3090 914 3096 915
rect 3574 916 3580 917
rect 2638 903 2644 904
rect 2638 899 2639 903
rect 2643 899 2644 903
rect 2638 898 2644 899
rect 2534 891 2540 892
rect 2534 887 2535 891
rect 2539 887 2540 891
rect 2640 887 2642 898
rect 2716 892 2718 914
rect 2766 903 2772 904
rect 2766 899 2767 903
rect 2771 899 2772 903
rect 2766 898 2772 899
rect 2714 891 2720 892
rect 2714 887 2715 891
rect 2719 887 2720 891
rect 2768 887 2770 898
rect 2856 892 2858 914
rect 2894 903 2900 904
rect 2894 899 2895 903
rect 2899 899 2900 903
rect 2894 898 2900 899
rect 3030 903 3036 904
rect 3030 899 3031 903
rect 3035 899 3036 903
rect 3030 898 3036 899
rect 2854 891 2860 892
rect 2854 887 2855 891
rect 2859 887 2860 891
rect 2896 887 2898 898
rect 3032 887 3034 898
rect 2055 886 2059 887
rect 2055 881 2059 882
rect 2167 886 2171 887
rect 2167 881 2171 882
rect 2207 886 2211 887
rect 2266 886 2272 887
rect 2319 886 2323 887
rect 2207 881 2211 882
rect 2319 881 2323 882
rect 2359 886 2363 887
rect 2390 886 2396 887
rect 2487 886 2491 887
rect 2359 881 2363 882
rect 2038 879 2044 880
rect 2038 875 2039 879
rect 2043 875 2044 879
rect 2038 874 2044 875
rect 2168 870 2170 881
rect 2206 875 2212 876
rect 2206 871 2207 875
rect 2211 871 2212 875
rect 2206 870 2212 871
rect 2320 870 2322 881
rect 2382 879 2388 880
rect 2382 875 2383 879
rect 2387 875 2388 879
rect 2382 874 2388 875
rect 2014 869 2020 870
rect 2014 865 2015 869
rect 2019 865 2020 869
rect 2014 864 2020 865
rect 2166 869 2172 870
rect 2166 865 2167 869
rect 2171 865 2172 869
rect 2166 864 2172 865
rect 1862 851 1868 852
rect 1966 851 1972 852
rect 1518 847 1524 848
rect 1822 847 1828 848
rect 1966 847 1967 851
rect 1971 847 1972 851
rect 1518 843 1519 847
rect 1523 843 1524 847
rect 1966 846 1972 847
rect 1518 842 1524 843
rect 1862 839 1868 840
rect 1822 835 1828 836
rect 1822 831 1823 835
rect 1827 831 1828 835
rect 1862 835 1863 839
rect 1867 835 1868 839
rect 1862 834 1868 835
rect 1822 830 1828 831
rect 1254 825 1260 826
rect 1254 821 1255 825
rect 1259 821 1260 825
rect 1254 820 1260 821
rect 1438 825 1444 826
rect 1438 821 1439 825
rect 1443 821 1444 825
rect 1438 820 1444 821
rect 1622 825 1628 826
rect 1622 821 1623 825
rect 1627 821 1628 825
rect 1622 820 1628 821
rect 1256 815 1258 820
rect 1440 815 1442 820
rect 1478 819 1484 820
rect 1478 815 1479 819
rect 1483 815 1484 819
rect 1624 815 1626 820
rect 1824 815 1826 830
rect 1864 819 1866 834
rect 1886 829 1892 830
rect 1886 825 1887 829
rect 1891 825 1892 829
rect 1886 824 1892 825
rect 2006 829 2012 830
rect 2006 825 2007 829
rect 2011 825 2012 829
rect 2006 824 2012 825
rect 2158 829 2164 830
rect 2158 825 2159 829
rect 2163 825 2164 829
rect 2158 824 2164 825
rect 1888 819 1890 824
rect 1926 823 1932 824
rect 1926 819 1927 823
rect 1931 819 1932 823
rect 2008 819 2010 824
rect 2160 819 2162 824
rect 1863 818 1867 819
rect 1255 814 1259 815
rect 1255 809 1259 810
rect 1279 814 1283 815
rect 1279 809 1283 810
rect 1439 814 1443 815
rect 1478 814 1484 815
rect 1599 814 1603 815
rect 1439 809 1443 810
rect 1280 804 1282 809
rect 1440 804 1442 809
rect 1278 803 1284 804
rect 1278 799 1279 803
rect 1283 799 1284 803
rect 1278 798 1284 799
rect 1438 803 1444 804
rect 1438 799 1439 803
rect 1443 799 1444 803
rect 1438 798 1444 799
rect 474 795 480 796
rect 474 791 475 795
rect 479 791 480 795
rect 474 790 480 791
rect 814 795 820 796
rect 814 791 815 795
rect 819 791 820 795
rect 814 790 820 791
rect 1222 795 1228 796
rect 1222 791 1223 795
rect 1227 791 1228 795
rect 1222 790 1228 791
rect 476 760 478 790
rect 542 763 548 764
rect 474 759 480 760
rect 474 755 475 759
rect 479 755 480 759
rect 542 759 543 763
rect 547 759 548 763
rect 542 758 548 759
rect 686 763 692 764
rect 686 759 687 763
rect 691 759 692 763
rect 686 758 692 759
rect 830 763 836 764
rect 830 759 831 763
rect 835 759 836 763
rect 830 758 836 759
rect 982 763 988 764
rect 982 759 983 763
rect 987 759 988 763
rect 982 758 988 759
rect 1134 763 1140 764
rect 1134 759 1135 763
rect 1139 759 1140 763
rect 1134 758 1140 759
rect 1286 763 1292 764
rect 1286 759 1287 763
rect 1291 759 1292 763
rect 1286 758 1292 759
rect 1446 763 1452 764
rect 1446 759 1447 763
rect 1451 759 1452 763
rect 1446 758 1452 759
rect 474 754 480 755
rect 430 751 436 752
rect 430 747 431 751
rect 435 747 436 751
rect 430 746 436 747
rect 544 743 546 758
rect 688 743 690 758
rect 706 751 712 752
rect 706 747 707 751
rect 711 747 712 751
rect 706 746 712 747
rect 295 742 299 743
rect 295 737 299 738
rect 359 742 363 743
rect 359 737 363 738
rect 415 742 419 743
rect 415 737 419 738
rect 503 742 507 743
rect 503 737 507 738
rect 543 742 547 743
rect 543 737 547 738
rect 647 742 651 743
rect 647 737 651 738
rect 687 742 691 743
rect 687 737 691 738
rect 246 735 252 736
rect 246 731 247 735
rect 251 731 252 735
rect 246 730 252 731
rect 326 735 332 736
rect 326 731 327 735
rect 331 731 332 735
rect 326 730 332 731
rect 214 725 220 726
rect 214 721 215 725
rect 219 721 220 725
rect 214 720 220 721
rect 110 712 116 713
rect 328 712 330 730
rect 360 726 362 737
rect 504 726 506 737
rect 648 726 650 737
rect 358 725 364 726
rect 358 721 359 725
rect 363 721 364 725
rect 358 720 364 721
rect 502 725 508 726
rect 502 721 503 725
rect 507 721 508 725
rect 502 720 508 721
rect 646 725 652 726
rect 646 721 647 725
rect 651 721 652 725
rect 646 720 652 721
rect 708 712 710 746
rect 832 743 834 758
rect 984 743 986 758
rect 1136 743 1138 758
rect 1162 743 1168 744
rect 1288 743 1290 758
rect 1315 756 1319 757
rect 1314 751 1320 752
rect 1314 747 1315 751
rect 1319 747 1320 751
rect 1314 746 1320 747
rect 1448 743 1450 758
rect 1480 752 1482 814
rect 1599 809 1603 810
rect 1623 814 1627 815
rect 1623 809 1627 810
rect 1823 814 1827 815
rect 1863 813 1867 814
rect 1887 818 1891 819
rect 1926 818 1932 819
rect 1991 818 1995 819
rect 1887 813 1891 814
rect 1823 809 1827 810
rect 1600 804 1602 809
rect 1598 803 1604 804
rect 1598 799 1599 803
rect 1603 799 1604 803
rect 1598 798 1604 799
rect 1518 795 1524 796
rect 1518 791 1519 795
rect 1523 791 1524 795
rect 1824 794 1826 809
rect 1864 798 1866 813
rect 1888 808 1890 813
rect 1886 807 1892 808
rect 1886 803 1887 807
rect 1891 803 1892 807
rect 1886 802 1892 803
rect 1862 797 1868 798
rect 1518 790 1524 791
rect 1822 793 1828 794
rect 1520 757 1522 790
rect 1822 789 1823 793
rect 1827 789 1828 793
rect 1862 793 1863 797
rect 1867 793 1868 797
rect 1862 792 1868 793
rect 1822 788 1828 789
rect 1862 780 1868 781
rect 1822 776 1828 777
rect 1822 772 1823 776
rect 1827 772 1828 776
rect 1862 776 1863 780
rect 1867 776 1868 780
rect 1862 775 1868 776
rect 1822 771 1828 772
rect 1606 763 1612 764
rect 1606 759 1607 763
rect 1611 759 1612 763
rect 1606 758 1612 759
rect 1519 756 1523 757
rect 1478 751 1484 752
rect 1519 751 1523 752
rect 1478 747 1479 751
rect 1483 747 1484 751
rect 1478 746 1484 747
rect 1608 743 1610 758
rect 1824 743 1826 771
rect 1864 747 1866 775
rect 1894 767 1900 768
rect 1894 763 1895 767
rect 1899 763 1900 767
rect 1894 762 1900 763
rect 1896 747 1898 762
rect 1928 756 1930 818
rect 1991 813 1995 814
rect 2007 818 2011 819
rect 2007 813 2011 814
rect 2135 818 2139 819
rect 2135 813 2139 814
rect 2159 818 2163 819
rect 2159 813 2163 814
rect 1992 808 1994 813
rect 2136 808 2138 813
rect 1990 807 1996 808
rect 1990 803 1991 807
rect 1995 803 1996 807
rect 1990 802 1996 803
rect 2134 807 2140 808
rect 2134 803 2135 807
rect 2139 803 2140 807
rect 2134 802 2140 803
rect 2208 800 2210 870
rect 2318 869 2324 870
rect 2318 865 2319 869
rect 2323 865 2324 869
rect 2318 864 2324 865
rect 2384 856 2386 874
rect 2382 855 2388 856
rect 2382 851 2383 855
rect 2387 851 2388 855
rect 2392 852 2394 886
rect 2487 881 2491 882
rect 2503 886 2507 887
rect 2534 886 2540 887
rect 2639 886 2643 887
rect 2503 881 2507 882
rect 2639 881 2643 882
rect 2663 886 2667 887
rect 2714 886 2720 887
rect 2767 886 2771 887
rect 2663 881 2667 882
rect 2767 881 2771 882
rect 2847 886 2851 887
rect 2854 886 2860 887
rect 2895 886 2899 887
rect 2847 881 2851 882
rect 2895 881 2899 882
rect 3031 886 3035 887
rect 3031 881 3035 882
rect 3039 886 3043 887
rect 3039 881 3043 882
rect 2488 870 2490 881
rect 2664 870 2666 881
rect 2848 870 2850 881
rect 2878 879 2884 880
rect 2878 875 2879 879
rect 2883 875 2884 879
rect 2878 874 2884 875
rect 2486 869 2492 870
rect 2486 865 2487 869
rect 2491 865 2492 869
rect 2486 864 2492 865
rect 2662 869 2668 870
rect 2662 865 2663 869
rect 2667 865 2668 869
rect 2662 864 2668 865
rect 2846 869 2852 870
rect 2846 865 2847 869
rect 2851 865 2852 869
rect 2846 864 2852 865
rect 2382 850 2388 851
rect 2390 851 2396 852
rect 2390 847 2391 851
rect 2395 847 2396 851
rect 2390 846 2396 847
rect 2662 839 2668 840
rect 2662 835 2663 839
rect 2667 835 2668 839
rect 2662 834 2668 835
rect 2310 829 2316 830
rect 2310 825 2311 829
rect 2315 825 2316 829
rect 2310 824 2316 825
rect 2478 829 2484 830
rect 2478 825 2479 829
rect 2483 825 2484 829
rect 2478 824 2484 825
rect 2654 829 2660 830
rect 2654 825 2655 829
rect 2659 825 2660 829
rect 2654 824 2660 825
rect 2312 819 2314 824
rect 2480 819 2482 824
rect 2656 819 2658 824
rect 2287 818 2291 819
rect 2287 813 2291 814
rect 2311 818 2315 819
rect 2311 813 2315 814
rect 2455 818 2459 819
rect 2455 813 2459 814
rect 2479 818 2483 819
rect 2479 813 2483 814
rect 2623 818 2627 819
rect 2623 813 2627 814
rect 2655 818 2659 819
rect 2655 813 2659 814
rect 2288 808 2290 813
rect 2456 808 2458 813
rect 2624 808 2626 813
rect 2286 807 2292 808
rect 2286 803 2287 807
rect 2291 803 2292 807
rect 2286 802 2292 803
rect 2454 807 2460 808
rect 2454 803 2455 807
rect 2459 803 2460 807
rect 2454 802 2460 803
rect 2622 807 2628 808
rect 2622 803 2623 807
rect 2627 803 2628 807
rect 2622 802 2628 803
rect 2206 799 2212 800
rect 2206 795 2207 799
rect 2211 795 2212 799
rect 2206 794 2212 795
rect 1954 783 1960 784
rect 1954 779 1955 783
rect 1959 779 1960 783
rect 1954 778 1960 779
rect 2202 783 2208 784
rect 2202 779 2203 783
rect 2207 779 2208 783
rect 2202 778 2208 779
rect 2354 783 2360 784
rect 2354 779 2355 783
rect 2359 779 2360 783
rect 2354 778 2360 779
rect 1926 755 1932 756
rect 1926 751 1927 755
rect 1931 751 1932 755
rect 1926 750 1932 751
rect 1863 746 1867 747
rect 791 742 795 743
rect 791 737 795 738
rect 831 742 835 743
rect 831 737 835 738
rect 935 742 939 743
rect 935 737 939 738
rect 983 742 987 743
rect 983 737 987 738
rect 1087 742 1091 743
rect 1087 737 1091 738
rect 1135 742 1139 743
rect 1162 739 1163 743
rect 1167 739 1168 743
rect 1162 738 1168 739
rect 1247 742 1251 743
rect 1135 737 1139 738
rect 738 735 744 736
rect 738 731 739 735
rect 743 731 744 735
rect 738 730 744 731
rect 110 708 111 712
rect 115 708 116 712
rect 110 707 116 708
rect 326 711 332 712
rect 326 707 327 711
rect 331 707 332 711
rect 326 706 332 707
rect 706 711 712 712
rect 706 707 707 711
rect 711 707 712 711
rect 740 708 742 730
rect 792 726 794 737
rect 842 735 848 736
rect 842 731 843 735
rect 847 731 848 735
rect 842 730 848 731
rect 790 725 796 726
rect 790 721 791 725
rect 795 721 796 725
rect 790 720 796 721
rect 706 706 712 707
rect 738 707 744 708
rect 738 703 739 707
rect 743 703 744 707
rect 738 702 744 703
rect 110 695 116 696
rect 110 691 111 695
rect 115 691 116 695
rect 110 690 116 691
rect 502 695 508 696
rect 502 691 503 695
rect 507 691 508 695
rect 502 690 508 691
rect 112 675 114 690
rect 206 685 212 686
rect 206 681 207 685
rect 211 681 212 685
rect 206 680 212 681
rect 350 685 356 686
rect 350 681 351 685
rect 355 681 356 685
rect 350 680 356 681
rect 494 685 500 686
rect 494 681 495 685
rect 499 681 500 685
rect 494 680 500 681
rect 208 675 210 680
rect 352 675 354 680
rect 496 675 498 680
rect 111 674 115 675
rect 111 669 115 670
rect 135 674 139 675
rect 135 669 139 670
rect 207 674 211 675
rect 207 669 211 670
rect 295 674 299 675
rect 295 669 299 670
rect 351 674 355 675
rect 351 669 355 670
rect 463 674 467 675
rect 463 669 467 670
rect 495 674 499 675
rect 495 669 499 670
rect 112 654 114 669
rect 136 664 138 669
rect 296 664 298 669
rect 464 664 466 669
rect 134 663 140 664
rect 134 659 135 663
rect 139 659 140 663
rect 134 658 140 659
rect 294 663 300 664
rect 294 659 295 663
rect 299 659 300 663
rect 294 658 300 659
rect 462 663 468 664
rect 462 659 463 663
rect 467 659 468 663
rect 462 658 468 659
rect 110 653 116 654
rect 110 649 111 653
rect 115 649 116 653
rect 110 648 116 649
rect 202 639 208 640
rect 110 636 116 637
rect 110 632 111 636
rect 115 632 116 636
rect 202 635 203 639
rect 207 635 208 639
rect 202 634 208 635
rect 362 639 368 640
rect 362 635 363 639
rect 367 635 368 639
rect 362 634 368 635
rect 110 631 116 632
rect 112 603 114 631
rect 142 623 148 624
rect 142 619 143 623
rect 147 619 148 623
rect 142 618 148 619
rect 144 603 146 618
rect 204 612 206 634
rect 302 623 308 624
rect 302 619 303 623
rect 307 619 308 623
rect 302 618 308 619
rect 202 611 208 612
rect 202 607 203 611
rect 207 607 208 611
rect 202 606 208 607
rect 304 603 306 618
rect 364 612 366 634
rect 470 623 476 624
rect 470 619 471 623
rect 475 619 476 623
rect 470 618 476 619
rect 362 611 368 612
rect 362 607 363 611
rect 367 607 368 611
rect 362 606 368 607
rect 472 603 474 618
rect 504 612 506 690
rect 638 685 644 686
rect 638 681 639 685
rect 643 681 644 685
rect 638 680 644 681
rect 782 685 788 686
rect 782 681 783 685
rect 787 681 788 685
rect 782 680 788 681
rect 640 675 642 680
rect 784 675 786 680
rect 623 674 627 675
rect 623 669 627 670
rect 639 674 643 675
rect 639 669 643 670
rect 775 674 779 675
rect 775 669 779 670
rect 783 674 787 675
rect 783 669 787 670
rect 624 664 626 669
rect 776 664 778 669
rect 622 663 628 664
rect 622 659 623 663
rect 627 659 628 663
rect 622 658 628 659
rect 774 663 780 664
rect 774 659 775 663
rect 779 659 780 663
rect 774 658 780 659
rect 844 656 846 730
rect 936 726 938 737
rect 1088 726 1090 737
rect 1142 735 1148 736
rect 1142 731 1143 735
rect 1147 731 1148 735
rect 1142 730 1148 731
rect 934 725 940 726
rect 934 721 935 725
rect 939 721 940 725
rect 934 720 940 721
rect 1086 725 1092 726
rect 1086 721 1087 725
rect 1091 721 1092 725
rect 1086 720 1092 721
rect 926 685 932 686
rect 926 681 927 685
rect 931 681 932 685
rect 926 680 932 681
rect 1078 685 1084 686
rect 1078 681 1079 685
rect 1083 681 1084 685
rect 1078 680 1084 681
rect 928 675 930 680
rect 1080 675 1082 680
rect 927 674 931 675
rect 927 669 931 670
rect 1071 674 1075 675
rect 1071 669 1075 670
rect 1079 674 1083 675
rect 1079 669 1083 670
rect 928 664 930 669
rect 1072 664 1074 669
rect 926 663 932 664
rect 926 659 927 663
rect 931 659 932 663
rect 926 658 932 659
rect 1070 663 1076 664
rect 1070 659 1071 663
rect 1075 659 1076 663
rect 1070 658 1076 659
rect 1144 656 1146 730
rect 1164 696 1166 738
rect 1247 737 1251 738
rect 1287 742 1291 743
rect 1287 737 1291 738
rect 1415 742 1419 743
rect 1415 737 1419 738
rect 1447 742 1451 743
rect 1447 737 1451 738
rect 1583 742 1587 743
rect 1583 737 1587 738
rect 1607 742 1611 743
rect 1607 737 1611 738
rect 1735 742 1739 743
rect 1735 737 1739 738
rect 1823 742 1827 743
rect 1863 741 1867 742
rect 1895 746 1899 747
rect 1895 741 1899 742
rect 1823 737 1827 738
rect 1248 726 1250 737
rect 1416 726 1418 737
rect 1584 726 1586 737
rect 1736 726 1738 737
rect 1246 725 1252 726
rect 1246 721 1247 725
rect 1251 721 1252 725
rect 1246 720 1252 721
rect 1414 725 1420 726
rect 1414 721 1415 725
rect 1419 721 1420 725
rect 1414 720 1420 721
rect 1582 725 1588 726
rect 1582 721 1583 725
rect 1587 721 1588 725
rect 1582 720 1588 721
rect 1734 725 1740 726
rect 1734 721 1735 725
rect 1739 721 1740 725
rect 1734 720 1740 721
rect 1824 713 1826 737
rect 1864 717 1866 741
rect 1870 735 1876 736
rect 1870 731 1871 735
rect 1875 731 1876 735
rect 1870 730 1876 731
rect 1896 730 1898 741
rect 1956 740 1958 778
rect 1998 767 2004 768
rect 1998 763 1999 767
rect 2003 763 2004 767
rect 1998 762 2004 763
rect 2142 767 2148 768
rect 2142 763 2143 767
rect 2147 763 2148 767
rect 2142 762 2148 763
rect 2000 747 2002 762
rect 2144 747 2146 762
rect 2204 748 2206 778
rect 2294 767 2300 768
rect 2294 763 2295 767
rect 2299 763 2300 767
rect 2294 762 2300 763
rect 2202 747 2208 748
rect 2296 747 2298 762
rect 2356 756 2358 778
rect 2462 767 2468 768
rect 2462 763 2463 767
rect 2467 763 2468 767
rect 2462 762 2468 763
rect 2630 767 2636 768
rect 2630 763 2631 767
rect 2635 763 2636 767
rect 2630 762 2636 763
rect 2354 755 2360 756
rect 2354 751 2355 755
rect 2359 751 2360 755
rect 2354 750 2360 751
rect 2464 747 2466 762
rect 2506 755 2512 756
rect 2506 751 2507 755
rect 2511 751 2512 755
rect 2506 750 2512 751
rect 1999 746 2003 747
rect 1999 741 2003 742
rect 2063 746 2067 747
rect 2063 741 2067 742
rect 2143 746 2147 747
rect 2202 743 2203 747
rect 2207 743 2208 747
rect 2202 742 2208 743
rect 2255 746 2259 747
rect 2143 741 2147 742
rect 2255 741 2259 742
rect 2295 746 2299 747
rect 2295 741 2299 742
rect 2447 746 2451 747
rect 2447 741 2451 742
rect 2463 746 2467 747
rect 2463 741 2467 742
rect 1954 739 1960 740
rect 1954 735 1955 739
rect 1959 735 1960 739
rect 1954 734 1960 735
rect 2064 730 2066 741
rect 2094 739 2100 740
rect 2094 735 2095 739
rect 2099 735 2100 739
rect 2094 734 2100 735
rect 1862 716 1868 717
rect 1822 712 1828 713
rect 1822 708 1823 712
rect 1827 708 1828 712
rect 1862 712 1863 716
rect 1867 712 1868 716
rect 1872 712 1874 730
rect 1894 729 1900 730
rect 1894 725 1895 729
rect 1899 725 1900 729
rect 1894 724 1900 725
rect 2062 729 2068 730
rect 2062 725 2063 729
rect 2067 725 2068 729
rect 2062 724 2068 725
rect 1862 711 1868 712
rect 1870 711 1876 712
rect 1822 707 1828 708
rect 1870 707 1871 711
rect 1875 707 1876 711
rect 1870 706 1876 707
rect 1862 699 1868 700
rect 1162 695 1168 696
rect 1162 691 1163 695
rect 1167 691 1168 695
rect 1162 690 1168 691
rect 1518 695 1524 696
rect 1518 691 1519 695
rect 1523 691 1524 695
rect 1518 690 1524 691
rect 1822 695 1828 696
rect 1822 691 1823 695
rect 1827 691 1828 695
rect 1862 695 1863 699
rect 1867 695 1868 699
rect 1862 694 1868 695
rect 1822 690 1828 691
rect 1238 685 1244 686
rect 1238 681 1239 685
rect 1243 681 1244 685
rect 1238 680 1244 681
rect 1406 685 1412 686
rect 1406 681 1407 685
rect 1411 681 1412 685
rect 1406 680 1412 681
rect 1240 675 1242 680
rect 1408 675 1410 680
rect 1207 674 1211 675
rect 1207 669 1211 670
rect 1239 674 1243 675
rect 1239 669 1243 670
rect 1343 674 1347 675
rect 1343 669 1347 670
rect 1407 674 1411 675
rect 1407 669 1411 670
rect 1479 674 1483 675
rect 1479 669 1483 670
rect 1208 664 1210 669
rect 1344 664 1346 669
rect 1480 664 1482 669
rect 1206 663 1212 664
rect 1206 659 1207 663
rect 1211 659 1212 663
rect 1206 658 1212 659
rect 1342 663 1348 664
rect 1342 659 1343 663
rect 1347 659 1348 663
rect 1342 658 1348 659
rect 1478 663 1484 664
rect 1478 659 1479 663
rect 1483 659 1484 663
rect 1478 658 1484 659
rect 842 655 848 656
rect 842 651 843 655
rect 847 651 848 655
rect 842 650 848 651
rect 1142 655 1148 656
rect 1142 651 1143 655
rect 1147 651 1148 655
rect 1142 650 1148 651
rect 1410 639 1416 640
rect 1410 635 1411 639
rect 1415 635 1416 639
rect 1410 634 1416 635
rect 1418 639 1424 640
rect 1418 635 1419 639
rect 1423 635 1424 639
rect 1418 634 1424 635
rect 630 623 636 624
rect 630 619 631 623
rect 635 619 636 623
rect 630 618 636 619
rect 782 623 788 624
rect 782 619 783 623
rect 787 619 788 623
rect 782 618 788 619
rect 934 623 940 624
rect 934 619 935 623
rect 939 619 940 623
rect 934 618 940 619
rect 1078 623 1084 624
rect 1078 619 1079 623
rect 1083 619 1084 623
rect 1078 618 1084 619
rect 1214 623 1220 624
rect 1214 619 1215 623
rect 1219 619 1220 623
rect 1214 618 1220 619
rect 1350 623 1356 624
rect 1350 619 1351 623
rect 1355 619 1356 623
rect 1350 618 1356 619
rect 502 611 508 612
rect 502 607 503 611
rect 507 607 508 611
rect 502 606 508 607
rect 632 603 634 618
rect 662 611 668 612
rect 662 607 663 611
rect 667 607 668 611
rect 662 606 668 607
rect 111 602 115 603
rect 111 597 115 598
rect 143 602 147 603
rect 143 597 147 598
rect 303 602 307 603
rect 303 597 307 598
rect 471 602 475 603
rect 471 597 475 598
rect 487 602 491 603
rect 487 597 491 598
rect 631 602 635 603
rect 631 597 635 598
rect 112 573 114 597
rect 144 586 146 597
rect 304 586 306 597
rect 488 586 490 597
rect 142 585 148 586
rect 142 581 143 585
rect 147 581 148 585
rect 142 580 148 581
rect 302 585 308 586
rect 302 581 303 585
rect 307 581 308 585
rect 302 580 308 581
rect 486 585 492 586
rect 486 581 487 585
rect 491 581 492 585
rect 486 580 492 581
rect 110 572 116 573
rect 110 568 111 572
rect 115 568 116 572
rect 664 568 666 606
rect 784 603 786 618
rect 936 603 938 618
rect 1080 603 1082 618
rect 1216 603 1218 618
rect 1352 603 1354 618
rect 671 602 675 603
rect 671 597 675 598
rect 783 602 787 603
rect 783 597 787 598
rect 847 602 851 603
rect 847 597 851 598
rect 935 602 939 603
rect 935 597 939 598
rect 1023 602 1027 603
rect 1023 597 1027 598
rect 1079 602 1083 603
rect 1079 597 1083 598
rect 1199 602 1203 603
rect 1199 597 1203 598
rect 1215 602 1219 603
rect 1215 597 1219 598
rect 1351 602 1355 603
rect 1351 597 1355 598
rect 1375 602 1379 603
rect 1375 597 1379 598
rect 672 586 674 597
rect 754 595 760 596
rect 754 591 755 595
rect 759 591 760 595
rect 754 590 760 591
rect 790 595 796 596
rect 790 591 791 595
rect 795 591 796 595
rect 790 590 796 591
rect 670 585 676 586
rect 670 581 671 585
rect 675 581 676 585
rect 670 580 676 581
rect 756 568 758 590
rect 110 567 116 568
rect 662 567 668 568
rect 662 563 663 567
rect 667 563 668 567
rect 662 562 668 563
rect 754 567 760 568
rect 754 563 755 567
rect 759 563 760 567
rect 754 562 760 563
rect 110 555 116 556
rect 110 551 111 555
rect 115 551 116 555
rect 110 550 116 551
rect 112 531 114 550
rect 134 545 140 546
rect 134 541 135 545
rect 139 541 140 545
rect 134 540 140 541
rect 294 545 300 546
rect 294 541 295 545
rect 299 541 300 545
rect 294 540 300 541
rect 478 545 484 546
rect 478 541 479 545
rect 483 541 484 545
rect 478 540 484 541
rect 662 545 668 546
rect 662 541 663 545
rect 667 541 668 545
rect 662 540 668 541
rect 136 531 138 540
rect 296 531 298 540
rect 480 531 482 540
rect 530 539 536 540
rect 530 535 531 539
rect 535 535 536 539
rect 530 534 536 535
rect 111 530 115 531
rect 111 525 115 526
rect 135 530 139 531
rect 135 525 139 526
rect 295 530 299 531
rect 295 525 299 526
rect 303 530 307 531
rect 303 525 307 526
rect 479 530 483 531
rect 479 525 483 526
rect 495 530 499 531
rect 495 525 499 526
rect 112 510 114 525
rect 136 520 138 525
rect 304 520 306 525
rect 496 520 498 525
rect 134 519 140 520
rect 134 515 135 519
rect 139 515 140 519
rect 134 514 140 515
rect 302 519 308 520
rect 302 515 303 519
rect 307 515 308 519
rect 302 514 308 515
rect 494 519 500 520
rect 494 515 495 519
rect 499 515 500 519
rect 494 514 500 515
rect 110 509 116 510
rect 110 505 111 509
rect 115 505 116 509
rect 110 504 116 505
rect 202 495 208 496
rect 110 492 116 493
rect 110 488 111 492
rect 115 488 116 492
rect 202 491 203 495
rect 207 491 208 495
rect 202 490 208 491
rect 370 495 376 496
rect 370 491 371 495
rect 375 491 376 495
rect 370 490 376 491
rect 110 487 116 488
rect 112 459 114 487
rect 142 479 148 480
rect 142 475 143 479
rect 147 475 148 479
rect 142 474 148 475
rect 144 459 146 474
rect 204 468 206 490
rect 310 479 316 480
rect 310 475 311 479
rect 315 475 316 479
rect 310 474 316 475
rect 202 467 208 468
rect 202 463 203 467
rect 207 463 208 467
rect 202 462 208 463
rect 312 459 314 474
rect 372 468 374 490
rect 502 479 508 480
rect 502 475 503 479
rect 507 475 508 479
rect 502 474 508 475
rect 370 467 376 468
rect 370 463 371 467
rect 375 463 376 467
rect 370 462 376 463
rect 504 459 506 474
rect 532 468 534 534
rect 664 531 666 540
rect 663 530 667 531
rect 663 525 667 526
rect 679 530 683 531
rect 679 525 683 526
rect 680 520 682 525
rect 678 519 684 520
rect 678 515 679 519
rect 683 515 684 519
rect 678 514 684 515
rect 792 512 794 590
rect 848 586 850 597
rect 1024 586 1026 597
rect 1038 595 1044 596
rect 1038 591 1039 595
rect 1043 591 1044 595
rect 1038 590 1044 591
rect 846 585 852 586
rect 846 581 847 585
rect 851 581 852 585
rect 846 580 852 581
rect 1022 585 1028 586
rect 1022 581 1023 585
rect 1027 581 1028 585
rect 1022 580 1028 581
rect 838 545 844 546
rect 838 541 839 545
rect 843 541 844 545
rect 838 540 844 541
rect 1014 545 1020 546
rect 1014 541 1015 545
rect 1019 541 1020 545
rect 1014 540 1020 541
rect 840 531 842 540
rect 1016 531 1018 540
rect 839 530 843 531
rect 839 525 843 526
rect 863 530 867 531
rect 863 525 867 526
rect 1015 530 1019 531
rect 1015 525 1019 526
rect 1031 530 1035 531
rect 1031 525 1035 526
rect 864 520 866 525
rect 1032 520 1034 525
rect 862 519 868 520
rect 862 515 863 519
rect 867 515 868 519
rect 862 514 868 515
rect 1030 519 1036 520
rect 1030 515 1031 519
rect 1035 515 1036 519
rect 1030 514 1036 515
rect 790 511 796 512
rect 790 507 791 511
rect 795 507 796 511
rect 1040 508 1042 590
rect 1200 586 1202 597
rect 1306 595 1312 596
rect 1306 591 1307 595
rect 1311 591 1312 595
rect 1306 590 1312 591
rect 1198 585 1204 586
rect 1198 581 1199 585
rect 1203 581 1204 585
rect 1198 580 1204 581
rect 1308 568 1310 590
rect 1376 586 1378 597
rect 1412 596 1414 634
rect 1420 620 1422 634
rect 1486 623 1492 624
rect 1418 619 1424 620
rect 1418 615 1419 619
rect 1423 615 1424 619
rect 1486 619 1487 623
rect 1491 619 1492 623
rect 1486 618 1492 619
rect 1418 614 1424 615
rect 1488 603 1490 618
rect 1520 612 1522 690
rect 1574 685 1580 686
rect 1574 681 1575 685
rect 1579 681 1580 685
rect 1574 680 1580 681
rect 1726 685 1732 686
rect 1726 681 1727 685
rect 1731 681 1732 685
rect 1726 680 1732 681
rect 1576 675 1578 680
rect 1728 675 1730 680
rect 1766 679 1772 680
rect 1766 675 1767 679
rect 1771 675 1772 679
rect 1824 675 1826 690
rect 1864 675 1866 694
rect 1886 689 1892 690
rect 1886 685 1887 689
rect 1891 685 1892 689
rect 1886 684 1892 685
rect 2054 689 2060 690
rect 2054 685 2055 689
rect 2059 685 2060 689
rect 2054 684 2060 685
rect 1888 675 1890 684
rect 2056 675 2058 684
rect 1575 674 1579 675
rect 1575 669 1579 670
rect 1615 674 1619 675
rect 1615 669 1619 670
rect 1727 674 1731 675
rect 1766 674 1772 675
rect 1823 674 1827 675
rect 1727 669 1731 670
rect 1616 664 1618 669
rect 1728 664 1730 669
rect 1614 663 1620 664
rect 1614 659 1615 663
rect 1619 659 1620 663
rect 1614 658 1620 659
rect 1726 663 1732 664
rect 1726 659 1727 663
rect 1731 659 1732 663
rect 1726 658 1732 659
rect 1590 639 1596 640
rect 1590 635 1591 639
rect 1595 635 1596 639
rect 1590 634 1596 635
rect 1682 639 1688 640
rect 1682 635 1683 639
rect 1687 635 1688 639
rect 1682 634 1688 635
rect 1518 611 1524 612
rect 1518 607 1519 611
rect 1523 607 1524 611
rect 1518 606 1524 607
rect 1487 602 1491 603
rect 1487 597 1491 598
rect 1559 602 1563 603
rect 1559 597 1563 598
rect 1406 595 1414 596
rect 1406 591 1407 595
rect 1411 592 1414 595
rect 1411 591 1412 592
rect 1406 590 1412 591
rect 1560 586 1562 597
rect 1592 596 1594 634
rect 1622 623 1628 624
rect 1622 619 1623 623
rect 1627 619 1628 623
rect 1622 618 1628 619
rect 1624 603 1626 618
rect 1684 612 1686 634
rect 1734 623 1740 624
rect 1734 619 1735 623
rect 1739 619 1740 623
rect 1734 618 1740 619
rect 1682 611 1688 612
rect 1682 607 1683 611
rect 1687 607 1688 611
rect 1682 606 1688 607
rect 1736 603 1738 618
rect 1768 612 1770 674
rect 1823 669 1827 670
rect 1863 674 1867 675
rect 1863 669 1867 670
rect 1887 674 1891 675
rect 1887 669 1891 670
rect 2055 674 2059 675
rect 2055 669 2059 670
rect 1824 654 1826 669
rect 1864 654 1866 669
rect 2096 656 2098 734
rect 2256 730 2258 741
rect 2448 730 2450 741
rect 2254 729 2260 730
rect 2254 725 2255 729
rect 2259 725 2260 729
rect 2254 724 2260 725
rect 2446 729 2452 730
rect 2446 725 2447 729
rect 2451 725 2452 729
rect 2446 724 2452 725
rect 2508 716 2510 750
rect 2632 747 2634 762
rect 2664 756 2666 834
rect 2838 829 2844 830
rect 2838 825 2839 829
rect 2843 825 2844 829
rect 2838 824 2844 825
rect 2880 824 2882 874
rect 3040 870 3042 881
rect 3092 880 3094 914
rect 3574 912 3575 916
rect 3579 912 3580 916
rect 3574 911 3580 912
rect 3576 887 3578 911
rect 3239 886 3243 887
rect 3239 881 3243 882
rect 3439 886 3443 887
rect 3439 881 3443 882
rect 3575 886 3579 887
rect 3575 881 3579 882
rect 3090 879 3096 880
rect 3090 875 3091 879
rect 3095 875 3096 879
rect 3090 874 3096 875
rect 3240 870 3242 881
rect 3406 879 3412 880
rect 3406 875 3407 879
rect 3411 875 3412 879
rect 3406 874 3412 875
rect 3038 869 3044 870
rect 3038 865 3039 869
rect 3043 865 3044 869
rect 3038 864 3044 865
rect 3238 869 3244 870
rect 3238 865 3239 869
rect 3243 865 3244 869
rect 3238 864 3244 865
rect 3030 829 3036 830
rect 3030 825 3031 829
rect 3035 825 3036 829
rect 3030 824 3036 825
rect 3230 829 3236 830
rect 3230 825 3231 829
rect 3235 825 3236 829
rect 3230 824 3236 825
rect 2840 819 2842 824
rect 2878 823 2884 824
rect 2878 819 2879 823
rect 2883 819 2884 823
rect 3032 819 3034 824
rect 3232 819 3234 824
rect 2799 818 2803 819
rect 2799 813 2803 814
rect 2839 818 2843 819
rect 2878 818 2884 819
rect 2967 818 2971 819
rect 2839 813 2843 814
rect 2967 813 2971 814
rect 3031 818 3035 819
rect 3031 813 3035 814
rect 3143 818 3147 819
rect 3143 813 3147 814
rect 3231 818 3235 819
rect 3231 813 3235 814
rect 3319 818 3323 819
rect 3319 813 3323 814
rect 2800 808 2802 813
rect 2968 808 2970 813
rect 3144 808 3146 813
rect 3320 808 3322 813
rect 2798 807 2804 808
rect 2798 803 2799 807
rect 2803 803 2804 807
rect 2798 802 2804 803
rect 2966 807 2972 808
rect 2966 803 2967 807
rect 2971 803 2972 807
rect 2966 802 2972 803
rect 3142 807 3148 808
rect 3142 803 3143 807
rect 3147 803 3148 807
rect 3142 802 3148 803
rect 3318 807 3324 808
rect 3318 803 3319 807
rect 3323 803 3324 807
rect 3318 802 3324 803
rect 3408 800 3410 874
rect 3440 870 3442 881
rect 3438 869 3444 870
rect 3438 865 3439 869
rect 3443 865 3444 869
rect 3438 864 3444 865
rect 3576 857 3578 881
rect 3574 856 3580 857
rect 3574 852 3575 856
rect 3579 852 3580 856
rect 3574 851 3580 852
rect 3514 839 3520 840
rect 3514 835 3515 839
rect 3519 835 3520 839
rect 3514 834 3520 835
rect 3574 839 3580 840
rect 3574 835 3575 839
rect 3579 835 3580 839
rect 3574 834 3580 835
rect 3430 829 3436 830
rect 3430 825 3431 829
rect 3435 825 3436 829
rect 3430 824 3436 825
rect 3432 819 3434 824
rect 3431 818 3435 819
rect 3431 813 3435 814
rect 3479 818 3483 819
rect 3479 813 3483 814
rect 3480 808 3482 813
rect 3478 807 3484 808
rect 3478 803 3479 807
rect 3483 803 3484 807
rect 3478 802 3484 803
rect 3406 799 3412 800
rect 3406 795 3407 799
rect 3411 795 3412 799
rect 3406 794 3412 795
rect 2866 783 2872 784
rect 2866 779 2867 783
rect 2871 779 2872 783
rect 2866 778 2872 779
rect 2806 767 2812 768
rect 2806 763 2807 767
rect 2811 763 2812 767
rect 2806 762 2812 763
rect 2662 755 2668 756
rect 2662 751 2663 755
rect 2667 751 2668 755
rect 2662 750 2668 751
rect 2808 747 2810 762
rect 2631 746 2635 747
rect 2631 741 2635 742
rect 2639 746 2643 747
rect 2639 741 2643 742
rect 2807 746 2811 747
rect 2807 741 2811 742
rect 2823 746 2827 747
rect 2823 741 2827 742
rect 2640 730 2642 741
rect 2730 739 2736 740
rect 2730 735 2731 739
rect 2735 735 2736 739
rect 2730 734 2736 735
rect 2638 729 2644 730
rect 2638 725 2639 729
rect 2643 725 2644 729
rect 2638 724 2644 725
rect 2506 715 2512 716
rect 2506 711 2507 715
rect 2511 711 2512 715
rect 2732 712 2734 734
rect 2824 730 2826 741
rect 2868 740 2870 778
rect 2974 767 2980 768
rect 2974 763 2975 767
rect 2979 763 2980 767
rect 2974 762 2980 763
rect 3150 767 3156 768
rect 3150 763 3151 767
rect 3155 763 3156 767
rect 3150 762 3156 763
rect 3326 767 3332 768
rect 3326 763 3327 767
rect 3331 763 3332 767
rect 3326 762 3332 763
rect 3486 767 3492 768
rect 3486 763 3487 767
rect 3491 763 3492 767
rect 3486 762 3492 763
rect 2976 747 2978 762
rect 3152 747 3154 762
rect 3234 755 3240 756
rect 3234 751 3235 755
rect 3239 751 3240 755
rect 3234 750 3240 751
rect 2975 746 2979 747
rect 2975 741 2979 742
rect 2999 746 3003 747
rect 2999 741 3003 742
rect 3151 746 3155 747
rect 3151 741 3155 742
rect 3167 746 3171 747
rect 3167 741 3171 742
rect 2866 739 2872 740
rect 2866 735 2867 739
rect 2871 735 2872 739
rect 2866 734 2872 735
rect 3000 730 3002 741
rect 3058 739 3064 740
rect 3058 735 3059 739
rect 3063 735 3064 739
rect 3058 734 3064 735
rect 2822 729 2828 730
rect 2822 725 2823 729
rect 2827 725 2828 729
rect 2822 724 2828 725
rect 2998 729 3004 730
rect 2998 725 2999 729
rect 3003 725 3004 729
rect 2998 724 3004 725
rect 2506 710 2512 711
rect 2730 711 2736 712
rect 2730 707 2731 711
rect 2735 707 2736 711
rect 2730 706 2736 707
rect 2706 699 2712 700
rect 2706 695 2707 699
rect 2711 695 2712 699
rect 2706 694 2712 695
rect 2246 689 2252 690
rect 2246 685 2247 689
rect 2251 685 2252 689
rect 2246 684 2252 685
rect 2438 689 2444 690
rect 2438 685 2439 689
rect 2443 685 2444 689
rect 2438 684 2444 685
rect 2630 689 2636 690
rect 2630 685 2631 689
rect 2635 685 2636 689
rect 2630 684 2636 685
rect 2248 675 2250 684
rect 2440 675 2442 684
rect 2632 675 2634 684
rect 2215 674 2219 675
rect 2215 669 2219 670
rect 2247 674 2251 675
rect 2247 669 2251 670
rect 2359 674 2363 675
rect 2359 669 2363 670
rect 2439 674 2443 675
rect 2439 669 2443 670
rect 2511 674 2515 675
rect 2511 669 2515 670
rect 2631 674 2635 675
rect 2631 669 2635 670
rect 2671 674 2675 675
rect 2671 669 2675 670
rect 2216 664 2218 669
rect 2360 664 2362 669
rect 2512 664 2514 669
rect 2672 664 2674 669
rect 2214 663 2220 664
rect 2214 659 2215 663
rect 2219 659 2220 663
rect 2214 658 2220 659
rect 2358 663 2364 664
rect 2358 659 2359 663
rect 2363 659 2364 663
rect 2358 658 2364 659
rect 2510 663 2516 664
rect 2510 659 2511 663
rect 2515 659 2516 663
rect 2510 658 2516 659
rect 2670 663 2676 664
rect 2670 659 2671 663
rect 2675 659 2676 663
rect 2670 658 2676 659
rect 2094 655 2100 656
rect 1822 653 1828 654
rect 1822 649 1823 653
rect 1827 649 1828 653
rect 1822 648 1828 649
rect 1862 653 1868 654
rect 1862 649 1863 653
rect 1867 649 1868 653
rect 2094 651 2095 655
rect 2099 651 2100 655
rect 2094 650 2100 651
rect 1862 648 1868 649
rect 2282 639 2288 640
rect 1822 636 1828 637
rect 1822 632 1823 636
rect 1827 632 1828 636
rect 1822 631 1828 632
rect 1862 636 1868 637
rect 1862 632 1863 636
rect 1867 632 1868 636
rect 2282 635 2283 639
rect 2287 635 2288 639
rect 2282 634 2288 635
rect 2426 639 2432 640
rect 2426 635 2427 639
rect 2431 635 2432 639
rect 2426 634 2432 635
rect 1862 631 1868 632
rect 1766 611 1772 612
rect 1766 607 1767 611
rect 1771 607 1772 611
rect 1766 606 1772 607
rect 1824 603 1826 631
rect 1864 603 1866 631
rect 2222 623 2228 624
rect 2222 619 2223 623
rect 2227 619 2228 623
rect 2222 618 2228 619
rect 2224 603 2226 618
rect 2284 612 2286 634
rect 2366 623 2372 624
rect 2366 619 2367 623
rect 2371 619 2372 623
rect 2366 618 2372 619
rect 2282 611 2288 612
rect 2282 607 2283 611
rect 2287 607 2288 611
rect 2282 606 2288 607
rect 2368 603 2370 618
rect 2428 612 2430 634
rect 2518 623 2524 624
rect 2518 619 2519 623
rect 2523 619 2524 623
rect 2518 618 2524 619
rect 2678 623 2684 624
rect 2678 619 2679 623
rect 2683 619 2684 623
rect 2678 618 2684 619
rect 2426 611 2432 612
rect 2426 607 2427 611
rect 2431 607 2432 611
rect 2426 606 2432 607
rect 2520 603 2522 618
rect 2680 603 2682 618
rect 2708 612 2710 694
rect 2814 689 2820 690
rect 2814 685 2815 689
rect 2819 685 2820 689
rect 2814 684 2820 685
rect 2990 689 2996 690
rect 2990 685 2991 689
rect 2995 685 2996 689
rect 2990 684 2996 685
rect 2816 675 2818 684
rect 2992 675 2994 684
rect 2815 674 2819 675
rect 2815 669 2819 670
rect 2831 674 2835 675
rect 2831 669 2835 670
rect 2991 674 2995 675
rect 2991 669 2995 670
rect 2832 664 2834 669
rect 2992 664 2994 669
rect 2830 663 2836 664
rect 2830 659 2831 663
rect 2835 659 2836 663
rect 2830 658 2836 659
rect 2990 663 2996 664
rect 2990 659 2991 663
rect 2995 659 2996 663
rect 2990 658 2996 659
rect 3060 656 3062 734
rect 3168 730 3170 741
rect 3226 739 3232 740
rect 3226 735 3227 739
rect 3231 735 3232 739
rect 3226 734 3232 735
rect 3166 729 3172 730
rect 3166 725 3167 729
rect 3171 725 3172 729
rect 3166 724 3172 725
rect 3228 716 3230 734
rect 3226 715 3232 716
rect 3226 711 3227 715
rect 3231 711 3232 715
rect 3236 712 3238 750
rect 3328 747 3330 762
rect 3488 747 3490 762
rect 3516 756 3518 834
rect 3576 819 3578 834
rect 3575 818 3579 819
rect 3575 813 3579 814
rect 3576 798 3578 813
rect 3574 797 3580 798
rect 3574 793 3575 797
rect 3579 793 3580 797
rect 3574 792 3580 793
rect 3546 783 3552 784
rect 3546 779 3547 783
rect 3551 779 3552 783
rect 3546 778 3552 779
rect 3574 780 3580 781
rect 3514 755 3520 756
rect 3514 751 3515 755
rect 3519 751 3520 755
rect 3514 750 3520 751
rect 3327 746 3331 747
rect 3327 741 3331 742
rect 3335 746 3339 747
rect 3335 741 3339 742
rect 3487 746 3491 747
rect 3487 741 3491 742
rect 3336 730 3338 741
rect 3488 730 3490 741
rect 3548 740 3550 778
rect 3574 776 3575 780
rect 3579 776 3580 780
rect 3574 775 3580 776
rect 3576 747 3578 775
rect 3575 746 3579 747
rect 3575 741 3579 742
rect 3546 739 3552 740
rect 3546 735 3547 739
rect 3551 735 3552 739
rect 3546 734 3552 735
rect 3334 729 3340 730
rect 3334 725 3335 729
rect 3339 725 3340 729
rect 3334 724 3340 725
rect 3486 729 3492 730
rect 3486 725 3487 729
rect 3491 725 3492 729
rect 3486 724 3492 725
rect 3576 717 3578 741
rect 3574 716 3580 717
rect 3574 712 3575 716
rect 3579 712 3580 716
rect 3226 710 3232 711
rect 3234 711 3240 712
rect 3574 711 3580 712
rect 3234 707 3235 711
rect 3239 707 3240 711
rect 3234 706 3240 707
rect 3574 699 3580 700
rect 3574 695 3575 699
rect 3579 695 3580 699
rect 3574 694 3580 695
rect 3158 689 3164 690
rect 3158 685 3159 689
rect 3163 685 3164 689
rect 3158 684 3164 685
rect 3326 689 3332 690
rect 3326 685 3327 689
rect 3331 685 3332 689
rect 3326 684 3332 685
rect 3478 689 3484 690
rect 3478 685 3479 689
rect 3483 685 3484 689
rect 3478 684 3484 685
rect 3160 675 3162 684
rect 3328 675 3330 684
rect 3480 675 3482 684
rect 3518 683 3524 684
rect 3518 679 3519 683
rect 3523 679 3524 683
rect 3518 678 3524 679
rect 3159 674 3163 675
rect 3159 669 3163 670
rect 3327 674 3331 675
rect 3327 669 3331 670
rect 3479 674 3483 675
rect 3479 669 3483 670
rect 3160 664 3162 669
rect 3328 664 3330 669
rect 3480 664 3482 669
rect 3158 663 3164 664
rect 3158 659 3159 663
rect 3163 659 3164 663
rect 3158 658 3164 659
rect 3326 663 3332 664
rect 3326 659 3327 663
rect 3331 659 3332 663
rect 3326 658 3332 659
rect 3478 663 3484 664
rect 3478 659 3479 663
rect 3483 659 3484 663
rect 3478 658 3484 659
rect 3058 655 3064 656
rect 3058 651 3059 655
rect 3063 651 3064 655
rect 3058 650 3064 651
rect 2822 639 2828 640
rect 2822 635 2823 639
rect 2827 635 2828 639
rect 2822 634 2828 635
rect 2982 639 2988 640
rect 2982 635 2983 639
rect 2987 635 2988 639
rect 2982 634 2988 635
rect 3058 639 3064 640
rect 3058 635 3059 639
rect 3063 635 3064 639
rect 3058 634 3064 635
rect 3226 639 3232 640
rect 3226 635 3227 639
rect 3231 635 3232 639
rect 3226 634 3232 635
rect 2824 612 2826 634
rect 2838 623 2844 624
rect 2838 619 2839 623
rect 2843 619 2844 623
rect 2838 618 2844 619
rect 2706 611 2712 612
rect 2706 607 2707 611
rect 2711 607 2712 611
rect 2706 606 2712 607
rect 2822 611 2828 612
rect 2822 607 2823 611
rect 2827 607 2828 611
rect 2822 606 2828 607
rect 2746 603 2752 604
rect 2840 603 2842 618
rect 1623 602 1627 603
rect 1623 597 1627 598
rect 1735 602 1739 603
rect 1735 597 1739 598
rect 1823 602 1827 603
rect 1823 597 1827 598
rect 1863 602 1867 603
rect 1863 597 1867 598
rect 2199 602 2203 603
rect 2199 597 2203 598
rect 2223 602 2227 603
rect 2223 597 2227 598
rect 2287 602 2291 603
rect 2287 597 2291 598
rect 2367 602 2371 603
rect 2367 597 2371 598
rect 2375 602 2379 603
rect 2375 597 2379 598
rect 2463 602 2467 603
rect 2463 597 2467 598
rect 2519 602 2523 603
rect 2519 597 2523 598
rect 2567 602 2571 603
rect 2567 597 2571 598
rect 2679 602 2683 603
rect 2746 599 2747 603
rect 2751 599 2752 603
rect 2746 598 2752 599
rect 2815 602 2819 603
rect 2679 597 2683 598
rect 1590 595 1596 596
rect 1590 591 1591 595
rect 1595 591 1596 595
rect 1590 590 1596 591
rect 1736 586 1738 597
rect 1374 585 1380 586
rect 1374 581 1375 585
rect 1379 581 1380 585
rect 1374 580 1380 581
rect 1558 585 1564 586
rect 1558 581 1559 585
rect 1563 581 1564 585
rect 1558 580 1564 581
rect 1734 585 1740 586
rect 1734 581 1735 585
rect 1739 581 1740 585
rect 1734 580 1740 581
rect 1824 573 1826 597
rect 1864 573 1866 597
rect 2200 586 2202 597
rect 2230 595 2236 596
rect 2230 591 2231 595
rect 2235 591 2236 595
rect 2230 590 2236 591
rect 2198 585 2204 586
rect 2198 581 2199 585
rect 2203 581 2204 585
rect 2198 580 2204 581
rect 1822 572 1828 573
rect 1822 568 1823 572
rect 1827 568 1828 572
rect 1306 567 1312 568
rect 1822 567 1828 568
rect 1862 572 1868 573
rect 1862 568 1863 572
rect 1867 568 1868 572
rect 1862 567 1868 568
rect 1306 563 1307 567
rect 1311 563 1312 567
rect 1306 562 1312 563
rect 1702 555 1708 556
rect 1702 551 1703 555
rect 1707 551 1708 555
rect 1702 550 1708 551
rect 1822 555 1828 556
rect 1822 551 1823 555
rect 1827 551 1828 555
rect 1822 550 1828 551
rect 1862 555 1868 556
rect 1862 551 1863 555
rect 1867 551 1868 555
rect 1862 550 1868 551
rect 1190 545 1196 546
rect 1190 541 1191 545
rect 1195 541 1196 545
rect 1190 540 1196 541
rect 1366 545 1372 546
rect 1366 541 1367 545
rect 1371 541 1372 545
rect 1366 540 1372 541
rect 1550 545 1556 546
rect 1550 541 1551 545
rect 1555 541 1556 545
rect 1550 540 1556 541
rect 1192 531 1194 540
rect 1230 539 1236 540
rect 1230 535 1231 539
rect 1235 535 1236 539
rect 1230 534 1236 535
rect 1191 530 1195 531
rect 1191 525 1195 526
rect 1192 520 1194 525
rect 1190 519 1196 520
rect 1190 515 1191 519
rect 1195 515 1196 519
rect 1190 514 1196 515
rect 790 506 796 507
rect 1038 507 1044 508
rect 1038 503 1039 507
rect 1043 503 1044 507
rect 1038 502 1044 503
rect 746 495 752 496
rect 746 491 747 495
rect 751 491 752 495
rect 746 490 752 491
rect 686 479 692 480
rect 686 475 687 479
rect 691 475 692 479
rect 686 474 692 475
rect 530 467 536 468
rect 530 463 531 467
rect 535 463 536 467
rect 530 462 536 463
rect 688 459 690 474
rect 748 468 750 490
rect 870 479 876 480
rect 870 475 871 479
rect 875 475 876 479
rect 870 474 876 475
rect 1038 479 1044 480
rect 1038 475 1039 479
rect 1043 475 1044 479
rect 1038 474 1044 475
rect 1198 479 1204 480
rect 1198 475 1199 479
rect 1203 475 1204 479
rect 1198 474 1204 475
rect 746 467 752 468
rect 746 463 747 467
rect 751 463 752 467
rect 746 462 752 463
rect 872 459 874 474
rect 938 467 944 468
rect 938 463 939 467
rect 943 463 944 467
rect 938 462 944 463
rect 111 458 115 459
rect 111 453 115 454
rect 143 458 147 459
rect 143 453 147 454
rect 303 458 307 459
rect 303 453 307 454
rect 311 458 315 459
rect 311 453 315 454
rect 495 458 499 459
rect 495 453 499 454
rect 503 458 507 459
rect 503 453 507 454
rect 687 458 691 459
rect 687 453 691 454
rect 871 458 875 459
rect 871 453 875 454
rect 879 458 883 459
rect 879 453 883 454
rect 112 429 114 453
rect 144 442 146 453
rect 304 442 306 453
rect 496 442 498 453
rect 688 442 690 453
rect 880 442 882 453
rect 142 441 148 442
rect 142 437 143 441
rect 147 437 148 441
rect 142 436 148 437
rect 302 441 308 442
rect 302 437 303 441
rect 307 437 308 441
rect 302 436 308 437
rect 494 441 500 442
rect 494 437 495 441
rect 499 437 500 441
rect 494 436 500 437
rect 686 441 692 442
rect 686 437 687 441
rect 691 437 692 441
rect 686 436 692 437
rect 878 441 884 442
rect 878 437 879 441
rect 883 437 884 441
rect 878 436 884 437
rect 110 428 116 429
rect 940 428 942 462
rect 1040 459 1042 474
rect 1046 467 1052 468
rect 1046 463 1047 467
rect 1051 463 1052 467
rect 1046 462 1052 463
rect 1039 458 1043 459
rect 1039 453 1043 454
rect 110 424 111 428
rect 115 424 116 428
rect 110 423 116 424
rect 938 427 944 428
rect 938 423 939 427
rect 943 423 944 427
rect 1048 424 1050 462
rect 1200 459 1202 474
rect 1232 468 1234 534
rect 1368 531 1370 540
rect 1552 531 1554 540
rect 1351 530 1355 531
rect 1351 525 1355 526
rect 1367 530 1371 531
rect 1367 525 1371 526
rect 1503 530 1507 531
rect 1503 525 1507 526
rect 1551 530 1555 531
rect 1551 525 1555 526
rect 1663 530 1667 531
rect 1663 525 1667 526
rect 1352 520 1354 525
rect 1504 520 1506 525
rect 1664 520 1666 525
rect 1350 519 1356 520
rect 1350 515 1351 519
rect 1355 515 1356 519
rect 1350 514 1356 515
rect 1502 519 1508 520
rect 1502 515 1503 519
rect 1507 515 1508 519
rect 1502 514 1508 515
rect 1662 519 1668 520
rect 1662 515 1663 519
rect 1667 515 1668 519
rect 1662 514 1668 515
rect 1418 495 1424 496
rect 1418 491 1419 495
rect 1423 491 1424 495
rect 1418 490 1424 491
rect 1570 495 1576 496
rect 1570 491 1571 495
rect 1575 491 1576 495
rect 1570 490 1576 491
rect 1358 479 1364 480
rect 1358 475 1359 479
rect 1363 475 1364 479
rect 1358 474 1364 475
rect 1230 467 1236 468
rect 1230 463 1231 467
rect 1235 463 1236 467
rect 1230 462 1236 463
rect 1360 459 1362 474
rect 1055 458 1059 459
rect 1055 453 1059 454
rect 1199 458 1203 459
rect 1199 453 1203 454
rect 1223 458 1227 459
rect 1223 453 1227 454
rect 1359 458 1363 459
rect 1359 453 1363 454
rect 1391 458 1395 459
rect 1391 453 1395 454
rect 1056 442 1058 453
rect 1094 451 1100 452
rect 1094 447 1095 451
rect 1099 447 1100 451
rect 1094 446 1100 447
rect 1054 441 1060 442
rect 1054 437 1055 441
rect 1059 437 1060 441
rect 1054 436 1060 437
rect 938 422 944 423
rect 1046 423 1052 424
rect 1046 419 1047 423
rect 1051 419 1052 423
rect 1046 418 1052 419
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 110 406 116 407
rect 462 411 468 412
rect 462 407 463 411
rect 467 407 468 411
rect 462 406 468 407
rect 112 391 114 406
rect 134 401 140 402
rect 134 397 135 401
rect 139 397 140 401
rect 134 396 140 397
rect 294 401 300 402
rect 294 397 295 401
rect 299 397 300 401
rect 294 396 300 397
rect 136 391 138 396
rect 296 391 298 396
rect 111 390 115 391
rect 111 385 115 386
rect 135 390 139 391
rect 135 385 139 386
rect 263 390 267 391
rect 263 385 267 386
rect 295 390 299 391
rect 295 385 299 386
rect 423 390 427 391
rect 423 385 427 386
rect 112 370 114 385
rect 136 380 138 385
rect 264 380 266 385
rect 424 380 426 385
rect 134 379 140 380
rect 134 375 135 379
rect 139 375 140 379
rect 134 374 140 375
rect 262 379 268 380
rect 262 375 263 379
rect 267 375 268 379
rect 262 374 268 375
rect 422 379 428 380
rect 422 375 423 379
rect 427 375 428 379
rect 422 374 428 375
rect 110 369 116 370
rect 110 365 111 369
rect 115 365 116 369
rect 110 364 116 365
rect 330 355 336 356
rect 110 352 116 353
rect 110 348 111 352
rect 115 348 116 352
rect 330 351 331 355
rect 335 351 336 355
rect 330 350 336 351
rect 110 347 116 348
rect 242 347 248 348
rect 112 323 114 347
rect 242 343 243 347
rect 247 343 248 347
rect 242 342 248 343
rect 142 339 148 340
rect 142 335 143 339
rect 147 335 148 339
rect 142 334 148 335
rect 144 323 146 334
rect 111 322 115 323
rect 111 317 115 318
rect 143 322 147 323
rect 143 317 147 318
rect 215 322 219 323
rect 215 317 219 318
rect 112 293 114 317
rect 216 306 218 317
rect 244 316 246 342
rect 270 339 276 340
rect 270 335 271 339
rect 275 335 276 339
rect 270 334 276 335
rect 272 323 274 334
rect 332 328 334 350
rect 430 339 436 340
rect 430 335 431 339
rect 435 335 436 339
rect 430 334 436 335
rect 330 327 336 328
rect 330 323 331 327
rect 335 323 336 327
rect 432 323 434 334
rect 464 328 466 406
rect 486 401 492 402
rect 486 397 487 401
rect 491 397 492 401
rect 486 396 492 397
rect 678 401 684 402
rect 678 397 679 401
rect 683 397 684 401
rect 678 396 684 397
rect 870 401 876 402
rect 870 397 871 401
rect 875 397 876 401
rect 870 396 876 397
rect 1046 401 1052 402
rect 1046 397 1047 401
rect 1051 397 1052 401
rect 1046 396 1052 397
rect 488 391 490 396
rect 680 391 682 396
rect 872 391 874 396
rect 1048 391 1050 396
rect 487 390 491 391
rect 487 385 491 386
rect 591 390 595 391
rect 591 385 595 386
rect 679 390 683 391
rect 679 385 683 386
rect 767 390 771 391
rect 767 385 771 386
rect 871 390 875 391
rect 871 385 875 386
rect 935 390 939 391
rect 935 385 939 386
rect 1047 390 1051 391
rect 1047 385 1051 386
rect 592 380 594 385
rect 768 380 770 385
rect 936 380 938 385
rect 590 379 596 380
rect 590 375 591 379
rect 595 375 596 379
rect 590 374 596 375
rect 766 379 772 380
rect 766 375 767 379
rect 771 375 772 379
rect 766 374 772 375
rect 934 379 940 380
rect 934 375 935 379
rect 939 375 940 379
rect 934 374 940 375
rect 1096 372 1098 446
rect 1224 442 1226 453
rect 1290 451 1296 452
rect 1290 447 1291 451
rect 1295 447 1296 451
rect 1290 446 1296 447
rect 1222 441 1228 442
rect 1222 437 1223 441
rect 1227 437 1228 441
rect 1222 436 1228 437
rect 1292 424 1294 446
rect 1392 442 1394 453
rect 1420 452 1422 490
rect 1510 479 1516 480
rect 1510 475 1511 479
rect 1515 475 1516 479
rect 1510 474 1516 475
rect 1512 459 1514 474
rect 1572 468 1574 490
rect 1586 487 1592 488
rect 1586 483 1587 487
rect 1591 483 1592 487
rect 1586 482 1592 483
rect 1570 467 1576 468
rect 1570 463 1571 467
rect 1575 463 1576 467
rect 1570 462 1576 463
rect 1511 458 1515 459
rect 1511 453 1515 454
rect 1559 458 1563 459
rect 1559 453 1563 454
rect 1418 451 1424 452
rect 1418 447 1419 451
rect 1423 447 1424 451
rect 1418 446 1424 447
rect 1560 442 1562 453
rect 1588 452 1590 482
rect 1670 479 1676 480
rect 1670 475 1671 479
rect 1675 475 1676 479
rect 1670 474 1676 475
rect 1672 459 1674 474
rect 1704 468 1706 550
rect 1726 545 1732 546
rect 1726 541 1727 545
rect 1731 541 1732 545
rect 1726 540 1732 541
rect 1728 531 1730 540
rect 1824 531 1826 550
rect 1864 531 1866 550
rect 2190 545 2196 546
rect 2190 541 2191 545
rect 2195 541 2196 545
rect 2190 540 2196 541
rect 2192 531 2194 540
rect 1727 530 1731 531
rect 1727 525 1731 526
rect 1823 530 1827 531
rect 1823 525 1827 526
rect 1863 530 1867 531
rect 1863 525 1867 526
rect 2191 530 2195 531
rect 2191 525 2195 526
rect 1824 510 1826 525
rect 1864 510 1866 525
rect 2232 512 2234 590
rect 2288 586 2290 597
rect 2376 586 2378 597
rect 2464 586 2466 597
rect 2568 586 2570 597
rect 2680 586 2682 597
rect 2286 585 2292 586
rect 2286 581 2287 585
rect 2291 581 2292 585
rect 2286 580 2292 581
rect 2374 585 2380 586
rect 2374 581 2375 585
rect 2379 581 2380 585
rect 2374 580 2380 581
rect 2462 585 2468 586
rect 2462 581 2463 585
rect 2467 581 2468 585
rect 2462 580 2468 581
rect 2566 585 2572 586
rect 2566 581 2567 585
rect 2571 581 2572 585
rect 2566 580 2572 581
rect 2678 585 2684 586
rect 2678 581 2679 585
rect 2683 581 2684 585
rect 2678 580 2684 581
rect 2748 568 2750 598
rect 2815 597 2819 598
rect 2839 602 2843 603
rect 2839 597 2843 598
rect 2975 602 2979 603
rect 2975 597 2979 598
rect 2816 586 2818 597
rect 2914 595 2920 596
rect 2914 591 2915 595
rect 2919 591 2920 595
rect 2914 590 2920 591
rect 2814 585 2820 586
rect 2814 581 2815 585
rect 2819 581 2820 585
rect 2814 580 2820 581
rect 2916 568 2918 590
rect 2976 586 2978 597
rect 2984 596 2986 634
rect 2998 623 3004 624
rect 2998 619 2999 623
rect 3003 619 3004 623
rect 2998 618 3004 619
rect 3000 603 3002 618
rect 3060 612 3062 634
rect 3166 623 3172 624
rect 3166 619 3167 623
rect 3171 619 3172 623
rect 3166 618 3172 619
rect 3058 611 3064 612
rect 3058 607 3059 611
rect 3063 607 3064 611
rect 3058 606 3064 607
rect 3168 603 3170 618
rect 3228 612 3230 634
rect 3334 623 3340 624
rect 3334 619 3335 623
rect 3339 619 3340 623
rect 3334 618 3340 619
rect 3486 623 3492 624
rect 3486 619 3487 623
rect 3491 619 3492 623
rect 3486 618 3492 619
rect 3226 611 3232 612
rect 3226 607 3227 611
rect 3231 607 3232 611
rect 3226 606 3232 607
rect 3336 603 3338 618
rect 3386 611 3392 612
rect 3386 607 3387 611
rect 3391 607 3392 611
rect 3386 606 3392 607
rect 2999 602 3003 603
rect 2999 597 3003 598
rect 3143 602 3147 603
rect 3143 597 3147 598
rect 3167 602 3171 603
rect 3167 597 3171 598
rect 3327 602 3331 603
rect 3327 597 3331 598
rect 3335 602 3339 603
rect 3335 597 3339 598
rect 2982 595 2988 596
rect 2982 591 2983 595
rect 2987 591 2988 595
rect 2982 590 2988 591
rect 3144 586 3146 597
rect 3174 595 3180 596
rect 3174 591 3175 595
rect 3179 591 3180 595
rect 3174 590 3180 591
rect 2974 585 2980 586
rect 2974 581 2975 585
rect 2979 581 2980 585
rect 2974 580 2980 581
rect 3142 585 3148 586
rect 3142 581 3143 585
rect 3147 581 3148 585
rect 3142 580 3148 581
rect 2746 567 2752 568
rect 2746 563 2747 567
rect 2751 563 2752 567
rect 2746 562 2752 563
rect 2914 567 2920 568
rect 2914 563 2915 567
rect 2919 563 2920 567
rect 2914 562 2920 563
rect 2754 555 2760 556
rect 2754 551 2755 555
rect 2759 551 2760 555
rect 2754 550 2760 551
rect 2278 545 2284 546
rect 2278 541 2279 545
rect 2283 541 2284 545
rect 2278 540 2284 541
rect 2366 545 2372 546
rect 2366 541 2367 545
rect 2371 541 2372 545
rect 2366 540 2372 541
rect 2454 545 2460 546
rect 2454 541 2455 545
rect 2459 541 2460 545
rect 2454 540 2460 541
rect 2558 545 2564 546
rect 2558 541 2559 545
rect 2563 541 2564 545
rect 2558 540 2564 541
rect 2670 545 2676 546
rect 2670 541 2671 545
rect 2675 541 2676 545
rect 2670 540 2676 541
rect 2280 531 2282 540
rect 2368 531 2370 540
rect 2456 531 2458 540
rect 2560 531 2562 540
rect 2672 531 2674 540
rect 2279 530 2283 531
rect 2279 525 2283 526
rect 2303 530 2307 531
rect 2303 525 2307 526
rect 2367 530 2371 531
rect 2367 525 2371 526
rect 2399 530 2403 531
rect 2399 525 2403 526
rect 2455 530 2459 531
rect 2455 525 2459 526
rect 2503 530 2507 531
rect 2503 525 2507 526
rect 2559 530 2563 531
rect 2559 525 2563 526
rect 2607 530 2611 531
rect 2607 525 2611 526
rect 2671 530 2675 531
rect 2671 525 2675 526
rect 2719 530 2723 531
rect 2719 525 2723 526
rect 2304 520 2306 525
rect 2400 520 2402 525
rect 2504 520 2506 525
rect 2608 520 2610 525
rect 2720 520 2722 525
rect 2302 519 2308 520
rect 2302 515 2303 519
rect 2307 515 2308 519
rect 2302 514 2308 515
rect 2398 519 2404 520
rect 2398 515 2399 519
rect 2403 515 2404 519
rect 2398 514 2404 515
rect 2502 519 2508 520
rect 2502 515 2503 519
rect 2507 515 2508 519
rect 2502 514 2508 515
rect 2606 519 2612 520
rect 2606 515 2607 519
rect 2611 515 2612 519
rect 2606 514 2612 515
rect 2718 519 2724 520
rect 2718 515 2719 519
rect 2723 515 2724 519
rect 2718 514 2724 515
rect 2230 511 2236 512
rect 1822 509 1828 510
rect 1822 505 1823 509
rect 1827 505 1828 509
rect 1822 504 1828 505
rect 1862 509 1868 510
rect 1862 505 1863 509
rect 1867 505 1868 509
rect 2230 507 2231 511
rect 2235 507 2236 511
rect 2230 506 2236 507
rect 1862 504 1868 505
rect 2370 495 2376 496
rect 1822 492 1828 493
rect 1822 488 1823 492
rect 1827 488 1828 492
rect 1822 487 1828 488
rect 1862 492 1868 493
rect 1862 488 1863 492
rect 1867 488 1868 492
rect 2370 491 2371 495
rect 2375 491 2376 495
rect 2370 490 2376 491
rect 2466 495 2472 496
rect 2466 491 2467 495
rect 2471 491 2472 495
rect 2466 490 2472 491
rect 2570 495 2576 496
rect 2570 491 2571 495
rect 2575 491 2576 495
rect 2570 490 2576 491
rect 1862 487 1868 488
rect 1702 467 1708 468
rect 1702 463 1703 467
rect 1707 463 1708 467
rect 1702 462 1708 463
rect 1824 459 1826 487
rect 1864 463 1866 487
rect 2310 479 2316 480
rect 2310 475 2311 479
rect 2315 475 2316 479
rect 2310 474 2316 475
rect 2312 463 2314 474
rect 2372 468 2374 490
rect 2406 479 2412 480
rect 2406 475 2407 479
rect 2411 475 2412 479
rect 2406 474 2412 475
rect 2370 467 2376 468
rect 2370 463 2371 467
rect 2375 463 2376 467
rect 2408 463 2410 474
rect 2468 468 2470 490
rect 2510 479 2516 480
rect 2510 475 2511 479
rect 2515 475 2516 479
rect 2510 474 2516 475
rect 2466 467 2472 468
rect 2466 463 2467 467
rect 2471 463 2472 467
rect 2512 463 2514 474
rect 2572 468 2574 490
rect 2614 479 2620 480
rect 2614 475 2615 479
rect 2619 475 2620 479
rect 2614 474 2620 475
rect 2726 479 2732 480
rect 2726 475 2727 479
rect 2731 475 2732 479
rect 2726 474 2732 475
rect 2570 467 2576 468
rect 2570 463 2571 467
rect 2575 463 2576 467
rect 2616 463 2618 474
rect 2646 467 2652 468
rect 2646 463 2647 467
rect 2651 463 2652 467
rect 2728 463 2730 474
rect 2756 468 2758 550
rect 2806 545 2812 546
rect 2806 541 2807 545
rect 2811 541 2812 545
rect 2806 540 2812 541
rect 2966 545 2972 546
rect 2966 541 2967 545
rect 2971 541 2972 545
rect 2966 540 2972 541
rect 3134 545 3140 546
rect 3134 541 3135 545
rect 3139 541 3140 545
rect 3134 540 3140 541
rect 2808 531 2810 540
rect 2968 531 2970 540
rect 3136 531 3138 540
rect 2807 530 2811 531
rect 2807 525 2811 526
rect 2839 530 2843 531
rect 2839 525 2843 526
rect 2967 530 2971 531
rect 2967 525 2971 526
rect 3095 530 3099 531
rect 3095 525 3099 526
rect 3135 530 3139 531
rect 3135 525 3139 526
rect 2840 520 2842 525
rect 2968 520 2970 525
rect 3096 520 3098 525
rect 2838 519 2844 520
rect 2838 515 2839 519
rect 2843 515 2844 519
rect 2838 514 2844 515
rect 2966 519 2972 520
rect 2966 515 2967 519
rect 2971 515 2972 519
rect 2966 514 2972 515
rect 3094 519 3100 520
rect 3094 515 3095 519
rect 3099 515 3100 519
rect 3094 514 3100 515
rect 3176 512 3178 590
rect 3328 586 3330 597
rect 3326 585 3332 586
rect 3326 581 3327 585
rect 3331 581 3332 585
rect 3326 580 3332 581
rect 3388 572 3390 606
rect 3488 603 3490 618
rect 3520 612 3522 678
rect 3576 675 3578 694
rect 3575 674 3579 675
rect 3575 669 3579 670
rect 3576 654 3578 669
rect 3574 653 3580 654
rect 3574 649 3575 653
rect 3579 649 3580 653
rect 3574 648 3580 649
rect 3546 639 3552 640
rect 3546 635 3547 639
rect 3551 635 3552 639
rect 3546 634 3552 635
rect 3574 636 3580 637
rect 3518 611 3524 612
rect 3518 607 3519 611
rect 3523 607 3524 611
rect 3518 606 3524 607
rect 3487 602 3491 603
rect 3487 597 3491 598
rect 3488 586 3490 597
rect 3548 596 3550 634
rect 3574 632 3575 636
rect 3579 632 3580 636
rect 3574 631 3580 632
rect 3576 603 3578 631
rect 3575 602 3579 603
rect 3575 597 3579 598
rect 3546 595 3552 596
rect 3546 591 3547 595
rect 3551 591 3552 595
rect 3546 590 3552 591
rect 3486 585 3492 586
rect 3486 581 3487 585
rect 3491 581 3492 585
rect 3486 580 3492 581
rect 3576 573 3578 597
rect 3574 572 3580 573
rect 3386 571 3392 572
rect 3386 567 3387 571
rect 3391 567 3392 571
rect 3574 568 3575 572
rect 3579 568 3580 572
rect 3574 567 3580 568
rect 3386 566 3392 567
rect 3574 555 3580 556
rect 3574 551 3575 555
rect 3579 551 3580 555
rect 3574 550 3580 551
rect 3318 545 3324 546
rect 3318 541 3319 545
rect 3323 541 3324 545
rect 3318 540 3324 541
rect 3478 545 3484 546
rect 3478 541 3479 545
rect 3483 541 3484 545
rect 3478 540 3484 541
rect 3320 531 3322 540
rect 3480 531 3482 540
rect 3518 539 3524 540
rect 3518 535 3519 539
rect 3523 535 3524 539
rect 3518 534 3524 535
rect 3223 530 3227 531
rect 3223 525 3227 526
rect 3319 530 3323 531
rect 3319 525 3323 526
rect 3351 530 3355 531
rect 3351 525 3355 526
rect 3479 530 3483 531
rect 3479 525 3483 526
rect 3224 520 3226 525
rect 3352 520 3354 525
rect 3480 520 3482 525
rect 3222 519 3228 520
rect 3222 515 3223 519
rect 3227 515 3228 519
rect 3222 514 3228 515
rect 3350 519 3356 520
rect 3350 515 3351 519
rect 3355 515 3356 519
rect 3350 514 3356 515
rect 3478 519 3484 520
rect 3478 515 3479 519
rect 3483 515 3484 519
rect 3478 514 3484 515
rect 3174 511 3180 512
rect 3174 507 3175 511
rect 3179 507 3180 511
rect 3174 506 3180 507
rect 3290 511 3296 512
rect 3290 507 3291 511
rect 3295 507 3296 511
rect 3290 506 3296 507
rect 2810 495 2816 496
rect 2810 491 2811 495
rect 2815 491 2816 495
rect 2810 490 2816 491
rect 2906 495 2912 496
rect 2906 491 2907 495
rect 2911 491 2912 495
rect 2906 490 2912 491
rect 2812 468 2814 490
rect 2846 479 2852 480
rect 2846 475 2847 479
rect 2851 475 2852 479
rect 2846 474 2852 475
rect 2754 467 2760 468
rect 2754 463 2755 467
rect 2759 463 2760 467
rect 1863 462 1867 463
rect 1671 458 1675 459
rect 1671 453 1675 454
rect 1727 458 1731 459
rect 1727 453 1731 454
rect 1823 458 1827 459
rect 1863 457 1867 458
rect 2239 462 2243 463
rect 2239 457 2243 458
rect 2311 462 2315 463
rect 2311 457 2315 458
rect 2327 462 2331 463
rect 2370 462 2376 463
rect 2407 462 2411 463
rect 2327 457 2331 458
rect 2407 457 2411 458
rect 2431 462 2435 463
rect 2466 462 2472 463
rect 2511 462 2515 463
rect 2431 457 2435 458
rect 2511 457 2515 458
rect 2559 462 2563 463
rect 2570 462 2576 463
rect 2615 462 2619 463
rect 2646 462 2652 463
rect 2695 462 2699 463
rect 2559 457 2563 458
rect 2615 457 2619 458
rect 1823 453 1827 454
rect 1586 451 1592 452
rect 1586 447 1587 451
rect 1591 447 1592 451
rect 1586 446 1592 447
rect 1728 442 1730 453
rect 1390 441 1396 442
rect 1390 437 1391 441
rect 1395 437 1396 441
rect 1390 436 1396 437
rect 1558 441 1564 442
rect 1558 437 1559 441
rect 1563 437 1564 441
rect 1558 436 1564 437
rect 1726 441 1732 442
rect 1726 437 1727 441
rect 1731 437 1732 441
rect 1726 436 1732 437
rect 1824 429 1826 453
rect 1864 433 1866 457
rect 2240 446 2242 457
rect 2270 455 2276 456
rect 2270 451 2271 455
rect 2275 451 2276 455
rect 2270 450 2276 451
rect 2238 445 2244 446
rect 2238 441 2239 445
rect 2243 441 2244 445
rect 2238 440 2244 441
rect 1862 432 1868 433
rect 1822 428 1828 429
rect 1822 424 1823 428
rect 1827 424 1828 428
rect 1862 428 1863 432
rect 1867 428 1868 432
rect 1862 427 1868 428
rect 1290 423 1296 424
rect 1822 423 1828 424
rect 1290 419 1291 423
rect 1295 419 1296 423
rect 1290 418 1296 419
rect 1862 415 1868 416
rect 1298 411 1304 412
rect 1298 407 1299 411
rect 1303 407 1304 411
rect 1298 406 1304 407
rect 1822 411 1828 412
rect 1822 407 1823 411
rect 1827 407 1828 411
rect 1862 411 1863 415
rect 1867 411 1868 415
rect 1862 410 1868 411
rect 1822 406 1828 407
rect 1214 401 1220 402
rect 1214 397 1215 401
rect 1219 397 1220 401
rect 1214 396 1220 397
rect 1216 391 1218 396
rect 1103 390 1107 391
rect 1103 385 1107 386
rect 1215 390 1219 391
rect 1215 385 1219 386
rect 1263 390 1267 391
rect 1263 385 1267 386
rect 1104 380 1106 385
rect 1264 380 1266 385
rect 1102 379 1108 380
rect 1102 375 1103 379
rect 1107 375 1108 379
rect 1102 374 1108 375
rect 1262 379 1268 380
rect 1262 375 1263 379
rect 1267 375 1268 379
rect 1262 374 1268 375
rect 1094 371 1100 372
rect 1094 367 1095 371
rect 1099 367 1100 371
rect 1094 366 1100 367
rect 658 355 664 356
rect 658 351 659 355
rect 663 351 664 355
rect 658 350 664 351
rect 1034 355 1040 356
rect 1034 351 1035 355
rect 1039 351 1040 355
rect 1034 350 1040 351
rect 1254 355 1260 356
rect 1254 351 1255 355
rect 1259 351 1260 355
rect 1254 350 1260 351
rect 598 339 604 340
rect 598 335 599 339
rect 603 335 604 339
rect 598 334 604 335
rect 462 327 468 328
rect 462 323 463 327
rect 467 323 468 327
rect 600 323 602 334
rect 660 328 662 350
rect 774 339 780 340
rect 774 335 775 339
rect 779 335 780 339
rect 774 334 780 335
rect 942 339 948 340
rect 942 335 943 339
rect 947 335 948 339
rect 942 334 948 335
rect 658 327 664 328
rect 658 323 659 327
rect 663 323 664 327
rect 776 323 778 334
rect 782 327 788 328
rect 782 323 783 327
rect 787 323 788 327
rect 944 323 946 334
rect 1036 328 1038 350
rect 1110 339 1116 340
rect 1110 335 1111 339
rect 1115 335 1116 339
rect 1110 334 1116 335
rect 994 327 1000 328
rect 994 323 995 327
rect 999 323 1000 327
rect 271 322 275 323
rect 330 322 336 323
rect 351 322 355 323
rect 271 317 275 318
rect 351 317 355 318
rect 431 322 435 323
rect 462 322 468 323
rect 495 322 499 323
rect 431 317 435 318
rect 495 317 499 318
rect 599 322 603 323
rect 599 317 603 318
rect 639 322 643 323
rect 658 322 664 323
rect 775 322 779 323
rect 782 322 788 323
rect 791 322 795 323
rect 639 317 643 318
rect 775 317 779 318
rect 242 315 248 316
rect 242 311 243 315
rect 247 311 248 315
rect 242 310 248 311
rect 352 306 354 317
rect 496 306 498 317
rect 554 315 560 316
rect 554 311 555 315
rect 559 311 560 315
rect 554 310 560 311
rect 214 305 220 306
rect 214 301 215 305
rect 219 301 220 305
rect 214 300 220 301
rect 350 305 356 306
rect 350 301 351 305
rect 355 301 356 305
rect 350 300 356 301
rect 494 305 500 306
rect 494 301 495 305
rect 499 301 500 305
rect 494 300 500 301
rect 110 292 116 293
rect 110 288 111 292
rect 115 288 116 292
rect 110 287 116 288
rect 110 275 116 276
rect 110 271 111 275
rect 115 271 116 275
rect 110 270 116 271
rect 112 247 114 270
rect 206 265 212 266
rect 206 261 207 265
rect 211 261 212 265
rect 206 260 212 261
rect 342 265 348 266
rect 342 261 343 265
rect 347 261 348 265
rect 342 260 348 261
rect 486 265 492 266
rect 486 261 487 265
rect 491 261 492 265
rect 486 260 492 261
rect 208 247 210 260
rect 344 247 346 260
rect 394 259 400 260
rect 394 255 395 259
rect 399 255 400 259
rect 394 254 400 255
rect 111 246 115 247
rect 111 241 115 242
rect 207 246 211 247
rect 207 241 211 242
rect 231 246 235 247
rect 231 241 235 242
rect 343 246 347 247
rect 343 241 347 242
rect 359 246 363 247
rect 359 241 363 242
rect 112 226 114 241
rect 232 236 234 241
rect 360 236 362 241
rect 230 235 236 236
rect 230 231 231 235
rect 235 231 236 235
rect 230 230 236 231
rect 358 235 364 236
rect 358 231 359 235
rect 363 231 364 235
rect 358 230 364 231
rect 110 225 116 226
rect 110 221 111 225
rect 115 221 116 225
rect 110 220 116 221
rect 206 211 212 212
rect 110 208 116 209
rect 110 204 111 208
rect 115 204 116 208
rect 206 207 207 211
rect 211 207 212 211
rect 206 206 212 207
rect 110 203 116 204
rect 112 155 114 203
rect 111 154 115 155
rect 111 149 115 150
rect 175 154 179 155
rect 175 149 179 150
rect 112 125 114 149
rect 176 138 178 149
rect 208 148 210 206
rect 238 195 244 196
rect 238 191 239 195
rect 243 191 244 195
rect 238 190 244 191
rect 366 195 372 196
rect 366 191 367 195
rect 371 191 372 195
rect 366 190 372 191
rect 240 155 242 190
rect 368 155 370 190
rect 396 184 398 254
rect 488 247 490 260
rect 487 246 491 247
rect 487 241 491 242
rect 488 236 490 241
rect 486 235 492 236
rect 486 231 487 235
rect 491 231 492 235
rect 486 230 492 231
rect 556 228 558 310
rect 640 306 642 317
rect 638 305 644 306
rect 638 301 639 305
rect 643 301 644 305
rect 638 300 644 301
rect 784 288 786 322
rect 791 317 795 318
rect 935 322 939 323
rect 935 317 939 318
rect 943 322 947 323
rect 994 322 1000 323
rect 1034 327 1040 328
rect 1034 323 1035 327
rect 1039 323 1040 327
rect 1112 323 1114 334
rect 1034 322 1040 323
rect 1079 322 1083 323
rect 943 317 947 318
rect 792 306 794 317
rect 936 306 938 317
rect 790 305 796 306
rect 790 301 791 305
rect 795 301 796 305
rect 790 300 796 301
rect 934 305 940 306
rect 934 301 935 305
rect 939 301 940 305
rect 934 300 940 301
rect 996 292 998 322
rect 1079 317 1083 318
rect 1111 322 1115 323
rect 1111 317 1115 318
rect 1223 322 1227 323
rect 1223 317 1227 318
rect 1080 306 1082 317
rect 1098 315 1104 316
rect 1098 311 1099 315
rect 1103 311 1104 315
rect 1098 310 1104 311
rect 1078 305 1084 306
rect 1078 301 1079 305
rect 1083 301 1084 305
rect 1078 300 1084 301
rect 994 291 1000 292
rect 782 287 788 288
rect 782 283 783 287
rect 787 283 788 287
rect 994 287 995 291
rect 999 287 1000 291
rect 994 286 1000 287
rect 782 282 788 283
rect 630 265 636 266
rect 630 261 631 265
rect 635 261 636 265
rect 630 260 636 261
rect 782 265 788 266
rect 782 261 783 265
rect 787 261 788 265
rect 782 260 788 261
rect 926 265 932 266
rect 926 261 927 265
rect 931 261 932 265
rect 926 260 932 261
rect 1070 265 1076 266
rect 1070 261 1071 265
rect 1075 261 1076 265
rect 1070 260 1076 261
rect 632 247 634 260
rect 784 247 786 260
rect 928 247 930 260
rect 1072 247 1074 260
rect 623 246 627 247
rect 623 241 627 242
rect 631 246 635 247
rect 631 241 635 242
rect 759 246 763 247
rect 759 241 763 242
rect 783 246 787 247
rect 783 241 787 242
rect 895 246 899 247
rect 895 241 899 242
rect 927 246 931 247
rect 927 241 931 242
rect 1031 246 1035 247
rect 1031 241 1035 242
rect 1071 246 1075 247
rect 1071 241 1075 242
rect 624 236 626 241
rect 760 236 762 241
rect 896 236 898 241
rect 1032 236 1034 241
rect 622 235 628 236
rect 622 231 623 235
rect 627 231 628 235
rect 622 230 628 231
rect 758 235 764 236
rect 758 231 759 235
rect 763 231 764 235
rect 758 230 764 231
rect 894 235 900 236
rect 894 231 895 235
rect 899 231 900 235
rect 894 230 900 231
rect 1030 235 1036 236
rect 1030 231 1031 235
rect 1035 231 1036 235
rect 1030 230 1036 231
rect 1100 228 1102 310
rect 1224 306 1226 317
rect 1256 316 1258 350
rect 1270 339 1276 340
rect 1270 335 1271 339
rect 1275 335 1276 339
rect 1270 334 1276 335
rect 1272 323 1274 334
rect 1300 328 1302 406
rect 1382 401 1388 402
rect 1382 397 1383 401
rect 1387 397 1388 401
rect 1382 396 1388 397
rect 1550 401 1556 402
rect 1550 397 1551 401
rect 1555 397 1556 401
rect 1550 396 1556 397
rect 1718 401 1724 402
rect 1718 397 1719 401
rect 1723 397 1724 401
rect 1718 396 1724 397
rect 1384 391 1386 396
rect 1552 391 1554 396
rect 1720 391 1722 396
rect 1766 395 1772 396
rect 1766 391 1767 395
rect 1771 391 1772 395
rect 1824 391 1826 406
rect 1864 395 1866 410
rect 2230 405 2236 406
rect 2230 401 2231 405
rect 2235 401 2236 405
rect 2230 400 2236 401
rect 2232 395 2234 400
rect 1863 394 1867 395
rect 1383 390 1387 391
rect 1383 385 1387 386
rect 1423 390 1427 391
rect 1423 385 1427 386
rect 1551 390 1555 391
rect 1551 385 1555 386
rect 1583 390 1587 391
rect 1583 385 1587 386
rect 1719 390 1723 391
rect 1719 385 1723 386
rect 1727 390 1731 391
rect 1766 390 1772 391
rect 1823 390 1827 391
rect 1727 385 1731 386
rect 1424 380 1426 385
rect 1584 380 1586 385
rect 1728 380 1730 385
rect 1422 379 1428 380
rect 1422 375 1423 379
rect 1427 375 1428 379
rect 1422 374 1428 375
rect 1582 379 1588 380
rect 1582 375 1583 379
rect 1587 375 1588 379
rect 1582 374 1588 375
rect 1726 379 1732 380
rect 1726 375 1727 379
rect 1731 375 1732 379
rect 1726 374 1732 375
rect 1650 355 1656 356
rect 1650 351 1651 355
rect 1655 351 1656 355
rect 1650 350 1656 351
rect 1658 355 1664 356
rect 1658 351 1659 355
rect 1663 351 1664 355
rect 1658 350 1664 351
rect 1430 339 1436 340
rect 1430 335 1431 339
rect 1435 335 1436 339
rect 1430 334 1436 335
rect 1590 339 1596 340
rect 1590 335 1591 339
rect 1595 335 1596 339
rect 1590 334 1596 335
rect 1298 327 1304 328
rect 1298 323 1299 327
rect 1303 323 1304 327
rect 1432 323 1434 334
rect 1592 323 1594 334
rect 1271 322 1275 323
rect 1298 322 1304 323
rect 1359 322 1363 323
rect 1271 317 1275 318
rect 1359 317 1363 318
rect 1431 322 1435 323
rect 1431 317 1435 318
rect 1487 322 1491 323
rect 1487 317 1491 318
rect 1591 322 1595 323
rect 1591 317 1595 318
rect 1623 322 1627 323
rect 1623 317 1627 318
rect 1254 315 1260 316
rect 1254 311 1255 315
rect 1259 311 1260 315
rect 1254 310 1260 311
rect 1360 306 1362 317
rect 1488 306 1490 317
rect 1624 306 1626 317
rect 1652 316 1654 350
rect 1660 336 1662 350
rect 1734 339 1740 340
rect 1658 335 1664 336
rect 1658 331 1659 335
rect 1663 331 1664 335
rect 1734 335 1735 339
rect 1739 335 1740 339
rect 1734 334 1740 335
rect 1658 330 1664 331
rect 1736 323 1738 334
rect 1768 328 1770 390
rect 1863 389 1867 390
rect 2183 394 2187 395
rect 2183 389 2187 390
rect 2231 394 2235 395
rect 2272 392 2274 450
rect 2328 446 2330 457
rect 2432 446 2434 457
rect 2560 446 2562 457
rect 2326 445 2332 446
rect 2326 441 2327 445
rect 2331 441 2332 445
rect 2326 440 2332 441
rect 2430 445 2436 446
rect 2430 441 2431 445
rect 2435 441 2436 445
rect 2430 440 2436 441
rect 2558 445 2564 446
rect 2558 441 2559 445
rect 2563 441 2564 445
rect 2558 440 2564 441
rect 2648 428 2650 462
rect 2695 457 2699 458
rect 2727 462 2731 463
rect 2754 462 2760 463
rect 2810 467 2816 468
rect 2810 463 2811 467
rect 2815 463 2816 467
rect 2848 463 2850 474
rect 2810 462 2816 463
rect 2847 462 2851 463
rect 2727 457 2731 458
rect 2847 457 2851 458
rect 2696 446 2698 457
rect 2848 446 2850 457
rect 2908 456 2910 490
rect 2974 479 2980 480
rect 2974 475 2975 479
rect 2979 475 2980 479
rect 3102 479 3108 480
rect 2974 474 2980 475
rect 3007 476 3011 477
rect 2976 463 2978 474
rect 3102 475 3103 479
rect 3107 475 3108 479
rect 3102 474 3108 475
rect 3230 479 3236 480
rect 3230 475 3231 479
rect 3235 475 3236 479
rect 3292 477 3294 506
rect 3358 479 3364 480
rect 3230 474 3236 475
rect 3291 476 3295 477
rect 3007 471 3011 472
rect 3008 468 3010 471
rect 3006 467 3012 468
rect 3006 463 3007 467
rect 3011 463 3012 467
rect 3104 463 3106 474
rect 3218 467 3224 468
rect 3218 463 3219 467
rect 3223 463 3224 467
rect 3232 463 3234 474
rect 3358 475 3359 479
rect 3363 475 3364 479
rect 3358 474 3364 475
rect 3486 479 3492 480
rect 3486 475 3487 479
rect 3491 475 3492 479
rect 3486 474 3492 475
rect 3291 471 3295 472
rect 3360 463 3362 474
rect 3488 463 3490 474
rect 3520 468 3522 534
rect 3576 531 3578 550
rect 3575 530 3579 531
rect 3575 525 3579 526
rect 3576 510 3578 525
rect 3574 509 3580 510
rect 3574 505 3575 509
rect 3579 505 3580 509
rect 3574 504 3580 505
rect 3546 495 3552 496
rect 3546 491 3547 495
rect 3551 491 3552 495
rect 3546 490 3552 491
rect 3574 492 3580 493
rect 3518 467 3524 468
rect 3518 463 3519 467
rect 3523 463 3524 467
rect 2975 462 2979 463
rect 2975 457 2979 458
rect 2999 462 3003 463
rect 3006 462 3012 463
rect 3103 462 3107 463
rect 2999 457 3003 458
rect 3103 457 3107 458
rect 3159 462 3163 463
rect 3218 462 3224 463
rect 3231 462 3235 463
rect 3159 457 3163 458
rect 2906 455 2912 456
rect 2906 451 2907 455
rect 2911 451 2912 455
rect 2906 450 2912 451
rect 3000 446 3002 457
rect 3160 446 3162 457
rect 2694 445 2700 446
rect 2694 441 2695 445
rect 2699 441 2700 445
rect 2694 440 2700 441
rect 2846 445 2852 446
rect 2846 441 2847 445
rect 2851 441 2852 445
rect 2846 440 2852 441
rect 2998 445 3004 446
rect 2998 441 2999 445
rect 3003 441 3004 445
rect 2998 440 3004 441
rect 3158 445 3164 446
rect 3158 441 3159 445
rect 3163 441 3164 445
rect 3158 440 3164 441
rect 3220 432 3222 462
rect 3231 457 3235 458
rect 3327 462 3331 463
rect 3327 457 3331 458
rect 3359 462 3363 463
rect 3359 457 3363 458
rect 3487 462 3491 463
rect 3518 462 3524 463
rect 3487 457 3491 458
rect 3262 455 3268 456
rect 3262 451 3263 455
rect 3267 451 3268 455
rect 3262 450 3268 451
rect 3218 431 3224 432
rect 2646 427 2652 428
rect 2646 423 2647 427
rect 2651 423 2652 427
rect 3218 427 3219 431
rect 3223 427 3224 431
rect 3264 428 3266 450
rect 3328 446 3330 457
rect 3488 446 3490 457
rect 3548 456 3550 490
rect 3574 488 3575 492
rect 3579 488 3580 492
rect 3574 487 3580 488
rect 3576 463 3578 487
rect 3575 462 3579 463
rect 3575 457 3579 458
rect 3546 455 3552 456
rect 3546 451 3547 455
rect 3551 451 3552 455
rect 3546 450 3552 451
rect 3326 445 3332 446
rect 3326 441 3327 445
rect 3331 441 3332 445
rect 3326 440 3332 441
rect 3486 445 3492 446
rect 3486 441 3487 445
rect 3491 441 3492 445
rect 3486 440 3492 441
rect 3576 433 3578 457
rect 3574 432 3580 433
rect 3574 428 3575 432
rect 3579 428 3580 432
rect 3218 426 3224 427
rect 3262 427 3268 428
rect 3574 427 3580 428
rect 2646 422 2652 423
rect 3262 423 3263 427
rect 3267 423 3268 427
rect 3262 422 3268 423
rect 2998 415 3004 416
rect 2998 411 2999 415
rect 3003 411 3004 415
rect 2998 410 3004 411
rect 3574 415 3580 416
rect 3574 411 3575 415
rect 3579 411 3580 415
rect 3574 410 3580 411
rect 2318 405 2324 406
rect 2318 401 2319 405
rect 2323 401 2324 405
rect 2318 400 2324 401
rect 2422 405 2428 406
rect 2422 401 2423 405
rect 2427 401 2428 405
rect 2422 400 2428 401
rect 2550 405 2556 406
rect 2550 401 2551 405
rect 2555 401 2556 405
rect 2550 400 2556 401
rect 2686 405 2692 406
rect 2686 401 2687 405
rect 2691 401 2692 405
rect 2686 400 2692 401
rect 2838 405 2844 406
rect 2838 401 2839 405
rect 2843 401 2844 405
rect 2838 400 2844 401
rect 2990 405 2996 406
rect 2990 401 2991 405
rect 2995 401 2996 405
rect 2990 400 2996 401
rect 2320 395 2322 400
rect 2424 395 2426 400
rect 2552 395 2554 400
rect 2688 395 2690 400
rect 2840 395 2842 400
rect 2992 395 2994 400
rect 2287 394 2291 395
rect 2231 389 2235 390
rect 2270 391 2276 392
rect 1823 385 1827 386
rect 1824 370 1826 385
rect 1864 374 1866 389
rect 2184 384 2186 389
rect 2270 387 2271 391
rect 2275 387 2276 391
rect 2287 389 2291 390
rect 2319 394 2323 395
rect 2319 389 2323 390
rect 2399 394 2403 395
rect 2399 389 2403 390
rect 2423 394 2427 395
rect 2423 389 2427 390
rect 2527 394 2531 395
rect 2527 389 2531 390
rect 2551 394 2555 395
rect 2551 389 2555 390
rect 2671 394 2675 395
rect 2671 389 2675 390
rect 2687 394 2691 395
rect 2687 389 2691 390
rect 2815 394 2819 395
rect 2815 389 2819 390
rect 2839 394 2843 395
rect 2839 389 2843 390
rect 2967 394 2971 395
rect 2967 389 2971 390
rect 2991 394 2995 395
rect 2991 389 2995 390
rect 2270 386 2276 387
rect 2288 384 2290 389
rect 2400 384 2402 389
rect 2528 384 2530 389
rect 2672 384 2674 389
rect 2816 384 2818 389
rect 2968 384 2970 389
rect 2182 383 2188 384
rect 2182 379 2183 383
rect 2187 379 2188 383
rect 2182 378 2188 379
rect 2286 383 2292 384
rect 2286 379 2287 383
rect 2291 379 2292 383
rect 2286 378 2292 379
rect 2398 383 2404 384
rect 2398 379 2399 383
rect 2403 379 2404 383
rect 2398 378 2404 379
rect 2526 383 2532 384
rect 2526 379 2527 383
rect 2531 379 2532 383
rect 2526 378 2532 379
rect 2670 383 2676 384
rect 2670 379 2671 383
rect 2675 379 2676 383
rect 2670 378 2676 379
rect 2814 383 2820 384
rect 2814 379 2815 383
rect 2819 379 2820 383
rect 2814 378 2820 379
rect 2966 383 2972 384
rect 2966 379 2967 383
rect 2971 379 2972 383
rect 2966 378 2972 379
rect 1862 373 1868 374
rect 1822 369 1828 370
rect 1822 365 1823 369
rect 1827 365 1828 369
rect 1862 369 1863 373
rect 1867 369 1868 373
rect 1862 368 1868 369
rect 1822 364 1828 365
rect 2594 359 2600 360
rect 1862 356 1868 357
rect 1822 352 1828 353
rect 1822 348 1823 352
rect 1827 348 1828 352
rect 1862 352 1863 356
rect 1867 352 1868 356
rect 2594 355 2595 359
rect 2599 355 2600 359
rect 2594 354 2600 355
rect 2882 359 2888 360
rect 2882 355 2883 359
rect 2887 355 2888 359
rect 2882 354 2888 355
rect 1862 351 1868 352
rect 1822 347 1828 348
rect 1766 327 1772 328
rect 1766 323 1767 327
rect 1771 323 1772 327
rect 1824 323 1826 347
rect 1735 322 1739 323
rect 1766 322 1772 323
rect 1823 322 1827 323
rect 1735 317 1739 318
rect 1864 319 1866 351
rect 2190 343 2196 344
rect 2190 339 2191 343
rect 2195 339 2196 343
rect 2190 338 2196 339
rect 2294 343 2300 344
rect 2294 339 2295 343
rect 2299 339 2300 343
rect 2294 338 2300 339
rect 2406 343 2412 344
rect 2406 339 2407 343
rect 2411 339 2412 343
rect 2406 338 2412 339
rect 2534 343 2540 344
rect 2534 339 2535 343
rect 2539 339 2540 343
rect 2534 338 2540 339
rect 2192 319 2194 338
rect 2296 319 2298 338
rect 2408 319 2410 338
rect 2536 319 2538 338
rect 1823 317 1827 318
rect 1863 318 1867 319
rect 1650 315 1656 316
rect 1650 311 1651 315
rect 1655 311 1656 315
rect 1650 310 1656 311
rect 1736 306 1738 317
rect 1222 305 1228 306
rect 1222 301 1223 305
rect 1227 301 1228 305
rect 1222 300 1228 301
rect 1358 305 1364 306
rect 1358 301 1359 305
rect 1363 301 1364 305
rect 1358 300 1364 301
rect 1486 305 1492 306
rect 1486 301 1487 305
rect 1491 301 1492 305
rect 1486 300 1492 301
rect 1622 305 1628 306
rect 1622 301 1623 305
rect 1627 301 1628 305
rect 1622 300 1628 301
rect 1734 305 1740 306
rect 1734 301 1735 305
rect 1739 301 1740 305
rect 1734 300 1740 301
rect 1824 293 1826 317
rect 1863 313 1867 314
rect 1895 318 1899 319
rect 1895 313 1899 314
rect 2087 318 2091 319
rect 2087 313 2091 314
rect 2191 318 2195 319
rect 2191 313 2195 314
rect 2295 318 2299 319
rect 2295 313 2299 314
rect 2303 318 2307 319
rect 2303 313 2307 314
rect 2407 318 2411 319
rect 2407 313 2411 314
rect 2511 318 2515 319
rect 2511 313 2515 314
rect 2535 318 2539 319
rect 2535 313 2539 314
rect 1822 292 1828 293
rect 1822 288 1823 292
rect 1827 288 1828 292
rect 1864 289 1866 313
rect 1896 302 1898 313
rect 2088 302 2090 313
rect 2154 311 2160 312
rect 2154 307 2155 311
rect 2159 307 2160 311
rect 2154 306 2160 307
rect 1894 301 1900 302
rect 1894 297 1895 301
rect 1899 297 1900 301
rect 1894 296 1900 297
rect 2086 301 2092 302
rect 2086 297 2087 301
rect 2091 297 2092 301
rect 2086 296 2092 297
rect 1822 287 1828 288
rect 1862 288 1868 289
rect 1862 284 1863 288
rect 1867 284 1868 288
rect 2156 284 2158 306
rect 2304 302 2306 313
rect 2362 311 2368 312
rect 2362 307 2363 311
rect 2367 307 2368 311
rect 2362 306 2368 307
rect 2302 301 2308 302
rect 2302 297 2303 301
rect 2307 297 2308 301
rect 2302 296 2308 297
rect 1862 283 1868 284
rect 2154 283 2160 284
rect 2154 279 2155 283
rect 2159 279 2160 283
rect 2154 278 2160 279
rect 1470 275 1476 276
rect 1470 271 1471 275
rect 1475 271 1476 275
rect 1470 270 1476 271
rect 1822 275 1828 276
rect 1822 271 1823 275
rect 1827 271 1828 275
rect 1822 270 1828 271
rect 1862 271 1868 272
rect 1214 265 1220 266
rect 1214 261 1215 265
rect 1219 261 1220 265
rect 1214 260 1220 261
rect 1350 265 1356 266
rect 1350 261 1351 265
rect 1355 261 1356 265
rect 1350 260 1356 261
rect 1216 247 1218 260
rect 1352 247 1354 260
rect 1159 246 1163 247
rect 1159 241 1163 242
rect 1215 246 1219 247
rect 1215 241 1219 242
rect 1295 246 1299 247
rect 1295 241 1299 242
rect 1351 246 1355 247
rect 1351 241 1355 242
rect 1431 246 1435 247
rect 1431 241 1435 242
rect 1160 236 1162 241
rect 1296 236 1298 241
rect 1432 236 1434 241
rect 1158 235 1164 236
rect 1158 231 1159 235
rect 1163 231 1164 235
rect 1158 230 1164 231
rect 1294 235 1300 236
rect 1294 231 1295 235
rect 1299 231 1300 235
rect 1294 230 1300 231
rect 1430 235 1436 236
rect 1430 231 1431 235
rect 1435 231 1436 235
rect 1430 230 1436 231
rect 426 227 432 228
rect 426 223 427 227
rect 431 223 432 227
rect 426 222 432 223
rect 554 227 560 228
rect 554 223 555 227
rect 559 223 560 227
rect 554 222 560 223
rect 1098 227 1104 228
rect 1098 223 1099 227
rect 1103 223 1104 227
rect 1098 222 1104 223
rect 428 192 430 222
rect 690 211 696 212
rect 690 207 691 211
rect 695 207 696 211
rect 690 206 696 207
rect 1362 211 1368 212
rect 1362 207 1363 211
rect 1367 207 1368 211
rect 1362 206 1368 207
rect 1370 211 1376 212
rect 1370 207 1371 211
rect 1375 207 1376 211
rect 1370 206 1376 207
rect 494 195 500 196
rect 426 191 432 192
rect 426 187 427 191
rect 431 187 432 191
rect 494 191 495 195
rect 499 191 500 195
rect 494 190 500 191
rect 630 195 636 196
rect 630 191 631 195
rect 635 191 636 195
rect 630 190 636 191
rect 426 186 432 187
rect 394 183 400 184
rect 394 179 395 183
rect 399 179 400 183
rect 394 178 400 179
rect 496 155 498 190
rect 632 155 634 190
rect 692 184 694 206
rect 766 195 772 196
rect 766 191 767 195
rect 771 191 772 195
rect 766 190 772 191
rect 902 195 908 196
rect 902 191 903 195
rect 907 191 908 195
rect 902 190 908 191
rect 1038 195 1044 196
rect 1038 191 1039 195
rect 1043 191 1044 195
rect 1038 190 1044 191
rect 1166 195 1172 196
rect 1166 191 1167 195
rect 1171 191 1172 195
rect 1166 190 1172 191
rect 1302 195 1308 196
rect 1302 191 1303 195
rect 1307 191 1308 195
rect 1302 190 1308 191
rect 690 183 696 184
rect 690 179 691 183
rect 695 179 696 183
rect 690 178 696 179
rect 768 155 770 190
rect 782 183 788 184
rect 782 179 783 183
rect 787 179 788 183
rect 782 178 788 179
rect 239 154 243 155
rect 239 149 243 150
rect 263 154 267 155
rect 263 149 267 150
rect 351 154 355 155
rect 351 149 355 150
rect 367 154 371 155
rect 367 149 371 150
rect 439 154 443 155
rect 439 149 443 150
rect 495 154 499 155
rect 495 149 499 150
rect 527 154 531 155
rect 527 149 531 150
rect 615 154 619 155
rect 615 149 619 150
rect 631 154 635 155
rect 631 149 635 150
rect 703 154 707 155
rect 703 149 707 150
rect 767 154 771 155
rect 767 149 771 150
rect 206 147 212 148
rect 206 143 207 147
rect 211 143 212 147
rect 206 142 212 143
rect 264 138 266 149
rect 352 138 354 149
rect 440 138 442 149
rect 528 138 530 149
rect 616 138 618 149
rect 704 138 706 149
rect 174 137 180 138
rect 174 133 175 137
rect 179 133 180 137
rect 174 132 180 133
rect 262 137 268 138
rect 262 133 263 137
rect 267 133 268 137
rect 262 132 268 133
rect 350 137 356 138
rect 350 133 351 137
rect 355 133 356 137
rect 350 132 356 133
rect 438 137 444 138
rect 438 133 439 137
rect 443 133 444 137
rect 438 132 444 133
rect 526 137 532 138
rect 526 133 527 137
rect 531 133 532 137
rect 526 132 532 133
rect 614 137 620 138
rect 614 133 615 137
rect 619 133 620 137
rect 614 132 620 133
rect 702 137 708 138
rect 702 133 703 137
rect 707 133 708 137
rect 702 132 708 133
rect 110 124 116 125
rect 110 120 111 124
rect 115 120 116 124
rect 784 120 786 178
rect 904 155 906 190
rect 934 183 940 184
rect 934 179 935 183
rect 939 179 940 183
rect 934 178 940 179
rect 791 154 795 155
rect 791 149 795 150
rect 879 154 883 155
rect 879 149 883 150
rect 903 154 907 155
rect 903 149 907 150
rect 792 138 794 149
rect 880 138 882 149
rect 790 137 796 138
rect 790 133 791 137
rect 795 133 796 137
rect 790 132 796 133
rect 878 137 884 138
rect 878 133 879 137
rect 883 133 884 137
rect 878 132 884 133
rect 936 132 938 178
rect 1040 155 1042 190
rect 1168 155 1170 190
rect 1304 155 1306 190
rect 967 154 971 155
rect 967 149 971 150
rect 1039 154 1043 155
rect 1039 149 1043 150
rect 1055 154 1059 155
rect 1055 149 1059 150
rect 1143 154 1147 155
rect 1143 149 1147 150
rect 1167 154 1171 155
rect 1167 149 1171 150
rect 1231 154 1235 155
rect 1231 149 1235 150
rect 1303 154 1307 155
rect 1303 149 1307 150
rect 1319 154 1323 155
rect 1319 149 1323 150
rect 946 147 952 148
rect 946 143 947 147
rect 951 143 952 147
rect 946 142 952 143
rect 934 131 940 132
rect 934 127 935 131
rect 939 127 940 131
rect 934 126 940 127
rect 948 120 950 142
rect 968 138 970 149
rect 1056 138 1058 149
rect 1122 147 1128 148
rect 1122 143 1123 147
rect 1127 143 1128 147
rect 1122 142 1128 143
rect 966 137 972 138
rect 966 133 967 137
rect 971 133 972 137
rect 966 132 972 133
rect 1054 137 1060 138
rect 1054 133 1055 137
rect 1059 133 1060 137
rect 1054 132 1060 133
rect 1124 120 1126 142
rect 1144 138 1146 149
rect 1210 147 1216 148
rect 1210 143 1211 147
rect 1215 143 1216 147
rect 1210 142 1216 143
rect 1142 137 1148 138
rect 1142 133 1143 137
rect 1147 133 1148 137
rect 1142 132 1148 133
rect 1212 120 1214 142
rect 1232 138 1234 149
rect 1320 138 1322 149
rect 1364 148 1366 206
rect 1372 176 1374 206
rect 1438 195 1444 196
rect 1438 191 1439 195
rect 1443 191 1444 195
rect 1438 190 1444 191
rect 1370 175 1376 176
rect 1370 171 1371 175
rect 1375 171 1376 175
rect 1370 170 1376 171
rect 1440 155 1442 190
rect 1472 184 1474 270
rect 1478 265 1484 266
rect 1478 261 1479 265
rect 1483 261 1484 265
rect 1478 260 1484 261
rect 1614 265 1620 266
rect 1614 261 1615 265
rect 1619 261 1620 265
rect 1614 260 1620 261
rect 1726 265 1732 266
rect 1726 261 1727 265
rect 1731 261 1732 265
rect 1726 260 1732 261
rect 1480 247 1482 260
rect 1616 247 1618 260
rect 1728 247 1730 260
rect 1824 247 1826 270
rect 1862 267 1863 271
rect 1867 267 1868 271
rect 1862 266 1868 267
rect 1864 251 1866 266
rect 1886 261 1892 262
rect 1886 257 1887 261
rect 1891 257 1892 261
rect 1886 256 1892 257
rect 2078 261 2084 262
rect 2078 257 2079 261
rect 2083 257 2084 261
rect 2078 256 2084 257
rect 2294 261 2300 262
rect 2294 257 2295 261
rect 2299 257 2300 261
rect 2294 256 2300 257
rect 1888 251 1890 256
rect 1926 255 1932 256
rect 1926 251 1927 255
rect 1931 251 1932 255
rect 2080 251 2082 256
rect 2296 251 2298 256
rect 1863 250 1867 251
rect 1479 246 1483 247
rect 1479 241 1483 242
rect 1615 246 1619 247
rect 1615 241 1619 242
rect 1727 246 1731 247
rect 1727 241 1731 242
rect 1823 246 1827 247
rect 1863 245 1867 246
rect 1887 250 1891 251
rect 1926 250 1932 251
rect 1999 250 2003 251
rect 1887 245 1891 246
rect 1823 241 1827 242
rect 1824 226 1826 241
rect 1864 230 1866 245
rect 1888 240 1890 245
rect 1886 239 1892 240
rect 1886 235 1887 239
rect 1891 235 1892 239
rect 1886 234 1892 235
rect 1862 229 1868 230
rect 1822 225 1828 226
rect 1822 221 1823 225
rect 1827 221 1828 225
rect 1862 225 1863 229
rect 1867 225 1868 229
rect 1862 224 1868 225
rect 1822 220 1828 221
rect 1862 212 1868 213
rect 1822 208 1828 209
rect 1822 204 1823 208
rect 1827 204 1828 208
rect 1862 208 1863 212
rect 1867 208 1868 212
rect 1862 207 1868 208
rect 1822 203 1828 204
rect 1470 183 1476 184
rect 1470 179 1471 183
rect 1475 179 1476 183
rect 1470 178 1476 179
rect 1824 155 1826 203
rect 1864 155 1866 207
rect 1894 199 1900 200
rect 1894 195 1895 199
rect 1899 195 1900 199
rect 1894 194 1900 195
rect 1896 155 1898 194
rect 1928 188 1930 250
rect 1999 245 2003 246
rect 2079 250 2083 251
rect 2079 245 2083 246
rect 2143 250 2147 251
rect 2143 245 2147 246
rect 2295 250 2299 251
rect 2295 245 2299 246
rect 2000 240 2002 245
rect 2144 240 2146 245
rect 2296 240 2298 245
rect 1998 239 2004 240
rect 1998 235 1999 239
rect 2003 235 2004 239
rect 1998 234 2004 235
rect 2142 239 2148 240
rect 2142 235 2143 239
rect 2147 235 2148 239
rect 2142 234 2148 235
rect 2294 239 2300 240
rect 2294 235 2295 239
rect 2299 235 2300 239
rect 2294 234 2300 235
rect 2364 232 2366 306
rect 2512 302 2514 313
rect 2596 312 2598 354
rect 2678 343 2684 344
rect 2678 339 2679 343
rect 2683 339 2684 343
rect 2678 338 2684 339
rect 2822 343 2828 344
rect 2822 339 2823 343
rect 2827 339 2828 343
rect 2822 338 2828 339
rect 2680 319 2682 338
rect 2824 319 2826 338
rect 2884 332 2886 354
rect 2974 343 2980 344
rect 2974 339 2975 343
rect 2979 339 2980 343
rect 2974 338 2980 339
rect 2882 331 2888 332
rect 2882 327 2883 331
rect 2887 327 2888 331
rect 2882 326 2888 327
rect 2976 319 2978 338
rect 3000 332 3002 410
rect 3150 405 3156 406
rect 3150 401 3151 405
rect 3155 401 3156 405
rect 3150 400 3156 401
rect 3318 405 3324 406
rect 3318 401 3319 405
rect 3323 401 3324 405
rect 3318 400 3324 401
rect 3478 405 3484 406
rect 3478 401 3479 405
rect 3483 401 3484 405
rect 3478 400 3484 401
rect 3152 395 3154 400
rect 3320 395 3322 400
rect 3480 395 3482 400
rect 3518 399 3524 400
rect 3518 395 3519 399
rect 3523 395 3524 399
rect 3576 395 3578 410
rect 3127 394 3131 395
rect 3127 389 3131 390
rect 3151 394 3155 395
rect 3151 389 3155 390
rect 3295 394 3299 395
rect 3295 389 3299 390
rect 3319 394 3323 395
rect 3319 389 3323 390
rect 3463 394 3467 395
rect 3463 389 3467 390
rect 3479 394 3483 395
rect 3518 394 3524 395
rect 3575 394 3579 395
rect 3479 389 3483 390
rect 3128 384 3130 389
rect 3296 384 3298 389
rect 3464 384 3466 389
rect 3126 383 3132 384
rect 3126 379 3127 383
rect 3131 379 3132 383
rect 3126 378 3132 379
rect 3294 383 3300 384
rect 3294 379 3295 383
rect 3299 379 3300 383
rect 3294 378 3300 379
rect 3462 383 3468 384
rect 3462 379 3463 383
rect 3467 379 3468 383
rect 3462 378 3468 379
rect 3134 343 3140 344
rect 3134 339 3135 343
rect 3139 339 3140 343
rect 3134 338 3140 339
rect 3302 343 3308 344
rect 3302 339 3303 343
rect 3307 339 3308 343
rect 3302 338 3308 339
rect 3470 343 3476 344
rect 3470 339 3471 343
rect 3475 339 3476 343
rect 3470 338 3476 339
rect 2998 331 3004 332
rect 2998 327 2999 331
rect 3003 327 3004 331
rect 2998 326 3004 327
rect 3136 319 3138 338
rect 3154 331 3160 332
rect 3154 327 3155 331
rect 3159 327 3160 331
rect 3154 326 3160 327
rect 2679 318 2683 319
rect 2679 313 2683 314
rect 2711 318 2715 319
rect 2711 313 2715 314
rect 2823 318 2827 319
rect 2823 313 2827 314
rect 2903 318 2907 319
rect 2903 313 2907 314
rect 2975 318 2979 319
rect 2975 313 2979 314
rect 3095 318 3099 319
rect 3095 313 3099 314
rect 3135 318 3139 319
rect 3135 313 3139 314
rect 2594 311 2600 312
rect 2594 307 2595 311
rect 2599 307 2600 311
rect 2594 306 2600 307
rect 2712 302 2714 313
rect 2854 311 2860 312
rect 2854 307 2855 311
rect 2859 307 2860 311
rect 2854 306 2860 307
rect 2510 301 2516 302
rect 2510 297 2511 301
rect 2515 297 2516 301
rect 2510 296 2516 297
rect 2710 301 2716 302
rect 2710 297 2711 301
rect 2715 297 2716 301
rect 2710 296 2716 297
rect 2856 288 2858 306
rect 2904 302 2906 313
rect 3096 302 3098 313
rect 2902 301 2908 302
rect 2902 297 2903 301
rect 2907 297 2908 301
rect 2902 296 2908 297
rect 3094 301 3100 302
rect 3094 297 3095 301
rect 3099 297 3100 301
rect 3094 296 3100 297
rect 3156 288 3158 326
rect 3304 319 3306 338
rect 3472 319 3474 338
rect 3295 318 3299 319
rect 3295 313 3299 314
rect 3303 318 3307 319
rect 3303 313 3307 314
rect 3471 318 3475 319
rect 3471 313 3475 314
rect 3487 318 3491 319
rect 3487 313 3491 314
rect 3238 311 3244 312
rect 3238 307 3239 311
rect 3243 307 3244 311
rect 3238 306 3244 307
rect 2854 287 2860 288
rect 2854 283 2855 287
rect 2859 283 2860 287
rect 2854 282 2860 283
rect 3154 287 3160 288
rect 3154 283 3155 287
rect 3159 283 3160 287
rect 3154 282 3160 283
rect 2986 271 2992 272
rect 2986 267 2987 271
rect 2991 267 2992 271
rect 2986 266 2992 267
rect 2502 261 2508 262
rect 2502 257 2503 261
rect 2507 257 2508 261
rect 2502 256 2508 257
rect 2702 261 2708 262
rect 2702 257 2703 261
rect 2707 257 2708 261
rect 2702 256 2708 257
rect 2894 261 2900 262
rect 2894 257 2895 261
rect 2899 257 2900 261
rect 2894 256 2900 257
rect 2504 251 2506 256
rect 2704 251 2706 256
rect 2896 251 2898 256
rect 2455 250 2459 251
rect 2455 245 2459 246
rect 2503 250 2507 251
rect 2503 245 2507 246
rect 2615 250 2619 251
rect 2615 245 2619 246
rect 2703 250 2707 251
rect 2703 245 2707 246
rect 2783 250 2787 251
rect 2783 245 2787 246
rect 2895 250 2899 251
rect 2895 245 2899 246
rect 2951 250 2955 251
rect 2951 245 2955 246
rect 2456 240 2458 245
rect 2616 240 2618 245
rect 2784 240 2786 245
rect 2952 240 2954 245
rect 2454 239 2460 240
rect 2454 235 2455 239
rect 2459 235 2460 239
rect 2454 234 2460 235
rect 2614 239 2620 240
rect 2614 235 2615 239
rect 2619 235 2620 239
rect 2614 234 2620 235
rect 2782 239 2788 240
rect 2782 235 2783 239
rect 2787 235 2788 239
rect 2782 234 2788 235
rect 2950 239 2956 240
rect 2950 235 2951 239
rect 2955 235 2956 239
rect 2950 234 2956 235
rect 2078 231 2084 232
rect 2078 227 2079 231
rect 2083 227 2084 231
rect 2078 226 2084 227
rect 2362 231 2368 232
rect 2362 227 2363 231
rect 2367 227 2368 231
rect 2362 226 2368 227
rect 2006 199 2012 200
rect 2006 195 2007 199
rect 2011 195 2012 199
rect 2006 194 2012 195
rect 1926 187 1932 188
rect 1926 183 1927 187
rect 1931 183 1932 187
rect 1926 182 1932 183
rect 2008 155 2010 194
rect 2080 156 2082 226
rect 2362 215 2368 216
rect 2362 211 2363 215
rect 2367 211 2368 215
rect 2362 210 2368 211
rect 2682 215 2688 216
rect 2682 211 2683 215
rect 2687 211 2688 215
rect 2682 210 2688 211
rect 2850 215 2856 216
rect 2850 211 2851 215
rect 2855 211 2856 215
rect 2850 210 2856 211
rect 2150 199 2156 200
rect 2150 195 2151 199
rect 2155 195 2156 199
rect 2150 194 2156 195
rect 2302 199 2308 200
rect 2302 195 2303 199
rect 2307 195 2308 199
rect 2302 194 2308 195
rect 2078 155 2084 156
rect 2152 155 2154 194
rect 2304 155 2306 194
rect 2364 188 2366 210
rect 2462 199 2468 200
rect 2462 195 2463 199
rect 2467 195 2468 199
rect 2462 194 2468 195
rect 2622 199 2628 200
rect 2622 195 2623 199
rect 2627 195 2628 199
rect 2622 194 2628 195
rect 2362 187 2368 188
rect 2362 183 2363 187
rect 2367 183 2368 187
rect 2362 182 2368 183
rect 2464 155 2466 194
rect 2506 187 2512 188
rect 2506 183 2507 187
rect 2511 183 2512 187
rect 2506 182 2512 183
rect 1407 154 1411 155
rect 1407 149 1411 150
rect 1439 154 1443 155
rect 1439 149 1443 150
rect 1503 154 1507 155
rect 1503 149 1507 150
rect 1823 154 1827 155
rect 1823 149 1827 150
rect 1863 154 1867 155
rect 1863 149 1867 150
rect 1895 154 1899 155
rect 1895 149 1899 150
rect 1983 154 1987 155
rect 1983 149 1987 150
rect 2007 154 2011 155
rect 2007 149 2011 150
rect 2071 154 2075 155
rect 2078 151 2079 155
rect 2083 151 2084 155
rect 2078 150 2084 151
rect 2151 154 2155 155
rect 2071 149 2075 150
rect 2151 149 2155 150
rect 2159 154 2163 155
rect 2159 149 2163 150
rect 2247 154 2251 155
rect 2247 149 2251 150
rect 2303 154 2307 155
rect 2303 149 2307 150
rect 2335 154 2339 155
rect 2335 149 2339 150
rect 2439 154 2443 155
rect 2439 149 2443 150
rect 2463 154 2467 155
rect 2463 149 2467 150
rect 1362 147 1368 148
rect 1362 143 1363 147
rect 1367 143 1368 147
rect 1362 142 1368 143
rect 1408 138 1410 149
rect 1504 138 1506 149
rect 1230 137 1236 138
rect 1230 133 1231 137
rect 1235 133 1236 137
rect 1230 132 1236 133
rect 1318 137 1324 138
rect 1318 133 1319 137
rect 1323 133 1324 137
rect 1318 132 1324 133
rect 1406 137 1412 138
rect 1406 133 1407 137
rect 1411 133 1412 137
rect 1406 132 1412 133
rect 1502 137 1508 138
rect 1502 133 1503 137
rect 1507 133 1508 137
rect 1502 132 1508 133
rect 1824 125 1826 149
rect 1864 125 1866 149
rect 1896 138 1898 149
rect 1984 138 1986 149
rect 2072 138 2074 149
rect 2160 138 2162 149
rect 2248 138 2250 149
rect 2336 138 2338 149
rect 2440 138 2442 149
rect 2498 147 2504 148
rect 2498 143 2499 147
rect 2503 143 2504 147
rect 2498 142 2504 143
rect 1894 137 1900 138
rect 1894 133 1895 137
rect 1899 133 1900 137
rect 1894 132 1900 133
rect 1982 137 1988 138
rect 1982 133 1983 137
rect 1987 133 1988 137
rect 1982 132 1988 133
rect 2070 137 2076 138
rect 2070 133 2071 137
rect 2075 133 2076 137
rect 2070 132 2076 133
rect 2158 137 2164 138
rect 2158 133 2159 137
rect 2163 133 2164 137
rect 2158 132 2164 133
rect 2246 137 2252 138
rect 2246 133 2247 137
rect 2251 133 2252 137
rect 2246 132 2252 133
rect 2334 137 2340 138
rect 2334 133 2335 137
rect 2339 133 2340 137
rect 2334 132 2340 133
rect 2438 137 2444 138
rect 2438 133 2439 137
rect 2443 133 2444 137
rect 2438 132 2444 133
rect 1822 124 1828 125
rect 1822 120 1823 124
rect 1827 120 1828 124
rect 110 119 116 120
rect 782 119 788 120
rect 782 115 783 119
rect 787 115 788 119
rect 782 114 788 115
rect 946 119 952 120
rect 946 115 947 119
rect 951 115 952 119
rect 946 114 952 115
rect 1122 119 1128 120
rect 1122 115 1123 119
rect 1127 115 1128 119
rect 1122 114 1128 115
rect 1210 119 1216 120
rect 1822 119 1828 120
rect 1862 124 1868 125
rect 2500 124 2502 142
rect 1862 120 1863 124
rect 1867 120 1868 124
rect 1862 119 1868 120
rect 2498 123 2504 124
rect 2498 119 2499 123
rect 2503 119 2504 123
rect 2508 120 2510 182
rect 2624 155 2626 194
rect 2684 188 2686 210
rect 2790 199 2796 200
rect 2790 195 2791 199
rect 2795 195 2796 199
rect 2790 194 2796 195
rect 2682 187 2688 188
rect 2682 183 2683 187
rect 2687 183 2688 187
rect 2682 182 2688 183
rect 2792 155 2794 194
rect 2852 188 2854 210
rect 2958 199 2964 200
rect 2958 195 2959 199
rect 2963 195 2964 199
rect 2958 194 2964 195
rect 2850 187 2856 188
rect 2850 183 2851 187
rect 2855 183 2856 187
rect 2850 182 2856 183
rect 2960 155 2962 194
rect 2988 188 2990 266
rect 3086 261 3092 262
rect 3086 257 3087 261
rect 3091 257 3092 261
rect 3086 256 3092 257
rect 3088 251 3090 256
rect 3087 250 3091 251
rect 3087 245 3091 246
rect 3127 250 3131 251
rect 3127 245 3131 246
rect 3128 240 3130 245
rect 3126 239 3132 240
rect 3126 235 3127 239
rect 3131 235 3132 239
rect 3126 234 3132 235
rect 3240 232 3242 306
rect 3296 302 3298 313
rect 3488 302 3490 313
rect 3520 312 3522 394
rect 3575 389 3579 390
rect 3576 374 3578 389
rect 3574 373 3580 374
rect 3574 369 3575 373
rect 3579 369 3580 373
rect 3574 368 3580 369
rect 3574 356 3580 357
rect 3574 352 3575 356
rect 3579 352 3580 356
rect 3574 351 3580 352
rect 3576 319 3578 351
rect 3575 318 3579 319
rect 3575 313 3579 314
rect 3518 311 3524 312
rect 3518 307 3519 311
rect 3523 307 3524 311
rect 3518 306 3524 307
rect 3294 301 3300 302
rect 3294 297 3295 301
rect 3299 297 3300 301
rect 3294 296 3300 297
rect 3486 301 3492 302
rect 3486 297 3487 301
rect 3491 297 3492 301
rect 3486 296 3492 297
rect 3576 289 3578 313
rect 3574 288 3580 289
rect 3574 284 3575 288
rect 3579 284 3580 288
rect 3574 283 3580 284
rect 3574 271 3580 272
rect 3574 267 3575 271
rect 3579 267 3580 271
rect 3574 266 3580 267
rect 3286 261 3292 262
rect 3286 257 3287 261
rect 3291 257 3292 261
rect 3286 256 3292 257
rect 3478 261 3484 262
rect 3478 257 3479 261
rect 3483 257 3484 261
rect 3478 256 3484 257
rect 3288 251 3290 256
rect 3480 251 3482 256
rect 3518 255 3524 256
rect 3518 251 3519 255
rect 3523 251 3524 255
rect 3576 251 3578 266
rect 3287 250 3291 251
rect 3287 245 3291 246
rect 3311 250 3315 251
rect 3311 245 3315 246
rect 3479 250 3483 251
rect 3518 250 3524 251
rect 3575 250 3579 251
rect 3479 245 3483 246
rect 3312 240 3314 245
rect 3480 240 3482 245
rect 3310 239 3316 240
rect 3310 235 3311 239
rect 3315 235 3316 239
rect 3310 234 3316 235
rect 3478 239 3484 240
rect 3478 235 3479 239
rect 3483 235 3484 239
rect 3478 234 3484 235
rect 3238 231 3244 232
rect 3238 227 3239 231
rect 3243 227 3244 231
rect 3238 226 3244 227
rect 3194 215 3200 216
rect 3194 211 3195 215
rect 3199 211 3200 215
rect 3194 210 3200 211
rect 3134 199 3140 200
rect 3134 195 3135 199
rect 3139 195 3140 199
rect 3134 194 3140 195
rect 2986 187 2992 188
rect 2986 183 2987 187
rect 2991 183 2992 187
rect 2986 182 2992 183
rect 3136 155 3138 194
rect 3196 188 3198 210
rect 3318 199 3324 200
rect 3318 195 3319 199
rect 3323 195 3324 199
rect 3318 194 3324 195
rect 3486 199 3492 200
rect 3486 195 3487 199
rect 3491 195 3492 199
rect 3486 194 3492 195
rect 3194 187 3200 188
rect 3194 183 3195 187
rect 3199 183 3200 187
rect 3194 182 3200 183
rect 3320 155 3322 194
rect 3370 187 3376 188
rect 3370 183 3371 187
rect 3375 183 3376 187
rect 3370 182 3376 183
rect 2543 154 2547 155
rect 2543 149 2547 150
rect 2623 154 2627 155
rect 2623 149 2627 150
rect 2647 154 2651 155
rect 2647 149 2651 150
rect 2743 154 2747 155
rect 2743 149 2747 150
rect 2791 154 2795 155
rect 2791 149 2795 150
rect 2839 154 2843 155
rect 2839 149 2843 150
rect 2935 154 2939 155
rect 2935 149 2939 150
rect 2959 154 2963 155
rect 2959 149 2963 150
rect 3031 154 3035 155
rect 3031 149 3035 150
rect 3127 154 3131 155
rect 3127 149 3131 150
rect 3135 154 3139 155
rect 3135 149 3139 150
rect 3223 154 3227 155
rect 3223 149 3227 150
rect 3311 154 3315 155
rect 3311 149 3315 150
rect 3319 154 3323 155
rect 3319 149 3323 150
rect 2544 138 2546 149
rect 2648 138 2650 149
rect 2744 138 2746 149
rect 2840 138 2842 149
rect 2936 138 2938 149
rect 3032 138 3034 149
rect 3128 138 3130 149
rect 3224 138 3226 149
rect 3312 138 3314 149
rect 2542 137 2548 138
rect 2542 133 2543 137
rect 2547 133 2548 137
rect 2542 132 2548 133
rect 2646 137 2652 138
rect 2646 133 2647 137
rect 2651 133 2652 137
rect 2646 132 2652 133
rect 2742 137 2748 138
rect 2742 133 2743 137
rect 2747 133 2748 137
rect 2742 132 2748 133
rect 2838 137 2844 138
rect 2838 133 2839 137
rect 2843 133 2844 137
rect 2838 132 2844 133
rect 2934 137 2940 138
rect 2934 133 2935 137
rect 2939 133 2940 137
rect 2934 132 2940 133
rect 3030 137 3036 138
rect 3030 133 3031 137
rect 3035 133 3036 137
rect 3030 132 3036 133
rect 3126 137 3132 138
rect 3126 133 3127 137
rect 3131 133 3132 137
rect 3126 132 3132 133
rect 3222 137 3228 138
rect 3222 133 3223 137
rect 3227 133 3228 137
rect 3222 132 3228 133
rect 3310 137 3316 138
rect 3310 133 3311 137
rect 3315 133 3316 137
rect 3310 132 3316 133
rect 3372 124 3374 182
rect 3488 155 3490 194
rect 3520 188 3522 250
rect 3575 245 3579 246
rect 3576 230 3578 245
rect 3574 229 3580 230
rect 3574 225 3575 229
rect 3579 225 3580 229
rect 3574 224 3580 225
rect 3546 215 3552 216
rect 3546 211 3547 215
rect 3551 211 3552 215
rect 3546 210 3552 211
rect 3574 212 3580 213
rect 3518 187 3524 188
rect 3518 183 3519 187
rect 3523 183 3524 187
rect 3518 182 3524 183
rect 3399 154 3403 155
rect 3399 149 3403 150
rect 3487 154 3491 155
rect 3487 149 3491 150
rect 3400 138 3402 149
rect 3466 147 3472 148
rect 3466 143 3467 147
rect 3471 143 3472 147
rect 3466 142 3472 143
rect 3398 137 3404 138
rect 3398 133 3399 137
rect 3403 133 3404 137
rect 3398 132 3404 133
rect 3370 123 3376 124
rect 1210 115 1211 119
rect 1215 115 1216 119
rect 2498 118 2504 119
rect 2506 119 2512 120
rect 1210 114 1216 115
rect 2506 115 2507 119
rect 2511 115 2512 119
rect 3370 119 3371 123
rect 3375 119 3376 123
rect 3468 120 3470 142
rect 3488 138 3490 149
rect 3548 148 3550 210
rect 3574 208 3575 212
rect 3579 208 3580 212
rect 3574 207 3580 208
rect 3576 155 3578 207
rect 3575 154 3579 155
rect 3575 149 3579 150
rect 3546 147 3552 148
rect 3546 143 3547 147
rect 3551 143 3552 147
rect 3546 142 3552 143
rect 3486 137 3492 138
rect 3486 133 3487 137
rect 3491 133 3492 137
rect 3486 132 3492 133
rect 3576 125 3578 149
rect 3574 124 3580 125
rect 3574 120 3575 124
rect 3579 120 3580 124
rect 3370 118 3376 119
rect 3466 119 3472 120
rect 3574 119 3580 120
rect 2506 114 2512 115
rect 3466 115 3467 119
rect 3471 115 3472 119
rect 3466 114 3472 115
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 110 102 116 103
rect 1822 107 1828 108
rect 1822 103 1823 107
rect 1827 103 1828 107
rect 1822 102 1828 103
rect 1862 107 1868 108
rect 1862 103 1863 107
rect 1867 103 1868 107
rect 1862 102 1868 103
rect 3574 107 3580 108
rect 3574 103 3575 107
rect 3579 103 3580 107
rect 3574 102 3580 103
rect 112 87 114 102
rect 166 97 172 98
rect 166 93 167 97
rect 171 93 172 97
rect 166 92 172 93
rect 254 97 260 98
rect 254 93 255 97
rect 259 93 260 97
rect 254 92 260 93
rect 342 97 348 98
rect 342 93 343 97
rect 347 93 348 97
rect 342 92 348 93
rect 430 97 436 98
rect 430 93 431 97
rect 435 93 436 97
rect 430 92 436 93
rect 518 97 524 98
rect 518 93 519 97
rect 523 93 524 97
rect 518 92 524 93
rect 606 97 612 98
rect 606 93 607 97
rect 611 93 612 97
rect 606 92 612 93
rect 694 97 700 98
rect 694 93 695 97
rect 699 93 700 97
rect 694 92 700 93
rect 782 97 788 98
rect 782 93 783 97
rect 787 93 788 97
rect 782 92 788 93
rect 870 97 876 98
rect 870 93 871 97
rect 875 93 876 97
rect 870 92 876 93
rect 958 97 964 98
rect 958 93 959 97
rect 963 93 964 97
rect 958 92 964 93
rect 1046 97 1052 98
rect 1046 93 1047 97
rect 1051 93 1052 97
rect 1046 92 1052 93
rect 1134 97 1140 98
rect 1134 93 1135 97
rect 1139 93 1140 97
rect 1134 92 1140 93
rect 1222 97 1228 98
rect 1222 93 1223 97
rect 1227 93 1228 97
rect 1222 92 1228 93
rect 1310 97 1316 98
rect 1310 93 1311 97
rect 1315 93 1316 97
rect 1310 92 1316 93
rect 1398 97 1404 98
rect 1398 93 1399 97
rect 1403 93 1404 97
rect 1398 92 1404 93
rect 1494 97 1500 98
rect 1494 93 1495 97
rect 1499 93 1500 97
rect 1494 92 1500 93
rect 168 87 170 92
rect 256 87 258 92
rect 344 87 346 92
rect 432 87 434 92
rect 520 87 522 92
rect 608 87 610 92
rect 696 87 698 92
rect 784 87 786 92
rect 872 87 874 92
rect 960 87 962 92
rect 1048 87 1050 92
rect 1136 87 1138 92
rect 1224 87 1226 92
rect 1312 87 1314 92
rect 1400 87 1402 92
rect 1496 87 1498 92
rect 1824 87 1826 102
rect 1864 87 1866 102
rect 1886 97 1892 98
rect 1886 93 1887 97
rect 1891 93 1892 97
rect 1886 92 1892 93
rect 1974 97 1980 98
rect 1974 93 1975 97
rect 1979 93 1980 97
rect 1974 92 1980 93
rect 2062 97 2068 98
rect 2062 93 2063 97
rect 2067 93 2068 97
rect 2062 92 2068 93
rect 2150 97 2156 98
rect 2150 93 2151 97
rect 2155 93 2156 97
rect 2150 92 2156 93
rect 2238 97 2244 98
rect 2238 93 2239 97
rect 2243 93 2244 97
rect 2238 92 2244 93
rect 2326 97 2332 98
rect 2326 93 2327 97
rect 2331 93 2332 97
rect 2326 92 2332 93
rect 2430 97 2436 98
rect 2430 93 2431 97
rect 2435 93 2436 97
rect 2430 92 2436 93
rect 2534 97 2540 98
rect 2534 93 2535 97
rect 2539 93 2540 97
rect 2534 92 2540 93
rect 2638 97 2644 98
rect 2638 93 2639 97
rect 2643 93 2644 97
rect 2638 92 2644 93
rect 2734 97 2740 98
rect 2734 93 2735 97
rect 2739 93 2740 97
rect 2734 92 2740 93
rect 2830 97 2836 98
rect 2830 93 2831 97
rect 2835 93 2836 97
rect 2830 92 2836 93
rect 2926 97 2932 98
rect 2926 93 2927 97
rect 2931 93 2932 97
rect 2926 92 2932 93
rect 3022 97 3028 98
rect 3022 93 3023 97
rect 3027 93 3028 97
rect 3022 92 3028 93
rect 3118 97 3124 98
rect 3118 93 3119 97
rect 3123 93 3124 97
rect 3118 92 3124 93
rect 3214 97 3220 98
rect 3214 93 3215 97
rect 3219 93 3220 97
rect 3214 92 3220 93
rect 3302 97 3308 98
rect 3302 93 3303 97
rect 3307 93 3308 97
rect 3302 92 3308 93
rect 3390 97 3396 98
rect 3390 93 3391 97
rect 3395 93 3396 97
rect 3390 92 3396 93
rect 3478 97 3484 98
rect 3478 93 3479 97
rect 3483 93 3484 97
rect 3478 92 3484 93
rect 1888 87 1890 92
rect 1976 87 1978 92
rect 2064 87 2066 92
rect 2152 87 2154 92
rect 2240 87 2242 92
rect 2328 87 2330 92
rect 2432 87 2434 92
rect 2536 87 2538 92
rect 2640 87 2642 92
rect 2736 87 2738 92
rect 2832 87 2834 92
rect 2928 87 2930 92
rect 3024 87 3026 92
rect 3120 87 3122 92
rect 3216 87 3218 92
rect 3304 87 3306 92
rect 3392 87 3394 92
rect 3480 87 3482 92
rect 3576 87 3578 102
rect 111 86 115 87
rect 111 81 115 82
rect 167 86 171 87
rect 167 81 171 82
rect 255 86 259 87
rect 255 81 259 82
rect 343 86 347 87
rect 343 81 347 82
rect 431 86 435 87
rect 431 81 435 82
rect 519 86 523 87
rect 519 81 523 82
rect 607 86 611 87
rect 607 81 611 82
rect 695 86 699 87
rect 695 81 699 82
rect 783 86 787 87
rect 783 81 787 82
rect 871 86 875 87
rect 871 81 875 82
rect 959 86 963 87
rect 959 81 963 82
rect 1047 86 1051 87
rect 1047 81 1051 82
rect 1135 86 1139 87
rect 1135 81 1139 82
rect 1223 86 1227 87
rect 1223 81 1227 82
rect 1311 86 1315 87
rect 1311 81 1315 82
rect 1399 86 1403 87
rect 1399 81 1403 82
rect 1495 86 1499 87
rect 1495 81 1499 82
rect 1823 86 1827 87
rect 1823 81 1827 82
rect 1863 86 1867 87
rect 1863 81 1867 82
rect 1887 86 1891 87
rect 1887 81 1891 82
rect 1975 86 1979 87
rect 1975 81 1979 82
rect 2063 86 2067 87
rect 2063 81 2067 82
rect 2151 86 2155 87
rect 2151 81 2155 82
rect 2239 86 2243 87
rect 2239 81 2243 82
rect 2327 86 2331 87
rect 2327 81 2331 82
rect 2431 86 2435 87
rect 2431 81 2435 82
rect 2535 86 2539 87
rect 2535 81 2539 82
rect 2639 86 2643 87
rect 2639 81 2643 82
rect 2735 86 2739 87
rect 2735 81 2739 82
rect 2831 86 2835 87
rect 2831 81 2835 82
rect 2927 86 2931 87
rect 2927 81 2931 82
rect 3023 86 3027 87
rect 3023 81 3027 82
rect 3119 86 3123 87
rect 3119 81 3123 82
rect 3215 86 3219 87
rect 3215 81 3219 82
rect 3303 86 3307 87
rect 3303 81 3307 82
rect 3391 86 3395 87
rect 3391 81 3395 82
rect 3479 86 3483 87
rect 3479 81 3483 82
rect 3575 86 3579 87
rect 3575 81 3579 82
<< m4c >>
rect 111 3646 115 3650
rect 239 3646 243 3650
rect 327 3646 331 3650
rect 415 3646 419 3650
rect 503 3646 507 3650
rect 591 3646 595 3650
rect 679 3646 683 3650
rect 1823 3646 1827 3650
rect 111 3570 115 3574
rect 231 3570 235 3574
rect 247 3570 251 3574
rect 1863 3582 1867 3586
rect 1887 3582 1891 3586
rect 1975 3582 1979 3586
rect 2063 3582 2067 3586
rect 2151 3582 2155 3586
rect 2239 3582 2243 3586
rect 2327 3582 2331 3586
rect 2415 3582 2419 3586
rect 2503 3582 2507 3586
rect 2591 3582 2595 3586
rect 2679 3582 2683 3586
rect 2767 3582 2771 3586
rect 2855 3582 2859 3586
rect 2943 3582 2947 3586
rect 3031 3582 3035 3586
rect 3119 3582 3123 3586
rect 3207 3582 3211 3586
rect 3295 3582 3299 3586
rect 3575 3582 3579 3586
rect 319 3570 323 3574
rect 399 3570 403 3574
rect 407 3570 411 3574
rect 495 3570 499 3574
rect 543 3570 547 3574
rect 583 3570 587 3574
rect 671 3570 675 3574
rect 687 3570 691 3574
rect 823 3570 827 3574
rect 951 3570 955 3574
rect 1079 3570 1083 3574
rect 1199 3570 1203 3574
rect 1311 3570 1315 3574
rect 1423 3570 1427 3574
rect 1543 3570 1547 3574
rect 1823 3570 1827 3574
rect 111 3502 115 3506
rect 183 3502 187 3506
rect 255 3502 259 3506
rect 351 3502 355 3506
rect 407 3502 411 3506
rect 519 3502 523 3506
rect 551 3502 555 3506
rect 679 3502 683 3506
rect 695 3502 699 3506
rect 1247 3512 1251 3516
rect 831 3502 835 3506
rect 959 3502 963 3506
rect 967 3502 971 3506
rect 1087 3502 1091 3506
rect 1095 3502 1099 3506
rect 1207 3502 1211 3506
rect 1215 3502 1219 3506
rect 111 3434 115 3438
rect 135 3434 139 3438
rect 175 3434 179 3438
rect 255 3434 259 3438
rect 343 3434 347 3438
rect 415 3434 419 3438
rect 511 3434 515 3438
rect 583 3434 587 3438
rect 671 3434 675 3438
rect 759 3434 763 3438
rect 823 3434 827 3438
rect 935 3434 939 3438
rect 959 3434 963 3438
rect 1491 3512 1495 3516
rect 1319 3502 1323 3506
rect 1335 3502 1339 3506
rect 1431 3502 1435 3506
rect 1455 3502 1459 3506
rect 1551 3502 1555 3506
rect 1575 3502 1579 3506
rect 1823 3502 1827 3506
rect 1863 3506 1867 3510
rect 1895 3506 1899 3510
rect 1911 3506 1915 3510
rect 1983 3506 1987 3510
rect 2015 3506 2019 3510
rect 2071 3506 2075 3510
rect 2135 3506 2139 3510
rect 2159 3506 2163 3510
rect 2247 3506 2251 3510
rect 2263 3506 2267 3510
rect 2335 3506 2339 3510
rect 2391 3506 2395 3510
rect 2423 3506 2427 3510
rect 2511 3506 2515 3510
rect 2527 3506 2531 3510
rect 1087 3434 1091 3438
rect 1111 3434 1115 3438
rect 1207 3434 1211 3438
rect 1295 3434 1299 3438
rect 1327 3434 1331 3438
rect 111 3358 115 3362
rect 143 3358 147 3362
rect 207 3358 211 3362
rect 263 3358 267 3362
rect 367 3358 371 3362
rect 423 3358 427 3362
rect 535 3358 539 3362
rect 591 3358 595 3362
rect 695 3358 699 3362
rect 767 3358 771 3362
rect 855 3358 859 3362
rect 943 3358 947 3362
rect 999 3358 1003 3362
rect 1119 3358 1123 3362
rect 111 3286 115 3290
rect 199 3286 203 3290
rect 255 3286 259 3290
rect 359 3286 363 3290
rect 375 3286 379 3290
rect 511 3286 515 3290
rect 527 3286 531 3290
rect 663 3286 667 3290
rect 687 3286 691 3290
rect 823 3286 827 3290
rect 847 3286 851 3290
rect 1447 3434 1451 3438
rect 1479 3434 1483 3438
rect 1567 3434 1571 3438
rect 1823 3434 1827 3438
rect 1863 3430 1867 3434
rect 1903 3430 1907 3434
rect 1911 3430 1915 3434
rect 2007 3430 2011 3434
rect 2071 3430 2075 3434
rect 2127 3430 2131 3434
rect 2599 3506 2603 3510
rect 2663 3506 2667 3510
rect 2687 3506 2691 3510
rect 2775 3506 2779 3510
rect 2799 3506 2803 3510
rect 2863 3506 2867 3510
rect 2943 3506 2947 3510
rect 2951 3506 2955 3510
rect 3039 3506 3043 3510
rect 3087 3506 3091 3510
rect 3127 3506 3131 3510
rect 3215 3506 3219 3510
rect 2223 3430 2227 3434
rect 2255 3430 2259 3434
rect 2367 3430 2371 3434
rect 2383 3430 2387 3434
rect 1143 3358 1147 3362
rect 1279 3358 1283 3362
rect 1303 3358 1307 3362
rect 1415 3358 1419 3362
rect 1487 3358 1491 3362
rect 1559 3358 1563 3362
rect 1823 3358 1827 3362
rect 1863 3358 1867 3362
rect 1895 3358 1899 3362
rect 1919 3358 1923 3362
rect 2047 3358 2051 3362
rect 2079 3358 2083 3362
rect 2207 3358 2211 3362
rect 991 3286 995 3290
rect 1135 3286 1139 3290
rect 1167 3286 1171 3290
rect 1271 3286 1275 3290
rect 1343 3286 1347 3290
rect 295 3264 299 3268
rect 619 3264 623 3268
rect 463 3232 467 3236
rect 111 3214 115 3218
rect 263 3214 267 3218
rect 383 3214 387 3218
rect 431 3214 435 3218
rect 739 3232 743 3236
rect 519 3214 523 3218
rect 551 3214 555 3218
rect 671 3214 675 3218
rect 799 3214 803 3218
rect 831 3214 835 3218
rect 935 3214 939 3218
rect 999 3214 1003 3218
rect 1079 3214 1083 3218
rect 1175 3214 1179 3218
rect 111 3142 115 3146
rect 423 3142 427 3146
rect 463 3142 467 3146
rect 543 3142 547 3146
rect 551 3142 555 3146
rect 639 3142 643 3146
rect 663 3142 667 3146
rect 735 3142 739 3146
rect 791 3142 795 3146
rect 847 3142 851 3146
rect 927 3142 931 3146
rect 967 3142 971 3146
rect 1407 3286 1411 3290
rect 1519 3286 1523 3290
rect 1551 3286 1555 3290
rect 1823 3286 1827 3290
rect 1863 3286 1867 3290
rect 1887 3286 1891 3290
rect 2039 3286 2043 3290
rect 2063 3286 2067 3290
rect 2503 3430 2507 3434
rect 2519 3430 2523 3434
rect 2631 3430 2635 3434
rect 2655 3430 2659 3434
rect 3303 3506 3307 3510
rect 3575 3506 3579 3510
rect 2759 3430 2763 3434
rect 2791 3430 2795 3434
rect 2231 3358 2235 3362
rect 2367 3358 2371 3362
rect 2375 3358 2379 3362
rect 2511 3358 2515 3362
rect 2535 3358 2539 3362
rect 2887 3430 2891 3434
rect 2935 3430 2939 3434
rect 3023 3430 3027 3434
rect 3079 3430 3083 3434
rect 3575 3430 3579 3434
rect 2639 3358 2643 3362
rect 2703 3358 2707 3362
rect 2767 3358 2771 3362
rect 2879 3358 2883 3362
rect 2895 3358 2899 3362
rect 3031 3358 3035 3362
rect 3055 3358 3059 3362
rect 2199 3286 2203 3290
rect 2263 3286 2267 3290
rect 2359 3286 2363 3290
rect 2455 3286 2459 3290
rect 1231 3214 1235 3218
rect 1351 3214 1355 3218
rect 1383 3214 1387 3218
rect 1527 3214 1531 3218
rect 1535 3214 1539 3218
rect 1823 3214 1827 3218
rect 1863 3218 1867 3222
rect 1895 3218 1899 3222
rect 2071 3218 2075 3222
rect 2087 3218 2091 3222
rect 2271 3218 2275 3222
rect 2303 3218 2307 3222
rect 1071 3142 1075 3146
rect 1095 3142 1099 3146
rect 1223 3142 1227 3146
rect 1231 3142 1235 3146
rect 1375 3142 1379 3146
rect 111 3066 115 3070
rect 151 3066 155 3070
rect 239 3066 243 3070
rect 327 3066 331 3070
rect 415 3066 419 3070
rect 471 3066 475 3070
rect 503 3066 507 3070
rect 559 3066 563 3070
rect 591 3066 595 3070
rect 647 3066 651 3070
rect 679 3066 683 3070
rect 743 3066 747 3070
rect 767 3066 771 3070
rect 855 3066 859 3070
rect 223 3059 227 3060
rect 223 3056 227 3059
rect 1519 3142 1523 3146
rect 1527 3142 1531 3146
rect 1823 3142 1827 3146
rect 1863 3146 1867 3150
rect 1887 3146 1891 3150
rect 2079 3146 2083 3150
rect 2527 3286 2531 3290
rect 2639 3286 2643 3290
rect 2695 3286 2699 3290
rect 3575 3358 3579 3362
rect 2815 3286 2819 3290
rect 2871 3286 2875 3290
rect 2983 3286 2987 3290
rect 3047 3286 3051 3290
rect 3151 3286 3155 3290
rect 3319 3286 3323 3290
rect 3479 3286 3483 3290
rect 3575 3286 3579 3290
rect 2463 3218 2467 3222
rect 2511 3218 2515 3222
rect 2647 3218 2651 3222
rect 2703 3218 2707 3222
rect 2823 3218 2827 3222
rect 2879 3218 2883 3222
rect 2991 3218 2995 3222
rect 3039 3218 3043 3222
rect 2295 3146 2299 3150
rect 2503 3146 2507 3150
rect 943 3066 947 3070
rect 975 3066 979 3070
rect 1031 3066 1035 3070
rect 1103 3066 1107 3070
rect 1119 3066 1123 3070
rect 1207 3066 1211 3070
rect 1239 3066 1243 3070
rect 1295 3066 1299 3070
rect 1383 3066 1387 3070
rect 1471 3066 1475 3070
rect 1527 3066 1531 3070
rect 1559 3066 1563 3070
rect 915 3056 919 3060
rect 1647 3066 1651 3070
rect 1735 3066 1739 3070
rect 1823 3066 1827 3070
rect 1863 3066 1867 3070
rect 1895 3066 1899 3070
rect 2087 3066 2091 3070
rect 2255 3066 2259 3070
rect 111 2990 115 2994
rect 143 2990 147 2994
rect 231 2990 235 2994
rect 319 2990 323 2994
rect 407 2990 411 2994
rect 495 2990 499 2994
rect 583 2990 587 2994
rect 671 2990 675 2994
rect 759 2990 763 2994
rect 847 2990 851 2994
rect 935 2990 939 2994
rect 1023 2990 1027 2994
rect 1111 2990 1115 2994
rect 1199 2990 1203 2994
rect 1287 2990 1291 2994
rect 1375 2990 1379 2994
rect 1407 2990 1411 2994
rect 1463 2990 1467 2994
rect 1519 2990 1523 2994
rect 111 2922 115 2926
rect 1359 2922 1363 2926
rect 1415 2922 1419 2926
rect 1471 2922 1475 2926
rect 1551 2990 1555 2994
rect 1631 2990 1635 2994
rect 1639 2990 1643 2994
rect 2695 3146 2699 3150
rect 3159 3218 3163 3222
rect 3199 3218 3203 3222
rect 3327 3218 3331 3222
rect 3351 3218 3355 3222
rect 3487 3218 3491 3222
rect 2871 3146 2875 3150
rect 3031 3146 3035 3150
rect 3039 3146 3043 3150
rect 3191 3146 3195 3150
rect 3343 3146 3347 3150
rect 3575 3218 3579 3222
rect 3479 3146 3483 3150
rect 3575 3146 3579 3150
rect 2303 3066 2307 3070
rect 2423 3066 2427 3070
rect 2511 3066 2515 3070
rect 2591 3066 2595 3070
rect 2703 3066 2707 3070
rect 2751 3066 2755 3070
rect 2879 3066 2883 3070
rect 2919 3066 2923 3070
rect 3047 3066 3051 3070
rect 3087 3066 3091 3070
rect 3199 3066 3203 3070
rect 3351 3066 3355 3070
rect 3487 3066 3491 3070
rect 2783 3059 2787 3060
rect 2783 3056 2787 3059
rect 1727 2990 1731 2994
rect 1823 2990 1827 2994
rect 1863 2994 1867 2998
rect 2239 2994 2243 2998
rect 2247 2994 2251 2998
rect 2415 2994 2419 2998
rect 2463 2994 2467 2998
rect 1527 2922 1531 2926
rect 1583 2922 1587 2926
rect 1639 2922 1643 2926
rect 1703 2922 1707 2926
rect 1735 2922 1739 2926
rect 111 2850 115 2854
rect 135 2850 139 2854
rect 223 2850 227 2854
rect 311 2850 315 2854
rect 399 2850 403 2854
rect 487 2850 491 2854
rect 599 2850 603 2854
rect 727 2850 731 2854
rect 863 2850 867 2854
rect 999 2850 1003 2854
rect 1135 2850 1139 2854
rect 1263 2850 1267 2854
rect 1351 2850 1355 2854
rect 1383 2850 1387 2854
rect 111 2782 115 2786
rect 143 2782 147 2786
rect 191 2782 195 2786
rect 231 2782 235 2786
rect 295 2782 299 2786
rect 319 2782 323 2786
rect 407 2782 411 2786
rect 415 2782 419 2786
rect 495 2782 499 2786
rect 551 2782 555 2786
rect 607 2782 611 2786
rect 687 2782 691 2786
rect 735 2782 739 2786
rect 823 2782 827 2786
rect 871 2782 875 2786
rect 959 2782 963 2786
rect 1007 2782 1011 2786
rect 111 2706 115 2710
rect 167 2706 171 2710
rect 183 2706 187 2710
rect 279 2706 283 2710
rect 287 2706 291 2710
rect 391 2706 395 2710
rect 407 2706 411 2710
rect 111 2622 115 2626
rect 175 2622 179 2626
rect 223 2622 227 2626
rect 503 2706 507 2710
rect 543 2706 547 2710
rect 1463 2850 1467 2854
rect 1503 2850 1507 2854
rect 1575 2850 1579 2854
rect 1623 2850 1627 2854
rect 1695 2850 1699 2854
rect 1823 2922 1827 2926
rect 1863 2910 1867 2914
rect 2239 2910 2243 2914
rect 2247 2910 2251 2914
rect 2583 2994 2587 2998
rect 2671 2994 2675 2998
rect 2743 2994 2747 2998
rect 2863 2994 2867 2998
rect 2911 2994 2915 2998
rect 3035 3056 3039 3060
rect 3031 2994 3035 2998
rect 3079 2994 3083 2998
rect 3191 2994 3195 2998
rect 3343 2994 3347 2998
rect 3479 2994 3483 2998
rect 2711 2936 2715 2940
rect 2959 2936 2963 2940
rect 2463 2910 2467 2914
rect 2471 2910 2475 2914
rect 2671 2910 2675 2914
rect 2679 2910 2683 2914
rect 2855 2910 2859 2914
rect 2871 2910 2875 2914
rect 3023 2910 3027 2914
rect 3039 2910 3043 2914
rect 3183 2910 3187 2914
rect 3199 2910 3203 2914
rect 3335 2910 3339 2914
rect 3351 2910 3355 2914
rect 3487 2910 3491 2914
rect 3575 3066 3579 3070
rect 3575 2994 3579 2998
rect 3575 2910 3579 2914
rect 2751 2864 2755 2868
rect 3099 2864 3103 2868
rect 1727 2850 1731 2854
rect 1823 2850 1827 2854
rect 1863 2838 1867 2842
rect 1895 2838 1899 2842
rect 1983 2838 1987 2842
rect 2071 2838 2075 2842
rect 2159 2838 2163 2842
rect 2231 2838 2235 2842
rect 2247 2838 2251 2842
rect 2335 2838 2339 2842
rect 2423 2838 2427 2842
rect 2455 2838 2459 2842
rect 2511 2838 2515 2842
rect 1087 2782 1091 2786
rect 1143 2782 1147 2786
rect 1207 2782 1211 2786
rect 1271 2782 1275 2786
rect 1319 2782 1323 2786
rect 1391 2782 1395 2786
rect 1431 2782 1435 2786
rect 1511 2782 1515 2786
rect 1535 2782 1539 2786
rect 1631 2782 1635 2786
rect 1647 2782 1651 2786
rect 1735 2782 1739 2786
rect 1823 2782 1827 2786
rect 1863 2758 1867 2762
rect 1903 2758 1907 2762
rect 1991 2758 1995 2762
rect 2047 2758 2051 2762
rect 2079 2758 2083 2762
rect 2167 2758 2171 2762
rect 2255 2758 2259 2762
rect 2295 2758 2299 2762
rect 2343 2758 2347 2762
rect 2431 2758 2435 2762
rect 2447 2758 2451 2762
rect 615 2706 619 2710
rect 679 2706 683 2710
rect 815 2706 819 2710
rect 951 2706 955 2710
rect 1079 2706 1083 2710
rect 1199 2706 1203 2710
rect 1311 2706 1315 2710
rect 1423 2706 1427 2710
rect 1527 2706 1531 2710
rect 1639 2706 1643 2710
rect 1727 2706 1731 2710
rect 1823 2706 1827 2710
rect 1863 2690 1867 2694
rect 1943 2690 1947 2694
rect 2599 2838 2603 2842
rect 2663 2838 2667 2842
rect 2687 2838 2691 2842
rect 2791 2838 2795 2842
rect 2847 2838 2851 2842
rect 2903 2838 2907 2842
rect 3015 2838 3019 2842
rect 3031 2838 3035 2842
rect 3175 2838 3179 2842
rect 3327 2838 3331 2842
rect 3479 2838 3483 2842
rect 2519 2758 2523 2762
rect 2607 2758 2611 2762
rect 2623 2758 2627 2762
rect 2695 2758 2699 2762
rect 2799 2758 2803 2762
rect 2823 2758 2827 2762
rect 2911 2758 2915 2762
rect 3039 2758 3043 2762
rect 3575 2838 3579 2842
rect 3183 2758 3187 2762
rect 3271 2758 3275 2762
rect 3335 2758 3339 2762
rect 3487 2758 3491 2762
rect 2039 2690 2043 2694
rect 2055 2690 2059 2694
rect 2159 2690 2163 2694
rect 2167 2690 2171 2694
rect 2287 2690 2291 2694
rect 287 2622 291 2626
rect 351 2622 355 2626
rect 399 2622 403 2626
rect 495 2622 499 2626
rect 511 2622 515 2626
rect 623 2622 627 2626
rect 663 2622 667 2626
rect 839 2622 843 2626
rect 1023 2622 1027 2626
rect 1215 2622 1219 2626
rect 1407 2622 1411 2626
rect 1607 2622 1611 2626
rect 1823 2622 1827 2626
rect 111 2554 115 2558
rect 215 2554 219 2558
rect 271 2554 275 2558
rect 343 2554 347 2558
rect 471 2554 475 2558
rect 487 2554 491 2558
rect 111 2482 115 2486
rect 183 2482 187 2486
rect 655 2554 659 2558
rect 671 2554 675 2558
rect 831 2554 835 2558
rect 855 2554 859 2558
rect 1015 2554 1019 2558
rect 1023 2554 1027 2558
rect 1175 2554 1179 2558
rect 1207 2554 1211 2558
rect 1863 2618 1867 2622
rect 1895 2618 1899 2622
rect 1951 2618 1955 2622
rect 2063 2618 2067 2622
rect 2071 2618 2075 2622
rect 2175 2618 2179 2622
rect 1319 2554 1323 2558
rect 1399 2554 1403 2558
rect 1455 2554 1459 2558
rect 1591 2554 1595 2558
rect 1599 2554 1603 2558
rect 1727 2554 1731 2558
rect 279 2482 283 2486
rect 319 2482 323 2486
rect 463 2482 467 2486
rect 479 2482 483 2486
rect 607 2482 611 2486
rect 679 2482 683 2486
rect 743 2482 747 2486
rect 863 2482 867 2486
rect 879 2482 883 2486
rect 1007 2482 1011 2486
rect 1031 2482 1035 2486
rect 1823 2554 1827 2558
rect 1863 2550 1867 2554
rect 1887 2550 1891 2554
rect 2407 2690 2411 2694
rect 2439 2690 2443 2694
rect 2519 2690 2523 2694
rect 2263 2618 2267 2622
rect 2295 2618 2299 2622
rect 2415 2618 2419 2622
rect 2463 2618 2467 2622
rect 2615 2690 2619 2694
rect 2631 2690 2635 2694
rect 2735 2690 2739 2694
rect 2815 2690 2819 2694
rect 2847 2690 2851 2694
rect 2959 2690 2963 2694
rect 3031 2690 3035 2694
rect 3071 2690 3075 2694
rect 3575 2758 3579 2762
rect 3263 2690 3267 2694
rect 3479 2690 3483 2694
rect 2527 2618 2531 2622
rect 2639 2618 2643 2622
rect 2663 2618 2667 2622
rect 2743 2618 2747 2622
rect 2855 2618 2859 2622
rect 2871 2618 2875 2622
rect 2967 2618 2971 2622
rect 3079 2618 3083 2622
rect 3295 2618 3299 2622
rect 3487 2618 3491 2622
rect 3575 2690 3579 2694
rect 3575 2618 3579 2622
rect 2039 2550 2043 2554
rect 2063 2550 2067 2554
rect 2215 2550 2219 2554
rect 2255 2550 2259 2554
rect 2399 2550 2403 2554
rect 2455 2550 2459 2554
rect 2575 2550 2579 2554
rect 2655 2550 2659 2554
rect 2743 2550 2747 2554
rect 1127 2482 1131 2486
rect 1183 2482 1187 2486
rect 1239 2482 1243 2486
rect 1327 2482 1331 2486
rect 1343 2482 1347 2486
rect 1447 2482 1451 2486
rect 1463 2482 1467 2486
rect 1551 2482 1555 2486
rect 1599 2482 1603 2486
rect 1647 2482 1651 2486
rect 1735 2482 1739 2486
rect 1823 2482 1827 2486
rect 1863 2482 1867 2486
rect 1895 2482 1899 2486
rect 1991 2482 1995 2486
rect 2047 2482 2051 2486
rect 2127 2482 2131 2486
rect 2223 2482 2227 2486
rect 111 2406 115 2410
rect 151 2406 155 2410
rect 175 2406 179 2410
rect 311 2406 315 2410
rect 319 2406 323 2410
rect 111 2334 115 2338
rect 143 2334 147 2338
rect 159 2334 163 2338
rect 455 2406 459 2410
rect 479 2406 483 2410
rect 599 2406 603 2410
rect 639 2406 643 2410
rect 735 2406 739 2410
rect 783 2406 787 2410
rect 871 2406 875 2410
rect 919 2406 923 2410
rect 999 2406 1003 2410
rect 1047 2406 1051 2410
rect 1119 2406 1123 2410
rect 2279 2482 2283 2486
rect 2407 2482 2411 2486
rect 2439 2482 2443 2486
rect 2583 2482 2587 2486
rect 2599 2482 2603 2486
rect 2863 2550 2867 2554
rect 2903 2550 2907 2554
rect 3055 2550 3059 2554
rect 3071 2550 3075 2554
rect 3199 2550 3203 2554
rect 3287 2550 3291 2554
rect 3343 2550 3347 2554
rect 3479 2550 3483 2554
rect 2751 2482 2755 2486
rect 2767 2482 2771 2486
rect 2911 2482 2915 2486
rect 2943 2482 2947 2486
rect 3063 2482 3067 2486
rect 3119 2482 3123 2486
rect 3575 2550 3579 2554
rect 3207 2482 3211 2486
rect 3295 2482 3299 2486
rect 3351 2482 3355 2486
rect 3471 2482 3475 2486
rect 3487 2482 3491 2486
rect 1175 2406 1179 2410
rect 1231 2406 1235 2410
rect 1303 2406 1307 2410
rect 1335 2406 1339 2410
rect 1431 2406 1435 2410
rect 1439 2406 1443 2410
rect 1543 2406 1547 2410
rect 1639 2406 1643 2410
rect 1727 2406 1731 2410
rect 1823 2406 1827 2410
rect 1863 2406 1867 2410
rect 1887 2406 1891 2410
rect 1983 2406 1987 2410
rect 2119 2406 2123 2410
rect 2271 2406 2275 2410
rect 2351 2406 2355 2410
rect 263 2334 267 2338
rect 327 2334 331 2338
rect 407 2334 411 2338
rect 487 2334 491 2338
rect 543 2334 547 2338
rect 647 2334 651 2338
rect 679 2334 683 2338
rect 791 2334 795 2338
rect 807 2334 811 2338
rect 927 2334 931 2338
rect 111 2266 115 2270
rect 135 2266 139 2270
rect 231 2266 235 2270
rect 255 2266 259 2270
rect 351 2266 355 2270
rect 399 2266 403 2270
rect 2431 2406 2435 2410
rect 2503 2406 2507 2410
rect 2591 2406 2595 2410
rect 2655 2406 2659 2410
rect 1039 2334 1043 2338
rect 1055 2334 1059 2338
rect 1159 2334 1163 2338
rect 1183 2334 1187 2338
rect 1279 2334 1283 2338
rect 1311 2334 1315 2338
rect 1439 2334 1443 2338
rect 1823 2334 1827 2338
rect 1863 2334 1867 2338
rect 2351 2334 2355 2338
rect 2359 2334 2363 2338
rect 2447 2334 2451 2338
rect 2511 2334 2515 2338
rect 2559 2334 2563 2338
rect 1027 2312 1031 2316
rect 1227 2312 1231 2316
rect 2759 2406 2763 2410
rect 2807 2406 2811 2410
rect 2935 2406 2939 2410
rect 2967 2406 2971 2410
rect 3111 2406 3115 2410
rect 3135 2406 3139 2410
rect 3287 2406 3291 2410
rect 3303 2406 3307 2410
rect 3575 2482 3579 2486
rect 3463 2406 3467 2410
rect 3471 2406 3475 2410
rect 2663 2334 2667 2338
rect 2703 2334 2707 2338
rect 2815 2334 2819 2338
rect 2879 2334 2883 2338
rect 2975 2334 2979 2338
rect 3079 2334 3083 2338
rect 3143 2334 3147 2338
rect 3287 2334 3291 2338
rect 3311 2334 3315 2338
rect 471 2266 475 2270
rect 535 2266 539 2270
rect 591 2266 595 2270
rect 671 2266 675 2270
rect 711 2266 715 2270
rect 799 2266 803 2270
rect 823 2266 827 2270
rect 919 2266 923 2270
rect 935 2266 939 2270
rect 1031 2266 1035 2270
rect 1055 2266 1059 2270
rect 1151 2266 1155 2270
rect 1175 2266 1179 2270
rect 1271 2266 1275 2270
rect 1823 2266 1827 2270
rect 1863 2266 1867 2270
rect 2335 2266 2339 2270
rect 2343 2266 2347 2270
rect 111 2194 115 2198
rect 143 2194 147 2198
rect 239 2194 243 2198
rect 247 2194 251 2198
rect 359 2194 363 2198
rect 383 2194 387 2198
rect 479 2194 483 2198
rect 519 2194 523 2198
rect 599 2194 603 2198
rect 111 2118 115 2122
rect 135 2118 139 2122
rect 231 2118 235 2122
rect 239 2118 243 2122
rect 359 2118 363 2122
rect 375 2118 379 2122
rect 655 2194 659 2198
rect 719 2194 723 2198
rect 783 2194 787 2198
rect 831 2194 835 2198
rect 911 2194 915 2198
rect 943 2194 947 2198
rect 2439 2266 2443 2270
rect 2447 2266 2451 2270
rect 2551 2266 2555 2270
rect 2583 2266 2587 2270
rect 2695 2266 2699 2270
rect 2735 2266 2739 2270
rect 2871 2266 2875 2270
rect 2911 2266 2915 2270
rect 1031 2194 1035 2198
rect 1063 2194 1067 2198
rect 1159 2194 1163 2198
rect 1183 2194 1187 2198
rect 1287 2194 1291 2198
rect 1823 2194 1827 2198
rect 1863 2198 1867 2202
rect 2255 2198 2259 2202
rect 2343 2198 2347 2202
rect 2439 2198 2443 2202
rect 2455 2198 2459 2202
rect 2551 2198 2555 2202
rect 2591 2198 2595 2202
rect 2695 2198 2699 2202
rect 3071 2266 3075 2270
rect 3103 2266 3107 2270
rect 3279 2266 3283 2270
rect 3303 2266 3307 2270
rect 3575 2406 3579 2410
rect 3479 2334 3483 2338
rect 3487 2334 3491 2338
rect 3575 2334 3579 2338
rect 3479 2266 3483 2270
rect 2743 2198 2747 2202
rect 2871 2198 2875 2202
rect 3575 2266 3579 2270
rect 2919 2198 2923 2202
rect 3071 2198 3075 2202
rect 3111 2198 3115 2202
rect 3287 2198 3291 2202
rect 3311 2198 3315 2202
rect 479 2118 483 2122
rect 511 2118 515 2122
rect 599 2118 603 2122
rect 647 2118 651 2122
rect 719 2118 723 2122
rect 775 2118 779 2122
rect 831 2118 835 2122
rect 903 2118 907 2122
rect 943 2118 947 2122
rect 1023 2118 1027 2122
rect 1055 2118 1059 2122
rect 1151 2118 1155 2122
rect 1175 2118 1179 2122
rect 1279 2118 1283 2122
rect 1823 2118 1827 2122
rect 1863 2122 1867 2126
rect 2151 2122 2155 2126
rect 2239 2122 2243 2126
rect 2247 2122 2251 2126
rect 2327 2122 2331 2126
rect 2335 2122 2339 2126
rect 111 2038 115 2042
rect 143 2038 147 2042
rect 167 2038 171 2042
rect 239 2038 243 2042
rect 311 2038 315 2042
rect 367 2038 371 2042
rect 447 2038 451 2042
rect 487 2038 491 2042
rect 575 2038 579 2042
rect 607 2038 611 2042
rect 111 1970 115 1974
rect 159 1970 163 1974
rect 295 1970 299 1974
rect 303 1970 307 1974
rect 695 2038 699 2042
rect 727 2038 731 2042
rect 439 1970 443 1974
rect 567 1970 571 1974
rect 583 1970 587 1974
rect 687 1970 691 1974
rect 719 1970 723 1974
rect 2191 2064 2195 2068
rect 1863 2050 1867 2054
rect 1999 2050 2003 2054
rect 2127 2050 2131 2054
rect 2159 2050 2163 2054
rect 2247 2050 2251 2054
rect 2255 2050 2259 2054
rect 807 2038 811 2042
rect 839 2038 843 2042
rect 911 2038 915 2042
rect 951 2038 955 2042
rect 1015 2038 1019 2042
rect 1063 2038 1067 2042
rect 1119 2038 1123 2042
rect 1183 2038 1187 2042
rect 1223 2038 1227 2042
rect 1327 2038 1331 2042
rect 1823 2038 1827 2042
rect 799 1970 803 1974
rect 855 1970 859 1974
rect 903 1970 907 1974
rect 991 1970 995 1974
rect 1007 1970 1011 1974
rect 111 1894 115 1898
rect 167 1894 171 1898
rect 223 1894 227 1898
rect 303 1894 307 1898
rect 447 1894 451 1898
rect 479 1894 483 1898
rect 591 1894 595 1898
rect 719 1894 723 1898
rect 727 1894 731 1898
rect 111 1826 115 1830
rect 215 1826 219 1830
rect 247 1826 251 1830
rect 415 1826 419 1830
rect 471 1826 475 1830
rect 591 1826 595 1830
rect 711 1826 715 1830
rect 1111 1970 1115 1974
rect 1119 1970 1123 1974
rect 1215 1970 1219 1974
rect 1239 1970 1243 1974
rect 2415 2122 2419 2126
rect 2431 2122 2435 2126
rect 2503 2122 2507 2126
rect 2543 2122 2547 2126
rect 2615 2122 2619 2126
rect 2687 2122 2691 2126
rect 2751 2122 2755 2126
rect 2863 2122 2867 2126
rect 2919 2122 2923 2126
rect 3063 2122 3067 2126
rect 3103 2122 3107 2126
rect 3279 2122 3283 2126
rect 3303 2122 3307 2126
rect 2663 2104 2667 2108
rect 3199 2104 3203 2108
rect 2483 2064 2487 2068
rect 2335 2050 2339 2054
rect 2399 2050 2403 2054
rect 2423 2050 2427 2054
rect 2511 2050 2515 2054
rect 2551 2050 2555 2054
rect 2623 2050 2627 2054
rect 2711 2050 2715 2054
rect 2759 2050 2763 2054
rect 2879 2050 2883 2054
rect 2927 2050 2931 2054
rect 3063 2050 3067 2054
rect 3111 2050 3115 2054
rect 3247 2050 3251 2054
rect 3311 2050 3315 2054
rect 2071 2016 2075 2020
rect 2479 2019 2483 2020
rect 2479 2016 2483 2019
rect 3487 2198 3491 2202
rect 3575 2198 3579 2202
rect 3479 2122 3483 2126
rect 3575 2122 3579 2126
rect 3439 2050 3443 2054
rect 3487 2050 3491 2054
rect 1319 1970 1323 1974
rect 1359 1970 1363 1974
rect 1479 1970 1483 1974
rect 1599 1970 1603 1974
rect 1823 1970 1827 1974
rect 1863 1974 1867 1978
rect 1903 1974 1907 1978
rect 1991 1974 1995 1978
rect 2119 1974 2123 1978
rect 2159 1974 2163 1978
rect 863 1894 867 1898
rect 935 1894 939 1898
rect 999 1894 1003 1898
rect 1127 1894 1131 1898
rect 1247 1894 1251 1898
rect 1295 1894 1299 1898
rect 1367 1894 1371 1898
rect 1455 1894 1459 1898
rect 1487 1894 1491 1898
rect 1607 1894 1611 1898
rect 759 1826 763 1830
rect 927 1826 931 1830
rect 1863 1906 1867 1910
rect 1895 1906 1899 1910
rect 1911 1906 1915 1910
rect 1735 1894 1739 1898
rect 1823 1894 1827 1898
rect 1983 1906 1987 1910
rect 2247 1974 2251 1978
rect 2391 1974 2395 1978
rect 2399 1974 2403 1978
rect 2543 1974 2547 1978
rect 2615 1974 2619 1978
rect 2703 1974 2707 1978
rect 2815 1974 2819 1978
rect 2871 1974 2875 1978
rect 2999 1974 3003 1978
rect 3055 1974 3059 1978
rect 3167 1974 3171 1978
rect 3239 1974 3243 1978
rect 3335 1974 3339 1978
rect 2655 1936 2659 1940
rect 3151 1936 3155 1940
rect 2951 1920 2955 1924
rect 2071 1906 2075 1910
rect 2167 1906 2171 1910
rect 2295 1906 2299 1910
rect 2407 1906 2411 1910
rect 2447 1906 2451 1910
rect 2607 1906 2611 1910
rect 2623 1906 2627 1910
rect 2767 1906 2771 1910
rect 2823 1906 2827 1910
rect 2919 1906 2923 1910
rect 1943 1880 1947 1884
rect 1863 1834 1867 1838
rect 1887 1834 1891 1838
rect 1975 1834 1979 1838
rect 1999 1834 2003 1838
rect 2063 1834 2067 1838
rect 1079 1826 1083 1830
rect 1119 1826 1123 1830
rect 1223 1826 1227 1830
rect 1287 1826 1291 1830
rect 1359 1826 1363 1830
rect 1447 1826 1451 1830
rect 1487 1826 1491 1830
rect 1599 1826 1603 1830
rect 1615 1826 1619 1830
rect 1727 1826 1731 1830
rect 111 1754 115 1758
rect 255 1754 259 1758
rect 327 1754 331 1758
rect 423 1754 427 1758
rect 471 1754 475 1758
rect 599 1754 603 1758
rect 615 1754 619 1758
rect 767 1754 771 1758
rect 919 1754 923 1758
rect 935 1754 939 1758
rect 111 1682 115 1686
rect 311 1682 315 1686
rect 319 1682 323 1686
rect 447 1682 451 1686
rect 463 1682 467 1686
rect 591 1682 595 1686
rect 607 1682 611 1686
rect 111 1606 115 1610
rect 223 1606 227 1610
rect 735 1682 739 1686
rect 759 1682 763 1686
rect 1071 1754 1075 1758
rect 1087 1754 1091 1758
rect 1223 1754 1227 1758
rect 1231 1754 1235 1758
rect 1367 1754 1371 1758
rect 1375 1754 1379 1758
rect 887 1682 891 1686
rect 911 1682 915 1686
rect 1039 1682 1043 1686
rect 1063 1682 1067 1686
rect 1495 1754 1499 1758
rect 1527 1754 1531 1758
rect 1823 1826 1827 1830
rect 3259 1920 3263 1924
rect 3007 1906 3011 1910
rect 3071 1906 3075 1910
rect 3175 1906 3179 1910
rect 3215 1906 3219 1910
rect 3343 1906 3347 1910
rect 3359 1906 3363 1910
rect 2403 1880 2407 1884
rect 3431 1974 3435 1978
rect 3479 1974 3483 1978
rect 3487 1906 3491 1910
rect 3575 2050 3579 2054
rect 3575 1974 3579 1978
rect 3575 1906 3579 1910
rect 2159 1834 2163 1838
rect 2223 1834 2227 1838
rect 2287 1834 2291 1838
rect 2439 1834 2443 1838
rect 2599 1834 2603 1838
rect 2639 1834 2643 1838
rect 2759 1834 2763 1838
rect 2831 1834 2835 1838
rect 2911 1834 2915 1838
rect 3015 1834 3019 1838
rect 3063 1834 3067 1838
rect 3199 1834 3203 1838
rect 3207 1834 3211 1838
rect 3351 1834 3355 1838
rect 3391 1834 3395 1838
rect 3479 1834 3483 1838
rect 3575 1834 3579 1838
rect 2263 1792 2267 1796
rect 2675 1792 2679 1796
rect 2479 1776 2483 1780
rect 2719 1776 2723 1780
rect 1863 1762 1867 1766
rect 1943 1762 1947 1766
rect 2007 1762 2011 1766
rect 2087 1762 2091 1766
rect 2231 1762 2235 1766
rect 2247 1762 2251 1766
rect 2415 1762 2419 1766
rect 2447 1762 2451 1766
rect 2599 1762 2603 1766
rect 2647 1762 2651 1766
rect 2791 1762 2795 1766
rect 1623 1754 1627 1758
rect 1687 1754 1691 1758
rect 1735 1754 1739 1758
rect 1823 1754 1827 1758
rect 2839 1762 2843 1766
rect 2991 1762 2995 1766
rect 3023 1762 3027 1766
rect 3199 1762 3203 1766
rect 3207 1762 3211 1766
rect 1191 1682 1195 1686
rect 1215 1682 1219 1686
rect 1343 1682 1347 1686
rect 1367 1682 1371 1686
rect 1495 1682 1499 1686
rect 1519 1682 1523 1686
rect 1647 1682 1651 1686
rect 1679 1682 1683 1686
rect 319 1606 323 1610
rect 351 1606 355 1610
rect 455 1606 459 1610
rect 487 1606 491 1610
rect 599 1606 603 1610
rect 623 1606 627 1610
rect 743 1606 747 1610
rect 111 1534 115 1538
rect 135 1534 139 1538
rect 215 1534 219 1538
rect 271 1534 275 1538
rect 343 1534 347 1538
rect 423 1534 427 1538
rect 111 1458 115 1462
rect 143 1458 147 1462
rect 479 1534 483 1538
rect 583 1534 587 1538
rect 615 1534 619 1538
rect 759 1606 763 1610
rect 895 1606 899 1610
rect 903 1606 907 1610
rect 1047 1606 1051 1610
rect 1055 1606 1059 1610
rect 1199 1606 1203 1610
rect 735 1534 739 1538
rect 751 1534 755 1538
rect 887 1534 891 1538
rect 895 1534 899 1538
rect 1863 1690 1867 1694
rect 1911 1690 1915 1694
rect 1935 1690 1939 1694
rect 2031 1690 2035 1694
rect 2079 1690 2083 1694
rect 2151 1690 2155 1694
rect 2239 1690 2243 1694
rect 2271 1690 2275 1694
rect 1823 1682 1827 1686
rect 1863 1614 1867 1618
rect 1895 1614 1899 1618
rect 1919 1614 1923 1618
rect 1215 1606 1219 1610
rect 1351 1606 1355 1610
rect 1375 1606 1379 1610
rect 1503 1606 1507 1610
rect 1543 1606 1547 1610
rect 1655 1606 1659 1610
rect 1823 1606 1827 1610
rect 2399 1690 2403 1694
rect 2407 1690 2411 1694
rect 2543 1690 2547 1694
rect 2591 1690 2595 1694
rect 2695 1690 2699 1694
rect 2783 1690 2787 1694
rect 2863 1690 2867 1694
rect 2983 1690 2987 1694
rect 3047 1690 3051 1694
rect 2015 1614 2019 1618
rect 2039 1614 2043 1618
rect 2151 1614 2155 1618
rect 2159 1614 2163 1618
rect 2279 1614 2283 1618
rect 2287 1614 2291 1618
rect 2407 1614 2411 1618
rect 2431 1614 2435 1618
rect 2551 1614 2555 1618
rect 2583 1614 2587 1618
rect 3191 1690 3195 1694
rect 3399 1762 3403 1766
rect 3415 1762 3419 1766
rect 3575 1762 3579 1766
rect 3239 1690 3243 1694
rect 3407 1690 3411 1694
rect 3431 1690 3435 1694
rect 2703 1614 2707 1618
rect 2743 1614 2747 1618
rect 2871 1614 2875 1618
rect 2911 1614 2915 1618
rect 3055 1614 3059 1618
rect 3095 1614 3099 1618
rect 3247 1614 3251 1618
rect 3575 1690 3579 1694
rect 3279 1614 3283 1618
rect 3439 1614 3443 1618
rect 3471 1614 3475 1618
rect 1039 1534 1043 1538
rect 1047 1534 1051 1538
rect 1191 1534 1195 1538
rect 1207 1534 1211 1538
rect 1343 1534 1347 1538
rect 1367 1534 1371 1538
rect 1495 1534 1499 1538
rect 1535 1534 1539 1538
rect 263 1458 267 1462
rect 279 1458 283 1462
rect 399 1458 403 1462
rect 431 1458 435 1462
rect 535 1458 539 1462
rect 591 1458 595 1462
rect 663 1458 667 1462
rect 743 1458 747 1462
rect 791 1458 795 1462
rect 895 1458 899 1462
rect 911 1458 915 1462
rect 1023 1458 1027 1462
rect 1047 1458 1051 1462
rect 111 1390 115 1394
rect 135 1390 139 1394
rect 255 1390 259 1394
rect 327 1390 331 1394
rect 391 1390 395 1394
rect 527 1390 531 1394
rect 111 1314 115 1318
rect 143 1314 147 1318
rect 551 1390 555 1394
rect 1143 1458 1147 1462
rect 1199 1458 1203 1462
rect 1263 1458 1267 1462
rect 1351 1458 1355 1462
rect 1383 1458 1387 1462
rect 1823 1534 1827 1538
rect 1863 1538 1867 1542
rect 1887 1538 1891 1542
rect 2007 1538 2011 1542
rect 2023 1538 2027 1542
rect 2143 1538 2147 1542
rect 2183 1538 2187 1542
rect 2279 1538 2283 1542
rect 2343 1538 2347 1542
rect 2423 1538 2427 1542
rect 2503 1538 2507 1542
rect 2575 1538 2579 1542
rect 2663 1538 2667 1542
rect 2735 1538 2739 1542
rect 2823 1538 2827 1542
rect 2903 1538 2907 1542
rect 2983 1538 2987 1542
rect 3087 1538 3091 1542
rect 3151 1538 3155 1542
rect 3271 1538 3275 1542
rect 2703 1528 2707 1532
rect 1503 1458 1507 1462
rect 1631 1458 1635 1462
rect 1735 1458 1739 1462
rect 1823 1458 1827 1462
rect 1863 1462 1867 1466
rect 1895 1462 1899 1466
rect 2031 1462 2035 1466
rect 2183 1462 2187 1466
rect 2191 1462 2195 1466
rect 2351 1462 2355 1466
rect 2359 1462 2363 1466
rect 2511 1462 2515 1466
rect 2527 1462 2531 1466
rect 3019 1528 3023 1532
rect 3575 1614 3579 1618
rect 3319 1538 3323 1542
rect 3463 1538 3467 1542
rect 3479 1538 3483 1542
rect 2719 1480 2723 1484
rect 2671 1462 2675 1466
rect 2687 1462 2691 1466
rect 3079 1480 3083 1484
rect 2831 1462 2835 1466
rect 2847 1462 2851 1466
rect 2991 1462 2995 1466
rect 3007 1462 3011 1466
rect 3159 1462 3163 1466
rect 3175 1462 3179 1466
rect 3327 1462 3331 1466
rect 3343 1462 3347 1466
rect 2223 1432 2227 1436
rect 2427 1432 2431 1436
rect 655 1390 659 1394
rect 783 1390 787 1394
rect 903 1390 907 1394
rect 1015 1390 1019 1394
rect 1023 1390 1027 1394
rect 1135 1390 1139 1394
rect 1255 1390 1259 1394
rect 1263 1390 1267 1394
rect 1375 1390 1379 1394
rect 1495 1390 1499 1394
rect 1503 1390 1507 1394
rect 1623 1390 1627 1394
rect 1727 1390 1731 1394
rect 1823 1390 1827 1394
rect 1863 1386 1867 1390
rect 2079 1386 2083 1390
rect 2175 1386 2179 1390
rect 2263 1386 2267 1390
rect 2351 1386 2355 1390
rect 2439 1386 2443 1390
rect 1303 1336 1307 1340
rect 1639 1336 1643 1340
rect 2119 1328 2123 1332
rect 327 1314 331 1318
rect 335 1314 339 1318
rect 527 1314 531 1318
rect 559 1314 563 1318
rect 719 1314 723 1318
rect 791 1314 795 1318
rect 903 1314 907 1318
rect 1031 1314 1035 1318
rect 1071 1314 1075 1318
rect 1231 1314 1235 1318
rect 1271 1314 1275 1318
rect 1383 1314 1387 1318
rect 1511 1314 1515 1318
rect 111 1242 115 1246
rect 135 1242 139 1246
rect 295 1242 299 1246
rect 319 1242 323 1246
rect 479 1242 483 1246
rect 519 1242 523 1246
rect 655 1242 659 1246
rect 711 1242 715 1246
rect 815 1242 819 1246
rect 895 1242 899 1246
rect 967 1242 971 1246
rect 1063 1242 1067 1246
rect 1111 1242 1115 1246
rect 1223 1242 1227 1246
rect 1247 1242 1251 1246
rect 1375 1242 1379 1246
rect 1383 1242 1387 1246
rect 1535 1314 1539 1318
rect 1687 1314 1691 1318
rect 1735 1314 1739 1318
rect 1823 1314 1827 1318
rect 1863 1318 1867 1322
rect 2087 1318 2091 1322
rect 2271 1318 2275 1322
rect 2311 1318 2315 1322
rect 2519 1386 2523 1390
rect 2615 1386 2619 1390
rect 2679 1386 2683 1390
rect 2783 1386 2787 1390
rect 2839 1386 2843 1390
rect 2935 1386 2939 1390
rect 2999 1386 3003 1390
rect 3079 1386 3083 1390
rect 3167 1386 3171 1390
rect 3223 1386 3227 1390
rect 3335 1386 3339 1390
rect 3575 1538 3579 1542
rect 3487 1462 3491 1466
rect 3575 1462 3579 1466
rect 3359 1386 3363 1390
rect 3479 1386 3483 1390
rect 2823 1336 2827 1340
rect 2539 1328 2543 1332
rect 3259 1336 3263 1340
rect 3575 1386 3579 1390
rect 2447 1318 2451 1322
rect 2519 1318 2523 1322
rect 2623 1318 2627 1322
rect 2711 1318 2715 1322
rect 2791 1318 2795 1322
rect 2887 1318 2891 1322
rect 2943 1318 2947 1322
rect 3047 1318 3051 1322
rect 3087 1318 3091 1322
rect 3199 1318 3203 1322
rect 3231 1318 3235 1322
rect 3351 1318 3355 1322
rect 3367 1318 3371 1322
rect 2295 1288 2299 1292
rect 2443 1288 2447 1292
rect 1527 1242 1531 1246
rect 1679 1242 1683 1246
rect 1823 1242 1827 1246
rect 1863 1246 1867 1250
rect 1903 1246 1907 1250
rect 1991 1246 1995 1250
rect 2079 1246 2083 1250
rect 2095 1246 2099 1250
rect 111 1170 115 1174
rect 143 1170 147 1174
rect 167 1170 171 1174
rect 303 1170 307 1174
rect 319 1170 323 1174
rect 471 1170 475 1174
rect 487 1170 491 1174
rect 615 1170 619 1174
rect 663 1170 667 1174
rect 759 1170 763 1174
rect 823 1170 827 1174
rect 911 1170 915 1174
rect 975 1170 979 1174
rect 111 1098 115 1102
rect 159 1098 163 1102
rect 215 1098 219 1102
rect 311 1098 315 1102
rect 327 1098 331 1102
rect 439 1098 443 1102
rect 463 1098 467 1102
rect 559 1098 563 1102
rect 607 1098 611 1102
rect 1063 1170 1067 1174
rect 1119 1170 1123 1174
rect 1231 1170 1235 1174
rect 1255 1170 1259 1174
rect 1391 1170 1395 1174
rect 1399 1170 1403 1174
rect 1535 1170 1539 1174
rect 1575 1170 1579 1174
rect 1735 1170 1739 1174
rect 1823 1170 1827 1174
rect 1863 1174 1867 1178
rect 1895 1174 1899 1178
rect 1911 1174 1915 1178
rect 679 1098 683 1102
rect 751 1098 755 1102
rect 807 1098 811 1102
rect 903 1098 907 1102
rect 943 1098 947 1102
rect 1051 1160 1055 1164
rect 1539 1160 1543 1164
rect 1999 1174 2003 1178
rect 2063 1174 2067 1178
rect 2215 1246 2219 1250
rect 2303 1246 2307 1250
rect 2351 1246 2355 1250
rect 2487 1246 2491 1250
rect 2511 1246 2515 1250
rect 2631 1246 2635 1250
rect 2703 1246 2707 1250
rect 2775 1246 2779 1250
rect 2879 1246 2883 1250
rect 2919 1246 2923 1250
rect 2103 1174 2107 1178
rect 2223 1174 2227 1178
rect 2255 1174 2259 1178
rect 2359 1174 2363 1178
rect 2439 1174 2443 1178
rect 2495 1174 2499 1178
rect 2615 1174 2619 1178
rect 2639 1174 2643 1178
rect 1055 1098 1059 1102
rect 1087 1098 1091 1102
rect 1223 1098 1227 1102
rect 1247 1098 1251 1102
rect 1391 1098 1395 1102
rect 1407 1098 1411 1102
rect 1567 1098 1571 1102
rect 1575 1098 1579 1102
rect 1727 1098 1731 1102
rect 999 1080 1003 1084
rect 1339 1083 1343 1084
rect 1339 1080 1343 1083
rect 111 1022 115 1026
rect 223 1022 227 1026
rect 335 1022 339 1026
rect 343 1022 347 1026
rect 431 1022 435 1026
rect 447 1022 451 1026
rect 535 1022 539 1026
rect 567 1022 571 1026
rect 655 1022 659 1026
rect 687 1022 691 1026
rect 791 1022 795 1026
rect 815 1022 819 1026
rect 111 950 115 954
rect 335 950 339 954
rect 367 950 371 954
rect 423 950 427 954
rect 463 950 467 954
rect 527 950 531 954
rect 575 950 579 954
rect 647 950 651 954
rect 703 950 707 954
rect 783 950 787 954
rect 951 1022 955 1026
rect 1095 1022 1099 1026
rect 1135 1022 1139 1026
rect 1255 1022 1259 1026
rect 1327 1022 1331 1026
rect 1415 1022 1419 1026
rect 1535 1022 1539 1026
rect 847 950 851 954
rect 943 950 947 954
rect 1007 950 1011 954
rect 1127 950 1131 954
rect 1175 950 1179 954
rect 1823 1098 1827 1102
rect 1863 1094 1867 1098
rect 1887 1094 1891 1098
rect 1935 1094 1939 1098
rect 2055 1094 2059 1098
rect 2095 1094 2099 1098
rect 1583 1022 1587 1026
rect 1735 1022 1739 1026
rect 1823 1022 1827 1026
rect 1863 1022 1867 1026
rect 1943 1022 1947 1026
rect 2247 1094 2251 1098
rect 2407 1094 2411 1098
rect 2431 1094 2435 1098
rect 2815 1192 2819 1196
rect 3039 1246 3043 1250
rect 3063 1246 3067 1250
rect 3191 1246 3195 1250
rect 3207 1246 3211 1250
rect 3343 1246 3347 1250
rect 3351 1246 3355 1250
rect 3487 1318 3491 1322
rect 3575 1318 3579 1322
rect 3479 1246 3483 1250
rect 3139 1192 3143 1196
rect 2783 1174 2787 1178
rect 2791 1174 2795 1178
rect 2927 1174 2931 1178
rect 2967 1174 2971 1178
rect 3071 1174 3075 1178
rect 3143 1174 3147 1178
rect 3215 1174 3219 1178
rect 3327 1174 3331 1178
rect 3359 1174 3363 1178
rect 2567 1094 2571 1098
rect 2607 1094 2611 1098
rect 2735 1094 2739 1098
rect 2783 1094 2787 1098
rect 2911 1094 2915 1098
rect 2959 1094 2963 1098
rect 3095 1094 3099 1098
rect 3135 1094 3139 1098
rect 2071 1022 2075 1026
rect 2103 1022 2107 1026
rect 2191 1022 2195 1026
rect 2255 1022 2259 1026
rect 2311 1022 2315 1026
rect 1319 950 1323 954
rect 1351 950 1355 954
rect 1527 950 1531 954
rect 1711 950 1715 954
rect 1727 950 1731 954
rect 111 878 115 882
rect 343 878 347 882
rect 375 878 379 882
rect 431 878 435 882
rect 471 878 475 882
rect 535 878 539 882
rect 583 878 587 882
rect 1391 896 1395 900
rect 647 878 651 882
rect 711 878 715 882
rect 783 878 787 882
rect 855 878 859 882
rect 927 878 931 882
rect 1015 878 1019 882
rect 1087 878 1091 882
rect 1183 878 1187 882
rect 1263 878 1267 882
rect 1359 878 1363 882
rect 1447 878 1451 882
rect 1535 878 1539 882
rect 1631 878 1635 882
rect 111 810 115 814
rect 287 810 291 814
rect 335 810 339 814
rect 407 810 411 814
rect 423 810 427 814
rect 111 738 115 742
rect 215 738 219 742
rect 527 810 531 814
rect 535 810 539 814
rect 639 810 643 814
rect 679 810 683 814
rect 775 810 779 814
rect 823 810 827 814
rect 919 810 923 814
rect 975 810 979 814
rect 1079 810 1083 814
rect 1127 810 1131 814
rect 1667 896 1671 900
rect 1823 950 1827 954
rect 1863 950 1867 954
rect 1887 950 1891 954
rect 1935 950 1939 954
rect 2047 950 2051 954
rect 2063 950 2067 954
rect 2415 1022 2419 1026
rect 2439 1022 2443 1026
rect 2575 1022 2579 1026
rect 3287 1094 3291 1098
rect 3319 1094 3323 1098
rect 3575 1246 3579 1250
rect 3487 1174 3491 1178
rect 3575 1174 3579 1178
rect 3479 1094 3483 1098
rect 3575 1094 3579 1098
rect 2719 1022 2723 1026
rect 2743 1022 2747 1026
rect 2871 1022 2875 1026
rect 2919 1022 2923 1026
rect 3031 1022 3035 1026
rect 3103 1022 3107 1026
rect 3191 1022 3195 1026
rect 3295 1022 3299 1026
rect 3351 1022 3355 1026
rect 3487 1022 3491 1026
rect 3575 1022 3579 1026
rect 2183 950 2187 954
rect 2199 950 2203 954
rect 2303 950 2307 954
rect 2351 950 2355 954
rect 2431 950 2435 954
rect 2495 950 2499 954
rect 2567 950 2571 954
rect 1719 878 1723 882
rect 1823 878 1827 882
rect 1863 882 1867 886
rect 1895 882 1899 886
rect 2015 882 2019 886
rect 2631 950 2635 954
rect 2711 950 2715 954
rect 2759 950 2763 954
rect 2863 950 2867 954
rect 2887 950 2891 954
rect 3023 950 3027 954
rect 3183 950 3187 954
rect 3343 950 3347 954
rect 3479 950 3483 954
rect 3575 950 3579 954
rect 2055 882 2059 886
rect 2167 882 2171 886
rect 2207 882 2211 886
rect 2319 882 2323 886
rect 2359 882 2363 886
rect 1255 810 1259 814
rect 1279 810 1283 814
rect 1439 810 1443 814
rect 295 738 299 742
rect 359 738 363 742
rect 415 738 419 742
rect 503 738 507 742
rect 543 738 547 742
rect 647 738 651 742
rect 687 738 691 742
rect 1315 752 1319 756
rect 1599 810 1603 814
rect 1623 810 1627 814
rect 1823 810 1827 814
rect 1863 814 1867 818
rect 1887 814 1891 818
rect 1519 752 1523 756
rect 1991 814 1995 818
rect 2007 814 2011 818
rect 2135 814 2139 818
rect 2159 814 2163 818
rect 2487 882 2491 886
rect 2503 882 2507 886
rect 2639 882 2643 886
rect 2663 882 2667 886
rect 2767 882 2771 886
rect 2847 882 2851 886
rect 2895 882 2899 886
rect 3031 882 3035 886
rect 3039 882 3043 886
rect 2287 814 2291 818
rect 2311 814 2315 818
rect 2455 814 2459 818
rect 2479 814 2483 818
rect 2623 814 2627 818
rect 2655 814 2659 818
rect 791 738 795 742
rect 831 738 835 742
rect 935 738 939 742
rect 983 738 987 742
rect 1087 738 1091 742
rect 1135 738 1139 742
rect 1247 738 1251 742
rect 111 670 115 674
rect 135 670 139 674
rect 207 670 211 674
rect 295 670 299 674
rect 351 670 355 674
rect 463 670 467 674
rect 495 670 499 674
rect 623 670 627 674
rect 639 670 643 674
rect 775 670 779 674
rect 783 670 787 674
rect 927 670 931 674
rect 1071 670 1075 674
rect 1079 670 1083 674
rect 1287 738 1291 742
rect 1415 738 1419 742
rect 1447 738 1451 742
rect 1583 738 1587 742
rect 1607 738 1611 742
rect 1735 738 1739 742
rect 1823 738 1827 742
rect 1863 742 1867 746
rect 1895 742 1899 746
rect 1999 742 2003 746
rect 2063 742 2067 746
rect 2143 742 2147 746
rect 2255 742 2259 746
rect 2295 742 2299 746
rect 2447 742 2451 746
rect 2463 742 2467 746
rect 1207 670 1211 674
rect 1239 670 1243 674
rect 1343 670 1347 674
rect 1407 670 1411 674
rect 1479 670 1483 674
rect 111 598 115 602
rect 143 598 147 602
rect 303 598 307 602
rect 471 598 475 602
rect 487 598 491 602
rect 631 598 635 602
rect 671 598 675 602
rect 783 598 787 602
rect 847 598 851 602
rect 935 598 939 602
rect 1023 598 1027 602
rect 1079 598 1083 602
rect 1199 598 1203 602
rect 1215 598 1219 602
rect 1351 598 1355 602
rect 1375 598 1379 602
rect 111 526 115 530
rect 135 526 139 530
rect 295 526 299 530
rect 303 526 307 530
rect 479 526 483 530
rect 495 526 499 530
rect 663 526 667 530
rect 679 526 683 530
rect 839 526 843 530
rect 863 526 867 530
rect 1015 526 1019 530
rect 1031 526 1035 530
rect 1575 670 1579 674
rect 1615 670 1619 674
rect 1727 670 1731 674
rect 1487 598 1491 602
rect 1559 598 1563 602
rect 1823 670 1827 674
rect 1863 670 1867 674
rect 1887 670 1891 674
rect 2055 670 2059 674
rect 3239 882 3243 886
rect 3439 882 3443 886
rect 3575 882 3579 886
rect 2799 814 2803 818
rect 2839 814 2843 818
rect 2967 814 2971 818
rect 3031 814 3035 818
rect 3143 814 3147 818
rect 3231 814 3235 818
rect 3319 814 3323 818
rect 3431 814 3435 818
rect 3479 814 3483 818
rect 2631 742 2635 746
rect 2639 742 2643 746
rect 2807 742 2811 746
rect 2823 742 2827 746
rect 2975 742 2979 746
rect 2999 742 3003 746
rect 3151 742 3155 746
rect 3167 742 3171 746
rect 2215 670 2219 674
rect 2247 670 2251 674
rect 2359 670 2363 674
rect 2439 670 2443 674
rect 2511 670 2515 674
rect 2631 670 2635 674
rect 2671 670 2675 674
rect 2815 670 2819 674
rect 2831 670 2835 674
rect 2991 670 2995 674
rect 3575 814 3579 818
rect 3327 742 3331 746
rect 3335 742 3339 746
rect 3487 742 3491 746
rect 3575 742 3579 746
rect 3159 670 3163 674
rect 3327 670 3331 674
rect 3479 670 3483 674
rect 1623 598 1627 602
rect 1735 598 1739 602
rect 1823 598 1827 602
rect 1863 598 1867 602
rect 2199 598 2203 602
rect 2223 598 2227 602
rect 2287 598 2291 602
rect 2367 598 2371 602
rect 2375 598 2379 602
rect 2463 598 2467 602
rect 2519 598 2523 602
rect 2567 598 2571 602
rect 2679 598 2683 602
rect 2815 598 2819 602
rect 1191 526 1195 530
rect 111 454 115 458
rect 143 454 147 458
rect 303 454 307 458
rect 311 454 315 458
rect 495 454 499 458
rect 503 454 507 458
rect 687 454 691 458
rect 871 454 875 458
rect 879 454 883 458
rect 1039 454 1043 458
rect 1351 526 1355 530
rect 1367 526 1371 530
rect 1503 526 1507 530
rect 1551 526 1555 530
rect 1663 526 1667 530
rect 1055 454 1059 458
rect 1199 454 1203 458
rect 1223 454 1227 458
rect 1359 454 1363 458
rect 1391 454 1395 458
rect 111 386 115 390
rect 135 386 139 390
rect 263 386 267 390
rect 295 386 299 390
rect 423 386 427 390
rect 111 318 115 322
rect 143 318 147 322
rect 215 318 219 322
rect 487 386 491 390
rect 591 386 595 390
rect 679 386 683 390
rect 767 386 771 390
rect 871 386 875 390
rect 935 386 939 390
rect 1047 386 1051 390
rect 1511 454 1515 458
rect 1559 454 1563 458
rect 1727 526 1731 530
rect 1823 526 1827 530
rect 1863 526 1867 530
rect 2191 526 2195 530
rect 2839 598 2843 602
rect 2975 598 2979 602
rect 2999 598 3003 602
rect 3143 598 3147 602
rect 3167 598 3171 602
rect 3327 598 3331 602
rect 3335 598 3339 602
rect 2279 526 2283 530
rect 2303 526 2307 530
rect 2367 526 2371 530
rect 2399 526 2403 530
rect 2455 526 2459 530
rect 2503 526 2507 530
rect 2559 526 2563 530
rect 2607 526 2611 530
rect 2671 526 2675 530
rect 2719 526 2723 530
rect 2807 526 2811 530
rect 2839 526 2843 530
rect 2967 526 2971 530
rect 3095 526 3099 530
rect 3135 526 3139 530
rect 3575 670 3579 674
rect 3487 598 3491 602
rect 3575 598 3579 602
rect 3223 526 3227 530
rect 3319 526 3323 530
rect 3351 526 3355 530
rect 3479 526 3483 530
rect 1671 454 1675 458
rect 1727 454 1731 458
rect 1823 454 1827 458
rect 1863 458 1867 462
rect 2239 458 2243 462
rect 2311 458 2315 462
rect 2327 458 2331 462
rect 2407 458 2411 462
rect 2431 458 2435 462
rect 2511 458 2515 462
rect 2559 458 2563 462
rect 2615 458 2619 462
rect 1103 386 1107 390
rect 1215 386 1219 390
rect 1263 386 1267 390
rect 271 318 275 322
rect 351 318 355 322
rect 431 318 435 322
rect 495 318 499 322
rect 599 318 603 322
rect 639 318 643 322
rect 775 318 779 322
rect 111 242 115 246
rect 207 242 211 246
rect 231 242 235 246
rect 343 242 347 246
rect 359 242 363 246
rect 111 150 115 154
rect 175 150 179 154
rect 487 242 491 246
rect 791 318 795 322
rect 935 318 939 322
rect 943 318 947 322
rect 1079 318 1083 322
rect 1111 318 1115 322
rect 1223 318 1227 322
rect 623 242 627 246
rect 631 242 635 246
rect 759 242 763 246
rect 783 242 787 246
rect 895 242 899 246
rect 927 242 931 246
rect 1031 242 1035 246
rect 1071 242 1075 246
rect 1383 386 1387 390
rect 1423 386 1427 390
rect 1551 386 1555 390
rect 1583 386 1587 390
rect 1719 386 1723 390
rect 1727 386 1731 390
rect 1271 318 1275 322
rect 1359 318 1363 322
rect 1431 318 1435 322
rect 1487 318 1491 322
rect 1591 318 1595 322
rect 1623 318 1627 322
rect 1823 386 1827 390
rect 1863 390 1867 394
rect 2183 390 2187 394
rect 2231 390 2235 394
rect 2695 458 2699 462
rect 2727 458 2731 462
rect 2847 458 2851 462
rect 3007 472 3011 476
rect 3291 472 3295 476
rect 3575 526 3579 530
rect 2975 458 2979 462
rect 2999 458 3003 462
rect 3103 458 3107 462
rect 3159 458 3163 462
rect 3231 458 3235 462
rect 3327 458 3331 462
rect 3359 458 3363 462
rect 3487 458 3491 462
rect 3575 458 3579 462
rect 2287 390 2291 394
rect 2319 390 2323 394
rect 2399 390 2403 394
rect 2423 390 2427 394
rect 2527 390 2531 394
rect 2551 390 2555 394
rect 2671 390 2675 394
rect 2687 390 2691 394
rect 2815 390 2819 394
rect 2839 390 2843 394
rect 2967 390 2971 394
rect 2991 390 2995 394
rect 1735 318 1739 322
rect 1823 318 1827 322
rect 1863 314 1867 318
rect 1895 314 1899 318
rect 2087 314 2091 318
rect 2191 314 2195 318
rect 2295 314 2299 318
rect 2303 314 2307 318
rect 2407 314 2411 318
rect 2511 314 2515 318
rect 2535 314 2539 318
rect 1159 242 1163 246
rect 1215 242 1219 246
rect 1295 242 1299 246
rect 1351 242 1355 246
rect 1431 242 1435 246
rect 239 150 243 154
rect 263 150 267 154
rect 351 150 355 154
rect 367 150 371 154
rect 439 150 443 154
rect 495 150 499 154
rect 527 150 531 154
rect 615 150 619 154
rect 631 150 635 154
rect 703 150 707 154
rect 767 150 771 154
rect 791 150 795 154
rect 879 150 883 154
rect 903 150 907 154
rect 967 150 971 154
rect 1039 150 1043 154
rect 1055 150 1059 154
rect 1143 150 1147 154
rect 1167 150 1171 154
rect 1231 150 1235 154
rect 1303 150 1307 154
rect 1319 150 1323 154
rect 1479 242 1483 246
rect 1615 242 1619 246
rect 1727 242 1731 246
rect 1823 242 1827 246
rect 1863 246 1867 250
rect 1887 246 1891 250
rect 1999 246 2003 250
rect 2079 246 2083 250
rect 2143 246 2147 250
rect 2295 246 2299 250
rect 3127 390 3131 394
rect 3151 390 3155 394
rect 3295 390 3299 394
rect 3319 390 3323 394
rect 3463 390 3467 394
rect 3479 390 3483 394
rect 2679 314 2683 318
rect 2711 314 2715 318
rect 2823 314 2827 318
rect 2903 314 2907 318
rect 2975 314 2979 318
rect 3095 314 3099 318
rect 3135 314 3139 318
rect 3295 314 3299 318
rect 3303 314 3307 318
rect 3471 314 3475 318
rect 3487 314 3491 318
rect 2455 246 2459 250
rect 2503 246 2507 250
rect 2615 246 2619 250
rect 2703 246 2707 250
rect 2783 246 2787 250
rect 2895 246 2899 250
rect 2951 246 2955 250
rect 1407 150 1411 154
rect 1439 150 1443 154
rect 1503 150 1507 154
rect 1823 150 1827 154
rect 1863 150 1867 154
rect 1895 150 1899 154
rect 1983 150 1987 154
rect 2007 150 2011 154
rect 2071 150 2075 154
rect 2151 150 2155 154
rect 2159 150 2163 154
rect 2247 150 2251 154
rect 2303 150 2307 154
rect 2335 150 2339 154
rect 2439 150 2443 154
rect 2463 150 2467 154
rect 3087 246 3091 250
rect 3127 246 3131 250
rect 3575 390 3579 394
rect 3575 314 3579 318
rect 3287 246 3291 250
rect 3311 246 3315 250
rect 3479 246 3483 250
rect 2543 150 2547 154
rect 2623 150 2627 154
rect 2647 150 2651 154
rect 2743 150 2747 154
rect 2791 150 2795 154
rect 2839 150 2843 154
rect 2935 150 2939 154
rect 2959 150 2963 154
rect 3031 150 3035 154
rect 3127 150 3131 154
rect 3135 150 3139 154
rect 3223 150 3227 154
rect 3311 150 3315 154
rect 3319 150 3323 154
rect 3575 246 3579 250
rect 3399 150 3403 154
rect 3487 150 3491 154
rect 3575 150 3579 154
rect 111 82 115 86
rect 167 82 171 86
rect 255 82 259 86
rect 343 82 347 86
rect 431 82 435 86
rect 519 82 523 86
rect 607 82 611 86
rect 695 82 699 86
rect 783 82 787 86
rect 871 82 875 86
rect 959 82 963 86
rect 1047 82 1051 86
rect 1135 82 1139 86
rect 1223 82 1227 86
rect 1311 82 1315 86
rect 1399 82 1403 86
rect 1495 82 1499 86
rect 1823 82 1827 86
rect 1863 82 1867 86
rect 1887 82 1891 86
rect 1975 82 1979 86
rect 2063 82 2067 86
rect 2151 82 2155 86
rect 2239 82 2243 86
rect 2327 82 2331 86
rect 2431 82 2435 86
rect 2535 82 2539 86
rect 2639 82 2643 86
rect 2735 82 2739 86
rect 2831 82 2835 86
rect 2927 82 2931 86
rect 3023 82 3027 86
rect 3119 82 3123 86
rect 3215 82 3219 86
rect 3303 82 3307 86
rect 3391 82 3395 86
rect 3479 82 3483 86
rect 3575 82 3579 86
<< m4 >>
rect 96 3645 97 3651
rect 103 3650 1847 3651
rect 103 3646 111 3650
rect 115 3646 239 3650
rect 243 3646 327 3650
rect 331 3646 415 3650
rect 419 3646 503 3650
rect 507 3646 591 3650
rect 595 3646 679 3650
rect 683 3646 1823 3650
rect 1827 3646 1847 3650
rect 103 3645 1847 3646
rect 1853 3645 1854 3651
rect 1834 3581 1835 3587
rect 1841 3586 3599 3587
rect 1841 3582 1863 3586
rect 1867 3582 1887 3586
rect 1891 3582 1975 3586
rect 1979 3582 2063 3586
rect 2067 3582 2151 3586
rect 2155 3582 2239 3586
rect 2243 3582 2327 3586
rect 2331 3582 2415 3586
rect 2419 3582 2503 3586
rect 2507 3582 2591 3586
rect 2595 3582 2679 3586
rect 2683 3582 2767 3586
rect 2771 3582 2855 3586
rect 2859 3582 2943 3586
rect 2947 3582 3031 3586
rect 3035 3582 3119 3586
rect 3123 3582 3207 3586
rect 3211 3582 3295 3586
rect 3299 3582 3575 3586
rect 3579 3582 3599 3586
rect 1841 3581 3599 3582
rect 3605 3581 3606 3587
rect 84 3569 85 3575
rect 91 3574 1835 3575
rect 91 3570 111 3574
rect 115 3570 231 3574
rect 235 3570 247 3574
rect 251 3570 319 3574
rect 323 3570 399 3574
rect 403 3570 407 3574
rect 411 3570 495 3574
rect 499 3570 543 3574
rect 547 3570 583 3574
rect 587 3570 671 3574
rect 675 3570 687 3574
rect 691 3570 823 3574
rect 827 3570 951 3574
rect 955 3570 1079 3574
rect 1083 3570 1199 3574
rect 1203 3570 1311 3574
rect 1315 3570 1423 3574
rect 1427 3570 1543 3574
rect 1547 3570 1823 3574
rect 1827 3570 1835 3574
rect 91 3569 1835 3570
rect 1841 3569 1842 3575
rect 1246 3516 1252 3517
rect 1490 3516 1496 3517
rect 1246 3512 1247 3516
rect 1251 3512 1491 3516
rect 1495 3512 1496 3516
rect 1246 3511 1252 3512
rect 1490 3511 1496 3512
rect 1846 3510 3618 3511
rect 1846 3507 1863 3510
rect 96 3501 97 3507
rect 103 3506 1847 3507
rect 103 3502 111 3506
rect 115 3502 183 3506
rect 187 3502 255 3506
rect 259 3502 351 3506
rect 355 3502 407 3506
rect 411 3502 519 3506
rect 523 3502 551 3506
rect 555 3502 679 3506
rect 683 3502 695 3506
rect 699 3502 831 3506
rect 835 3502 959 3506
rect 963 3502 967 3506
rect 971 3502 1087 3506
rect 1091 3502 1095 3506
rect 1099 3502 1207 3506
rect 1211 3502 1215 3506
rect 1219 3502 1319 3506
rect 1323 3502 1335 3506
rect 1339 3502 1431 3506
rect 1435 3502 1455 3506
rect 1459 3502 1551 3506
rect 1555 3502 1575 3506
rect 1579 3502 1823 3506
rect 1827 3502 1847 3506
rect 103 3501 1847 3502
rect 1853 3506 1863 3507
rect 1867 3506 1895 3510
rect 1899 3506 1911 3510
rect 1915 3506 1983 3510
rect 1987 3506 2015 3510
rect 2019 3506 2071 3510
rect 2075 3506 2135 3510
rect 2139 3506 2159 3510
rect 2163 3506 2247 3510
rect 2251 3506 2263 3510
rect 2267 3506 2335 3510
rect 2339 3506 2391 3510
rect 2395 3506 2423 3510
rect 2427 3506 2511 3510
rect 2515 3506 2527 3510
rect 2531 3506 2599 3510
rect 2603 3506 2663 3510
rect 2667 3506 2687 3510
rect 2691 3506 2775 3510
rect 2779 3506 2799 3510
rect 2803 3506 2863 3510
rect 2867 3506 2943 3510
rect 2947 3506 2951 3510
rect 2955 3506 3039 3510
rect 3043 3506 3087 3510
rect 3091 3506 3127 3510
rect 3131 3506 3215 3510
rect 3219 3506 3303 3510
rect 3307 3506 3575 3510
rect 3579 3506 3618 3510
rect 1853 3505 3618 3506
rect 1853 3501 1854 3505
rect 84 3433 85 3439
rect 91 3438 1835 3439
rect 91 3434 111 3438
rect 115 3434 135 3438
rect 139 3434 175 3438
rect 179 3434 255 3438
rect 259 3434 343 3438
rect 347 3434 415 3438
rect 419 3434 511 3438
rect 515 3434 583 3438
rect 587 3434 671 3438
rect 675 3434 759 3438
rect 763 3434 823 3438
rect 827 3434 935 3438
rect 939 3434 959 3438
rect 963 3434 1087 3438
rect 1091 3434 1111 3438
rect 1115 3434 1207 3438
rect 1211 3434 1295 3438
rect 1299 3434 1327 3438
rect 1331 3434 1447 3438
rect 1451 3434 1479 3438
rect 1483 3434 1567 3438
rect 1571 3434 1823 3438
rect 1827 3434 1835 3438
rect 91 3433 1835 3434
rect 1841 3435 1842 3439
rect 1841 3434 3606 3435
rect 1841 3433 1863 3434
rect 1834 3430 1863 3433
rect 1867 3430 1903 3434
rect 1907 3430 1911 3434
rect 1915 3430 2007 3434
rect 2011 3430 2071 3434
rect 2075 3430 2127 3434
rect 2131 3430 2223 3434
rect 2227 3430 2255 3434
rect 2259 3430 2367 3434
rect 2371 3430 2383 3434
rect 2387 3430 2503 3434
rect 2507 3430 2519 3434
rect 2523 3430 2631 3434
rect 2635 3430 2655 3434
rect 2659 3430 2759 3434
rect 2763 3430 2791 3434
rect 2795 3430 2887 3434
rect 2891 3430 2935 3434
rect 2939 3430 3023 3434
rect 3027 3430 3079 3434
rect 3083 3430 3575 3434
rect 3579 3430 3606 3434
rect 1834 3429 3606 3430
rect 96 3357 97 3363
rect 103 3362 1847 3363
rect 103 3358 111 3362
rect 115 3358 143 3362
rect 147 3358 207 3362
rect 211 3358 263 3362
rect 267 3358 367 3362
rect 371 3358 423 3362
rect 427 3358 535 3362
rect 539 3358 591 3362
rect 595 3358 695 3362
rect 699 3358 767 3362
rect 771 3358 855 3362
rect 859 3358 943 3362
rect 947 3358 999 3362
rect 1003 3358 1119 3362
rect 1123 3358 1143 3362
rect 1147 3358 1279 3362
rect 1283 3358 1303 3362
rect 1307 3358 1415 3362
rect 1419 3358 1487 3362
rect 1491 3358 1559 3362
rect 1563 3358 1823 3362
rect 1827 3358 1847 3362
rect 103 3357 1847 3358
rect 1853 3362 3618 3363
rect 1853 3358 1863 3362
rect 1867 3358 1895 3362
rect 1899 3358 1919 3362
rect 1923 3358 2047 3362
rect 2051 3358 2079 3362
rect 2083 3358 2207 3362
rect 2211 3358 2231 3362
rect 2235 3358 2367 3362
rect 2371 3358 2375 3362
rect 2379 3358 2511 3362
rect 2515 3358 2535 3362
rect 2539 3358 2639 3362
rect 2643 3358 2703 3362
rect 2707 3358 2767 3362
rect 2771 3358 2879 3362
rect 2883 3358 2895 3362
rect 2899 3358 3031 3362
rect 3035 3358 3055 3362
rect 3059 3358 3575 3362
rect 3579 3358 3618 3362
rect 1853 3357 3618 3358
rect 84 3285 85 3291
rect 91 3290 1835 3291
rect 91 3286 111 3290
rect 115 3286 199 3290
rect 203 3286 255 3290
rect 259 3286 359 3290
rect 363 3286 375 3290
rect 379 3286 511 3290
rect 515 3286 527 3290
rect 531 3286 663 3290
rect 667 3286 687 3290
rect 691 3286 823 3290
rect 827 3286 847 3290
rect 851 3286 991 3290
rect 995 3286 1135 3290
rect 1139 3286 1167 3290
rect 1171 3286 1271 3290
rect 1275 3286 1343 3290
rect 1347 3286 1407 3290
rect 1411 3286 1519 3290
rect 1523 3286 1551 3290
rect 1555 3286 1823 3290
rect 1827 3286 1835 3290
rect 91 3285 1835 3286
rect 1841 3290 3606 3291
rect 1841 3286 1863 3290
rect 1867 3286 1887 3290
rect 1891 3286 2039 3290
rect 2043 3286 2063 3290
rect 2067 3286 2199 3290
rect 2203 3286 2263 3290
rect 2267 3286 2359 3290
rect 2363 3286 2455 3290
rect 2459 3286 2527 3290
rect 2531 3286 2639 3290
rect 2643 3286 2695 3290
rect 2699 3286 2815 3290
rect 2819 3286 2871 3290
rect 2875 3286 2983 3290
rect 2987 3286 3047 3290
rect 3051 3286 3151 3290
rect 3155 3286 3319 3290
rect 3323 3286 3479 3290
rect 3483 3286 3575 3290
rect 3579 3286 3606 3290
rect 1841 3285 3606 3286
rect 294 3268 300 3269
rect 618 3268 624 3269
rect 294 3264 295 3268
rect 299 3264 619 3268
rect 623 3264 624 3268
rect 294 3263 300 3264
rect 618 3263 624 3264
rect 462 3236 468 3237
rect 738 3236 744 3237
rect 462 3232 463 3236
rect 467 3232 739 3236
rect 743 3232 744 3236
rect 462 3231 468 3232
rect 738 3231 744 3232
rect 1846 3222 3618 3223
rect 1846 3219 1863 3222
rect 96 3213 97 3219
rect 103 3218 1847 3219
rect 103 3214 111 3218
rect 115 3214 263 3218
rect 267 3214 383 3218
rect 387 3214 431 3218
rect 435 3214 519 3218
rect 523 3214 551 3218
rect 555 3214 671 3218
rect 675 3214 799 3218
rect 803 3214 831 3218
rect 835 3214 935 3218
rect 939 3214 999 3218
rect 1003 3214 1079 3218
rect 1083 3214 1175 3218
rect 1179 3214 1231 3218
rect 1235 3214 1351 3218
rect 1355 3214 1383 3218
rect 1387 3214 1527 3218
rect 1531 3214 1535 3218
rect 1539 3214 1823 3218
rect 1827 3214 1847 3218
rect 103 3213 1847 3214
rect 1853 3218 1863 3219
rect 1867 3218 1895 3222
rect 1899 3218 2071 3222
rect 2075 3218 2087 3222
rect 2091 3218 2271 3222
rect 2275 3218 2303 3222
rect 2307 3218 2463 3222
rect 2467 3218 2511 3222
rect 2515 3218 2647 3222
rect 2651 3218 2703 3222
rect 2707 3218 2823 3222
rect 2827 3218 2879 3222
rect 2883 3218 2991 3222
rect 2995 3218 3039 3222
rect 3043 3218 3159 3222
rect 3163 3218 3199 3222
rect 3203 3218 3327 3222
rect 3331 3218 3351 3222
rect 3355 3218 3487 3222
rect 3491 3218 3575 3222
rect 3579 3218 3618 3222
rect 1853 3217 3618 3218
rect 1853 3213 1854 3217
rect 1834 3150 3606 3151
rect 1834 3147 1863 3150
rect 84 3141 85 3147
rect 91 3146 1835 3147
rect 91 3142 111 3146
rect 115 3142 423 3146
rect 427 3142 463 3146
rect 467 3142 543 3146
rect 547 3142 551 3146
rect 555 3142 639 3146
rect 643 3142 663 3146
rect 667 3142 735 3146
rect 739 3142 791 3146
rect 795 3142 847 3146
rect 851 3142 927 3146
rect 931 3142 967 3146
rect 971 3142 1071 3146
rect 1075 3142 1095 3146
rect 1099 3142 1223 3146
rect 1227 3142 1231 3146
rect 1235 3142 1375 3146
rect 1379 3142 1519 3146
rect 1523 3142 1527 3146
rect 1531 3142 1823 3146
rect 1827 3142 1835 3146
rect 91 3141 1835 3142
rect 1841 3146 1863 3147
rect 1867 3146 1887 3150
rect 1891 3146 2079 3150
rect 2083 3146 2295 3150
rect 2299 3146 2503 3150
rect 2507 3146 2695 3150
rect 2699 3146 2871 3150
rect 2875 3146 3031 3150
rect 3035 3146 3039 3150
rect 3043 3146 3191 3150
rect 3195 3146 3343 3150
rect 3347 3146 3479 3150
rect 3483 3146 3575 3150
rect 3579 3146 3606 3150
rect 1841 3145 3606 3146
rect 1841 3141 1842 3145
rect 96 3065 97 3071
rect 103 3070 1847 3071
rect 103 3066 111 3070
rect 115 3066 151 3070
rect 155 3066 239 3070
rect 243 3066 327 3070
rect 331 3066 415 3070
rect 419 3066 471 3070
rect 475 3066 503 3070
rect 507 3066 559 3070
rect 563 3066 591 3070
rect 595 3066 647 3070
rect 651 3066 679 3070
rect 683 3066 743 3070
rect 747 3066 767 3070
rect 771 3066 855 3070
rect 859 3066 943 3070
rect 947 3066 975 3070
rect 979 3066 1031 3070
rect 1035 3066 1103 3070
rect 1107 3066 1119 3070
rect 1123 3066 1207 3070
rect 1211 3066 1239 3070
rect 1243 3066 1295 3070
rect 1299 3066 1383 3070
rect 1387 3066 1471 3070
rect 1475 3066 1527 3070
rect 1531 3066 1559 3070
rect 1563 3066 1647 3070
rect 1651 3066 1735 3070
rect 1739 3066 1823 3070
rect 1827 3066 1847 3070
rect 103 3065 1847 3066
rect 1853 3070 3618 3071
rect 1853 3066 1863 3070
rect 1867 3066 1895 3070
rect 1899 3066 2087 3070
rect 2091 3066 2255 3070
rect 2259 3066 2303 3070
rect 2307 3066 2423 3070
rect 2427 3066 2511 3070
rect 2515 3066 2591 3070
rect 2595 3066 2703 3070
rect 2707 3066 2751 3070
rect 2755 3066 2879 3070
rect 2883 3066 2919 3070
rect 2923 3066 3047 3070
rect 3051 3066 3087 3070
rect 3091 3066 3199 3070
rect 3203 3066 3351 3070
rect 3355 3066 3487 3070
rect 3491 3066 3575 3070
rect 3579 3066 3618 3070
rect 1853 3065 3618 3066
rect 222 3060 228 3061
rect 914 3060 920 3061
rect 222 3056 223 3060
rect 227 3056 915 3060
rect 919 3056 920 3060
rect 222 3055 228 3056
rect 914 3055 920 3056
rect 2782 3060 2788 3061
rect 3034 3060 3040 3061
rect 2782 3056 2783 3060
rect 2787 3056 3035 3060
rect 3039 3056 3040 3060
rect 2782 3055 2788 3056
rect 3034 3055 3040 3056
rect 1834 2998 3606 2999
rect 1834 2995 1863 2998
rect 84 2989 85 2995
rect 91 2994 1835 2995
rect 91 2990 111 2994
rect 115 2990 143 2994
rect 147 2990 231 2994
rect 235 2990 319 2994
rect 323 2990 407 2994
rect 411 2990 495 2994
rect 499 2990 583 2994
rect 587 2990 671 2994
rect 675 2990 759 2994
rect 763 2990 847 2994
rect 851 2990 935 2994
rect 939 2990 1023 2994
rect 1027 2990 1111 2994
rect 1115 2990 1199 2994
rect 1203 2990 1287 2994
rect 1291 2990 1375 2994
rect 1379 2990 1407 2994
rect 1411 2990 1463 2994
rect 1467 2990 1519 2994
rect 1523 2990 1551 2994
rect 1555 2990 1631 2994
rect 1635 2990 1639 2994
rect 1643 2990 1727 2994
rect 1731 2990 1823 2994
rect 1827 2990 1835 2994
rect 91 2989 1835 2990
rect 1841 2994 1863 2995
rect 1867 2994 2239 2998
rect 2243 2994 2247 2998
rect 2251 2994 2415 2998
rect 2419 2994 2463 2998
rect 2467 2994 2583 2998
rect 2587 2994 2671 2998
rect 2675 2994 2743 2998
rect 2747 2994 2863 2998
rect 2867 2994 2911 2998
rect 2915 2994 3031 2998
rect 3035 2994 3079 2998
rect 3083 2994 3191 2998
rect 3195 2994 3343 2998
rect 3347 2994 3479 2998
rect 3483 2994 3575 2998
rect 3579 2994 3606 2998
rect 1841 2993 3606 2994
rect 1841 2989 1842 2993
rect 2710 2940 2716 2941
rect 2958 2940 2964 2941
rect 2710 2936 2711 2940
rect 2715 2936 2959 2940
rect 2963 2936 2964 2940
rect 2710 2935 2716 2936
rect 2958 2935 2964 2936
rect 96 2921 97 2927
rect 103 2926 1847 2927
rect 103 2922 111 2926
rect 115 2922 1359 2926
rect 1363 2922 1415 2926
rect 1419 2922 1471 2926
rect 1475 2922 1527 2926
rect 1531 2922 1583 2926
rect 1587 2922 1639 2926
rect 1643 2922 1703 2926
rect 1707 2922 1735 2926
rect 1739 2922 1823 2926
rect 1827 2922 1847 2926
rect 103 2921 1847 2922
rect 1853 2921 1854 2927
rect 1846 2909 1847 2915
rect 1853 2914 3611 2915
rect 1853 2910 1863 2914
rect 1867 2910 2239 2914
rect 2243 2910 2247 2914
rect 2251 2910 2463 2914
rect 2467 2910 2471 2914
rect 2475 2910 2671 2914
rect 2675 2910 2679 2914
rect 2683 2910 2855 2914
rect 2859 2910 2871 2914
rect 2875 2910 3023 2914
rect 3027 2910 3039 2914
rect 3043 2910 3183 2914
rect 3187 2910 3199 2914
rect 3203 2910 3335 2914
rect 3339 2910 3351 2914
rect 3355 2910 3487 2914
rect 3491 2910 3575 2914
rect 3579 2910 3611 2914
rect 1853 2909 3611 2910
rect 3617 2909 3618 2915
rect 2750 2868 2756 2869
rect 3098 2868 3104 2869
rect 2750 2864 2751 2868
rect 2755 2864 3099 2868
rect 3103 2864 3104 2868
rect 2750 2863 2756 2864
rect 3098 2863 3104 2864
rect 84 2849 85 2855
rect 91 2854 1835 2855
rect 91 2850 111 2854
rect 115 2850 135 2854
rect 139 2850 223 2854
rect 227 2850 311 2854
rect 315 2850 399 2854
rect 403 2850 487 2854
rect 491 2850 599 2854
rect 603 2850 727 2854
rect 731 2850 863 2854
rect 867 2850 999 2854
rect 1003 2850 1135 2854
rect 1139 2850 1263 2854
rect 1267 2850 1351 2854
rect 1355 2850 1383 2854
rect 1387 2850 1463 2854
rect 1467 2850 1503 2854
rect 1507 2850 1575 2854
rect 1579 2850 1623 2854
rect 1627 2850 1695 2854
rect 1699 2850 1727 2854
rect 1731 2850 1823 2854
rect 1827 2850 1835 2854
rect 91 2849 1835 2850
rect 1841 2849 1842 2855
rect 1834 2837 1835 2843
rect 1841 2842 3599 2843
rect 1841 2838 1863 2842
rect 1867 2838 1895 2842
rect 1899 2838 1983 2842
rect 1987 2838 2071 2842
rect 2075 2838 2159 2842
rect 2163 2838 2231 2842
rect 2235 2838 2247 2842
rect 2251 2838 2335 2842
rect 2339 2838 2423 2842
rect 2427 2838 2455 2842
rect 2459 2838 2511 2842
rect 2515 2838 2599 2842
rect 2603 2838 2663 2842
rect 2667 2838 2687 2842
rect 2691 2838 2791 2842
rect 2795 2838 2847 2842
rect 2851 2838 2903 2842
rect 2907 2838 3015 2842
rect 3019 2838 3031 2842
rect 3035 2838 3175 2842
rect 3179 2838 3327 2842
rect 3331 2838 3479 2842
rect 3483 2838 3575 2842
rect 3579 2838 3599 2842
rect 1841 2837 3599 2838
rect 3605 2837 3606 2843
rect 96 2781 97 2787
rect 103 2786 1847 2787
rect 103 2782 111 2786
rect 115 2782 143 2786
rect 147 2782 191 2786
rect 195 2782 231 2786
rect 235 2782 295 2786
rect 299 2782 319 2786
rect 323 2782 407 2786
rect 411 2782 415 2786
rect 419 2782 495 2786
rect 499 2782 551 2786
rect 555 2782 607 2786
rect 611 2782 687 2786
rect 691 2782 735 2786
rect 739 2782 823 2786
rect 827 2782 871 2786
rect 875 2782 959 2786
rect 963 2782 1007 2786
rect 1011 2782 1087 2786
rect 1091 2782 1143 2786
rect 1147 2782 1207 2786
rect 1211 2782 1271 2786
rect 1275 2782 1319 2786
rect 1323 2782 1391 2786
rect 1395 2782 1431 2786
rect 1435 2782 1511 2786
rect 1515 2782 1535 2786
rect 1539 2782 1631 2786
rect 1635 2782 1647 2786
rect 1651 2782 1735 2786
rect 1739 2782 1823 2786
rect 1827 2782 1847 2786
rect 103 2781 1847 2782
rect 1853 2781 1854 2787
rect 1846 2757 1847 2763
rect 1853 2762 3611 2763
rect 1853 2758 1863 2762
rect 1867 2758 1903 2762
rect 1907 2758 1991 2762
rect 1995 2758 2047 2762
rect 2051 2758 2079 2762
rect 2083 2758 2167 2762
rect 2171 2758 2255 2762
rect 2259 2758 2295 2762
rect 2299 2758 2343 2762
rect 2347 2758 2431 2762
rect 2435 2758 2447 2762
rect 2451 2758 2519 2762
rect 2523 2758 2607 2762
rect 2611 2758 2623 2762
rect 2627 2758 2695 2762
rect 2699 2758 2799 2762
rect 2803 2758 2823 2762
rect 2827 2758 2911 2762
rect 2915 2758 3039 2762
rect 3043 2758 3183 2762
rect 3187 2758 3271 2762
rect 3275 2758 3335 2762
rect 3339 2758 3487 2762
rect 3491 2758 3575 2762
rect 3579 2758 3611 2762
rect 1853 2757 3611 2758
rect 3617 2757 3618 2763
rect 84 2705 85 2711
rect 91 2710 1835 2711
rect 91 2706 111 2710
rect 115 2706 167 2710
rect 171 2706 183 2710
rect 187 2706 279 2710
rect 283 2706 287 2710
rect 291 2706 391 2710
rect 395 2706 407 2710
rect 411 2706 503 2710
rect 507 2706 543 2710
rect 547 2706 615 2710
rect 619 2706 679 2710
rect 683 2706 815 2710
rect 819 2706 951 2710
rect 955 2706 1079 2710
rect 1083 2706 1199 2710
rect 1203 2706 1311 2710
rect 1315 2706 1423 2710
rect 1427 2706 1527 2710
rect 1531 2706 1639 2710
rect 1643 2706 1727 2710
rect 1731 2706 1823 2710
rect 1827 2706 1835 2710
rect 91 2705 1835 2706
rect 1841 2705 1842 2711
rect 1834 2689 1835 2695
rect 1841 2694 3599 2695
rect 1841 2690 1863 2694
rect 1867 2690 1943 2694
rect 1947 2690 2039 2694
rect 2043 2690 2055 2694
rect 2059 2690 2159 2694
rect 2163 2690 2167 2694
rect 2171 2690 2287 2694
rect 2291 2690 2407 2694
rect 2411 2690 2439 2694
rect 2443 2690 2519 2694
rect 2523 2690 2615 2694
rect 2619 2690 2631 2694
rect 2635 2690 2735 2694
rect 2739 2690 2815 2694
rect 2819 2690 2847 2694
rect 2851 2690 2959 2694
rect 2963 2690 3031 2694
rect 3035 2690 3071 2694
rect 3075 2690 3263 2694
rect 3267 2690 3479 2694
rect 3483 2690 3575 2694
rect 3579 2690 3599 2694
rect 1841 2689 3599 2690
rect 3605 2689 3606 2695
rect 96 2621 97 2627
rect 103 2626 1847 2627
rect 103 2622 111 2626
rect 115 2622 175 2626
rect 179 2622 223 2626
rect 227 2622 287 2626
rect 291 2622 351 2626
rect 355 2622 399 2626
rect 403 2622 495 2626
rect 499 2622 511 2626
rect 515 2622 623 2626
rect 627 2622 663 2626
rect 667 2622 839 2626
rect 843 2622 1023 2626
rect 1027 2622 1215 2626
rect 1219 2622 1407 2626
rect 1411 2622 1607 2626
rect 1611 2622 1823 2626
rect 1827 2622 1847 2626
rect 103 2621 1847 2622
rect 1853 2623 1854 2627
rect 1853 2622 3618 2623
rect 1853 2621 1863 2622
rect 1846 2618 1863 2621
rect 1867 2618 1895 2622
rect 1899 2618 1951 2622
rect 1955 2618 2063 2622
rect 2067 2618 2071 2622
rect 2075 2618 2175 2622
rect 2179 2618 2263 2622
rect 2267 2618 2295 2622
rect 2299 2618 2415 2622
rect 2419 2618 2463 2622
rect 2467 2618 2527 2622
rect 2531 2618 2639 2622
rect 2643 2618 2663 2622
rect 2667 2618 2743 2622
rect 2747 2618 2855 2622
rect 2859 2618 2871 2622
rect 2875 2618 2967 2622
rect 2971 2618 3079 2622
rect 3083 2618 3295 2622
rect 3299 2618 3487 2622
rect 3491 2618 3575 2622
rect 3579 2618 3618 2622
rect 1846 2617 3618 2618
rect 84 2553 85 2559
rect 91 2558 1835 2559
rect 91 2554 111 2558
rect 115 2554 215 2558
rect 219 2554 271 2558
rect 275 2554 343 2558
rect 347 2554 471 2558
rect 475 2554 487 2558
rect 491 2554 655 2558
rect 659 2554 671 2558
rect 675 2554 831 2558
rect 835 2554 855 2558
rect 859 2554 1015 2558
rect 1019 2554 1023 2558
rect 1027 2554 1175 2558
rect 1179 2554 1207 2558
rect 1211 2554 1319 2558
rect 1323 2554 1399 2558
rect 1403 2554 1455 2558
rect 1459 2554 1591 2558
rect 1595 2554 1599 2558
rect 1603 2554 1727 2558
rect 1731 2554 1823 2558
rect 1827 2554 1835 2558
rect 91 2553 1835 2554
rect 1841 2555 1842 2559
rect 1841 2554 3606 2555
rect 1841 2553 1863 2554
rect 1834 2550 1863 2553
rect 1867 2550 1887 2554
rect 1891 2550 2039 2554
rect 2043 2550 2063 2554
rect 2067 2550 2215 2554
rect 2219 2550 2255 2554
rect 2259 2550 2399 2554
rect 2403 2550 2455 2554
rect 2459 2550 2575 2554
rect 2579 2550 2655 2554
rect 2659 2550 2743 2554
rect 2747 2550 2863 2554
rect 2867 2550 2903 2554
rect 2907 2550 3055 2554
rect 3059 2550 3071 2554
rect 3075 2550 3199 2554
rect 3203 2550 3287 2554
rect 3291 2550 3343 2554
rect 3347 2550 3479 2554
rect 3483 2550 3575 2554
rect 3579 2550 3606 2554
rect 1834 2549 3606 2550
rect 96 2481 97 2487
rect 103 2486 1847 2487
rect 103 2482 111 2486
rect 115 2482 183 2486
rect 187 2482 279 2486
rect 283 2482 319 2486
rect 323 2482 463 2486
rect 467 2482 479 2486
rect 483 2482 607 2486
rect 611 2482 679 2486
rect 683 2482 743 2486
rect 747 2482 863 2486
rect 867 2482 879 2486
rect 883 2482 1007 2486
rect 1011 2482 1031 2486
rect 1035 2482 1127 2486
rect 1131 2482 1183 2486
rect 1187 2482 1239 2486
rect 1243 2482 1327 2486
rect 1331 2482 1343 2486
rect 1347 2482 1447 2486
rect 1451 2482 1463 2486
rect 1467 2482 1551 2486
rect 1555 2482 1599 2486
rect 1603 2482 1647 2486
rect 1651 2482 1735 2486
rect 1739 2482 1823 2486
rect 1827 2482 1847 2486
rect 103 2481 1847 2482
rect 1853 2486 3618 2487
rect 1853 2482 1863 2486
rect 1867 2482 1895 2486
rect 1899 2482 1991 2486
rect 1995 2482 2047 2486
rect 2051 2482 2127 2486
rect 2131 2482 2223 2486
rect 2227 2482 2279 2486
rect 2283 2482 2407 2486
rect 2411 2482 2439 2486
rect 2443 2482 2583 2486
rect 2587 2482 2599 2486
rect 2603 2482 2751 2486
rect 2755 2482 2767 2486
rect 2771 2482 2911 2486
rect 2915 2482 2943 2486
rect 2947 2482 3063 2486
rect 3067 2482 3119 2486
rect 3123 2482 3207 2486
rect 3211 2482 3295 2486
rect 3299 2482 3351 2486
rect 3355 2482 3471 2486
rect 3475 2482 3487 2486
rect 3491 2482 3575 2486
rect 3579 2482 3618 2486
rect 1853 2481 3618 2482
rect 84 2405 85 2411
rect 91 2410 1835 2411
rect 91 2406 111 2410
rect 115 2406 151 2410
rect 155 2406 175 2410
rect 179 2406 311 2410
rect 315 2406 319 2410
rect 323 2406 455 2410
rect 459 2406 479 2410
rect 483 2406 599 2410
rect 603 2406 639 2410
rect 643 2406 735 2410
rect 739 2406 783 2410
rect 787 2406 871 2410
rect 875 2406 919 2410
rect 923 2406 999 2410
rect 1003 2406 1047 2410
rect 1051 2406 1119 2410
rect 1123 2406 1175 2410
rect 1179 2406 1231 2410
rect 1235 2406 1303 2410
rect 1307 2406 1335 2410
rect 1339 2406 1431 2410
rect 1435 2406 1439 2410
rect 1443 2406 1543 2410
rect 1547 2406 1639 2410
rect 1643 2406 1727 2410
rect 1731 2406 1823 2410
rect 1827 2406 1835 2410
rect 91 2405 1835 2406
rect 1841 2410 3606 2411
rect 1841 2406 1863 2410
rect 1867 2406 1887 2410
rect 1891 2406 1983 2410
rect 1987 2406 2119 2410
rect 2123 2406 2271 2410
rect 2275 2406 2351 2410
rect 2355 2406 2431 2410
rect 2435 2406 2503 2410
rect 2507 2406 2591 2410
rect 2595 2406 2655 2410
rect 2659 2406 2759 2410
rect 2763 2406 2807 2410
rect 2811 2406 2935 2410
rect 2939 2406 2967 2410
rect 2971 2406 3111 2410
rect 3115 2406 3135 2410
rect 3139 2406 3287 2410
rect 3291 2406 3303 2410
rect 3307 2406 3463 2410
rect 3467 2406 3471 2410
rect 3475 2406 3575 2410
rect 3579 2406 3606 2410
rect 1841 2405 3606 2406
rect 96 2333 97 2339
rect 103 2338 1847 2339
rect 103 2334 111 2338
rect 115 2334 143 2338
rect 147 2334 159 2338
rect 163 2334 263 2338
rect 267 2334 327 2338
rect 331 2334 407 2338
rect 411 2334 487 2338
rect 491 2334 543 2338
rect 547 2334 647 2338
rect 651 2334 679 2338
rect 683 2334 791 2338
rect 795 2334 807 2338
rect 811 2334 927 2338
rect 931 2334 1039 2338
rect 1043 2334 1055 2338
rect 1059 2334 1159 2338
rect 1163 2334 1183 2338
rect 1187 2334 1279 2338
rect 1283 2334 1311 2338
rect 1315 2334 1439 2338
rect 1443 2334 1823 2338
rect 1827 2334 1847 2338
rect 103 2333 1847 2334
rect 1853 2338 3618 2339
rect 1853 2334 1863 2338
rect 1867 2334 2351 2338
rect 2355 2334 2359 2338
rect 2363 2334 2447 2338
rect 2451 2334 2511 2338
rect 2515 2334 2559 2338
rect 2563 2334 2663 2338
rect 2667 2334 2703 2338
rect 2707 2334 2815 2338
rect 2819 2334 2879 2338
rect 2883 2334 2975 2338
rect 2979 2334 3079 2338
rect 3083 2334 3143 2338
rect 3147 2334 3287 2338
rect 3291 2334 3311 2338
rect 3315 2334 3479 2338
rect 3483 2334 3487 2338
rect 3491 2334 3575 2338
rect 3579 2334 3618 2338
rect 1853 2333 3618 2334
rect 1026 2316 1032 2317
rect 1226 2316 1232 2317
rect 1026 2312 1027 2316
rect 1031 2312 1227 2316
rect 1231 2312 1232 2316
rect 1026 2311 1032 2312
rect 1226 2311 1232 2312
rect 84 2265 85 2271
rect 91 2270 1835 2271
rect 91 2266 111 2270
rect 115 2266 135 2270
rect 139 2266 231 2270
rect 235 2266 255 2270
rect 259 2266 351 2270
rect 355 2266 399 2270
rect 403 2266 471 2270
rect 475 2266 535 2270
rect 539 2266 591 2270
rect 595 2266 671 2270
rect 675 2266 711 2270
rect 715 2266 799 2270
rect 803 2266 823 2270
rect 827 2266 919 2270
rect 923 2266 935 2270
rect 939 2266 1031 2270
rect 1035 2266 1055 2270
rect 1059 2266 1151 2270
rect 1155 2266 1175 2270
rect 1179 2266 1271 2270
rect 1275 2266 1823 2270
rect 1827 2266 1835 2270
rect 91 2265 1835 2266
rect 1841 2270 3606 2271
rect 1841 2266 1863 2270
rect 1867 2266 2335 2270
rect 2339 2266 2343 2270
rect 2347 2266 2439 2270
rect 2443 2266 2447 2270
rect 2451 2266 2551 2270
rect 2555 2266 2583 2270
rect 2587 2266 2695 2270
rect 2699 2266 2735 2270
rect 2739 2266 2871 2270
rect 2875 2266 2911 2270
rect 2915 2266 3071 2270
rect 3075 2266 3103 2270
rect 3107 2266 3279 2270
rect 3283 2266 3303 2270
rect 3307 2266 3479 2270
rect 3483 2266 3575 2270
rect 3579 2266 3606 2270
rect 1841 2265 3606 2266
rect 1846 2202 3618 2203
rect 1846 2199 1863 2202
rect 96 2193 97 2199
rect 103 2198 1847 2199
rect 103 2194 111 2198
rect 115 2194 143 2198
rect 147 2194 239 2198
rect 243 2194 247 2198
rect 251 2194 359 2198
rect 363 2194 383 2198
rect 387 2194 479 2198
rect 483 2194 519 2198
rect 523 2194 599 2198
rect 603 2194 655 2198
rect 659 2194 719 2198
rect 723 2194 783 2198
rect 787 2194 831 2198
rect 835 2194 911 2198
rect 915 2194 943 2198
rect 947 2194 1031 2198
rect 1035 2194 1063 2198
rect 1067 2194 1159 2198
rect 1163 2194 1183 2198
rect 1187 2194 1287 2198
rect 1291 2194 1823 2198
rect 1827 2194 1847 2198
rect 103 2193 1847 2194
rect 1853 2198 1863 2199
rect 1867 2198 2255 2202
rect 2259 2198 2343 2202
rect 2347 2198 2439 2202
rect 2443 2198 2455 2202
rect 2459 2198 2551 2202
rect 2555 2198 2591 2202
rect 2595 2198 2695 2202
rect 2699 2198 2743 2202
rect 2747 2198 2871 2202
rect 2875 2198 2919 2202
rect 2923 2198 3071 2202
rect 3075 2198 3111 2202
rect 3115 2198 3287 2202
rect 3291 2198 3311 2202
rect 3315 2198 3487 2202
rect 3491 2198 3575 2202
rect 3579 2198 3618 2202
rect 1853 2197 3618 2198
rect 1853 2193 1854 2197
rect 1834 2126 3606 2127
rect 1834 2123 1863 2126
rect 84 2117 85 2123
rect 91 2122 1835 2123
rect 91 2118 111 2122
rect 115 2118 135 2122
rect 139 2118 231 2122
rect 235 2118 239 2122
rect 243 2118 359 2122
rect 363 2118 375 2122
rect 379 2118 479 2122
rect 483 2118 511 2122
rect 515 2118 599 2122
rect 603 2118 647 2122
rect 651 2118 719 2122
rect 723 2118 775 2122
rect 779 2118 831 2122
rect 835 2118 903 2122
rect 907 2118 943 2122
rect 947 2118 1023 2122
rect 1027 2118 1055 2122
rect 1059 2118 1151 2122
rect 1155 2118 1175 2122
rect 1179 2118 1279 2122
rect 1283 2118 1823 2122
rect 1827 2118 1835 2122
rect 91 2117 1835 2118
rect 1841 2122 1863 2123
rect 1867 2122 2151 2126
rect 2155 2122 2239 2126
rect 2243 2122 2247 2126
rect 2251 2122 2327 2126
rect 2331 2122 2335 2126
rect 2339 2122 2415 2126
rect 2419 2122 2431 2126
rect 2435 2122 2503 2126
rect 2507 2122 2543 2126
rect 2547 2122 2615 2126
rect 2619 2122 2687 2126
rect 2691 2122 2751 2126
rect 2755 2122 2863 2126
rect 2867 2122 2919 2126
rect 2923 2122 3063 2126
rect 3067 2122 3103 2126
rect 3107 2122 3279 2126
rect 3283 2122 3303 2126
rect 3307 2122 3479 2126
rect 3483 2122 3575 2126
rect 3579 2122 3606 2126
rect 1841 2121 3606 2122
rect 1841 2117 1842 2121
rect 2662 2108 2668 2109
rect 3198 2108 3204 2109
rect 2662 2104 2663 2108
rect 2667 2104 3199 2108
rect 3203 2104 3204 2108
rect 2662 2103 2668 2104
rect 3198 2103 3204 2104
rect 2190 2068 2196 2069
rect 2482 2068 2488 2069
rect 2190 2064 2191 2068
rect 2195 2064 2483 2068
rect 2487 2064 2488 2068
rect 2190 2063 2196 2064
rect 2482 2063 2488 2064
rect 1846 2049 1847 2055
rect 1853 2054 3611 2055
rect 1853 2050 1863 2054
rect 1867 2050 1999 2054
rect 2003 2050 2127 2054
rect 2131 2050 2159 2054
rect 2163 2050 2247 2054
rect 2251 2050 2255 2054
rect 2259 2050 2335 2054
rect 2339 2050 2399 2054
rect 2403 2050 2423 2054
rect 2427 2050 2511 2054
rect 2515 2050 2551 2054
rect 2555 2050 2623 2054
rect 2627 2050 2711 2054
rect 2715 2050 2759 2054
rect 2763 2050 2879 2054
rect 2883 2050 2927 2054
rect 2931 2050 3063 2054
rect 3067 2050 3111 2054
rect 3115 2050 3247 2054
rect 3251 2050 3311 2054
rect 3315 2050 3439 2054
rect 3443 2050 3487 2054
rect 3491 2050 3575 2054
rect 3579 2050 3611 2054
rect 1853 2049 3611 2050
rect 3617 2049 3618 2055
rect 96 2037 97 2043
rect 103 2042 1847 2043
rect 103 2038 111 2042
rect 115 2038 143 2042
rect 147 2038 167 2042
rect 171 2038 239 2042
rect 243 2038 311 2042
rect 315 2038 367 2042
rect 371 2038 447 2042
rect 451 2038 487 2042
rect 491 2038 575 2042
rect 579 2038 607 2042
rect 611 2038 695 2042
rect 699 2038 727 2042
rect 731 2038 807 2042
rect 811 2038 839 2042
rect 843 2038 911 2042
rect 915 2038 951 2042
rect 955 2038 1015 2042
rect 1019 2038 1063 2042
rect 1067 2038 1119 2042
rect 1123 2038 1183 2042
rect 1187 2038 1223 2042
rect 1227 2038 1327 2042
rect 1331 2038 1823 2042
rect 1827 2038 1847 2042
rect 103 2037 1847 2038
rect 1853 2037 1854 2043
rect 2070 2020 2076 2021
rect 2478 2020 2484 2021
rect 2070 2016 2071 2020
rect 2075 2016 2479 2020
rect 2483 2016 2484 2020
rect 2070 2015 2076 2016
rect 2478 2015 2484 2016
rect 1834 1978 3606 1979
rect 1834 1975 1863 1978
rect 84 1969 85 1975
rect 91 1974 1835 1975
rect 91 1970 111 1974
rect 115 1970 159 1974
rect 163 1970 295 1974
rect 299 1970 303 1974
rect 307 1970 439 1974
rect 443 1970 567 1974
rect 571 1970 583 1974
rect 587 1970 687 1974
rect 691 1970 719 1974
rect 723 1970 799 1974
rect 803 1970 855 1974
rect 859 1970 903 1974
rect 907 1970 991 1974
rect 995 1970 1007 1974
rect 1011 1970 1111 1974
rect 1115 1970 1119 1974
rect 1123 1970 1215 1974
rect 1219 1970 1239 1974
rect 1243 1970 1319 1974
rect 1323 1970 1359 1974
rect 1363 1970 1479 1974
rect 1483 1970 1599 1974
rect 1603 1970 1823 1974
rect 1827 1970 1835 1974
rect 91 1969 1835 1970
rect 1841 1974 1863 1975
rect 1867 1974 1903 1978
rect 1907 1974 1991 1978
rect 1995 1974 2119 1978
rect 2123 1974 2159 1978
rect 2163 1974 2247 1978
rect 2251 1974 2391 1978
rect 2395 1974 2399 1978
rect 2403 1974 2543 1978
rect 2547 1974 2615 1978
rect 2619 1974 2703 1978
rect 2707 1974 2815 1978
rect 2819 1974 2871 1978
rect 2875 1974 2999 1978
rect 3003 1974 3055 1978
rect 3059 1974 3167 1978
rect 3171 1974 3239 1978
rect 3243 1974 3335 1978
rect 3339 1974 3431 1978
rect 3435 1974 3479 1978
rect 3483 1974 3575 1978
rect 3579 1974 3606 1978
rect 1841 1973 3606 1974
rect 1841 1969 1842 1973
rect 2654 1940 2660 1941
rect 3150 1940 3156 1941
rect 2654 1936 2655 1940
rect 2659 1936 3151 1940
rect 3155 1936 3156 1940
rect 2654 1935 2660 1936
rect 3150 1935 3156 1936
rect 2950 1924 2956 1925
rect 3258 1924 3264 1925
rect 2950 1920 2951 1924
rect 2955 1920 3259 1924
rect 3263 1920 3264 1924
rect 2950 1919 2956 1920
rect 3258 1919 3264 1920
rect 1846 1905 1847 1911
rect 1853 1910 3611 1911
rect 1853 1906 1863 1910
rect 1867 1906 1895 1910
rect 1899 1906 1911 1910
rect 1915 1906 1983 1910
rect 1987 1906 2071 1910
rect 2075 1906 2167 1910
rect 2171 1906 2295 1910
rect 2299 1906 2407 1910
rect 2411 1906 2447 1910
rect 2451 1906 2607 1910
rect 2611 1906 2623 1910
rect 2627 1906 2767 1910
rect 2771 1906 2823 1910
rect 2827 1906 2919 1910
rect 2923 1906 3007 1910
rect 3011 1906 3071 1910
rect 3075 1906 3175 1910
rect 3179 1906 3215 1910
rect 3219 1906 3343 1910
rect 3347 1906 3359 1910
rect 3363 1906 3487 1910
rect 3491 1906 3575 1910
rect 3579 1906 3611 1910
rect 1853 1905 3611 1906
rect 3617 1905 3618 1911
rect 96 1893 97 1899
rect 103 1898 1847 1899
rect 103 1894 111 1898
rect 115 1894 167 1898
rect 171 1894 223 1898
rect 227 1894 303 1898
rect 307 1894 447 1898
rect 451 1894 479 1898
rect 483 1894 591 1898
rect 595 1894 719 1898
rect 723 1894 727 1898
rect 731 1894 863 1898
rect 867 1894 935 1898
rect 939 1894 999 1898
rect 1003 1894 1127 1898
rect 1131 1894 1247 1898
rect 1251 1894 1295 1898
rect 1299 1894 1367 1898
rect 1371 1894 1455 1898
rect 1459 1894 1487 1898
rect 1491 1894 1607 1898
rect 1611 1894 1735 1898
rect 1739 1894 1823 1898
rect 1827 1894 1847 1898
rect 103 1893 1847 1894
rect 1853 1893 1854 1899
rect 1942 1884 1948 1885
rect 2402 1884 2408 1885
rect 1942 1880 1943 1884
rect 1947 1880 2403 1884
rect 2407 1880 2408 1884
rect 1942 1879 1948 1880
rect 2402 1879 2408 1880
rect 1834 1833 1835 1839
rect 1841 1838 3599 1839
rect 1841 1834 1863 1838
rect 1867 1834 1887 1838
rect 1891 1834 1975 1838
rect 1979 1834 1999 1838
rect 2003 1834 2063 1838
rect 2067 1834 2159 1838
rect 2163 1834 2223 1838
rect 2227 1834 2287 1838
rect 2291 1834 2439 1838
rect 2443 1834 2599 1838
rect 2603 1834 2639 1838
rect 2643 1834 2759 1838
rect 2763 1834 2831 1838
rect 2835 1834 2911 1838
rect 2915 1834 3015 1838
rect 3019 1834 3063 1838
rect 3067 1834 3199 1838
rect 3203 1834 3207 1838
rect 3211 1834 3351 1838
rect 3355 1834 3391 1838
rect 3395 1834 3479 1838
rect 3483 1834 3575 1838
rect 3579 1834 3599 1838
rect 1841 1833 3599 1834
rect 3605 1833 3606 1839
rect 1834 1831 1842 1833
rect 84 1825 85 1831
rect 91 1830 1835 1831
rect 91 1826 111 1830
rect 115 1826 215 1830
rect 219 1826 247 1830
rect 251 1826 415 1830
rect 419 1826 471 1830
rect 475 1826 591 1830
rect 595 1826 711 1830
rect 715 1826 759 1830
rect 763 1826 927 1830
rect 931 1826 1079 1830
rect 1083 1826 1119 1830
rect 1123 1826 1223 1830
rect 1227 1826 1287 1830
rect 1291 1826 1359 1830
rect 1363 1826 1447 1830
rect 1451 1826 1487 1830
rect 1491 1826 1599 1830
rect 1603 1826 1615 1830
rect 1619 1826 1727 1830
rect 1731 1826 1823 1830
rect 1827 1826 1835 1830
rect 91 1825 1835 1826
rect 1841 1825 1842 1831
rect 2262 1796 2268 1797
rect 2674 1796 2680 1797
rect 2262 1792 2263 1796
rect 2267 1792 2675 1796
rect 2679 1792 2680 1796
rect 2262 1791 2268 1792
rect 2674 1791 2680 1792
rect 2478 1780 2484 1781
rect 2718 1780 2724 1781
rect 2478 1776 2479 1780
rect 2483 1776 2719 1780
rect 2723 1776 2724 1780
rect 2478 1775 2484 1776
rect 2718 1775 2724 1776
rect 1846 1761 1847 1767
rect 1853 1766 3611 1767
rect 1853 1762 1863 1766
rect 1867 1762 1943 1766
rect 1947 1762 2007 1766
rect 2011 1762 2087 1766
rect 2091 1762 2231 1766
rect 2235 1762 2247 1766
rect 2251 1762 2415 1766
rect 2419 1762 2447 1766
rect 2451 1762 2599 1766
rect 2603 1762 2647 1766
rect 2651 1762 2791 1766
rect 2795 1762 2839 1766
rect 2843 1762 2991 1766
rect 2995 1762 3023 1766
rect 3027 1762 3199 1766
rect 3203 1762 3207 1766
rect 3211 1762 3399 1766
rect 3403 1762 3415 1766
rect 3419 1762 3575 1766
rect 3579 1762 3611 1766
rect 1853 1761 3611 1762
rect 3617 1761 3618 1767
rect 1846 1759 1854 1761
rect 96 1753 97 1759
rect 103 1758 1847 1759
rect 103 1754 111 1758
rect 115 1754 255 1758
rect 259 1754 327 1758
rect 331 1754 423 1758
rect 427 1754 471 1758
rect 475 1754 599 1758
rect 603 1754 615 1758
rect 619 1754 767 1758
rect 771 1754 919 1758
rect 923 1754 935 1758
rect 939 1754 1071 1758
rect 1075 1754 1087 1758
rect 1091 1754 1223 1758
rect 1227 1754 1231 1758
rect 1235 1754 1367 1758
rect 1371 1754 1375 1758
rect 1379 1754 1495 1758
rect 1499 1754 1527 1758
rect 1531 1754 1623 1758
rect 1627 1754 1687 1758
rect 1691 1754 1735 1758
rect 1739 1754 1823 1758
rect 1827 1754 1847 1758
rect 103 1753 1847 1754
rect 1853 1753 1854 1759
rect 1834 1689 1835 1695
rect 1841 1694 3599 1695
rect 1841 1690 1863 1694
rect 1867 1690 1911 1694
rect 1915 1690 1935 1694
rect 1939 1690 2031 1694
rect 2035 1690 2079 1694
rect 2083 1690 2151 1694
rect 2155 1690 2239 1694
rect 2243 1690 2271 1694
rect 2275 1690 2399 1694
rect 2403 1690 2407 1694
rect 2411 1690 2543 1694
rect 2547 1690 2591 1694
rect 2595 1690 2695 1694
rect 2699 1690 2783 1694
rect 2787 1690 2863 1694
rect 2867 1690 2983 1694
rect 2987 1690 3047 1694
rect 3051 1690 3191 1694
rect 3195 1690 3239 1694
rect 3243 1690 3407 1694
rect 3411 1690 3431 1694
rect 3435 1690 3575 1694
rect 3579 1690 3599 1694
rect 1841 1689 3599 1690
rect 3605 1689 3606 1695
rect 1834 1687 1842 1689
rect 84 1681 85 1687
rect 91 1686 1835 1687
rect 91 1682 111 1686
rect 115 1682 311 1686
rect 315 1682 319 1686
rect 323 1682 447 1686
rect 451 1682 463 1686
rect 467 1682 591 1686
rect 595 1682 607 1686
rect 611 1682 735 1686
rect 739 1682 759 1686
rect 763 1682 887 1686
rect 891 1682 911 1686
rect 915 1682 1039 1686
rect 1043 1682 1063 1686
rect 1067 1682 1191 1686
rect 1195 1682 1215 1686
rect 1219 1682 1343 1686
rect 1347 1682 1367 1686
rect 1371 1682 1495 1686
rect 1499 1682 1519 1686
rect 1523 1682 1647 1686
rect 1651 1682 1679 1686
rect 1683 1682 1823 1686
rect 1827 1682 1835 1686
rect 91 1681 1835 1682
rect 1841 1681 1842 1687
rect 1846 1613 1847 1619
rect 1853 1618 3611 1619
rect 1853 1614 1863 1618
rect 1867 1614 1895 1618
rect 1899 1614 1919 1618
rect 1923 1614 2015 1618
rect 2019 1614 2039 1618
rect 2043 1614 2151 1618
rect 2155 1614 2159 1618
rect 2163 1614 2279 1618
rect 2283 1614 2287 1618
rect 2291 1614 2407 1618
rect 2411 1614 2431 1618
rect 2435 1614 2551 1618
rect 2555 1614 2583 1618
rect 2587 1614 2703 1618
rect 2707 1614 2743 1618
rect 2747 1614 2871 1618
rect 2875 1614 2911 1618
rect 2915 1614 3055 1618
rect 3059 1614 3095 1618
rect 3099 1614 3247 1618
rect 3251 1614 3279 1618
rect 3283 1614 3439 1618
rect 3443 1614 3471 1618
rect 3475 1614 3575 1618
rect 3579 1614 3611 1618
rect 1853 1613 3611 1614
rect 3617 1613 3618 1619
rect 1846 1611 1854 1613
rect 96 1605 97 1611
rect 103 1610 1847 1611
rect 103 1606 111 1610
rect 115 1606 223 1610
rect 227 1606 319 1610
rect 323 1606 351 1610
rect 355 1606 455 1610
rect 459 1606 487 1610
rect 491 1606 599 1610
rect 603 1606 623 1610
rect 627 1606 743 1610
rect 747 1606 759 1610
rect 763 1606 895 1610
rect 899 1606 903 1610
rect 907 1606 1047 1610
rect 1051 1606 1055 1610
rect 1059 1606 1199 1610
rect 1203 1606 1215 1610
rect 1219 1606 1351 1610
rect 1355 1606 1375 1610
rect 1379 1606 1503 1610
rect 1507 1606 1543 1610
rect 1547 1606 1655 1610
rect 1659 1606 1823 1610
rect 1827 1606 1847 1610
rect 103 1605 1847 1606
rect 1853 1605 1854 1611
rect 1834 1542 3606 1543
rect 1834 1539 1863 1542
rect 84 1533 85 1539
rect 91 1538 1835 1539
rect 91 1534 111 1538
rect 115 1534 135 1538
rect 139 1534 215 1538
rect 219 1534 271 1538
rect 275 1534 343 1538
rect 347 1534 423 1538
rect 427 1534 479 1538
rect 483 1534 583 1538
rect 587 1534 615 1538
rect 619 1534 735 1538
rect 739 1534 751 1538
rect 755 1534 887 1538
rect 891 1534 895 1538
rect 899 1534 1039 1538
rect 1043 1534 1047 1538
rect 1051 1534 1191 1538
rect 1195 1534 1207 1538
rect 1211 1534 1343 1538
rect 1347 1534 1367 1538
rect 1371 1534 1495 1538
rect 1499 1534 1535 1538
rect 1539 1534 1823 1538
rect 1827 1534 1835 1538
rect 91 1533 1835 1534
rect 1841 1538 1863 1539
rect 1867 1538 1887 1542
rect 1891 1538 2007 1542
rect 2011 1538 2023 1542
rect 2027 1538 2143 1542
rect 2147 1538 2183 1542
rect 2187 1538 2279 1542
rect 2283 1538 2343 1542
rect 2347 1538 2423 1542
rect 2427 1538 2503 1542
rect 2507 1538 2575 1542
rect 2579 1538 2663 1542
rect 2667 1538 2735 1542
rect 2739 1538 2823 1542
rect 2827 1538 2903 1542
rect 2907 1538 2983 1542
rect 2987 1538 3087 1542
rect 3091 1538 3151 1542
rect 3155 1538 3271 1542
rect 3275 1538 3319 1542
rect 3323 1538 3463 1542
rect 3467 1538 3479 1542
rect 3483 1538 3575 1542
rect 3579 1538 3606 1542
rect 1841 1537 3606 1538
rect 1841 1533 1842 1537
rect 2702 1532 2708 1533
rect 3018 1532 3024 1533
rect 2702 1528 2703 1532
rect 2707 1528 3019 1532
rect 3023 1528 3024 1532
rect 2702 1527 2708 1528
rect 3018 1527 3024 1528
rect 2718 1484 2724 1485
rect 3078 1484 3084 1485
rect 2718 1480 2719 1484
rect 2723 1480 3079 1484
rect 3083 1480 3084 1484
rect 2718 1479 2724 1480
rect 3078 1479 3084 1480
rect 1846 1466 3618 1467
rect 1846 1463 1863 1466
rect 96 1457 97 1463
rect 103 1462 1847 1463
rect 103 1458 111 1462
rect 115 1458 143 1462
rect 147 1458 263 1462
rect 267 1458 279 1462
rect 283 1458 399 1462
rect 403 1458 431 1462
rect 435 1458 535 1462
rect 539 1458 591 1462
rect 595 1458 663 1462
rect 667 1458 743 1462
rect 747 1458 791 1462
rect 795 1458 895 1462
rect 899 1458 911 1462
rect 915 1458 1023 1462
rect 1027 1458 1047 1462
rect 1051 1458 1143 1462
rect 1147 1458 1199 1462
rect 1203 1458 1263 1462
rect 1267 1458 1351 1462
rect 1355 1458 1383 1462
rect 1387 1458 1503 1462
rect 1507 1458 1631 1462
rect 1635 1458 1735 1462
rect 1739 1458 1823 1462
rect 1827 1458 1847 1462
rect 103 1457 1847 1458
rect 1853 1462 1863 1463
rect 1867 1462 1895 1466
rect 1899 1462 2031 1466
rect 2035 1462 2183 1466
rect 2187 1462 2191 1466
rect 2195 1462 2351 1466
rect 2355 1462 2359 1466
rect 2363 1462 2511 1466
rect 2515 1462 2527 1466
rect 2531 1462 2671 1466
rect 2675 1462 2687 1466
rect 2691 1462 2831 1466
rect 2835 1462 2847 1466
rect 2851 1462 2991 1466
rect 2995 1462 3007 1466
rect 3011 1462 3159 1466
rect 3163 1462 3175 1466
rect 3179 1462 3327 1466
rect 3331 1462 3343 1466
rect 3347 1462 3487 1466
rect 3491 1462 3575 1466
rect 3579 1462 3618 1466
rect 1853 1461 3618 1462
rect 1853 1457 1854 1461
rect 2222 1436 2228 1437
rect 2426 1436 2432 1437
rect 2222 1432 2223 1436
rect 2227 1432 2427 1436
rect 2431 1432 2432 1436
rect 2222 1431 2228 1432
rect 2426 1431 2432 1432
rect 84 1389 85 1395
rect 91 1394 1835 1395
rect 91 1390 111 1394
rect 115 1390 135 1394
rect 139 1390 255 1394
rect 259 1390 327 1394
rect 331 1390 391 1394
rect 395 1390 527 1394
rect 531 1390 551 1394
rect 555 1390 655 1394
rect 659 1390 783 1394
rect 787 1390 903 1394
rect 907 1390 1015 1394
rect 1019 1390 1023 1394
rect 1027 1390 1135 1394
rect 1139 1390 1255 1394
rect 1259 1390 1263 1394
rect 1267 1390 1375 1394
rect 1379 1390 1495 1394
rect 1499 1390 1503 1394
rect 1507 1390 1623 1394
rect 1627 1390 1727 1394
rect 1731 1390 1823 1394
rect 1827 1390 1835 1394
rect 91 1389 1835 1390
rect 1841 1391 1842 1395
rect 1841 1390 3606 1391
rect 1841 1389 1863 1390
rect 1834 1386 1863 1389
rect 1867 1386 2079 1390
rect 2083 1386 2175 1390
rect 2179 1386 2263 1390
rect 2267 1386 2351 1390
rect 2355 1386 2439 1390
rect 2443 1386 2519 1390
rect 2523 1386 2615 1390
rect 2619 1386 2679 1390
rect 2683 1386 2783 1390
rect 2787 1386 2839 1390
rect 2843 1386 2935 1390
rect 2939 1386 2999 1390
rect 3003 1386 3079 1390
rect 3083 1386 3167 1390
rect 3171 1386 3223 1390
rect 3227 1386 3335 1390
rect 3339 1386 3359 1390
rect 3363 1386 3479 1390
rect 3483 1386 3575 1390
rect 3579 1386 3606 1390
rect 1834 1385 3606 1386
rect 1302 1340 1308 1341
rect 1638 1340 1644 1341
rect 1302 1336 1303 1340
rect 1307 1336 1639 1340
rect 1643 1336 1644 1340
rect 1302 1335 1308 1336
rect 1638 1335 1644 1336
rect 2822 1340 2828 1341
rect 3258 1340 3264 1341
rect 2822 1336 2823 1340
rect 2827 1336 3259 1340
rect 3263 1336 3264 1340
rect 2822 1335 2828 1336
rect 3258 1335 3264 1336
rect 2118 1332 2124 1333
rect 2538 1332 2544 1333
rect 2118 1328 2119 1332
rect 2123 1328 2539 1332
rect 2543 1328 2544 1332
rect 2118 1327 2124 1328
rect 2538 1327 2544 1328
rect 1846 1322 3618 1323
rect 1846 1319 1863 1322
rect 96 1313 97 1319
rect 103 1318 1847 1319
rect 103 1314 111 1318
rect 115 1314 143 1318
rect 147 1314 327 1318
rect 331 1314 335 1318
rect 339 1314 527 1318
rect 531 1314 559 1318
rect 563 1314 719 1318
rect 723 1314 791 1318
rect 795 1314 903 1318
rect 907 1314 1031 1318
rect 1035 1314 1071 1318
rect 1075 1314 1231 1318
rect 1235 1314 1271 1318
rect 1275 1314 1383 1318
rect 1387 1314 1511 1318
rect 1515 1314 1535 1318
rect 1539 1314 1687 1318
rect 1691 1314 1735 1318
rect 1739 1314 1823 1318
rect 1827 1314 1847 1318
rect 103 1313 1847 1314
rect 1853 1318 1863 1319
rect 1867 1318 2087 1322
rect 2091 1318 2271 1322
rect 2275 1318 2311 1322
rect 2315 1318 2447 1322
rect 2451 1318 2519 1322
rect 2523 1318 2623 1322
rect 2627 1318 2711 1322
rect 2715 1318 2791 1322
rect 2795 1318 2887 1322
rect 2891 1318 2943 1322
rect 2947 1318 3047 1322
rect 3051 1318 3087 1322
rect 3091 1318 3199 1322
rect 3203 1318 3231 1322
rect 3235 1318 3351 1322
rect 3355 1318 3367 1322
rect 3371 1318 3487 1322
rect 3491 1318 3575 1322
rect 3579 1318 3618 1322
rect 1853 1317 3618 1318
rect 1853 1313 1854 1317
rect 2294 1292 2300 1293
rect 2442 1292 2448 1293
rect 2294 1288 2295 1292
rect 2299 1288 2443 1292
rect 2447 1288 2448 1292
rect 2294 1287 2300 1288
rect 2442 1287 2448 1288
rect 1834 1250 3606 1251
rect 1834 1247 1863 1250
rect 84 1241 85 1247
rect 91 1246 1835 1247
rect 91 1242 111 1246
rect 115 1242 135 1246
rect 139 1242 295 1246
rect 299 1242 319 1246
rect 323 1242 479 1246
rect 483 1242 519 1246
rect 523 1242 655 1246
rect 659 1242 711 1246
rect 715 1242 815 1246
rect 819 1242 895 1246
rect 899 1242 967 1246
rect 971 1242 1063 1246
rect 1067 1242 1111 1246
rect 1115 1242 1223 1246
rect 1227 1242 1247 1246
rect 1251 1242 1375 1246
rect 1379 1242 1383 1246
rect 1387 1242 1527 1246
rect 1531 1242 1679 1246
rect 1683 1242 1823 1246
rect 1827 1242 1835 1246
rect 91 1241 1835 1242
rect 1841 1246 1863 1247
rect 1867 1246 1903 1250
rect 1907 1246 1991 1250
rect 1995 1246 2079 1250
rect 2083 1246 2095 1250
rect 2099 1246 2215 1250
rect 2219 1246 2303 1250
rect 2307 1246 2351 1250
rect 2355 1246 2487 1250
rect 2491 1246 2511 1250
rect 2515 1246 2631 1250
rect 2635 1246 2703 1250
rect 2707 1246 2775 1250
rect 2779 1246 2879 1250
rect 2883 1246 2919 1250
rect 2923 1246 3039 1250
rect 3043 1246 3063 1250
rect 3067 1246 3191 1250
rect 3195 1246 3207 1250
rect 3211 1246 3343 1250
rect 3347 1246 3351 1250
rect 3355 1246 3479 1250
rect 3483 1246 3575 1250
rect 3579 1246 3606 1250
rect 1841 1245 3606 1246
rect 1841 1241 1842 1245
rect 2814 1196 2820 1197
rect 3138 1196 3144 1197
rect 2814 1192 2815 1196
rect 2819 1192 3139 1196
rect 3143 1192 3144 1196
rect 2814 1191 2820 1192
rect 3138 1191 3144 1192
rect 1846 1178 3618 1179
rect 1846 1175 1863 1178
rect 96 1169 97 1175
rect 103 1174 1847 1175
rect 103 1170 111 1174
rect 115 1170 143 1174
rect 147 1170 167 1174
rect 171 1170 303 1174
rect 307 1170 319 1174
rect 323 1170 471 1174
rect 475 1170 487 1174
rect 491 1170 615 1174
rect 619 1170 663 1174
rect 667 1170 759 1174
rect 763 1170 823 1174
rect 827 1170 911 1174
rect 915 1170 975 1174
rect 979 1170 1063 1174
rect 1067 1170 1119 1174
rect 1123 1170 1231 1174
rect 1235 1170 1255 1174
rect 1259 1170 1391 1174
rect 1395 1170 1399 1174
rect 1403 1170 1535 1174
rect 1539 1170 1575 1174
rect 1579 1170 1735 1174
rect 1739 1170 1823 1174
rect 1827 1170 1847 1174
rect 103 1169 1847 1170
rect 1853 1174 1863 1175
rect 1867 1174 1895 1178
rect 1899 1174 1911 1178
rect 1915 1174 1999 1178
rect 2003 1174 2063 1178
rect 2067 1174 2103 1178
rect 2107 1174 2223 1178
rect 2227 1174 2255 1178
rect 2259 1174 2359 1178
rect 2363 1174 2439 1178
rect 2443 1174 2495 1178
rect 2499 1174 2615 1178
rect 2619 1174 2639 1178
rect 2643 1174 2783 1178
rect 2787 1174 2791 1178
rect 2795 1174 2927 1178
rect 2931 1174 2967 1178
rect 2971 1174 3071 1178
rect 3075 1174 3143 1178
rect 3147 1174 3215 1178
rect 3219 1174 3327 1178
rect 3331 1174 3359 1178
rect 3363 1174 3487 1178
rect 3491 1174 3575 1178
rect 3579 1174 3618 1178
rect 1853 1173 3618 1174
rect 1853 1169 1854 1173
rect 1050 1164 1056 1165
rect 1538 1164 1544 1165
rect 1050 1160 1051 1164
rect 1055 1160 1539 1164
rect 1543 1160 1544 1164
rect 1050 1159 1056 1160
rect 1538 1159 1544 1160
rect 84 1097 85 1103
rect 91 1102 1835 1103
rect 91 1098 111 1102
rect 115 1098 159 1102
rect 163 1098 215 1102
rect 219 1098 311 1102
rect 315 1098 327 1102
rect 331 1098 439 1102
rect 443 1098 463 1102
rect 467 1098 559 1102
rect 563 1098 607 1102
rect 611 1098 679 1102
rect 683 1098 751 1102
rect 755 1098 807 1102
rect 811 1098 903 1102
rect 907 1098 943 1102
rect 947 1098 1055 1102
rect 1059 1098 1087 1102
rect 1091 1098 1223 1102
rect 1227 1098 1247 1102
rect 1251 1098 1391 1102
rect 1395 1098 1407 1102
rect 1411 1098 1567 1102
rect 1571 1098 1575 1102
rect 1579 1098 1727 1102
rect 1731 1098 1823 1102
rect 1827 1098 1835 1102
rect 91 1097 1835 1098
rect 1841 1099 1842 1103
rect 1841 1098 3606 1099
rect 1841 1097 1863 1098
rect 1834 1094 1863 1097
rect 1867 1094 1887 1098
rect 1891 1094 1935 1098
rect 1939 1094 2055 1098
rect 2059 1094 2095 1098
rect 2099 1094 2247 1098
rect 2251 1094 2407 1098
rect 2411 1094 2431 1098
rect 2435 1094 2567 1098
rect 2571 1094 2607 1098
rect 2611 1094 2735 1098
rect 2739 1094 2783 1098
rect 2787 1094 2911 1098
rect 2915 1094 2959 1098
rect 2963 1094 3095 1098
rect 3099 1094 3135 1098
rect 3139 1094 3287 1098
rect 3291 1094 3319 1098
rect 3323 1094 3479 1098
rect 3483 1094 3575 1098
rect 3579 1094 3606 1098
rect 1834 1093 3606 1094
rect 998 1084 1004 1085
rect 1338 1084 1344 1085
rect 998 1080 999 1084
rect 1003 1080 1339 1084
rect 1343 1080 1344 1084
rect 998 1079 1004 1080
rect 1338 1079 1344 1080
rect 96 1021 97 1027
rect 103 1026 1847 1027
rect 103 1022 111 1026
rect 115 1022 223 1026
rect 227 1022 335 1026
rect 339 1022 343 1026
rect 347 1022 431 1026
rect 435 1022 447 1026
rect 451 1022 535 1026
rect 539 1022 567 1026
rect 571 1022 655 1026
rect 659 1022 687 1026
rect 691 1022 791 1026
rect 795 1022 815 1026
rect 819 1022 951 1026
rect 955 1022 1095 1026
rect 1099 1022 1135 1026
rect 1139 1022 1255 1026
rect 1259 1022 1327 1026
rect 1331 1022 1415 1026
rect 1419 1022 1535 1026
rect 1539 1022 1583 1026
rect 1587 1022 1735 1026
rect 1739 1022 1823 1026
rect 1827 1022 1847 1026
rect 103 1021 1847 1022
rect 1853 1026 3618 1027
rect 1853 1022 1863 1026
rect 1867 1022 1943 1026
rect 1947 1022 2071 1026
rect 2075 1022 2103 1026
rect 2107 1022 2191 1026
rect 2195 1022 2255 1026
rect 2259 1022 2311 1026
rect 2315 1022 2415 1026
rect 2419 1022 2439 1026
rect 2443 1022 2575 1026
rect 2579 1022 2719 1026
rect 2723 1022 2743 1026
rect 2747 1022 2871 1026
rect 2875 1022 2919 1026
rect 2923 1022 3031 1026
rect 3035 1022 3103 1026
rect 3107 1022 3191 1026
rect 3195 1022 3295 1026
rect 3299 1022 3351 1026
rect 3355 1022 3487 1026
rect 3491 1022 3575 1026
rect 3579 1022 3618 1026
rect 1853 1021 3618 1022
rect 84 949 85 955
rect 91 954 1835 955
rect 91 950 111 954
rect 115 950 335 954
rect 339 950 367 954
rect 371 950 423 954
rect 427 950 463 954
rect 467 950 527 954
rect 531 950 575 954
rect 579 950 647 954
rect 651 950 703 954
rect 707 950 783 954
rect 787 950 847 954
rect 851 950 943 954
rect 947 950 1007 954
rect 1011 950 1127 954
rect 1131 950 1175 954
rect 1179 950 1319 954
rect 1323 950 1351 954
rect 1355 950 1527 954
rect 1531 950 1711 954
rect 1715 950 1727 954
rect 1731 950 1823 954
rect 1827 950 1835 954
rect 91 949 1835 950
rect 1841 954 3606 955
rect 1841 950 1863 954
rect 1867 950 1887 954
rect 1891 950 1935 954
rect 1939 950 2047 954
rect 2051 950 2063 954
rect 2067 950 2183 954
rect 2187 950 2199 954
rect 2203 950 2303 954
rect 2307 950 2351 954
rect 2355 950 2431 954
rect 2435 950 2495 954
rect 2499 950 2567 954
rect 2571 950 2631 954
rect 2635 950 2711 954
rect 2715 950 2759 954
rect 2763 950 2863 954
rect 2867 950 2887 954
rect 2891 950 3023 954
rect 3027 950 3183 954
rect 3187 950 3343 954
rect 3347 950 3479 954
rect 3483 950 3575 954
rect 3579 950 3606 954
rect 1841 949 3606 950
rect 1390 900 1396 901
rect 1666 900 1672 901
rect 1390 896 1391 900
rect 1395 896 1667 900
rect 1671 896 1672 900
rect 1390 895 1396 896
rect 1666 895 1672 896
rect 1846 886 3618 887
rect 1846 883 1863 886
rect 96 877 97 883
rect 103 882 1847 883
rect 103 878 111 882
rect 115 878 343 882
rect 347 878 375 882
rect 379 878 431 882
rect 435 878 471 882
rect 475 878 535 882
rect 539 878 583 882
rect 587 878 647 882
rect 651 878 711 882
rect 715 878 783 882
rect 787 878 855 882
rect 859 878 927 882
rect 931 878 1015 882
rect 1019 878 1087 882
rect 1091 878 1183 882
rect 1187 878 1263 882
rect 1267 878 1359 882
rect 1363 878 1447 882
rect 1451 878 1535 882
rect 1539 878 1631 882
rect 1635 878 1719 882
rect 1723 878 1823 882
rect 1827 878 1847 882
rect 103 877 1847 878
rect 1853 882 1863 883
rect 1867 882 1895 886
rect 1899 882 2015 886
rect 2019 882 2055 886
rect 2059 882 2167 886
rect 2171 882 2207 886
rect 2211 882 2319 886
rect 2323 882 2359 886
rect 2363 882 2487 886
rect 2491 882 2503 886
rect 2507 882 2639 886
rect 2643 882 2663 886
rect 2667 882 2767 886
rect 2771 882 2847 886
rect 2851 882 2895 886
rect 2899 882 3031 886
rect 3035 882 3039 886
rect 3043 882 3239 886
rect 3243 882 3439 886
rect 3443 882 3575 886
rect 3579 882 3618 886
rect 1853 881 3618 882
rect 1853 877 1854 881
rect 1834 818 3606 819
rect 1834 815 1863 818
rect 84 809 85 815
rect 91 814 1835 815
rect 91 810 111 814
rect 115 810 287 814
rect 291 810 335 814
rect 339 810 407 814
rect 411 810 423 814
rect 427 810 527 814
rect 531 810 535 814
rect 539 810 639 814
rect 643 810 679 814
rect 683 810 775 814
rect 779 810 823 814
rect 827 810 919 814
rect 923 810 975 814
rect 979 810 1079 814
rect 1083 810 1127 814
rect 1131 810 1255 814
rect 1259 810 1279 814
rect 1283 810 1439 814
rect 1443 810 1599 814
rect 1603 810 1623 814
rect 1627 810 1823 814
rect 1827 810 1835 814
rect 91 809 1835 810
rect 1841 814 1863 815
rect 1867 814 1887 818
rect 1891 814 1991 818
rect 1995 814 2007 818
rect 2011 814 2135 818
rect 2139 814 2159 818
rect 2163 814 2287 818
rect 2291 814 2311 818
rect 2315 814 2455 818
rect 2459 814 2479 818
rect 2483 814 2623 818
rect 2627 814 2655 818
rect 2659 814 2799 818
rect 2803 814 2839 818
rect 2843 814 2967 818
rect 2971 814 3031 818
rect 3035 814 3143 818
rect 3147 814 3231 818
rect 3235 814 3319 818
rect 3323 814 3431 818
rect 3435 814 3479 818
rect 3483 814 3575 818
rect 3579 814 3606 818
rect 1841 813 3606 814
rect 1841 809 1842 813
rect 1314 756 1320 757
rect 1518 756 1524 757
rect 1314 752 1315 756
rect 1319 752 1519 756
rect 1523 752 1524 756
rect 1314 751 1320 752
rect 1518 751 1524 752
rect 1846 746 3618 747
rect 1846 743 1863 746
rect 96 737 97 743
rect 103 742 1847 743
rect 103 738 111 742
rect 115 738 215 742
rect 219 738 295 742
rect 299 738 359 742
rect 363 738 415 742
rect 419 738 503 742
rect 507 738 543 742
rect 547 738 647 742
rect 651 738 687 742
rect 691 738 791 742
rect 795 738 831 742
rect 835 738 935 742
rect 939 738 983 742
rect 987 738 1087 742
rect 1091 738 1135 742
rect 1139 738 1247 742
rect 1251 738 1287 742
rect 1291 738 1415 742
rect 1419 738 1447 742
rect 1451 738 1583 742
rect 1587 738 1607 742
rect 1611 738 1735 742
rect 1739 738 1823 742
rect 1827 738 1847 742
rect 103 737 1847 738
rect 1853 742 1863 743
rect 1867 742 1895 746
rect 1899 742 1999 746
rect 2003 742 2063 746
rect 2067 742 2143 746
rect 2147 742 2255 746
rect 2259 742 2295 746
rect 2299 742 2447 746
rect 2451 742 2463 746
rect 2467 742 2631 746
rect 2635 742 2639 746
rect 2643 742 2807 746
rect 2811 742 2823 746
rect 2827 742 2975 746
rect 2979 742 2999 746
rect 3003 742 3151 746
rect 3155 742 3167 746
rect 3171 742 3327 746
rect 3331 742 3335 746
rect 3339 742 3487 746
rect 3491 742 3575 746
rect 3579 742 3618 746
rect 1853 741 3618 742
rect 1853 737 1854 741
rect 84 669 85 675
rect 91 674 1835 675
rect 91 670 111 674
rect 115 670 135 674
rect 139 670 207 674
rect 211 670 295 674
rect 299 670 351 674
rect 355 670 463 674
rect 467 670 495 674
rect 499 670 623 674
rect 627 670 639 674
rect 643 670 775 674
rect 779 670 783 674
rect 787 670 927 674
rect 931 670 1071 674
rect 1075 670 1079 674
rect 1083 670 1207 674
rect 1211 670 1239 674
rect 1243 670 1343 674
rect 1347 670 1407 674
rect 1411 670 1479 674
rect 1483 670 1575 674
rect 1579 670 1615 674
rect 1619 670 1727 674
rect 1731 670 1823 674
rect 1827 670 1835 674
rect 91 669 1835 670
rect 1841 674 3606 675
rect 1841 670 1863 674
rect 1867 670 1887 674
rect 1891 670 2055 674
rect 2059 670 2215 674
rect 2219 670 2247 674
rect 2251 670 2359 674
rect 2363 670 2439 674
rect 2443 670 2511 674
rect 2515 670 2631 674
rect 2635 670 2671 674
rect 2675 670 2815 674
rect 2819 670 2831 674
rect 2835 670 2991 674
rect 2995 670 3159 674
rect 3163 670 3327 674
rect 3331 670 3479 674
rect 3483 670 3575 674
rect 3579 670 3606 674
rect 1841 669 3606 670
rect 96 597 97 603
rect 103 602 1847 603
rect 103 598 111 602
rect 115 598 143 602
rect 147 598 303 602
rect 307 598 471 602
rect 475 598 487 602
rect 491 598 631 602
rect 635 598 671 602
rect 675 598 783 602
rect 787 598 847 602
rect 851 598 935 602
rect 939 598 1023 602
rect 1027 598 1079 602
rect 1083 598 1199 602
rect 1203 598 1215 602
rect 1219 598 1351 602
rect 1355 598 1375 602
rect 1379 598 1487 602
rect 1491 598 1559 602
rect 1563 598 1623 602
rect 1627 598 1735 602
rect 1739 598 1823 602
rect 1827 598 1847 602
rect 103 597 1847 598
rect 1853 602 3618 603
rect 1853 598 1863 602
rect 1867 598 2199 602
rect 2203 598 2223 602
rect 2227 598 2287 602
rect 2291 598 2367 602
rect 2371 598 2375 602
rect 2379 598 2463 602
rect 2467 598 2519 602
rect 2523 598 2567 602
rect 2571 598 2679 602
rect 2683 598 2815 602
rect 2819 598 2839 602
rect 2843 598 2975 602
rect 2979 598 2999 602
rect 3003 598 3143 602
rect 3147 598 3167 602
rect 3171 598 3327 602
rect 3331 598 3335 602
rect 3339 598 3487 602
rect 3491 598 3575 602
rect 3579 598 3618 602
rect 1853 597 3618 598
rect 84 525 85 531
rect 91 530 1835 531
rect 91 526 111 530
rect 115 526 135 530
rect 139 526 295 530
rect 299 526 303 530
rect 307 526 479 530
rect 483 526 495 530
rect 499 526 663 530
rect 667 526 679 530
rect 683 526 839 530
rect 843 526 863 530
rect 867 526 1015 530
rect 1019 526 1031 530
rect 1035 526 1191 530
rect 1195 526 1351 530
rect 1355 526 1367 530
rect 1371 526 1503 530
rect 1507 526 1551 530
rect 1555 526 1663 530
rect 1667 526 1727 530
rect 1731 526 1823 530
rect 1827 526 1835 530
rect 91 525 1835 526
rect 1841 530 3606 531
rect 1841 526 1863 530
rect 1867 526 2191 530
rect 2195 526 2279 530
rect 2283 526 2303 530
rect 2307 526 2367 530
rect 2371 526 2399 530
rect 2403 526 2455 530
rect 2459 526 2503 530
rect 2507 526 2559 530
rect 2563 526 2607 530
rect 2611 526 2671 530
rect 2675 526 2719 530
rect 2723 526 2807 530
rect 2811 526 2839 530
rect 2843 526 2967 530
rect 2971 526 3095 530
rect 3099 526 3135 530
rect 3139 526 3223 530
rect 3227 526 3319 530
rect 3323 526 3351 530
rect 3355 526 3479 530
rect 3483 526 3575 530
rect 3579 526 3606 530
rect 1841 525 3606 526
rect 3006 476 3012 477
rect 3290 476 3296 477
rect 3006 472 3007 476
rect 3011 472 3291 476
rect 3295 472 3296 476
rect 3006 471 3012 472
rect 3290 471 3296 472
rect 1846 462 3618 463
rect 1846 459 1863 462
rect 96 453 97 459
rect 103 458 1847 459
rect 103 454 111 458
rect 115 454 143 458
rect 147 454 303 458
rect 307 454 311 458
rect 315 454 495 458
rect 499 454 503 458
rect 507 454 687 458
rect 691 454 871 458
rect 875 454 879 458
rect 883 454 1039 458
rect 1043 454 1055 458
rect 1059 454 1199 458
rect 1203 454 1223 458
rect 1227 454 1359 458
rect 1363 454 1391 458
rect 1395 454 1511 458
rect 1515 454 1559 458
rect 1563 454 1671 458
rect 1675 454 1727 458
rect 1731 454 1823 458
rect 1827 454 1847 458
rect 103 453 1847 454
rect 1853 458 1863 459
rect 1867 458 2239 462
rect 2243 458 2311 462
rect 2315 458 2327 462
rect 2331 458 2407 462
rect 2411 458 2431 462
rect 2435 458 2511 462
rect 2515 458 2559 462
rect 2563 458 2615 462
rect 2619 458 2695 462
rect 2699 458 2727 462
rect 2731 458 2847 462
rect 2851 458 2975 462
rect 2979 458 2999 462
rect 3003 458 3103 462
rect 3107 458 3159 462
rect 3163 458 3231 462
rect 3235 458 3327 462
rect 3331 458 3359 462
rect 3363 458 3487 462
rect 3491 458 3575 462
rect 3579 458 3618 462
rect 1853 457 3618 458
rect 1853 453 1854 457
rect 1834 394 3606 395
rect 1834 391 1863 394
rect 84 385 85 391
rect 91 390 1835 391
rect 91 386 111 390
rect 115 386 135 390
rect 139 386 263 390
rect 267 386 295 390
rect 299 386 423 390
rect 427 386 487 390
rect 491 386 591 390
rect 595 386 679 390
rect 683 386 767 390
rect 771 386 871 390
rect 875 386 935 390
rect 939 386 1047 390
rect 1051 386 1103 390
rect 1107 386 1215 390
rect 1219 386 1263 390
rect 1267 386 1383 390
rect 1387 386 1423 390
rect 1427 386 1551 390
rect 1555 386 1583 390
rect 1587 386 1719 390
rect 1723 386 1727 390
rect 1731 386 1823 390
rect 1827 386 1835 390
rect 91 385 1835 386
rect 1841 390 1863 391
rect 1867 390 2183 394
rect 2187 390 2231 394
rect 2235 390 2287 394
rect 2291 390 2319 394
rect 2323 390 2399 394
rect 2403 390 2423 394
rect 2427 390 2527 394
rect 2531 390 2551 394
rect 2555 390 2671 394
rect 2675 390 2687 394
rect 2691 390 2815 394
rect 2819 390 2839 394
rect 2843 390 2967 394
rect 2971 390 2991 394
rect 2995 390 3127 394
rect 3131 390 3151 394
rect 3155 390 3295 394
rect 3299 390 3319 394
rect 3323 390 3463 394
rect 3467 390 3479 394
rect 3483 390 3575 394
rect 3579 390 3606 394
rect 1841 389 3606 390
rect 1841 385 1842 389
rect 96 317 97 323
rect 103 322 1847 323
rect 103 318 111 322
rect 115 318 143 322
rect 147 318 215 322
rect 219 318 271 322
rect 275 318 351 322
rect 355 318 431 322
rect 435 318 495 322
rect 499 318 599 322
rect 603 318 639 322
rect 643 318 775 322
rect 779 318 791 322
rect 795 318 935 322
rect 939 318 943 322
rect 947 318 1079 322
rect 1083 318 1111 322
rect 1115 318 1223 322
rect 1227 318 1271 322
rect 1275 318 1359 322
rect 1363 318 1431 322
rect 1435 318 1487 322
rect 1491 318 1591 322
rect 1595 318 1623 322
rect 1627 318 1735 322
rect 1739 318 1823 322
rect 1827 318 1847 322
rect 103 317 1847 318
rect 1853 319 1854 323
rect 1853 318 3618 319
rect 1853 317 1863 318
rect 1846 314 1863 317
rect 1867 314 1895 318
rect 1899 314 2087 318
rect 2091 314 2191 318
rect 2195 314 2295 318
rect 2299 314 2303 318
rect 2307 314 2407 318
rect 2411 314 2511 318
rect 2515 314 2535 318
rect 2539 314 2679 318
rect 2683 314 2711 318
rect 2715 314 2823 318
rect 2827 314 2903 318
rect 2907 314 2975 318
rect 2979 314 3095 318
rect 3099 314 3135 318
rect 3139 314 3295 318
rect 3299 314 3303 318
rect 3307 314 3471 318
rect 3475 314 3487 318
rect 3491 314 3575 318
rect 3579 314 3618 318
rect 1846 313 3618 314
rect 1834 250 3606 251
rect 1834 247 1863 250
rect 84 241 85 247
rect 91 246 1835 247
rect 91 242 111 246
rect 115 242 207 246
rect 211 242 231 246
rect 235 242 343 246
rect 347 242 359 246
rect 363 242 487 246
rect 491 242 623 246
rect 627 242 631 246
rect 635 242 759 246
rect 763 242 783 246
rect 787 242 895 246
rect 899 242 927 246
rect 931 242 1031 246
rect 1035 242 1071 246
rect 1075 242 1159 246
rect 1163 242 1215 246
rect 1219 242 1295 246
rect 1299 242 1351 246
rect 1355 242 1431 246
rect 1435 242 1479 246
rect 1483 242 1615 246
rect 1619 242 1727 246
rect 1731 242 1823 246
rect 1827 242 1835 246
rect 91 241 1835 242
rect 1841 246 1863 247
rect 1867 246 1887 250
rect 1891 246 1999 250
rect 2003 246 2079 250
rect 2083 246 2143 250
rect 2147 246 2295 250
rect 2299 246 2455 250
rect 2459 246 2503 250
rect 2507 246 2615 250
rect 2619 246 2703 250
rect 2707 246 2783 250
rect 2787 246 2895 250
rect 2899 246 2951 250
rect 2955 246 3087 250
rect 3091 246 3127 250
rect 3131 246 3287 250
rect 3291 246 3311 250
rect 3315 246 3479 250
rect 3483 246 3575 250
rect 3579 246 3606 250
rect 1841 245 3606 246
rect 1841 241 1842 245
rect 96 149 97 155
rect 103 154 1847 155
rect 103 150 111 154
rect 115 150 175 154
rect 179 150 239 154
rect 243 150 263 154
rect 267 150 351 154
rect 355 150 367 154
rect 371 150 439 154
rect 443 150 495 154
rect 499 150 527 154
rect 531 150 615 154
rect 619 150 631 154
rect 635 150 703 154
rect 707 150 767 154
rect 771 150 791 154
rect 795 150 879 154
rect 883 150 903 154
rect 907 150 967 154
rect 971 150 1039 154
rect 1043 150 1055 154
rect 1059 150 1143 154
rect 1147 150 1167 154
rect 1171 150 1231 154
rect 1235 150 1303 154
rect 1307 150 1319 154
rect 1323 150 1407 154
rect 1411 150 1439 154
rect 1443 150 1503 154
rect 1507 150 1823 154
rect 1827 150 1847 154
rect 103 149 1847 150
rect 1853 154 3618 155
rect 1853 150 1863 154
rect 1867 150 1895 154
rect 1899 150 1983 154
rect 1987 150 2007 154
rect 2011 150 2071 154
rect 2075 150 2151 154
rect 2155 150 2159 154
rect 2163 150 2247 154
rect 2251 150 2303 154
rect 2307 150 2335 154
rect 2339 150 2439 154
rect 2443 150 2463 154
rect 2467 150 2543 154
rect 2547 150 2623 154
rect 2627 150 2647 154
rect 2651 150 2743 154
rect 2747 150 2791 154
rect 2795 150 2839 154
rect 2843 150 2935 154
rect 2939 150 2959 154
rect 2963 150 3031 154
rect 3035 150 3127 154
rect 3131 150 3135 154
rect 3139 150 3223 154
rect 3227 150 3311 154
rect 3315 150 3319 154
rect 3323 150 3399 154
rect 3403 150 3487 154
rect 3491 150 3575 154
rect 3579 150 3618 154
rect 1853 149 3618 150
rect 84 81 85 87
rect 91 86 1835 87
rect 91 82 111 86
rect 115 82 167 86
rect 171 82 255 86
rect 259 82 343 86
rect 347 82 431 86
rect 435 82 519 86
rect 523 82 607 86
rect 611 82 695 86
rect 699 82 783 86
rect 787 82 871 86
rect 875 82 959 86
rect 963 82 1047 86
rect 1051 82 1135 86
rect 1139 82 1223 86
rect 1227 82 1311 86
rect 1315 82 1399 86
rect 1403 82 1495 86
rect 1499 82 1823 86
rect 1827 82 1835 86
rect 91 81 1835 82
rect 1841 86 3606 87
rect 1841 82 1863 86
rect 1867 82 1887 86
rect 1891 82 1975 86
rect 1979 82 2063 86
rect 2067 82 2151 86
rect 2155 82 2239 86
rect 2243 82 2327 86
rect 2331 82 2431 86
rect 2435 82 2535 86
rect 2539 82 2639 86
rect 2643 82 2735 86
rect 2739 82 2831 86
rect 2835 82 2927 86
rect 2931 82 3023 86
rect 3027 82 3119 86
rect 3123 82 3215 86
rect 3219 82 3303 86
rect 3307 82 3391 86
rect 3395 82 3479 86
rect 3483 82 3575 86
rect 3579 82 3606 86
rect 1841 81 3606 82
<< m5c >>
rect 97 3645 103 3651
rect 1847 3645 1853 3651
rect 1835 3581 1841 3587
rect 3599 3581 3605 3587
rect 85 3569 91 3575
rect 1835 3569 1841 3575
rect 97 3501 103 3507
rect 1847 3501 1853 3507
rect 85 3433 91 3439
rect 1835 3433 1841 3439
rect 97 3357 103 3363
rect 1847 3357 1853 3363
rect 85 3285 91 3291
rect 1835 3285 1841 3291
rect 97 3213 103 3219
rect 1847 3213 1853 3219
rect 85 3141 91 3147
rect 1835 3141 1841 3147
rect 97 3065 103 3071
rect 1847 3065 1853 3071
rect 85 2989 91 2995
rect 1835 2989 1841 2995
rect 97 2921 103 2927
rect 1847 2921 1853 2927
rect 1847 2909 1853 2915
rect 3611 2909 3617 2915
rect 85 2849 91 2855
rect 1835 2849 1841 2855
rect 1835 2837 1841 2843
rect 3599 2837 3605 2843
rect 97 2781 103 2787
rect 1847 2781 1853 2787
rect 1847 2757 1853 2763
rect 3611 2757 3617 2763
rect 85 2705 91 2711
rect 1835 2705 1841 2711
rect 1835 2689 1841 2695
rect 3599 2689 3605 2695
rect 97 2621 103 2627
rect 1847 2621 1853 2627
rect 85 2553 91 2559
rect 1835 2553 1841 2559
rect 97 2481 103 2487
rect 1847 2481 1853 2487
rect 85 2405 91 2411
rect 1835 2405 1841 2411
rect 97 2333 103 2339
rect 1847 2333 1853 2339
rect 85 2265 91 2271
rect 1835 2265 1841 2271
rect 97 2193 103 2199
rect 1847 2193 1853 2199
rect 85 2117 91 2123
rect 1835 2117 1841 2123
rect 1847 2049 1853 2055
rect 3611 2049 3617 2055
rect 97 2037 103 2043
rect 1847 2037 1853 2043
rect 85 1969 91 1975
rect 1835 1969 1841 1975
rect 1847 1905 1853 1911
rect 3611 1905 3617 1911
rect 97 1893 103 1899
rect 1847 1893 1853 1899
rect 1835 1833 1841 1839
rect 3599 1833 3605 1839
rect 85 1825 91 1831
rect 1835 1825 1841 1831
rect 1847 1761 1853 1767
rect 3611 1761 3617 1767
rect 97 1753 103 1759
rect 1847 1753 1853 1759
rect 1835 1689 1841 1695
rect 3599 1689 3605 1695
rect 85 1681 91 1687
rect 1835 1681 1841 1687
rect 1847 1613 1853 1619
rect 3611 1613 3617 1619
rect 97 1605 103 1611
rect 1847 1605 1853 1611
rect 85 1533 91 1539
rect 1835 1533 1841 1539
rect 97 1457 103 1463
rect 1847 1457 1853 1463
rect 85 1389 91 1395
rect 1835 1389 1841 1395
rect 97 1313 103 1319
rect 1847 1313 1853 1319
rect 85 1241 91 1247
rect 1835 1241 1841 1247
rect 97 1169 103 1175
rect 1847 1169 1853 1175
rect 85 1097 91 1103
rect 1835 1097 1841 1103
rect 97 1021 103 1027
rect 1847 1021 1853 1027
rect 85 949 91 955
rect 1835 949 1841 955
rect 97 877 103 883
rect 1847 877 1853 883
rect 85 809 91 815
rect 1835 809 1841 815
rect 97 737 103 743
rect 1847 737 1853 743
rect 85 669 91 675
rect 1835 669 1841 675
rect 97 597 103 603
rect 1847 597 1853 603
rect 85 525 91 531
rect 1835 525 1841 531
rect 97 453 103 459
rect 1847 453 1853 459
rect 85 385 91 391
rect 1835 385 1841 391
rect 97 317 103 323
rect 1847 317 1853 323
rect 85 241 91 247
rect 1835 241 1841 247
rect 97 149 103 155
rect 1847 149 1853 155
rect 85 81 91 87
rect 1835 81 1841 87
<< m5 >>
rect 84 3575 92 3672
rect 84 3569 85 3575
rect 91 3569 92 3575
rect 84 3439 92 3569
rect 84 3433 85 3439
rect 91 3433 92 3439
rect 84 3291 92 3433
rect 84 3285 85 3291
rect 91 3285 92 3291
rect 84 3147 92 3285
rect 84 3141 85 3147
rect 91 3141 92 3147
rect 84 2995 92 3141
rect 84 2989 85 2995
rect 91 2989 92 2995
rect 84 2855 92 2989
rect 84 2849 85 2855
rect 91 2849 92 2855
rect 84 2711 92 2849
rect 84 2705 85 2711
rect 91 2705 92 2711
rect 84 2559 92 2705
rect 84 2553 85 2559
rect 91 2553 92 2559
rect 84 2411 92 2553
rect 84 2405 85 2411
rect 91 2405 92 2411
rect 84 2271 92 2405
rect 84 2265 85 2271
rect 91 2265 92 2271
rect 84 2123 92 2265
rect 84 2117 85 2123
rect 91 2117 92 2123
rect 84 1975 92 2117
rect 84 1969 85 1975
rect 91 1969 92 1975
rect 84 1831 92 1969
rect 84 1825 85 1831
rect 91 1825 92 1831
rect 84 1687 92 1825
rect 84 1681 85 1687
rect 91 1681 92 1687
rect 84 1539 92 1681
rect 84 1533 85 1539
rect 91 1533 92 1539
rect 84 1395 92 1533
rect 84 1389 85 1395
rect 91 1389 92 1395
rect 84 1247 92 1389
rect 84 1241 85 1247
rect 91 1241 92 1247
rect 84 1103 92 1241
rect 84 1097 85 1103
rect 91 1097 92 1103
rect 84 955 92 1097
rect 84 949 85 955
rect 91 949 92 955
rect 84 815 92 949
rect 84 809 85 815
rect 91 809 92 815
rect 84 675 92 809
rect 84 669 85 675
rect 91 669 92 675
rect 84 531 92 669
rect 84 525 85 531
rect 91 525 92 531
rect 84 391 92 525
rect 84 385 85 391
rect 91 385 92 391
rect 84 247 92 385
rect 84 241 85 247
rect 91 241 92 247
rect 84 87 92 241
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 3651 104 3672
rect 96 3645 97 3651
rect 103 3645 104 3651
rect 96 3507 104 3645
rect 96 3501 97 3507
rect 103 3501 104 3507
rect 96 3363 104 3501
rect 96 3357 97 3363
rect 103 3357 104 3363
rect 96 3219 104 3357
rect 96 3213 97 3219
rect 103 3213 104 3219
rect 96 3071 104 3213
rect 96 3065 97 3071
rect 103 3065 104 3071
rect 96 2927 104 3065
rect 96 2921 97 2927
rect 103 2921 104 2927
rect 96 2787 104 2921
rect 96 2781 97 2787
rect 103 2781 104 2787
rect 96 2627 104 2781
rect 96 2621 97 2627
rect 103 2621 104 2627
rect 96 2487 104 2621
rect 96 2481 97 2487
rect 103 2481 104 2487
rect 96 2339 104 2481
rect 96 2333 97 2339
rect 103 2333 104 2339
rect 96 2199 104 2333
rect 96 2193 97 2199
rect 103 2193 104 2199
rect 96 2043 104 2193
rect 96 2037 97 2043
rect 103 2037 104 2043
rect 96 1899 104 2037
rect 96 1893 97 1899
rect 103 1893 104 1899
rect 96 1759 104 1893
rect 96 1753 97 1759
rect 103 1753 104 1759
rect 96 1611 104 1753
rect 96 1605 97 1611
rect 103 1605 104 1611
rect 96 1463 104 1605
rect 96 1457 97 1463
rect 103 1457 104 1463
rect 96 1319 104 1457
rect 96 1313 97 1319
rect 103 1313 104 1319
rect 96 1175 104 1313
rect 96 1169 97 1175
rect 103 1169 104 1175
rect 96 1027 104 1169
rect 96 1021 97 1027
rect 103 1021 104 1027
rect 96 883 104 1021
rect 96 877 97 883
rect 103 877 104 883
rect 96 743 104 877
rect 96 737 97 743
rect 103 737 104 743
rect 96 603 104 737
rect 96 597 97 603
rect 103 597 104 603
rect 96 459 104 597
rect 96 453 97 459
rect 103 453 104 459
rect 96 323 104 453
rect 96 317 97 323
rect 103 317 104 323
rect 96 155 104 317
rect 96 149 97 155
rect 103 149 104 155
rect 96 72 104 149
rect 1834 3587 1842 3672
rect 1834 3581 1835 3587
rect 1841 3581 1842 3587
rect 1834 3575 1842 3581
rect 1834 3569 1835 3575
rect 1841 3569 1842 3575
rect 1834 3439 1842 3569
rect 1834 3433 1835 3439
rect 1841 3433 1842 3439
rect 1834 3291 1842 3433
rect 1834 3285 1835 3291
rect 1841 3285 1842 3291
rect 1834 3147 1842 3285
rect 1834 3141 1835 3147
rect 1841 3141 1842 3147
rect 1834 2995 1842 3141
rect 1834 2989 1835 2995
rect 1841 2989 1842 2995
rect 1834 2855 1842 2989
rect 1834 2849 1835 2855
rect 1841 2849 1842 2855
rect 1834 2843 1842 2849
rect 1834 2837 1835 2843
rect 1841 2837 1842 2843
rect 1834 2711 1842 2837
rect 1834 2705 1835 2711
rect 1841 2705 1842 2711
rect 1834 2695 1842 2705
rect 1834 2689 1835 2695
rect 1841 2689 1842 2695
rect 1834 2559 1842 2689
rect 1834 2553 1835 2559
rect 1841 2553 1842 2559
rect 1834 2411 1842 2553
rect 1834 2405 1835 2411
rect 1841 2405 1842 2411
rect 1834 2271 1842 2405
rect 1834 2265 1835 2271
rect 1841 2265 1842 2271
rect 1834 2123 1842 2265
rect 1834 2117 1835 2123
rect 1841 2117 1842 2123
rect 1834 1975 1842 2117
rect 1834 1969 1835 1975
rect 1841 1969 1842 1975
rect 1834 1839 1842 1969
rect 1834 1833 1835 1839
rect 1841 1833 1842 1839
rect 1834 1831 1842 1833
rect 1834 1825 1835 1831
rect 1841 1825 1842 1831
rect 1834 1695 1842 1825
rect 1834 1689 1835 1695
rect 1841 1689 1842 1695
rect 1834 1687 1842 1689
rect 1834 1681 1835 1687
rect 1841 1681 1842 1687
rect 1834 1539 1842 1681
rect 1834 1533 1835 1539
rect 1841 1533 1842 1539
rect 1834 1395 1842 1533
rect 1834 1389 1835 1395
rect 1841 1389 1842 1395
rect 1834 1247 1842 1389
rect 1834 1241 1835 1247
rect 1841 1241 1842 1247
rect 1834 1103 1842 1241
rect 1834 1097 1835 1103
rect 1841 1097 1842 1103
rect 1834 955 1842 1097
rect 1834 949 1835 955
rect 1841 949 1842 955
rect 1834 815 1842 949
rect 1834 809 1835 815
rect 1841 809 1842 815
rect 1834 675 1842 809
rect 1834 669 1835 675
rect 1841 669 1842 675
rect 1834 531 1842 669
rect 1834 525 1835 531
rect 1841 525 1842 531
rect 1834 391 1842 525
rect 1834 385 1835 391
rect 1841 385 1842 391
rect 1834 247 1842 385
rect 1834 241 1835 247
rect 1841 241 1842 247
rect 1834 87 1842 241
rect 1834 81 1835 87
rect 1841 81 1842 87
rect 1834 72 1842 81
rect 1846 3651 1854 3672
rect 1846 3645 1847 3651
rect 1853 3645 1854 3651
rect 1846 3507 1854 3645
rect 1846 3501 1847 3507
rect 1853 3501 1854 3507
rect 1846 3363 1854 3501
rect 1846 3357 1847 3363
rect 1853 3357 1854 3363
rect 1846 3219 1854 3357
rect 1846 3213 1847 3219
rect 1853 3213 1854 3219
rect 1846 3071 1854 3213
rect 1846 3065 1847 3071
rect 1853 3065 1854 3071
rect 1846 2927 1854 3065
rect 1846 2921 1847 2927
rect 1853 2921 1854 2927
rect 1846 2915 1854 2921
rect 1846 2909 1847 2915
rect 1853 2909 1854 2915
rect 1846 2787 1854 2909
rect 1846 2781 1847 2787
rect 1853 2781 1854 2787
rect 1846 2763 1854 2781
rect 1846 2757 1847 2763
rect 1853 2757 1854 2763
rect 1846 2627 1854 2757
rect 1846 2621 1847 2627
rect 1853 2621 1854 2627
rect 1846 2487 1854 2621
rect 1846 2481 1847 2487
rect 1853 2481 1854 2487
rect 1846 2339 1854 2481
rect 1846 2333 1847 2339
rect 1853 2333 1854 2339
rect 1846 2199 1854 2333
rect 1846 2193 1847 2199
rect 1853 2193 1854 2199
rect 1846 2055 1854 2193
rect 1846 2049 1847 2055
rect 1853 2049 1854 2055
rect 1846 2043 1854 2049
rect 1846 2037 1847 2043
rect 1853 2037 1854 2043
rect 1846 1911 1854 2037
rect 1846 1905 1847 1911
rect 1853 1905 1854 1911
rect 1846 1899 1854 1905
rect 1846 1893 1847 1899
rect 1853 1893 1854 1899
rect 1846 1767 1854 1893
rect 1846 1761 1847 1767
rect 1853 1761 1854 1767
rect 1846 1759 1854 1761
rect 1846 1753 1847 1759
rect 1853 1753 1854 1759
rect 1846 1619 1854 1753
rect 1846 1613 1847 1619
rect 1853 1613 1854 1619
rect 1846 1611 1854 1613
rect 1846 1605 1847 1611
rect 1853 1605 1854 1611
rect 1846 1463 1854 1605
rect 1846 1457 1847 1463
rect 1853 1457 1854 1463
rect 1846 1319 1854 1457
rect 1846 1313 1847 1319
rect 1853 1313 1854 1319
rect 1846 1175 1854 1313
rect 1846 1169 1847 1175
rect 1853 1169 1854 1175
rect 1846 1027 1854 1169
rect 1846 1021 1847 1027
rect 1853 1021 1854 1027
rect 1846 883 1854 1021
rect 1846 877 1847 883
rect 1853 877 1854 883
rect 1846 743 1854 877
rect 1846 737 1847 743
rect 1853 737 1854 743
rect 1846 603 1854 737
rect 1846 597 1847 603
rect 1853 597 1854 603
rect 1846 459 1854 597
rect 1846 453 1847 459
rect 1853 453 1854 459
rect 1846 323 1854 453
rect 1846 317 1847 323
rect 1853 317 1854 323
rect 1846 155 1854 317
rect 1846 149 1847 155
rect 1853 149 1854 155
rect 1846 72 1854 149
rect 3598 3587 3606 3672
rect 3598 3581 3599 3587
rect 3605 3581 3606 3587
rect 3598 2843 3606 3581
rect 3598 2837 3599 2843
rect 3605 2837 3606 2843
rect 3598 2695 3606 2837
rect 3598 2689 3599 2695
rect 3605 2689 3606 2695
rect 3598 1839 3606 2689
rect 3598 1833 3599 1839
rect 3605 1833 3606 1839
rect 3598 1695 3606 1833
rect 3598 1689 3599 1695
rect 3605 1689 3606 1695
rect 3598 72 3606 1689
rect 3610 2915 3618 3672
rect 3610 2909 3611 2915
rect 3617 2909 3618 2915
rect 3610 2763 3618 2909
rect 3610 2757 3611 2763
rect 3617 2757 3618 2763
rect 3610 2055 3618 2757
rect 3610 2049 3611 2055
rect 3617 2049 3618 2055
rect 3610 1911 3618 2049
rect 3610 1905 3611 1911
rect 3617 1905 3618 1911
rect 3610 1767 3618 1905
rect 3610 1761 3611 1767
rect 3617 1761 3618 1767
rect 3610 1619 3618 1761
rect 3610 1613 3611 1619
rect 3617 1613 3618 1619
rect 3610 72 3618 1613
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__193
timestamp 1731220607
transform 1 0 3568 0 -1 3568
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220607
transform 1 0 1856 0 -1 3568
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220607
transform 1 0 3568 0 1 3456
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220607
transform 1 0 1856 0 1 3456
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220607
transform 1 0 3568 0 -1 3416
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220607
transform 1 0 1856 0 -1 3416
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220607
transform 1 0 3568 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220607
transform 1 0 1856 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220607
transform 1 0 3568 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220607
transform 1 0 1856 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220607
transform 1 0 3568 0 1 3168
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220607
transform 1 0 1856 0 1 3168
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220607
transform 1 0 3568 0 -1 3132
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220607
transform 1 0 1856 0 -1 3132
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220607
transform 1 0 3568 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220607
transform 1 0 1856 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220607
transform 1 0 3568 0 -1 2980
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220607
transform 1 0 1856 0 -1 2980
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220607
transform 1 0 3568 0 1 2860
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220607
transform 1 0 1856 0 1 2860
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220607
transform 1 0 3568 0 -1 2824
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220607
transform 1 0 1856 0 -1 2824
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220607
transform 1 0 3568 0 1 2708
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220607
transform 1 0 1856 0 1 2708
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220607
transform 1 0 3568 0 -1 2676
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220607
transform 1 0 1856 0 -1 2676
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220607
transform 1 0 3568 0 1 2568
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220607
transform 1 0 1856 0 1 2568
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220607
transform 1 0 3568 0 -1 2536
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220607
transform 1 0 1856 0 -1 2536
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220607
transform 1 0 3568 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220607
transform 1 0 1856 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220607
transform 1 0 3568 0 -1 2392
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220607
transform 1 0 1856 0 -1 2392
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220607
transform 1 0 3568 0 1 2284
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220607
transform 1 0 1856 0 1 2284
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220607
transform 1 0 3568 0 -1 2252
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220607
transform 1 0 1856 0 -1 2252
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220607
transform 1 0 3568 0 1 2148
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220607
transform 1 0 1856 0 1 2148
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220607
transform 1 0 3568 0 -1 2108
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220607
transform 1 0 1856 0 -1 2108
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220607
transform 1 0 3568 0 1 2000
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220607
transform 1 0 1856 0 1 2000
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220607
transform 1 0 3568 0 -1 1960
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220607
transform 1 0 1856 0 -1 1960
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220607
transform 1 0 3568 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220607
transform 1 0 1856 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220607
transform 1 0 3568 0 -1 1820
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220607
transform 1 0 1856 0 -1 1820
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220607
transform 1 0 3568 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220607
transform 1 0 1856 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220607
transform 1 0 3568 0 -1 1676
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220607
transform 1 0 1856 0 -1 1676
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220607
transform 1 0 3568 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220607
transform 1 0 1856 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220607
transform 1 0 3568 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220607
transform 1 0 1856 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220607
transform 1 0 3568 0 1 1412
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220607
transform 1 0 1856 0 1 1412
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220607
transform 1 0 3568 0 -1 1372
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220607
transform 1 0 1856 0 -1 1372
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220607
transform 1 0 3568 0 1 1268
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220607
transform 1 0 1856 0 1 1268
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220607
transform 1 0 3568 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220607
transform 1 0 1856 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220607
transform 1 0 3568 0 1 1124
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220607
transform 1 0 1856 0 1 1124
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220607
transform 1 0 3568 0 -1 1080
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220607
transform 1 0 1856 0 -1 1080
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220607
transform 1 0 3568 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220607
transform 1 0 1856 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220607
transform 1 0 3568 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220607
transform 1 0 1856 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220607
transform 1 0 3568 0 1 832
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220607
transform 1 0 1856 0 1 832
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220607
transform 1 0 3568 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220607
transform 1 0 1856 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220607
transform 1 0 3568 0 1 692
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220607
transform 1 0 1856 0 1 692
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220607
transform 1 0 3568 0 -1 656
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220607
transform 1 0 1856 0 -1 656
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220607
transform 1 0 3568 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220607
transform 1 0 1856 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220607
transform 1 0 3568 0 -1 512
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220607
transform 1 0 1856 0 -1 512
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220607
transform 1 0 3568 0 1 408
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220607
transform 1 0 1856 0 1 408
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220607
transform 1 0 3568 0 -1 376
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220607
transform 1 0 1856 0 -1 376
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220607
transform 1 0 3568 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220607
transform 1 0 1856 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220607
transform 1 0 3568 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220607
transform 1 0 1856 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220607
transform 1 0 3568 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220607
transform 1 0 1856 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220607
transform 1 0 1816 0 1 3596
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220607
transform 1 0 104 0 1 3596
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220607
transform 1 0 1816 0 -1 3556
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220607
transform 1 0 104 0 -1 3556
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220607
transform 1 0 1816 0 1 3452
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220607
transform 1 0 104 0 1 3452
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220607
transform 1 0 1816 0 -1 3420
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220607
transform 1 0 104 0 -1 3420
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220607
transform 1 0 1816 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220607
transform 1 0 104 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220607
transform 1 0 1816 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220607
transform 1 0 104 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220607
transform 1 0 1816 0 1 3164
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220607
transform 1 0 104 0 1 3164
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220607
transform 1 0 1816 0 -1 3128
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220607
transform 1 0 104 0 -1 3128
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220607
transform 1 0 1816 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220607
transform 1 0 104 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220607
transform 1 0 1816 0 -1 2976
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220607
transform 1 0 104 0 -1 2976
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220607
transform 1 0 1816 0 1 2872
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220607
transform 1 0 104 0 1 2872
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220607
transform 1 0 1816 0 -1 2836
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220607
transform 1 0 104 0 -1 2836
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220607
transform 1 0 1816 0 1 2732
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220607
transform 1 0 104 0 1 2732
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220607
transform 1 0 1816 0 -1 2692
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220607
transform 1 0 104 0 -1 2692
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220607
transform 1 0 1816 0 1 2572
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220607
transform 1 0 104 0 1 2572
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220607
transform 1 0 1816 0 -1 2540
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220607
transform 1 0 104 0 -1 2540
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220607
transform 1 0 1816 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220607
transform 1 0 104 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220607
transform 1 0 1816 0 -1 2392
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220607
transform 1 0 104 0 -1 2392
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220607
transform 1 0 1816 0 1 2284
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220607
transform 1 0 104 0 1 2284
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220607
transform 1 0 1816 0 -1 2252
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220607
transform 1 0 104 0 -1 2252
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220607
transform 1 0 1816 0 1 2144
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220607
transform 1 0 104 0 1 2144
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220607
transform 1 0 1816 0 -1 2104
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220607
transform 1 0 104 0 -1 2104
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220607
transform 1 0 1816 0 1 1988
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220607
transform 1 0 104 0 1 1988
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220607
transform 1 0 1816 0 -1 1956
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220607
transform 1 0 104 0 -1 1956
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220607
transform 1 0 1816 0 1 1844
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220607
transform 1 0 104 0 1 1844
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220607
transform 1 0 1816 0 -1 1812
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220607
transform 1 0 104 0 -1 1812
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220607
transform 1 0 1816 0 1 1704
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220607
transform 1 0 104 0 1 1704
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220607
transform 1 0 1816 0 -1 1668
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220607
transform 1 0 104 0 -1 1668
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220607
transform 1 0 1816 0 1 1556
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220607
transform 1 0 104 0 1 1556
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220607
transform 1 0 1816 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220607
transform 1 0 104 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220607
transform 1 0 1816 0 1 1408
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220607
transform 1 0 104 0 1 1408
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220607
transform 1 0 1816 0 -1 1376
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220607
transform 1 0 104 0 -1 1376
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220607
transform 1 0 1816 0 1 1264
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220607
transform 1 0 104 0 1 1264
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220607
transform 1 0 1816 0 -1 1228
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220607
transform 1 0 104 0 -1 1228
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220607
transform 1 0 1816 0 1 1120
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220607
transform 1 0 104 0 1 1120
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220607
transform 1 0 1816 0 -1 1084
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220607
transform 1 0 104 0 -1 1084
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220607
transform 1 0 1816 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220607
transform 1 0 104 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220607
transform 1 0 1816 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220607
transform 1 0 104 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220607
transform 1 0 1816 0 1 828
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220607
transform 1 0 104 0 1 828
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220607
transform 1 0 1816 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220607
transform 1 0 104 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220607
transform 1 0 1816 0 1 688
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220607
transform 1 0 104 0 1 688
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220607
transform 1 0 1816 0 -1 656
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220607
transform 1 0 104 0 -1 656
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220607
transform 1 0 1816 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220607
transform 1 0 104 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220607
transform 1 0 1816 0 -1 512
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220607
transform 1 0 104 0 -1 512
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220607
transform 1 0 1816 0 1 404
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220607
transform 1 0 104 0 1 404
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220607
transform 1 0 1816 0 -1 372
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220607
transform 1 0 104 0 -1 372
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220607
transform 1 0 1816 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220607
transform 1 0 104 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220607
transform 1 0 1816 0 -1 228
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220607
transform 1 0 104 0 -1 228
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220607
transform 1 0 1816 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220607
transform 1 0 104 0 1 100
box 7 3 12 24
use _0_0std_0_0cells_0_0MUX2X1  tst_5999_6
timestamp 1731220607
transform 1 0 3384 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5998_6
timestamp 1731220607
transform 1 0 3472 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5997_6
timestamp 1731220607
transform 1 0 3472 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5996_6
timestamp 1731220607
transform 1 0 3472 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5995_6
timestamp 1731220607
transform 1 0 3472 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5994_6
timestamp 1731220607
transform 1 0 3472 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5993_6
timestamp 1731220607
transform 1 0 3472 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5992_6
timestamp 1731220607
transform 1 0 3472 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5991_6
timestamp 1731220607
transform 1 0 3472 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5990_6
timestamp 1731220607
transform 1 0 3472 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5989_6
timestamp 1731220607
transform 1 0 3424 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5988_6
timestamp 1731220607
transform 1 0 3312 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5987_6
timestamp 1731220607
transform 1 0 3136 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5986_6
timestamp 1731220607
transform 1 0 3320 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5985_6
timestamp 1731220607
transform 1 0 3152 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5984_6
timestamp 1731220607
transform 1 0 2984 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5983_6
timestamp 1731220607
transform 1 0 2984 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5982_6
timestamp 1731220607
transform 1 0 3152 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5981_6
timestamp 1731220607
transform 1 0 3320 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5980_6
timestamp 1731220607
transform 1 0 3312 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5979_6
timestamp 1731220607
transform 1 0 3128 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5978_6
timestamp 1731220607
transform 1 0 3088 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5977_6
timestamp 1731220607
transform 1 0 2960 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5976_6
timestamp 1731220607
transform 1 0 3344 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5975_6
timestamp 1731220607
transform 1 0 3216 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5974_6
timestamp 1731220607
transform 1 0 3144 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5973_6
timestamp 1731220607
transform 1 0 3312 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5972_6
timestamp 1731220607
transform 1 0 3456 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5971_6
timestamp 1731220607
transform 1 0 3288 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5970_6
timestamp 1731220607
transform 1 0 3120 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5969_6
timestamp 1731220607
transform 1 0 3080 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5968_6
timestamp 1731220607
transform 1 0 3280 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5967_6
timestamp 1731220607
transform 1 0 3120 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5966_6
timestamp 1731220607
transform 1 0 3304 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5965_6
timestamp 1731220607
transform 1 0 3296 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5964_6
timestamp 1731220607
transform 1 0 3208 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5963_6
timestamp 1731220607
transform 1 0 3112 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5962_6
timestamp 1731220607
transform 1 0 3016 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5961_6
timestamp 1731220607
transform 1 0 2920 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5960_6
timestamp 1731220607
transform 1 0 2824 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5959_6
timestamp 1731220607
transform 1 0 2728 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5958_6
timestamp 1731220607
transform 1 0 2632 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5957_6
timestamp 1731220607
transform 1 0 2608 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5956_6
timestamp 1731220607
transform 1 0 2776 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5955_6
timestamp 1731220607
transform 1 0 2944 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5954_6
timestamp 1731220607
transform 1 0 2888 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5953_6
timestamp 1731220607
transform 1 0 2696 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5952_6
timestamp 1731220607
transform 1 0 2496 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5951_6
timestamp 1731220607
transform 1 0 2664 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5950_6
timestamp 1731220607
transform 1 0 2808 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5949_6
timestamp 1731220607
transform 1 0 2960 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5948_6
timestamp 1731220607
transform 1 0 2984 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5947_6
timestamp 1731220607
transform 1 0 2832 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5946_6
timestamp 1731220607
transform 1 0 2832 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5945_6
timestamp 1731220607
transform 1 0 2712 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5944_6
timestamp 1731220607
transform 1 0 2664 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5943_6
timestamp 1731220607
transform 1 0 2552 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5942_6
timestamp 1731220607
transform 1 0 2800 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5941_6
timestamp 1731220607
transform 1 0 2960 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5940_6
timestamp 1731220607
transform 1 0 2824 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5939_6
timestamp 1731220607
transform 1 0 2664 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5938_6
timestamp 1731220607
transform 1 0 2624 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5937_6
timestamp 1731220607
transform 1 0 2808 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5936_6
timestamp 1731220607
transform 1 0 2960 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5935_6
timestamp 1731220607
transform 1 0 2792 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5934_6
timestamp 1731220607
transform 1 0 2616 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5933_6
timestamp 1731220607
transform 1 0 2648 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5932_6
timestamp 1731220607
transform 1 0 2832 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5931_6
timestamp 1731220607
transform 1 0 3224 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5930_6
timestamp 1731220607
transform 1 0 3024 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5929_6
timestamp 1731220607
transform 1 0 3016 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5928_6
timestamp 1731220607
transform 1 0 2880 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5927_6
timestamp 1731220607
transform 1 0 2752 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5926_6
timestamp 1731220607
transform 1 0 2624 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5925_6
timestamp 1731220607
transform 1 0 2488 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5924_6
timestamp 1731220607
transform 1 0 3016 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5923_6
timestamp 1731220607
transform 1 0 2856 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5922_6
timestamp 1731220607
transform 1 0 2704 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5921_6
timestamp 1731220607
transform 1 0 2560 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5920_6
timestamp 1731220607
transform 1 0 2560 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5919_6
timestamp 1731220607
transform 1 0 2728 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5918_6
timestamp 1731220607
transform 1 0 2904 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5917_6
timestamp 1731220607
transform 1 0 3088 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5916_6
timestamp 1731220607
transform 1 0 3128 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5915_6
timestamp 1731220607
transform 1 0 2952 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5914_6
timestamp 1731220607
transform 1 0 2776 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5913_6
timestamp 1731220607
transform 1 0 2600 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5912_6
timestamp 1731220607
transform 1 0 2768 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5911_6
timestamp 1731220607
transform 1 0 3200 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5910_6
timestamp 1731220607
transform 1 0 3056 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5909_6
timestamp 1731220607
transform 1 0 2912 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5908_6
timestamp 1731220607
transform 1 0 2872 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5907_6
timestamp 1731220607
transform 1 0 2696 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5906_6
timestamp 1731220607
transform 1 0 3032 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5905_6
timestamp 1731220607
transform 1 0 3184 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5904_6
timestamp 1731220607
transform 1 0 3336 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5903_6
timestamp 1731220607
transform 1 0 3216 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5902_6
timestamp 1731220607
transform 1 0 3072 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5901_6
timestamp 1731220607
transform 1 0 2928 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5900_6
timestamp 1731220607
transform 1 0 2776 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5899_6
timestamp 1731220607
transform 1 0 3328 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5898_6
timestamp 1731220607
transform 1 0 3160 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5897_6
timestamp 1731220607
transform 1 0 2992 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5896_6
timestamp 1731220607
transform 1 0 2832 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5895_6
timestamp 1731220607
transform 1 0 2672 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5894_6
timestamp 1731220607
transform 1 0 3144 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5893_6
timestamp 1731220607
transform 1 0 2976 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5892_6
timestamp 1731220607
transform 1 0 2816 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5891_6
timestamp 1731220607
transform 1 0 2656 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5890_6
timestamp 1731220607
transform 1 0 3080 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5889_6
timestamp 1731220607
transform 1 0 2896 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5888_6
timestamp 1731220607
transform 1 0 2728 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5887_6
timestamp 1731220607
transform 1 0 2568 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5886_6
timestamp 1731220607
transform 1 0 2536 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5885_6
timestamp 1731220607
transform 1 0 2688 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5884_6
timestamp 1731220607
transform 1 0 2856 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5883_6
timestamp 1731220607
transform 1 0 3040 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5882_6
timestamp 1731220607
transform 1 0 2976 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5881_6
timestamp 1731220607
transform 1 0 2776 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5880_6
timestamp 1731220607
transform 1 0 2632 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5879_6
timestamp 1731220607
transform 1 0 2432 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5878_6
timestamp 1731220607
transform 1 0 2824 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5877_6
timestamp 1731220607
transform 1 0 3008 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5876_6
timestamp 1731220607
transform 1 0 3192 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5875_6
timestamp 1731220607
transform 1 0 3184 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5874_6
timestamp 1731220607
transform 1 0 3232 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5873_6
timestamp 1731220607
transform 1 0 3264 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5872_6
timestamp 1731220607
transform 1 0 3312 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5871_6
timestamp 1731220607
transform 1 0 3352 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5870_6
timestamp 1731220607
transform 1 0 3344 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5869_6
timestamp 1731220607
transform 1 0 3312 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5868_6
timestamp 1731220607
transform 1 0 3280 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5867_6
timestamp 1731220607
transform 1 0 3176 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5866_6
timestamp 1731220607
transform 1 0 3336 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5865_6
timestamp 1731220607
transform 1 0 3472 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5864_6
timestamp 1731220607
transform 1 0 3472 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5863_6
timestamp 1731220607
transform 1 0 3472 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5862_6
timestamp 1731220607
transform 1 0 3472 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5861_6
timestamp 1731220607
transform 1 0 3472 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5860_6
timestamp 1731220607
transform 1 0 3472 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5859_6
timestamp 1731220607
transform 1 0 3472 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5858_6
timestamp 1731220607
transform 1 0 3472 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5857_6
timestamp 1731220607
transform 1 0 3456 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5856_6
timestamp 1731220607
transform 1 0 3424 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5855_6
timestamp 1731220607
transform 1 0 3400 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5854_6
timestamp 1731220607
transform 1 0 3384 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5853_6
timestamp 1731220607
transform 1 0 3200 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5852_6
timestamp 1731220607
transform 1 0 3056 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5851_6
timestamp 1731220607
transform 1 0 2904 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5850_6
timestamp 1731220607
transform 1 0 3328 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5849_6
timestamp 1731220607
transform 1 0 3160 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5848_6
timestamp 1731220607
transform 1 0 2992 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5847_6
timestamp 1731220607
transform 1 0 2808 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5846_6
timestamp 1731220607
transform 1 0 2608 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5845_6
timestamp 1731220607
transform 1 0 3232 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5844_6
timestamp 1731220607
transform 1 0 3048 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5843_6
timestamp 1731220607
transform 1 0 2864 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5842_6
timestamp 1731220607
transform 1 0 2696 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5841_6
timestamp 1731220607
transform 1 0 3296 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5840_6
timestamp 1731220607
transform 1 0 3096 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5839_6
timestamp 1731220607
transform 1 0 2912 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5838_6
timestamp 1731220607
transform 1 0 2744 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5837_6
timestamp 1731220607
transform 1 0 2608 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5836_6
timestamp 1731220607
transform 1 0 3272 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5835_6
timestamp 1731220607
transform 1 0 3056 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5834_6
timestamp 1731220607
transform 1 0 2856 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5833_6
timestamp 1731220607
transform 1 0 2680 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5832_6
timestamp 1731220607
transform 1 0 2728 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5831_6
timestamp 1731220607
transform 1 0 3096 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5830_6
timestamp 1731220607
transform 1 0 2904 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5829_6
timestamp 1731220607
transform 1 0 2864 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5828_6
timestamp 1731220607
transform 1 0 2688 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5827_6
timestamp 1731220607
transform 1 0 3064 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5826_6
timestamp 1731220607
transform 1 0 3272 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5825_6
timestamp 1731220607
transform 1 0 3128 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5824_6
timestamp 1731220607
transform 1 0 2960 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5823_6
timestamp 1731220607
transform 1 0 2800 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5822_6
timestamp 1731220607
transform 1 0 2648 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5821_6
timestamp 1731220607
transform 1 0 2752 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5820_6
timestamp 1731220607
transform 1 0 2928 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5819_6
timestamp 1731220607
transform 1 0 3104 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5818_6
timestamp 1731220607
transform 1 0 3048 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5817_6
timestamp 1731220607
transform 1 0 2896 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5816_6
timestamp 1731220607
transform 1 0 2736 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5815_6
timestamp 1731220607
transform 1 0 2856 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5814_6
timestamp 1731220607
transform 1 0 3064 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5813_6
timestamp 1731220607
transform 1 0 3280 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5812_6
timestamp 1731220607
transform 1 0 3192 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5811_6
timestamp 1731220607
transform 1 0 3336 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5810_6
timestamp 1731220607
transform 1 0 3280 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5809_6
timestamp 1731220607
transform 1 0 3296 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5808_6
timestamp 1731220607
transform 1 0 3296 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5807_6
timestamp 1731220607
transform 1 0 3424 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5806_6
timestamp 1731220607
transform 1 0 3344 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5805_6
timestamp 1731220607
transform 1 0 3472 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5804_6
timestamp 1731220607
transform 1 0 3472 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5803_6
timestamp 1731220607
transform 1 0 3472 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5802_6
timestamp 1731220607
transform 1 0 3472 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5801_6
timestamp 1731220607
transform 1 0 3472 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5800_6
timestamp 1731220607
transform 1 0 3472 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5799_6
timestamp 1731220607
transform 1 0 3464 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5798_6
timestamp 1731220607
transform 1 0 3456 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5797_6
timestamp 1731220607
transform 1 0 3472 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5796_6
timestamp 1731220607
transform 1 0 3472 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5795_6
timestamp 1731220607
transform 1 0 3472 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5794_6
timestamp 1731220607
transform 1 0 3472 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5793_6
timestamp 1731220607
transform 1 0 3472 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5792_6
timestamp 1731220607
transform 1 0 3472 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5791_6
timestamp 1731220607
transform 1 0 3472 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5790_6
timestamp 1731220607
transform 1 0 3472 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5789_6
timestamp 1731220607
transform 1 0 3472 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5788_6
timestamp 1731220607
transform 1 0 3312 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5787_6
timestamp 1731220607
transform 1 0 3184 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5786_6
timestamp 1731220607
transform 1 0 3336 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5785_6
timestamp 1731220607
transform 1 0 3336 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5784_6
timestamp 1731220607
transform 1 0 3184 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5783_6
timestamp 1731220607
transform 1 0 3032 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5782_6
timestamp 1731220607
transform 1 0 2864 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5781_6
timestamp 1731220607
transform 1 0 2864 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5780_6
timestamp 1731220607
transform 1 0 3024 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5779_6
timestamp 1731220607
transform 1 0 3144 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5778_6
timestamp 1731220607
transform 1 0 2976 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5777_6
timestamp 1731220607
transform 1 0 2808 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5776_6
timestamp 1731220607
transform 1 0 2864 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5775_6
timestamp 1731220607
transform 1 0 3040 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5774_6
timestamp 1731220607
transform 1 0 3016 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5773_6
timestamp 1731220607
transform 1 0 2880 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5772_6
timestamp 1731220607
transform 1 0 2752 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5771_6
timestamp 1731220607
transform 1 0 2784 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5770_6
timestamp 1731220607
transform 1 0 2928 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5769_6
timestamp 1731220607
transform 1 0 3072 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5768_6
timestamp 1731220607
transform 1 0 3288 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5767_6
timestamp 1731220607
transform 1 0 3200 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5766_6
timestamp 1731220607
transform 1 0 3112 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5765_6
timestamp 1731220607
transform 1 0 3024 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5764_6
timestamp 1731220607
transform 1 0 2936 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5763_6
timestamp 1731220607
transform 1 0 2848 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5762_6
timestamp 1731220607
transform 1 0 2760 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5761_6
timestamp 1731220607
transform 1 0 2672 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5760_6
timestamp 1731220607
transform 1 0 2584 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5759_6
timestamp 1731220607
transform 1 0 2648 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5758_6
timestamp 1731220607
transform 1 0 2624 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5757_6
timestamp 1731220607
transform 1 0 2496 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5756_6
timestamp 1731220607
transform 1 0 2688 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5755_6
timestamp 1731220607
transform 1 0 2632 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5754_6
timestamp 1731220607
transform 1 0 2688 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5753_6
timestamp 1731220607
transform 1 0 2688 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5752_6
timestamp 1731220607
transform 1 0 2576 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5751_6
timestamp 1731220607
transform 1 0 2736 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5750_6
timestamp 1731220607
transform 1 0 3072 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5749_6
timestamp 1731220607
transform 1 0 2904 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5748_6
timestamp 1731220607
transform 1 0 2856 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5747_6
timestamp 1731220607
transform 1 0 2664 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5746_6
timestamp 1731220607
transform 1 0 3024 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5745_6
timestamp 1731220607
transform 1 0 3184 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5744_6
timestamp 1731220607
transform 1 0 3336 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5743_6
timestamp 1731220607
transform 1 0 3320 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5742_6
timestamp 1731220607
transform 1 0 3168 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5741_6
timestamp 1731220607
transform 1 0 3008 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5740_6
timestamp 1731220607
transform 1 0 2840 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5739_6
timestamp 1731220607
transform 1 0 2656 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5738_6
timestamp 1731220607
transform 1 0 3168 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5737_6
timestamp 1731220607
transform 1 0 3320 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5736_6
timestamp 1731220607
transform 1 0 3256 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5735_6
timestamp 1731220607
transform 1 0 3064 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5734_6
timestamp 1731220607
transform 1 0 2952 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5733_6
timestamp 1731220607
transform 1 0 2840 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5732_6
timestamp 1731220607
transform 1 0 2728 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5731_6
timestamp 1731220607
transform 1 0 2624 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5730_6
timestamp 1731220607
transform 1 0 2512 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5729_6
timestamp 1731220607
transform 1 0 2608 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5728_6
timestamp 1731220607
transform 1 0 2808 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5727_6
timestamp 1731220607
transform 1 0 3024 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5726_6
timestamp 1731220607
transform 1 0 3024 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5725_6
timestamp 1731220607
transform 1 0 2896 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5724_6
timestamp 1731220607
transform 1 0 2784 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5723_6
timestamp 1731220607
transform 1 0 2680 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5722_6
timestamp 1731220607
transform 1 0 2592 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5721_6
timestamp 1731220607
transform 1 0 2328 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5720_6
timestamp 1731220607
transform 1 0 2240 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5719_6
timestamp 1731220607
transform 1 0 2152 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5718_6
timestamp 1731220607
transform 1 0 2064 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5717_6
timestamp 1731220607
transform 1 0 1976 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5716_6
timestamp 1731220607
transform 1 0 1888 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5715_6
timestamp 1731220607
transform 1 0 2280 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5714_6
timestamp 1731220607
transform 1 0 2152 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5713_6
timestamp 1731220607
transform 1 0 2032 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5712_6
timestamp 1731220607
transform 1 0 1936 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5711_6
timestamp 1731220607
transform 1 0 2048 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5710_6
timestamp 1731220607
transform 1 0 2160 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5709_6
timestamp 1731220607
transform 1 0 2248 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5708_6
timestamp 1731220607
transform 1 0 2056 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5707_6
timestamp 1731220607
transform 1 0 1880 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5706_6
timestamp 1731220607
transform 1 0 1880 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5705_6
timestamp 1731220607
transform 1 0 2032 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5704_6
timestamp 1731220607
transform 1 0 2208 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5703_6
timestamp 1731220607
transform 1 0 2264 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5702_6
timestamp 1731220607
transform 1 0 2112 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5701_6
timestamp 1731220607
transform 1 0 1976 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5700_6
timestamp 1731220607
transform 1 0 1880 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5699_6
timestamp 1731220607
transform 1 0 1720 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5698_6
timestamp 1731220607
transform 1 0 1632 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5697_6
timestamp 1731220607
transform 1 0 1536 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5696_6
timestamp 1731220607
transform 1 0 1432 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5695_6
timestamp 1731220607
transform 1 0 1328 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5694_6
timestamp 1731220607
transform 1 0 1224 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5693_6
timestamp 1731220607
transform 1 0 1448 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5692_6
timestamp 1731220607
transform 1 0 1584 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5691_6
timestamp 1731220607
transform 1 0 1720 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5690_6
timestamp 1731220607
transform 1 0 1592 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5689_6
timestamp 1731220607
transform 1 0 1392 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5688_6
timestamp 1731220607
transform 1 0 1200 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5687_6
timestamp 1731220607
transform 1 0 1312 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5686_6
timestamp 1731220607
transform 1 0 1168 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5685_6
timestamp 1731220607
transform 1 0 1016 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5684_6
timestamp 1731220607
transform 1 0 992 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5683_6
timestamp 1731220607
transform 1 0 1112 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5682_6
timestamp 1731220607
transform 1 0 1424 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5681_6
timestamp 1731220607
transform 1 0 1296 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5680_6
timestamp 1731220607
transform 1 0 1168 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5679_6
timestamp 1731220607
transform 1 0 1040 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5678_6
timestamp 1731220607
transform 1 0 912 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5677_6
timestamp 1731220607
transform 1 0 1264 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5676_6
timestamp 1731220607
transform 1 0 1144 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5675_6
timestamp 1731220607
transform 1 0 1024 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5674_6
timestamp 1731220607
transform 1 0 912 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5673_6
timestamp 1731220607
transform 1 0 792 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5672_6
timestamp 1731220607
transform 1 0 704 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5671_6
timestamp 1731220607
transform 1 0 816 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5670_6
timestamp 1731220607
transform 1 0 1168 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5669_6
timestamp 1731220607
transform 1 0 1048 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5668_6
timestamp 1731220607
transform 1 0 928 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5667_6
timestamp 1731220607
transform 1 0 896 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5666_6
timestamp 1731220607
transform 1 0 768 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5665_6
timestamp 1731220607
transform 1 0 1016 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5664_6
timestamp 1731220607
transform 1 0 1144 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5663_6
timestamp 1731220607
transform 1 0 1272 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5662_6
timestamp 1731220607
transform 1 0 1168 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5661_6
timestamp 1731220607
transform 1 0 1048 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5660_6
timestamp 1731220607
transform 1 0 936 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5659_6
timestamp 1731220607
transform 1 0 824 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5658_6
timestamp 1731220607
transform 1 0 712 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5657_6
timestamp 1731220607
transform 1 0 792 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5656_6
timestamp 1731220607
transform 1 0 680 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5655_6
timestamp 1731220607
transform 1 0 712 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5654_6
timestamp 1731220607
transform 1 0 704 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5653_6
timestamp 1731220607
transform 1 0 752 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5652_6
timestamp 1731220607
transform 1 0 920 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5651_6
timestamp 1731220607
transform 1 0 904 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5650_6
timestamp 1731220607
transform 1 0 752 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5649_6
timestamp 1731220607
transform 1 0 880 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5648_6
timestamp 1731220607
transform 1 0 728 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5647_6
timestamp 1731220607
transform 1 0 744 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5646_6
timestamp 1731220607
transform 1 0 608 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5645_6
timestamp 1731220607
transform 1 0 576 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5644_6
timestamp 1731220607
transform 1 0 728 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5643_6
timestamp 1731220607
transform 1 0 648 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5642_6
timestamp 1731220607
transform 1 0 520 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5641_6
timestamp 1731220607
transform 1 0 776 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5640_6
timestamp 1731220607
transform 1 0 1016 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5639_6
timestamp 1731220607
transform 1 0 888 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5638_6
timestamp 1731220607
transform 1 0 704 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5637_6
timestamp 1731220607
transform 1 0 512 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5636_6
timestamp 1731220607
transform 1 0 648 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5635_6
timestamp 1731220607
transform 1 0 808 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5634_6
timestamp 1731220607
transform 1 0 744 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5633_6
timestamp 1731220607
transform 1 0 600 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5632_6
timestamp 1731220607
transform 1 0 672 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5631_6
timestamp 1731220607
transform 1 0 640 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5630_6
timestamp 1731220607
transform 1 0 776 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5629_6
timestamp 1731220607
transform 1 0 840 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5628_6
timestamp 1731220607
transform 1 0 696 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5627_6
timestamp 1731220607
transform 1 0 568 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5626_6
timestamp 1731220607
transform 1 0 632 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5625_6
timestamp 1731220607
transform 1 0 768 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5624_6
timestamp 1731220607
transform 1 0 816 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5623_6
timestamp 1731220607
transform 1 0 672 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5622_6
timestamp 1731220607
transform 1 0 632 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5621_6
timestamp 1731220607
transform 1 0 776 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5620_6
timestamp 1731220607
transform 1 0 768 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5619_6
timestamp 1731220607
transform 1 0 616 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5618_6
timestamp 1731220607
transform 1 0 656 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5617_6
timestamp 1731220607
transform 1 0 832 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5616_6
timestamp 1731220607
transform 1 0 672 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5615_6
timestamp 1731220607
transform 1 0 856 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5614_6
timestamp 1731220607
transform 1 0 864 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5613_6
timestamp 1731220607
transform 1 0 672 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5612_6
timestamp 1731220607
transform 1 0 584 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5611_6
timestamp 1731220607
transform 1 0 760 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5610_6
timestamp 1731220607
transform 1 0 776 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5609_6
timestamp 1731220607
transform 1 0 624 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5608_6
timestamp 1731220607
transform 1 0 480 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5607_6
timestamp 1731220607
transform 1 0 616 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5606_6
timestamp 1731220607
transform 1 0 752 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5605_6
timestamp 1731220607
transform 1 0 776 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5604_6
timestamp 1731220607
transform 1 0 688 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5603_6
timestamp 1731220607
transform 1 0 600 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5602_6
timestamp 1731220607
transform 1 0 512 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5601_6
timestamp 1731220607
transform 1 0 424 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5600_6
timestamp 1731220607
transform 1 0 336 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5599_6
timestamp 1731220607
transform 1 0 248 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5598_6
timestamp 1731220607
transform 1 0 160 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5597_6
timestamp 1731220607
transform 1 0 224 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5596_6
timestamp 1731220607
transform 1 0 480 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5595_6
timestamp 1731220607
transform 1 0 352 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5594_6
timestamp 1731220607
transform 1 0 336 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5593_6
timestamp 1731220607
transform 1 0 200 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5592_6
timestamp 1731220607
transform 1 0 128 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5591_6
timestamp 1731220607
transform 1 0 256 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5590_6
timestamp 1731220607
transform 1 0 416 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5589_6
timestamp 1731220607
transform 1 0 480 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5588_6
timestamp 1731220607
transform 1 0 288 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5587_6
timestamp 1731220607
transform 1 0 128 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5586_6
timestamp 1731220607
transform 1 0 128 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5585_6
timestamp 1731220607
transform 1 0 296 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5584_6
timestamp 1731220607
transform 1 0 488 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5583_6
timestamp 1731220607
transform 1 0 472 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5582_6
timestamp 1731220607
transform 1 0 288 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5581_6
timestamp 1731220607
transform 1 0 128 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5580_6
timestamp 1731220607
transform 1 0 128 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5579_6
timestamp 1731220607
transform 1 0 288 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5578_6
timestamp 1731220607
transform 1 0 456 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5577_6
timestamp 1731220607
transform 1 0 488 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5576_6
timestamp 1731220607
transform 1 0 344 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5575_6
timestamp 1731220607
transform 1 0 200 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5574_6
timestamp 1731220607
transform 1 0 280 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5573_6
timestamp 1731220607
transform 1 0 528 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5572_6
timestamp 1731220607
transform 1 0 400 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5571_6
timestamp 1731220607
transform 1 0 328 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5570_6
timestamp 1731220607
transform 1 0 416 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5569_6
timestamp 1731220607
transform 1 0 520 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5568_6
timestamp 1731220607
transform 1 0 456 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5567_6
timestamp 1731220607
transform 1 0 360 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5566_6
timestamp 1731220607
transform 1 0 328 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5565_6
timestamp 1731220607
transform 1 0 416 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5564_6
timestamp 1731220607
transform 1 0 520 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5563_6
timestamp 1731220607
transform 1 0 552 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5562_6
timestamp 1731220607
transform 1 0 432 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5561_6
timestamp 1731220607
transform 1 0 320 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5560_6
timestamp 1731220607
transform 1 0 208 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5559_6
timestamp 1731220607
transform 1 0 152 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5558_6
timestamp 1731220607
transform 1 0 304 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5557_6
timestamp 1731220607
transform 1 0 456 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5556_6
timestamp 1731220607
transform 1 0 472 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5555_6
timestamp 1731220607
transform 1 0 288 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5554_6
timestamp 1731220607
transform 1 0 128 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5553_6
timestamp 1731220607
transform 1 0 312 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5552_6
timestamp 1731220607
transform 1 0 128 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5551_6
timestamp 1731220607
transform 1 0 128 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5550_6
timestamp 1731220607
transform 1 0 320 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5549_6
timestamp 1731220607
transform 1 0 544 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5548_6
timestamp 1731220607
transform 1 0 384 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5547_6
timestamp 1731220607
transform 1 0 248 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5546_6
timestamp 1731220607
transform 1 0 128 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5545_6
timestamp 1731220607
transform 1 0 128 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5544_6
timestamp 1731220607
transform 1 0 264 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5543_6
timestamp 1731220607
transform 1 0 416 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5542_6
timestamp 1731220607
transform 1 0 472 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5541_6
timestamp 1731220607
transform 1 0 336 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5540_6
timestamp 1731220607
transform 1 0 208 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5539_6
timestamp 1731220607
transform 1 0 304 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5538_6
timestamp 1731220607
transform 1 0 440 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5537_6
timestamp 1731220607
transform 1 0 584 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5536_6
timestamp 1731220607
transform 1 0 456 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5535_6
timestamp 1731220607
transform 1 0 312 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5534_6
timestamp 1731220607
transform 1 0 600 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5533_6
timestamp 1731220607
transform 1 0 584 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5532_6
timestamp 1731220607
transform 1 0 408 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5531_6
timestamp 1731220607
transform 1 0 240 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5530_6
timestamp 1731220607
transform 1 0 208 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5529_6
timestamp 1731220607
transform 1 0 464 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5528_6
timestamp 1731220607
transform 1 0 288 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5527_6
timestamp 1731220607
transform 1 0 152 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5526_6
timestamp 1731220607
transform 1 0 152 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5525_6
timestamp 1731220607
transform 1 0 128 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5524_6
timestamp 1731220607
transform 1 0 224 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5523_6
timestamp 1731220607
transform 1 0 232 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5522_6
timestamp 1731220607
transform 1 0 128 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5521_6
timestamp 1731220607
transform 1 0 128 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5520_6
timestamp 1731220607
transform 1 0 224 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5519_6
timestamp 1731220607
transform 1 0 344 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5518_6
timestamp 1731220607
transform 1 0 248 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5517_6
timestamp 1731220607
transform 1 0 128 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5516_6
timestamp 1731220607
transform 1 0 144 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5515_6
timestamp 1731220607
transform 1 0 312 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5514_6
timestamp 1731220607
transform 1 0 448 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5513_6
timestamp 1731220607
transform 1 0 304 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5512_6
timestamp 1731220607
transform 1 0 168 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5511_6
timestamp 1731220607
transform 1 0 264 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5510_6
timestamp 1731220607
transform 1 0 464 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5509_6
timestamp 1731220607
transform 1 0 480 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5508_6
timestamp 1731220607
transform 1 0 336 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5507_6
timestamp 1731220607
transform 1 0 208 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5506_6
timestamp 1731220607
transform 1 0 160 0 -1 2708
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5505_6
timestamp 1731220607
transform 1 0 272 0 -1 2708
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5504_6
timestamp 1731220607
transform 1 0 384 0 -1 2708
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5503_6
timestamp 1731220607
transform 1 0 400 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5502_6
timestamp 1731220607
transform 1 0 280 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5501_6
timestamp 1731220607
transform 1 0 176 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5500_6
timestamp 1731220607
transform 1 0 128 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5499_6
timestamp 1731220607
transform 1 0 216 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5498_6
timestamp 1731220607
transform 1 0 304 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5497_6
timestamp 1731220607
transform 1 0 392 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5496_6
timestamp 1731220607
transform 1 0 480 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5495_6
timestamp 1731220607
transform 1 0 592 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5494_6
timestamp 1731220607
transform 1 0 720 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5493_6
timestamp 1731220607
transform 1 0 992 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5492_6
timestamp 1731220607
transform 1 0 856 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5491_6
timestamp 1731220607
transform 1 0 808 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5490_6
timestamp 1731220607
transform 1 0 672 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5489_6
timestamp 1731220607
transform 1 0 536 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5488_6
timestamp 1731220607
transform 1 0 496 0 -1 2708
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5487_6
timestamp 1731220607
transform 1 0 608 0 -1 2708
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5486_6
timestamp 1731220607
transform 1 0 648 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5485_6
timestamp 1731220607
transform 1 0 824 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5484_6
timestamp 1731220607
transform 1 0 1008 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5483_6
timestamp 1731220607
transform 1 0 848 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5482_6
timestamp 1731220607
transform 1 0 664 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5481_6
timestamp 1731220607
transform 1 0 864 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5480_6
timestamp 1731220607
transform 1 0 728 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5479_6
timestamp 1731220607
transform 1 0 592 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5478_6
timestamp 1731220607
transform 1 0 472 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5477_6
timestamp 1731220607
transform 1 0 632 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5476_6
timestamp 1731220607
transform 1 0 776 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5475_6
timestamp 1731220607
transform 1 0 664 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5474_6
timestamp 1731220607
transform 1 0 528 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5473_6
timestamp 1731220607
transform 1 0 392 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5472_6
timestamp 1731220607
transform 1 0 464 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5471_6
timestamp 1731220607
transform 1 0 584 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5470_6
timestamp 1731220607
transform 1 0 640 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5469_6
timestamp 1731220607
transform 1 0 504 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5468_6
timestamp 1731220607
transform 1 0 368 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5467_6
timestamp 1731220607
transform 1 0 352 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5466_6
timestamp 1731220607
transform 1 0 472 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5465_6
timestamp 1731220607
transform 1 0 592 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5464_6
timestamp 1731220607
transform 1 0 560 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5463_6
timestamp 1731220607
transform 1 0 432 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5462_6
timestamp 1731220607
transform 1 0 296 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5461_6
timestamp 1731220607
transform 1 0 432 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5460_6
timestamp 1731220607
transform 1 0 576 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5459_6
timestamp 1731220607
transform 1 0 848 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5458_6
timestamp 1731220607
transform 1 0 984 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5457_6
timestamp 1731220607
transform 1 0 896 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5456_6
timestamp 1731220607
transform 1 0 1000 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5455_6
timestamp 1731220607
transform 1 0 1104 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5454_6
timestamp 1731220607
transform 1 0 1208 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5453_6
timestamp 1731220607
transform 1 0 1312 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5452_6
timestamp 1731220607
transform 1 0 1232 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5451_6
timestamp 1731220607
transform 1 0 1112 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5450_6
timestamp 1731220607
transform 1 0 1352 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5449_6
timestamp 1731220607
transform 1 0 1472 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5448_6
timestamp 1731220607
transform 1 0 1592 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5447_6
timestamp 1731220607
transform 1 0 1592 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5446_6
timestamp 1731220607
transform 1 0 1440 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5445_6
timestamp 1731220607
transform 1 0 1280 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5444_6
timestamp 1731220607
transform 1 0 1112 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5443_6
timestamp 1731220607
transform 1 0 920 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5442_6
timestamp 1731220607
transform 1 0 1072 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5441_6
timestamp 1731220607
transform 1 0 1216 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5440_6
timestamp 1731220607
transform 1 0 1352 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5439_6
timestamp 1731220607
transform 1 0 1360 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5438_6
timestamp 1731220607
transform 1 0 1208 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5437_6
timestamp 1731220607
transform 1 0 1056 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5436_6
timestamp 1731220607
transform 1 0 1032 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5435_6
timestamp 1731220607
transform 1 0 1184 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5434_6
timestamp 1731220607
transform 1 0 1200 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5433_6
timestamp 1731220607
transform 1 0 1040 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5432_6
timestamp 1731220607
transform 1 0 888 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5431_6
timestamp 1731220607
transform 1 0 880 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5430_6
timestamp 1731220607
transform 1 0 1032 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5429_6
timestamp 1731220607
transform 1 0 1008 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5428_6
timestamp 1731220607
transform 1 0 896 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5427_6
timestamp 1731220607
transform 1 0 776 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5426_6
timestamp 1731220607
transform 1 0 1128 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5425_6
timestamp 1731220607
transform 1 0 1248 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5424_6
timestamp 1731220607
transform 1 0 1488 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5423_6
timestamp 1731220607
transform 1 0 1368 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5422_6
timestamp 1731220607
transform 1 0 1336 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5421_6
timestamp 1731220607
transform 1 0 1184 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5420_6
timestamp 1731220607
transform 1 0 1488 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5419_6
timestamp 1731220607
transform 1 0 1528 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5418_6
timestamp 1731220607
transform 1 0 1360 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5417_6
timestamp 1731220607
transform 1 0 1336 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5416_6
timestamp 1731220607
transform 1 0 1488 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5415_6
timestamp 1731220607
transform 1 0 1640 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5414_6
timestamp 1731220607
transform 1 0 1672 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5413_6
timestamp 1731220607
transform 1 0 1512 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5412_6
timestamp 1731220607
transform 1 0 1480 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5411_6
timestamp 1731220607
transform 1 0 1608 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5410_6
timestamp 1731220607
transform 1 0 1720 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5409_6
timestamp 1731220607
transform 1 0 1720 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5408_6
timestamp 1731220607
transform 1 0 1880 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5407_6
timestamp 1731220607
transform 1 0 2056 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5406_6
timestamp 1731220607
transform 1 0 1968 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5405_6
timestamp 1731220607
transform 1 0 1896 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5404_6
timestamp 1731220607
transform 1 0 2432 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5403_6
timestamp 1731220607
transform 1 0 2280 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5402_6
timestamp 1731220607
transform 1 0 2152 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5401_6
timestamp 1731220607
transform 1 0 1992 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5400_6
timestamp 1731220607
transform 1 0 1928 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5399_6
timestamp 1731220607
transform 1 0 2072 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5398_6
timestamp 1731220607
transform 1 0 2232 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5397_6
timestamp 1731220607
transform 1 0 2144 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5396_6
timestamp 1731220607
transform 1 0 2024 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5395_6
timestamp 1731220607
transform 1 0 1904 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5394_6
timestamp 1731220607
transform 1 0 1880 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5393_6
timestamp 1731220607
transform 1 0 2000 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5392_6
timestamp 1731220607
transform 1 0 2136 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5391_6
timestamp 1731220607
transform 1 0 2016 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5390_6
timestamp 1731220607
transform 1 0 1880 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5389_6
timestamp 1731220607
transform 1 0 1720 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5388_6
timestamp 1731220607
transform 1 0 1616 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5387_6
timestamp 1731220607
transform 1 0 1496 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5386_6
timestamp 1731220607
transform 1 0 1256 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5385_6
timestamp 1731220607
transform 1 0 1720 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5384_6
timestamp 1731220607
transform 1 0 1672 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5383_6
timestamp 1731220607
transform 1 0 1520 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5382_6
timestamp 1731220607
transform 1 0 1368 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5381_6
timestamp 1731220607
transform 1 0 1216 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5380_6
timestamp 1731220607
transform 1 0 1056 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5379_6
timestamp 1731220607
transform 1 0 1520 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5378_6
timestamp 1731220607
transform 1 0 1376 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5377_6
timestamp 1731220607
transform 1 0 1240 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5376_6
timestamp 1731220607
transform 1 0 1104 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5375_6
timestamp 1731220607
transform 1 0 960 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5374_6
timestamp 1731220607
transform 1 0 1560 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5373_6
timestamp 1731220607
transform 1 0 1384 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5372_6
timestamp 1731220607
transform 1 0 1216 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5371_6
timestamp 1731220607
transform 1 0 1048 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5370_6
timestamp 1731220607
transform 1 0 896 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5369_6
timestamp 1731220607
transform 1 0 1400 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5368_6
timestamp 1731220607
transform 1 0 1240 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5367_6
timestamp 1731220607
transform 1 0 1080 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5366_6
timestamp 1731220607
transform 1 0 936 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5365_6
timestamp 1731220607
transform 1 0 800 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5364_6
timestamp 1731220607
transform 1 0 936 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5363_6
timestamp 1731220607
transform 1 0 1120 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5362_6
timestamp 1731220607
transform 1 0 1312 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5361_6
timestamp 1731220607
transform 1 0 1168 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5360_6
timestamp 1731220607
transform 1 0 1000 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5359_6
timestamp 1731220607
transform 1 0 912 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5358_6
timestamp 1731220607
transform 1 0 1072 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5357_6
timestamp 1731220607
transform 1 0 1248 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5356_6
timestamp 1731220607
transform 1 0 1120 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5355_6
timestamp 1731220607
transform 1 0 968 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5354_6
timestamp 1731220607
transform 1 0 920 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5353_6
timestamp 1731220607
transform 1 0 1232 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5352_6
timestamp 1731220607
transform 1 0 1072 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5351_6
timestamp 1731220607
transform 1 0 1064 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5350_6
timestamp 1731220607
transform 1 0 920 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5349_6
timestamp 1731220607
transform 1 0 1008 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5348_6
timestamp 1731220607
transform 1 0 1024 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5347_6
timestamp 1731220607
transform 1 0 1040 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5346_6
timestamp 1731220607
transform 1 0 1096 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5345_6
timestamp 1731220607
transform 1 0 928 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5344_6
timestamp 1731220607
transform 1 0 920 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5343_6
timestamp 1731220607
transform 1 0 1064 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5342_6
timestamp 1731220607
transform 1 0 1024 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5341_6
timestamp 1731220607
transform 1 0 888 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5340_6
timestamp 1731220607
transform 1 0 864 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5339_6
timestamp 1731220607
transform 1 0 952 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5338_6
timestamp 1731220607
transform 1 0 1040 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5337_6
timestamp 1731220607
transform 1 0 1128 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5336_6
timestamp 1731220607
transform 1 0 1216 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5335_6
timestamp 1731220607
transform 1 0 1488 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5334_6
timestamp 1731220607
transform 1 0 1392 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5333_6
timestamp 1731220607
transform 1 0 1304 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5332_6
timestamp 1731220607
transform 1 0 1288 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5331_6
timestamp 1731220607
transform 1 0 1152 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5330_6
timestamp 1731220607
transform 1 0 1424 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5329_6
timestamp 1731220607
transform 1 0 1472 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5328_6
timestamp 1731220607
transform 1 0 1344 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5327_6
timestamp 1731220607
transform 1 0 1208 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5326_6
timestamp 1731220607
transform 1 0 1256 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5325_6
timestamp 1731220607
transform 1 0 1208 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5324_6
timestamp 1731220607
transform 1 0 1376 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5323_6
timestamp 1731220607
transform 1 0 1344 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5322_6
timestamp 1731220607
transform 1 0 1184 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5321_6
timestamp 1731220607
transform 1 0 1184 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5320_6
timestamp 1731220607
transform 1 0 1360 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5319_6
timestamp 1731220607
transform 1 0 1336 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5318_6
timestamp 1731220607
transform 1 0 1200 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5317_6
timestamp 1731220607
transform 1 0 1472 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5316_6
timestamp 1731220607
transform 1 0 1568 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5315_6
timestamp 1731220607
transform 1 0 1400 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5314_6
timestamp 1731220607
transform 1 0 1272 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5313_6
timestamp 1731220607
transform 1 0 1592 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5312_6
timestamp 1731220607
transform 1 0 1432 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5311_6
timestamp 1731220607
transform 1 0 1432 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5310_6
timestamp 1731220607
transform 1 0 1616 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5309_6
timestamp 1731220607
transform 1 0 1520 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5308_6
timestamp 1731220607
transform 1 0 1344 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5307_6
timestamp 1731220607
transform 1 0 1704 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5306_6
timestamp 1731220607
transform 1 0 1720 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5305_6
timestamp 1731220607
transform 1 0 1520 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5304_6
timestamp 1731220607
transform 1 0 1568 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5303_6
timestamp 1731220607
transform 1 0 1720 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5302_6
timestamp 1731220607
transform 1 0 1720 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5301_6
timestamp 1731220607
transform 1 0 1880 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5300_6
timestamp 1731220607
transform 1 0 1896 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5299_6
timestamp 1731220607
transform 1 0 1984 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5298_6
timestamp 1731220607
transform 1 0 2208 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5297_6
timestamp 1731220607
transform 1 0 2344 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5296_6
timestamp 1731220607
transform 1 0 2624 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5295_6
timestamp 1731220607
transform 1 0 2480 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5294_6
timestamp 1731220607
transform 1 0 2424 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5293_6
timestamp 1731220607
transform 1 0 2400 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5292_6
timestamp 1731220607
transform 1 0 2240 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5291_6
timestamp 1731220607
transform 1 0 2424 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5290_6
timestamp 1731220607
transform 1 0 2296 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5289_6
timestamp 1731220607
transform 1 0 2176 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5288_6
timestamp 1731220607
transform 1 0 2056 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5287_6
timestamp 1731220607
transform 1 0 2192 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5286_6
timestamp 1731220607
transform 1 0 2344 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5285_6
timestamp 1731220607
transform 1 0 2472 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5284_6
timestamp 1731220607
transform 1 0 2304 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5283_6
timestamp 1731220607
transform 1 0 2152 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5282_6
timestamp 1731220607
transform 1 0 2128 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5281_6
timestamp 1731220607
transform 1 0 1984 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5280_6
timestamp 1731220607
transform 1 0 2280 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5279_6
timestamp 1731220607
transform 1 0 2448 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5278_6
timestamp 1731220607
transform 1 0 2432 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5277_6
timestamp 1731220607
transform 1 0 2240 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5276_6
timestamp 1731220607
transform 1 0 2048 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5275_6
timestamp 1731220607
transform 1 0 2208 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5274_6
timestamp 1731220607
transform 1 0 2352 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5273_6
timestamp 1731220607
transform 1 0 2504 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5272_6
timestamp 1731220607
transform 1 0 2448 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5271_6
timestamp 1731220607
transform 1 0 2360 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5270_6
timestamp 1731220607
transform 1 0 2272 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5269_6
timestamp 1731220607
transform 1 0 2184 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5268_6
timestamp 1731220607
transform 1 0 2296 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5267_6
timestamp 1731220607
transform 1 0 2392 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5266_6
timestamp 1731220607
transform 1 0 2496 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5265_6
timestamp 1731220607
transform 1 0 2600 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5264_6
timestamp 1731220607
transform 1 0 2680 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5263_6
timestamp 1731220607
transform 1 0 2544 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5262_6
timestamp 1731220607
transform 1 0 2416 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5261_6
timestamp 1731220607
transform 1 0 2312 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5260_6
timestamp 1731220607
transform 1 0 2224 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5259_6
timestamp 1731220607
transform 1 0 2520 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5258_6
timestamp 1731220607
transform 1 0 2392 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5257_6
timestamp 1731220607
transform 1 0 2280 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5256_6
timestamp 1731220607
transform 1 0 2176 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5255_6
timestamp 1731220607
transform 1 0 2072 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5254_6
timestamp 1731220607
transform 1 0 2288 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5253_6
timestamp 1731220607
transform 1 0 2288 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5252_6
timestamp 1731220607
transform 1 0 2448 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5251_6
timestamp 1731220607
transform 1 0 2528 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5250_6
timestamp 1731220607
transform 1 0 2424 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5249_6
timestamp 1731220607
transform 1 0 2320 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5248_6
timestamp 1731220607
transform 1 0 2232 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5247_6
timestamp 1731220607
transform 1 0 2144 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5246_6
timestamp 1731220607
transform 1 0 2056 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5245_6
timestamp 1731220607
transform 1 0 1968 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5244_6
timestamp 1731220607
transform 1 0 1880 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5243_6
timestamp 1731220607
transform 1 0 2136 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5242_6
timestamp 1731220607
transform 1 0 1992 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5241_6
timestamp 1731220607
transform 1 0 1880 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5240_6
timestamp 1731220607
transform 1 0 1880 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5239_6
timestamp 1731220607
transform 1 0 1720 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5238_6
timestamp 1731220607
transform 1 0 1608 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5237_6
timestamp 1731220607
transform 1 0 1576 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5236_6
timestamp 1731220607
transform 1 0 1416 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5235_6
timestamp 1731220607
transform 1 0 1720 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5234_6
timestamp 1731220607
transform 1 0 1712 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5233_6
timestamp 1731220607
transform 1 0 1544 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5232_6
timestamp 1731220607
transform 1 0 1496 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5231_6
timestamp 1731220607
transform 1 0 1656 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5230_6
timestamp 1731220607
transform 1 0 1720 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5229_6
timestamp 1731220607
transform 1 0 1544 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5228_6
timestamp 1731220607
transform 1 0 1608 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5227_6
timestamp 1731220607
transform 1 0 1720 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5226_6
timestamp 1731220607
transform 1 0 1720 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5225_6
timestamp 1731220607
transform 1 0 1880 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5224_6
timestamp 1731220607
transform 1 0 1880 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5223_6
timestamp 1731220607
transform 1 0 1880 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5222_6
timestamp 1731220607
transform 1 0 2000 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5221_6
timestamp 1731220607
transform 1 0 2040 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5220_6
timestamp 1731220607
transform 1 0 1880 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5219_6
timestamp 1731220607
transform 1 0 1928 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5218_6
timestamp 1731220607
transform 1 0 1928 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5217_6
timestamp 1731220607
transform 1 0 2088 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5216_6
timestamp 1731220607
transform 1 0 2240 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5215_6
timestamp 1731220607
transform 1 0 2048 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5214_6
timestamp 1731220607
transform 1 0 2088 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5213_6
timestamp 1731220607
transform 1 0 2072 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5212_6
timestamp 1731220607
transform 1 0 2504 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5211_6
timestamp 1731220607
transform 1 0 2296 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5210_6
timestamp 1731220607
transform 1 0 2256 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5209_6
timestamp 1731220607
transform 1 0 2072 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5208_6
timestamp 1731220607
transform 1 0 2608 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5207_6
timestamp 1731220607
transform 1 0 2432 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5206_6
timestamp 1731220607
transform 1 0 2344 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5205_6
timestamp 1731220607
transform 1 0 2168 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5204_6
timestamp 1731220607
transform 1 0 2512 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5203_6
timestamp 1731220607
transform 1 0 2496 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5202_6
timestamp 1731220607
transform 1 0 2336 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5201_6
timestamp 1731220607
transform 1 0 2176 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5200_6
timestamp 1731220607
transform 1 0 2272 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5199_6
timestamp 1731220607
transform 1 0 2416 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5198_6
timestamp 1731220607
transform 1 0 2392 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5197_6
timestamp 1731220607
transform 1 0 2264 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5196_6
timestamp 1731220607
transform 1 0 2584 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5195_6
timestamp 1731220607
transform 1 0 2400 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5194_6
timestamp 1731220607
transform 1 0 2216 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5193_6
timestamp 1731220607
transform 1 0 2752 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5192_6
timestamp 1731220607
transform 1 0 2592 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5191_6
timestamp 1731220607
transform 1 0 2392 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5190_6
timestamp 1731220607
transform 1 0 2152 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5189_6
timestamp 1731220607
transform 1 0 2112 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5188_6
timestamp 1731220607
transform 1 0 1984 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5187_6
timestamp 1731220607
transform 1 0 2536 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5186_6
timestamp 1731220607
transform 1 0 2384 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5185_6
timestamp 1731220607
transform 1 0 2240 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5184_6
timestamp 1731220607
transform 1 0 2232 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5183_6
timestamp 1731220607
transform 1 0 2144 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5182_6
timestamp 1731220607
transform 1 0 2496 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5181_6
timestamp 1731220607
transform 1 0 2408 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5180_6
timestamp 1731220607
transform 1 0 2320 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5179_6
timestamp 1731220607
transform 1 0 2240 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5178_6
timestamp 1731220607
transform 1 0 2328 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5177_6
timestamp 1731220607
transform 1 0 2424 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5176_6
timestamp 1731220607
transform 1 0 2536 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5175_6
timestamp 1731220607
transform 1 0 2576 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5174_6
timestamp 1731220607
transform 1 0 2440 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5173_6
timestamp 1731220607
transform 1 0 2328 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5172_6
timestamp 1731220607
transform 1 0 2336 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5171_6
timestamp 1731220607
transform 1 0 2432 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5170_6
timestamp 1731220607
transform 1 0 2544 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5169_6
timestamp 1731220607
transform 1 0 2496 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5168_6
timestamp 1731220607
transform 1 0 2344 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5167_6
timestamp 1731220607
transform 1 0 2424 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5166_6
timestamp 1731220607
transform 1 0 2584 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5165_6
timestamp 1731220607
transform 1 0 2568 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5164_6
timestamp 1731220607
transform 1 0 2392 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5163_6
timestamp 1731220607
transform 1 0 2648 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5162_6
timestamp 1731220607
transform 1 0 2448 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5161_6
timestamp 1731220607
transform 1 0 2400 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5160_6
timestamp 1731220607
transform 1 0 2280 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5159_6
timestamp 1731220607
transform 1 0 2432 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5158_6
timestamp 1731220607
transform 1 0 2416 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5157_6
timestamp 1731220607
transform 1 0 2504 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5156_6
timestamp 1731220607
transform 1 0 2448 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5155_6
timestamp 1731220607
transform 1 0 2224 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5154_6
timestamp 1731220607
transform 1 0 2232 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5153_6
timestamp 1731220607
transform 1 0 2456 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5152_6
timestamp 1731220607
transform 1 0 2408 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5151_6
timestamp 1731220607
transform 1 0 2240 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5150_6
timestamp 1731220607
transform 1 0 2288 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5149_6
timestamp 1731220607
transform 1 0 2496 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5148_6
timestamp 1731220607
transform 1 0 2496 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5147_6
timestamp 1731220607
transform 1 0 2288 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5146_6
timestamp 1731220607
transform 1 0 2256 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5145_6
timestamp 1731220607
transform 1 0 2448 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5144_6
timestamp 1731220607
transform 1 0 2520 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5143_6
timestamp 1731220607
transform 1 0 2352 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5142_6
timestamp 1731220607
transform 1 0 2192 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5141_6
timestamp 1731220607
transform 1 0 2216 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5140_6
timestamp 1731220607
transform 1 0 2360 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5139_6
timestamp 1731220607
transform 1 0 2248 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5138_6
timestamp 1731220607
transform 1 0 2376 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5137_6
timestamp 1731220607
transform 1 0 2512 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5136_6
timestamp 1731220607
transform 1 0 2496 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5135_6
timestamp 1731220607
transform 1 0 2408 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5134_6
timestamp 1731220607
transform 1 0 2320 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5133_6
timestamp 1731220607
transform 1 0 2232 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5132_6
timestamp 1731220607
transform 1 0 2144 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5131_6
timestamp 1731220607
transform 1 0 2056 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5130_6
timestamp 1731220607
transform 1 0 1968 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5129_6
timestamp 1731220607
transform 1 0 1880 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5128_6
timestamp 1731220607
transform 1 0 1896 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5127_6
timestamp 1731220607
transform 1 0 2000 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5126_6
timestamp 1731220607
transform 1 0 2120 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5125_6
timestamp 1731220607
transform 1 0 2064 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5124_6
timestamp 1731220607
transform 1 0 1904 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5123_6
timestamp 1731220607
transform 1 0 1880 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5122_6
timestamp 1731220607
transform 1 0 2032 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5121_6
timestamp 1731220607
transform 1 0 2056 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5120_6
timestamp 1731220607
transform 1 0 1880 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5119_6
timestamp 1731220607
transform 1 0 1880 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5118_6
timestamp 1731220607
transform 1 0 2072 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5117_6
timestamp 1731220607
transform 1 0 2072 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5116_6
timestamp 1731220607
transform 1 0 1880 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5115_6
timestamp 1731220607
transform 1 0 1720 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5114_6
timestamp 1731220607
transform 1 0 1632 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5113_6
timestamp 1731220607
transform 1 0 1624 0 -1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5112_6
timestamp 1731220607
transform 1 0 1720 0 -1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5111_6
timestamp 1731220607
transform 1 0 1688 0 1 2856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5110_6
timestamp 1731220607
transform 1 0 1616 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5109_6
timestamp 1731220607
transform 1 0 1496 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5108_6
timestamp 1731220607
transform 1 0 1720 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5107_6
timestamp 1731220607
transform 1 0 1720 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5106_6
timestamp 1731220607
transform 1 0 1632 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5105_6
timestamp 1731220607
transform 1 0 1520 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5104_6
timestamp 1731220607
transform 1 0 1416 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5103_6
timestamp 1731220607
transform 1 0 1304 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5102_6
timestamp 1731220607
transform 1 0 1192 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5101_6
timestamp 1731220607
transform 1 0 1072 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5100_6
timestamp 1731220607
transform 1 0 944 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_599_6
timestamp 1731220607
transform 1 0 1128 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_598_6
timestamp 1731220607
transform 1 0 1256 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_597_6
timestamp 1731220607
transform 1 0 1376 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_596_6
timestamp 1731220607
transform 1 0 1344 0 1 2856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_595_6
timestamp 1731220607
transform 1 0 1568 0 1 2856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_594_6
timestamp 1731220607
transform 1 0 1456 0 1 2856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_593_6
timestamp 1731220607
transform 1 0 1400 0 -1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_592_6
timestamp 1731220607
transform 1 0 1512 0 -1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_591_6
timestamp 1731220607
transform 1 0 1456 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_590_6
timestamp 1731220607
transform 1 0 1544 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_589_6
timestamp 1731220607
transform 1 0 1512 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_588_6
timestamp 1731220607
transform 1 0 1368 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_587_6
timestamp 1731220607
transform 1 0 1368 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_586_6
timestamp 1731220607
transform 1 0 1520 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_585_6
timestamp 1731220607
transform 1 0 1512 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_584_6
timestamp 1731220607
transform 1 0 1336 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_583_6
timestamp 1731220607
transform 1 0 1264 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_582_6
timestamp 1731220607
transform 1 0 1400 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_581_6
timestamp 1731220607
transform 1 0 1544 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_580_6
timestamp 1731220607
transform 1 0 1472 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_579_6
timestamp 1731220607
transform 1 0 1288 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_578_6
timestamp 1731220607
transform 1 0 1560 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_577_6
timestamp 1731220607
transform 1 0 1440 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_576_6
timestamp 1731220607
transform 1 0 1320 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_575_6
timestamp 1731220607
transform 1 0 1200 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_574_6
timestamp 1731220607
transform 1 0 1536 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_573_6
timestamp 1731220607
transform 1 0 1416 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_572_6
timestamp 1731220607
transform 1 0 1304 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_571_6
timestamp 1731220607
transform 1 0 1192 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_570_6
timestamp 1731220607
transform 1 0 1072 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_569_6
timestamp 1731220607
transform 1 0 944 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_568_6
timestamp 1731220607
transform 1 0 816 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_567_6
timestamp 1731220607
transform 1 0 816 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_566_6
timestamp 1731220607
transform 1 0 1080 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_565_6
timestamp 1731220607
transform 1 0 952 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_564_6
timestamp 1731220607
transform 1 0 928 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_563_6
timestamp 1731220607
transform 1 0 1104 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_562_6
timestamp 1731220607
transform 1 0 1128 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_561_6
timestamp 1731220607
transform 1 0 984 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_560_6
timestamp 1731220607
transform 1 0 840 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_559_6
timestamp 1731220607
transform 1 0 984 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_558_6
timestamp 1731220607
transform 1 0 1160 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_557_6
timestamp 1731220607
transform 1 0 1216 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_556_6
timestamp 1731220607
transform 1 0 1064 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_555_6
timestamp 1731220607
transform 1 0 920 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_554_6
timestamp 1731220607
transform 1 0 1088 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_553_6
timestamp 1731220607
transform 1 0 1224 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_552_6
timestamp 1731220607
transform 1 0 1368 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_551_6
timestamp 1731220607
transform 1 0 1280 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_550_6
timestamp 1731220607
transform 1 0 1192 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_549_6
timestamp 1731220607
transform 1 0 1104 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_548_6
timestamp 1731220607
transform 1 0 1016 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_547_6
timestamp 1731220607
transform 1 0 928 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_546_6
timestamp 1731220607
transform 1 0 840 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_545_6
timestamp 1731220607
transform 1 0 752 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_544_6
timestamp 1731220607
transform 1 0 664 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_543_6
timestamp 1731220607
transform 1 0 576 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_542_6
timestamp 1731220607
transform 1 0 488 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_541_6
timestamp 1731220607
transform 1 0 400 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_540_6
timestamp 1731220607
transform 1 0 312 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_539_6
timestamp 1731220607
transform 1 0 224 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_538_6
timestamp 1731220607
transform 1 0 136 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_537_6
timestamp 1731220607
transform 1 0 960 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_536_6
timestamp 1731220607
transform 1 0 840 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_535_6
timestamp 1731220607
transform 1 0 728 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_534_6
timestamp 1731220607
transform 1 0 632 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_533_6
timestamp 1731220607
transform 1 0 544 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_532_6
timestamp 1731220607
transform 1 0 456 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_531_6
timestamp 1731220607
transform 1 0 784 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_530_6
timestamp 1731220607
transform 1 0 656 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_529_6
timestamp 1731220607
transform 1 0 536 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_528_6
timestamp 1731220607
transform 1 0 416 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_527_6
timestamp 1731220607
transform 1 0 816 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_526_6
timestamp 1731220607
transform 1 0 656 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_525_6
timestamp 1731220607
transform 1 0 504 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_524_6
timestamp 1731220607
transform 1 0 368 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_523_6
timestamp 1731220607
transform 1 0 248 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_522_6
timestamp 1731220607
transform 1 0 680 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_521_6
timestamp 1731220607
transform 1 0 520 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_520_6
timestamp 1731220607
transform 1 0 352 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_519_6
timestamp 1731220607
transform 1 0 192 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_518_6
timestamp 1731220607
transform 1 0 752 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_517_6
timestamp 1731220607
transform 1 0 576 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_516_6
timestamp 1731220607
transform 1 0 408 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_515_6
timestamp 1731220607
transform 1 0 248 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_514_6
timestamp 1731220607
transform 1 0 128 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_513_6
timestamp 1731220607
transform 1 0 168 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_512_6
timestamp 1731220607
transform 1 0 336 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_511_6
timestamp 1731220607
transform 1 0 504 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_510_6
timestamp 1731220607
transform 1 0 664 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_59_6
timestamp 1731220607
transform 1 0 680 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_58_6
timestamp 1731220607
transform 1 0 536 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_57_6
timestamp 1731220607
transform 1 0 392 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_56_6
timestamp 1731220607
transform 1 0 240 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_55_6
timestamp 1731220607
transform 1 0 224 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_54_6
timestamp 1731220607
transform 1 0 312 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_53_6
timestamp 1731220607
transform 1 0 400 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_52_6
timestamp 1731220607
transform 1 0 488 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_51_6
timestamp 1731220607
transform 1 0 576 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_50_6
timestamp 1731220607
transform 1 0 664 0 1 3580
box 8 4 80 64
<< end >>
