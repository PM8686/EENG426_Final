magic
tech sky130l
timestamp 1731220477
<< m1 >>
rect 400 5699 404 5731
rect 2152 5631 2156 5663
rect 2368 5631 2372 5663
rect 2536 5631 2540 5663
rect 4600 5635 4604 5667
rect 4736 5635 4740 5667
rect 4872 5635 4876 5667
rect 1392 5511 1396 5527
rect 1008 5475 1012 5507
rect 1536 5511 1540 5587
rect 1576 5559 1580 5587
rect 1752 5559 1756 5587
rect 1144 5475 1148 5507
rect 4576 5411 4580 5443
rect 4896 5411 4900 5443
rect 5040 5411 5044 5443
rect 824 5335 828 5363
rect 960 5335 964 5363
rect 1096 5335 1100 5363
rect 1488 5251 1492 5283
rect 3304 5175 3308 5207
rect 4720 5199 4724 5291
rect 5120 5263 5124 5291
rect 4744 5163 4748 5195
rect 4904 5163 4908 5195
rect 5048 5163 5052 5195
rect 5200 5163 5204 5195
rect 5368 5163 5372 5195
rect 5512 5163 5516 5195
rect 944 5111 948 5139
rect 2472 5019 2476 5047
rect 1952 4963 1956 5015
rect 3320 4963 3324 5047
rect 2128 4927 2132 4959
rect 2264 4927 2268 4959
rect 4264 4931 4268 4963
rect 4400 4931 4404 4963
rect 4536 4931 4540 4963
rect 4672 4931 4676 4963
rect 4944 4931 4948 4963
rect 5080 4931 5084 4963
rect 5512 4931 5516 4963
rect 264 4851 268 4879
rect 3312 4779 3316 4807
rect 4672 4631 4676 4663
rect 4808 4631 4812 4663
rect 4960 4631 4964 4663
rect 5104 4631 5108 4663
rect 5240 4631 5244 4663
rect 5512 4631 5516 4663
rect 1704 4515 1708 4547
rect 4480 4403 4484 4435
rect 4616 4403 4620 4435
rect 4752 4403 4756 4435
rect 4888 4403 4892 4435
rect 848 4287 852 4319
rect 984 4287 988 4319
rect 1120 4287 1124 4319
rect 1256 4287 1260 4319
rect 2152 4291 2156 4319
rect 2376 4203 2380 4235
rect 3280 4203 3284 4235
rect 1104 4139 1108 4167
rect 1240 4139 1244 4167
rect 4104 4151 4108 4183
rect 4376 4151 4380 4183
rect 4512 4151 4516 4183
rect 696 4055 700 4087
rect 832 4055 836 4087
rect 1104 4055 1108 4087
rect 1376 4055 1380 4087
rect 1648 4055 1652 4087
rect 1784 4055 1788 4079
rect 3512 4051 3516 4079
rect 3648 4051 3652 4079
rect 4264 3939 4268 4007
rect 1448 3711 1452 3863
rect 2136 3679 2140 3747
rect 2144 3643 2148 3675
rect 3152 3643 3156 3675
rect 4968 3631 4972 3663
rect 5104 3631 5108 3663
rect 5240 3631 5244 3663
rect 5376 3631 5380 3663
rect 5512 3631 5516 3663
rect 632 3579 636 3611
rect 3024 3495 3028 3523
rect 456 3327 460 3359
rect 864 3327 868 3359
rect 4096 3351 4100 3383
rect 5200 3351 5204 3383
rect 3088 3195 3092 3263
rect 320 3079 324 3111
rect 3200 2971 3204 3039
rect 2936 2935 2940 2967
rect 3208 2935 3212 2967
rect 3344 2935 3348 2967
rect 3480 2935 3484 2967
rect 528 2851 532 2883
rect 1304 2851 1308 2935
rect 1480 2851 1484 2883
rect 1632 2851 1636 2883
rect 1784 2851 1788 2883
rect 2136 2743 2140 2771
rect 2272 2743 2276 2771
rect 2456 2743 2460 2771
rect 776 2699 780 2727
rect 936 2699 940 2727
rect 2512 2659 2516 2691
rect 904 2615 908 2647
rect 1176 2615 1180 2647
rect 1312 2615 1316 2647
rect 1584 2615 1588 2647
rect 1720 2615 1724 2647
rect 2616 2515 2620 2543
rect 2752 2515 2756 2543
rect 1584 2459 1588 2487
rect 4968 2379 4972 2411
rect 5104 2379 5108 2411
rect 5240 2379 5244 2411
rect 288 2219 292 2287
rect 2288 2183 2292 2215
rect 872 2111 876 2143
rect 4128 2139 4132 2171
rect 4264 2139 4268 2171
rect 4400 2139 4404 2171
rect 5232 2139 5236 2171
rect 1216 1967 1220 1995
rect 1360 1967 1364 1995
rect 3992 1979 3996 2007
rect 4128 1979 4132 2007
rect 4264 1979 4268 2007
rect 4400 1979 4404 2007
rect 4536 1943 4540 2007
rect 5032 1979 5036 2007
rect 5224 1979 5228 2007
rect 3512 1843 3516 1871
rect 3648 1843 3652 1871
rect 2128 1747 2132 1779
rect 2264 1747 2268 1779
rect 2416 1747 2420 1779
rect 2568 1747 2572 1779
rect 3032 1747 3036 1779
rect 3648 1747 3652 1779
rect 384 1719 388 1747
rect 4696 1655 4700 1687
rect 4832 1655 4836 1679
rect 816 1623 820 1655
rect 3216 1535 3220 1623
rect 2128 1499 2132 1531
rect 2264 1499 2268 1523
rect 2808 1499 2812 1531
rect 2944 1499 2948 1531
rect 3080 1499 3084 1531
rect 3352 1499 3356 1531
rect 5328 1531 5332 1671
rect 3488 1499 3492 1531
rect 5480 1379 5484 1519
rect 2272 1347 2276 1375
rect 4944 1343 4948 1375
rect 5080 1343 5084 1375
rect 5476 1375 5484 1379
rect 5216 1343 5220 1375
rect 2400 1263 2404 1295
rect 3024 1263 3028 1295
rect 3264 1263 3268 1295
rect 1200 1163 1204 1263
rect 992 1127 996 1159
rect 1192 1127 1196 1159
rect 392 987 396 1015
rect 1240 899 1244 983
rect 1392 899 1396 931
rect 1776 899 1780 931
rect 1968 879 1972 931
rect 5376 883 5380 915
rect 584 659 588 675
rect 1320 659 1324 691
rect 1472 659 1476 691
rect 1640 659 1644 691
rect 1784 659 1788 691
rect 4504 687 4508 771
rect 4128 651 4132 683
rect 4264 651 4268 683
rect 4400 651 4404 683
rect 760 519 764 547
rect 944 519 948 547
rect 1632 519 1636 547
rect 4128 511 4132 539
rect 4408 511 4412 607
rect 1960 407 1964 467
rect 2144 407 2148 439
rect 832 279 836 307
rect 992 279 996 307
rect 5368 303 5372 435
rect 2696 243 2700 271
rect 280 163 284 195
rect 416 163 420 195
rect 552 163 556 195
rect 688 163 692 195
rect 960 163 964 195
rect 1096 163 1100 195
rect 4416 183 4420 299
rect 2128 143 2132 175
rect 2264 143 2268 175
rect 2400 143 2404 175
rect 2672 143 2676 175
rect 2808 143 2812 175
rect 3080 143 3084 175
rect 3216 143 3220 175
rect 3488 143 3492 175
rect 3624 143 3628 175
rect 4424 147 4428 179
rect 4560 147 4564 179
rect 4696 147 4700 179
rect 4968 147 4972 179
rect 5104 147 5108 179
rect 5240 147 5244 179
<< m2c >>
rect 400 5731 404 5735
rect 256 5695 260 5699
rect 392 5695 396 5699
rect 400 5695 404 5699
rect 528 5695 532 5699
rect 4600 5667 4604 5671
rect 2152 5663 2156 5667
rect 2368 5663 2372 5667
rect 2536 5663 2540 5667
rect 4736 5667 4740 5671
rect 4872 5667 4876 5671
rect 4592 5631 4596 5635
rect 4600 5631 4604 5635
rect 4728 5631 4732 5635
rect 4736 5631 4740 5635
rect 4864 5631 4868 5635
rect 4872 5631 4876 5635
rect 5000 5631 5004 5635
rect 2120 5627 2124 5631
rect 2152 5627 2156 5631
rect 2296 5627 2300 5631
rect 2368 5627 2372 5631
rect 2496 5627 2500 5631
rect 2536 5627 2540 5631
rect 2688 5627 2692 5631
rect 2872 5627 2876 5631
rect 3056 5627 3060 5631
rect 3232 5627 3236 5631
rect 3400 5627 3404 5631
rect 3568 5627 3572 5631
rect 3744 5627 3748 5631
rect 440 5587 444 5591
rect 632 5587 636 5591
rect 832 5587 836 5591
rect 1040 5587 1044 5591
rect 1256 5587 1260 5591
rect 1480 5587 1484 5591
rect 1536 5587 1540 5591
rect 1392 5527 1396 5531
rect 1008 5507 1012 5511
rect 1144 5507 1148 5511
rect 1392 5507 1396 5511
rect 1576 5587 1580 5591
rect 1704 5587 1708 5591
rect 1752 5587 1756 5591
rect 1912 5587 1916 5591
rect 1576 5555 1580 5559
rect 1752 5555 1756 5559
rect 4528 5523 4532 5527
rect 4664 5523 4668 5527
rect 4800 5523 4804 5527
rect 4936 5523 4940 5527
rect 5072 5523 5076 5527
rect 5208 5523 5212 5527
rect 2472 5519 2476 5523
rect 2704 5519 2708 5523
rect 2928 5519 2932 5523
rect 3144 5519 3148 5523
rect 3360 5519 3364 5523
rect 3576 5519 3580 5523
rect 3776 5519 3780 5523
rect 1536 5507 1540 5511
rect 1000 5471 1004 5475
rect 1008 5471 1012 5475
rect 1136 5471 1140 5475
rect 1144 5471 1148 5475
rect 1272 5471 1276 5475
rect 1416 5471 1420 5475
rect 1560 5471 1564 5475
rect 1704 5471 1708 5475
rect 1848 5471 1852 5475
rect 4576 5443 4580 5447
rect 4896 5443 4900 5447
rect 5040 5443 5044 5447
rect 4552 5407 4556 5411
rect 4576 5407 4580 5411
rect 4712 5407 4716 5411
rect 4872 5407 4876 5411
rect 4896 5407 4900 5411
rect 5032 5407 5036 5411
rect 5040 5407 5044 5411
rect 5200 5407 5204 5411
rect 2576 5399 2580 5403
rect 2824 5399 2828 5403
rect 3072 5399 3076 5403
rect 3312 5399 3316 5403
rect 3552 5399 3556 5403
rect 3776 5399 3780 5403
rect 816 5363 820 5367
rect 824 5363 828 5367
rect 952 5363 956 5367
rect 960 5363 964 5367
rect 1088 5363 1092 5367
rect 1096 5363 1100 5367
rect 1224 5363 1228 5367
rect 1360 5363 1364 5367
rect 1496 5363 1500 5367
rect 1632 5363 1636 5367
rect 1768 5363 1772 5367
rect 1904 5363 1908 5367
rect 824 5331 828 5335
rect 960 5331 964 5335
rect 1096 5331 1100 5335
rect 2416 5291 2420 5295
rect 2616 5291 2620 5295
rect 2816 5291 2820 5295
rect 3016 5291 3020 5295
rect 3216 5291 3220 5295
rect 3424 5291 3428 5295
rect 3632 5291 3636 5295
rect 4528 5291 4532 5295
rect 4712 5291 4716 5295
rect 4720 5291 4724 5295
rect 4896 5291 4900 5295
rect 5080 5291 5084 5295
rect 5120 5291 5124 5295
rect 5272 5291 5276 5295
rect 1488 5283 1492 5287
rect 848 5247 852 5251
rect 1000 5247 1004 5251
rect 1152 5247 1156 5251
rect 1312 5247 1316 5251
rect 1480 5247 1484 5251
rect 1488 5247 1492 5251
rect 1648 5247 1652 5251
rect 3304 5207 3308 5211
rect 5120 5259 5124 5263
rect 4720 5195 4724 5199
rect 4744 5195 4748 5199
rect 2400 5171 2404 5175
rect 2600 5171 2604 5175
rect 2808 5171 2812 5175
rect 3016 5171 3020 5175
rect 3224 5171 3228 5175
rect 3304 5171 3308 5175
rect 3432 5171 3436 5175
rect 4904 5195 4908 5199
rect 5048 5195 5052 5199
rect 5200 5195 5204 5199
rect 5368 5195 5372 5199
rect 5512 5195 5516 5199
rect 4560 5159 4564 5163
rect 4720 5159 4724 5163
rect 4744 5159 4748 5163
rect 4880 5159 4884 5163
rect 4904 5159 4908 5163
rect 5040 5159 5044 5163
rect 5048 5159 5052 5163
rect 5192 5159 5196 5163
rect 5200 5159 5204 5163
rect 5344 5159 5348 5163
rect 5368 5159 5372 5163
rect 5504 5159 5508 5163
rect 5512 5159 5516 5163
rect 5640 5159 5644 5163
rect 544 5139 548 5143
rect 720 5139 724 5143
rect 904 5139 908 5143
rect 944 5139 948 5143
rect 1096 5139 1100 5143
rect 1296 5139 1300 5143
rect 1496 5139 1500 5143
rect 1704 5139 1708 5143
rect 1912 5139 1916 5143
rect 944 5107 948 5111
rect 2216 5047 2220 5051
rect 2424 5047 2428 5051
rect 2472 5047 2476 5051
rect 2632 5047 2636 5051
rect 2848 5047 2852 5051
rect 3072 5047 3076 5051
rect 3304 5047 3308 5051
rect 3320 5047 3324 5051
rect 280 5015 284 5019
rect 504 5015 508 5019
rect 752 5015 756 5019
rect 1024 5015 1028 5019
rect 1320 5015 1324 5019
rect 1624 5015 1628 5019
rect 1912 5015 1916 5019
rect 1952 5015 1956 5019
rect 2472 5015 2476 5019
rect 3984 5043 3988 5047
rect 4184 5043 4188 5047
rect 4424 5043 4428 5047
rect 4664 5043 4668 5047
rect 4912 5043 4916 5047
rect 5160 5043 5164 5047
rect 5408 5043 5412 5047
rect 5640 5043 5644 5047
rect 1952 4959 1956 4963
rect 2128 4959 2132 4963
rect 2264 4959 2268 4963
rect 3320 4959 3324 4963
rect 4264 4963 4268 4967
rect 4400 4963 4404 4967
rect 4536 4963 4540 4967
rect 4672 4963 4676 4967
rect 4944 4963 4948 4967
rect 5080 4963 5084 4967
rect 5512 4963 5516 4967
rect 3984 4927 3988 4931
rect 4120 4927 4124 4931
rect 4256 4927 4260 4931
rect 4264 4927 4268 4931
rect 4392 4927 4396 4931
rect 4400 4927 4404 4931
rect 4528 4927 4532 4931
rect 4536 4927 4540 4931
rect 4664 4927 4668 4931
rect 4672 4927 4676 4931
rect 4800 4927 4804 4931
rect 4936 4927 4940 4931
rect 4944 4927 4948 4931
rect 5072 4927 5076 4931
rect 5080 4927 5084 4931
rect 5208 4927 5212 4931
rect 5352 4927 5356 4931
rect 5504 4927 5508 4931
rect 5512 4927 5516 4931
rect 5640 4927 5644 4931
rect 2120 4923 2124 4927
rect 2128 4923 2132 4927
rect 2256 4923 2260 4927
rect 2264 4923 2268 4927
rect 2392 4923 2396 4927
rect 2544 4923 2548 4927
rect 2744 4923 2748 4927
rect 2984 4923 2988 4927
rect 3248 4923 3252 4927
rect 3520 4923 3524 4927
rect 3776 4923 3780 4927
rect 256 4879 260 4883
rect 264 4879 268 4883
rect 392 4879 396 4883
rect 528 4879 532 4883
rect 664 4879 668 4883
rect 800 4879 804 4883
rect 264 4847 268 4851
rect 2424 4807 2428 4811
rect 2656 4807 2660 4811
rect 2920 4807 2924 4811
rect 3200 4807 3204 4811
rect 3312 4807 3316 4811
rect 3496 4807 3500 4811
rect 3776 4807 3780 4811
rect 3312 4775 3316 4779
rect 256 4751 260 4755
rect 392 4751 396 4755
rect 528 4751 532 4755
rect 664 4751 668 4755
rect 800 4751 804 4755
rect 3984 4743 3988 4747
rect 4168 4743 4172 4747
rect 4392 4743 4396 4747
rect 4632 4743 4636 4747
rect 4880 4743 4884 4747
rect 5136 4743 5140 4747
rect 5400 4743 5404 4747
rect 5640 4743 5644 4747
rect 2144 4679 2148 4683
rect 2320 4679 2324 4683
rect 2496 4679 2500 4683
rect 2672 4679 2676 4683
rect 2848 4679 2852 4683
rect 4672 4663 4676 4667
rect 256 4639 260 4643
rect 392 4639 396 4643
rect 528 4639 532 4643
rect 664 4639 668 4643
rect 800 4639 804 4643
rect 4808 4663 4812 4667
rect 4960 4663 4964 4667
rect 5104 4663 5108 4667
rect 5240 4663 5244 4667
rect 5512 4663 5516 4667
rect 3984 4627 3988 4631
rect 4120 4627 4124 4631
rect 4256 4627 4260 4631
rect 4392 4627 4396 4631
rect 4528 4627 4532 4631
rect 4664 4627 4668 4631
rect 4672 4627 4676 4631
rect 4800 4627 4804 4631
rect 4808 4627 4812 4631
rect 4944 4627 4948 4631
rect 4960 4627 4964 4631
rect 5088 4627 5092 4631
rect 5104 4627 5108 4631
rect 5232 4627 5236 4631
rect 5240 4627 5244 4631
rect 5368 4627 5372 4631
rect 5504 4627 5508 4631
rect 5512 4627 5516 4631
rect 5640 4627 5644 4631
rect 2120 4567 2124 4571
rect 2360 4567 2364 4571
rect 2624 4567 2628 4571
rect 2872 4567 2876 4571
rect 3112 4567 3116 4571
rect 3344 4567 3348 4571
rect 3568 4567 3572 4571
rect 3776 4567 3780 4571
rect 1704 4547 1708 4551
rect 4768 4519 4772 4523
rect 4904 4519 4908 4523
rect 5040 4519 5044 4523
rect 5176 4519 5180 4523
rect 376 4511 380 4515
rect 568 4511 572 4515
rect 776 4511 780 4515
rect 1000 4511 1004 4515
rect 1224 4511 1228 4515
rect 1456 4511 1460 4515
rect 1696 4511 1700 4515
rect 1704 4511 1708 4515
rect 1912 4511 1916 4515
rect 2392 4439 2396 4443
rect 2640 4439 2644 4443
rect 2872 4439 2876 4443
rect 3096 4439 3100 4443
rect 3312 4439 3316 4443
rect 3520 4439 3524 4443
rect 3736 4439 3740 4443
rect 4480 4435 4484 4439
rect 608 4403 612 4407
rect 784 4403 788 4407
rect 968 4403 972 4407
rect 1168 4403 1172 4407
rect 1376 4403 1380 4407
rect 1592 4403 1596 4407
rect 1816 4403 1820 4407
rect 4616 4435 4620 4439
rect 4752 4435 4756 4439
rect 4888 4435 4892 4439
rect 4472 4399 4476 4403
rect 4480 4399 4484 4403
rect 4608 4399 4612 4403
rect 4616 4399 4620 4403
rect 4744 4399 4748 4403
rect 4752 4399 4756 4403
rect 4880 4399 4884 4403
rect 4888 4399 4892 4403
rect 5016 4399 5020 4403
rect 848 4319 852 4323
rect 984 4319 988 4323
rect 1120 4319 1124 4323
rect 1256 4319 1260 4323
rect 2120 4319 2124 4323
rect 2152 4319 2156 4323
rect 2296 4319 2300 4323
rect 2496 4319 2500 4323
rect 2688 4319 2692 4323
rect 2872 4319 2876 4323
rect 3048 4319 3052 4323
rect 3232 4319 3236 4323
rect 3416 4319 3420 4323
rect 2152 4287 2156 4291
rect 840 4283 844 4287
rect 848 4283 852 4287
rect 976 4283 980 4287
rect 984 4283 988 4287
rect 1112 4283 1116 4287
rect 1120 4283 1124 4287
rect 1248 4283 1252 4287
rect 1256 4283 1260 4287
rect 1384 4283 1388 4287
rect 1520 4283 1524 4287
rect 1656 4283 1660 4287
rect 1792 4283 1796 4287
rect 4232 4275 4236 4279
rect 4368 4275 4372 4279
rect 4504 4275 4508 4279
rect 4640 4275 4644 4279
rect 4776 4275 4780 4279
rect 2376 4235 2380 4239
rect 3280 4235 3284 4239
rect 2120 4199 2124 4203
rect 2368 4199 2372 4203
rect 2376 4199 2380 4203
rect 2632 4199 2636 4203
rect 2888 4199 2892 4203
rect 3144 4199 3148 4203
rect 3280 4199 3284 4203
rect 3408 4199 3412 4203
rect 4104 4183 4108 4187
rect 824 4167 828 4171
rect 960 4167 964 4171
rect 1096 4167 1100 4171
rect 1104 4167 1108 4171
rect 1232 4167 1236 4171
rect 1240 4167 1244 4171
rect 1368 4167 1372 4171
rect 1504 4167 1508 4171
rect 1640 4167 1644 4171
rect 1776 4167 1780 4171
rect 1912 4167 1916 4171
rect 1104 4135 1108 4139
rect 4376 4183 4380 4187
rect 4512 4183 4516 4187
rect 4096 4147 4100 4151
rect 4104 4147 4108 4151
rect 4232 4147 4236 4151
rect 4368 4147 4372 4151
rect 4376 4147 4380 4151
rect 4504 4147 4508 4151
rect 4512 4147 4516 4151
rect 4640 4147 4644 4151
rect 1240 4135 1244 4139
rect 696 4087 700 4091
rect 832 4087 836 4091
rect 1104 4087 1108 4091
rect 1376 4087 1380 4091
rect 1648 4087 1652 4091
rect 1784 4079 1788 4083
rect 3232 4079 3236 4083
rect 3368 4079 3372 4083
rect 3504 4079 3508 4083
rect 3512 4079 3516 4083
rect 3640 4079 3644 4083
rect 3648 4079 3652 4083
rect 3776 4079 3780 4083
rect 688 4051 692 4055
rect 696 4051 700 4055
rect 824 4051 828 4055
rect 832 4051 836 4055
rect 960 4051 964 4055
rect 1096 4051 1100 4055
rect 1104 4051 1108 4055
rect 1232 4051 1236 4055
rect 1368 4051 1372 4055
rect 1376 4051 1380 4055
rect 1504 4051 1508 4055
rect 1640 4051 1644 4055
rect 1648 4051 1652 4055
rect 1776 4051 1780 4055
rect 1784 4051 1788 4055
rect 1912 4051 1916 4055
rect 3512 4047 3516 4051
rect 3648 4047 3652 4051
rect 3984 4015 3988 4019
rect 4120 4015 4124 4019
rect 4256 4015 4260 4019
rect 4392 4015 4396 4019
rect 4528 4015 4532 4019
rect 4664 4015 4668 4019
rect 4800 4015 4804 4019
rect 4936 4015 4940 4019
rect 4264 4007 4268 4011
rect 256 3943 260 3947
rect 424 3943 428 3947
rect 632 3943 636 3947
rect 848 3943 852 3947
rect 1064 3943 1068 3947
rect 1280 3943 1284 3947
rect 1496 3943 1500 3947
rect 1712 3943 1716 3947
rect 1912 3943 1916 3947
rect 4264 3935 4268 3939
rect 3984 3899 3988 3903
rect 4120 3899 4124 3903
rect 4272 3899 4276 3903
rect 4424 3899 4428 3903
rect 4584 3899 4588 3903
rect 4744 3899 4748 3903
rect 4904 3899 4908 3903
rect 2120 3871 2124 3875
rect 2528 3871 2532 3875
rect 2952 3871 2956 3875
rect 3376 3871 3380 3875
rect 3776 3871 3780 3875
rect 1448 3863 1452 3867
rect 256 3827 260 3831
rect 480 3827 484 3831
rect 744 3827 748 3831
rect 1024 3827 1028 3831
rect 1320 3827 1324 3831
rect 1624 3827 1628 3831
rect 1912 3827 1916 3831
rect 2120 3763 2124 3767
rect 2272 3763 2276 3767
rect 2448 3763 2452 3767
rect 2632 3763 2636 3767
rect 2816 3763 2820 3767
rect 2992 3763 2996 3767
rect 3168 3763 3172 3767
rect 3344 3763 3348 3767
rect 3520 3763 3524 3767
rect 3704 3763 3708 3767
rect 4600 3763 4604 3767
rect 4736 3763 4740 3767
rect 4872 3763 4876 3767
rect 5008 3763 5012 3767
rect 5144 3763 5148 3767
rect 344 3707 348 3711
rect 616 3707 620 3711
rect 888 3707 892 3711
rect 1160 3707 1164 3711
rect 1440 3707 1444 3711
rect 1448 3707 1452 3711
rect 2136 3747 2140 3751
rect 2136 3675 2140 3679
rect 2144 3675 2148 3679
rect 3152 3675 3156 3679
rect 4968 3663 4972 3667
rect 2136 3639 2140 3643
rect 2144 3639 2148 3643
rect 2272 3639 2276 3643
rect 2416 3639 2420 3643
rect 2560 3639 2564 3643
rect 2704 3639 2708 3643
rect 2848 3639 2852 3643
rect 2992 3639 2996 3643
rect 3136 3639 3140 3643
rect 3152 3639 3156 3643
rect 3280 3639 3284 3643
rect 3424 3639 3428 3643
rect 5104 3663 5108 3667
rect 5240 3663 5244 3667
rect 5376 3663 5380 3667
rect 5512 3663 5516 3667
rect 4144 3627 4148 3631
rect 4280 3627 4284 3631
rect 4416 3627 4420 3631
rect 4552 3627 4556 3631
rect 4688 3627 4692 3631
rect 4824 3627 4828 3631
rect 4960 3627 4964 3631
rect 4968 3627 4972 3631
rect 5096 3627 5100 3631
rect 5104 3627 5108 3631
rect 5232 3627 5236 3631
rect 5240 3627 5244 3631
rect 5368 3627 5372 3631
rect 5376 3627 5380 3631
rect 5504 3627 5508 3631
rect 5512 3627 5516 3631
rect 5640 3627 5644 3631
rect 632 3611 636 3615
rect 616 3575 620 3579
rect 632 3575 636 3579
rect 760 3575 764 3579
rect 904 3575 908 3579
rect 1048 3575 1052 3579
rect 1192 3575 1196 3579
rect 1336 3575 1340 3579
rect 2336 3523 2340 3527
rect 2472 3523 2476 3527
rect 2608 3523 2612 3527
rect 2744 3523 2748 3527
rect 2880 3523 2884 3527
rect 3016 3523 3020 3527
rect 3024 3523 3028 3527
rect 3152 3523 3156 3527
rect 3288 3523 3292 3527
rect 3424 3523 3428 3527
rect 3560 3523 3564 3527
rect 3024 3491 3028 3495
rect 5504 3471 5508 3475
rect 5640 3471 5644 3475
rect 528 3447 532 3451
rect 664 3447 668 3451
rect 800 3447 804 3451
rect 936 3447 940 3451
rect 1072 3447 1076 3451
rect 2296 3403 2300 3407
rect 2472 3403 2476 3407
rect 2656 3403 2660 3407
rect 2840 3403 2844 3407
rect 3032 3403 3036 3407
rect 3224 3403 3228 3407
rect 3416 3403 3420 3407
rect 3608 3403 3612 3407
rect 3776 3403 3780 3407
rect 4096 3383 4100 3387
rect 456 3359 460 3363
rect 864 3359 868 3363
rect 5200 3383 5204 3387
rect 3984 3347 3988 3351
rect 4096 3347 4100 3351
rect 4224 3347 4228 3351
rect 4472 3347 4476 3351
rect 4712 3347 4716 3351
rect 4936 3347 4940 3351
rect 5152 3347 5156 3351
rect 5200 3347 5204 3351
rect 5360 3347 5364 3351
rect 5576 3347 5580 3351
rect 448 3323 452 3327
rect 456 3323 460 3327
rect 584 3323 588 3327
rect 720 3323 724 3327
rect 856 3323 860 3327
rect 864 3323 868 3327
rect 992 3323 996 3327
rect 2248 3271 2252 3275
rect 2496 3271 2500 3275
rect 2784 3271 2788 3275
rect 3112 3271 3116 3275
rect 3456 3271 3460 3275
rect 3776 3271 3780 3275
rect 3088 3263 3092 3267
rect 256 3207 260 3211
rect 432 3207 436 3211
rect 640 3207 644 3211
rect 848 3207 852 3211
rect 1056 3207 1060 3211
rect 3984 3239 3988 3243
rect 4224 3239 4228 3243
rect 4472 3239 4476 3243
rect 4704 3239 4708 3243
rect 4912 3239 4916 3243
rect 5112 3239 5116 3243
rect 5296 3239 5300 3243
rect 5480 3239 5484 3243
rect 5640 3239 5644 3243
rect 3088 3191 3092 3195
rect 2120 3155 2124 3159
rect 2272 3155 2276 3159
rect 2472 3155 2476 3159
rect 2680 3155 2684 3159
rect 2896 3155 2900 3159
rect 3112 3155 3116 3159
rect 3336 3155 3340 3159
rect 3568 3155 3572 3159
rect 3776 3155 3780 3159
rect 320 3111 324 3115
rect 4592 3107 4596 3111
rect 4776 3107 4780 3111
rect 4984 3107 4988 3111
rect 5200 3107 5204 3111
rect 5432 3107 5436 3111
rect 5640 3107 5644 3111
rect 256 3075 260 3079
rect 320 3075 324 3079
rect 496 3075 500 3079
rect 752 3075 756 3079
rect 1000 3075 1004 3079
rect 1240 3075 1244 3079
rect 1472 3075 1476 3079
rect 1704 3075 1708 3079
rect 1912 3075 1916 3079
rect 2744 3047 2748 3051
rect 2880 3047 2884 3051
rect 3024 3047 3028 3051
rect 3176 3047 3180 3051
rect 3336 3047 3340 3051
rect 3496 3047 3500 3051
rect 3664 3047 3668 3051
rect 3200 3039 3204 3043
rect 4352 2999 4356 3003
rect 4552 2999 4556 3003
rect 4768 2999 4772 3003
rect 5008 2999 5012 3003
rect 5264 2999 5268 3003
rect 5520 2999 5524 3003
rect 272 2967 276 2971
rect 504 2967 508 2971
rect 720 2967 724 2971
rect 920 2967 924 2971
rect 1104 2967 1108 2971
rect 1280 2967 1284 2971
rect 1448 2967 1452 2971
rect 1608 2967 1612 2971
rect 1768 2967 1772 2971
rect 1912 2967 1916 2971
rect 2936 2967 2940 2971
rect 3200 2967 3204 2971
rect 3208 2967 3212 2971
rect 1304 2935 1308 2939
rect 3344 2967 3348 2971
rect 3480 2967 3484 2971
rect 528 2883 532 2887
rect 2928 2931 2932 2935
rect 2936 2931 2940 2935
rect 3064 2931 3068 2935
rect 3200 2931 3204 2935
rect 3208 2931 3212 2935
rect 3336 2931 3340 2935
rect 3344 2931 3348 2935
rect 3472 2931 3476 2935
rect 3480 2931 3484 2935
rect 3608 2931 3612 2935
rect 1480 2883 1484 2887
rect 1632 2883 1636 2887
rect 1784 2883 1788 2887
rect 4120 2859 4124 2863
rect 4336 2859 4340 2863
rect 4568 2859 4572 2863
rect 4824 2859 4828 2863
rect 5096 2859 5100 2863
rect 5376 2859 5380 2863
rect 5640 2859 5644 2863
rect 520 2847 524 2851
rect 528 2847 532 2851
rect 720 2847 724 2851
rect 912 2847 916 2851
rect 1096 2847 1100 2851
rect 1272 2847 1276 2851
rect 1304 2847 1308 2851
rect 1440 2847 1444 2851
rect 1480 2847 1484 2851
rect 1608 2847 1612 2851
rect 1632 2847 1636 2851
rect 1768 2847 1772 2851
rect 1784 2847 1788 2851
rect 1912 2847 1916 2851
rect 2120 2771 2124 2775
rect 2136 2771 2140 2775
rect 2264 2771 2268 2775
rect 2272 2771 2276 2775
rect 2432 2771 2436 2775
rect 2456 2771 2460 2775
rect 2592 2771 2596 2775
rect 2760 2771 2764 2775
rect 2928 2771 2932 2775
rect 3096 2771 3100 2775
rect 3264 2771 3268 2775
rect 2136 2739 2140 2743
rect 2272 2739 2276 2743
rect 4016 2747 4020 2751
rect 4152 2747 4156 2751
rect 4288 2747 4292 2751
rect 4424 2747 4428 2751
rect 4560 2747 4564 2751
rect 2456 2739 2460 2743
rect 752 2727 756 2731
rect 776 2727 780 2731
rect 912 2727 916 2731
rect 936 2727 940 2731
rect 1072 2727 1076 2731
rect 1240 2727 1244 2731
rect 1408 2727 1412 2731
rect 1576 2727 1580 2731
rect 776 2695 780 2699
rect 936 2695 940 2699
rect 2512 2691 2516 2695
rect 2504 2655 2508 2659
rect 2512 2655 2516 2659
rect 2640 2655 2644 2659
rect 2784 2655 2788 2659
rect 2928 2655 2932 2659
rect 3072 2655 3076 2659
rect 3216 2655 3220 2659
rect 3360 2655 3364 2659
rect 904 2647 908 2651
rect 1176 2647 1180 2651
rect 1312 2647 1316 2651
rect 1584 2647 1588 2651
rect 1720 2647 1724 2651
rect 4224 2619 4228 2623
rect 4424 2619 4428 2623
rect 4640 2619 4644 2623
rect 4880 2619 4884 2623
rect 5136 2619 5140 2623
rect 5400 2619 5404 2623
rect 5640 2619 5644 2623
rect 896 2611 900 2615
rect 904 2611 908 2615
rect 1032 2611 1036 2615
rect 1168 2611 1172 2615
rect 1176 2611 1180 2615
rect 1304 2611 1308 2615
rect 1312 2611 1316 2615
rect 1440 2611 1444 2615
rect 1576 2611 1580 2615
rect 1584 2611 1588 2615
rect 1712 2611 1716 2615
rect 1720 2611 1724 2615
rect 1848 2611 1852 2615
rect 2608 2543 2612 2547
rect 2616 2543 2620 2547
rect 2744 2543 2748 2547
rect 2752 2543 2756 2547
rect 2880 2543 2884 2547
rect 3016 2543 3020 2547
rect 3152 2543 3156 2547
rect 3288 2543 3292 2547
rect 3424 2543 3428 2547
rect 3560 2543 3564 2547
rect 2616 2511 2620 2515
rect 2752 2511 2756 2515
rect 4592 2507 4596 2511
rect 4728 2507 4732 2511
rect 4864 2507 4868 2511
rect 5000 2507 5004 2511
rect 5136 2507 5140 2511
rect 648 2487 652 2491
rect 784 2487 788 2491
rect 928 2487 932 2491
rect 1080 2487 1084 2491
rect 1232 2487 1236 2491
rect 1392 2487 1396 2491
rect 1552 2487 1556 2491
rect 1584 2487 1588 2491
rect 1712 2487 1716 2491
rect 1880 2487 1884 2491
rect 1584 2455 1588 2459
rect 2432 2411 2436 2415
rect 2640 2411 2644 2415
rect 2840 2411 2844 2415
rect 3032 2411 3036 2415
rect 3224 2411 3228 2415
rect 3408 2411 3412 2415
rect 3592 2411 3596 2415
rect 3776 2411 3780 2415
rect 4968 2411 4972 2415
rect 5104 2411 5108 2415
rect 5240 2411 5244 2415
rect 4824 2375 4828 2379
rect 4960 2375 4964 2379
rect 4968 2375 4972 2379
rect 5096 2375 5100 2379
rect 5104 2375 5108 2379
rect 5232 2375 5236 2379
rect 5240 2375 5244 2379
rect 5368 2375 5372 2379
rect 5504 2375 5508 2379
rect 5640 2375 5644 2379
rect 256 2359 260 2363
rect 464 2359 468 2363
rect 688 2359 692 2363
rect 928 2359 932 2363
rect 1168 2359 1172 2363
rect 1416 2359 1420 2363
rect 1672 2359 1676 2363
rect 1912 2359 1916 2363
rect 2320 2295 2324 2299
rect 2600 2295 2604 2299
rect 2864 2295 2868 2299
rect 3104 2295 3108 2299
rect 3336 2295 3340 2299
rect 3568 2295 3572 2299
rect 3776 2295 3780 2299
rect 288 2287 292 2291
rect 256 2247 260 2251
rect 3984 2255 3988 2259
rect 4280 2255 4284 2259
rect 4592 2255 4596 2259
rect 4888 2255 4892 2259
rect 5184 2255 5188 2259
rect 5480 2255 5484 2259
rect 416 2247 420 2251
rect 648 2247 652 2251
rect 928 2247 932 2251
rect 1248 2247 1252 2251
rect 1592 2247 1596 2251
rect 1912 2247 1916 2251
rect 288 2215 292 2219
rect 2288 2215 2292 2219
rect 2120 2179 2124 2183
rect 2280 2179 2284 2183
rect 2288 2179 2292 2183
rect 2512 2179 2516 2183
rect 2792 2179 2796 2183
rect 3112 2179 3116 2183
rect 3456 2179 3460 2183
rect 3776 2179 3780 2183
rect 4128 2171 4132 2175
rect 872 2143 876 2147
rect 4264 2171 4268 2175
rect 4400 2171 4404 2175
rect 5232 2171 5236 2175
rect 3984 2135 3988 2139
rect 4120 2135 4124 2139
rect 4128 2135 4132 2139
rect 4256 2135 4260 2139
rect 4264 2135 4268 2139
rect 4392 2135 4396 2139
rect 4400 2135 4404 2139
rect 4528 2135 4532 2139
rect 4664 2135 4668 2139
rect 4824 2135 4828 2139
rect 5016 2135 5020 2139
rect 5224 2135 5228 2139
rect 5232 2135 5236 2139
rect 5440 2135 5444 2139
rect 5640 2135 5644 2139
rect 416 2107 420 2111
rect 608 2107 612 2111
rect 816 2107 820 2111
rect 872 2107 876 2111
rect 1040 2107 1044 2111
rect 1272 2107 1276 2111
rect 1512 2107 1516 2111
rect 1760 2107 1764 2111
rect 3984 2007 3988 2011
rect 3992 2007 3996 2011
rect 4120 2007 4124 2011
rect 4128 2007 4132 2011
rect 4256 2007 4260 2011
rect 4264 2007 4268 2011
rect 4392 2007 4396 2011
rect 4400 2007 4404 2011
rect 4528 2007 4532 2011
rect 4536 2007 4540 2011
rect 4664 2007 4668 2011
rect 4816 2007 4820 2011
rect 4992 2007 4996 2011
rect 5032 2007 5036 2011
rect 5184 2007 5188 2011
rect 5224 2007 5228 2011
rect 5376 2007 5380 2011
rect 5576 2007 5580 2011
rect 360 1995 364 1999
rect 496 1995 500 1999
rect 632 1995 636 1999
rect 776 1995 780 1999
rect 920 1995 924 1999
rect 1064 1995 1068 1999
rect 1208 1995 1212 1999
rect 1216 1995 1220 1999
rect 1352 1995 1356 1999
rect 1360 1995 1364 1999
rect 1496 1995 1500 1999
rect 1640 1995 1644 1999
rect 1776 1995 1780 1999
rect 1912 1995 1916 1999
rect 1216 1963 1220 1967
rect 3992 1975 3996 1979
rect 4128 1975 4132 1979
rect 4264 1975 4268 1979
rect 4400 1975 4404 1979
rect 1360 1963 1364 1967
rect 5032 1975 5036 1979
rect 5224 1975 5228 1979
rect 4536 1939 4540 1943
rect 3984 1891 3988 1895
rect 4168 1891 4172 1895
rect 4408 1891 4412 1895
rect 4688 1891 4692 1895
rect 5000 1891 5004 1895
rect 5328 1891 5332 1895
rect 5640 1891 5644 1895
rect 3232 1871 3236 1875
rect 3368 1871 3372 1875
rect 3504 1871 3508 1875
rect 3512 1871 3516 1875
rect 3640 1871 3644 1875
rect 3648 1871 3652 1875
rect 3776 1871 3780 1875
rect 360 1867 364 1871
rect 560 1867 564 1871
rect 752 1867 756 1871
rect 936 1867 940 1871
rect 1112 1867 1116 1871
rect 1280 1867 1284 1871
rect 1448 1867 1452 1871
rect 1608 1867 1612 1871
rect 1768 1867 1772 1871
rect 1912 1867 1916 1871
rect 3512 1839 3516 1843
rect 3648 1839 3652 1843
rect 4504 1783 4508 1787
rect 4640 1783 4644 1787
rect 4776 1783 4780 1787
rect 4912 1783 4916 1787
rect 5048 1783 5052 1787
rect 2128 1779 2132 1783
rect 320 1747 324 1751
rect 384 1747 388 1751
rect 560 1747 564 1751
rect 792 1747 796 1751
rect 1024 1747 1028 1751
rect 1256 1747 1260 1751
rect 1488 1747 1492 1751
rect 2264 1779 2268 1783
rect 2416 1779 2420 1783
rect 2568 1779 2572 1783
rect 3032 1779 3036 1783
rect 3648 1779 3652 1783
rect 2120 1743 2124 1747
rect 2128 1743 2132 1747
rect 2256 1743 2260 1747
rect 2264 1743 2268 1747
rect 2392 1743 2396 1747
rect 2416 1743 2420 1747
rect 2544 1743 2548 1747
rect 2568 1743 2572 1747
rect 2704 1743 2708 1747
rect 2864 1743 2868 1747
rect 3024 1743 3028 1747
rect 3032 1743 3036 1747
rect 3176 1743 3180 1747
rect 3328 1743 3332 1747
rect 3480 1743 3484 1747
rect 3640 1743 3644 1747
rect 3648 1743 3652 1747
rect 3776 1743 3780 1747
rect 384 1715 388 1719
rect 4696 1687 4700 1691
rect 816 1655 820 1659
rect 4832 1679 4836 1683
rect 5328 1671 5332 1675
rect 4688 1651 4692 1655
rect 4696 1651 4700 1655
rect 4824 1651 4828 1655
rect 4832 1651 4836 1655
rect 4960 1651 4964 1655
rect 5096 1651 5100 1655
rect 5232 1651 5236 1655
rect 2120 1623 2124 1627
rect 2264 1623 2268 1627
rect 2416 1623 2420 1627
rect 2576 1623 2580 1627
rect 2736 1623 2740 1627
rect 2888 1623 2892 1627
rect 3040 1623 3044 1627
rect 3200 1623 3204 1627
rect 3216 1623 3220 1627
rect 3360 1623 3364 1627
rect 3520 1623 3524 1627
rect 256 1619 260 1623
rect 488 1619 492 1623
rect 744 1619 748 1623
rect 816 1619 820 1623
rect 1000 1619 1004 1623
rect 1264 1619 1268 1623
rect 2128 1531 2132 1535
rect 256 1499 260 1503
rect 424 1499 428 1503
rect 608 1499 612 1503
rect 792 1499 796 1503
rect 984 1499 988 1503
rect 1176 1499 1180 1503
rect 2808 1531 2812 1535
rect 2264 1523 2268 1527
rect 2944 1531 2948 1535
rect 3080 1531 3084 1535
rect 3216 1531 3220 1535
rect 3352 1531 3356 1535
rect 3488 1531 3492 1535
rect 5368 1651 5372 1655
rect 5504 1651 5508 1655
rect 5640 1651 5644 1655
rect 4688 1527 4692 1531
rect 4824 1527 4828 1531
rect 4960 1527 4964 1531
rect 5096 1527 5100 1531
rect 5232 1527 5236 1531
rect 5328 1527 5332 1531
rect 5368 1527 5372 1531
rect 5504 1527 5508 1531
rect 5640 1527 5644 1531
rect 5480 1519 5484 1523
rect 2120 1495 2124 1499
rect 2128 1495 2132 1499
rect 2256 1495 2260 1499
rect 2264 1495 2268 1499
rect 2392 1495 2396 1499
rect 2528 1495 2532 1499
rect 2664 1495 2668 1499
rect 2800 1495 2804 1499
rect 2808 1495 2812 1499
rect 2936 1495 2940 1499
rect 2944 1495 2948 1499
rect 3072 1495 3076 1499
rect 3080 1495 3084 1499
rect 3208 1495 3212 1499
rect 3344 1495 3348 1499
rect 3352 1495 3356 1499
rect 3480 1495 3484 1499
rect 3488 1495 3492 1499
rect 3616 1495 3620 1499
rect 2264 1375 2268 1379
rect 2272 1375 2276 1379
rect 2400 1375 2404 1379
rect 2536 1375 2540 1379
rect 2672 1375 2676 1379
rect 2808 1375 2812 1379
rect 2944 1375 2948 1379
rect 3080 1375 3084 1379
rect 3216 1375 3220 1379
rect 3352 1375 3356 1379
rect 4944 1375 4948 1379
rect 256 1371 260 1375
rect 520 1371 524 1375
rect 808 1371 812 1375
rect 1096 1371 1100 1375
rect 1384 1371 1388 1375
rect 2272 1343 2276 1347
rect 5080 1375 5084 1379
rect 5216 1375 5220 1379
rect 5472 1375 5476 1379
rect 4936 1339 4940 1343
rect 4944 1339 4948 1343
rect 5072 1339 5076 1343
rect 5080 1339 5084 1343
rect 5208 1339 5212 1343
rect 5216 1339 5220 1343
rect 5344 1339 5348 1343
rect 5480 1339 5484 1343
rect 5616 1339 5620 1343
rect 2400 1295 2404 1299
rect 256 1263 260 1267
rect 552 1263 556 1267
rect 872 1263 876 1267
rect 1192 1263 1196 1267
rect 1200 1263 1204 1267
rect 1520 1263 1524 1267
rect 3024 1295 3028 1299
rect 3264 1295 3268 1299
rect 2256 1259 2260 1263
rect 2392 1259 2396 1263
rect 2400 1259 2404 1263
rect 2528 1259 2532 1263
rect 2680 1259 2684 1263
rect 2840 1259 2844 1263
rect 3016 1259 3020 1263
rect 3024 1259 3028 1263
rect 3200 1259 3204 1263
rect 3264 1259 3268 1263
rect 3392 1259 3396 1263
rect 3592 1259 3596 1263
rect 3776 1259 3780 1263
rect 4832 1227 4836 1231
rect 4976 1227 4980 1231
rect 5128 1227 5132 1231
rect 5288 1227 5292 1231
rect 5456 1227 5460 1231
rect 5624 1227 5628 1231
rect 992 1159 996 1163
rect 1192 1159 1196 1163
rect 1200 1159 1204 1163
rect 2120 1151 2124 1155
rect 2336 1151 2340 1155
rect 2576 1151 2580 1155
rect 2816 1151 2820 1155
rect 3056 1151 3060 1155
rect 3304 1151 3308 1155
rect 3552 1151 3556 1155
rect 3776 1151 3780 1155
rect 256 1123 260 1127
rect 456 1123 460 1127
rect 688 1123 692 1127
rect 928 1123 932 1127
rect 992 1123 996 1127
rect 1168 1123 1172 1127
rect 1192 1123 1196 1127
rect 1408 1123 1412 1127
rect 1648 1123 1652 1127
rect 1896 1123 1900 1127
rect 3984 1103 3988 1107
rect 4192 1103 4196 1107
rect 4424 1103 4428 1107
rect 4664 1103 4668 1107
rect 4904 1103 4908 1107
rect 5152 1103 5156 1107
rect 5408 1103 5412 1107
rect 5640 1103 5644 1107
rect 360 1015 364 1019
rect 392 1015 396 1019
rect 536 1015 540 1019
rect 712 1015 716 1019
rect 880 1015 884 1019
rect 1048 1015 1052 1019
rect 1208 1015 1212 1019
rect 1368 1015 1372 1019
rect 1528 1015 1532 1019
rect 1688 1015 1692 1019
rect 1848 1015 1852 1019
rect 3216 1011 3220 1015
rect 3368 1011 3372 1015
rect 3520 1011 3524 1015
rect 3984 995 3988 999
rect 4168 995 4172 999
rect 4376 995 4380 999
rect 4608 995 4612 999
rect 4856 995 4860 999
rect 5120 995 5124 999
rect 5392 995 5396 999
rect 5640 995 5644 999
rect 392 983 396 987
rect 1240 983 1244 987
rect 1392 931 1396 935
rect 1776 931 1780 935
rect 1968 931 1972 935
rect 352 895 356 899
rect 504 895 508 899
rect 664 895 668 899
rect 840 895 844 899
rect 1016 895 1020 899
rect 1200 895 1204 899
rect 1240 895 1244 899
rect 1384 895 1388 899
rect 1392 895 1396 899
rect 1568 895 1572 899
rect 1752 895 1756 899
rect 1776 895 1780 899
rect 1912 895 1916 899
rect 5376 915 5380 919
rect 4096 879 4100 883
rect 4304 879 4308 883
rect 4528 879 4532 883
rect 4768 879 4772 883
rect 5024 879 5028 883
rect 5296 879 5300 883
rect 5376 879 5380 883
rect 5568 879 5572 883
rect 1968 875 1972 879
rect 2144 875 2148 879
rect 2448 875 2452 879
rect 2744 875 2748 879
rect 3024 875 3028 879
rect 3304 875 3308 879
rect 3592 875 3596 879
rect 472 771 476 775
rect 752 771 756 775
rect 1040 771 1044 775
rect 1336 771 1340 775
rect 1632 771 1636 775
rect 1912 771 1916 775
rect 3984 771 3988 775
rect 4144 771 4148 775
rect 4376 771 4380 775
rect 4504 771 4508 775
rect 4656 771 4660 775
rect 4976 771 4980 775
rect 5320 771 5324 775
rect 5640 771 5644 775
rect 2120 759 2124 763
rect 2376 759 2380 763
rect 2648 759 2652 763
rect 2896 759 2900 763
rect 3128 759 3132 763
rect 3352 759 3356 763
rect 3576 759 3580 763
rect 3776 759 3780 763
rect 1320 691 1324 695
rect 584 675 588 679
rect 1472 691 1476 695
rect 1640 691 1644 695
rect 1784 691 1788 695
rect 4128 683 4132 687
rect 256 655 260 659
rect 432 655 436 659
rect 584 655 588 659
rect 624 655 628 659
rect 808 655 812 659
rect 984 655 988 659
rect 1152 655 1156 659
rect 1312 655 1316 659
rect 1320 655 1324 659
rect 1464 655 1468 659
rect 1472 655 1476 659
rect 1616 655 1620 659
rect 1640 655 1644 659
rect 1776 655 1780 659
rect 1784 655 1788 659
rect 1912 655 1916 659
rect 4264 683 4268 687
rect 4400 683 4404 687
rect 4504 683 4508 687
rect 3984 647 3988 651
rect 4120 647 4124 651
rect 4128 647 4132 651
rect 4256 647 4260 651
rect 4264 647 4268 651
rect 4392 647 4396 651
rect 4400 647 4404 651
rect 4528 647 4532 651
rect 4696 647 4700 651
rect 4896 647 4900 651
rect 5120 647 5124 651
rect 5352 647 5356 651
rect 5584 647 5588 651
rect 4408 607 4412 611
rect 256 547 260 551
rect 472 547 476 551
rect 696 547 700 551
rect 760 547 764 551
rect 904 547 908 551
rect 944 547 948 551
rect 1096 547 1100 551
rect 1272 547 1276 551
rect 1440 547 1444 551
rect 1608 547 1612 551
rect 1632 547 1636 551
rect 1768 547 1772 551
rect 1912 547 1916 551
rect 760 515 764 519
rect 944 515 948 519
rect 3984 539 3988 543
rect 4120 539 4124 543
rect 4128 539 4132 543
rect 4256 539 4260 543
rect 4392 539 4396 543
rect 3408 519 3412 523
rect 3544 519 3548 523
rect 3680 519 3684 523
rect 1632 515 1636 519
rect 4128 507 4132 511
rect 4576 539 4580 543
rect 4792 539 4796 543
rect 5032 539 5036 543
rect 5288 539 5292 543
rect 5544 539 5548 543
rect 4408 507 4412 511
rect 1960 467 1964 471
rect 256 431 260 435
rect 552 431 556 435
rect 888 431 892 435
rect 1232 431 1236 435
rect 1584 431 1588 435
rect 1912 431 1916 435
rect 2144 439 2148 443
rect 5368 435 5372 439
rect 4576 411 4580 415
rect 4776 411 4780 415
rect 4984 411 4988 415
rect 5192 411 5196 415
rect 1960 403 1964 407
rect 2120 403 2124 407
rect 2144 403 2148 407
rect 2280 403 2284 407
rect 2472 403 2476 407
rect 2664 403 2668 407
rect 2856 403 2860 407
rect 3048 403 3052 407
rect 3240 403 3244 407
rect 3424 403 3428 407
rect 3608 403 3612 407
rect 3776 403 3780 407
rect 336 307 340 311
rect 488 307 492 311
rect 648 307 652 311
rect 808 307 812 311
rect 832 307 836 311
rect 968 307 972 311
rect 992 307 996 311
rect 1128 307 1132 311
rect 832 275 836 279
rect 5408 411 5412 415
rect 5632 411 5636 415
rect 992 275 996 279
rect 4416 299 4420 303
rect 4848 299 4852 303
rect 5008 299 5012 303
rect 5168 299 5172 303
rect 5328 299 5332 303
rect 5368 299 5372 303
rect 5496 299 5500 303
rect 5640 299 5644 303
rect 2144 271 2148 275
rect 2280 271 2284 275
rect 2416 271 2420 275
rect 2552 271 2556 275
rect 2688 271 2692 275
rect 2696 271 2700 275
rect 2824 271 2828 275
rect 2960 271 2964 275
rect 3096 271 3100 275
rect 3232 271 3236 275
rect 3368 271 3372 275
rect 3504 271 3508 275
rect 3640 271 3644 275
rect 3776 271 3780 275
rect 2696 239 2700 243
rect 280 195 284 199
rect 416 195 420 199
rect 552 195 556 199
rect 688 195 692 199
rect 960 195 964 199
rect 1096 195 1100 199
rect 4416 179 4420 183
rect 4424 179 4428 183
rect 2128 175 2132 179
rect 272 159 276 163
rect 280 159 284 163
rect 408 159 412 163
rect 416 159 420 163
rect 544 159 548 163
rect 552 159 556 163
rect 680 159 684 163
rect 688 159 692 163
rect 816 159 820 163
rect 952 159 956 163
rect 960 159 964 163
rect 1088 159 1092 163
rect 1096 159 1100 163
rect 1224 159 1228 163
rect 2264 175 2268 179
rect 2400 175 2404 179
rect 2672 175 2676 179
rect 2808 175 2812 179
rect 3080 175 3084 179
rect 3216 175 3220 179
rect 3488 175 3492 179
rect 3624 175 3628 179
rect 4560 179 4564 183
rect 4696 179 4700 183
rect 4968 179 4972 183
rect 5104 179 5108 183
rect 5240 179 5244 183
rect 4416 143 4420 147
rect 4424 143 4428 147
rect 4552 143 4556 147
rect 4560 143 4564 147
rect 4688 143 4692 147
rect 4696 143 4700 147
rect 4824 143 4828 147
rect 4960 143 4964 147
rect 4968 143 4972 147
rect 5096 143 5100 147
rect 5104 143 5108 147
rect 5232 143 5236 147
rect 5240 143 5244 147
rect 5368 143 5372 147
rect 5640 143 5644 147
rect 2120 139 2124 143
rect 2128 139 2132 143
rect 2256 139 2260 143
rect 2264 139 2268 143
rect 2392 139 2396 143
rect 2400 139 2404 143
rect 2528 139 2532 143
rect 2664 139 2668 143
rect 2672 139 2676 143
rect 2800 139 2804 143
rect 2808 139 2812 143
rect 2936 139 2940 143
rect 3072 139 3076 143
rect 3080 139 3084 143
rect 3208 139 3212 143
rect 3216 139 3220 143
rect 3344 139 3348 143
rect 3480 139 3484 143
rect 3488 139 3492 143
rect 3616 139 3620 143
rect 3624 139 3628 143
rect 3752 139 3756 143
<< m2 >>
rect 258 5735 264 5736
rect 258 5731 259 5735
rect 263 5734 264 5735
rect 399 5735 405 5736
rect 263 5732 285 5734
rect 263 5731 264 5732
rect 258 5730 264 5731
rect 399 5731 400 5735
rect 404 5734 405 5735
rect 404 5732 421 5734
rect 404 5731 405 5732
rect 399 5730 405 5731
rect 255 5699 264 5700
rect 255 5695 256 5699
rect 263 5695 264 5699
rect 255 5694 264 5695
rect 391 5699 397 5700
rect 391 5695 392 5699
rect 396 5698 397 5699
rect 399 5699 405 5700
rect 399 5698 400 5699
rect 396 5696 400 5698
rect 396 5695 397 5696
rect 391 5694 397 5695
rect 399 5695 400 5696
rect 404 5695 405 5699
rect 399 5694 405 5695
rect 422 5699 428 5700
rect 422 5695 423 5699
rect 427 5698 428 5699
rect 527 5699 533 5700
rect 527 5698 528 5699
rect 427 5696 528 5698
rect 427 5695 428 5696
rect 422 5694 428 5695
rect 527 5695 528 5696
rect 532 5695 533 5699
rect 527 5694 533 5695
rect 110 5692 116 5693
rect 1934 5692 1940 5693
rect 110 5688 111 5692
rect 115 5688 116 5692
rect 110 5687 116 5688
rect 130 5691 136 5692
rect 130 5687 131 5691
rect 135 5687 136 5691
rect 130 5686 136 5687
rect 266 5691 272 5692
rect 266 5687 267 5691
rect 271 5687 272 5691
rect 266 5686 272 5687
rect 402 5691 408 5692
rect 402 5687 403 5691
rect 407 5687 408 5691
rect 1934 5688 1935 5692
rect 1939 5688 1940 5692
rect 1934 5687 1940 5688
rect 402 5686 408 5687
rect 158 5676 164 5677
rect 110 5675 116 5676
rect 110 5671 111 5675
rect 115 5671 116 5675
rect 158 5672 159 5676
rect 163 5672 164 5676
rect 158 5671 164 5672
rect 294 5676 300 5677
rect 294 5672 295 5676
rect 299 5672 300 5676
rect 294 5671 300 5672
rect 430 5676 436 5677
rect 430 5672 431 5676
rect 435 5672 436 5676
rect 430 5671 436 5672
rect 1934 5675 1940 5676
rect 1934 5671 1935 5675
rect 1939 5671 1940 5675
rect 110 5670 116 5671
rect 1934 5670 1940 5671
rect 4599 5671 4605 5672
rect 2151 5667 2157 5668
rect 2151 5666 2152 5667
rect 2085 5664 2152 5666
rect 2151 5663 2152 5664
rect 2156 5663 2157 5667
rect 2367 5667 2373 5668
rect 2367 5666 2368 5667
rect 2261 5664 2368 5666
rect 2151 5662 2157 5663
rect 2367 5663 2368 5664
rect 2372 5663 2373 5667
rect 2535 5667 2541 5668
rect 2535 5666 2536 5667
rect 2461 5664 2536 5666
rect 2367 5662 2373 5663
rect 2535 5663 2536 5664
rect 2540 5663 2541 5667
rect 2874 5667 2880 5668
rect 2535 5662 2541 5663
rect 2650 5663 2656 5664
rect 2650 5659 2651 5663
rect 2655 5659 2656 5663
rect 2874 5663 2875 5667
rect 2879 5666 2880 5667
rect 3058 5667 3064 5668
rect 2879 5664 2949 5666
rect 2879 5663 2880 5664
rect 2874 5662 2880 5663
rect 3058 5663 3059 5667
rect 3063 5666 3064 5667
rect 3234 5667 3240 5668
rect 3063 5664 3125 5666
rect 3063 5663 3064 5664
rect 3058 5662 3064 5663
rect 3234 5663 3235 5667
rect 3239 5666 3240 5667
rect 3402 5667 3408 5668
rect 3239 5664 3293 5666
rect 3239 5663 3240 5664
rect 3234 5662 3240 5663
rect 3402 5663 3403 5667
rect 3407 5666 3408 5667
rect 3570 5667 3576 5668
rect 3407 5664 3461 5666
rect 3407 5663 3408 5664
rect 3402 5662 3408 5663
rect 3570 5663 3571 5667
rect 3575 5666 3576 5667
rect 4554 5667 4560 5668
rect 3575 5664 3637 5666
rect 3575 5663 3576 5664
rect 3570 5662 3576 5663
rect 4554 5663 4555 5667
rect 4559 5663 4560 5667
rect 4599 5667 4600 5671
rect 4604 5670 4605 5671
rect 4735 5671 4741 5672
rect 4604 5668 4621 5670
rect 4604 5667 4605 5668
rect 4599 5666 4605 5667
rect 4735 5667 4736 5671
rect 4740 5670 4741 5671
rect 4871 5671 4877 5672
rect 4740 5668 4757 5670
rect 4740 5667 4741 5668
rect 4735 5666 4741 5667
rect 4871 5667 4872 5671
rect 4876 5670 4877 5671
rect 4876 5668 4893 5670
rect 4876 5667 4877 5668
rect 4871 5666 4877 5667
rect 4554 5662 4560 5663
rect 2650 5658 2656 5659
rect 2832 5650 2834 5661
rect 3066 5651 3072 5652
rect 3066 5650 3067 5651
rect 2832 5648 3067 5650
rect 3066 5647 3067 5648
rect 3071 5647 3072 5651
rect 3066 5646 3072 5647
rect 4591 5635 4597 5636
rect 1942 5631 1948 5632
rect 1942 5627 1943 5631
rect 1947 5630 1948 5631
rect 2119 5631 2125 5632
rect 2119 5630 2120 5631
rect 1947 5628 2120 5630
rect 1947 5627 1948 5628
rect 1942 5626 1948 5627
rect 2119 5627 2120 5628
rect 2124 5627 2125 5631
rect 2119 5626 2125 5627
rect 2151 5631 2157 5632
rect 2151 5627 2152 5631
rect 2156 5630 2157 5631
rect 2295 5631 2301 5632
rect 2295 5630 2296 5631
rect 2156 5628 2296 5630
rect 2156 5627 2157 5628
rect 2151 5626 2157 5627
rect 2295 5627 2296 5628
rect 2300 5627 2301 5631
rect 2295 5626 2301 5627
rect 2367 5631 2373 5632
rect 2367 5627 2368 5631
rect 2372 5630 2373 5631
rect 2495 5631 2501 5632
rect 2495 5630 2496 5631
rect 2372 5628 2496 5630
rect 2372 5627 2373 5628
rect 2367 5626 2373 5627
rect 2495 5627 2496 5628
rect 2500 5627 2501 5631
rect 2495 5626 2501 5627
rect 2535 5631 2541 5632
rect 2535 5627 2536 5631
rect 2540 5630 2541 5631
rect 2687 5631 2693 5632
rect 2687 5630 2688 5631
rect 2540 5628 2688 5630
rect 2540 5627 2541 5628
rect 2535 5626 2541 5627
rect 2687 5627 2688 5628
rect 2692 5627 2693 5631
rect 2687 5626 2693 5627
rect 2871 5631 2880 5632
rect 2871 5627 2872 5631
rect 2879 5627 2880 5631
rect 2871 5626 2880 5627
rect 3055 5631 3064 5632
rect 3055 5627 3056 5631
rect 3063 5627 3064 5631
rect 3055 5626 3064 5627
rect 3231 5631 3240 5632
rect 3231 5627 3232 5631
rect 3239 5627 3240 5631
rect 3231 5626 3240 5627
rect 3399 5631 3408 5632
rect 3399 5627 3400 5631
rect 3407 5627 3408 5631
rect 3399 5626 3408 5627
rect 3567 5631 3576 5632
rect 3567 5627 3568 5631
rect 3575 5627 3576 5631
rect 3567 5626 3576 5627
rect 3738 5631 3749 5632
rect 3738 5627 3739 5631
rect 3743 5627 3744 5631
rect 3748 5627 3749 5631
rect 4591 5631 4592 5635
rect 4596 5634 4597 5635
rect 4599 5635 4605 5636
rect 4599 5634 4600 5635
rect 4596 5632 4600 5634
rect 4596 5631 4597 5632
rect 4591 5630 4597 5631
rect 4599 5631 4600 5632
rect 4604 5631 4605 5635
rect 4599 5630 4605 5631
rect 4727 5635 4733 5636
rect 4727 5631 4728 5635
rect 4732 5634 4733 5635
rect 4735 5635 4741 5636
rect 4735 5634 4736 5635
rect 4732 5632 4736 5634
rect 4732 5631 4733 5632
rect 4727 5630 4733 5631
rect 4735 5631 4736 5632
rect 4740 5631 4741 5635
rect 4735 5630 4741 5631
rect 4863 5635 4869 5636
rect 4863 5631 4864 5635
rect 4868 5634 4869 5635
rect 4871 5635 4877 5636
rect 4871 5634 4872 5635
rect 4868 5632 4872 5634
rect 4868 5631 4869 5632
rect 4863 5630 4869 5631
rect 4871 5631 4872 5632
rect 4876 5631 4877 5635
rect 4871 5630 4877 5631
rect 4910 5635 4916 5636
rect 4910 5631 4911 5635
rect 4915 5634 4916 5635
rect 4999 5635 5005 5636
rect 4999 5634 5000 5635
rect 4915 5632 5000 5634
rect 4915 5631 4916 5632
rect 4910 5630 4916 5631
rect 4999 5631 5000 5632
rect 5004 5631 5005 5635
rect 4999 5630 5005 5631
rect 3738 5626 3749 5627
rect 3838 5628 3844 5629
rect 5662 5628 5668 5629
rect 1974 5624 1980 5625
rect 3798 5624 3804 5625
rect 1974 5620 1975 5624
rect 1979 5620 1980 5624
rect 1974 5619 1980 5620
rect 1994 5623 2000 5624
rect 1994 5619 1995 5623
rect 1999 5619 2000 5623
rect 1994 5618 2000 5619
rect 2170 5623 2176 5624
rect 2170 5619 2171 5623
rect 2175 5619 2176 5623
rect 2170 5618 2176 5619
rect 2370 5623 2376 5624
rect 2370 5619 2371 5623
rect 2375 5619 2376 5623
rect 2370 5618 2376 5619
rect 2562 5623 2568 5624
rect 2562 5619 2563 5623
rect 2567 5619 2568 5623
rect 2562 5618 2568 5619
rect 2746 5623 2752 5624
rect 2746 5619 2747 5623
rect 2751 5619 2752 5623
rect 2746 5618 2752 5619
rect 2930 5623 2936 5624
rect 2930 5619 2931 5623
rect 2935 5619 2936 5623
rect 2930 5618 2936 5619
rect 3106 5623 3112 5624
rect 3106 5619 3107 5623
rect 3111 5619 3112 5623
rect 3106 5618 3112 5619
rect 3274 5623 3280 5624
rect 3274 5619 3275 5623
rect 3279 5619 3280 5623
rect 3274 5618 3280 5619
rect 3442 5623 3448 5624
rect 3442 5619 3443 5623
rect 3447 5619 3448 5623
rect 3442 5618 3448 5619
rect 3618 5623 3624 5624
rect 3618 5619 3619 5623
rect 3623 5619 3624 5623
rect 3798 5620 3799 5624
rect 3803 5620 3804 5624
rect 3838 5624 3839 5628
rect 3843 5624 3844 5628
rect 3838 5623 3844 5624
rect 4466 5627 4472 5628
rect 4466 5623 4467 5627
rect 4471 5623 4472 5627
rect 4466 5622 4472 5623
rect 4602 5627 4608 5628
rect 4602 5623 4603 5627
rect 4607 5623 4608 5627
rect 4602 5622 4608 5623
rect 4738 5627 4744 5628
rect 4738 5623 4739 5627
rect 4743 5623 4744 5627
rect 4738 5622 4744 5623
rect 4874 5627 4880 5628
rect 4874 5623 4875 5627
rect 4879 5623 4880 5627
rect 5662 5624 5663 5628
rect 5667 5624 5668 5628
rect 5662 5623 5668 5624
rect 4874 5622 4880 5623
rect 3798 5619 3804 5620
rect 3618 5618 3624 5619
rect 110 5617 116 5618
rect 1934 5617 1940 5618
rect 110 5613 111 5617
rect 115 5613 116 5617
rect 110 5612 116 5613
rect 342 5616 348 5617
rect 342 5612 343 5616
rect 347 5612 348 5616
rect 342 5611 348 5612
rect 534 5616 540 5617
rect 534 5612 535 5616
rect 539 5612 540 5616
rect 534 5611 540 5612
rect 734 5616 740 5617
rect 734 5612 735 5616
rect 739 5612 740 5616
rect 734 5611 740 5612
rect 942 5616 948 5617
rect 942 5612 943 5616
rect 947 5612 948 5616
rect 942 5611 948 5612
rect 1158 5616 1164 5617
rect 1158 5612 1159 5616
rect 1163 5612 1164 5616
rect 1158 5611 1164 5612
rect 1382 5616 1388 5617
rect 1382 5612 1383 5616
rect 1387 5612 1388 5616
rect 1382 5611 1388 5612
rect 1606 5616 1612 5617
rect 1606 5612 1607 5616
rect 1611 5612 1612 5616
rect 1606 5611 1612 5612
rect 1814 5616 1820 5617
rect 1814 5612 1815 5616
rect 1819 5612 1820 5616
rect 1934 5613 1935 5617
rect 1939 5613 1940 5617
rect 1934 5612 1940 5613
rect 4494 5612 4500 5613
rect 1814 5611 1820 5612
rect 3838 5611 3844 5612
rect 2022 5608 2028 5609
rect 1974 5607 1980 5608
rect 1974 5603 1975 5607
rect 1979 5603 1980 5607
rect 2022 5604 2023 5608
rect 2027 5604 2028 5608
rect 2022 5603 2028 5604
rect 2198 5608 2204 5609
rect 2198 5604 2199 5608
rect 2203 5604 2204 5608
rect 2198 5603 2204 5604
rect 2398 5608 2404 5609
rect 2398 5604 2399 5608
rect 2403 5604 2404 5608
rect 2398 5603 2404 5604
rect 2590 5608 2596 5609
rect 2590 5604 2591 5608
rect 2595 5604 2596 5608
rect 2590 5603 2596 5604
rect 2774 5608 2780 5609
rect 2774 5604 2775 5608
rect 2779 5604 2780 5608
rect 2774 5603 2780 5604
rect 2958 5608 2964 5609
rect 2958 5604 2959 5608
rect 2963 5604 2964 5608
rect 2958 5603 2964 5604
rect 3134 5608 3140 5609
rect 3134 5604 3135 5608
rect 3139 5604 3140 5608
rect 3134 5603 3140 5604
rect 3302 5608 3308 5609
rect 3302 5604 3303 5608
rect 3307 5604 3308 5608
rect 3302 5603 3308 5604
rect 3470 5608 3476 5609
rect 3470 5604 3471 5608
rect 3475 5604 3476 5608
rect 3470 5603 3476 5604
rect 3646 5608 3652 5609
rect 3646 5604 3647 5608
rect 3651 5604 3652 5608
rect 3646 5603 3652 5604
rect 3798 5607 3804 5608
rect 3798 5603 3799 5607
rect 3803 5603 3804 5607
rect 3838 5607 3839 5611
rect 3843 5607 3844 5611
rect 4494 5608 4495 5612
rect 4499 5608 4500 5612
rect 4494 5607 4500 5608
rect 4630 5612 4636 5613
rect 4630 5608 4631 5612
rect 4635 5608 4636 5612
rect 4630 5607 4636 5608
rect 4766 5612 4772 5613
rect 4766 5608 4767 5612
rect 4771 5608 4772 5612
rect 4766 5607 4772 5608
rect 4902 5612 4908 5613
rect 4902 5608 4903 5612
rect 4907 5608 4908 5612
rect 4902 5607 4908 5608
rect 5662 5611 5668 5612
rect 5662 5607 5663 5611
rect 5667 5607 5668 5611
rect 3838 5606 3844 5607
rect 5662 5606 5668 5607
rect 1974 5602 1980 5603
rect 3798 5602 3804 5603
rect 314 5601 320 5602
rect 110 5600 116 5601
rect 110 5596 111 5600
rect 115 5596 116 5600
rect 314 5597 315 5601
rect 319 5597 320 5601
rect 314 5596 320 5597
rect 506 5601 512 5602
rect 506 5597 507 5601
rect 511 5597 512 5601
rect 506 5596 512 5597
rect 706 5601 712 5602
rect 706 5597 707 5601
rect 711 5597 712 5601
rect 706 5596 712 5597
rect 914 5601 920 5602
rect 914 5597 915 5601
rect 919 5597 920 5601
rect 914 5596 920 5597
rect 1130 5601 1136 5602
rect 1130 5597 1131 5601
rect 1135 5597 1136 5601
rect 1130 5596 1136 5597
rect 1354 5601 1360 5602
rect 1354 5597 1355 5601
rect 1359 5597 1360 5601
rect 1354 5596 1360 5597
rect 1578 5601 1584 5602
rect 1578 5597 1579 5601
rect 1583 5597 1584 5601
rect 1578 5596 1584 5597
rect 1786 5601 1792 5602
rect 1786 5597 1787 5601
rect 1791 5597 1792 5601
rect 1786 5596 1792 5597
rect 1934 5600 1940 5601
rect 1934 5596 1935 5600
rect 1939 5596 1940 5600
rect 110 5595 116 5596
rect 1934 5595 1940 5596
rect 439 5591 445 5592
rect 439 5587 440 5591
rect 444 5590 445 5591
rect 522 5591 528 5592
rect 522 5590 523 5591
rect 444 5588 523 5590
rect 444 5587 445 5588
rect 439 5586 445 5587
rect 522 5587 523 5588
rect 527 5587 528 5591
rect 522 5586 528 5587
rect 631 5591 637 5592
rect 631 5587 632 5591
rect 636 5590 637 5591
rect 722 5591 728 5592
rect 722 5590 723 5591
rect 636 5588 723 5590
rect 636 5587 637 5588
rect 631 5586 637 5587
rect 722 5587 723 5588
rect 727 5587 728 5591
rect 722 5586 728 5587
rect 831 5591 837 5592
rect 831 5587 832 5591
rect 836 5590 837 5591
rect 930 5591 936 5592
rect 930 5590 931 5591
rect 836 5588 931 5590
rect 836 5587 837 5588
rect 831 5586 837 5587
rect 930 5587 931 5588
rect 935 5587 936 5591
rect 930 5586 936 5587
rect 1039 5591 1045 5592
rect 1039 5587 1040 5591
rect 1044 5590 1045 5591
rect 1146 5591 1152 5592
rect 1146 5590 1147 5591
rect 1044 5588 1147 5590
rect 1044 5587 1045 5588
rect 1039 5586 1045 5587
rect 1146 5587 1147 5588
rect 1151 5587 1152 5591
rect 1255 5591 1261 5592
rect 1255 5590 1256 5591
rect 1146 5586 1152 5587
rect 1156 5588 1256 5590
rect 998 5583 1004 5584
rect 998 5579 999 5583
rect 1003 5582 1004 5583
rect 1156 5582 1158 5588
rect 1255 5587 1256 5588
rect 1260 5587 1261 5591
rect 1255 5586 1261 5587
rect 1479 5591 1485 5592
rect 1479 5587 1480 5591
rect 1484 5590 1485 5591
rect 1535 5591 1541 5592
rect 1535 5590 1536 5591
rect 1484 5588 1536 5590
rect 1484 5587 1485 5588
rect 1479 5586 1485 5587
rect 1535 5587 1536 5588
rect 1540 5587 1541 5591
rect 1535 5586 1541 5587
rect 1575 5591 1581 5592
rect 1575 5587 1576 5591
rect 1580 5590 1581 5591
rect 1703 5591 1709 5592
rect 1703 5590 1704 5591
rect 1580 5588 1704 5590
rect 1580 5587 1581 5588
rect 1575 5586 1581 5587
rect 1703 5587 1704 5588
rect 1708 5587 1709 5591
rect 1703 5586 1709 5587
rect 1751 5591 1757 5592
rect 1751 5587 1752 5591
rect 1756 5590 1757 5591
rect 1911 5591 1917 5592
rect 1911 5590 1912 5591
rect 1756 5588 1912 5590
rect 1756 5587 1757 5588
rect 1751 5586 1757 5587
rect 1911 5587 1912 5588
rect 1916 5587 1917 5591
rect 1911 5586 1917 5587
rect 1003 5580 1158 5582
rect 1003 5579 1004 5580
rect 998 5578 1004 5579
rect 422 5559 428 5560
rect 422 5558 423 5559
rect 405 5556 423 5558
rect 422 5555 423 5556
rect 427 5555 428 5559
rect 422 5554 428 5555
rect 522 5559 528 5560
rect 522 5555 523 5559
rect 527 5555 528 5559
rect 522 5554 528 5555
rect 722 5559 728 5560
rect 722 5555 723 5559
rect 727 5555 728 5559
rect 722 5554 728 5555
rect 930 5559 936 5560
rect 930 5555 931 5559
rect 935 5555 936 5559
rect 930 5554 936 5555
rect 1146 5559 1152 5560
rect 1146 5555 1147 5559
rect 1151 5555 1152 5559
rect 1575 5559 1581 5560
rect 1575 5558 1576 5559
rect 1445 5556 1576 5558
rect 1146 5554 1152 5555
rect 1575 5555 1576 5556
rect 1580 5555 1581 5559
rect 1751 5559 1757 5560
rect 1751 5558 1752 5559
rect 1669 5556 1752 5558
rect 1575 5554 1581 5555
rect 1751 5555 1752 5556
rect 1756 5555 1757 5559
rect 1942 5559 1948 5560
rect 1942 5558 1943 5559
rect 1877 5556 1943 5558
rect 1751 5554 1757 5555
rect 1942 5555 1943 5556
rect 1947 5555 1948 5559
rect 1942 5554 1948 5555
rect 3838 5553 3844 5554
rect 5662 5553 5668 5554
rect 1974 5549 1980 5550
rect 3798 5549 3804 5550
rect 1974 5545 1975 5549
rect 1979 5545 1980 5549
rect 1974 5544 1980 5545
rect 2374 5548 2380 5549
rect 2374 5544 2375 5548
rect 2379 5544 2380 5548
rect 2374 5543 2380 5544
rect 2606 5548 2612 5549
rect 2606 5544 2607 5548
rect 2611 5544 2612 5548
rect 2606 5543 2612 5544
rect 2830 5548 2836 5549
rect 2830 5544 2831 5548
rect 2835 5544 2836 5548
rect 2830 5543 2836 5544
rect 3046 5548 3052 5549
rect 3046 5544 3047 5548
rect 3051 5544 3052 5548
rect 3046 5543 3052 5544
rect 3262 5548 3268 5549
rect 3262 5544 3263 5548
rect 3267 5544 3268 5548
rect 3262 5543 3268 5544
rect 3478 5548 3484 5549
rect 3478 5544 3479 5548
rect 3483 5544 3484 5548
rect 3478 5543 3484 5544
rect 3678 5548 3684 5549
rect 3678 5544 3679 5548
rect 3683 5544 3684 5548
rect 3798 5545 3799 5549
rect 3803 5545 3804 5549
rect 3838 5549 3839 5553
rect 3843 5549 3844 5553
rect 3838 5548 3844 5549
rect 4430 5552 4436 5553
rect 4430 5548 4431 5552
rect 4435 5548 4436 5552
rect 4430 5547 4436 5548
rect 4566 5552 4572 5553
rect 4566 5548 4567 5552
rect 4571 5548 4572 5552
rect 4566 5547 4572 5548
rect 4702 5552 4708 5553
rect 4702 5548 4703 5552
rect 4707 5548 4708 5552
rect 4702 5547 4708 5548
rect 4838 5552 4844 5553
rect 4838 5548 4839 5552
rect 4843 5548 4844 5552
rect 4838 5547 4844 5548
rect 4974 5552 4980 5553
rect 4974 5548 4975 5552
rect 4979 5548 4980 5552
rect 4974 5547 4980 5548
rect 5110 5552 5116 5553
rect 5110 5548 5111 5552
rect 5115 5548 5116 5552
rect 5662 5549 5663 5553
rect 5667 5549 5668 5553
rect 5662 5548 5668 5549
rect 5110 5547 5116 5548
rect 3798 5544 3804 5545
rect 3678 5543 3684 5544
rect 4402 5537 4408 5538
rect 3838 5536 3844 5537
rect 2346 5533 2352 5534
rect 1974 5532 1980 5533
rect 1391 5531 1397 5532
rect 1391 5527 1392 5531
rect 1396 5530 1397 5531
rect 1846 5531 1852 5532
rect 1846 5530 1847 5531
rect 1396 5528 1847 5530
rect 1396 5527 1397 5528
rect 1391 5526 1397 5527
rect 1846 5527 1847 5528
rect 1851 5527 1852 5531
rect 1974 5528 1975 5532
rect 1979 5528 1980 5532
rect 2346 5529 2347 5533
rect 2351 5529 2352 5533
rect 2346 5528 2352 5529
rect 2578 5533 2584 5534
rect 2578 5529 2579 5533
rect 2583 5529 2584 5533
rect 2578 5528 2584 5529
rect 2802 5533 2808 5534
rect 2802 5529 2803 5533
rect 2807 5529 2808 5533
rect 2802 5528 2808 5529
rect 3018 5533 3024 5534
rect 3018 5529 3019 5533
rect 3023 5529 3024 5533
rect 3018 5528 3024 5529
rect 3234 5533 3240 5534
rect 3234 5529 3235 5533
rect 3239 5529 3240 5533
rect 3234 5528 3240 5529
rect 3450 5533 3456 5534
rect 3450 5529 3451 5533
rect 3455 5529 3456 5533
rect 3450 5528 3456 5529
rect 3650 5533 3656 5534
rect 3650 5529 3651 5533
rect 3655 5529 3656 5533
rect 3650 5528 3656 5529
rect 3798 5532 3804 5533
rect 3798 5528 3799 5532
rect 3803 5528 3804 5532
rect 3838 5532 3839 5536
rect 3843 5532 3844 5536
rect 4402 5533 4403 5537
rect 4407 5533 4408 5537
rect 4402 5532 4408 5533
rect 4538 5537 4544 5538
rect 4538 5533 4539 5537
rect 4543 5533 4544 5537
rect 4538 5532 4544 5533
rect 4674 5537 4680 5538
rect 4674 5533 4675 5537
rect 4679 5533 4680 5537
rect 4674 5532 4680 5533
rect 4810 5537 4816 5538
rect 4810 5533 4811 5537
rect 4815 5533 4816 5537
rect 4810 5532 4816 5533
rect 4946 5537 4952 5538
rect 4946 5533 4947 5537
rect 4951 5533 4952 5537
rect 4946 5532 4952 5533
rect 5082 5537 5088 5538
rect 5082 5533 5083 5537
rect 5087 5533 5088 5537
rect 5082 5532 5088 5533
rect 5662 5536 5668 5537
rect 5662 5532 5663 5536
rect 5667 5532 5668 5536
rect 3838 5531 3844 5532
rect 5662 5531 5668 5532
rect 1974 5527 1980 5528
rect 3798 5527 3804 5528
rect 4527 5527 4533 5528
rect 1846 5526 1852 5527
rect 2471 5523 2477 5524
rect 2471 5519 2472 5523
rect 2476 5522 2477 5523
rect 2594 5523 2600 5524
rect 2594 5522 2595 5523
rect 2476 5520 2595 5522
rect 2476 5519 2477 5520
rect 2471 5518 2477 5519
rect 2594 5519 2595 5520
rect 2599 5519 2600 5523
rect 2594 5518 2600 5519
rect 2650 5523 2656 5524
rect 2650 5519 2651 5523
rect 2655 5522 2656 5523
rect 2703 5523 2709 5524
rect 2703 5522 2704 5523
rect 2655 5520 2704 5522
rect 2655 5519 2656 5520
rect 2650 5518 2656 5519
rect 2703 5519 2704 5520
rect 2708 5519 2709 5523
rect 2703 5518 2709 5519
rect 2927 5523 2933 5524
rect 2927 5519 2928 5523
rect 2932 5522 2933 5523
rect 3034 5523 3040 5524
rect 3034 5522 3035 5523
rect 2932 5520 3035 5522
rect 2932 5519 2933 5520
rect 2927 5518 2933 5519
rect 3034 5519 3035 5520
rect 3039 5519 3040 5523
rect 3034 5518 3040 5519
rect 3066 5523 3072 5524
rect 3066 5519 3067 5523
rect 3071 5522 3072 5523
rect 3143 5523 3149 5524
rect 3143 5522 3144 5523
rect 3071 5520 3144 5522
rect 3071 5519 3072 5520
rect 3066 5518 3072 5519
rect 3143 5519 3144 5520
rect 3148 5519 3149 5523
rect 3143 5518 3149 5519
rect 3359 5523 3365 5524
rect 3359 5519 3360 5523
rect 3364 5522 3365 5523
rect 3466 5523 3472 5524
rect 3466 5522 3467 5523
rect 3364 5520 3467 5522
rect 3364 5519 3365 5520
rect 3359 5518 3365 5519
rect 3466 5519 3467 5520
rect 3471 5519 3472 5523
rect 3466 5518 3472 5519
rect 3575 5523 3584 5524
rect 3575 5519 3576 5523
rect 3583 5519 3584 5523
rect 3775 5523 3781 5524
rect 3775 5522 3776 5523
rect 3575 5518 3584 5519
rect 3588 5520 3776 5522
rect 3322 5515 3328 5516
rect 998 5511 1004 5512
rect 998 5510 999 5511
rect 965 5508 999 5510
rect 998 5507 999 5508
rect 1003 5507 1004 5511
rect 998 5506 1004 5507
rect 1007 5511 1013 5512
rect 1007 5507 1008 5511
rect 1012 5510 1013 5511
rect 1143 5511 1149 5512
rect 1012 5508 1029 5510
rect 1012 5507 1013 5508
rect 1007 5506 1013 5507
rect 1143 5507 1144 5511
rect 1148 5510 1149 5511
rect 1391 5511 1397 5512
rect 1391 5510 1392 5511
rect 1148 5508 1165 5510
rect 1381 5508 1392 5510
rect 1148 5507 1149 5508
rect 1143 5506 1149 5507
rect 1391 5507 1392 5508
rect 1396 5507 1397 5511
rect 1391 5506 1397 5507
rect 1418 5511 1424 5512
rect 1418 5507 1419 5511
rect 1423 5510 1424 5511
rect 1535 5511 1541 5512
rect 1423 5508 1453 5510
rect 1423 5507 1424 5508
rect 1418 5506 1424 5507
rect 1535 5507 1536 5511
rect 1540 5510 1541 5511
rect 1706 5511 1712 5512
rect 1540 5508 1597 5510
rect 1540 5507 1541 5508
rect 1535 5506 1541 5507
rect 1706 5507 1707 5511
rect 1711 5510 1712 5511
rect 3322 5511 3323 5515
rect 3327 5514 3328 5515
rect 3588 5514 3590 5520
rect 3775 5519 3776 5520
rect 3780 5519 3781 5523
rect 4527 5523 4528 5527
rect 4532 5526 4533 5527
rect 4554 5527 4560 5528
rect 4554 5526 4555 5527
rect 4532 5524 4555 5526
rect 4532 5523 4533 5524
rect 4527 5522 4533 5523
rect 4554 5523 4555 5524
rect 4559 5523 4560 5527
rect 4663 5527 4669 5528
rect 4663 5526 4664 5527
rect 4554 5522 4560 5523
rect 4564 5524 4664 5526
rect 3775 5518 3781 5519
rect 4490 5519 4496 5520
rect 4490 5515 4491 5519
rect 4495 5518 4496 5519
rect 4564 5518 4566 5524
rect 4663 5523 4664 5524
rect 4668 5523 4669 5527
rect 4663 5522 4669 5523
rect 4799 5527 4805 5528
rect 4799 5523 4800 5527
rect 4804 5526 4805 5527
rect 4826 5527 4832 5528
rect 4826 5526 4827 5527
rect 4804 5524 4827 5526
rect 4804 5523 4805 5524
rect 4799 5522 4805 5523
rect 4826 5523 4827 5524
rect 4831 5523 4832 5527
rect 4826 5522 4832 5523
rect 4935 5527 4941 5528
rect 4935 5523 4936 5527
rect 4940 5526 4941 5527
rect 4962 5527 4968 5528
rect 4962 5526 4963 5527
rect 4940 5524 4963 5526
rect 4940 5523 4941 5524
rect 4935 5522 4941 5523
rect 4962 5523 4963 5524
rect 4967 5523 4968 5527
rect 4962 5522 4968 5523
rect 5071 5527 5077 5528
rect 5071 5523 5072 5527
rect 5076 5526 5077 5527
rect 5098 5527 5104 5528
rect 5098 5526 5099 5527
rect 5076 5524 5099 5526
rect 5076 5523 5077 5524
rect 5071 5522 5077 5523
rect 5098 5523 5099 5524
rect 5103 5523 5104 5527
rect 5207 5527 5213 5528
rect 5207 5526 5208 5527
rect 5098 5522 5104 5523
rect 5108 5524 5208 5526
rect 4495 5516 4566 5518
rect 4886 5519 4892 5520
rect 4495 5515 4496 5516
rect 4490 5514 4496 5515
rect 4886 5515 4887 5519
rect 4891 5518 4892 5519
rect 5108 5518 5110 5524
rect 5207 5523 5208 5524
rect 5212 5523 5213 5527
rect 5207 5522 5213 5523
rect 4891 5516 5110 5518
rect 4891 5515 4892 5516
rect 4886 5514 4892 5515
rect 3327 5512 3590 5514
rect 3327 5511 3328 5512
rect 3322 5510 3328 5511
rect 4910 5511 4916 5512
rect 4910 5510 4911 5511
rect 1711 5508 1741 5510
rect 4768 5508 4911 5510
rect 1711 5507 1712 5508
rect 1706 5506 1712 5507
rect 4490 5495 4496 5496
rect 2434 5491 2440 5492
rect 2434 5487 2435 5491
rect 2439 5487 2440 5491
rect 2434 5486 2440 5487
rect 2594 5491 2600 5492
rect 2594 5487 2595 5491
rect 2599 5487 2600 5491
rect 2594 5486 2600 5487
rect 2822 5491 2828 5492
rect 2822 5487 2823 5491
rect 2827 5487 2828 5491
rect 2822 5486 2828 5487
rect 3034 5491 3040 5492
rect 3034 5487 3035 5491
rect 3039 5487 3040 5491
rect 3034 5486 3040 5487
rect 3322 5491 3328 5492
rect 3322 5487 3323 5491
rect 3327 5487 3328 5491
rect 3322 5486 3328 5487
rect 3466 5491 3472 5492
rect 3466 5487 3467 5491
rect 3471 5487 3472 5491
rect 3466 5486 3472 5487
rect 3738 5491 3744 5492
rect 3738 5487 3739 5491
rect 3743 5487 3744 5491
rect 4490 5491 4491 5495
rect 4495 5491 4496 5495
rect 4490 5490 4496 5491
rect 4626 5495 4632 5496
rect 4626 5491 4627 5495
rect 4631 5491 4632 5495
rect 4768 5494 4770 5508
rect 4910 5507 4911 5508
rect 4915 5507 4916 5511
rect 4910 5506 4916 5507
rect 4765 5492 4770 5494
rect 4826 5495 4832 5496
rect 4626 5490 4632 5491
rect 4826 5491 4827 5495
rect 4831 5491 4832 5495
rect 4826 5490 4832 5491
rect 4962 5495 4968 5496
rect 4962 5491 4963 5495
rect 4967 5491 4968 5495
rect 4962 5490 4968 5491
rect 5098 5495 5104 5496
rect 5098 5491 5099 5495
rect 5103 5491 5104 5495
rect 5098 5490 5104 5491
rect 3738 5486 3744 5487
rect 999 5475 1005 5476
rect 999 5471 1000 5475
rect 1004 5474 1005 5475
rect 1007 5475 1013 5476
rect 1007 5474 1008 5475
rect 1004 5472 1008 5474
rect 1004 5471 1005 5472
rect 999 5470 1005 5471
rect 1007 5471 1008 5472
rect 1012 5471 1013 5475
rect 1007 5470 1013 5471
rect 1135 5475 1141 5476
rect 1135 5471 1136 5475
rect 1140 5474 1141 5475
rect 1143 5475 1149 5476
rect 1143 5474 1144 5475
rect 1140 5472 1144 5474
rect 1140 5471 1141 5472
rect 1135 5470 1141 5471
rect 1143 5471 1144 5472
rect 1148 5471 1149 5475
rect 1143 5470 1149 5471
rect 1270 5475 1277 5476
rect 1270 5471 1271 5475
rect 1276 5471 1277 5475
rect 1270 5470 1277 5471
rect 1415 5475 1424 5476
rect 1415 5471 1416 5475
rect 1423 5471 1424 5475
rect 1415 5470 1424 5471
rect 1558 5475 1565 5476
rect 1558 5471 1559 5475
rect 1564 5471 1565 5475
rect 1558 5470 1565 5471
rect 1703 5475 1712 5476
rect 1703 5471 1704 5475
rect 1711 5471 1712 5475
rect 1703 5470 1712 5471
rect 1846 5475 1853 5476
rect 1846 5471 1847 5475
rect 1852 5471 1853 5475
rect 1846 5470 1853 5471
rect 110 5468 116 5469
rect 1934 5468 1940 5469
rect 110 5464 111 5468
rect 115 5464 116 5468
rect 110 5463 116 5464
rect 874 5467 880 5468
rect 874 5463 875 5467
rect 879 5463 880 5467
rect 874 5462 880 5463
rect 1010 5467 1016 5468
rect 1010 5463 1011 5467
rect 1015 5463 1016 5467
rect 1010 5462 1016 5463
rect 1146 5467 1152 5468
rect 1146 5463 1147 5467
rect 1151 5463 1152 5467
rect 1146 5462 1152 5463
rect 1290 5467 1296 5468
rect 1290 5463 1291 5467
rect 1295 5463 1296 5467
rect 1290 5462 1296 5463
rect 1434 5467 1440 5468
rect 1434 5463 1435 5467
rect 1439 5463 1440 5467
rect 1434 5462 1440 5463
rect 1578 5467 1584 5468
rect 1578 5463 1579 5467
rect 1583 5463 1584 5467
rect 1578 5462 1584 5463
rect 1722 5467 1728 5468
rect 1722 5463 1723 5467
rect 1727 5463 1728 5467
rect 1934 5464 1935 5468
rect 1939 5464 1940 5468
rect 1934 5463 1940 5464
rect 1722 5462 1728 5463
rect 902 5452 908 5453
rect 110 5451 116 5452
rect 110 5447 111 5451
rect 115 5447 116 5451
rect 902 5448 903 5452
rect 907 5448 908 5452
rect 902 5447 908 5448
rect 1038 5452 1044 5453
rect 1038 5448 1039 5452
rect 1043 5448 1044 5452
rect 1038 5447 1044 5448
rect 1174 5452 1180 5453
rect 1174 5448 1175 5452
rect 1179 5448 1180 5452
rect 1174 5447 1180 5448
rect 1318 5452 1324 5453
rect 1318 5448 1319 5452
rect 1323 5448 1324 5452
rect 1318 5447 1324 5448
rect 1462 5452 1468 5453
rect 1462 5448 1463 5452
rect 1467 5448 1468 5452
rect 1462 5447 1468 5448
rect 1606 5452 1612 5453
rect 1606 5448 1607 5452
rect 1611 5448 1612 5452
rect 1606 5447 1612 5448
rect 1750 5452 1756 5453
rect 1750 5448 1751 5452
rect 1755 5448 1756 5452
rect 1750 5447 1756 5448
rect 1934 5451 1940 5452
rect 1934 5447 1935 5451
rect 1939 5447 1940 5451
rect 110 5446 116 5447
rect 1934 5446 1940 5447
rect 4575 5447 4581 5448
rect 4514 5443 4520 5444
rect 2418 5439 2424 5440
rect 2418 5435 2419 5439
rect 2423 5438 2424 5439
rect 2894 5439 2900 5440
rect 2894 5438 2895 5439
rect 2423 5436 2469 5438
rect 2789 5436 2895 5438
rect 2423 5435 2424 5436
rect 2418 5434 2424 5435
rect 2894 5435 2895 5436
rect 2899 5435 2900 5439
rect 3314 5439 3320 5440
rect 2894 5434 2900 5435
rect 3034 5435 3040 5436
rect 3034 5431 3035 5435
rect 3039 5431 3040 5435
rect 3034 5430 3040 5431
rect 3274 5435 3280 5436
rect 3274 5431 3275 5435
rect 3279 5431 3280 5435
rect 3314 5435 3315 5439
rect 3319 5438 3320 5439
rect 3578 5439 3584 5440
rect 3319 5436 3445 5438
rect 3319 5435 3320 5436
rect 3314 5434 3320 5435
rect 3578 5435 3579 5439
rect 3583 5438 3584 5439
rect 4514 5439 4515 5443
rect 4519 5439 4520 5443
rect 4575 5443 4576 5447
rect 4580 5446 4581 5447
rect 4886 5447 4892 5448
rect 4886 5446 4887 5447
rect 4580 5444 4605 5446
rect 4837 5444 4887 5446
rect 4580 5443 4581 5444
rect 4575 5442 4581 5443
rect 4886 5443 4887 5444
rect 4891 5443 4892 5447
rect 4886 5442 4892 5443
rect 4895 5447 4901 5448
rect 4895 5443 4896 5447
rect 4900 5446 4901 5447
rect 5039 5447 5045 5448
rect 4900 5444 4925 5446
rect 4900 5443 4901 5444
rect 4895 5442 4901 5443
rect 5039 5443 5040 5447
rect 5044 5446 5045 5447
rect 5044 5444 5093 5446
rect 5044 5443 5045 5444
rect 5039 5442 5045 5443
rect 4514 5438 4520 5439
rect 3583 5436 3669 5438
rect 3583 5435 3584 5436
rect 3578 5434 3584 5435
rect 3274 5430 3280 5431
rect 3274 5415 3280 5416
rect 3274 5411 3275 5415
rect 3279 5414 3280 5415
rect 3279 5412 3682 5414
rect 3279 5411 3280 5412
rect 3274 5410 3280 5411
rect 2434 5403 2440 5404
rect 2434 5399 2435 5403
rect 2439 5402 2440 5403
rect 2575 5403 2581 5404
rect 2575 5402 2576 5403
rect 2439 5400 2576 5402
rect 2439 5399 2440 5400
rect 2434 5398 2440 5399
rect 2575 5399 2576 5400
rect 2580 5399 2581 5403
rect 2575 5398 2581 5399
rect 2822 5403 2829 5404
rect 2822 5399 2823 5403
rect 2828 5399 2829 5403
rect 2822 5398 2829 5399
rect 2894 5403 2900 5404
rect 2894 5399 2895 5403
rect 2899 5402 2900 5403
rect 3071 5403 3077 5404
rect 3071 5402 3072 5403
rect 2899 5400 3072 5402
rect 2899 5399 2900 5400
rect 2894 5398 2900 5399
rect 3071 5399 3072 5400
rect 3076 5399 3077 5403
rect 3071 5398 3077 5399
rect 3311 5403 3320 5404
rect 3311 5399 3312 5403
rect 3319 5399 3320 5403
rect 3311 5398 3320 5399
rect 3550 5403 3557 5404
rect 3550 5399 3551 5403
rect 3556 5399 3557 5403
rect 3680 5402 3682 5412
rect 4551 5411 4557 5412
rect 4551 5407 4552 5411
rect 4556 5410 4557 5411
rect 4575 5411 4581 5412
rect 4575 5410 4576 5411
rect 4556 5408 4576 5410
rect 4556 5407 4557 5408
rect 4551 5406 4557 5407
rect 4575 5407 4576 5408
rect 4580 5407 4581 5411
rect 4575 5406 4581 5407
rect 4626 5411 4632 5412
rect 4626 5407 4627 5411
rect 4631 5410 4632 5411
rect 4711 5411 4717 5412
rect 4711 5410 4712 5411
rect 4631 5408 4712 5410
rect 4631 5407 4632 5408
rect 4626 5406 4632 5407
rect 4711 5407 4712 5408
rect 4716 5407 4717 5411
rect 4711 5406 4717 5407
rect 4871 5411 4877 5412
rect 4871 5407 4872 5411
rect 4876 5410 4877 5411
rect 4895 5411 4901 5412
rect 4895 5410 4896 5411
rect 4876 5408 4896 5410
rect 4876 5407 4877 5408
rect 4871 5406 4877 5407
rect 4895 5407 4896 5408
rect 4900 5407 4901 5411
rect 4895 5406 4901 5407
rect 5031 5411 5037 5412
rect 5031 5407 5032 5411
rect 5036 5410 5037 5411
rect 5039 5411 5045 5412
rect 5039 5410 5040 5411
rect 5036 5408 5040 5410
rect 5036 5407 5037 5408
rect 5031 5406 5037 5407
rect 5039 5407 5040 5408
rect 5044 5407 5045 5411
rect 5039 5406 5045 5407
rect 5198 5411 5205 5412
rect 5198 5407 5199 5411
rect 5204 5407 5205 5411
rect 5198 5406 5205 5407
rect 3838 5404 3844 5405
rect 5662 5404 5668 5405
rect 3775 5403 3781 5404
rect 3775 5402 3776 5403
rect 3680 5400 3776 5402
rect 3550 5398 3557 5399
rect 3775 5399 3776 5400
rect 3780 5399 3781 5403
rect 3838 5400 3839 5404
rect 3843 5400 3844 5404
rect 3838 5399 3844 5400
rect 4426 5403 4432 5404
rect 4426 5399 4427 5403
rect 4431 5399 4432 5403
rect 3775 5398 3781 5399
rect 4426 5398 4432 5399
rect 4586 5403 4592 5404
rect 4586 5399 4587 5403
rect 4591 5399 4592 5403
rect 4586 5398 4592 5399
rect 4746 5403 4752 5404
rect 4746 5399 4747 5403
rect 4751 5399 4752 5403
rect 4746 5398 4752 5399
rect 4906 5403 4912 5404
rect 4906 5399 4907 5403
rect 4911 5399 4912 5403
rect 4906 5398 4912 5399
rect 5074 5403 5080 5404
rect 5074 5399 5075 5403
rect 5079 5399 5080 5403
rect 5662 5400 5663 5404
rect 5667 5400 5668 5404
rect 5662 5399 5668 5400
rect 5074 5398 5080 5399
rect 1974 5396 1980 5397
rect 3798 5396 3804 5397
rect 110 5393 116 5394
rect 1934 5393 1940 5394
rect 110 5389 111 5393
rect 115 5389 116 5393
rect 110 5388 116 5389
rect 718 5392 724 5393
rect 718 5388 719 5392
rect 723 5388 724 5392
rect 718 5387 724 5388
rect 854 5392 860 5393
rect 854 5388 855 5392
rect 859 5388 860 5392
rect 854 5387 860 5388
rect 990 5392 996 5393
rect 990 5388 991 5392
rect 995 5388 996 5392
rect 990 5387 996 5388
rect 1126 5392 1132 5393
rect 1126 5388 1127 5392
rect 1131 5388 1132 5392
rect 1126 5387 1132 5388
rect 1262 5392 1268 5393
rect 1262 5388 1263 5392
rect 1267 5388 1268 5392
rect 1262 5387 1268 5388
rect 1398 5392 1404 5393
rect 1398 5388 1399 5392
rect 1403 5388 1404 5392
rect 1398 5387 1404 5388
rect 1534 5392 1540 5393
rect 1534 5388 1535 5392
rect 1539 5388 1540 5392
rect 1534 5387 1540 5388
rect 1670 5392 1676 5393
rect 1670 5388 1671 5392
rect 1675 5388 1676 5392
rect 1670 5387 1676 5388
rect 1806 5392 1812 5393
rect 1806 5388 1807 5392
rect 1811 5388 1812 5392
rect 1934 5389 1935 5393
rect 1939 5389 1940 5393
rect 1974 5392 1975 5396
rect 1979 5392 1980 5396
rect 1974 5391 1980 5392
rect 2450 5395 2456 5396
rect 2450 5391 2451 5395
rect 2455 5391 2456 5395
rect 2450 5390 2456 5391
rect 2698 5395 2704 5396
rect 2698 5391 2699 5395
rect 2703 5391 2704 5395
rect 2698 5390 2704 5391
rect 2946 5395 2952 5396
rect 2946 5391 2947 5395
rect 2951 5391 2952 5395
rect 2946 5390 2952 5391
rect 3186 5395 3192 5396
rect 3186 5391 3187 5395
rect 3191 5391 3192 5395
rect 3186 5390 3192 5391
rect 3426 5395 3432 5396
rect 3426 5391 3427 5395
rect 3431 5391 3432 5395
rect 3426 5390 3432 5391
rect 3650 5395 3656 5396
rect 3650 5391 3651 5395
rect 3655 5391 3656 5395
rect 3798 5392 3799 5396
rect 3803 5392 3804 5396
rect 3798 5391 3804 5392
rect 3650 5390 3656 5391
rect 1934 5388 1940 5389
rect 4454 5388 4460 5389
rect 1806 5387 1812 5388
rect 3838 5387 3844 5388
rect 3838 5383 3839 5387
rect 3843 5383 3844 5387
rect 4454 5384 4455 5388
rect 4459 5384 4460 5388
rect 4454 5383 4460 5384
rect 4614 5388 4620 5389
rect 4614 5384 4615 5388
rect 4619 5384 4620 5388
rect 4614 5383 4620 5384
rect 4774 5388 4780 5389
rect 4774 5384 4775 5388
rect 4779 5384 4780 5388
rect 4774 5383 4780 5384
rect 4934 5388 4940 5389
rect 4934 5384 4935 5388
rect 4939 5384 4940 5388
rect 4934 5383 4940 5384
rect 5102 5388 5108 5389
rect 5102 5384 5103 5388
rect 5107 5384 5108 5388
rect 5102 5383 5108 5384
rect 5662 5387 5668 5388
rect 5662 5383 5663 5387
rect 5667 5383 5668 5387
rect 3838 5382 3844 5383
rect 5662 5382 5668 5383
rect 2478 5380 2484 5381
rect 1974 5379 1980 5380
rect 690 5377 696 5378
rect 110 5376 116 5377
rect 110 5372 111 5376
rect 115 5372 116 5376
rect 690 5373 691 5377
rect 695 5373 696 5377
rect 690 5372 696 5373
rect 826 5377 832 5378
rect 826 5373 827 5377
rect 831 5373 832 5377
rect 826 5372 832 5373
rect 962 5377 968 5378
rect 962 5373 963 5377
rect 967 5373 968 5377
rect 962 5372 968 5373
rect 1098 5377 1104 5378
rect 1098 5373 1099 5377
rect 1103 5373 1104 5377
rect 1098 5372 1104 5373
rect 1234 5377 1240 5378
rect 1234 5373 1235 5377
rect 1239 5373 1240 5377
rect 1234 5372 1240 5373
rect 1370 5377 1376 5378
rect 1370 5373 1371 5377
rect 1375 5373 1376 5377
rect 1370 5372 1376 5373
rect 1506 5377 1512 5378
rect 1506 5373 1507 5377
rect 1511 5373 1512 5377
rect 1506 5372 1512 5373
rect 1642 5377 1648 5378
rect 1642 5373 1643 5377
rect 1647 5373 1648 5377
rect 1642 5372 1648 5373
rect 1778 5377 1784 5378
rect 1778 5373 1779 5377
rect 1783 5373 1784 5377
rect 1778 5372 1784 5373
rect 1934 5376 1940 5377
rect 1934 5372 1935 5376
rect 1939 5372 1940 5376
rect 1974 5375 1975 5379
rect 1979 5375 1980 5379
rect 2478 5376 2479 5380
rect 2483 5376 2484 5380
rect 2478 5375 2484 5376
rect 2726 5380 2732 5381
rect 2726 5376 2727 5380
rect 2731 5376 2732 5380
rect 2726 5375 2732 5376
rect 2974 5380 2980 5381
rect 2974 5376 2975 5380
rect 2979 5376 2980 5380
rect 2974 5375 2980 5376
rect 3214 5380 3220 5381
rect 3214 5376 3215 5380
rect 3219 5376 3220 5380
rect 3214 5375 3220 5376
rect 3454 5380 3460 5381
rect 3454 5376 3455 5380
rect 3459 5376 3460 5380
rect 3454 5375 3460 5376
rect 3678 5380 3684 5381
rect 3678 5376 3679 5380
rect 3683 5376 3684 5380
rect 3678 5375 3684 5376
rect 3798 5379 3804 5380
rect 3798 5375 3799 5379
rect 3803 5375 3804 5379
rect 1974 5374 1980 5375
rect 3798 5374 3804 5375
rect 110 5371 116 5372
rect 1934 5371 1940 5372
rect 810 5367 821 5368
rect 810 5363 811 5367
rect 815 5363 816 5367
rect 820 5363 821 5367
rect 810 5362 821 5363
rect 823 5367 829 5368
rect 823 5363 824 5367
rect 828 5366 829 5367
rect 951 5367 957 5368
rect 951 5366 952 5367
rect 828 5364 952 5366
rect 828 5363 829 5364
rect 823 5362 829 5363
rect 951 5363 952 5364
rect 956 5363 957 5367
rect 951 5362 957 5363
rect 959 5367 965 5368
rect 959 5363 960 5367
rect 964 5366 965 5367
rect 1087 5367 1093 5368
rect 1087 5366 1088 5367
rect 964 5364 1088 5366
rect 964 5363 965 5364
rect 959 5362 965 5363
rect 1087 5363 1088 5364
rect 1092 5363 1093 5367
rect 1087 5362 1093 5363
rect 1095 5367 1101 5368
rect 1095 5363 1096 5367
rect 1100 5366 1101 5367
rect 1223 5367 1229 5368
rect 1223 5366 1224 5367
rect 1100 5364 1224 5366
rect 1100 5363 1101 5364
rect 1095 5362 1101 5363
rect 1223 5363 1224 5364
rect 1228 5363 1229 5367
rect 1223 5362 1229 5363
rect 1359 5367 1365 5368
rect 1359 5363 1360 5367
rect 1364 5366 1365 5367
rect 1386 5367 1392 5368
rect 1386 5366 1387 5367
rect 1364 5364 1387 5366
rect 1364 5363 1365 5364
rect 1359 5362 1365 5363
rect 1386 5363 1387 5364
rect 1391 5363 1392 5367
rect 1386 5362 1392 5363
rect 1474 5367 1480 5368
rect 1474 5363 1475 5367
rect 1479 5366 1480 5367
rect 1495 5367 1501 5368
rect 1495 5366 1496 5367
rect 1479 5364 1496 5366
rect 1479 5363 1480 5364
rect 1474 5362 1480 5363
rect 1495 5363 1496 5364
rect 1500 5363 1501 5367
rect 1495 5362 1501 5363
rect 1631 5367 1637 5368
rect 1631 5363 1632 5367
rect 1636 5366 1637 5367
rect 1658 5367 1664 5368
rect 1658 5366 1659 5367
rect 1636 5364 1659 5366
rect 1636 5363 1637 5364
rect 1631 5362 1637 5363
rect 1658 5363 1659 5364
rect 1663 5363 1664 5367
rect 1658 5362 1664 5363
rect 1767 5367 1773 5368
rect 1767 5363 1768 5367
rect 1772 5366 1773 5367
rect 1794 5367 1800 5368
rect 1794 5366 1795 5367
rect 1772 5364 1795 5366
rect 1772 5363 1773 5364
rect 1767 5362 1773 5363
rect 1794 5363 1795 5364
rect 1799 5363 1800 5367
rect 1903 5367 1909 5368
rect 1903 5366 1904 5367
rect 1794 5362 1800 5363
rect 1804 5364 1904 5366
rect 1186 5355 1192 5356
rect 1186 5351 1187 5355
rect 1191 5354 1192 5355
rect 1804 5354 1806 5364
rect 1903 5363 1904 5364
rect 1908 5363 1909 5367
rect 1903 5362 1909 5363
rect 1191 5352 1806 5354
rect 1191 5351 1192 5352
rect 1186 5350 1192 5351
rect 823 5335 829 5336
rect 823 5334 824 5335
rect 781 5332 824 5334
rect 823 5331 824 5332
rect 828 5331 829 5335
rect 959 5335 965 5336
rect 959 5334 960 5335
rect 917 5332 960 5334
rect 823 5330 829 5331
rect 959 5331 960 5332
rect 964 5331 965 5335
rect 1095 5335 1101 5336
rect 1095 5334 1096 5335
rect 1053 5332 1096 5334
rect 959 5330 965 5331
rect 1095 5331 1096 5332
rect 1100 5331 1101 5335
rect 1095 5330 1101 5331
rect 1186 5335 1192 5336
rect 1186 5331 1187 5335
rect 1191 5331 1192 5335
rect 1186 5330 1192 5331
rect 1270 5335 1276 5336
rect 1270 5331 1271 5335
rect 1275 5331 1276 5335
rect 1270 5330 1276 5331
rect 1386 5335 1392 5336
rect 1386 5331 1387 5335
rect 1391 5331 1392 5335
rect 1386 5330 1392 5331
rect 1558 5335 1564 5336
rect 1558 5331 1559 5335
rect 1563 5331 1564 5335
rect 1558 5330 1564 5331
rect 1658 5335 1664 5336
rect 1658 5331 1659 5335
rect 1663 5331 1664 5335
rect 1658 5330 1664 5331
rect 1794 5335 1800 5336
rect 1794 5331 1795 5335
rect 1799 5331 1800 5335
rect 1794 5330 1800 5331
rect 1974 5321 1980 5322
rect 3798 5321 3804 5322
rect 1974 5317 1975 5321
rect 1979 5317 1980 5321
rect 1974 5316 1980 5317
rect 2318 5320 2324 5321
rect 2318 5316 2319 5320
rect 2323 5316 2324 5320
rect 2318 5315 2324 5316
rect 2518 5320 2524 5321
rect 2518 5316 2519 5320
rect 2523 5316 2524 5320
rect 2518 5315 2524 5316
rect 2718 5320 2724 5321
rect 2718 5316 2719 5320
rect 2723 5316 2724 5320
rect 2718 5315 2724 5316
rect 2918 5320 2924 5321
rect 2918 5316 2919 5320
rect 2923 5316 2924 5320
rect 2918 5315 2924 5316
rect 3118 5320 3124 5321
rect 3118 5316 3119 5320
rect 3123 5316 3124 5320
rect 3118 5315 3124 5316
rect 3326 5320 3332 5321
rect 3326 5316 3327 5320
rect 3331 5316 3332 5320
rect 3326 5315 3332 5316
rect 3534 5320 3540 5321
rect 3534 5316 3535 5320
rect 3539 5316 3540 5320
rect 3798 5317 3799 5321
rect 3803 5317 3804 5321
rect 3798 5316 3804 5317
rect 3838 5321 3844 5322
rect 5662 5321 5668 5322
rect 3838 5317 3839 5321
rect 3843 5317 3844 5321
rect 3838 5316 3844 5317
rect 4430 5320 4436 5321
rect 4430 5316 4431 5320
rect 4435 5316 4436 5320
rect 3534 5315 3540 5316
rect 4430 5315 4436 5316
rect 4614 5320 4620 5321
rect 4614 5316 4615 5320
rect 4619 5316 4620 5320
rect 4614 5315 4620 5316
rect 4798 5320 4804 5321
rect 4798 5316 4799 5320
rect 4803 5316 4804 5320
rect 4798 5315 4804 5316
rect 4982 5320 4988 5321
rect 4982 5316 4983 5320
rect 4987 5316 4988 5320
rect 4982 5315 4988 5316
rect 5174 5320 5180 5321
rect 5174 5316 5175 5320
rect 5179 5316 5180 5320
rect 5662 5317 5663 5321
rect 5667 5317 5668 5321
rect 5662 5316 5668 5317
rect 5174 5315 5180 5316
rect 2290 5305 2296 5306
rect 1974 5304 1980 5305
rect 1974 5300 1975 5304
rect 1979 5300 1980 5304
rect 2290 5301 2291 5305
rect 2295 5301 2296 5305
rect 2290 5300 2296 5301
rect 2490 5305 2496 5306
rect 2490 5301 2491 5305
rect 2495 5301 2496 5305
rect 2490 5300 2496 5301
rect 2690 5305 2696 5306
rect 2690 5301 2691 5305
rect 2695 5301 2696 5305
rect 2690 5300 2696 5301
rect 2890 5305 2896 5306
rect 2890 5301 2891 5305
rect 2895 5301 2896 5305
rect 2890 5300 2896 5301
rect 3090 5305 3096 5306
rect 3090 5301 3091 5305
rect 3095 5301 3096 5305
rect 3090 5300 3096 5301
rect 3298 5305 3304 5306
rect 3298 5301 3299 5305
rect 3303 5301 3304 5305
rect 3298 5300 3304 5301
rect 3506 5305 3512 5306
rect 4402 5305 4408 5306
rect 3506 5301 3507 5305
rect 3511 5301 3512 5305
rect 3506 5300 3512 5301
rect 3798 5304 3804 5305
rect 3798 5300 3799 5304
rect 3803 5300 3804 5304
rect 1974 5299 1980 5300
rect 3798 5299 3804 5300
rect 3838 5304 3844 5305
rect 3838 5300 3839 5304
rect 3843 5300 3844 5304
rect 4402 5301 4403 5305
rect 4407 5301 4408 5305
rect 4402 5300 4408 5301
rect 4586 5305 4592 5306
rect 4586 5301 4587 5305
rect 4591 5301 4592 5305
rect 4586 5300 4592 5301
rect 4770 5305 4776 5306
rect 4770 5301 4771 5305
rect 4775 5301 4776 5305
rect 4770 5300 4776 5301
rect 4954 5305 4960 5306
rect 4954 5301 4955 5305
rect 4959 5301 4960 5305
rect 4954 5300 4960 5301
rect 5146 5305 5152 5306
rect 5146 5301 5147 5305
rect 5151 5301 5152 5305
rect 5146 5300 5152 5301
rect 5662 5304 5668 5305
rect 5662 5300 5663 5304
rect 5667 5300 5668 5304
rect 3838 5299 3844 5300
rect 5662 5299 5668 5300
rect 2415 5295 2424 5296
rect 2415 5291 2416 5295
rect 2423 5291 2424 5295
rect 2415 5290 2424 5291
rect 2615 5295 2621 5296
rect 2615 5291 2616 5295
rect 2620 5294 2621 5295
rect 2706 5295 2712 5296
rect 2706 5294 2707 5295
rect 2620 5292 2707 5294
rect 2620 5291 2621 5292
rect 2615 5290 2621 5291
rect 2706 5291 2707 5292
rect 2711 5291 2712 5295
rect 2815 5295 2821 5296
rect 2815 5294 2816 5295
rect 2706 5290 2712 5291
rect 2716 5292 2816 5294
rect 850 5287 856 5288
rect 810 5283 816 5284
rect 810 5279 811 5283
rect 815 5279 816 5283
rect 850 5283 851 5287
rect 855 5286 856 5287
rect 1002 5287 1008 5288
rect 855 5284 893 5286
rect 855 5283 856 5284
rect 850 5282 856 5283
rect 1002 5283 1003 5287
rect 1007 5286 1008 5287
rect 1154 5287 1160 5288
rect 1007 5284 1045 5286
rect 1007 5283 1008 5284
rect 1002 5282 1008 5283
rect 1154 5283 1155 5287
rect 1159 5286 1160 5287
rect 1474 5287 1480 5288
rect 1474 5286 1475 5287
rect 1159 5284 1205 5286
rect 1445 5284 1475 5286
rect 1159 5283 1160 5284
rect 1154 5282 1160 5283
rect 1474 5283 1475 5284
rect 1479 5283 1480 5287
rect 1474 5282 1480 5283
rect 1487 5287 1493 5288
rect 1487 5283 1488 5287
rect 1492 5286 1493 5287
rect 2378 5287 2384 5288
rect 1492 5284 1541 5286
rect 1492 5283 1493 5284
rect 1487 5282 1493 5283
rect 2378 5283 2379 5287
rect 2383 5286 2384 5287
rect 2716 5286 2718 5292
rect 2815 5291 2816 5292
rect 2820 5291 2821 5295
rect 2815 5290 2821 5291
rect 3015 5295 3021 5296
rect 3015 5291 3016 5295
rect 3020 5294 3021 5295
rect 3034 5295 3040 5296
rect 3034 5294 3035 5295
rect 3020 5292 3035 5294
rect 3020 5291 3021 5292
rect 3015 5290 3021 5291
rect 3034 5291 3035 5292
rect 3039 5291 3040 5295
rect 3034 5290 3040 5291
rect 3215 5295 3221 5296
rect 3215 5291 3216 5295
rect 3220 5294 3221 5295
rect 3314 5295 3320 5296
rect 3314 5294 3315 5295
rect 3220 5292 3315 5294
rect 3220 5291 3221 5292
rect 3215 5290 3221 5291
rect 3314 5291 3315 5292
rect 3319 5291 3320 5295
rect 3314 5290 3320 5291
rect 3410 5295 3416 5296
rect 3410 5291 3411 5295
rect 3415 5294 3416 5295
rect 3423 5295 3429 5296
rect 3423 5294 3424 5295
rect 3415 5292 3424 5294
rect 3415 5291 3416 5292
rect 3410 5290 3416 5291
rect 3423 5291 3424 5292
rect 3428 5291 3429 5295
rect 3631 5295 3637 5296
rect 3631 5294 3632 5295
rect 3423 5290 3429 5291
rect 3432 5292 3632 5294
rect 2383 5284 2718 5286
rect 3178 5287 3184 5288
rect 2383 5283 2384 5284
rect 2378 5282 2384 5283
rect 3178 5283 3179 5287
rect 3183 5286 3184 5287
rect 3432 5286 3434 5292
rect 3631 5291 3632 5292
rect 3636 5291 3637 5295
rect 3631 5290 3637 5291
rect 4514 5295 4520 5296
rect 4514 5291 4515 5295
rect 4519 5294 4520 5295
rect 4527 5295 4533 5296
rect 4527 5294 4528 5295
rect 4519 5292 4528 5294
rect 4519 5291 4520 5292
rect 4514 5290 4520 5291
rect 4527 5291 4528 5292
rect 4532 5291 4533 5295
rect 4527 5290 4533 5291
rect 4566 5295 4572 5296
rect 4566 5291 4567 5295
rect 4571 5294 4572 5295
rect 4711 5295 4717 5296
rect 4711 5294 4712 5295
rect 4571 5292 4712 5294
rect 4571 5291 4572 5292
rect 4566 5290 4572 5291
rect 4711 5291 4712 5292
rect 4716 5291 4717 5295
rect 4711 5290 4717 5291
rect 4719 5295 4725 5296
rect 4719 5291 4720 5295
rect 4724 5294 4725 5295
rect 4895 5295 4901 5296
rect 4895 5294 4896 5295
rect 4724 5292 4896 5294
rect 4724 5291 4725 5292
rect 4719 5290 4725 5291
rect 4895 5291 4896 5292
rect 4900 5291 4901 5295
rect 4895 5290 4901 5291
rect 4946 5295 4952 5296
rect 4946 5291 4947 5295
rect 4951 5294 4952 5295
rect 5079 5295 5085 5296
rect 5079 5294 5080 5295
rect 4951 5292 5080 5294
rect 4951 5291 4952 5292
rect 4946 5290 4952 5291
rect 5079 5291 5080 5292
rect 5084 5291 5085 5295
rect 5079 5290 5085 5291
rect 5119 5295 5125 5296
rect 5119 5291 5120 5295
rect 5124 5294 5125 5295
rect 5271 5295 5277 5296
rect 5271 5294 5272 5295
rect 5124 5292 5272 5294
rect 5124 5291 5125 5292
rect 5119 5290 5125 5291
rect 5271 5291 5272 5292
rect 5276 5291 5277 5295
rect 5271 5290 5277 5291
rect 3183 5284 3434 5286
rect 3183 5283 3184 5284
rect 3178 5282 3184 5283
rect 810 5278 816 5279
rect 2378 5263 2384 5264
rect 2378 5259 2379 5263
rect 2383 5259 2384 5263
rect 2378 5258 2384 5259
rect 2578 5263 2584 5264
rect 2578 5259 2579 5263
rect 2583 5259 2584 5263
rect 2578 5258 2584 5259
rect 2706 5263 2712 5264
rect 2706 5259 2707 5263
rect 2711 5259 2712 5263
rect 2706 5258 2712 5259
rect 2978 5263 2984 5264
rect 2978 5259 2979 5263
rect 2983 5259 2984 5263
rect 2978 5258 2984 5259
rect 3178 5263 3184 5264
rect 3178 5259 3179 5263
rect 3183 5259 3184 5263
rect 3178 5258 3184 5259
rect 3314 5263 3320 5264
rect 3314 5259 3315 5263
rect 3319 5259 3320 5263
rect 3314 5258 3320 5259
rect 3550 5263 3556 5264
rect 3550 5259 3551 5263
rect 3555 5259 3556 5263
rect 4566 5263 4572 5264
rect 4566 5262 4567 5263
rect 4493 5260 4567 5262
rect 3550 5258 3556 5259
rect 4566 5259 4567 5260
rect 4571 5259 4572 5263
rect 4566 5258 4572 5259
rect 4602 5263 4608 5264
rect 4602 5259 4603 5263
rect 4607 5259 4608 5263
rect 4946 5263 4952 5264
rect 4946 5262 4947 5263
rect 4861 5260 4947 5262
rect 4602 5258 4608 5259
rect 4946 5259 4947 5260
rect 4951 5259 4952 5263
rect 5119 5263 5125 5264
rect 5119 5262 5120 5263
rect 5045 5260 5120 5262
rect 4946 5258 4952 5259
rect 5119 5259 5120 5260
rect 5124 5259 5125 5263
rect 5119 5258 5125 5259
rect 5198 5263 5204 5264
rect 5198 5259 5199 5263
rect 5203 5259 5204 5263
rect 5198 5258 5204 5259
rect 847 5251 856 5252
rect 847 5247 848 5251
rect 855 5247 856 5251
rect 847 5246 856 5247
rect 999 5251 1008 5252
rect 999 5247 1000 5251
rect 1007 5247 1008 5251
rect 999 5246 1008 5247
rect 1151 5251 1160 5252
rect 1151 5247 1152 5251
rect 1159 5247 1160 5251
rect 1151 5246 1160 5247
rect 1258 5251 1264 5252
rect 1258 5247 1259 5251
rect 1263 5250 1264 5251
rect 1311 5251 1317 5252
rect 1311 5250 1312 5251
rect 1263 5248 1312 5250
rect 1263 5247 1264 5248
rect 1258 5246 1264 5247
rect 1311 5247 1312 5248
rect 1316 5247 1317 5251
rect 1311 5246 1317 5247
rect 1479 5251 1485 5252
rect 1479 5247 1480 5251
rect 1484 5250 1485 5251
rect 1487 5251 1493 5252
rect 1487 5250 1488 5251
rect 1484 5248 1488 5250
rect 1484 5247 1485 5248
rect 1479 5246 1485 5247
rect 1487 5247 1488 5248
rect 1492 5247 1493 5251
rect 1487 5246 1493 5247
rect 1646 5251 1653 5252
rect 1646 5247 1647 5251
rect 1652 5247 1653 5251
rect 1646 5246 1653 5247
rect 110 5244 116 5245
rect 1934 5244 1940 5245
rect 110 5240 111 5244
rect 115 5240 116 5244
rect 110 5239 116 5240
rect 722 5243 728 5244
rect 722 5239 723 5243
rect 727 5239 728 5243
rect 722 5238 728 5239
rect 874 5243 880 5244
rect 874 5239 875 5243
rect 879 5239 880 5243
rect 874 5238 880 5239
rect 1026 5243 1032 5244
rect 1026 5239 1027 5243
rect 1031 5239 1032 5243
rect 1026 5238 1032 5239
rect 1186 5243 1192 5244
rect 1186 5239 1187 5243
rect 1191 5239 1192 5243
rect 1186 5238 1192 5239
rect 1354 5243 1360 5244
rect 1354 5239 1355 5243
rect 1359 5239 1360 5243
rect 1354 5238 1360 5239
rect 1522 5243 1528 5244
rect 1522 5239 1523 5243
rect 1527 5239 1528 5243
rect 1934 5240 1935 5244
rect 1939 5240 1940 5244
rect 1934 5239 1940 5240
rect 1522 5238 1528 5239
rect 750 5228 756 5229
rect 110 5227 116 5228
rect 110 5223 111 5227
rect 115 5223 116 5227
rect 750 5224 751 5228
rect 755 5224 756 5228
rect 750 5223 756 5224
rect 902 5228 908 5229
rect 902 5224 903 5228
rect 907 5224 908 5228
rect 902 5223 908 5224
rect 1054 5228 1060 5229
rect 1054 5224 1055 5228
rect 1059 5224 1060 5228
rect 1054 5223 1060 5224
rect 1214 5228 1220 5229
rect 1214 5224 1215 5228
rect 1219 5224 1220 5228
rect 1214 5223 1220 5224
rect 1382 5228 1388 5229
rect 1382 5224 1383 5228
rect 1387 5224 1388 5228
rect 1382 5223 1388 5224
rect 1550 5228 1556 5229
rect 1550 5224 1551 5228
rect 1555 5224 1556 5228
rect 1550 5223 1556 5224
rect 1934 5227 1940 5228
rect 1934 5223 1935 5227
rect 1939 5223 1940 5227
rect 110 5222 116 5223
rect 1934 5222 1940 5223
rect 2402 5211 2408 5212
rect 2362 5207 2368 5208
rect 2362 5203 2363 5207
rect 2367 5203 2368 5207
rect 2402 5207 2403 5211
rect 2407 5210 2408 5211
rect 2810 5211 2816 5212
rect 2407 5208 2493 5210
rect 2407 5207 2408 5208
rect 2402 5206 2408 5207
rect 2770 5207 2776 5208
rect 2362 5202 2368 5203
rect 2770 5203 2771 5207
rect 2775 5203 2776 5207
rect 2810 5207 2811 5211
rect 2815 5210 2816 5211
rect 3303 5211 3309 5212
rect 3303 5210 3304 5211
rect 2815 5208 2909 5210
rect 3189 5208 3304 5210
rect 2815 5207 2816 5208
rect 2810 5206 2816 5207
rect 3303 5207 3304 5208
rect 3308 5207 3309 5211
rect 3410 5211 3416 5212
rect 3410 5210 3411 5211
rect 3397 5208 3411 5210
rect 3303 5206 3309 5207
rect 3410 5207 3411 5208
rect 3415 5207 3416 5211
rect 3410 5206 3416 5207
rect 2770 5202 2776 5203
rect 4426 5199 4432 5200
rect 4426 5195 4427 5199
rect 4431 5198 4432 5199
rect 4719 5199 4725 5200
rect 4719 5198 4720 5199
rect 4431 5196 4453 5198
rect 4685 5196 4720 5198
rect 4431 5195 4432 5196
rect 4426 5194 4432 5195
rect 4719 5195 4720 5196
rect 4724 5195 4725 5199
rect 4719 5194 4725 5195
rect 4743 5199 4749 5200
rect 4743 5195 4744 5199
rect 4748 5198 4749 5199
rect 4903 5199 4909 5200
rect 4748 5196 4773 5198
rect 4748 5195 4749 5196
rect 4743 5194 4749 5195
rect 4903 5195 4904 5199
rect 4908 5198 4909 5199
rect 5047 5199 5053 5200
rect 4908 5196 4933 5198
rect 4908 5195 4909 5196
rect 4903 5194 4909 5195
rect 5047 5195 5048 5199
rect 5052 5198 5053 5199
rect 5199 5199 5205 5200
rect 5052 5196 5085 5198
rect 5052 5195 5053 5196
rect 5047 5194 5053 5195
rect 5199 5195 5200 5199
rect 5204 5198 5205 5199
rect 5367 5199 5373 5200
rect 5204 5196 5237 5198
rect 5204 5195 5205 5196
rect 5199 5194 5205 5195
rect 5367 5195 5368 5199
rect 5372 5198 5373 5199
rect 5511 5199 5517 5200
rect 5372 5196 5397 5198
rect 5372 5195 5373 5196
rect 5367 5194 5373 5195
rect 5511 5195 5512 5199
rect 5516 5198 5517 5199
rect 5516 5196 5533 5198
rect 5516 5195 5517 5196
rect 5511 5194 5517 5195
rect 2399 5175 2408 5176
rect 2399 5171 2400 5175
rect 2407 5171 2408 5175
rect 2399 5170 2408 5171
rect 2578 5175 2584 5176
rect 2578 5171 2579 5175
rect 2583 5174 2584 5175
rect 2599 5175 2605 5176
rect 2599 5174 2600 5175
rect 2583 5172 2600 5174
rect 2583 5171 2584 5172
rect 2578 5170 2584 5171
rect 2599 5171 2600 5172
rect 2604 5171 2605 5175
rect 2599 5170 2605 5171
rect 2807 5175 2816 5176
rect 2807 5171 2808 5175
rect 2815 5171 2816 5175
rect 2807 5170 2816 5171
rect 2978 5175 2984 5176
rect 2978 5171 2979 5175
rect 2983 5174 2984 5175
rect 3015 5175 3021 5176
rect 3015 5174 3016 5175
rect 2983 5172 3016 5174
rect 2983 5171 2984 5172
rect 2978 5170 2984 5171
rect 3015 5171 3016 5172
rect 3020 5171 3021 5175
rect 3015 5170 3021 5171
rect 3078 5175 3084 5176
rect 3078 5171 3079 5175
rect 3083 5174 3084 5175
rect 3223 5175 3229 5176
rect 3223 5174 3224 5175
rect 3083 5172 3224 5174
rect 3083 5171 3084 5172
rect 3078 5170 3084 5171
rect 3223 5171 3224 5172
rect 3228 5171 3229 5175
rect 3223 5170 3229 5171
rect 3303 5175 3309 5176
rect 3303 5171 3304 5175
rect 3308 5174 3309 5175
rect 3431 5175 3437 5176
rect 3431 5174 3432 5175
rect 3308 5172 3432 5174
rect 3308 5171 3309 5172
rect 3303 5170 3309 5171
rect 3431 5171 3432 5172
rect 3436 5171 3437 5175
rect 3431 5170 3437 5171
rect 110 5169 116 5170
rect 1934 5169 1940 5170
rect 110 5165 111 5169
rect 115 5165 116 5169
rect 110 5164 116 5165
rect 446 5168 452 5169
rect 446 5164 447 5168
rect 451 5164 452 5168
rect 446 5163 452 5164
rect 622 5168 628 5169
rect 622 5164 623 5168
rect 627 5164 628 5168
rect 622 5163 628 5164
rect 806 5168 812 5169
rect 806 5164 807 5168
rect 811 5164 812 5168
rect 806 5163 812 5164
rect 998 5168 1004 5169
rect 998 5164 999 5168
rect 1003 5164 1004 5168
rect 998 5163 1004 5164
rect 1198 5168 1204 5169
rect 1198 5164 1199 5168
rect 1203 5164 1204 5168
rect 1198 5163 1204 5164
rect 1398 5168 1404 5169
rect 1398 5164 1399 5168
rect 1403 5164 1404 5168
rect 1398 5163 1404 5164
rect 1606 5168 1612 5169
rect 1606 5164 1607 5168
rect 1611 5164 1612 5168
rect 1606 5163 1612 5164
rect 1814 5168 1820 5169
rect 1814 5164 1815 5168
rect 1819 5164 1820 5168
rect 1934 5165 1935 5169
rect 1939 5165 1940 5169
rect 1934 5164 1940 5165
rect 1974 5168 1980 5169
rect 3798 5168 3804 5169
rect 1974 5164 1975 5168
rect 1979 5164 1980 5168
rect 1814 5163 1820 5164
rect 1974 5163 1980 5164
rect 2274 5167 2280 5168
rect 2274 5163 2275 5167
rect 2279 5163 2280 5167
rect 2274 5162 2280 5163
rect 2474 5167 2480 5168
rect 2474 5163 2475 5167
rect 2479 5163 2480 5167
rect 2474 5162 2480 5163
rect 2682 5167 2688 5168
rect 2682 5163 2683 5167
rect 2687 5163 2688 5167
rect 2682 5162 2688 5163
rect 2890 5167 2896 5168
rect 2890 5163 2891 5167
rect 2895 5163 2896 5167
rect 2890 5162 2896 5163
rect 3098 5167 3104 5168
rect 3098 5163 3099 5167
rect 3103 5163 3104 5167
rect 3098 5162 3104 5163
rect 3306 5167 3312 5168
rect 3306 5163 3307 5167
rect 3311 5163 3312 5167
rect 3798 5164 3799 5168
rect 3803 5164 3804 5168
rect 3798 5163 3804 5164
rect 4559 5163 4565 5164
rect 3306 5162 3312 5163
rect 4559 5159 4560 5163
rect 4564 5162 4565 5163
rect 4602 5163 4608 5164
rect 4602 5162 4603 5163
rect 4564 5160 4603 5162
rect 4564 5159 4565 5160
rect 4559 5158 4565 5159
rect 4602 5159 4603 5160
rect 4607 5159 4608 5163
rect 4602 5158 4608 5159
rect 4719 5163 4725 5164
rect 4719 5159 4720 5163
rect 4724 5162 4725 5163
rect 4743 5163 4749 5164
rect 4743 5162 4744 5163
rect 4724 5160 4744 5162
rect 4724 5159 4725 5160
rect 4719 5158 4725 5159
rect 4743 5159 4744 5160
rect 4748 5159 4749 5163
rect 4743 5158 4749 5159
rect 4879 5163 4885 5164
rect 4879 5159 4880 5163
rect 4884 5162 4885 5163
rect 4903 5163 4909 5164
rect 4903 5162 4904 5163
rect 4884 5160 4904 5162
rect 4884 5159 4885 5160
rect 4879 5158 4885 5159
rect 4903 5159 4904 5160
rect 4908 5159 4909 5163
rect 4903 5158 4909 5159
rect 5039 5163 5045 5164
rect 5039 5159 5040 5163
rect 5044 5162 5045 5163
rect 5047 5163 5053 5164
rect 5047 5162 5048 5163
rect 5044 5160 5048 5162
rect 5044 5159 5045 5160
rect 5039 5158 5045 5159
rect 5047 5159 5048 5160
rect 5052 5159 5053 5163
rect 5047 5158 5053 5159
rect 5191 5163 5197 5164
rect 5191 5159 5192 5163
rect 5196 5162 5197 5163
rect 5199 5163 5205 5164
rect 5199 5162 5200 5163
rect 5196 5160 5200 5162
rect 5196 5159 5197 5160
rect 5191 5158 5197 5159
rect 5199 5159 5200 5160
rect 5204 5159 5205 5163
rect 5199 5158 5205 5159
rect 5343 5163 5349 5164
rect 5343 5159 5344 5163
rect 5348 5162 5349 5163
rect 5367 5163 5373 5164
rect 5367 5162 5368 5163
rect 5348 5160 5368 5162
rect 5348 5159 5349 5160
rect 5343 5158 5349 5159
rect 5367 5159 5368 5160
rect 5372 5159 5373 5163
rect 5367 5158 5373 5159
rect 5503 5163 5509 5164
rect 5503 5159 5504 5163
rect 5508 5162 5509 5163
rect 5511 5163 5517 5164
rect 5511 5162 5512 5163
rect 5508 5160 5512 5162
rect 5508 5159 5509 5160
rect 5503 5158 5509 5159
rect 5511 5159 5512 5160
rect 5516 5159 5517 5163
rect 5511 5158 5517 5159
rect 5602 5163 5608 5164
rect 5602 5159 5603 5163
rect 5607 5162 5608 5163
rect 5639 5163 5645 5164
rect 5639 5162 5640 5163
rect 5607 5160 5640 5162
rect 5607 5159 5608 5160
rect 5602 5158 5608 5159
rect 5639 5159 5640 5160
rect 5644 5159 5645 5163
rect 5639 5158 5645 5159
rect 3838 5156 3844 5157
rect 5662 5156 5668 5157
rect 418 5153 424 5154
rect 110 5152 116 5153
rect 110 5148 111 5152
rect 115 5148 116 5152
rect 418 5149 419 5153
rect 423 5149 424 5153
rect 418 5148 424 5149
rect 594 5153 600 5154
rect 594 5149 595 5153
rect 599 5149 600 5153
rect 594 5148 600 5149
rect 778 5153 784 5154
rect 778 5149 779 5153
rect 783 5149 784 5153
rect 778 5148 784 5149
rect 970 5153 976 5154
rect 970 5149 971 5153
rect 975 5149 976 5153
rect 970 5148 976 5149
rect 1170 5153 1176 5154
rect 1170 5149 1171 5153
rect 1175 5149 1176 5153
rect 1170 5148 1176 5149
rect 1370 5153 1376 5154
rect 1370 5149 1371 5153
rect 1375 5149 1376 5153
rect 1370 5148 1376 5149
rect 1578 5153 1584 5154
rect 1578 5149 1579 5153
rect 1583 5149 1584 5153
rect 1578 5148 1584 5149
rect 1786 5153 1792 5154
rect 1786 5149 1787 5153
rect 1791 5149 1792 5153
rect 1786 5148 1792 5149
rect 1934 5152 1940 5153
rect 2302 5152 2308 5153
rect 1934 5148 1935 5152
rect 1939 5148 1940 5152
rect 110 5147 116 5148
rect 1934 5147 1940 5148
rect 1974 5151 1980 5152
rect 1974 5147 1975 5151
rect 1979 5147 1980 5151
rect 2302 5148 2303 5152
rect 2307 5148 2308 5152
rect 2302 5147 2308 5148
rect 2502 5152 2508 5153
rect 2502 5148 2503 5152
rect 2507 5148 2508 5152
rect 2502 5147 2508 5148
rect 2710 5152 2716 5153
rect 2710 5148 2711 5152
rect 2715 5148 2716 5152
rect 2710 5147 2716 5148
rect 2918 5152 2924 5153
rect 2918 5148 2919 5152
rect 2923 5148 2924 5152
rect 2918 5147 2924 5148
rect 3126 5152 3132 5153
rect 3126 5148 3127 5152
rect 3131 5148 3132 5152
rect 3126 5147 3132 5148
rect 3334 5152 3340 5153
rect 3838 5152 3839 5156
rect 3843 5152 3844 5156
rect 3334 5148 3335 5152
rect 3339 5148 3340 5152
rect 3334 5147 3340 5148
rect 3798 5151 3804 5152
rect 3838 5151 3844 5152
rect 4434 5155 4440 5156
rect 4434 5151 4435 5155
rect 4439 5151 4440 5155
rect 3798 5147 3799 5151
rect 3803 5147 3804 5151
rect 4434 5150 4440 5151
rect 4594 5155 4600 5156
rect 4594 5151 4595 5155
rect 4599 5151 4600 5155
rect 4594 5150 4600 5151
rect 4754 5155 4760 5156
rect 4754 5151 4755 5155
rect 4759 5151 4760 5155
rect 4754 5150 4760 5151
rect 4914 5155 4920 5156
rect 4914 5151 4915 5155
rect 4919 5151 4920 5155
rect 4914 5150 4920 5151
rect 5066 5155 5072 5156
rect 5066 5151 5067 5155
rect 5071 5151 5072 5155
rect 5066 5150 5072 5151
rect 5218 5155 5224 5156
rect 5218 5151 5219 5155
rect 5223 5151 5224 5155
rect 5218 5150 5224 5151
rect 5378 5155 5384 5156
rect 5378 5151 5379 5155
rect 5383 5151 5384 5155
rect 5378 5150 5384 5151
rect 5514 5155 5520 5156
rect 5514 5151 5515 5155
rect 5519 5151 5520 5155
rect 5662 5152 5663 5156
rect 5667 5152 5668 5156
rect 5662 5151 5668 5152
rect 5514 5150 5520 5151
rect 1974 5146 1980 5147
rect 3798 5146 3804 5147
rect 543 5143 549 5144
rect 543 5139 544 5143
rect 548 5142 549 5143
rect 610 5143 616 5144
rect 610 5142 611 5143
rect 548 5140 611 5142
rect 548 5139 549 5140
rect 543 5138 549 5139
rect 610 5139 611 5140
rect 615 5139 616 5143
rect 610 5138 616 5139
rect 714 5143 725 5144
rect 714 5139 715 5143
rect 719 5139 720 5143
rect 724 5139 725 5143
rect 714 5138 725 5139
rect 734 5143 740 5144
rect 734 5139 735 5143
rect 739 5142 740 5143
rect 903 5143 909 5144
rect 903 5142 904 5143
rect 739 5140 904 5142
rect 739 5139 740 5140
rect 734 5138 740 5139
rect 903 5139 904 5140
rect 908 5139 909 5143
rect 903 5138 909 5139
rect 943 5143 949 5144
rect 943 5139 944 5143
rect 948 5142 949 5143
rect 1095 5143 1101 5144
rect 1095 5142 1096 5143
rect 948 5140 1096 5142
rect 948 5139 949 5140
rect 943 5138 949 5139
rect 1095 5139 1096 5140
rect 1100 5139 1101 5143
rect 1095 5138 1101 5139
rect 1142 5143 1148 5144
rect 1142 5139 1143 5143
rect 1147 5142 1148 5143
rect 1295 5143 1301 5144
rect 1295 5142 1296 5143
rect 1147 5140 1296 5142
rect 1147 5139 1148 5140
rect 1142 5138 1148 5139
rect 1295 5139 1296 5140
rect 1300 5139 1301 5143
rect 1295 5138 1301 5139
rect 1490 5143 1501 5144
rect 1490 5139 1491 5143
rect 1495 5139 1496 5143
rect 1500 5139 1501 5143
rect 1490 5138 1501 5139
rect 1703 5143 1709 5144
rect 1703 5139 1704 5143
rect 1708 5142 1709 5143
rect 1802 5143 1808 5144
rect 1802 5142 1803 5143
rect 1708 5140 1803 5142
rect 1708 5139 1709 5140
rect 1703 5138 1709 5139
rect 1802 5139 1803 5140
rect 1807 5139 1808 5143
rect 1911 5143 1917 5144
rect 1911 5142 1912 5143
rect 1802 5138 1808 5139
rect 1812 5140 1912 5142
rect 1458 5135 1464 5136
rect 1458 5131 1459 5135
rect 1463 5134 1464 5135
rect 1812 5134 1814 5140
rect 1911 5139 1912 5140
rect 1916 5139 1917 5143
rect 4462 5140 4468 5141
rect 1911 5138 1917 5139
rect 3838 5139 3844 5140
rect 3838 5135 3839 5139
rect 3843 5135 3844 5139
rect 4462 5136 4463 5140
rect 4467 5136 4468 5140
rect 4462 5135 4468 5136
rect 4622 5140 4628 5141
rect 4622 5136 4623 5140
rect 4627 5136 4628 5140
rect 4622 5135 4628 5136
rect 4782 5140 4788 5141
rect 4782 5136 4783 5140
rect 4787 5136 4788 5140
rect 4782 5135 4788 5136
rect 4942 5140 4948 5141
rect 4942 5136 4943 5140
rect 4947 5136 4948 5140
rect 4942 5135 4948 5136
rect 5094 5140 5100 5141
rect 5094 5136 5095 5140
rect 5099 5136 5100 5140
rect 5094 5135 5100 5136
rect 5246 5140 5252 5141
rect 5246 5136 5247 5140
rect 5251 5136 5252 5140
rect 5246 5135 5252 5136
rect 5406 5140 5412 5141
rect 5406 5136 5407 5140
rect 5411 5136 5412 5140
rect 5406 5135 5412 5136
rect 5542 5140 5548 5141
rect 5542 5136 5543 5140
rect 5547 5136 5548 5140
rect 5542 5135 5548 5136
rect 5662 5139 5668 5140
rect 5662 5135 5663 5139
rect 5667 5135 5668 5139
rect 3838 5134 3844 5135
rect 5662 5134 5668 5135
rect 1463 5132 1814 5134
rect 1463 5131 1464 5132
rect 1458 5130 1464 5131
rect 610 5111 616 5112
rect 509 5108 530 5110
rect 528 5094 530 5108
rect 610 5107 611 5111
rect 615 5107 616 5111
rect 943 5111 949 5112
rect 943 5110 944 5111
rect 869 5108 944 5110
rect 610 5106 616 5107
rect 943 5107 944 5108
rect 948 5107 949 5111
rect 1142 5111 1148 5112
rect 1142 5110 1143 5111
rect 1061 5108 1143 5110
rect 943 5106 949 5107
rect 1142 5107 1143 5108
rect 1147 5107 1148 5111
rect 1142 5106 1148 5107
rect 1258 5111 1264 5112
rect 1258 5107 1259 5111
rect 1263 5107 1264 5111
rect 1258 5106 1264 5107
rect 1458 5111 1464 5112
rect 1458 5107 1459 5111
rect 1463 5107 1464 5111
rect 1458 5106 1464 5107
rect 1646 5111 1652 5112
rect 1646 5107 1647 5111
rect 1651 5107 1652 5111
rect 1646 5106 1652 5107
rect 1802 5111 1808 5112
rect 1802 5107 1803 5111
rect 1807 5107 1808 5111
rect 1802 5106 1808 5107
rect 734 5095 740 5096
rect 734 5094 735 5095
rect 528 5092 735 5094
rect 734 5091 735 5092
rect 739 5091 740 5095
rect 734 5090 740 5091
rect 274 5079 280 5080
rect 274 5075 275 5079
rect 279 5078 280 5079
rect 1318 5079 1324 5080
rect 1318 5078 1319 5079
rect 279 5076 1319 5078
rect 279 5075 280 5076
rect 274 5074 280 5075
rect 1318 5075 1319 5076
rect 1323 5075 1324 5079
rect 1318 5074 1324 5075
rect 1974 5077 1980 5078
rect 3798 5077 3804 5078
rect 1974 5073 1975 5077
rect 1979 5073 1980 5077
rect 1974 5072 1980 5073
rect 2118 5076 2124 5077
rect 2118 5072 2119 5076
rect 2123 5072 2124 5076
rect 2118 5071 2124 5072
rect 2326 5076 2332 5077
rect 2326 5072 2327 5076
rect 2331 5072 2332 5076
rect 2326 5071 2332 5072
rect 2534 5076 2540 5077
rect 2534 5072 2535 5076
rect 2539 5072 2540 5076
rect 2534 5071 2540 5072
rect 2750 5076 2756 5077
rect 2750 5072 2751 5076
rect 2755 5072 2756 5076
rect 2750 5071 2756 5072
rect 2974 5076 2980 5077
rect 2974 5072 2975 5076
rect 2979 5072 2980 5076
rect 2974 5071 2980 5072
rect 3206 5076 3212 5077
rect 3206 5072 3207 5076
rect 3211 5072 3212 5076
rect 3798 5073 3799 5077
rect 3803 5073 3804 5077
rect 3798 5072 3804 5073
rect 3838 5073 3844 5074
rect 5662 5073 5668 5074
rect 3206 5071 3212 5072
rect 3838 5069 3839 5073
rect 3843 5069 3844 5073
rect 3838 5068 3844 5069
rect 3886 5072 3892 5073
rect 3886 5068 3887 5072
rect 3891 5068 3892 5072
rect 3886 5067 3892 5068
rect 4086 5072 4092 5073
rect 4086 5068 4087 5072
rect 4091 5068 4092 5072
rect 4086 5067 4092 5068
rect 4326 5072 4332 5073
rect 4326 5068 4327 5072
rect 4331 5068 4332 5072
rect 4326 5067 4332 5068
rect 4566 5072 4572 5073
rect 4566 5068 4567 5072
rect 4571 5068 4572 5072
rect 4566 5067 4572 5068
rect 4814 5072 4820 5073
rect 4814 5068 4815 5072
rect 4819 5068 4820 5072
rect 4814 5067 4820 5068
rect 5062 5072 5068 5073
rect 5062 5068 5063 5072
rect 5067 5068 5068 5072
rect 5062 5067 5068 5068
rect 5310 5072 5316 5073
rect 5310 5068 5311 5072
rect 5315 5068 5316 5072
rect 5310 5067 5316 5068
rect 5542 5072 5548 5073
rect 5542 5068 5543 5072
rect 5547 5068 5548 5072
rect 5662 5069 5663 5073
rect 5667 5069 5668 5073
rect 5662 5068 5668 5069
rect 5542 5067 5548 5068
rect 2090 5061 2096 5062
rect 1974 5060 1980 5061
rect 1974 5056 1975 5060
rect 1979 5056 1980 5060
rect 2090 5057 2091 5061
rect 2095 5057 2096 5061
rect 2090 5056 2096 5057
rect 2298 5061 2304 5062
rect 2298 5057 2299 5061
rect 2303 5057 2304 5061
rect 2298 5056 2304 5057
rect 2506 5061 2512 5062
rect 2506 5057 2507 5061
rect 2511 5057 2512 5061
rect 2506 5056 2512 5057
rect 2722 5061 2728 5062
rect 2722 5057 2723 5061
rect 2727 5057 2728 5061
rect 2722 5056 2728 5057
rect 2946 5061 2952 5062
rect 2946 5057 2947 5061
rect 2951 5057 2952 5061
rect 2946 5056 2952 5057
rect 3178 5061 3184 5062
rect 3178 5057 3179 5061
rect 3183 5057 3184 5061
rect 3178 5056 3184 5057
rect 3798 5060 3804 5061
rect 3798 5056 3799 5060
rect 3803 5056 3804 5060
rect 3858 5057 3864 5058
rect 274 5055 280 5056
rect 274 5054 275 5055
rect 245 5052 275 5054
rect 274 5051 275 5052
rect 279 5051 280 5055
rect 274 5050 280 5051
rect 282 5055 288 5056
rect 282 5051 283 5055
rect 287 5054 288 5055
rect 754 5055 760 5056
rect 287 5052 397 5054
rect 287 5051 288 5052
rect 282 5050 288 5051
rect 714 5051 720 5052
rect 714 5047 715 5051
rect 719 5047 720 5051
rect 754 5051 755 5055
rect 759 5054 760 5055
rect 1118 5055 1124 5056
rect 759 5052 917 5054
rect 759 5051 760 5052
rect 754 5050 760 5051
rect 1118 5051 1119 5055
rect 1123 5054 1124 5055
rect 1490 5055 1496 5056
rect 1123 5052 1213 5054
rect 1123 5051 1124 5052
rect 1118 5050 1124 5051
rect 1490 5051 1491 5055
rect 1495 5054 1496 5055
rect 1626 5055 1632 5056
rect 1974 5055 1980 5056
rect 3798 5055 3804 5056
rect 3838 5056 3844 5057
rect 1495 5052 1517 5054
rect 1495 5051 1496 5052
rect 1490 5050 1496 5051
rect 1626 5051 1627 5055
rect 1631 5054 1632 5055
rect 1631 5052 1805 5054
rect 3838 5052 3839 5056
rect 3843 5052 3844 5056
rect 3858 5053 3859 5057
rect 3863 5053 3864 5057
rect 3858 5052 3864 5053
rect 4058 5057 4064 5058
rect 4058 5053 4059 5057
rect 4063 5053 4064 5057
rect 4058 5052 4064 5053
rect 4298 5057 4304 5058
rect 4298 5053 4299 5057
rect 4303 5053 4304 5057
rect 4298 5052 4304 5053
rect 4538 5057 4544 5058
rect 4538 5053 4539 5057
rect 4543 5053 4544 5057
rect 4538 5052 4544 5053
rect 4786 5057 4792 5058
rect 4786 5053 4787 5057
rect 4791 5053 4792 5057
rect 4786 5052 4792 5053
rect 5034 5057 5040 5058
rect 5034 5053 5035 5057
rect 5039 5053 5040 5057
rect 5034 5052 5040 5053
rect 5282 5057 5288 5058
rect 5282 5053 5283 5057
rect 5287 5053 5288 5057
rect 5282 5052 5288 5053
rect 5514 5057 5520 5058
rect 5514 5053 5515 5057
rect 5519 5053 5520 5057
rect 5514 5052 5520 5053
rect 5662 5056 5668 5057
rect 5662 5052 5663 5056
rect 5667 5052 5668 5056
rect 1631 5051 1632 5052
rect 1626 5050 1632 5051
rect 2215 5051 2221 5052
rect 714 5046 720 5047
rect 2215 5047 2216 5051
rect 2220 5050 2221 5051
rect 2354 5051 2360 5052
rect 2354 5050 2355 5051
rect 2220 5048 2355 5050
rect 2220 5047 2221 5048
rect 2215 5046 2221 5047
rect 2354 5047 2355 5048
rect 2359 5047 2360 5051
rect 2423 5051 2429 5052
rect 2423 5050 2424 5051
rect 2354 5046 2360 5047
rect 2364 5048 2424 5050
rect 2178 5043 2184 5044
rect 2178 5039 2179 5043
rect 2183 5042 2184 5043
rect 2364 5042 2366 5048
rect 2423 5047 2424 5048
rect 2428 5047 2429 5051
rect 2423 5046 2429 5047
rect 2471 5051 2477 5052
rect 2471 5047 2472 5051
rect 2476 5050 2477 5051
rect 2631 5051 2637 5052
rect 2631 5050 2632 5051
rect 2476 5048 2632 5050
rect 2476 5047 2477 5048
rect 2471 5046 2477 5047
rect 2631 5047 2632 5048
rect 2636 5047 2637 5051
rect 2631 5046 2637 5047
rect 2770 5051 2776 5052
rect 2770 5047 2771 5051
rect 2775 5050 2776 5051
rect 2847 5051 2853 5052
rect 2847 5050 2848 5051
rect 2775 5048 2848 5050
rect 2775 5047 2776 5048
rect 2770 5046 2776 5047
rect 2847 5047 2848 5048
rect 2852 5047 2853 5051
rect 2847 5046 2853 5047
rect 3071 5051 3077 5052
rect 3071 5047 3072 5051
rect 3076 5050 3077 5051
rect 3194 5051 3200 5052
rect 3194 5050 3195 5051
rect 3076 5048 3195 5050
rect 3076 5047 3077 5048
rect 3071 5046 3077 5047
rect 3194 5047 3195 5048
rect 3199 5047 3200 5051
rect 3194 5046 3200 5047
rect 3303 5051 3309 5052
rect 3303 5047 3304 5051
rect 3308 5050 3309 5051
rect 3319 5051 3325 5052
rect 3838 5051 3844 5052
rect 5662 5051 5668 5052
rect 3319 5050 3320 5051
rect 3308 5048 3320 5050
rect 3308 5047 3309 5048
rect 3303 5046 3309 5047
rect 3319 5047 3320 5048
rect 3324 5047 3325 5051
rect 3319 5046 3325 5047
rect 3983 5047 3989 5048
rect 3983 5043 3984 5047
rect 3988 5046 3989 5047
rect 4074 5047 4080 5048
rect 4074 5046 4075 5047
rect 3988 5044 4075 5046
rect 3988 5043 3989 5044
rect 3983 5042 3989 5043
rect 4074 5043 4075 5044
rect 4079 5043 4080 5047
rect 4074 5042 4080 5043
rect 4183 5047 4189 5048
rect 4183 5043 4184 5047
rect 4188 5046 4189 5047
rect 4218 5047 4224 5048
rect 4218 5046 4219 5047
rect 4188 5044 4219 5046
rect 4188 5043 4189 5044
rect 4183 5042 4189 5043
rect 4218 5043 4219 5044
rect 4223 5043 4224 5047
rect 4218 5042 4224 5043
rect 4423 5047 4432 5048
rect 4423 5043 4424 5047
rect 4431 5043 4432 5047
rect 4423 5042 4432 5043
rect 4458 5047 4464 5048
rect 4458 5043 4459 5047
rect 4463 5046 4464 5047
rect 4663 5047 4669 5048
rect 4663 5046 4664 5047
rect 4463 5044 4664 5046
rect 4463 5043 4464 5044
rect 4458 5042 4464 5043
rect 4663 5043 4664 5044
rect 4668 5043 4669 5047
rect 4663 5042 4669 5043
rect 4682 5047 4688 5048
rect 4682 5043 4683 5047
rect 4687 5046 4688 5047
rect 4911 5047 4917 5048
rect 4911 5046 4912 5047
rect 4687 5044 4912 5046
rect 4687 5043 4688 5044
rect 4682 5042 4688 5043
rect 4911 5043 4912 5044
rect 4916 5043 4917 5047
rect 4911 5042 4917 5043
rect 5159 5047 5165 5048
rect 5159 5043 5160 5047
rect 5164 5046 5165 5047
rect 5298 5047 5304 5048
rect 5298 5046 5299 5047
rect 5164 5044 5299 5046
rect 5164 5043 5165 5044
rect 5159 5042 5165 5043
rect 5298 5043 5299 5044
rect 5303 5043 5304 5047
rect 5298 5042 5304 5043
rect 5370 5047 5376 5048
rect 5370 5043 5371 5047
rect 5375 5046 5376 5047
rect 5407 5047 5413 5048
rect 5407 5046 5408 5047
rect 5375 5044 5408 5046
rect 5375 5043 5376 5044
rect 5370 5042 5376 5043
rect 5407 5043 5408 5044
rect 5412 5043 5413 5047
rect 5639 5047 5645 5048
rect 5639 5046 5640 5047
rect 5407 5042 5413 5043
rect 5416 5044 5640 5046
rect 2183 5040 2366 5042
rect 2183 5039 2184 5040
rect 2178 5038 2184 5039
rect 5122 5039 5128 5040
rect 5122 5035 5123 5039
rect 5127 5038 5128 5039
rect 5416 5038 5418 5044
rect 5639 5043 5640 5044
rect 5644 5043 5645 5047
rect 5639 5042 5645 5043
rect 5127 5036 5418 5038
rect 5127 5035 5128 5036
rect 5122 5034 5128 5035
rect 279 5019 288 5020
rect 279 5015 280 5019
rect 287 5015 288 5019
rect 279 5014 288 5015
rect 490 5019 496 5020
rect 490 5015 491 5019
rect 495 5018 496 5019
rect 503 5019 509 5020
rect 503 5018 504 5019
rect 495 5016 504 5018
rect 495 5015 496 5016
rect 490 5014 496 5015
rect 503 5015 504 5016
rect 508 5015 509 5019
rect 503 5014 509 5015
rect 751 5019 760 5020
rect 751 5015 752 5019
rect 759 5015 760 5019
rect 751 5014 760 5015
rect 1023 5019 1029 5020
rect 1023 5015 1024 5019
rect 1028 5018 1029 5019
rect 1118 5019 1124 5020
rect 1118 5018 1119 5019
rect 1028 5016 1119 5018
rect 1028 5015 1029 5016
rect 1023 5014 1029 5015
rect 1118 5015 1119 5016
rect 1123 5015 1124 5019
rect 1118 5014 1124 5015
rect 1318 5019 1325 5020
rect 1318 5015 1319 5019
rect 1324 5015 1325 5019
rect 1318 5014 1325 5015
rect 1623 5019 1632 5020
rect 1623 5015 1624 5019
rect 1631 5015 1632 5019
rect 1623 5014 1632 5015
rect 1911 5019 1917 5020
rect 1911 5015 1912 5019
rect 1916 5018 1917 5019
rect 1951 5019 1957 5020
rect 1951 5018 1952 5019
rect 1916 5016 1952 5018
rect 1916 5015 1917 5016
rect 1911 5014 1917 5015
rect 1951 5015 1952 5016
rect 1956 5015 1957 5019
rect 1951 5014 1957 5015
rect 2178 5019 2184 5020
rect 2178 5015 2179 5019
rect 2183 5015 2184 5019
rect 2471 5019 2477 5020
rect 2471 5018 2472 5019
rect 2389 5016 2472 5018
rect 2178 5014 2184 5015
rect 2471 5015 2472 5016
rect 2476 5015 2477 5019
rect 3078 5019 3084 5020
rect 3078 5018 3079 5019
rect 2597 5016 2662 5018
rect 2813 5016 2942 5018
rect 3037 5016 3079 5018
rect 2471 5014 2477 5015
rect 110 5012 116 5013
rect 1934 5012 1940 5013
rect 110 5008 111 5012
rect 115 5008 116 5012
rect 110 5007 116 5008
rect 154 5011 160 5012
rect 154 5007 155 5011
rect 159 5007 160 5011
rect 154 5006 160 5007
rect 378 5011 384 5012
rect 378 5007 379 5011
rect 383 5007 384 5011
rect 378 5006 384 5007
rect 626 5011 632 5012
rect 626 5007 627 5011
rect 631 5007 632 5011
rect 626 5006 632 5007
rect 898 5011 904 5012
rect 898 5007 899 5011
rect 903 5007 904 5011
rect 898 5006 904 5007
rect 1194 5011 1200 5012
rect 1194 5007 1195 5011
rect 1199 5007 1200 5011
rect 1194 5006 1200 5007
rect 1498 5011 1504 5012
rect 1498 5007 1499 5011
rect 1503 5007 1504 5011
rect 1498 5006 1504 5007
rect 1786 5011 1792 5012
rect 1786 5007 1787 5011
rect 1791 5007 1792 5011
rect 1934 5008 1935 5012
rect 1939 5008 1940 5012
rect 1934 5007 1940 5008
rect 1786 5006 1792 5007
rect 2660 5002 2662 5016
rect 2838 5003 2844 5004
rect 2838 5002 2839 5003
rect 2660 5000 2839 5002
rect 2838 4999 2839 5000
rect 2843 4999 2844 5003
rect 2940 5002 2942 5016
rect 3078 5015 3079 5016
rect 3083 5015 3084 5019
rect 3078 5014 3084 5015
rect 3194 5019 3200 5020
rect 3194 5015 3195 5019
rect 3199 5015 3200 5019
rect 3194 5014 3200 5015
rect 4066 5015 4072 5016
rect 4066 5014 4067 5015
rect 3949 5012 4067 5014
rect 4066 5011 4067 5012
rect 4071 5011 4072 5015
rect 4066 5010 4072 5011
rect 4074 5015 4080 5016
rect 4074 5011 4075 5015
rect 4079 5011 4080 5015
rect 4458 5015 4464 5016
rect 4458 5014 4459 5015
rect 4389 5012 4459 5014
rect 4074 5010 4080 5011
rect 4458 5011 4459 5012
rect 4463 5011 4464 5015
rect 4682 5015 4688 5016
rect 4682 5014 4683 5015
rect 4629 5012 4683 5014
rect 4458 5010 4464 5011
rect 4682 5011 4683 5012
rect 4687 5011 4688 5015
rect 4682 5010 4688 5011
rect 4874 5015 4880 5016
rect 4874 5011 4875 5015
rect 4879 5011 4880 5015
rect 4874 5010 4880 5011
rect 5122 5015 5128 5016
rect 5122 5011 5123 5015
rect 5127 5011 5128 5015
rect 5122 5010 5128 5011
rect 5298 5015 5304 5016
rect 5298 5011 5299 5015
rect 5303 5011 5304 5015
rect 5298 5010 5304 5011
rect 5602 5015 5608 5016
rect 5602 5011 5603 5015
rect 5607 5011 5608 5015
rect 5602 5010 5608 5011
rect 3246 5003 3252 5004
rect 3246 5002 3247 5003
rect 2940 5000 3247 5002
rect 2838 4998 2844 4999
rect 3246 4999 3247 5000
rect 3251 4999 3252 5003
rect 3246 4998 3252 4999
rect 182 4996 188 4997
rect 110 4995 116 4996
rect 110 4991 111 4995
rect 115 4991 116 4995
rect 182 4992 183 4996
rect 187 4992 188 4996
rect 182 4991 188 4992
rect 406 4996 412 4997
rect 406 4992 407 4996
rect 411 4992 412 4996
rect 406 4991 412 4992
rect 654 4996 660 4997
rect 654 4992 655 4996
rect 659 4992 660 4996
rect 654 4991 660 4992
rect 926 4996 932 4997
rect 926 4992 927 4996
rect 931 4992 932 4996
rect 926 4991 932 4992
rect 1222 4996 1228 4997
rect 1222 4992 1223 4996
rect 1227 4992 1228 4996
rect 1222 4991 1228 4992
rect 1526 4996 1532 4997
rect 1526 4992 1527 4996
rect 1531 4992 1532 4996
rect 1526 4991 1532 4992
rect 1814 4996 1820 4997
rect 1814 4992 1815 4996
rect 1819 4992 1820 4996
rect 1814 4991 1820 4992
rect 1934 4995 1940 4996
rect 1934 4991 1935 4995
rect 1939 4991 1940 4995
rect 110 4990 116 4991
rect 1934 4990 1940 4991
rect 3790 4967 3796 4968
rect 1951 4963 1957 4964
rect 1951 4959 1952 4963
rect 1956 4962 1957 4963
rect 2127 4963 2133 4964
rect 1956 4960 2013 4962
rect 1956 4959 1957 4960
rect 1951 4958 1957 4959
rect 2127 4959 2128 4963
rect 2132 4962 2133 4963
rect 2263 4963 2269 4964
rect 2132 4960 2149 4962
rect 2132 4959 2133 4960
rect 2127 4958 2133 4959
rect 2263 4959 2264 4963
rect 2268 4962 2269 4963
rect 2394 4963 2400 4964
rect 2268 4960 2285 4962
rect 2268 4959 2269 4960
rect 2263 4958 2269 4959
rect 2394 4959 2395 4963
rect 2399 4962 2400 4963
rect 2546 4963 2552 4964
rect 2399 4960 2437 4962
rect 2399 4959 2400 4960
rect 2394 4958 2400 4959
rect 2546 4959 2547 4963
rect 2551 4962 2552 4963
rect 2746 4963 2752 4964
rect 2551 4960 2637 4962
rect 2551 4959 2552 4960
rect 2546 4958 2552 4959
rect 2746 4959 2747 4963
rect 2751 4962 2752 4963
rect 2962 4963 2968 4964
rect 2751 4960 2877 4962
rect 2751 4959 2752 4960
rect 2746 4958 2752 4959
rect 2962 4959 2963 4963
rect 2967 4962 2968 4963
rect 3319 4963 3325 4964
rect 2967 4960 3141 4962
rect 2967 4959 2968 4960
rect 2962 4958 2968 4959
rect 3319 4959 3320 4963
rect 3324 4962 3325 4963
rect 3790 4963 3791 4967
rect 3795 4966 3796 4967
rect 3986 4967 3992 4968
rect 3795 4964 3877 4966
rect 3795 4963 3796 4964
rect 3790 4962 3796 4963
rect 3986 4963 3987 4967
rect 3991 4966 3992 4967
rect 4263 4967 4269 4968
rect 3991 4964 4013 4966
rect 3991 4963 3992 4964
rect 3986 4962 3992 4963
rect 4218 4963 4224 4964
rect 3324 4960 3413 4962
rect 3324 4959 3325 4960
rect 3319 4958 3325 4959
rect 3738 4959 3744 4960
rect 3738 4955 3739 4959
rect 3743 4955 3744 4959
rect 4218 4959 4219 4963
rect 4223 4959 4224 4963
rect 4263 4963 4264 4967
rect 4268 4966 4269 4967
rect 4399 4967 4405 4968
rect 4268 4964 4285 4966
rect 4268 4963 4269 4964
rect 4263 4962 4269 4963
rect 4399 4963 4400 4967
rect 4404 4966 4405 4967
rect 4535 4967 4541 4968
rect 4404 4964 4421 4966
rect 4404 4963 4405 4964
rect 4399 4962 4405 4963
rect 4535 4963 4536 4967
rect 4540 4966 4541 4967
rect 4671 4967 4677 4968
rect 4540 4964 4557 4966
rect 4540 4963 4541 4964
rect 4535 4962 4541 4963
rect 4671 4963 4672 4967
rect 4676 4966 4677 4967
rect 4802 4967 4808 4968
rect 4676 4964 4693 4966
rect 4676 4963 4677 4964
rect 4671 4962 4677 4963
rect 4802 4963 4803 4967
rect 4807 4966 4808 4967
rect 4943 4967 4949 4968
rect 4807 4964 4829 4966
rect 4807 4963 4808 4964
rect 4802 4962 4808 4963
rect 4943 4963 4944 4967
rect 4948 4966 4949 4967
rect 5079 4967 5085 4968
rect 4948 4964 4965 4966
rect 4948 4963 4949 4964
rect 4943 4962 4949 4963
rect 5079 4963 5080 4967
rect 5084 4966 5085 4967
rect 5210 4967 5216 4968
rect 5084 4964 5101 4966
rect 5084 4963 5085 4964
rect 5079 4962 5085 4963
rect 5210 4963 5211 4967
rect 5215 4966 5216 4967
rect 5370 4967 5376 4968
rect 5215 4964 5245 4966
rect 5215 4963 5216 4964
rect 5210 4962 5216 4963
rect 5370 4963 5371 4967
rect 5375 4966 5376 4967
rect 5511 4967 5517 4968
rect 5375 4964 5397 4966
rect 5375 4963 5376 4964
rect 5370 4962 5376 4963
rect 5511 4963 5512 4967
rect 5516 4966 5517 4967
rect 5516 4964 5533 4966
rect 5516 4963 5517 4964
rect 5511 4962 5517 4963
rect 4218 4958 4224 4959
rect 3738 4954 3744 4955
rect 3983 4931 3992 4932
rect 2119 4927 2125 4928
rect 2119 4923 2120 4927
rect 2124 4926 2125 4927
rect 2127 4927 2133 4928
rect 2127 4926 2128 4927
rect 2124 4924 2128 4926
rect 2124 4923 2125 4924
rect 2119 4922 2125 4923
rect 2127 4923 2128 4924
rect 2132 4923 2133 4927
rect 2127 4922 2133 4923
rect 2255 4927 2261 4928
rect 2255 4923 2256 4927
rect 2260 4926 2261 4927
rect 2263 4927 2269 4928
rect 2263 4926 2264 4927
rect 2260 4924 2264 4926
rect 2260 4923 2261 4924
rect 2255 4922 2261 4923
rect 2263 4923 2264 4924
rect 2268 4923 2269 4927
rect 2263 4922 2269 4923
rect 2391 4927 2400 4928
rect 2391 4923 2392 4927
rect 2399 4923 2400 4927
rect 2391 4922 2400 4923
rect 2543 4927 2552 4928
rect 2543 4923 2544 4927
rect 2551 4923 2552 4927
rect 2543 4922 2552 4923
rect 2743 4927 2752 4928
rect 2743 4923 2744 4927
rect 2751 4923 2752 4927
rect 2743 4922 2752 4923
rect 2838 4927 2844 4928
rect 2838 4923 2839 4927
rect 2843 4926 2844 4927
rect 2983 4927 2989 4928
rect 2983 4926 2984 4927
rect 2843 4924 2984 4926
rect 2843 4923 2844 4924
rect 2838 4922 2844 4923
rect 2983 4923 2984 4924
rect 2988 4923 2989 4927
rect 2983 4922 2989 4923
rect 3246 4927 3253 4928
rect 3246 4923 3247 4927
rect 3252 4923 3253 4927
rect 3246 4922 3253 4923
rect 3458 4927 3464 4928
rect 3458 4923 3459 4927
rect 3463 4926 3464 4927
rect 3519 4927 3525 4928
rect 3519 4926 3520 4927
rect 3463 4924 3520 4926
rect 3463 4923 3464 4924
rect 3458 4922 3464 4923
rect 3519 4923 3520 4924
rect 3524 4923 3525 4927
rect 3519 4922 3525 4923
rect 3775 4927 3781 4928
rect 3775 4923 3776 4927
rect 3780 4926 3781 4927
rect 3790 4927 3796 4928
rect 3790 4926 3791 4927
rect 3780 4924 3791 4926
rect 3780 4923 3781 4924
rect 3775 4922 3781 4923
rect 3790 4923 3791 4924
rect 3795 4923 3796 4927
rect 3983 4927 3984 4931
rect 3991 4927 3992 4931
rect 3983 4926 3992 4927
rect 4066 4931 4072 4932
rect 4066 4927 4067 4931
rect 4071 4930 4072 4931
rect 4119 4931 4125 4932
rect 4119 4930 4120 4931
rect 4071 4928 4120 4930
rect 4071 4927 4072 4928
rect 4066 4926 4072 4927
rect 4119 4927 4120 4928
rect 4124 4927 4125 4931
rect 4119 4926 4125 4927
rect 4255 4931 4261 4932
rect 4255 4927 4256 4931
rect 4260 4930 4261 4931
rect 4263 4931 4269 4932
rect 4263 4930 4264 4931
rect 4260 4928 4264 4930
rect 4260 4927 4261 4928
rect 4255 4926 4261 4927
rect 4263 4927 4264 4928
rect 4268 4927 4269 4931
rect 4263 4926 4269 4927
rect 4391 4931 4397 4932
rect 4391 4927 4392 4931
rect 4396 4930 4397 4931
rect 4399 4931 4405 4932
rect 4399 4930 4400 4931
rect 4396 4928 4400 4930
rect 4396 4927 4397 4928
rect 4391 4926 4397 4927
rect 4399 4927 4400 4928
rect 4404 4927 4405 4931
rect 4399 4926 4405 4927
rect 4527 4931 4533 4932
rect 4527 4927 4528 4931
rect 4532 4930 4533 4931
rect 4535 4931 4541 4932
rect 4535 4930 4536 4931
rect 4532 4928 4536 4930
rect 4532 4927 4533 4928
rect 4527 4926 4533 4927
rect 4535 4927 4536 4928
rect 4540 4927 4541 4931
rect 4535 4926 4541 4927
rect 4663 4931 4669 4932
rect 4663 4927 4664 4931
rect 4668 4930 4669 4931
rect 4671 4931 4677 4932
rect 4671 4930 4672 4931
rect 4668 4928 4672 4930
rect 4668 4927 4669 4928
rect 4663 4926 4669 4927
rect 4671 4927 4672 4928
rect 4676 4927 4677 4931
rect 4671 4926 4677 4927
rect 4799 4931 4808 4932
rect 4799 4927 4800 4931
rect 4807 4927 4808 4931
rect 4799 4926 4808 4927
rect 4935 4931 4941 4932
rect 4935 4927 4936 4931
rect 4940 4930 4941 4931
rect 4943 4931 4949 4932
rect 4943 4930 4944 4931
rect 4940 4928 4944 4930
rect 4940 4927 4941 4928
rect 4935 4926 4941 4927
rect 4943 4927 4944 4928
rect 4948 4927 4949 4931
rect 4943 4926 4949 4927
rect 5071 4931 5077 4932
rect 5071 4927 5072 4931
rect 5076 4930 5077 4931
rect 5079 4931 5085 4932
rect 5079 4930 5080 4931
rect 5076 4928 5080 4930
rect 5076 4927 5077 4928
rect 5071 4926 5077 4927
rect 5079 4927 5080 4928
rect 5084 4927 5085 4931
rect 5079 4926 5085 4927
rect 5207 4931 5216 4932
rect 5207 4927 5208 4931
rect 5215 4927 5216 4931
rect 5207 4926 5216 4927
rect 5238 4931 5244 4932
rect 5238 4927 5239 4931
rect 5243 4930 5244 4931
rect 5351 4931 5357 4932
rect 5351 4930 5352 4931
rect 5243 4928 5352 4930
rect 5243 4927 5244 4928
rect 5238 4926 5244 4927
rect 5351 4927 5352 4928
rect 5356 4927 5357 4931
rect 5351 4926 5357 4927
rect 5503 4931 5509 4932
rect 5503 4927 5504 4931
rect 5508 4930 5509 4931
rect 5511 4931 5517 4932
rect 5511 4930 5512 4931
rect 5508 4928 5512 4930
rect 5508 4927 5509 4928
rect 5503 4926 5509 4927
rect 5511 4927 5512 4928
rect 5516 4927 5517 4931
rect 5511 4926 5517 4927
rect 5602 4931 5608 4932
rect 5602 4927 5603 4931
rect 5607 4930 5608 4931
rect 5639 4931 5645 4932
rect 5639 4930 5640 4931
rect 5607 4928 5640 4930
rect 5607 4927 5608 4928
rect 5602 4926 5608 4927
rect 5639 4927 5640 4928
rect 5644 4927 5645 4931
rect 5639 4926 5645 4927
rect 3790 4922 3796 4923
rect 3838 4924 3844 4925
rect 5662 4924 5668 4925
rect 1974 4920 1980 4921
rect 3798 4920 3804 4921
rect 1974 4916 1975 4920
rect 1979 4916 1980 4920
rect 1974 4915 1980 4916
rect 1994 4919 2000 4920
rect 1994 4915 1995 4919
rect 1999 4915 2000 4919
rect 1994 4914 2000 4915
rect 2130 4919 2136 4920
rect 2130 4915 2131 4919
rect 2135 4915 2136 4919
rect 2130 4914 2136 4915
rect 2266 4919 2272 4920
rect 2266 4915 2267 4919
rect 2271 4915 2272 4919
rect 2266 4914 2272 4915
rect 2418 4919 2424 4920
rect 2418 4915 2419 4919
rect 2423 4915 2424 4919
rect 2418 4914 2424 4915
rect 2618 4919 2624 4920
rect 2618 4915 2619 4919
rect 2623 4915 2624 4919
rect 2618 4914 2624 4915
rect 2858 4919 2864 4920
rect 2858 4915 2859 4919
rect 2863 4915 2864 4919
rect 2858 4914 2864 4915
rect 3122 4919 3128 4920
rect 3122 4915 3123 4919
rect 3127 4915 3128 4919
rect 3122 4914 3128 4915
rect 3394 4919 3400 4920
rect 3394 4915 3395 4919
rect 3399 4915 3400 4919
rect 3394 4914 3400 4915
rect 3650 4919 3656 4920
rect 3650 4915 3651 4919
rect 3655 4915 3656 4919
rect 3798 4916 3799 4920
rect 3803 4916 3804 4920
rect 3838 4920 3839 4924
rect 3843 4920 3844 4924
rect 3838 4919 3844 4920
rect 3858 4923 3864 4924
rect 3858 4919 3859 4923
rect 3863 4919 3864 4923
rect 3858 4918 3864 4919
rect 3994 4923 4000 4924
rect 3994 4919 3995 4923
rect 3999 4919 4000 4923
rect 3994 4918 4000 4919
rect 4130 4923 4136 4924
rect 4130 4919 4131 4923
rect 4135 4919 4136 4923
rect 4130 4918 4136 4919
rect 4266 4923 4272 4924
rect 4266 4919 4267 4923
rect 4271 4919 4272 4923
rect 4266 4918 4272 4919
rect 4402 4923 4408 4924
rect 4402 4919 4403 4923
rect 4407 4919 4408 4923
rect 4402 4918 4408 4919
rect 4538 4923 4544 4924
rect 4538 4919 4539 4923
rect 4543 4919 4544 4923
rect 4538 4918 4544 4919
rect 4674 4923 4680 4924
rect 4674 4919 4675 4923
rect 4679 4919 4680 4923
rect 4674 4918 4680 4919
rect 4810 4923 4816 4924
rect 4810 4919 4811 4923
rect 4815 4919 4816 4923
rect 4810 4918 4816 4919
rect 4946 4923 4952 4924
rect 4946 4919 4947 4923
rect 4951 4919 4952 4923
rect 4946 4918 4952 4919
rect 5082 4923 5088 4924
rect 5082 4919 5083 4923
rect 5087 4919 5088 4923
rect 5082 4918 5088 4919
rect 5226 4923 5232 4924
rect 5226 4919 5227 4923
rect 5231 4919 5232 4923
rect 5226 4918 5232 4919
rect 5378 4923 5384 4924
rect 5378 4919 5379 4923
rect 5383 4919 5384 4923
rect 5378 4918 5384 4919
rect 5514 4923 5520 4924
rect 5514 4919 5515 4923
rect 5519 4919 5520 4923
rect 5662 4920 5663 4924
rect 5667 4920 5668 4924
rect 5662 4919 5668 4920
rect 5514 4918 5520 4919
rect 3798 4915 3804 4916
rect 3650 4914 3656 4915
rect 110 4909 116 4910
rect 1934 4909 1940 4910
rect 110 4905 111 4909
rect 115 4905 116 4909
rect 110 4904 116 4905
rect 158 4908 164 4909
rect 158 4904 159 4908
rect 163 4904 164 4908
rect 158 4903 164 4904
rect 294 4908 300 4909
rect 294 4904 295 4908
rect 299 4904 300 4908
rect 294 4903 300 4904
rect 430 4908 436 4909
rect 430 4904 431 4908
rect 435 4904 436 4908
rect 430 4903 436 4904
rect 566 4908 572 4909
rect 566 4904 567 4908
rect 571 4904 572 4908
rect 566 4903 572 4904
rect 702 4908 708 4909
rect 702 4904 703 4908
rect 707 4904 708 4908
rect 1934 4905 1935 4909
rect 1939 4905 1940 4909
rect 3886 4908 3892 4909
rect 3838 4907 3844 4908
rect 1934 4904 1940 4905
rect 2022 4904 2028 4905
rect 702 4903 708 4904
rect 1974 4903 1980 4904
rect 1974 4899 1975 4903
rect 1979 4899 1980 4903
rect 2022 4900 2023 4904
rect 2027 4900 2028 4904
rect 2022 4899 2028 4900
rect 2158 4904 2164 4905
rect 2158 4900 2159 4904
rect 2163 4900 2164 4904
rect 2158 4899 2164 4900
rect 2294 4904 2300 4905
rect 2294 4900 2295 4904
rect 2299 4900 2300 4904
rect 2294 4899 2300 4900
rect 2446 4904 2452 4905
rect 2446 4900 2447 4904
rect 2451 4900 2452 4904
rect 2446 4899 2452 4900
rect 2646 4904 2652 4905
rect 2646 4900 2647 4904
rect 2651 4900 2652 4904
rect 2646 4899 2652 4900
rect 2886 4904 2892 4905
rect 2886 4900 2887 4904
rect 2891 4900 2892 4904
rect 2886 4899 2892 4900
rect 3150 4904 3156 4905
rect 3150 4900 3151 4904
rect 3155 4900 3156 4904
rect 3150 4899 3156 4900
rect 3422 4904 3428 4905
rect 3422 4900 3423 4904
rect 3427 4900 3428 4904
rect 3422 4899 3428 4900
rect 3678 4904 3684 4905
rect 3678 4900 3679 4904
rect 3683 4900 3684 4904
rect 3678 4899 3684 4900
rect 3798 4903 3804 4904
rect 3798 4899 3799 4903
rect 3803 4899 3804 4903
rect 3838 4903 3839 4907
rect 3843 4903 3844 4907
rect 3886 4904 3887 4908
rect 3891 4904 3892 4908
rect 3886 4903 3892 4904
rect 4022 4908 4028 4909
rect 4022 4904 4023 4908
rect 4027 4904 4028 4908
rect 4022 4903 4028 4904
rect 4158 4908 4164 4909
rect 4158 4904 4159 4908
rect 4163 4904 4164 4908
rect 4158 4903 4164 4904
rect 4294 4908 4300 4909
rect 4294 4904 4295 4908
rect 4299 4904 4300 4908
rect 4294 4903 4300 4904
rect 4430 4908 4436 4909
rect 4430 4904 4431 4908
rect 4435 4904 4436 4908
rect 4430 4903 4436 4904
rect 4566 4908 4572 4909
rect 4566 4904 4567 4908
rect 4571 4904 4572 4908
rect 4566 4903 4572 4904
rect 4702 4908 4708 4909
rect 4702 4904 4703 4908
rect 4707 4904 4708 4908
rect 4702 4903 4708 4904
rect 4838 4908 4844 4909
rect 4838 4904 4839 4908
rect 4843 4904 4844 4908
rect 4838 4903 4844 4904
rect 4974 4908 4980 4909
rect 4974 4904 4975 4908
rect 4979 4904 4980 4908
rect 4974 4903 4980 4904
rect 5110 4908 5116 4909
rect 5110 4904 5111 4908
rect 5115 4904 5116 4908
rect 5110 4903 5116 4904
rect 5254 4908 5260 4909
rect 5254 4904 5255 4908
rect 5259 4904 5260 4908
rect 5254 4903 5260 4904
rect 5406 4908 5412 4909
rect 5406 4904 5407 4908
rect 5411 4904 5412 4908
rect 5406 4903 5412 4904
rect 5542 4908 5548 4909
rect 5542 4904 5543 4908
rect 5547 4904 5548 4908
rect 5542 4903 5548 4904
rect 5662 4907 5668 4908
rect 5662 4903 5663 4907
rect 5667 4903 5668 4907
rect 3838 4902 3844 4903
rect 5662 4902 5668 4903
rect 1974 4898 1980 4899
rect 3798 4898 3804 4899
rect 130 4893 136 4894
rect 110 4892 116 4893
rect 110 4888 111 4892
rect 115 4888 116 4892
rect 130 4889 131 4893
rect 135 4889 136 4893
rect 130 4888 136 4889
rect 266 4893 272 4894
rect 266 4889 267 4893
rect 271 4889 272 4893
rect 266 4888 272 4889
rect 402 4893 408 4894
rect 402 4889 403 4893
rect 407 4889 408 4893
rect 402 4888 408 4889
rect 538 4893 544 4894
rect 538 4889 539 4893
rect 543 4889 544 4893
rect 538 4888 544 4889
rect 674 4893 680 4894
rect 674 4889 675 4893
rect 679 4889 680 4893
rect 674 4888 680 4889
rect 1934 4892 1940 4893
rect 1934 4888 1935 4892
rect 1939 4888 1940 4892
rect 110 4887 116 4888
rect 1934 4887 1940 4888
rect 234 4883 240 4884
rect 234 4879 235 4883
rect 239 4882 240 4883
rect 255 4883 261 4884
rect 255 4882 256 4883
rect 239 4880 256 4882
rect 239 4879 240 4880
rect 234 4878 240 4879
rect 255 4879 256 4880
rect 260 4879 261 4883
rect 255 4878 261 4879
rect 263 4883 269 4884
rect 263 4879 264 4883
rect 268 4882 269 4883
rect 391 4883 397 4884
rect 391 4882 392 4883
rect 268 4880 392 4882
rect 268 4879 269 4880
rect 263 4878 269 4879
rect 391 4879 392 4880
rect 396 4879 397 4883
rect 391 4878 397 4879
rect 527 4883 533 4884
rect 527 4879 528 4883
rect 532 4882 533 4883
rect 554 4883 560 4884
rect 554 4882 555 4883
rect 532 4880 555 4882
rect 532 4879 533 4880
rect 527 4878 533 4879
rect 554 4879 555 4880
rect 559 4879 560 4883
rect 554 4878 560 4879
rect 663 4883 669 4884
rect 663 4879 664 4883
rect 668 4882 669 4883
rect 690 4883 696 4884
rect 690 4882 691 4883
rect 668 4880 691 4882
rect 668 4879 669 4880
rect 663 4878 669 4879
rect 690 4879 691 4880
rect 695 4879 696 4883
rect 799 4883 805 4884
rect 799 4882 800 4883
rect 690 4878 696 4879
rect 708 4880 800 4882
rect 354 4875 360 4876
rect 354 4871 355 4875
rect 359 4874 360 4875
rect 708 4874 710 4880
rect 799 4879 800 4880
rect 804 4879 805 4883
rect 799 4878 805 4879
rect 359 4872 710 4874
rect 359 4871 360 4872
rect 354 4870 360 4871
rect 263 4851 269 4852
rect 263 4850 264 4851
rect 221 4848 264 4850
rect 263 4847 264 4848
rect 268 4847 269 4851
rect 263 4846 269 4847
rect 354 4851 360 4852
rect 354 4847 355 4851
rect 359 4847 360 4851
rect 354 4846 360 4847
rect 490 4851 496 4852
rect 490 4847 491 4851
rect 495 4847 496 4851
rect 490 4846 496 4847
rect 554 4851 560 4852
rect 554 4847 555 4851
rect 559 4847 560 4851
rect 554 4846 560 4847
rect 690 4851 696 4852
rect 690 4847 691 4851
rect 695 4847 696 4851
rect 690 4846 696 4847
rect 1974 4837 1980 4838
rect 3798 4837 3804 4838
rect 1974 4833 1975 4837
rect 1979 4833 1980 4837
rect 1974 4832 1980 4833
rect 2326 4836 2332 4837
rect 2326 4832 2327 4836
rect 2331 4832 2332 4836
rect 2326 4831 2332 4832
rect 2558 4836 2564 4837
rect 2558 4832 2559 4836
rect 2563 4832 2564 4836
rect 2558 4831 2564 4832
rect 2822 4836 2828 4837
rect 2822 4832 2823 4836
rect 2827 4832 2828 4836
rect 2822 4831 2828 4832
rect 3102 4836 3108 4837
rect 3102 4832 3103 4836
rect 3107 4832 3108 4836
rect 3102 4831 3108 4832
rect 3398 4836 3404 4837
rect 3398 4832 3399 4836
rect 3403 4832 3404 4836
rect 3398 4831 3404 4832
rect 3678 4836 3684 4837
rect 3678 4832 3679 4836
rect 3683 4832 3684 4836
rect 3798 4833 3799 4837
rect 3803 4833 3804 4837
rect 3798 4832 3804 4833
rect 3678 4831 3684 4832
rect 2298 4821 2304 4822
rect 1974 4820 1980 4821
rect 1974 4816 1975 4820
rect 1979 4816 1980 4820
rect 2298 4817 2299 4821
rect 2303 4817 2304 4821
rect 2298 4816 2304 4817
rect 2530 4821 2536 4822
rect 2530 4817 2531 4821
rect 2535 4817 2536 4821
rect 2530 4816 2536 4817
rect 2794 4821 2800 4822
rect 2794 4817 2795 4821
rect 2799 4817 2800 4821
rect 2794 4816 2800 4817
rect 3074 4821 3080 4822
rect 3074 4817 3075 4821
rect 3079 4817 3080 4821
rect 3074 4816 3080 4817
rect 3370 4821 3376 4822
rect 3370 4817 3371 4821
rect 3375 4817 3376 4821
rect 3370 4816 3376 4817
rect 3650 4821 3656 4822
rect 3650 4817 3651 4821
rect 3655 4817 3656 4821
rect 3650 4816 3656 4817
rect 3798 4820 3804 4821
rect 3798 4816 3799 4820
rect 3803 4816 3804 4820
rect 1974 4815 1980 4816
rect 3798 4815 3804 4816
rect 2423 4811 2429 4812
rect 2423 4807 2424 4811
rect 2428 4810 2429 4811
rect 2546 4811 2552 4812
rect 2546 4810 2547 4811
rect 2428 4808 2547 4810
rect 2428 4807 2429 4808
rect 2423 4806 2429 4807
rect 2546 4807 2547 4808
rect 2551 4807 2552 4811
rect 2546 4806 2552 4807
rect 2655 4811 2661 4812
rect 2655 4807 2656 4811
rect 2660 4810 2661 4811
rect 2810 4811 2816 4812
rect 2810 4810 2811 4811
rect 2660 4808 2811 4810
rect 2660 4807 2661 4808
rect 2655 4806 2661 4807
rect 2810 4807 2811 4808
rect 2815 4807 2816 4811
rect 2810 4806 2816 4807
rect 2919 4811 2925 4812
rect 2919 4807 2920 4811
rect 2924 4810 2925 4811
rect 2962 4811 2968 4812
rect 2962 4810 2963 4811
rect 2924 4808 2963 4810
rect 2924 4807 2925 4808
rect 2919 4806 2925 4807
rect 2962 4807 2963 4808
rect 2967 4807 2968 4811
rect 3199 4811 3205 4812
rect 3199 4810 3200 4811
rect 2962 4806 2968 4807
rect 3139 4808 3200 4810
rect 2666 4803 2672 4804
rect 2666 4799 2667 4803
rect 2671 4802 2672 4803
rect 3139 4802 3141 4808
rect 3199 4807 3200 4808
rect 3204 4807 3205 4811
rect 3199 4806 3205 4807
rect 3311 4811 3317 4812
rect 3311 4807 3312 4811
rect 3316 4810 3317 4811
rect 3495 4811 3501 4812
rect 3495 4810 3496 4811
rect 3316 4808 3496 4810
rect 3316 4807 3317 4808
rect 3311 4806 3317 4807
rect 3495 4807 3496 4808
rect 3500 4807 3501 4811
rect 3495 4806 3501 4807
rect 3738 4811 3744 4812
rect 3738 4807 3739 4811
rect 3743 4810 3744 4811
rect 3775 4811 3781 4812
rect 3775 4810 3776 4811
rect 3743 4808 3776 4810
rect 3743 4807 3744 4808
rect 3738 4806 3744 4807
rect 3775 4807 3776 4808
rect 3780 4807 3781 4811
rect 3775 4806 3781 4807
rect 2671 4800 3141 4802
rect 2671 4799 2672 4800
rect 2666 4798 2672 4799
rect 234 4791 240 4792
rect 234 4790 235 4791
rect 221 4788 235 4790
rect 234 4787 235 4788
rect 239 4787 240 4791
rect 234 4786 240 4787
rect 258 4791 264 4792
rect 258 4787 259 4791
rect 263 4790 264 4791
rect 394 4791 400 4792
rect 263 4788 285 4790
rect 263 4787 264 4788
rect 258 4786 264 4787
rect 394 4787 395 4791
rect 399 4790 400 4791
rect 530 4791 536 4792
rect 399 4788 421 4790
rect 399 4787 400 4788
rect 394 4786 400 4787
rect 530 4787 531 4791
rect 535 4790 536 4791
rect 666 4791 672 4792
rect 535 4788 557 4790
rect 535 4787 536 4788
rect 530 4786 536 4787
rect 666 4787 667 4791
rect 671 4790 672 4791
rect 671 4788 693 4790
rect 671 4787 672 4788
rect 666 4786 672 4787
rect 2386 4779 2392 4780
rect 2386 4775 2387 4779
rect 2391 4775 2392 4779
rect 2386 4774 2392 4775
rect 2546 4779 2552 4780
rect 2546 4775 2547 4779
rect 2551 4775 2552 4779
rect 2546 4774 2552 4775
rect 2810 4779 2816 4780
rect 2810 4775 2811 4779
rect 2815 4775 2816 4779
rect 3311 4779 3317 4780
rect 3311 4778 3312 4779
rect 3165 4776 3312 4778
rect 2810 4774 2816 4775
rect 3311 4775 3312 4776
rect 3316 4775 3317 4779
rect 3311 4774 3317 4775
rect 3458 4779 3464 4780
rect 3458 4775 3459 4779
rect 3463 4775 3464 4779
rect 3458 4774 3464 4775
rect 3738 4779 3744 4780
rect 3738 4775 3739 4779
rect 3743 4775 3744 4779
rect 3738 4774 3744 4775
rect 3838 4773 3844 4774
rect 5662 4773 5668 4774
rect 3838 4769 3839 4773
rect 3843 4769 3844 4773
rect 3838 4768 3844 4769
rect 3886 4772 3892 4773
rect 3886 4768 3887 4772
rect 3891 4768 3892 4772
rect 3886 4767 3892 4768
rect 4070 4772 4076 4773
rect 4070 4768 4071 4772
rect 4075 4768 4076 4772
rect 4070 4767 4076 4768
rect 4294 4772 4300 4773
rect 4294 4768 4295 4772
rect 4299 4768 4300 4772
rect 4294 4767 4300 4768
rect 4534 4772 4540 4773
rect 4534 4768 4535 4772
rect 4539 4768 4540 4772
rect 4534 4767 4540 4768
rect 4782 4772 4788 4773
rect 4782 4768 4783 4772
rect 4787 4768 4788 4772
rect 4782 4767 4788 4768
rect 5038 4772 5044 4773
rect 5038 4768 5039 4772
rect 5043 4768 5044 4772
rect 5038 4767 5044 4768
rect 5302 4772 5308 4773
rect 5302 4768 5303 4772
rect 5307 4768 5308 4772
rect 5302 4767 5308 4768
rect 5542 4772 5548 4773
rect 5542 4768 5543 4772
rect 5547 4768 5548 4772
rect 5662 4769 5663 4773
rect 5667 4769 5668 4773
rect 5662 4768 5668 4769
rect 5542 4767 5548 4768
rect 218 4763 224 4764
rect 218 4759 219 4763
rect 223 4762 224 4763
rect 223 4760 803 4762
rect 223 4759 224 4760
rect 218 4758 224 4759
rect 801 4756 803 4760
rect 3858 4757 3864 4758
rect 3838 4756 3844 4757
rect 255 4755 264 4756
rect 255 4751 256 4755
rect 263 4751 264 4755
rect 255 4750 264 4751
rect 391 4755 400 4756
rect 391 4751 392 4755
rect 399 4751 400 4755
rect 391 4750 400 4751
rect 527 4755 536 4756
rect 527 4751 528 4755
rect 535 4751 536 4755
rect 527 4750 536 4751
rect 663 4755 672 4756
rect 663 4751 664 4755
rect 671 4751 672 4755
rect 663 4750 672 4751
rect 799 4755 805 4756
rect 799 4751 800 4755
rect 804 4751 805 4755
rect 3838 4752 3839 4756
rect 3843 4752 3844 4756
rect 3858 4753 3859 4757
rect 3863 4753 3864 4757
rect 3858 4752 3864 4753
rect 4042 4757 4048 4758
rect 4042 4753 4043 4757
rect 4047 4753 4048 4757
rect 4042 4752 4048 4753
rect 4266 4757 4272 4758
rect 4266 4753 4267 4757
rect 4271 4753 4272 4757
rect 4266 4752 4272 4753
rect 4506 4757 4512 4758
rect 4506 4753 4507 4757
rect 4511 4753 4512 4757
rect 4506 4752 4512 4753
rect 4754 4757 4760 4758
rect 4754 4753 4755 4757
rect 4759 4753 4760 4757
rect 4754 4752 4760 4753
rect 5010 4757 5016 4758
rect 5010 4753 5011 4757
rect 5015 4753 5016 4757
rect 5010 4752 5016 4753
rect 5274 4757 5280 4758
rect 5274 4753 5275 4757
rect 5279 4753 5280 4757
rect 5274 4752 5280 4753
rect 5514 4757 5520 4758
rect 5514 4753 5515 4757
rect 5519 4753 5520 4757
rect 5514 4752 5520 4753
rect 5662 4756 5668 4757
rect 5662 4752 5663 4756
rect 5667 4752 5668 4756
rect 3838 4751 3844 4752
rect 5662 4751 5668 4752
rect 799 4750 805 4751
rect 110 4748 116 4749
rect 1934 4748 1940 4749
rect 110 4744 111 4748
rect 115 4744 116 4748
rect 110 4743 116 4744
rect 130 4747 136 4748
rect 130 4743 131 4747
rect 135 4743 136 4747
rect 130 4742 136 4743
rect 266 4747 272 4748
rect 266 4743 267 4747
rect 271 4743 272 4747
rect 266 4742 272 4743
rect 402 4747 408 4748
rect 402 4743 403 4747
rect 407 4743 408 4747
rect 402 4742 408 4743
rect 538 4747 544 4748
rect 538 4743 539 4747
rect 543 4743 544 4747
rect 538 4742 544 4743
rect 674 4747 680 4748
rect 674 4743 675 4747
rect 679 4743 680 4747
rect 1934 4744 1935 4748
rect 1939 4744 1940 4748
rect 1934 4743 1940 4744
rect 3738 4747 3744 4748
rect 3738 4743 3739 4747
rect 3743 4746 3744 4747
rect 3983 4747 3989 4748
rect 3983 4746 3984 4747
rect 3743 4744 3984 4746
rect 3743 4743 3744 4744
rect 674 4742 680 4743
rect 3738 4742 3744 4743
rect 3983 4743 3984 4744
rect 3988 4743 3989 4747
rect 3983 4742 3989 4743
rect 4002 4747 4008 4748
rect 4002 4743 4003 4747
rect 4007 4746 4008 4747
rect 4167 4747 4173 4748
rect 4167 4746 4168 4747
rect 4007 4744 4168 4746
rect 4007 4743 4008 4744
rect 4002 4742 4008 4743
rect 4167 4743 4168 4744
rect 4172 4743 4173 4747
rect 4167 4742 4173 4743
rect 4391 4747 4397 4748
rect 4391 4743 4392 4747
rect 4396 4746 4397 4747
rect 4522 4747 4528 4748
rect 4522 4746 4523 4747
rect 4396 4744 4523 4746
rect 4396 4743 4397 4744
rect 4391 4742 4397 4743
rect 4522 4743 4523 4744
rect 4527 4743 4528 4747
rect 4522 4742 4528 4743
rect 4631 4747 4637 4748
rect 4631 4743 4632 4747
rect 4636 4746 4637 4747
rect 4770 4747 4776 4748
rect 4770 4746 4771 4747
rect 4636 4744 4771 4746
rect 4636 4743 4637 4744
rect 4631 4742 4637 4743
rect 4770 4743 4771 4744
rect 4775 4743 4776 4747
rect 4879 4747 4885 4748
rect 4879 4746 4880 4747
rect 4770 4742 4776 4743
rect 4819 4744 4880 4746
rect 4130 4739 4136 4740
rect 4130 4735 4131 4739
rect 4135 4738 4136 4739
rect 4819 4738 4821 4744
rect 4879 4743 4880 4744
rect 4884 4743 4885 4747
rect 4879 4742 4885 4743
rect 5135 4747 5141 4748
rect 5135 4743 5136 4747
rect 5140 4746 5141 4747
rect 5290 4747 5296 4748
rect 5290 4746 5291 4747
rect 5140 4744 5291 4746
rect 5140 4743 5141 4744
rect 5135 4742 5141 4743
rect 5290 4743 5291 4744
rect 5295 4743 5296 4747
rect 5290 4742 5296 4743
rect 5370 4747 5376 4748
rect 5370 4743 5371 4747
rect 5375 4746 5376 4747
rect 5399 4747 5405 4748
rect 5399 4746 5400 4747
rect 5375 4744 5400 4746
rect 5375 4743 5376 4744
rect 5370 4742 5376 4743
rect 5399 4743 5400 4744
rect 5404 4743 5405 4747
rect 5639 4747 5645 4748
rect 5639 4746 5640 4747
rect 5399 4742 5405 4743
rect 5408 4744 5640 4746
rect 4135 4736 4821 4738
rect 5098 4739 5104 4740
rect 4135 4735 4136 4736
rect 4130 4734 4136 4735
rect 5098 4735 5099 4739
rect 5103 4738 5104 4739
rect 5408 4738 5410 4744
rect 5639 4743 5640 4744
rect 5644 4743 5645 4747
rect 5639 4742 5645 4743
rect 5103 4736 5410 4738
rect 5103 4735 5104 4736
rect 5098 4734 5104 4735
rect 158 4732 164 4733
rect 110 4731 116 4732
rect 110 4727 111 4731
rect 115 4727 116 4731
rect 158 4728 159 4732
rect 163 4728 164 4732
rect 158 4727 164 4728
rect 294 4732 300 4733
rect 294 4728 295 4732
rect 299 4728 300 4732
rect 294 4727 300 4728
rect 430 4732 436 4733
rect 430 4728 431 4732
rect 435 4728 436 4732
rect 430 4727 436 4728
rect 566 4732 572 4733
rect 566 4728 567 4732
rect 571 4728 572 4732
rect 566 4727 572 4728
rect 702 4732 708 4733
rect 702 4728 703 4732
rect 707 4728 708 4732
rect 702 4727 708 4728
rect 1934 4731 1940 4732
rect 1934 4727 1935 4731
rect 1939 4727 1940 4731
rect 110 4726 116 4727
rect 1934 4726 1940 4727
rect 2146 4719 2152 4720
rect 2106 4715 2112 4716
rect 2106 4711 2107 4715
rect 2111 4711 2112 4715
rect 2146 4715 2147 4719
rect 2151 4718 2152 4719
rect 2322 4719 2328 4720
rect 2151 4716 2213 4718
rect 2151 4715 2152 4716
rect 2146 4714 2152 4715
rect 2322 4715 2323 4719
rect 2327 4718 2328 4719
rect 2666 4719 2672 4720
rect 2666 4718 2667 4719
rect 2327 4716 2389 4718
rect 2637 4716 2667 4718
rect 2327 4715 2328 4716
rect 2322 4714 2328 4715
rect 2666 4715 2667 4716
rect 2671 4715 2672 4719
rect 2666 4714 2672 4715
rect 2674 4719 2680 4720
rect 2674 4715 2675 4719
rect 2679 4718 2680 4719
rect 2679 4716 2741 4718
rect 2679 4715 2680 4716
rect 2674 4714 2680 4715
rect 4002 4715 4008 4716
rect 4002 4714 4003 4715
rect 3949 4712 4003 4714
rect 2106 4710 2112 4711
rect 4002 4711 4003 4712
rect 4007 4711 4008 4715
rect 4002 4710 4008 4711
rect 4130 4715 4136 4716
rect 4130 4711 4131 4715
rect 4135 4711 4136 4715
rect 4130 4710 4136 4711
rect 4138 4715 4144 4716
rect 4138 4711 4139 4715
rect 4143 4714 4144 4715
rect 4522 4715 4528 4716
rect 4143 4712 4285 4714
rect 4143 4711 4144 4712
rect 4138 4710 4144 4711
rect 4522 4711 4523 4715
rect 4527 4711 4528 4715
rect 4522 4710 4528 4711
rect 4770 4715 4776 4716
rect 4770 4711 4771 4715
rect 4775 4711 4776 4715
rect 4770 4710 4776 4711
rect 5098 4715 5104 4716
rect 5098 4711 5099 4715
rect 5103 4711 5104 4715
rect 5098 4710 5104 4711
rect 5290 4715 5296 4716
rect 5290 4711 5291 4715
rect 5295 4711 5296 4715
rect 5290 4710 5296 4711
rect 5602 4715 5608 4716
rect 5602 4711 5603 4715
rect 5607 4711 5608 4715
rect 5602 4710 5608 4711
rect 2143 4683 2152 4684
rect 2143 4679 2144 4683
rect 2151 4679 2152 4683
rect 2143 4678 2152 4679
rect 2319 4683 2328 4684
rect 2319 4679 2320 4683
rect 2327 4679 2328 4683
rect 2319 4678 2328 4679
rect 2386 4683 2392 4684
rect 2386 4679 2387 4683
rect 2391 4682 2392 4683
rect 2495 4683 2501 4684
rect 2495 4682 2496 4683
rect 2391 4680 2496 4682
rect 2391 4679 2392 4680
rect 2386 4678 2392 4679
rect 2495 4679 2496 4680
rect 2500 4679 2501 4683
rect 2495 4678 2501 4679
rect 2671 4683 2680 4684
rect 2671 4679 2672 4683
rect 2679 4679 2680 4683
rect 2671 4678 2680 4679
rect 2834 4683 2840 4684
rect 2834 4679 2835 4683
rect 2839 4682 2840 4683
rect 2847 4683 2853 4684
rect 2847 4682 2848 4683
rect 2839 4680 2848 4682
rect 2839 4679 2840 4680
rect 2834 4678 2840 4679
rect 2847 4679 2848 4680
rect 2852 4679 2853 4683
rect 2847 4678 2853 4679
rect 1974 4676 1980 4677
rect 3798 4676 3804 4677
rect 1974 4672 1975 4676
rect 1979 4672 1980 4676
rect 1974 4671 1980 4672
rect 2018 4675 2024 4676
rect 2018 4671 2019 4675
rect 2023 4671 2024 4675
rect 2018 4670 2024 4671
rect 2194 4675 2200 4676
rect 2194 4671 2195 4675
rect 2199 4671 2200 4675
rect 2194 4670 2200 4671
rect 2370 4675 2376 4676
rect 2370 4671 2371 4675
rect 2375 4671 2376 4675
rect 2370 4670 2376 4671
rect 2546 4675 2552 4676
rect 2546 4671 2547 4675
rect 2551 4671 2552 4675
rect 2546 4670 2552 4671
rect 2722 4675 2728 4676
rect 2722 4671 2723 4675
rect 2727 4671 2728 4675
rect 3798 4672 3799 4676
rect 3803 4672 3804 4676
rect 3798 4671 3804 4672
rect 2722 4670 2728 4671
rect 110 4669 116 4670
rect 1934 4669 1940 4670
rect 110 4665 111 4669
rect 115 4665 116 4669
rect 110 4664 116 4665
rect 158 4668 164 4669
rect 158 4664 159 4668
rect 163 4664 164 4668
rect 158 4663 164 4664
rect 294 4668 300 4669
rect 294 4664 295 4668
rect 299 4664 300 4668
rect 294 4663 300 4664
rect 430 4668 436 4669
rect 430 4664 431 4668
rect 435 4664 436 4668
rect 430 4663 436 4664
rect 566 4668 572 4669
rect 566 4664 567 4668
rect 571 4664 572 4668
rect 566 4663 572 4664
rect 702 4668 708 4669
rect 702 4664 703 4668
rect 707 4664 708 4668
rect 1934 4665 1935 4669
rect 1939 4665 1940 4669
rect 1934 4664 1940 4665
rect 3778 4667 3784 4668
rect 702 4663 708 4664
rect 3778 4663 3779 4667
rect 3783 4666 3784 4667
rect 3986 4667 3992 4668
rect 3783 4664 3877 4666
rect 3783 4663 3784 4664
rect 3778 4662 3784 4663
rect 3986 4663 3987 4667
rect 3991 4666 3992 4667
rect 4258 4667 4264 4668
rect 3991 4664 4013 4666
rect 3991 4663 3992 4664
rect 3986 4662 3992 4663
rect 4218 4663 4224 4664
rect 2046 4660 2052 4661
rect 1974 4659 1980 4660
rect 1974 4655 1975 4659
rect 1979 4655 1980 4659
rect 2046 4656 2047 4660
rect 2051 4656 2052 4660
rect 2046 4655 2052 4656
rect 2222 4660 2228 4661
rect 2222 4656 2223 4660
rect 2227 4656 2228 4660
rect 2222 4655 2228 4656
rect 2398 4660 2404 4661
rect 2398 4656 2399 4660
rect 2403 4656 2404 4660
rect 2398 4655 2404 4656
rect 2574 4660 2580 4661
rect 2574 4656 2575 4660
rect 2579 4656 2580 4660
rect 2574 4655 2580 4656
rect 2750 4660 2756 4661
rect 2750 4656 2751 4660
rect 2755 4656 2756 4660
rect 2750 4655 2756 4656
rect 3798 4659 3804 4660
rect 3798 4655 3799 4659
rect 3803 4655 3804 4659
rect 4218 4659 4219 4663
rect 4223 4659 4224 4663
rect 4258 4663 4259 4667
rect 4263 4666 4264 4667
rect 4394 4667 4400 4668
rect 4263 4664 4285 4666
rect 4263 4663 4264 4664
rect 4258 4662 4264 4663
rect 4394 4663 4395 4667
rect 4399 4666 4400 4667
rect 4671 4667 4677 4668
rect 4671 4666 4672 4667
rect 4399 4664 4421 4666
rect 4629 4664 4672 4666
rect 4399 4663 4400 4664
rect 4394 4662 4400 4663
rect 4671 4663 4672 4664
rect 4676 4663 4677 4667
rect 4807 4667 4813 4668
rect 4807 4666 4808 4667
rect 4765 4664 4808 4666
rect 4671 4662 4677 4663
rect 4807 4663 4808 4664
rect 4812 4663 4813 4667
rect 4959 4667 4965 4668
rect 4959 4666 4960 4667
rect 4909 4664 4960 4666
rect 4807 4662 4813 4663
rect 4959 4663 4960 4664
rect 4964 4663 4965 4667
rect 5103 4667 5109 4668
rect 5103 4666 5104 4667
rect 5053 4664 5104 4666
rect 4959 4662 4965 4663
rect 5103 4663 5104 4664
rect 5108 4663 5109 4667
rect 5239 4667 5245 4668
rect 5239 4666 5240 4667
rect 5197 4664 5240 4666
rect 5103 4662 5109 4663
rect 5239 4663 5240 4664
rect 5244 4663 5245 4667
rect 5370 4667 5376 4668
rect 5239 4662 5245 4663
rect 5330 4663 5336 4664
rect 4218 4658 4224 4659
rect 5330 4659 5331 4663
rect 5335 4659 5336 4663
rect 5370 4663 5371 4667
rect 5375 4666 5376 4667
rect 5511 4667 5517 4668
rect 5375 4664 5397 4666
rect 5375 4663 5376 4664
rect 5370 4662 5376 4663
rect 5511 4663 5512 4667
rect 5516 4666 5517 4667
rect 5516 4664 5533 4666
rect 5516 4663 5517 4664
rect 5511 4662 5517 4663
rect 5330 4658 5336 4659
rect 1974 4654 1980 4655
rect 3798 4654 3804 4655
rect 130 4653 136 4654
rect 110 4652 116 4653
rect 110 4648 111 4652
rect 115 4648 116 4652
rect 130 4649 131 4653
rect 135 4649 136 4653
rect 130 4648 136 4649
rect 266 4653 272 4654
rect 266 4649 267 4653
rect 271 4649 272 4653
rect 266 4648 272 4649
rect 402 4653 408 4654
rect 402 4649 403 4653
rect 407 4649 408 4653
rect 402 4648 408 4649
rect 538 4653 544 4654
rect 538 4649 539 4653
rect 543 4649 544 4653
rect 538 4648 544 4649
rect 674 4653 680 4654
rect 674 4649 675 4653
rect 679 4649 680 4653
rect 674 4648 680 4649
rect 1934 4652 1940 4653
rect 1934 4648 1935 4652
rect 1939 4648 1940 4652
rect 110 4647 116 4648
rect 1934 4647 1940 4648
rect 255 4643 261 4644
rect 255 4639 256 4643
rect 260 4642 261 4643
rect 282 4643 288 4644
rect 282 4642 283 4643
rect 260 4640 283 4642
rect 260 4639 261 4640
rect 255 4638 261 4639
rect 282 4639 283 4640
rect 287 4639 288 4643
rect 282 4638 288 4639
rect 391 4643 397 4644
rect 391 4639 392 4643
rect 396 4642 397 4643
rect 418 4643 424 4644
rect 418 4642 419 4643
rect 396 4640 419 4642
rect 396 4639 397 4640
rect 391 4638 397 4639
rect 418 4639 419 4640
rect 423 4639 424 4643
rect 418 4638 424 4639
rect 527 4643 533 4644
rect 527 4639 528 4643
rect 532 4642 533 4643
rect 554 4643 560 4644
rect 554 4642 555 4643
rect 532 4640 555 4642
rect 532 4639 533 4640
rect 527 4638 533 4639
rect 554 4639 555 4640
rect 559 4639 560 4643
rect 554 4638 560 4639
rect 663 4643 669 4644
rect 663 4639 664 4643
rect 668 4642 669 4643
rect 690 4643 696 4644
rect 690 4642 691 4643
rect 668 4640 691 4642
rect 668 4639 669 4640
rect 663 4638 669 4639
rect 690 4639 691 4640
rect 695 4639 696 4643
rect 690 4638 696 4639
rect 754 4643 760 4644
rect 754 4639 755 4643
rect 759 4642 760 4643
rect 799 4643 805 4644
rect 799 4642 800 4643
rect 759 4640 800 4642
rect 759 4639 760 4640
rect 754 4638 760 4639
rect 799 4639 800 4640
rect 804 4639 805 4643
rect 799 4638 805 4639
rect 4218 4639 4224 4640
rect 4218 4635 4219 4639
rect 4223 4638 4224 4639
rect 5330 4639 5336 4640
rect 4223 4636 4667 4638
rect 4223 4635 4224 4636
rect 4218 4634 4224 4635
rect 4665 4632 4667 4636
rect 5330 4635 5331 4639
rect 5335 4638 5336 4639
rect 5335 4636 5542 4638
rect 5335 4635 5336 4636
rect 5330 4634 5336 4635
rect 3983 4631 3992 4632
rect 3983 4627 3984 4631
rect 3991 4627 3992 4631
rect 3983 4626 3992 4627
rect 4119 4631 4125 4632
rect 4119 4627 4120 4631
rect 4124 4630 4125 4631
rect 4138 4631 4144 4632
rect 4138 4630 4139 4631
rect 4124 4628 4139 4630
rect 4124 4627 4125 4628
rect 4119 4626 4125 4627
rect 4138 4627 4139 4628
rect 4143 4627 4144 4631
rect 4138 4626 4144 4627
rect 4255 4631 4264 4632
rect 4255 4627 4256 4631
rect 4263 4627 4264 4631
rect 4255 4626 4264 4627
rect 4391 4631 4400 4632
rect 4391 4627 4392 4631
rect 4399 4627 4400 4631
rect 4391 4626 4400 4627
rect 4527 4631 4533 4632
rect 4527 4627 4528 4631
rect 4532 4630 4533 4631
rect 4594 4631 4600 4632
rect 4594 4630 4595 4631
rect 4532 4628 4595 4630
rect 4532 4627 4533 4628
rect 4527 4626 4533 4627
rect 4594 4627 4595 4628
rect 4599 4627 4600 4631
rect 4594 4626 4600 4627
rect 4663 4631 4669 4632
rect 4663 4627 4664 4631
rect 4668 4627 4669 4631
rect 4663 4626 4669 4627
rect 4671 4631 4677 4632
rect 4671 4627 4672 4631
rect 4676 4630 4677 4631
rect 4799 4631 4805 4632
rect 4799 4630 4800 4631
rect 4676 4628 4800 4630
rect 4676 4627 4677 4628
rect 4671 4626 4677 4627
rect 4799 4627 4800 4628
rect 4804 4627 4805 4631
rect 4799 4626 4805 4627
rect 4807 4631 4813 4632
rect 4807 4627 4808 4631
rect 4812 4630 4813 4631
rect 4943 4631 4949 4632
rect 4943 4630 4944 4631
rect 4812 4628 4944 4630
rect 4812 4627 4813 4628
rect 4807 4626 4813 4627
rect 4943 4627 4944 4628
rect 4948 4627 4949 4631
rect 4943 4626 4949 4627
rect 4959 4631 4965 4632
rect 4959 4627 4960 4631
rect 4964 4630 4965 4631
rect 5087 4631 5093 4632
rect 5087 4630 5088 4631
rect 4964 4628 5088 4630
rect 4964 4627 4965 4628
rect 4959 4626 4965 4627
rect 5087 4627 5088 4628
rect 5092 4627 5093 4631
rect 5087 4626 5093 4627
rect 5103 4631 5109 4632
rect 5103 4627 5104 4631
rect 5108 4630 5109 4631
rect 5231 4631 5237 4632
rect 5231 4630 5232 4631
rect 5108 4628 5232 4630
rect 5108 4627 5109 4628
rect 5103 4626 5109 4627
rect 5231 4627 5232 4628
rect 5236 4627 5237 4631
rect 5231 4626 5237 4627
rect 5239 4631 5245 4632
rect 5239 4627 5240 4631
rect 5244 4630 5245 4631
rect 5367 4631 5373 4632
rect 5367 4630 5368 4631
rect 5244 4628 5368 4630
rect 5244 4627 5245 4628
rect 5239 4626 5245 4627
rect 5367 4627 5368 4628
rect 5372 4627 5373 4631
rect 5367 4626 5373 4627
rect 5503 4631 5509 4632
rect 5503 4627 5504 4631
rect 5508 4630 5509 4631
rect 5511 4631 5517 4632
rect 5511 4630 5512 4631
rect 5508 4628 5512 4630
rect 5508 4627 5509 4628
rect 5503 4626 5509 4627
rect 5511 4627 5512 4628
rect 5516 4627 5517 4631
rect 5540 4630 5542 4636
rect 5639 4631 5645 4632
rect 5639 4630 5640 4631
rect 5540 4628 5640 4630
rect 5511 4626 5517 4627
rect 5639 4627 5640 4628
rect 5644 4627 5645 4631
rect 5639 4626 5645 4627
rect 3838 4624 3844 4625
rect 5662 4624 5668 4625
rect 3838 4620 3839 4624
rect 3843 4620 3844 4624
rect 3838 4619 3844 4620
rect 3858 4623 3864 4624
rect 3858 4619 3859 4623
rect 3863 4619 3864 4623
rect 3858 4618 3864 4619
rect 3994 4623 4000 4624
rect 3994 4619 3995 4623
rect 3999 4619 4000 4623
rect 3994 4618 4000 4619
rect 4130 4623 4136 4624
rect 4130 4619 4131 4623
rect 4135 4619 4136 4623
rect 4130 4618 4136 4619
rect 4266 4623 4272 4624
rect 4266 4619 4267 4623
rect 4271 4619 4272 4623
rect 4266 4618 4272 4619
rect 4402 4623 4408 4624
rect 4402 4619 4403 4623
rect 4407 4619 4408 4623
rect 4402 4618 4408 4619
rect 4538 4623 4544 4624
rect 4538 4619 4539 4623
rect 4543 4619 4544 4623
rect 4538 4618 4544 4619
rect 4674 4623 4680 4624
rect 4674 4619 4675 4623
rect 4679 4619 4680 4623
rect 4674 4618 4680 4619
rect 4818 4623 4824 4624
rect 4818 4619 4819 4623
rect 4823 4619 4824 4623
rect 4818 4618 4824 4619
rect 4962 4623 4968 4624
rect 4962 4619 4963 4623
rect 4967 4619 4968 4623
rect 4962 4618 4968 4619
rect 5106 4623 5112 4624
rect 5106 4619 5107 4623
rect 5111 4619 5112 4623
rect 5106 4618 5112 4619
rect 5242 4623 5248 4624
rect 5242 4619 5243 4623
rect 5247 4619 5248 4623
rect 5242 4618 5248 4619
rect 5378 4623 5384 4624
rect 5378 4619 5379 4623
rect 5383 4619 5384 4623
rect 5378 4618 5384 4619
rect 5514 4623 5520 4624
rect 5514 4619 5515 4623
rect 5519 4619 5520 4623
rect 5662 4620 5663 4624
rect 5667 4620 5668 4624
rect 5662 4619 5668 4620
rect 5514 4618 5520 4619
rect 218 4611 224 4612
rect 218 4607 219 4611
rect 223 4607 224 4611
rect 218 4606 224 4607
rect 282 4611 288 4612
rect 282 4607 283 4611
rect 287 4607 288 4611
rect 282 4606 288 4607
rect 418 4611 424 4612
rect 418 4607 419 4611
rect 423 4607 424 4611
rect 418 4606 424 4607
rect 554 4611 560 4612
rect 554 4607 555 4611
rect 559 4607 560 4611
rect 554 4606 560 4607
rect 690 4611 696 4612
rect 690 4607 691 4611
rect 695 4607 696 4611
rect 3886 4608 3892 4609
rect 690 4606 696 4607
rect 3838 4607 3844 4608
rect 3838 4603 3839 4607
rect 3843 4603 3844 4607
rect 3886 4604 3887 4608
rect 3891 4604 3892 4608
rect 3886 4603 3892 4604
rect 4022 4608 4028 4609
rect 4022 4604 4023 4608
rect 4027 4604 4028 4608
rect 4022 4603 4028 4604
rect 4158 4608 4164 4609
rect 4158 4604 4159 4608
rect 4163 4604 4164 4608
rect 4158 4603 4164 4604
rect 4294 4608 4300 4609
rect 4294 4604 4295 4608
rect 4299 4604 4300 4608
rect 4294 4603 4300 4604
rect 4430 4608 4436 4609
rect 4430 4604 4431 4608
rect 4435 4604 4436 4608
rect 4430 4603 4436 4604
rect 4566 4608 4572 4609
rect 4566 4604 4567 4608
rect 4571 4604 4572 4608
rect 4566 4603 4572 4604
rect 4702 4608 4708 4609
rect 4702 4604 4703 4608
rect 4707 4604 4708 4608
rect 4702 4603 4708 4604
rect 4846 4608 4852 4609
rect 4846 4604 4847 4608
rect 4851 4604 4852 4608
rect 4846 4603 4852 4604
rect 4990 4608 4996 4609
rect 4990 4604 4991 4608
rect 4995 4604 4996 4608
rect 4990 4603 4996 4604
rect 5134 4608 5140 4609
rect 5134 4604 5135 4608
rect 5139 4604 5140 4608
rect 5134 4603 5140 4604
rect 5270 4608 5276 4609
rect 5270 4604 5271 4608
rect 5275 4604 5276 4608
rect 5270 4603 5276 4604
rect 5406 4608 5412 4609
rect 5406 4604 5407 4608
rect 5411 4604 5412 4608
rect 5406 4603 5412 4604
rect 5542 4608 5548 4609
rect 5542 4604 5543 4608
rect 5547 4604 5548 4608
rect 5542 4603 5548 4604
rect 5662 4607 5668 4608
rect 5662 4603 5663 4607
rect 5667 4603 5668 4607
rect 3838 4602 3844 4603
rect 5662 4602 5668 4603
rect 1974 4597 1980 4598
rect 3798 4597 3804 4598
rect 1974 4593 1975 4597
rect 1979 4593 1980 4597
rect 1974 4592 1980 4593
rect 2022 4596 2028 4597
rect 2022 4592 2023 4596
rect 2027 4592 2028 4596
rect 2022 4591 2028 4592
rect 2262 4596 2268 4597
rect 2262 4592 2263 4596
rect 2267 4592 2268 4596
rect 2262 4591 2268 4592
rect 2526 4596 2532 4597
rect 2526 4592 2527 4596
rect 2531 4592 2532 4596
rect 2526 4591 2532 4592
rect 2774 4596 2780 4597
rect 2774 4592 2775 4596
rect 2779 4592 2780 4596
rect 2774 4591 2780 4592
rect 3014 4596 3020 4597
rect 3014 4592 3015 4596
rect 3019 4592 3020 4596
rect 3014 4591 3020 4592
rect 3246 4596 3252 4597
rect 3246 4592 3247 4596
rect 3251 4592 3252 4596
rect 3246 4591 3252 4592
rect 3470 4596 3476 4597
rect 3470 4592 3471 4596
rect 3475 4592 3476 4596
rect 3470 4591 3476 4592
rect 3678 4596 3684 4597
rect 3678 4592 3679 4596
rect 3683 4592 3684 4596
rect 3798 4593 3799 4597
rect 3803 4593 3804 4597
rect 3798 4592 3804 4593
rect 3678 4591 3684 4592
rect 1994 4581 2000 4582
rect 1974 4580 1980 4581
rect 1974 4576 1975 4580
rect 1979 4576 1980 4580
rect 1994 4577 1995 4581
rect 1999 4577 2000 4581
rect 1994 4576 2000 4577
rect 2234 4581 2240 4582
rect 2234 4577 2235 4581
rect 2239 4577 2240 4581
rect 2234 4576 2240 4577
rect 2498 4581 2504 4582
rect 2498 4577 2499 4581
rect 2503 4577 2504 4581
rect 2498 4576 2504 4577
rect 2746 4581 2752 4582
rect 2746 4577 2747 4581
rect 2751 4577 2752 4581
rect 2746 4576 2752 4577
rect 2986 4581 2992 4582
rect 2986 4577 2987 4581
rect 2991 4577 2992 4581
rect 2986 4576 2992 4577
rect 3218 4581 3224 4582
rect 3218 4577 3219 4581
rect 3223 4577 3224 4581
rect 3218 4576 3224 4577
rect 3442 4581 3448 4582
rect 3442 4577 3443 4581
rect 3447 4577 3448 4581
rect 3442 4576 3448 4577
rect 3650 4581 3656 4582
rect 3650 4577 3651 4581
rect 3655 4577 3656 4581
rect 3650 4576 3656 4577
rect 3798 4580 3804 4581
rect 3798 4576 3799 4580
rect 3803 4576 3804 4580
rect 1974 4575 1980 4576
rect 3798 4575 3804 4576
rect 578 4571 584 4572
rect 578 4567 579 4571
rect 583 4570 584 4571
rect 1222 4571 1228 4572
rect 1222 4570 1223 4571
rect 583 4568 1223 4570
rect 583 4567 584 4568
rect 578 4566 584 4567
rect 1222 4567 1223 4568
rect 1227 4567 1228 4571
rect 1222 4566 1228 4567
rect 2106 4571 2112 4572
rect 2106 4567 2107 4571
rect 2111 4570 2112 4571
rect 2119 4571 2125 4572
rect 2119 4570 2120 4571
rect 2111 4568 2120 4570
rect 2111 4567 2112 4568
rect 2106 4566 2112 4567
rect 2119 4567 2120 4568
rect 2124 4567 2125 4571
rect 2119 4566 2125 4567
rect 2359 4571 2365 4572
rect 2359 4567 2360 4571
rect 2364 4570 2365 4571
rect 2514 4571 2520 4572
rect 2514 4570 2515 4571
rect 2364 4568 2515 4570
rect 2364 4567 2365 4568
rect 2359 4566 2365 4567
rect 2514 4567 2515 4568
rect 2519 4567 2520 4571
rect 2514 4566 2520 4567
rect 2618 4571 2629 4572
rect 2618 4567 2619 4571
rect 2623 4567 2624 4571
rect 2628 4567 2629 4571
rect 2871 4571 2877 4572
rect 2871 4570 2872 4571
rect 2618 4566 2629 4567
rect 2632 4568 2872 4570
rect 754 4563 760 4564
rect 754 4562 755 4563
rect 368 4560 755 4562
rect 368 4550 370 4560
rect 754 4559 755 4560
rect 759 4559 760 4563
rect 754 4558 760 4559
rect 2322 4563 2328 4564
rect 2322 4559 2323 4563
rect 2327 4562 2328 4563
rect 2632 4562 2634 4568
rect 2871 4567 2872 4568
rect 2876 4567 2877 4571
rect 2871 4566 2877 4567
rect 3111 4571 3117 4572
rect 3111 4567 3112 4571
rect 3116 4570 3117 4571
rect 3234 4571 3240 4572
rect 3234 4570 3235 4571
rect 3116 4568 3235 4570
rect 3116 4567 3117 4568
rect 3111 4566 3117 4567
rect 3234 4567 3235 4568
rect 3239 4567 3240 4571
rect 3234 4566 3240 4567
rect 3343 4571 3349 4572
rect 3343 4567 3344 4571
rect 3348 4570 3349 4571
rect 3458 4571 3464 4572
rect 3458 4570 3459 4571
rect 3348 4568 3459 4570
rect 3348 4567 3349 4568
rect 3343 4566 3349 4567
rect 3458 4567 3459 4568
rect 3463 4567 3464 4571
rect 3458 4566 3464 4567
rect 3567 4571 3573 4572
rect 3567 4567 3568 4571
rect 3572 4570 3573 4571
rect 3666 4571 3672 4572
rect 3666 4570 3667 4571
rect 3572 4568 3667 4570
rect 3572 4567 3573 4568
rect 3567 4566 3573 4567
rect 3666 4567 3667 4568
rect 3671 4567 3672 4571
rect 3666 4566 3672 4567
rect 3775 4571 3784 4572
rect 3775 4567 3776 4571
rect 3783 4567 3784 4571
rect 3775 4566 3784 4567
rect 2327 4560 2634 4562
rect 2327 4559 2328 4560
rect 2322 4558 2328 4559
rect 341 4548 370 4550
rect 378 4551 384 4552
rect 378 4547 379 4551
rect 383 4550 384 4551
rect 566 4551 572 4552
rect 383 4548 461 4550
rect 383 4547 384 4548
rect 378 4546 384 4547
rect 566 4547 567 4551
rect 571 4550 572 4551
rect 778 4551 784 4552
rect 571 4548 669 4550
rect 571 4547 572 4548
rect 566 4546 572 4547
rect 778 4547 779 4551
rect 783 4550 784 4551
rect 1002 4551 1008 4552
rect 783 4548 893 4550
rect 783 4547 784 4548
rect 778 4546 784 4547
rect 1002 4547 1003 4551
rect 1007 4550 1008 4551
rect 1522 4551 1528 4552
rect 1007 4548 1117 4550
rect 1007 4547 1008 4548
rect 1002 4546 1008 4547
rect 1522 4547 1523 4551
rect 1527 4550 1528 4551
rect 1703 4551 1709 4552
rect 1527 4548 1589 4550
rect 1527 4547 1528 4548
rect 1522 4546 1528 4547
rect 1703 4547 1704 4551
rect 1708 4550 1709 4551
rect 1708 4548 1805 4550
rect 3838 4549 3844 4550
rect 5662 4549 5668 4550
rect 1708 4547 1709 4548
rect 1703 4546 1709 4547
rect 3838 4545 3839 4549
rect 3843 4545 3844 4549
rect 1416 4542 1418 4545
rect 3838 4544 3844 4545
rect 4670 4548 4676 4549
rect 4670 4544 4671 4548
rect 4675 4544 4676 4548
rect 1562 4543 1568 4544
rect 4670 4543 4676 4544
rect 4806 4548 4812 4549
rect 4806 4544 4807 4548
rect 4811 4544 4812 4548
rect 4806 4543 4812 4544
rect 4942 4548 4948 4549
rect 4942 4544 4943 4548
rect 4947 4544 4948 4548
rect 4942 4543 4948 4544
rect 5078 4548 5084 4549
rect 5078 4544 5079 4548
rect 5083 4544 5084 4548
rect 5662 4545 5663 4549
rect 5667 4545 5668 4549
rect 5662 4544 5668 4545
rect 5078 4543 5084 4544
rect 1562 4542 1563 4543
rect 1416 4540 1563 4542
rect 1562 4539 1563 4540
rect 1567 4539 1568 4543
rect 1562 4538 1568 4539
rect 2010 4539 2016 4540
rect 2010 4535 2011 4539
rect 2015 4535 2016 4539
rect 2010 4534 2016 4535
rect 2322 4539 2328 4540
rect 2322 4535 2323 4539
rect 2327 4535 2328 4539
rect 2322 4534 2328 4535
rect 2514 4539 2520 4540
rect 2514 4535 2515 4539
rect 2519 4535 2520 4539
rect 2514 4534 2520 4535
rect 2834 4539 2840 4540
rect 2834 4535 2835 4539
rect 2839 4535 2840 4539
rect 2834 4534 2840 4535
rect 3074 4539 3080 4540
rect 3074 4535 3075 4539
rect 3079 4535 3080 4539
rect 3074 4534 3080 4535
rect 3234 4539 3240 4540
rect 3234 4535 3235 4539
rect 3239 4535 3240 4539
rect 3234 4534 3240 4535
rect 3458 4539 3464 4540
rect 3458 4535 3459 4539
rect 3463 4535 3464 4539
rect 3458 4534 3464 4535
rect 3666 4539 3672 4540
rect 3666 4535 3667 4539
rect 3671 4535 3672 4539
rect 3666 4534 3672 4535
rect 4642 4533 4648 4534
rect 3838 4532 3844 4533
rect 3838 4528 3839 4532
rect 3843 4528 3844 4532
rect 4642 4529 4643 4533
rect 4647 4529 4648 4533
rect 4642 4528 4648 4529
rect 4778 4533 4784 4534
rect 4778 4529 4779 4533
rect 4783 4529 4784 4533
rect 4778 4528 4784 4529
rect 4914 4533 4920 4534
rect 4914 4529 4915 4533
rect 4919 4529 4920 4533
rect 4914 4528 4920 4529
rect 5050 4533 5056 4534
rect 5050 4529 5051 4533
rect 5055 4529 5056 4533
rect 5050 4528 5056 4529
rect 5662 4532 5668 4533
rect 5662 4528 5663 4532
rect 5667 4528 5668 4532
rect 3838 4527 3844 4528
rect 5662 4527 5668 4528
rect 4767 4523 4773 4524
rect 4767 4519 4768 4523
rect 4772 4522 4773 4523
rect 4794 4523 4800 4524
rect 4794 4522 4795 4523
rect 4772 4520 4795 4522
rect 4772 4519 4773 4520
rect 4767 4518 4773 4519
rect 4794 4519 4795 4520
rect 4799 4519 4800 4523
rect 4794 4518 4800 4519
rect 4903 4523 4909 4524
rect 4903 4519 4904 4523
rect 4908 4522 4909 4523
rect 4930 4523 4936 4524
rect 4930 4522 4931 4523
rect 4908 4520 4931 4522
rect 4908 4519 4909 4520
rect 4903 4518 4909 4519
rect 4930 4519 4931 4520
rect 4935 4519 4936 4523
rect 4930 4518 4936 4519
rect 5039 4523 5045 4524
rect 5039 4519 5040 4523
rect 5044 4522 5045 4523
rect 5066 4523 5072 4524
rect 5066 4522 5067 4523
rect 5044 4520 5067 4522
rect 5044 4519 5045 4520
rect 5039 4518 5045 4519
rect 5066 4519 5067 4520
rect 5071 4519 5072 4523
rect 5066 4518 5072 4519
rect 5074 4523 5080 4524
rect 5074 4519 5075 4523
rect 5079 4522 5080 4523
rect 5175 4523 5181 4524
rect 5175 4522 5176 4523
rect 5079 4520 5176 4522
rect 5079 4519 5080 4520
rect 5074 4518 5080 4519
rect 5175 4519 5176 4520
rect 5180 4519 5181 4523
rect 5175 4518 5181 4519
rect 375 4515 384 4516
rect 375 4511 376 4515
rect 383 4511 384 4515
rect 375 4510 384 4511
rect 566 4515 573 4516
rect 566 4511 567 4515
rect 572 4511 573 4515
rect 566 4510 573 4511
rect 775 4515 784 4516
rect 775 4511 776 4515
rect 783 4511 784 4515
rect 775 4510 784 4511
rect 999 4515 1008 4516
rect 999 4511 1000 4515
rect 1007 4511 1008 4515
rect 999 4510 1008 4511
rect 1222 4515 1229 4516
rect 1222 4511 1223 4515
rect 1228 4511 1229 4515
rect 1222 4510 1229 4511
rect 1455 4515 1461 4516
rect 1455 4511 1456 4515
rect 1460 4514 1461 4515
rect 1522 4515 1528 4516
rect 1522 4514 1523 4515
rect 1460 4512 1523 4514
rect 1460 4511 1461 4512
rect 1455 4510 1461 4511
rect 1522 4511 1523 4512
rect 1527 4511 1528 4515
rect 1522 4510 1528 4511
rect 1695 4515 1701 4516
rect 1695 4511 1696 4515
rect 1700 4514 1701 4515
rect 1703 4515 1709 4516
rect 1703 4514 1704 4515
rect 1700 4512 1704 4514
rect 1700 4511 1701 4512
rect 1695 4510 1701 4511
rect 1703 4511 1704 4512
rect 1708 4511 1709 4515
rect 1703 4510 1709 4511
rect 1911 4515 1917 4516
rect 1911 4511 1912 4515
rect 1916 4514 1917 4515
rect 2010 4515 2016 4516
rect 2010 4514 2011 4515
rect 1916 4512 2011 4514
rect 1916 4511 1917 4512
rect 1911 4510 1917 4511
rect 2010 4511 2011 4512
rect 2015 4511 2016 4515
rect 2010 4510 2016 4511
rect 110 4508 116 4509
rect 1934 4508 1940 4509
rect 110 4504 111 4508
rect 115 4504 116 4508
rect 110 4503 116 4504
rect 250 4507 256 4508
rect 250 4503 251 4507
rect 255 4503 256 4507
rect 250 4502 256 4503
rect 442 4507 448 4508
rect 442 4503 443 4507
rect 447 4503 448 4507
rect 442 4502 448 4503
rect 650 4507 656 4508
rect 650 4503 651 4507
rect 655 4503 656 4507
rect 650 4502 656 4503
rect 874 4507 880 4508
rect 874 4503 875 4507
rect 879 4503 880 4507
rect 874 4502 880 4503
rect 1098 4507 1104 4508
rect 1098 4503 1099 4507
rect 1103 4503 1104 4507
rect 1098 4502 1104 4503
rect 1330 4507 1336 4508
rect 1330 4503 1331 4507
rect 1335 4503 1336 4507
rect 1330 4502 1336 4503
rect 1570 4507 1576 4508
rect 1570 4503 1571 4507
rect 1575 4503 1576 4507
rect 1570 4502 1576 4503
rect 1786 4507 1792 4508
rect 1786 4503 1787 4507
rect 1791 4503 1792 4507
rect 1934 4504 1935 4508
rect 1939 4504 1940 4508
rect 1934 4503 1940 4504
rect 1786 4502 1792 4503
rect 278 4492 284 4493
rect 110 4491 116 4492
rect 110 4487 111 4491
rect 115 4487 116 4491
rect 278 4488 279 4492
rect 283 4488 284 4492
rect 278 4487 284 4488
rect 470 4492 476 4493
rect 470 4488 471 4492
rect 475 4488 476 4492
rect 470 4487 476 4488
rect 678 4492 684 4493
rect 678 4488 679 4492
rect 683 4488 684 4492
rect 678 4487 684 4488
rect 902 4492 908 4493
rect 902 4488 903 4492
rect 907 4488 908 4492
rect 902 4487 908 4488
rect 1126 4492 1132 4493
rect 1126 4488 1127 4492
rect 1131 4488 1132 4492
rect 1126 4487 1132 4488
rect 1358 4492 1364 4493
rect 1358 4488 1359 4492
rect 1363 4488 1364 4492
rect 1358 4487 1364 4488
rect 1598 4492 1604 4493
rect 1598 4488 1599 4492
rect 1603 4488 1604 4492
rect 1598 4487 1604 4488
rect 1814 4492 1820 4493
rect 1814 4488 1815 4492
rect 1819 4488 1820 4492
rect 1814 4487 1820 4488
rect 1934 4491 1940 4492
rect 1934 4487 1935 4491
rect 1939 4487 1940 4491
rect 110 4486 116 4487
rect 1934 4486 1940 4487
rect 4594 4491 4600 4492
rect 4594 4487 4595 4491
rect 4599 4490 4600 4491
rect 4794 4491 4800 4492
rect 4599 4488 4661 4490
rect 4599 4487 4600 4488
rect 4594 4486 4600 4487
rect 4794 4487 4795 4491
rect 4799 4487 4800 4491
rect 4794 4486 4800 4487
rect 4930 4491 4936 4492
rect 4930 4487 4931 4491
rect 4935 4487 4936 4491
rect 4930 4486 4936 4487
rect 5066 4491 5072 4492
rect 5066 4487 5067 4491
rect 5071 4487 5072 4491
rect 5066 4486 5072 4487
rect 2494 4479 2500 4480
rect 2494 4478 2495 4479
rect 2357 4476 2495 4478
rect 2494 4475 2495 4476
rect 2499 4475 2500 4479
rect 2618 4479 2624 4480
rect 2618 4478 2619 4479
rect 2605 4476 2619 4478
rect 2494 4474 2500 4475
rect 2618 4475 2619 4476
rect 2623 4475 2624 4479
rect 2874 4479 2880 4480
rect 2618 4474 2624 4475
rect 2834 4475 2840 4476
rect 2834 4471 2835 4475
rect 2839 4471 2840 4475
rect 2874 4475 2875 4479
rect 2879 4478 2880 4479
rect 3098 4479 3104 4480
rect 2879 4476 2989 4478
rect 2879 4475 2880 4476
rect 2874 4474 2880 4475
rect 3098 4475 3099 4479
rect 3103 4478 3104 4479
rect 3314 4479 3320 4480
rect 3103 4476 3205 4478
rect 3103 4475 3104 4476
rect 3098 4474 3104 4475
rect 3314 4475 3315 4479
rect 3319 4478 3320 4479
rect 3522 4479 3528 4480
rect 3319 4476 3413 4478
rect 3319 4475 3320 4476
rect 3314 4474 3320 4475
rect 3522 4475 3523 4479
rect 3527 4478 3528 4479
rect 3527 4476 3629 4478
rect 3527 4475 3528 4476
rect 3522 4474 3528 4475
rect 2834 4470 2840 4471
rect 2390 4443 2397 4444
rect 2390 4439 2391 4443
rect 2396 4439 2397 4443
rect 2390 4438 2397 4439
rect 2494 4443 2500 4444
rect 2494 4439 2495 4443
rect 2499 4442 2500 4443
rect 2639 4443 2645 4444
rect 2639 4442 2640 4443
rect 2499 4440 2640 4442
rect 2499 4439 2500 4440
rect 2494 4438 2500 4439
rect 2639 4439 2640 4440
rect 2644 4439 2645 4443
rect 2639 4438 2645 4439
rect 2871 4443 2880 4444
rect 2871 4439 2872 4443
rect 2879 4439 2880 4443
rect 2871 4438 2880 4439
rect 3095 4443 3104 4444
rect 3095 4439 3096 4443
rect 3103 4439 3104 4443
rect 3095 4438 3104 4439
rect 3311 4443 3320 4444
rect 3311 4439 3312 4443
rect 3319 4439 3320 4443
rect 3311 4438 3320 4439
rect 3519 4443 3528 4444
rect 3519 4439 3520 4443
rect 3527 4439 3528 4443
rect 3519 4438 3528 4439
rect 3734 4443 3741 4444
rect 3734 4439 3735 4443
rect 3740 4439 3741 4443
rect 3734 4438 3741 4439
rect 4479 4439 4485 4440
rect 4479 4438 4480 4439
rect 1974 4436 1980 4437
rect 3798 4436 3804 4437
rect 4437 4436 4480 4438
rect 110 4433 116 4434
rect 1934 4433 1940 4434
rect 110 4429 111 4433
rect 115 4429 116 4433
rect 110 4428 116 4429
rect 510 4432 516 4433
rect 510 4428 511 4432
rect 515 4428 516 4432
rect 510 4427 516 4428
rect 686 4432 692 4433
rect 686 4428 687 4432
rect 691 4428 692 4432
rect 686 4427 692 4428
rect 870 4432 876 4433
rect 870 4428 871 4432
rect 875 4428 876 4432
rect 870 4427 876 4428
rect 1070 4432 1076 4433
rect 1070 4428 1071 4432
rect 1075 4428 1076 4432
rect 1070 4427 1076 4428
rect 1278 4432 1284 4433
rect 1278 4428 1279 4432
rect 1283 4428 1284 4432
rect 1278 4427 1284 4428
rect 1494 4432 1500 4433
rect 1494 4428 1495 4432
rect 1499 4428 1500 4432
rect 1494 4427 1500 4428
rect 1718 4432 1724 4433
rect 1718 4428 1719 4432
rect 1723 4428 1724 4432
rect 1934 4429 1935 4433
rect 1939 4429 1940 4433
rect 1974 4432 1975 4436
rect 1979 4432 1980 4436
rect 1974 4431 1980 4432
rect 2266 4435 2272 4436
rect 2266 4431 2267 4435
rect 2271 4431 2272 4435
rect 2266 4430 2272 4431
rect 2514 4435 2520 4436
rect 2514 4431 2515 4435
rect 2519 4431 2520 4435
rect 2514 4430 2520 4431
rect 2746 4435 2752 4436
rect 2746 4431 2747 4435
rect 2751 4431 2752 4435
rect 2746 4430 2752 4431
rect 2970 4435 2976 4436
rect 2970 4431 2971 4435
rect 2975 4431 2976 4435
rect 2970 4430 2976 4431
rect 3186 4435 3192 4436
rect 3186 4431 3187 4435
rect 3191 4431 3192 4435
rect 3186 4430 3192 4431
rect 3394 4435 3400 4436
rect 3394 4431 3395 4435
rect 3399 4431 3400 4435
rect 3394 4430 3400 4431
rect 3610 4435 3616 4436
rect 3610 4431 3611 4435
rect 3615 4431 3616 4435
rect 3798 4432 3799 4436
rect 3803 4432 3804 4436
rect 4479 4435 4480 4436
rect 4484 4435 4485 4439
rect 4615 4439 4621 4440
rect 4615 4438 4616 4439
rect 4573 4436 4616 4438
rect 4479 4434 4485 4435
rect 4615 4435 4616 4436
rect 4620 4435 4621 4439
rect 4751 4439 4757 4440
rect 4751 4438 4752 4439
rect 4709 4436 4752 4438
rect 4615 4434 4621 4435
rect 4751 4435 4752 4436
rect 4756 4435 4757 4439
rect 4887 4439 4893 4440
rect 4887 4438 4888 4439
rect 4845 4436 4888 4438
rect 4751 4434 4757 4435
rect 4887 4435 4888 4436
rect 4892 4435 4893 4439
rect 5074 4439 5080 4440
rect 5074 4438 5075 4439
rect 4981 4436 5075 4438
rect 4887 4434 4893 4435
rect 5074 4435 5075 4436
rect 5079 4435 5080 4439
rect 5074 4434 5080 4435
rect 3798 4431 3804 4432
rect 3610 4430 3616 4431
rect 1934 4428 1940 4429
rect 1718 4427 1724 4428
rect 2294 4420 2300 4421
rect 1974 4419 1980 4420
rect 482 4417 488 4418
rect 110 4416 116 4417
rect 110 4412 111 4416
rect 115 4412 116 4416
rect 482 4413 483 4417
rect 487 4413 488 4417
rect 482 4412 488 4413
rect 658 4417 664 4418
rect 658 4413 659 4417
rect 663 4413 664 4417
rect 658 4412 664 4413
rect 842 4417 848 4418
rect 842 4413 843 4417
rect 847 4413 848 4417
rect 842 4412 848 4413
rect 1042 4417 1048 4418
rect 1042 4413 1043 4417
rect 1047 4413 1048 4417
rect 1042 4412 1048 4413
rect 1250 4417 1256 4418
rect 1250 4413 1251 4417
rect 1255 4413 1256 4417
rect 1250 4412 1256 4413
rect 1466 4417 1472 4418
rect 1466 4413 1467 4417
rect 1471 4413 1472 4417
rect 1466 4412 1472 4413
rect 1690 4417 1696 4418
rect 1690 4413 1691 4417
rect 1695 4413 1696 4417
rect 1690 4412 1696 4413
rect 1934 4416 1940 4417
rect 1934 4412 1935 4416
rect 1939 4412 1940 4416
rect 1974 4415 1975 4419
rect 1979 4415 1980 4419
rect 2294 4416 2295 4420
rect 2299 4416 2300 4420
rect 2294 4415 2300 4416
rect 2542 4420 2548 4421
rect 2542 4416 2543 4420
rect 2547 4416 2548 4420
rect 2542 4415 2548 4416
rect 2774 4420 2780 4421
rect 2774 4416 2775 4420
rect 2779 4416 2780 4420
rect 2774 4415 2780 4416
rect 2998 4420 3004 4421
rect 2998 4416 2999 4420
rect 3003 4416 3004 4420
rect 2998 4415 3004 4416
rect 3214 4420 3220 4421
rect 3214 4416 3215 4420
rect 3219 4416 3220 4420
rect 3214 4415 3220 4416
rect 3422 4420 3428 4421
rect 3422 4416 3423 4420
rect 3427 4416 3428 4420
rect 3422 4415 3428 4416
rect 3638 4420 3644 4421
rect 3638 4416 3639 4420
rect 3643 4416 3644 4420
rect 3638 4415 3644 4416
rect 3798 4419 3804 4420
rect 3798 4415 3799 4419
rect 3803 4415 3804 4419
rect 1974 4414 1980 4415
rect 3798 4414 3804 4415
rect 110 4411 116 4412
rect 1934 4411 1940 4412
rect 607 4407 613 4408
rect 607 4403 608 4407
rect 612 4406 613 4407
rect 674 4407 680 4408
rect 674 4406 675 4407
rect 612 4404 675 4406
rect 612 4403 613 4404
rect 607 4402 613 4403
rect 674 4403 675 4404
rect 679 4403 680 4407
rect 674 4402 680 4403
rect 783 4407 789 4408
rect 783 4403 784 4407
rect 788 4406 789 4407
rect 858 4407 864 4408
rect 858 4406 859 4407
rect 788 4404 859 4406
rect 788 4403 789 4404
rect 783 4402 789 4403
rect 858 4403 859 4404
rect 863 4403 864 4407
rect 858 4402 864 4403
rect 967 4407 973 4408
rect 967 4403 968 4407
rect 972 4406 973 4407
rect 1058 4407 1064 4408
rect 1058 4406 1059 4407
rect 972 4404 1059 4406
rect 972 4403 973 4404
rect 967 4402 973 4403
rect 1058 4403 1059 4404
rect 1063 4403 1064 4407
rect 1058 4402 1064 4403
rect 1167 4407 1173 4408
rect 1167 4403 1168 4407
rect 1172 4406 1173 4407
rect 1266 4407 1272 4408
rect 1266 4406 1267 4407
rect 1172 4404 1267 4406
rect 1172 4403 1173 4404
rect 1167 4402 1173 4403
rect 1266 4403 1267 4404
rect 1271 4403 1272 4407
rect 1266 4402 1272 4403
rect 1362 4407 1368 4408
rect 1362 4403 1363 4407
rect 1367 4406 1368 4407
rect 1375 4407 1381 4408
rect 1375 4406 1376 4407
rect 1367 4404 1376 4406
rect 1367 4403 1368 4404
rect 1362 4402 1368 4403
rect 1375 4403 1376 4404
rect 1380 4403 1381 4407
rect 1375 4402 1381 4403
rect 1562 4407 1568 4408
rect 1562 4403 1563 4407
rect 1567 4406 1568 4407
rect 1591 4407 1597 4408
rect 1591 4406 1592 4407
rect 1567 4404 1592 4406
rect 1567 4403 1568 4404
rect 1562 4402 1568 4403
rect 1591 4403 1592 4404
rect 1596 4403 1597 4407
rect 1591 4402 1597 4403
rect 1610 4407 1616 4408
rect 1610 4403 1611 4407
rect 1615 4406 1616 4407
rect 1815 4407 1821 4408
rect 1815 4406 1816 4407
rect 1615 4404 1816 4406
rect 1615 4403 1616 4404
rect 1610 4402 1616 4403
rect 1815 4403 1816 4404
rect 1820 4403 1821 4407
rect 1815 4402 1821 4403
rect 4466 4403 4477 4404
rect 4466 4399 4467 4403
rect 4471 4399 4472 4403
rect 4476 4399 4477 4403
rect 4466 4398 4477 4399
rect 4479 4403 4485 4404
rect 4479 4399 4480 4403
rect 4484 4402 4485 4403
rect 4607 4403 4613 4404
rect 4607 4402 4608 4403
rect 4484 4400 4608 4402
rect 4484 4399 4485 4400
rect 4479 4398 4485 4399
rect 4607 4399 4608 4400
rect 4612 4399 4613 4403
rect 4607 4398 4613 4399
rect 4615 4403 4621 4404
rect 4615 4399 4616 4403
rect 4620 4402 4621 4403
rect 4743 4403 4749 4404
rect 4743 4402 4744 4403
rect 4620 4400 4744 4402
rect 4620 4399 4621 4400
rect 4615 4398 4621 4399
rect 4743 4399 4744 4400
rect 4748 4399 4749 4403
rect 4743 4398 4749 4399
rect 4751 4403 4757 4404
rect 4751 4399 4752 4403
rect 4756 4402 4757 4403
rect 4879 4403 4885 4404
rect 4879 4402 4880 4403
rect 4756 4400 4880 4402
rect 4756 4399 4757 4400
rect 4751 4398 4757 4399
rect 4879 4399 4880 4400
rect 4884 4399 4885 4403
rect 4879 4398 4885 4399
rect 4887 4403 4893 4404
rect 4887 4399 4888 4403
rect 4892 4402 4893 4403
rect 5015 4403 5021 4404
rect 5015 4402 5016 4403
rect 4892 4400 5016 4402
rect 4892 4399 4893 4400
rect 4887 4398 4893 4399
rect 5015 4399 5016 4400
rect 5020 4399 5021 4403
rect 5015 4398 5021 4399
rect 3838 4396 3844 4397
rect 5662 4396 5668 4397
rect 3838 4392 3839 4396
rect 3843 4392 3844 4396
rect 3838 4391 3844 4392
rect 4346 4395 4352 4396
rect 4346 4391 4347 4395
rect 4351 4391 4352 4395
rect 4346 4390 4352 4391
rect 4482 4395 4488 4396
rect 4482 4391 4483 4395
rect 4487 4391 4488 4395
rect 4482 4390 4488 4391
rect 4618 4395 4624 4396
rect 4618 4391 4619 4395
rect 4623 4391 4624 4395
rect 4618 4390 4624 4391
rect 4754 4395 4760 4396
rect 4754 4391 4755 4395
rect 4759 4391 4760 4395
rect 4754 4390 4760 4391
rect 4890 4395 4896 4396
rect 4890 4391 4891 4395
rect 4895 4391 4896 4395
rect 5662 4392 5663 4396
rect 5667 4392 5668 4396
rect 5662 4391 5668 4392
rect 4890 4390 4896 4391
rect 4374 4380 4380 4381
rect 3838 4379 3844 4380
rect 578 4375 584 4376
rect 578 4374 579 4375
rect 573 4372 579 4374
rect 578 4371 579 4372
rect 583 4371 584 4375
rect 578 4370 584 4371
rect 674 4375 680 4376
rect 674 4371 675 4375
rect 679 4371 680 4375
rect 674 4370 680 4371
rect 858 4375 864 4376
rect 858 4371 859 4375
rect 863 4371 864 4375
rect 858 4370 864 4371
rect 1058 4375 1064 4376
rect 1058 4371 1059 4375
rect 1063 4371 1064 4375
rect 1058 4370 1064 4371
rect 1266 4375 1272 4376
rect 1266 4371 1267 4375
rect 1271 4371 1272 4375
rect 1610 4375 1616 4376
rect 1610 4374 1611 4375
rect 1557 4372 1611 4374
rect 1266 4370 1272 4371
rect 1610 4371 1611 4372
rect 1615 4371 1616 4375
rect 1610 4370 1616 4371
rect 1778 4375 1784 4376
rect 1778 4371 1779 4375
rect 1783 4371 1784 4375
rect 3838 4375 3839 4379
rect 3843 4375 3844 4379
rect 4374 4376 4375 4380
rect 4379 4376 4380 4380
rect 4374 4375 4380 4376
rect 4510 4380 4516 4381
rect 4510 4376 4511 4380
rect 4515 4376 4516 4380
rect 4510 4375 4516 4376
rect 4646 4380 4652 4381
rect 4646 4376 4647 4380
rect 4651 4376 4652 4380
rect 4646 4375 4652 4376
rect 4782 4380 4788 4381
rect 4782 4376 4783 4380
rect 4787 4376 4788 4380
rect 4782 4375 4788 4376
rect 4918 4380 4924 4381
rect 4918 4376 4919 4380
rect 4923 4376 4924 4380
rect 4918 4375 4924 4376
rect 5662 4379 5668 4380
rect 5662 4375 5663 4379
rect 5667 4375 5668 4379
rect 3838 4374 3844 4375
rect 5662 4374 5668 4375
rect 1778 4370 1784 4371
rect 1974 4349 1980 4350
rect 3798 4349 3804 4350
rect 1974 4345 1975 4349
rect 1979 4345 1980 4349
rect 1974 4344 1980 4345
rect 2022 4348 2028 4349
rect 2022 4344 2023 4348
rect 2027 4344 2028 4348
rect 2022 4343 2028 4344
rect 2198 4348 2204 4349
rect 2198 4344 2199 4348
rect 2203 4344 2204 4348
rect 2198 4343 2204 4344
rect 2398 4348 2404 4349
rect 2398 4344 2399 4348
rect 2403 4344 2404 4348
rect 2398 4343 2404 4344
rect 2590 4348 2596 4349
rect 2590 4344 2591 4348
rect 2595 4344 2596 4348
rect 2590 4343 2596 4344
rect 2774 4348 2780 4349
rect 2774 4344 2775 4348
rect 2779 4344 2780 4348
rect 2774 4343 2780 4344
rect 2950 4348 2956 4349
rect 2950 4344 2951 4348
rect 2955 4344 2956 4348
rect 2950 4343 2956 4344
rect 3134 4348 3140 4349
rect 3134 4344 3135 4348
rect 3139 4344 3140 4348
rect 3134 4343 3140 4344
rect 3318 4348 3324 4349
rect 3318 4344 3319 4348
rect 3323 4344 3324 4348
rect 3798 4345 3799 4349
rect 3803 4345 3804 4349
rect 3798 4344 3804 4345
rect 3318 4343 3324 4344
rect 1362 4335 1368 4336
rect 1362 4334 1363 4335
rect 840 4332 1363 4334
rect 840 4322 842 4332
rect 1362 4331 1363 4332
rect 1367 4331 1368 4335
rect 1994 4333 2000 4334
rect 1362 4330 1368 4331
rect 1974 4332 1980 4333
rect 1974 4328 1975 4332
rect 1979 4328 1980 4332
rect 1994 4329 1995 4333
rect 1999 4329 2000 4333
rect 1994 4328 2000 4329
rect 2170 4333 2176 4334
rect 2170 4329 2171 4333
rect 2175 4329 2176 4333
rect 2170 4328 2176 4329
rect 2370 4333 2376 4334
rect 2370 4329 2371 4333
rect 2375 4329 2376 4333
rect 2370 4328 2376 4329
rect 2562 4333 2568 4334
rect 2562 4329 2563 4333
rect 2567 4329 2568 4333
rect 2562 4328 2568 4329
rect 2746 4333 2752 4334
rect 2746 4329 2747 4333
rect 2751 4329 2752 4333
rect 2746 4328 2752 4329
rect 2922 4333 2928 4334
rect 2922 4329 2923 4333
rect 2927 4329 2928 4333
rect 2922 4328 2928 4329
rect 3106 4333 3112 4334
rect 3106 4329 3107 4333
rect 3111 4329 3112 4333
rect 3106 4328 3112 4329
rect 3290 4333 3296 4334
rect 3290 4329 3291 4333
rect 3295 4329 3296 4333
rect 3290 4328 3296 4329
rect 3798 4332 3804 4333
rect 3798 4328 3799 4332
rect 3803 4328 3804 4332
rect 1974 4327 1980 4328
rect 3798 4327 3804 4328
rect 805 4320 842 4322
rect 847 4323 853 4324
rect 847 4319 848 4323
rect 852 4322 853 4323
rect 983 4323 989 4324
rect 852 4320 869 4322
rect 852 4319 853 4320
rect 847 4318 853 4319
rect 983 4319 984 4323
rect 988 4322 989 4323
rect 1119 4323 1125 4324
rect 988 4320 1005 4322
rect 988 4319 989 4320
rect 983 4318 989 4319
rect 1119 4319 1120 4323
rect 1124 4322 1125 4323
rect 1255 4323 1261 4324
rect 1124 4320 1141 4322
rect 1124 4319 1125 4320
rect 1119 4318 1125 4319
rect 1255 4319 1256 4323
rect 1260 4322 1261 4323
rect 1522 4323 1528 4324
rect 1260 4320 1277 4322
rect 1260 4319 1261 4320
rect 1255 4318 1261 4319
rect 1522 4319 1523 4323
rect 1527 4322 1528 4323
rect 1658 4323 1664 4324
rect 1527 4320 1549 4322
rect 1527 4319 1528 4320
rect 1522 4318 1528 4319
rect 1658 4319 1659 4323
rect 1663 4322 1664 4323
rect 2098 4323 2104 4324
rect 1663 4320 1685 4322
rect 1663 4319 1664 4320
rect 1658 4318 1664 4319
rect 2098 4319 2099 4323
rect 2103 4322 2104 4323
rect 2119 4323 2125 4324
rect 2119 4322 2120 4323
rect 2103 4320 2120 4322
rect 2103 4319 2104 4320
rect 2098 4318 2104 4319
rect 2119 4319 2120 4320
rect 2124 4319 2125 4323
rect 2119 4318 2125 4319
rect 2151 4323 2157 4324
rect 2151 4319 2152 4323
rect 2156 4322 2157 4323
rect 2295 4323 2301 4324
rect 2295 4322 2296 4323
rect 2156 4320 2296 4322
rect 2156 4319 2157 4320
rect 2151 4318 2157 4319
rect 2295 4319 2296 4320
rect 2300 4319 2301 4323
rect 2295 4318 2301 4319
rect 2310 4323 2316 4324
rect 2310 4319 2311 4323
rect 2315 4322 2316 4323
rect 2495 4323 2501 4324
rect 2495 4322 2496 4323
rect 2315 4320 2496 4322
rect 2315 4319 2316 4320
rect 2310 4318 2316 4319
rect 2495 4319 2496 4320
rect 2500 4319 2501 4323
rect 2495 4318 2501 4319
rect 2687 4323 2693 4324
rect 2687 4319 2688 4323
rect 2692 4322 2693 4323
rect 2762 4323 2768 4324
rect 2762 4322 2763 4323
rect 2692 4320 2763 4322
rect 2692 4319 2693 4320
rect 2687 4318 2693 4319
rect 2762 4319 2763 4320
rect 2767 4319 2768 4323
rect 2762 4318 2768 4319
rect 2871 4323 2877 4324
rect 2871 4319 2872 4323
rect 2876 4322 2877 4323
rect 2938 4323 2944 4324
rect 2938 4322 2939 4323
rect 2876 4320 2939 4322
rect 2876 4319 2877 4320
rect 2871 4318 2877 4319
rect 2938 4319 2939 4320
rect 2943 4319 2944 4323
rect 2938 4318 2944 4319
rect 3047 4323 3053 4324
rect 3047 4319 3048 4323
rect 3052 4322 3053 4323
rect 3122 4323 3128 4324
rect 3122 4322 3123 4323
rect 3052 4320 3123 4322
rect 3052 4319 3053 4320
rect 3047 4318 3053 4319
rect 3122 4319 3123 4320
rect 3127 4319 3128 4323
rect 3122 4318 3128 4319
rect 3231 4323 3237 4324
rect 3231 4319 3232 4323
rect 3236 4322 3237 4323
rect 3306 4323 3312 4324
rect 3306 4322 3307 4323
rect 3236 4320 3307 4322
rect 3236 4319 3237 4320
rect 3231 4318 3237 4319
rect 3306 4319 3307 4320
rect 3311 4319 3312 4323
rect 3415 4323 3421 4324
rect 3415 4322 3416 4323
rect 3306 4318 3312 4319
rect 3316 4320 3416 4322
rect 1480 4306 1482 4317
rect 2834 4315 2840 4316
rect 2834 4311 2835 4315
rect 2839 4314 2840 4315
rect 3316 4314 3318 4320
rect 3415 4319 3416 4320
rect 3420 4319 3421 4323
rect 3415 4318 3421 4319
rect 2839 4312 3318 4314
rect 2839 4311 2840 4312
rect 2834 4310 2840 4311
rect 1618 4307 1624 4308
rect 1618 4306 1619 4307
rect 1480 4304 1619 4306
rect 1618 4303 1619 4304
rect 1623 4303 1624 4307
rect 1618 4302 1624 4303
rect 3838 4305 3844 4306
rect 5662 4305 5668 4306
rect 3838 4301 3839 4305
rect 3843 4301 3844 4305
rect 3838 4300 3844 4301
rect 4134 4304 4140 4305
rect 4134 4300 4135 4304
rect 4139 4300 4140 4304
rect 4134 4299 4140 4300
rect 4270 4304 4276 4305
rect 4270 4300 4271 4304
rect 4275 4300 4276 4304
rect 4270 4299 4276 4300
rect 4406 4304 4412 4305
rect 4406 4300 4407 4304
rect 4411 4300 4412 4304
rect 4406 4299 4412 4300
rect 4542 4304 4548 4305
rect 4542 4300 4543 4304
rect 4547 4300 4548 4304
rect 4542 4299 4548 4300
rect 4678 4304 4684 4305
rect 4678 4300 4679 4304
rect 4683 4300 4684 4304
rect 5662 4301 5663 4305
rect 5667 4301 5668 4305
rect 5662 4300 5668 4301
rect 4678 4299 4684 4300
rect 2151 4291 2157 4292
rect 2151 4290 2152 4291
rect 2085 4288 2152 4290
rect 839 4287 845 4288
rect 839 4283 840 4287
rect 844 4286 845 4287
rect 847 4287 853 4288
rect 847 4286 848 4287
rect 844 4284 848 4286
rect 844 4283 845 4284
rect 839 4282 845 4283
rect 847 4283 848 4284
rect 852 4283 853 4287
rect 847 4282 853 4283
rect 975 4287 981 4288
rect 975 4283 976 4287
rect 980 4286 981 4287
rect 983 4287 989 4288
rect 983 4286 984 4287
rect 980 4284 984 4286
rect 980 4283 981 4284
rect 975 4282 981 4283
rect 983 4283 984 4284
rect 988 4283 989 4287
rect 983 4282 989 4283
rect 1111 4287 1117 4288
rect 1111 4283 1112 4287
rect 1116 4286 1117 4287
rect 1119 4287 1125 4288
rect 1119 4286 1120 4287
rect 1116 4284 1120 4286
rect 1116 4283 1117 4284
rect 1111 4282 1117 4283
rect 1119 4283 1120 4284
rect 1124 4283 1125 4287
rect 1119 4282 1125 4283
rect 1247 4287 1253 4288
rect 1247 4283 1248 4287
rect 1252 4286 1253 4287
rect 1255 4287 1261 4288
rect 1255 4286 1256 4287
rect 1252 4284 1256 4286
rect 1252 4283 1253 4284
rect 1247 4282 1253 4283
rect 1255 4283 1256 4284
rect 1260 4283 1261 4287
rect 1255 4282 1261 4283
rect 1330 4287 1336 4288
rect 1330 4283 1331 4287
rect 1335 4286 1336 4287
rect 1383 4287 1389 4288
rect 1383 4286 1384 4287
rect 1335 4284 1384 4286
rect 1335 4283 1336 4284
rect 1330 4282 1336 4283
rect 1383 4283 1384 4284
rect 1388 4283 1389 4287
rect 1383 4282 1389 4283
rect 1519 4287 1528 4288
rect 1519 4283 1520 4287
rect 1527 4283 1528 4287
rect 1519 4282 1528 4283
rect 1655 4287 1664 4288
rect 1655 4283 1656 4287
rect 1663 4283 1664 4287
rect 1655 4282 1664 4283
rect 1778 4287 1784 4288
rect 1778 4283 1779 4287
rect 1783 4286 1784 4287
rect 1791 4287 1797 4288
rect 1791 4286 1792 4287
rect 1783 4284 1792 4286
rect 1783 4283 1784 4284
rect 1778 4282 1784 4283
rect 1791 4283 1792 4284
rect 1796 4283 1797 4287
rect 2151 4287 2152 4288
rect 2156 4287 2157 4291
rect 2310 4291 2316 4292
rect 2310 4290 2311 4291
rect 2261 4288 2311 4290
rect 2151 4286 2157 4287
rect 2310 4287 2311 4288
rect 2315 4287 2316 4291
rect 2310 4286 2316 4287
rect 2390 4291 2396 4292
rect 2390 4287 2391 4291
rect 2395 4287 2396 4291
rect 2390 4286 2396 4287
rect 2630 4291 2636 4292
rect 2630 4287 2631 4291
rect 2635 4287 2636 4291
rect 2630 4286 2636 4287
rect 2762 4291 2768 4292
rect 2762 4287 2763 4291
rect 2767 4287 2768 4291
rect 2762 4286 2768 4287
rect 2938 4291 2944 4292
rect 2938 4287 2939 4291
rect 2943 4287 2944 4291
rect 2938 4286 2944 4287
rect 3122 4291 3128 4292
rect 3122 4287 3123 4291
rect 3127 4287 3128 4291
rect 3122 4286 3128 4287
rect 3306 4291 3312 4292
rect 3306 4287 3307 4291
rect 3311 4287 3312 4291
rect 4106 4289 4112 4290
rect 3306 4286 3312 4287
rect 3838 4288 3844 4289
rect 3838 4284 3839 4288
rect 3843 4284 3844 4288
rect 4106 4285 4107 4289
rect 4111 4285 4112 4289
rect 4106 4284 4112 4285
rect 4242 4289 4248 4290
rect 4242 4285 4243 4289
rect 4247 4285 4248 4289
rect 4242 4284 4248 4285
rect 4378 4289 4384 4290
rect 4378 4285 4379 4289
rect 4383 4285 4384 4289
rect 4378 4284 4384 4285
rect 4514 4289 4520 4290
rect 4514 4285 4515 4289
rect 4519 4285 4520 4289
rect 4514 4284 4520 4285
rect 4650 4289 4656 4290
rect 4650 4285 4651 4289
rect 4655 4285 4656 4289
rect 4650 4284 4656 4285
rect 5662 4288 5668 4289
rect 5662 4284 5663 4288
rect 5667 4284 5668 4288
rect 3838 4283 3844 4284
rect 5662 4283 5668 4284
rect 1791 4282 1797 4283
rect 110 4280 116 4281
rect 1934 4280 1940 4281
rect 110 4276 111 4280
rect 115 4276 116 4280
rect 110 4275 116 4276
rect 714 4279 720 4280
rect 714 4275 715 4279
rect 719 4275 720 4279
rect 714 4274 720 4275
rect 850 4279 856 4280
rect 850 4275 851 4279
rect 855 4275 856 4279
rect 850 4274 856 4275
rect 986 4279 992 4280
rect 986 4275 987 4279
rect 991 4275 992 4279
rect 986 4274 992 4275
rect 1122 4279 1128 4280
rect 1122 4275 1123 4279
rect 1127 4275 1128 4279
rect 1122 4274 1128 4275
rect 1258 4279 1264 4280
rect 1258 4275 1259 4279
rect 1263 4275 1264 4279
rect 1258 4274 1264 4275
rect 1394 4279 1400 4280
rect 1394 4275 1395 4279
rect 1399 4275 1400 4279
rect 1394 4274 1400 4275
rect 1530 4279 1536 4280
rect 1530 4275 1531 4279
rect 1535 4275 1536 4279
rect 1530 4274 1536 4275
rect 1666 4279 1672 4280
rect 1666 4275 1667 4279
rect 1671 4275 1672 4279
rect 1934 4276 1935 4280
rect 1939 4276 1940 4280
rect 1934 4275 1940 4276
rect 4231 4279 4240 4280
rect 4231 4275 4232 4279
rect 4239 4275 4240 4279
rect 1666 4274 1672 4275
rect 4231 4274 4240 4275
rect 4250 4279 4256 4280
rect 4250 4275 4251 4279
rect 4255 4278 4256 4279
rect 4367 4279 4373 4280
rect 4367 4278 4368 4279
rect 4255 4276 4368 4278
rect 4255 4275 4256 4276
rect 4250 4274 4256 4275
rect 4367 4275 4368 4276
rect 4372 4275 4373 4279
rect 4367 4274 4373 4275
rect 4503 4279 4509 4280
rect 4503 4275 4504 4279
rect 4508 4278 4509 4279
rect 4530 4279 4536 4280
rect 4530 4278 4531 4279
rect 4508 4276 4531 4278
rect 4508 4275 4509 4276
rect 4503 4274 4509 4275
rect 4530 4275 4531 4276
rect 4535 4275 4536 4279
rect 4530 4274 4536 4275
rect 4639 4279 4645 4280
rect 4639 4275 4640 4279
rect 4644 4278 4645 4279
rect 4666 4279 4672 4280
rect 4666 4278 4667 4279
rect 4644 4276 4667 4278
rect 4644 4275 4645 4276
rect 4639 4274 4645 4275
rect 4666 4275 4667 4276
rect 4671 4275 4672 4279
rect 4775 4279 4781 4280
rect 4775 4278 4776 4279
rect 4666 4274 4672 4275
rect 4676 4276 4776 4278
rect 4330 4271 4336 4272
rect 4330 4267 4331 4271
rect 4335 4270 4336 4271
rect 4676 4270 4678 4276
rect 4775 4275 4776 4276
rect 4780 4275 4781 4279
rect 4775 4274 4781 4275
rect 4335 4268 4678 4270
rect 4335 4267 4336 4268
rect 4330 4266 4336 4267
rect 742 4264 748 4265
rect 110 4263 116 4264
rect 110 4259 111 4263
rect 115 4259 116 4263
rect 742 4260 743 4264
rect 747 4260 748 4264
rect 742 4259 748 4260
rect 878 4264 884 4265
rect 878 4260 879 4264
rect 883 4260 884 4264
rect 878 4259 884 4260
rect 1014 4264 1020 4265
rect 1014 4260 1015 4264
rect 1019 4260 1020 4264
rect 1014 4259 1020 4260
rect 1150 4264 1156 4265
rect 1150 4260 1151 4264
rect 1155 4260 1156 4264
rect 1150 4259 1156 4260
rect 1286 4264 1292 4265
rect 1286 4260 1287 4264
rect 1291 4260 1292 4264
rect 1286 4259 1292 4260
rect 1422 4264 1428 4265
rect 1422 4260 1423 4264
rect 1427 4260 1428 4264
rect 1422 4259 1428 4260
rect 1558 4264 1564 4265
rect 1558 4260 1559 4264
rect 1563 4260 1564 4264
rect 1558 4259 1564 4260
rect 1694 4264 1700 4265
rect 1694 4260 1695 4264
rect 1699 4260 1700 4264
rect 1694 4259 1700 4260
rect 1934 4263 1940 4264
rect 1934 4259 1935 4263
rect 1939 4259 1940 4263
rect 110 4258 116 4259
rect 1934 4258 1940 4259
rect 4250 4247 4256 4248
rect 4250 4246 4251 4247
rect 4197 4244 4251 4246
rect 4250 4243 4251 4244
rect 4255 4243 4256 4247
rect 4250 4242 4256 4243
rect 4330 4247 4336 4248
rect 4330 4243 4331 4247
rect 4335 4243 4336 4247
rect 4330 4242 4336 4243
rect 4466 4247 4472 4248
rect 4466 4243 4467 4247
rect 4471 4243 4472 4247
rect 4466 4242 4472 4243
rect 4530 4247 4536 4248
rect 4530 4243 4531 4247
rect 4535 4243 4536 4247
rect 4530 4242 4536 4243
rect 4666 4247 4672 4248
rect 4666 4243 4667 4247
rect 4671 4243 4672 4247
rect 4666 4242 4672 4243
rect 2098 4239 2104 4240
rect 2098 4238 2099 4239
rect 2085 4236 2099 4238
rect 2098 4235 2099 4236
rect 2103 4235 2104 4239
rect 2375 4239 2381 4240
rect 2098 4234 2104 4235
rect 2330 4235 2336 4236
rect 2330 4231 2331 4235
rect 2335 4231 2336 4235
rect 2375 4235 2376 4239
rect 2380 4238 2381 4239
rect 2958 4239 2964 4240
rect 2958 4238 2959 4239
rect 2380 4236 2525 4238
rect 2853 4236 2959 4238
rect 2380 4235 2381 4236
rect 2375 4234 2381 4235
rect 2958 4235 2959 4236
rect 2963 4235 2964 4239
rect 3279 4239 3285 4240
rect 3279 4238 3280 4239
rect 3109 4236 3280 4238
rect 2958 4234 2964 4235
rect 3279 4235 3280 4236
rect 3284 4235 3285 4239
rect 3279 4234 3285 4235
rect 3370 4235 3376 4236
rect 2330 4230 2336 4231
rect 3370 4231 3371 4235
rect 3375 4231 3376 4235
rect 3370 4230 3376 4231
rect 2330 4211 2336 4212
rect 2330 4207 2331 4211
rect 2335 4210 2336 4211
rect 2335 4208 2642 4210
rect 2335 4207 2336 4208
rect 2330 4206 2336 4207
rect 1946 4203 1952 4204
rect 1946 4199 1947 4203
rect 1951 4202 1952 4203
rect 2119 4203 2125 4204
rect 2119 4202 2120 4203
rect 1951 4200 2120 4202
rect 1951 4199 1952 4200
rect 1946 4198 1952 4199
rect 2119 4199 2120 4200
rect 2124 4199 2125 4203
rect 2119 4198 2125 4199
rect 2367 4203 2373 4204
rect 2367 4199 2368 4203
rect 2372 4202 2373 4203
rect 2375 4203 2381 4204
rect 2375 4202 2376 4203
rect 2372 4200 2376 4202
rect 2372 4199 2373 4200
rect 2367 4198 2373 4199
rect 2375 4199 2376 4200
rect 2380 4199 2381 4203
rect 2375 4198 2381 4199
rect 2630 4203 2637 4204
rect 2630 4199 2631 4203
rect 2636 4199 2637 4203
rect 2640 4202 2642 4208
rect 2887 4203 2893 4204
rect 2887 4202 2888 4203
rect 2640 4200 2888 4202
rect 2630 4198 2637 4199
rect 2887 4199 2888 4200
rect 2892 4199 2893 4203
rect 2887 4198 2893 4199
rect 2958 4203 2964 4204
rect 2958 4199 2959 4203
rect 2963 4202 2964 4203
rect 3143 4203 3149 4204
rect 3143 4202 3144 4203
rect 2963 4200 3144 4202
rect 2963 4199 2964 4200
rect 2958 4198 2964 4199
rect 3143 4199 3144 4200
rect 3148 4199 3149 4203
rect 3143 4198 3149 4199
rect 3279 4203 3285 4204
rect 3279 4199 3280 4203
rect 3284 4202 3285 4203
rect 3407 4203 3413 4204
rect 3407 4202 3408 4203
rect 3284 4200 3408 4202
rect 3284 4199 3285 4200
rect 3279 4198 3285 4199
rect 3407 4199 3408 4200
rect 3412 4199 3413 4203
rect 3407 4198 3413 4199
rect 110 4197 116 4198
rect 1934 4197 1940 4198
rect 110 4193 111 4197
rect 115 4193 116 4197
rect 110 4192 116 4193
rect 726 4196 732 4197
rect 726 4192 727 4196
rect 731 4192 732 4196
rect 726 4191 732 4192
rect 862 4196 868 4197
rect 862 4192 863 4196
rect 867 4192 868 4196
rect 862 4191 868 4192
rect 998 4196 1004 4197
rect 998 4192 999 4196
rect 1003 4192 1004 4196
rect 998 4191 1004 4192
rect 1134 4196 1140 4197
rect 1134 4192 1135 4196
rect 1139 4192 1140 4196
rect 1134 4191 1140 4192
rect 1270 4196 1276 4197
rect 1270 4192 1271 4196
rect 1275 4192 1276 4196
rect 1270 4191 1276 4192
rect 1406 4196 1412 4197
rect 1406 4192 1407 4196
rect 1411 4192 1412 4196
rect 1406 4191 1412 4192
rect 1542 4196 1548 4197
rect 1542 4192 1543 4196
rect 1547 4192 1548 4196
rect 1542 4191 1548 4192
rect 1678 4196 1684 4197
rect 1678 4192 1679 4196
rect 1683 4192 1684 4196
rect 1678 4191 1684 4192
rect 1814 4196 1820 4197
rect 1814 4192 1815 4196
rect 1819 4192 1820 4196
rect 1934 4193 1935 4197
rect 1939 4193 1940 4197
rect 1934 4192 1940 4193
rect 1974 4196 1980 4197
rect 3798 4196 3804 4197
rect 1974 4192 1975 4196
rect 1979 4192 1980 4196
rect 1814 4191 1820 4192
rect 1974 4191 1980 4192
rect 1994 4195 2000 4196
rect 1994 4191 1995 4195
rect 1999 4191 2000 4195
rect 1994 4190 2000 4191
rect 2242 4195 2248 4196
rect 2242 4191 2243 4195
rect 2247 4191 2248 4195
rect 2242 4190 2248 4191
rect 2506 4195 2512 4196
rect 2506 4191 2507 4195
rect 2511 4191 2512 4195
rect 2506 4190 2512 4191
rect 2762 4195 2768 4196
rect 2762 4191 2763 4195
rect 2767 4191 2768 4195
rect 2762 4190 2768 4191
rect 3018 4195 3024 4196
rect 3018 4191 3019 4195
rect 3023 4191 3024 4195
rect 3018 4190 3024 4191
rect 3282 4195 3288 4196
rect 3282 4191 3283 4195
rect 3287 4191 3288 4195
rect 3798 4192 3799 4196
rect 3803 4192 3804 4196
rect 3798 4191 3804 4192
rect 3282 4190 3288 4191
rect 4103 4187 4109 4188
rect 4058 4183 4064 4184
rect 698 4181 704 4182
rect 110 4180 116 4181
rect 110 4176 111 4180
rect 115 4176 116 4180
rect 698 4177 699 4181
rect 703 4177 704 4181
rect 698 4176 704 4177
rect 834 4181 840 4182
rect 834 4177 835 4181
rect 839 4177 840 4181
rect 834 4176 840 4177
rect 970 4181 976 4182
rect 970 4177 971 4181
rect 975 4177 976 4181
rect 970 4176 976 4177
rect 1106 4181 1112 4182
rect 1106 4177 1107 4181
rect 1111 4177 1112 4181
rect 1106 4176 1112 4177
rect 1242 4181 1248 4182
rect 1242 4177 1243 4181
rect 1247 4177 1248 4181
rect 1242 4176 1248 4177
rect 1378 4181 1384 4182
rect 1378 4177 1379 4181
rect 1383 4177 1384 4181
rect 1378 4176 1384 4177
rect 1514 4181 1520 4182
rect 1514 4177 1515 4181
rect 1519 4177 1520 4181
rect 1514 4176 1520 4177
rect 1650 4181 1656 4182
rect 1650 4177 1651 4181
rect 1655 4177 1656 4181
rect 1650 4176 1656 4177
rect 1786 4181 1792 4182
rect 1786 4177 1787 4181
rect 1791 4177 1792 4181
rect 1786 4176 1792 4177
rect 1934 4180 1940 4181
rect 2022 4180 2028 4181
rect 1934 4176 1935 4180
rect 1939 4176 1940 4180
rect 110 4175 116 4176
rect 1934 4175 1940 4176
rect 1974 4179 1980 4180
rect 1974 4175 1975 4179
rect 1979 4175 1980 4179
rect 2022 4176 2023 4180
rect 2027 4176 2028 4180
rect 2022 4175 2028 4176
rect 2270 4180 2276 4181
rect 2270 4176 2271 4180
rect 2275 4176 2276 4180
rect 2270 4175 2276 4176
rect 2534 4180 2540 4181
rect 2534 4176 2535 4180
rect 2539 4176 2540 4180
rect 2534 4175 2540 4176
rect 2790 4180 2796 4181
rect 2790 4176 2791 4180
rect 2795 4176 2796 4180
rect 2790 4175 2796 4176
rect 3046 4180 3052 4181
rect 3046 4176 3047 4180
rect 3051 4176 3052 4180
rect 3046 4175 3052 4176
rect 3310 4180 3316 4181
rect 3310 4176 3311 4180
rect 3315 4176 3316 4180
rect 3310 4175 3316 4176
rect 3798 4179 3804 4180
rect 3798 4175 3799 4179
rect 3803 4175 3804 4179
rect 4058 4179 4059 4183
rect 4063 4179 4064 4183
rect 4103 4183 4104 4187
rect 4108 4186 4109 4187
rect 4234 4187 4240 4188
rect 4108 4184 4125 4186
rect 4108 4183 4109 4184
rect 4103 4182 4109 4183
rect 4234 4183 4235 4187
rect 4239 4186 4240 4187
rect 4375 4187 4381 4188
rect 4239 4184 4261 4186
rect 4239 4183 4240 4184
rect 4234 4182 4240 4183
rect 4375 4183 4376 4187
rect 4380 4186 4381 4187
rect 4511 4187 4517 4188
rect 4380 4184 4397 4186
rect 4380 4183 4381 4184
rect 4375 4182 4381 4183
rect 4511 4183 4512 4187
rect 4516 4186 4517 4187
rect 4516 4184 4533 4186
rect 4516 4183 4517 4184
rect 4511 4182 4517 4183
rect 4058 4178 4064 4179
rect 1974 4174 1980 4175
rect 3798 4174 3804 4175
rect 823 4171 829 4172
rect 823 4167 824 4171
rect 828 4170 829 4171
rect 850 4171 856 4172
rect 850 4170 851 4171
rect 828 4168 851 4170
rect 828 4167 829 4168
rect 823 4166 829 4167
rect 850 4167 851 4168
rect 855 4167 856 4171
rect 850 4166 856 4167
rect 959 4171 968 4172
rect 959 4167 960 4171
rect 967 4167 968 4171
rect 1095 4171 1101 4172
rect 1095 4170 1096 4171
rect 959 4166 968 4167
rect 972 4168 1096 4170
rect 786 4163 792 4164
rect 786 4159 787 4163
rect 791 4162 792 4163
rect 972 4162 974 4168
rect 1095 4167 1096 4168
rect 1100 4167 1101 4171
rect 1095 4166 1101 4167
rect 1103 4171 1109 4172
rect 1103 4167 1104 4171
rect 1108 4170 1109 4171
rect 1231 4171 1237 4172
rect 1231 4170 1232 4171
rect 1108 4168 1232 4170
rect 1108 4167 1109 4168
rect 1103 4166 1109 4167
rect 1231 4167 1232 4168
rect 1236 4167 1237 4171
rect 1231 4166 1237 4167
rect 1239 4171 1245 4172
rect 1239 4167 1240 4171
rect 1244 4170 1245 4171
rect 1367 4171 1373 4172
rect 1367 4170 1368 4171
rect 1244 4168 1368 4170
rect 1244 4167 1245 4168
rect 1239 4166 1245 4167
rect 1367 4167 1368 4168
rect 1372 4167 1373 4171
rect 1367 4166 1373 4167
rect 1503 4171 1509 4172
rect 1503 4167 1504 4171
rect 1508 4170 1509 4171
rect 1530 4171 1536 4172
rect 1530 4170 1531 4171
rect 1508 4168 1531 4170
rect 1508 4167 1509 4168
rect 1503 4166 1509 4167
rect 1530 4167 1531 4168
rect 1535 4167 1536 4171
rect 1530 4166 1536 4167
rect 1618 4171 1624 4172
rect 1618 4167 1619 4171
rect 1623 4170 1624 4171
rect 1639 4171 1645 4172
rect 1639 4170 1640 4171
rect 1623 4168 1640 4170
rect 1623 4167 1624 4168
rect 1618 4166 1624 4167
rect 1639 4167 1640 4168
rect 1644 4167 1645 4171
rect 1639 4166 1645 4167
rect 1775 4171 1784 4172
rect 1775 4167 1776 4171
rect 1783 4167 1784 4171
rect 1775 4166 1784 4167
rect 1794 4171 1800 4172
rect 1794 4167 1795 4171
rect 1799 4170 1800 4171
rect 1911 4171 1917 4172
rect 1911 4170 1912 4171
rect 1799 4168 1912 4170
rect 1799 4167 1800 4168
rect 1794 4166 1800 4167
rect 1911 4167 1912 4168
rect 1916 4167 1917 4171
rect 1911 4166 1917 4167
rect 791 4160 974 4162
rect 791 4159 792 4160
rect 786 4158 792 4159
rect 4095 4151 4101 4152
rect 4095 4147 4096 4151
rect 4100 4150 4101 4151
rect 4103 4151 4109 4152
rect 4103 4150 4104 4151
rect 4100 4148 4104 4150
rect 4100 4147 4101 4148
rect 4095 4146 4101 4147
rect 4103 4147 4104 4148
rect 4108 4147 4109 4151
rect 4103 4146 4109 4147
rect 4231 4151 4237 4152
rect 4231 4147 4232 4151
rect 4236 4150 4237 4151
rect 4282 4151 4288 4152
rect 4282 4150 4283 4151
rect 4236 4148 4283 4150
rect 4236 4147 4237 4148
rect 4231 4146 4237 4147
rect 4282 4147 4283 4148
rect 4287 4147 4288 4151
rect 4282 4146 4288 4147
rect 4367 4151 4373 4152
rect 4367 4147 4368 4151
rect 4372 4150 4373 4151
rect 4375 4151 4381 4152
rect 4375 4150 4376 4151
rect 4372 4148 4376 4150
rect 4372 4147 4373 4148
rect 4367 4146 4373 4147
rect 4375 4147 4376 4148
rect 4380 4147 4381 4151
rect 4375 4146 4381 4147
rect 4503 4151 4509 4152
rect 4503 4147 4504 4151
rect 4508 4150 4509 4151
rect 4511 4151 4517 4152
rect 4511 4150 4512 4151
rect 4508 4148 4512 4150
rect 4508 4147 4509 4148
rect 4503 4146 4509 4147
rect 4511 4147 4512 4148
rect 4516 4147 4517 4151
rect 4511 4146 4517 4147
rect 4522 4151 4528 4152
rect 4522 4147 4523 4151
rect 4527 4150 4528 4151
rect 4639 4151 4645 4152
rect 4639 4150 4640 4151
rect 4527 4148 4640 4150
rect 4527 4147 4528 4148
rect 4522 4146 4528 4147
rect 4639 4147 4640 4148
rect 4644 4147 4645 4151
rect 4639 4146 4645 4147
rect 3838 4144 3844 4145
rect 5662 4144 5668 4145
rect 3838 4140 3839 4144
rect 3843 4140 3844 4144
rect 786 4139 792 4140
rect 786 4135 787 4139
rect 791 4135 792 4139
rect 786 4134 792 4135
rect 850 4139 856 4140
rect 850 4135 851 4139
rect 855 4135 856 4139
rect 1103 4139 1109 4140
rect 1103 4138 1104 4139
rect 1061 4136 1104 4138
rect 850 4134 856 4135
rect 1103 4135 1104 4136
rect 1108 4135 1109 4139
rect 1239 4139 1245 4140
rect 1239 4138 1240 4139
rect 1197 4136 1240 4138
rect 1103 4134 1109 4135
rect 1239 4135 1240 4136
rect 1244 4135 1245 4139
rect 1239 4134 1245 4135
rect 1330 4139 1336 4140
rect 1330 4135 1331 4139
rect 1335 4135 1336 4139
rect 1330 4134 1336 4135
rect 1466 4139 1472 4140
rect 1466 4135 1467 4139
rect 1471 4135 1472 4139
rect 1466 4134 1472 4135
rect 1530 4139 1536 4140
rect 1530 4135 1531 4139
rect 1535 4135 1536 4139
rect 1794 4139 1800 4140
rect 1794 4138 1795 4139
rect 1741 4136 1795 4138
rect 1530 4134 1536 4135
rect 1794 4135 1795 4136
rect 1799 4135 1800 4139
rect 1946 4139 1952 4140
rect 3838 4139 3844 4140
rect 3970 4143 3976 4144
rect 3970 4139 3971 4143
rect 3975 4139 3976 4143
rect 1946 4138 1947 4139
rect 1877 4136 1947 4138
rect 1794 4134 1800 4135
rect 1946 4135 1947 4136
rect 1951 4135 1952 4139
rect 3970 4138 3976 4139
rect 4106 4143 4112 4144
rect 4106 4139 4107 4143
rect 4111 4139 4112 4143
rect 4106 4138 4112 4139
rect 4242 4143 4248 4144
rect 4242 4139 4243 4143
rect 4247 4139 4248 4143
rect 4242 4138 4248 4139
rect 4378 4143 4384 4144
rect 4378 4139 4379 4143
rect 4383 4139 4384 4143
rect 4378 4138 4384 4139
rect 4514 4143 4520 4144
rect 4514 4139 4515 4143
rect 4519 4139 4520 4143
rect 5662 4140 5663 4144
rect 5667 4140 5668 4144
rect 5662 4139 5668 4140
rect 4514 4138 4520 4139
rect 1946 4134 1952 4135
rect 3998 4128 4004 4129
rect 3838 4127 3844 4128
rect 3838 4123 3839 4127
rect 3843 4123 3844 4127
rect 3998 4124 3999 4128
rect 4003 4124 4004 4128
rect 3998 4123 4004 4124
rect 4134 4128 4140 4129
rect 4134 4124 4135 4128
rect 4139 4124 4140 4128
rect 4134 4123 4140 4124
rect 4270 4128 4276 4129
rect 4270 4124 4271 4128
rect 4275 4124 4276 4128
rect 4270 4123 4276 4124
rect 4406 4128 4412 4129
rect 4406 4124 4407 4128
rect 4411 4124 4412 4128
rect 4406 4123 4412 4124
rect 4542 4128 4548 4129
rect 4542 4124 4543 4128
rect 4547 4124 4548 4128
rect 4542 4123 4548 4124
rect 5662 4127 5668 4128
rect 5662 4123 5663 4127
rect 5667 4123 5668 4127
rect 3838 4122 3844 4123
rect 5662 4122 5668 4123
rect 1974 4109 1980 4110
rect 3798 4109 3804 4110
rect 1974 4105 1975 4109
rect 1979 4105 1980 4109
rect 1974 4104 1980 4105
rect 3134 4108 3140 4109
rect 3134 4104 3135 4108
rect 3139 4104 3140 4108
rect 3134 4103 3140 4104
rect 3270 4108 3276 4109
rect 3270 4104 3271 4108
rect 3275 4104 3276 4108
rect 3270 4103 3276 4104
rect 3406 4108 3412 4109
rect 3406 4104 3407 4108
rect 3411 4104 3412 4108
rect 3406 4103 3412 4104
rect 3542 4108 3548 4109
rect 3542 4104 3543 4108
rect 3547 4104 3548 4108
rect 3542 4103 3548 4104
rect 3678 4108 3684 4109
rect 3678 4104 3679 4108
rect 3683 4104 3684 4108
rect 3798 4105 3799 4109
rect 3803 4105 3804 4109
rect 3798 4104 3804 4105
rect 3678 4103 3684 4104
rect 3106 4093 3112 4094
rect 1974 4092 1980 4093
rect 695 4091 701 4092
rect 650 4087 656 4088
rect 650 4083 651 4087
rect 655 4083 656 4087
rect 695 4087 696 4091
rect 700 4090 701 4091
rect 831 4091 837 4092
rect 700 4088 717 4090
rect 700 4087 701 4088
rect 695 4086 701 4087
rect 831 4087 832 4091
rect 836 4090 837 4091
rect 962 4091 968 4092
rect 836 4088 853 4090
rect 836 4087 837 4088
rect 831 4086 837 4087
rect 962 4087 963 4091
rect 967 4090 968 4091
rect 1103 4091 1109 4092
rect 967 4088 989 4090
rect 967 4087 968 4088
rect 962 4086 968 4087
rect 1103 4087 1104 4091
rect 1108 4090 1109 4091
rect 1375 4091 1381 4092
rect 1108 4088 1125 4090
rect 1108 4087 1109 4088
rect 1103 4086 1109 4087
rect 1375 4087 1376 4091
rect 1380 4090 1381 4091
rect 1647 4091 1653 4092
rect 1647 4090 1648 4091
rect 1380 4088 1397 4090
rect 1605 4088 1648 4090
rect 1380 4087 1381 4088
rect 1375 4086 1381 4087
rect 1647 4087 1648 4088
rect 1652 4087 1653 4091
rect 1647 4086 1653 4087
rect 1778 4091 1784 4092
rect 1778 4087 1779 4091
rect 1783 4090 1784 4091
rect 1783 4088 1805 4090
rect 1974 4088 1975 4092
rect 1979 4088 1980 4092
rect 3106 4089 3107 4093
rect 3111 4089 3112 4093
rect 3106 4088 3112 4089
rect 3242 4093 3248 4094
rect 3242 4089 3243 4093
rect 3247 4089 3248 4093
rect 3242 4088 3248 4089
rect 3378 4093 3384 4094
rect 3378 4089 3379 4093
rect 3383 4089 3384 4093
rect 3378 4088 3384 4089
rect 3514 4093 3520 4094
rect 3514 4089 3515 4093
rect 3519 4089 3520 4093
rect 3514 4088 3520 4089
rect 3650 4093 3656 4094
rect 3650 4089 3651 4093
rect 3655 4089 3656 4093
rect 3650 4088 3656 4089
rect 3798 4092 3804 4093
rect 3798 4088 3799 4092
rect 3803 4088 3804 4092
rect 1783 4087 1784 4088
rect 1974 4087 1980 4088
rect 3798 4087 3804 4088
rect 1778 4086 1784 4087
rect 650 4082 656 4083
rect 1328 4074 1330 4085
rect 1736 4082 1738 4085
rect 1783 4083 1789 4084
rect 1783 4082 1784 4083
rect 1736 4080 1784 4082
rect 1783 4079 1784 4080
rect 1788 4079 1789 4083
rect 1783 4078 1789 4079
rect 3231 4083 3237 4084
rect 3231 4079 3232 4083
rect 3236 4082 3237 4083
rect 3258 4083 3264 4084
rect 3258 4082 3259 4083
rect 3236 4080 3259 4082
rect 3236 4079 3237 4080
rect 3231 4078 3237 4079
rect 3258 4079 3259 4080
rect 3263 4079 3264 4083
rect 3258 4078 3264 4079
rect 3367 4083 3376 4084
rect 3367 4079 3368 4083
rect 3375 4079 3376 4083
rect 3503 4083 3509 4084
rect 3503 4082 3504 4083
rect 3367 4078 3376 4079
rect 3380 4080 3504 4082
rect 1474 4075 1480 4076
rect 1474 4074 1475 4075
rect 1328 4072 1475 4074
rect 1474 4071 1475 4072
rect 1479 4071 1480 4075
rect 1474 4070 1480 4071
rect 3194 4075 3200 4076
rect 3194 4071 3195 4075
rect 3199 4074 3200 4075
rect 3380 4074 3382 4080
rect 3503 4079 3504 4080
rect 3508 4079 3509 4083
rect 3503 4078 3509 4079
rect 3511 4083 3517 4084
rect 3511 4079 3512 4083
rect 3516 4082 3517 4083
rect 3639 4083 3645 4084
rect 3639 4082 3640 4083
rect 3516 4080 3640 4082
rect 3516 4079 3517 4080
rect 3511 4078 3517 4079
rect 3639 4079 3640 4080
rect 3644 4079 3645 4083
rect 3639 4078 3645 4079
rect 3647 4083 3653 4084
rect 3647 4079 3648 4083
rect 3652 4082 3653 4083
rect 3775 4083 3781 4084
rect 3775 4082 3776 4083
rect 3652 4080 3776 4082
rect 3652 4079 3653 4080
rect 3647 4078 3653 4079
rect 3775 4079 3776 4080
rect 3780 4079 3781 4083
rect 3775 4078 3781 4079
rect 3199 4072 3382 4074
rect 3199 4071 3200 4072
rect 3194 4070 3200 4071
rect 650 4063 656 4064
rect 650 4059 651 4063
rect 655 4062 656 4063
rect 655 4060 1114 4062
rect 655 4059 656 4060
rect 650 4058 656 4059
rect 687 4055 693 4056
rect 687 4051 688 4055
rect 692 4054 693 4055
rect 695 4055 701 4056
rect 695 4054 696 4055
rect 692 4052 696 4054
rect 692 4051 693 4052
rect 687 4050 693 4051
rect 695 4051 696 4052
rect 700 4051 701 4055
rect 695 4050 701 4051
rect 823 4055 829 4056
rect 823 4051 824 4055
rect 828 4054 829 4055
rect 831 4055 837 4056
rect 831 4054 832 4055
rect 828 4052 832 4054
rect 828 4051 829 4052
rect 823 4050 829 4051
rect 831 4051 832 4052
rect 836 4051 837 4055
rect 831 4050 837 4051
rect 958 4055 965 4056
rect 958 4051 959 4055
rect 964 4051 965 4055
rect 958 4050 965 4051
rect 1095 4055 1101 4056
rect 1095 4051 1096 4055
rect 1100 4054 1101 4055
rect 1103 4055 1109 4056
rect 1103 4054 1104 4055
rect 1100 4052 1104 4054
rect 1100 4051 1101 4052
rect 1095 4050 1101 4051
rect 1103 4051 1104 4052
rect 1108 4051 1109 4055
rect 1112 4054 1114 4060
rect 1231 4055 1237 4056
rect 1231 4054 1232 4055
rect 1112 4052 1232 4054
rect 1103 4050 1109 4051
rect 1231 4051 1232 4052
rect 1236 4051 1237 4055
rect 1231 4050 1237 4051
rect 1367 4055 1373 4056
rect 1367 4051 1368 4055
rect 1372 4054 1373 4055
rect 1375 4055 1381 4056
rect 1375 4054 1376 4055
rect 1372 4052 1376 4054
rect 1372 4051 1373 4052
rect 1367 4050 1373 4051
rect 1375 4051 1376 4052
rect 1380 4051 1381 4055
rect 1375 4050 1381 4051
rect 1466 4055 1472 4056
rect 1466 4051 1467 4055
rect 1471 4054 1472 4055
rect 1503 4055 1509 4056
rect 1503 4054 1504 4055
rect 1471 4052 1504 4054
rect 1471 4051 1472 4052
rect 1466 4050 1472 4051
rect 1503 4051 1504 4052
rect 1508 4051 1509 4055
rect 1503 4050 1509 4051
rect 1638 4055 1645 4056
rect 1638 4051 1639 4055
rect 1644 4051 1645 4055
rect 1638 4050 1645 4051
rect 1647 4055 1653 4056
rect 1647 4051 1648 4055
rect 1652 4054 1653 4055
rect 1775 4055 1781 4056
rect 1775 4054 1776 4055
rect 1652 4052 1776 4054
rect 1652 4051 1653 4052
rect 1647 4050 1653 4051
rect 1775 4051 1776 4052
rect 1780 4051 1781 4055
rect 1775 4050 1781 4051
rect 1783 4055 1789 4056
rect 1783 4051 1784 4055
rect 1788 4054 1789 4055
rect 1911 4055 1917 4056
rect 1911 4054 1912 4055
rect 1788 4052 1912 4054
rect 1788 4051 1789 4052
rect 1783 4050 1789 4051
rect 1911 4051 1912 4052
rect 1916 4051 1917 4055
rect 1911 4050 1917 4051
rect 3194 4051 3200 4052
rect 110 4048 116 4049
rect 1934 4048 1940 4049
rect 110 4044 111 4048
rect 115 4044 116 4048
rect 110 4043 116 4044
rect 562 4047 568 4048
rect 562 4043 563 4047
rect 567 4043 568 4047
rect 562 4042 568 4043
rect 698 4047 704 4048
rect 698 4043 699 4047
rect 703 4043 704 4047
rect 698 4042 704 4043
rect 834 4047 840 4048
rect 834 4043 835 4047
rect 839 4043 840 4047
rect 834 4042 840 4043
rect 970 4047 976 4048
rect 970 4043 971 4047
rect 975 4043 976 4047
rect 970 4042 976 4043
rect 1106 4047 1112 4048
rect 1106 4043 1107 4047
rect 1111 4043 1112 4047
rect 1106 4042 1112 4043
rect 1242 4047 1248 4048
rect 1242 4043 1243 4047
rect 1247 4043 1248 4047
rect 1242 4042 1248 4043
rect 1378 4047 1384 4048
rect 1378 4043 1379 4047
rect 1383 4043 1384 4047
rect 1378 4042 1384 4043
rect 1514 4047 1520 4048
rect 1514 4043 1515 4047
rect 1519 4043 1520 4047
rect 1514 4042 1520 4043
rect 1650 4047 1656 4048
rect 1650 4043 1651 4047
rect 1655 4043 1656 4047
rect 1650 4042 1656 4043
rect 1786 4047 1792 4048
rect 1786 4043 1787 4047
rect 1791 4043 1792 4047
rect 1934 4044 1935 4048
rect 1939 4044 1940 4048
rect 3194 4047 3195 4051
rect 3199 4047 3200 4051
rect 3194 4046 3200 4047
rect 3258 4051 3264 4052
rect 3258 4047 3259 4051
rect 3263 4047 3264 4051
rect 3511 4051 3517 4052
rect 3511 4050 3512 4051
rect 3469 4048 3512 4050
rect 3258 4046 3264 4047
rect 3511 4047 3512 4048
rect 3516 4047 3517 4051
rect 3647 4051 3653 4052
rect 3647 4050 3648 4051
rect 3605 4048 3648 4050
rect 3511 4046 3517 4047
rect 3647 4047 3648 4048
rect 3652 4047 3653 4051
rect 3647 4046 3653 4047
rect 3738 4051 3744 4052
rect 3738 4047 3739 4051
rect 3743 4047 3744 4051
rect 3738 4046 3744 4047
rect 1934 4043 1940 4044
rect 3838 4045 3844 4046
rect 5662 4045 5668 4046
rect 1786 4042 1792 4043
rect 3838 4041 3839 4045
rect 3843 4041 3844 4045
rect 3838 4040 3844 4041
rect 3886 4044 3892 4045
rect 3886 4040 3887 4044
rect 3891 4040 3892 4044
rect 3886 4039 3892 4040
rect 4022 4044 4028 4045
rect 4022 4040 4023 4044
rect 4027 4040 4028 4044
rect 4022 4039 4028 4040
rect 4158 4044 4164 4045
rect 4158 4040 4159 4044
rect 4163 4040 4164 4044
rect 4158 4039 4164 4040
rect 4294 4044 4300 4045
rect 4294 4040 4295 4044
rect 4299 4040 4300 4044
rect 4294 4039 4300 4040
rect 4430 4044 4436 4045
rect 4430 4040 4431 4044
rect 4435 4040 4436 4044
rect 4430 4039 4436 4040
rect 4566 4044 4572 4045
rect 4566 4040 4567 4044
rect 4571 4040 4572 4044
rect 4566 4039 4572 4040
rect 4702 4044 4708 4045
rect 4702 4040 4703 4044
rect 4707 4040 4708 4044
rect 4702 4039 4708 4040
rect 4838 4044 4844 4045
rect 4838 4040 4839 4044
rect 4843 4040 4844 4044
rect 5662 4041 5663 4045
rect 5667 4041 5668 4045
rect 5662 4040 5668 4041
rect 4838 4039 4844 4040
rect 590 4032 596 4033
rect 110 4031 116 4032
rect 110 4027 111 4031
rect 115 4027 116 4031
rect 590 4028 591 4032
rect 595 4028 596 4032
rect 590 4027 596 4028
rect 726 4032 732 4033
rect 726 4028 727 4032
rect 731 4028 732 4032
rect 726 4027 732 4028
rect 862 4032 868 4033
rect 862 4028 863 4032
rect 867 4028 868 4032
rect 862 4027 868 4028
rect 998 4032 1004 4033
rect 998 4028 999 4032
rect 1003 4028 1004 4032
rect 998 4027 1004 4028
rect 1134 4032 1140 4033
rect 1134 4028 1135 4032
rect 1139 4028 1140 4032
rect 1134 4027 1140 4028
rect 1270 4032 1276 4033
rect 1270 4028 1271 4032
rect 1275 4028 1276 4032
rect 1270 4027 1276 4028
rect 1406 4032 1412 4033
rect 1406 4028 1407 4032
rect 1411 4028 1412 4032
rect 1406 4027 1412 4028
rect 1542 4032 1548 4033
rect 1542 4028 1543 4032
rect 1547 4028 1548 4032
rect 1542 4027 1548 4028
rect 1678 4032 1684 4033
rect 1678 4028 1679 4032
rect 1683 4028 1684 4032
rect 1678 4027 1684 4028
rect 1814 4032 1820 4033
rect 1814 4028 1815 4032
rect 1819 4028 1820 4032
rect 1814 4027 1820 4028
rect 1934 4031 1940 4032
rect 1934 4027 1935 4031
rect 1939 4027 1940 4031
rect 3858 4029 3864 4030
rect 110 4026 116 4027
rect 1934 4026 1940 4027
rect 3838 4028 3844 4029
rect 3838 4024 3839 4028
rect 3843 4024 3844 4028
rect 3858 4025 3859 4029
rect 3863 4025 3864 4029
rect 3858 4024 3864 4025
rect 3994 4029 4000 4030
rect 3994 4025 3995 4029
rect 3999 4025 4000 4029
rect 3994 4024 4000 4025
rect 4130 4029 4136 4030
rect 4130 4025 4131 4029
rect 4135 4025 4136 4029
rect 4130 4024 4136 4025
rect 4266 4029 4272 4030
rect 4266 4025 4267 4029
rect 4271 4025 4272 4029
rect 4266 4024 4272 4025
rect 4402 4029 4408 4030
rect 4402 4025 4403 4029
rect 4407 4025 4408 4029
rect 4402 4024 4408 4025
rect 4538 4029 4544 4030
rect 4538 4025 4539 4029
rect 4543 4025 4544 4029
rect 4538 4024 4544 4025
rect 4674 4029 4680 4030
rect 4674 4025 4675 4029
rect 4679 4025 4680 4029
rect 4674 4024 4680 4025
rect 4810 4029 4816 4030
rect 4810 4025 4811 4029
rect 4815 4025 4816 4029
rect 4810 4024 4816 4025
rect 5662 4028 5668 4029
rect 5662 4024 5663 4028
rect 5667 4024 5668 4028
rect 3838 4023 3844 4024
rect 5662 4023 5668 4024
rect 3738 4019 3744 4020
rect 3738 4015 3739 4019
rect 3743 4018 3744 4019
rect 3983 4019 3989 4020
rect 3983 4018 3984 4019
rect 3743 4016 3984 4018
rect 3743 4015 3744 4016
rect 3738 4014 3744 4015
rect 3983 4015 3984 4016
rect 3988 4015 3989 4019
rect 3983 4014 3989 4015
rect 4002 4019 4008 4020
rect 4002 4015 4003 4019
rect 4007 4018 4008 4019
rect 4119 4019 4125 4020
rect 4119 4018 4120 4019
rect 4007 4016 4120 4018
rect 4007 4015 4008 4016
rect 4002 4014 4008 4015
rect 4119 4015 4120 4016
rect 4124 4015 4125 4019
rect 4255 4019 4261 4020
rect 4255 4018 4256 4019
rect 4119 4014 4125 4015
rect 4128 4016 4256 4018
rect 4082 4011 4088 4012
rect 4082 4007 4083 4011
rect 4087 4010 4088 4011
rect 4128 4010 4130 4016
rect 4255 4015 4256 4016
rect 4260 4015 4261 4019
rect 4255 4014 4261 4015
rect 4391 4019 4397 4020
rect 4391 4015 4392 4019
rect 4396 4018 4397 4019
rect 4418 4019 4424 4020
rect 4418 4018 4419 4019
rect 4396 4016 4419 4018
rect 4396 4015 4397 4016
rect 4391 4014 4397 4015
rect 4418 4015 4419 4016
rect 4423 4015 4424 4019
rect 4418 4014 4424 4015
rect 4527 4019 4533 4020
rect 4527 4015 4528 4019
rect 4532 4018 4533 4019
rect 4554 4019 4560 4020
rect 4554 4018 4555 4019
rect 4532 4016 4555 4018
rect 4532 4015 4533 4016
rect 4527 4014 4533 4015
rect 4554 4015 4555 4016
rect 4559 4015 4560 4019
rect 4554 4014 4560 4015
rect 4663 4019 4669 4020
rect 4663 4015 4664 4019
rect 4668 4018 4669 4019
rect 4690 4019 4696 4020
rect 4690 4018 4691 4019
rect 4668 4016 4691 4018
rect 4668 4015 4669 4016
rect 4663 4014 4669 4015
rect 4690 4015 4691 4016
rect 4695 4015 4696 4019
rect 4690 4014 4696 4015
rect 4799 4019 4805 4020
rect 4799 4015 4800 4019
rect 4804 4018 4805 4019
rect 4826 4019 4832 4020
rect 4826 4018 4827 4019
rect 4804 4016 4827 4018
rect 4804 4015 4805 4016
rect 4799 4014 4805 4015
rect 4826 4015 4827 4016
rect 4831 4015 4832 4019
rect 4935 4019 4941 4020
rect 4935 4018 4936 4019
rect 4826 4014 4832 4015
rect 4864 4016 4936 4018
rect 4087 4008 4130 4010
rect 4263 4011 4269 4012
rect 4087 4007 4088 4008
rect 4082 4006 4088 4007
rect 4263 4007 4264 4011
rect 4268 4010 4269 4011
rect 4864 4010 4866 4016
rect 4935 4015 4936 4016
rect 4940 4015 4941 4019
rect 4935 4014 4941 4015
rect 4268 4008 4866 4010
rect 4268 4007 4269 4008
rect 4263 4006 4269 4007
rect 4002 3987 4008 3988
rect 4002 3986 4003 3987
rect 3949 3984 4003 3986
rect 4002 3983 4003 3984
rect 4007 3983 4008 3987
rect 4002 3982 4008 3983
rect 4082 3987 4088 3988
rect 4082 3983 4083 3987
rect 4087 3983 4088 3987
rect 4082 3982 4088 3983
rect 4122 3987 4128 3988
rect 4122 3983 4123 3987
rect 4127 3986 4128 3987
rect 4282 3987 4288 3988
rect 4127 3984 4149 3986
rect 4127 3983 4128 3984
rect 4122 3982 4128 3983
rect 4282 3983 4283 3987
rect 4287 3983 4288 3987
rect 4282 3982 4288 3983
rect 4418 3987 4424 3988
rect 4418 3983 4419 3987
rect 4423 3983 4424 3987
rect 4418 3982 4424 3983
rect 4554 3987 4560 3988
rect 4554 3983 4555 3987
rect 4559 3983 4560 3987
rect 4554 3982 4560 3983
rect 4690 3987 4696 3988
rect 4690 3983 4691 3987
rect 4695 3983 4696 3987
rect 4690 3982 4696 3983
rect 4826 3987 4832 3988
rect 4826 3983 4827 3987
rect 4831 3983 4832 3987
rect 4826 3982 4832 3983
rect 110 3973 116 3974
rect 1934 3973 1940 3974
rect 110 3969 111 3973
rect 115 3969 116 3973
rect 110 3968 116 3969
rect 158 3972 164 3973
rect 158 3968 159 3972
rect 163 3968 164 3972
rect 158 3967 164 3968
rect 326 3972 332 3973
rect 326 3968 327 3972
rect 331 3968 332 3972
rect 326 3967 332 3968
rect 534 3972 540 3973
rect 534 3968 535 3972
rect 539 3968 540 3972
rect 534 3967 540 3968
rect 750 3972 756 3973
rect 750 3968 751 3972
rect 755 3968 756 3972
rect 750 3967 756 3968
rect 966 3972 972 3973
rect 966 3968 967 3972
rect 971 3968 972 3972
rect 966 3967 972 3968
rect 1182 3972 1188 3973
rect 1182 3968 1183 3972
rect 1187 3968 1188 3972
rect 1182 3967 1188 3968
rect 1398 3972 1404 3973
rect 1398 3968 1399 3972
rect 1403 3968 1404 3972
rect 1398 3967 1404 3968
rect 1614 3972 1620 3973
rect 1614 3968 1615 3972
rect 1619 3968 1620 3972
rect 1614 3967 1620 3968
rect 1814 3972 1820 3973
rect 1814 3968 1815 3972
rect 1819 3968 1820 3972
rect 1934 3969 1935 3973
rect 1939 3969 1940 3973
rect 1934 3968 1940 3969
rect 1814 3967 1820 3968
rect 130 3957 136 3958
rect 110 3956 116 3957
rect 110 3952 111 3956
rect 115 3952 116 3956
rect 130 3953 131 3957
rect 135 3953 136 3957
rect 130 3952 136 3953
rect 298 3957 304 3958
rect 298 3953 299 3957
rect 303 3953 304 3957
rect 298 3952 304 3953
rect 506 3957 512 3958
rect 506 3953 507 3957
rect 511 3953 512 3957
rect 506 3952 512 3953
rect 722 3957 728 3958
rect 722 3953 723 3957
rect 727 3953 728 3957
rect 722 3952 728 3953
rect 938 3957 944 3958
rect 938 3953 939 3957
rect 943 3953 944 3957
rect 938 3952 944 3953
rect 1154 3957 1160 3958
rect 1154 3953 1155 3957
rect 1159 3953 1160 3957
rect 1154 3952 1160 3953
rect 1370 3957 1376 3958
rect 1370 3953 1371 3957
rect 1375 3953 1376 3957
rect 1370 3952 1376 3953
rect 1586 3957 1592 3958
rect 1586 3953 1587 3957
rect 1591 3953 1592 3957
rect 1586 3952 1592 3953
rect 1786 3957 1792 3958
rect 1786 3953 1787 3957
rect 1791 3953 1792 3957
rect 1786 3952 1792 3953
rect 1934 3956 1940 3957
rect 1934 3952 1935 3956
rect 1939 3952 1940 3956
rect 110 3951 116 3952
rect 1934 3951 1940 3952
rect 234 3947 240 3948
rect 234 3943 235 3947
rect 239 3946 240 3947
rect 255 3947 261 3948
rect 255 3946 256 3947
rect 239 3944 256 3946
rect 239 3943 240 3944
rect 234 3942 240 3943
rect 255 3943 256 3944
rect 260 3943 261 3947
rect 255 3942 261 3943
rect 286 3947 292 3948
rect 286 3943 287 3947
rect 291 3946 292 3947
rect 423 3947 429 3948
rect 423 3946 424 3947
rect 291 3944 424 3946
rect 291 3943 292 3944
rect 286 3942 292 3943
rect 423 3943 424 3944
rect 428 3943 429 3947
rect 423 3942 429 3943
rect 450 3947 456 3948
rect 450 3943 451 3947
rect 455 3946 456 3947
rect 631 3947 637 3948
rect 631 3946 632 3947
rect 455 3944 632 3946
rect 455 3943 456 3944
rect 450 3942 456 3943
rect 631 3943 632 3944
rect 636 3943 637 3947
rect 631 3942 637 3943
rect 702 3947 708 3948
rect 702 3943 703 3947
rect 707 3946 708 3947
rect 847 3947 853 3948
rect 847 3946 848 3947
rect 707 3944 848 3946
rect 707 3943 708 3944
rect 702 3942 708 3943
rect 847 3943 848 3944
rect 852 3943 853 3947
rect 847 3942 853 3943
rect 878 3947 884 3948
rect 878 3943 879 3947
rect 883 3946 884 3947
rect 1063 3947 1069 3948
rect 1063 3946 1064 3947
rect 883 3944 1064 3946
rect 883 3943 884 3944
rect 878 3942 884 3943
rect 1063 3943 1064 3944
rect 1068 3943 1069 3947
rect 1063 3942 1069 3943
rect 1279 3947 1285 3948
rect 1279 3943 1280 3947
rect 1284 3946 1285 3947
rect 1386 3947 1392 3948
rect 1386 3946 1387 3947
rect 1284 3944 1387 3946
rect 1284 3943 1285 3944
rect 1279 3942 1285 3943
rect 1386 3943 1387 3944
rect 1391 3943 1392 3947
rect 1386 3942 1392 3943
rect 1474 3947 1480 3948
rect 1474 3943 1475 3947
rect 1479 3946 1480 3947
rect 1495 3947 1501 3948
rect 1495 3946 1496 3947
rect 1479 3944 1496 3946
rect 1479 3943 1480 3944
rect 1474 3942 1480 3943
rect 1495 3943 1496 3944
rect 1500 3943 1501 3947
rect 1495 3942 1501 3943
rect 1711 3947 1717 3948
rect 1711 3943 1712 3947
rect 1716 3946 1717 3947
rect 1802 3947 1808 3948
rect 1802 3946 1803 3947
rect 1716 3944 1803 3946
rect 1716 3943 1717 3944
rect 1711 3942 1717 3943
rect 1802 3943 1803 3944
rect 1807 3943 1808 3947
rect 1802 3942 1808 3943
rect 1890 3947 1896 3948
rect 1890 3943 1891 3947
rect 1895 3946 1896 3947
rect 1911 3947 1917 3948
rect 1911 3946 1912 3947
rect 1895 3944 1912 3946
rect 1895 3943 1896 3944
rect 1890 3942 1896 3943
rect 1911 3943 1912 3944
rect 1916 3943 1917 3947
rect 1911 3942 1917 3943
rect 3778 3939 3784 3940
rect 3778 3935 3779 3939
rect 3783 3938 3784 3939
rect 3986 3939 3992 3940
rect 3783 3936 3877 3938
rect 3783 3935 3784 3936
rect 3778 3934 3784 3935
rect 3986 3935 3987 3939
rect 3991 3938 3992 3939
rect 4263 3939 4269 3940
rect 4263 3938 4264 3939
rect 3991 3936 4013 3938
rect 4237 3936 4264 3938
rect 3991 3935 3992 3936
rect 3986 3934 3992 3935
rect 4263 3935 4264 3936
rect 4268 3935 4269 3939
rect 4263 3934 4269 3935
rect 4274 3939 4280 3940
rect 4274 3935 4275 3939
rect 4279 3938 4280 3939
rect 4450 3939 4456 3940
rect 4279 3936 4317 3938
rect 4279 3935 4280 3936
rect 4274 3934 4280 3935
rect 4450 3935 4451 3939
rect 4455 3938 4456 3939
rect 4610 3939 4616 3940
rect 4455 3936 4477 3938
rect 4455 3935 4456 3936
rect 4450 3934 4456 3935
rect 4610 3935 4611 3939
rect 4615 3938 4616 3939
rect 4770 3939 4776 3940
rect 4615 3936 4637 3938
rect 4615 3935 4616 3936
rect 4610 3934 4616 3935
rect 4770 3935 4771 3939
rect 4775 3938 4776 3939
rect 4775 3936 4797 3938
rect 4775 3935 4776 3936
rect 4770 3934 4776 3935
rect 286 3915 292 3916
rect 286 3914 287 3915
rect 221 3912 287 3914
rect 286 3911 287 3912
rect 291 3911 292 3915
rect 450 3915 456 3916
rect 450 3914 451 3915
rect 389 3912 451 3914
rect 286 3910 292 3911
rect 450 3911 451 3912
rect 455 3911 456 3915
rect 702 3915 708 3916
rect 702 3914 703 3915
rect 597 3912 703 3914
rect 450 3910 456 3911
rect 702 3911 703 3912
rect 707 3911 708 3915
rect 878 3915 884 3916
rect 878 3914 879 3915
rect 813 3912 879 3914
rect 702 3910 708 3911
rect 878 3911 879 3912
rect 883 3911 884 3915
rect 878 3910 884 3911
rect 958 3915 964 3916
rect 958 3911 959 3915
rect 963 3911 964 3915
rect 958 3910 964 3911
rect 1242 3915 1248 3916
rect 1242 3911 1243 3915
rect 1247 3911 1248 3915
rect 1242 3910 1248 3911
rect 1386 3915 1392 3916
rect 1386 3911 1387 3915
rect 1391 3911 1392 3915
rect 1386 3910 1392 3911
rect 1638 3915 1644 3916
rect 1638 3911 1639 3915
rect 1643 3911 1644 3915
rect 1638 3910 1644 3911
rect 1802 3915 1808 3916
rect 1802 3911 1803 3915
rect 1807 3911 1808 3915
rect 1802 3910 1808 3911
rect 1914 3911 1920 3912
rect 1914 3907 1915 3911
rect 1919 3910 1920 3911
rect 2522 3911 2528 3912
rect 2522 3910 2523 3911
rect 1919 3908 2013 3910
rect 2493 3908 2523 3910
rect 1919 3907 1920 3908
rect 1914 3906 1920 3907
rect 2522 3907 2523 3908
rect 2527 3907 2528 3911
rect 2522 3906 2528 3907
rect 2530 3911 2536 3912
rect 2530 3907 2531 3911
rect 2535 3910 2536 3911
rect 2954 3911 2960 3912
rect 2535 3908 2845 3910
rect 2535 3907 2536 3908
rect 2530 3906 2536 3907
rect 2954 3907 2955 3911
rect 2959 3910 2960 3911
rect 3378 3911 3384 3912
rect 2959 3908 3269 3910
rect 2959 3907 2960 3908
rect 2954 3906 2960 3907
rect 3378 3907 3379 3911
rect 3383 3910 3384 3911
rect 3383 3908 3669 3910
rect 3383 3907 3384 3908
rect 3378 3906 3384 3907
rect 3983 3903 3992 3904
rect 3983 3899 3984 3903
rect 3991 3899 3992 3903
rect 3983 3898 3992 3899
rect 4119 3903 4128 3904
rect 4119 3899 4120 3903
rect 4127 3899 4128 3903
rect 4119 3898 4128 3899
rect 4271 3903 4280 3904
rect 4271 3899 4272 3903
rect 4279 3899 4280 3903
rect 4271 3898 4280 3899
rect 4423 3903 4429 3904
rect 4423 3899 4424 3903
rect 4428 3902 4429 3903
rect 4450 3903 4456 3904
rect 4450 3902 4451 3903
rect 4428 3900 4451 3902
rect 4428 3899 4429 3900
rect 4423 3898 4429 3899
rect 4450 3899 4451 3900
rect 4455 3899 4456 3903
rect 4450 3898 4456 3899
rect 4583 3903 4589 3904
rect 4583 3899 4584 3903
rect 4588 3902 4589 3903
rect 4610 3903 4616 3904
rect 4610 3902 4611 3903
rect 4588 3900 4611 3902
rect 4588 3899 4589 3900
rect 4583 3898 4589 3899
rect 4610 3899 4611 3900
rect 4615 3899 4616 3903
rect 4610 3898 4616 3899
rect 4743 3903 4749 3904
rect 4743 3899 4744 3903
rect 4748 3902 4749 3903
rect 4770 3903 4776 3904
rect 4770 3902 4771 3903
rect 4748 3900 4771 3902
rect 4748 3899 4749 3900
rect 4743 3898 4749 3899
rect 4770 3899 4771 3900
rect 4775 3899 4776 3903
rect 4770 3898 4776 3899
rect 4786 3903 4792 3904
rect 4786 3899 4787 3903
rect 4791 3902 4792 3903
rect 4903 3903 4909 3904
rect 4903 3902 4904 3903
rect 4791 3900 4904 3902
rect 4791 3899 4792 3900
rect 4786 3898 4792 3899
rect 4903 3899 4904 3900
rect 4908 3899 4909 3903
rect 4903 3898 4909 3899
rect 3838 3896 3844 3897
rect 5662 3896 5668 3897
rect 3838 3892 3839 3896
rect 3843 3892 3844 3896
rect 3838 3891 3844 3892
rect 3858 3895 3864 3896
rect 3858 3891 3859 3895
rect 3863 3891 3864 3895
rect 3858 3890 3864 3891
rect 3994 3895 4000 3896
rect 3994 3891 3995 3895
rect 3999 3891 4000 3895
rect 3994 3890 4000 3891
rect 4146 3895 4152 3896
rect 4146 3891 4147 3895
rect 4151 3891 4152 3895
rect 4146 3890 4152 3891
rect 4298 3895 4304 3896
rect 4298 3891 4299 3895
rect 4303 3891 4304 3895
rect 4298 3890 4304 3891
rect 4458 3895 4464 3896
rect 4458 3891 4459 3895
rect 4463 3891 4464 3895
rect 4458 3890 4464 3891
rect 4618 3895 4624 3896
rect 4618 3891 4619 3895
rect 4623 3891 4624 3895
rect 4618 3890 4624 3891
rect 4778 3895 4784 3896
rect 4778 3891 4779 3895
rect 4783 3891 4784 3895
rect 5662 3892 5663 3896
rect 5667 3892 5668 3896
rect 5662 3891 5668 3892
rect 4778 3890 4784 3891
rect 3886 3880 3892 3881
rect 3838 3879 3844 3880
rect 2082 3875 2088 3876
rect 2082 3871 2083 3875
rect 2087 3874 2088 3875
rect 2119 3875 2125 3876
rect 2119 3874 2120 3875
rect 2087 3872 2120 3874
rect 2087 3871 2088 3872
rect 2082 3870 2088 3871
rect 2119 3871 2120 3872
rect 2124 3871 2125 3875
rect 2119 3870 2125 3871
rect 2527 3875 2536 3876
rect 2527 3871 2528 3875
rect 2535 3871 2536 3875
rect 2527 3870 2536 3871
rect 2951 3875 2960 3876
rect 2951 3871 2952 3875
rect 2959 3871 2960 3875
rect 2951 3870 2960 3871
rect 3375 3875 3384 3876
rect 3375 3871 3376 3875
rect 3383 3871 3384 3875
rect 3375 3870 3384 3871
rect 3775 3875 3784 3876
rect 3775 3871 3776 3875
rect 3783 3871 3784 3875
rect 3838 3875 3839 3879
rect 3843 3875 3844 3879
rect 3886 3876 3887 3880
rect 3891 3876 3892 3880
rect 3886 3875 3892 3876
rect 4022 3880 4028 3881
rect 4022 3876 4023 3880
rect 4027 3876 4028 3880
rect 4022 3875 4028 3876
rect 4174 3880 4180 3881
rect 4174 3876 4175 3880
rect 4179 3876 4180 3880
rect 4174 3875 4180 3876
rect 4326 3880 4332 3881
rect 4326 3876 4327 3880
rect 4331 3876 4332 3880
rect 4326 3875 4332 3876
rect 4486 3880 4492 3881
rect 4486 3876 4487 3880
rect 4491 3876 4492 3880
rect 4486 3875 4492 3876
rect 4646 3880 4652 3881
rect 4646 3876 4647 3880
rect 4651 3876 4652 3880
rect 4646 3875 4652 3876
rect 4806 3880 4812 3881
rect 4806 3876 4807 3880
rect 4811 3876 4812 3880
rect 4806 3875 4812 3876
rect 5662 3879 5668 3880
rect 5662 3875 5663 3879
rect 5667 3875 5668 3879
rect 3838 3874 3844 3875
rect 5662 3874 5668 3875
rect 3775 3870 3784 3871
rect 1974 3868 1980 3869
rect 3798 3868 3804 3869
rect 234 3867 240 3868
rect 234 3866 235 3867
rect 221 3864 235 3866
rect 234 3863 235 3864
rect 239 3863 240 3867
rect 234 3862 240 3863
rect 258 3867 264 3868
rect 258 3863 259 3867
rect 263 3866 264 3867
rect 482 3867 488 3868
rect 263 3864 373 3866
rect 263 3863 264 3864
rect 258 3862 264 3863
rect 482 3863 483 3867
rect 487 3866 488 3867
rect 746 3867 752 3868
rect 487 3864 637 3866
rect 487 3863 488 3864
rect 482 3862 488 3863
rect 746 3863 747 3867
rect 751 3866 752 3867
rect 1334 3867 1340 3868
rect 1334 3866 1335 3867
rect 751 3864 917 3866
rect 1285 3864 1335 3866
rect 751 3863 752 3864
rect 746 3862 752 3863
rect 1334 3863 1335 3864
rect 1339 3863 1340 3867
rect 1334 3862 1340 3863
rect 1447 3867 1453 3868
rect 1447 3863 1448 3867
rect 1452 3866 1453 3867
rect 1890 3867 1896 3868
rect 1890 3866 1891 3867
rect 1452 3864 1517 3866
rect 1877 3864 1891 3866
rect 1452 3863 1453 3864
rect 1447 3862 1453 3863
rect 1890 3863 1891 3864
rect 1895 3863 1896 3867
rect 1974 3864 1975 3868
rect 1979 3864 1980 3868
rect 1974 3863 1980 3864
rect 1994 3867 2000 3868
rect 1994 3863 1995 3867
rect 1999 3863 2000 3867
rect 1890 3862 1896 3863
rect 1994 3862 2000 3863
rect 2402 3867 2408 3868
rect 2402 3863 2403 3867
rect 2407 3863 2408 3867
rect 2402 3862 2408 3863
rect 2826 3867 2832 3868
rect 2826 3863 2827 3867
rect 2831 3863 2832 3867
rect 2826 3862 2832 3863
rect 3250 3867 3256 3868
rect 3250 3863 3251 3867
rect 3255 3863 3256 3867
rect 3250 3862 3256 3863
rect 3650 3867 3656 3868
rect 3650 3863 3651 3867
rect 3655 3863 3656 3867
rect 3798 3864 3799 3868
rect 3803 3864 3804 3868
rect 3798 3863 3804 3864
rect 3650 3862 3656 3863
rect 2022 3852 2028 3853
rect 1974 3851 1980 3852
rect 1974 3847 1975 3851
rect 1979 3847 1980 3851
rect 2022 3848 2023 3852
rect 2027 3848 2028 3852
rect 2022 3847 2028 3848
rect 2430 3852 2436 3853
rect 2430 3848 2431 3852
rect 2435 3848 2436 3852
rect 2430 3847 2436 3848
rect 2854 3852 2860 3853
rect 2854 3848 2855 3852
rect 2859 3848 2860 3852
rect 2854 3847 2860 3848
rect 3278 3852 3284 3853
rect 3278 3848 3279 3852
rect 3283 3848 3284 3852
rect 3278 3847 3284 3848
rect 3678 3852 3684 3853
rect 3678 3848 3679 3852
rect 3683 3848 3684 3852
rect 3678 3847 3684 3848
rect 3798 3851 3804 3852
rect 3798 3847 3799 3851
rect 3803 3847 3804 3851
rect 1974 3846 1980 3847
rect 3798 3846 3804 3847
rect 2522 3835 2528 3836
rect 255 3831 264 3832
rect 255 3827 256 3831
rect 263 3827 264 3831
rect 255 3826 264 3827
rect 479 3831 488 3832
rect 479 3827 480 3831
rect 487 3827 488 3831
rect 479 3826 488 3827
rect 743 3831 752 3832
rect 743 3827 744 3831
rect 751 3827 752 3831
rect 743 3826 752 3827
rect 850 3831 856 3832
rect 850 3827 851 3831
rect 855 3830 856 3831
rect 1023 3831 1029 3832
rect 1023 3830 1024 3831
rect 855 3828 1024 3830
rect 855 3827 856 3828
rect 850 3826 856 3827
rect 1023 3827 1024 3828
rect 1028 3827 1029 3831
rect 1023 3826 1029 3827
rect 1242 3831 1248 3832
rect 1242 3827 1243 3831
rect 1247 3830 1248 3831
rect 1319 3831 1325 3832
rect 1319 3830 1320 3831
rect 1247 3828 1320 3830
rect 1247 3827 1248 3828
rect 1242 3826 1248 3827
rect 1319 3827 1320 3828
rect 1324 3827 1325 3831
rect 1319 3826 1325 3827
rect 1334 3831 1340 3832
rect 1334 3827 1335 3831
rect 1339 3830 1340 3831
rect 1623 3831 1629 3832
rect 1623 3830 1624 3831
rect 1339 3828 1624 3830
rect 1339 3827 1340 3828
rect 1334 3826 1340 3827
rect 1623 3827 1624 3828
rect 1628 3827 1629 3831
rect 1623 3826 1629 3827
rect 1911 3831 1920 3832
rect 1911 3827 1912 3831
rect 1919 3827 1920 3831
rect 2522 3831 2523 3835
rect 2527 3834 2528 3835
rect 3654 3835 3660 3836
rect 3654 3834 3655 3835
rect 2527 3832 3655 3834
rect 2527 3831 2528 3832
rect 2522 3830 2528 3831
rect 3654 3831 3655 3832
rect 3659 3831 3660 3835
rect 3654 3830 3660 3831
rect 1911 3826 1920 3827
rect 110 3824 116 3825
rect 1934 3824 1940 3825
rect 110 3820 111 3824
rect 115 3820 116 3824
rect 110 3819 116 3820
rect 130 3823 136 3824
rect 130 3819 131 3823
rect 135 3819 136 3823
rect 130 3818 136 3819
rect 354 3823 360 3824
rect 354 3819 355 3823
rect 359 3819 360 3823
rect 354 3818 360 3819
rect 618 3823 624 3824
rect 618 3819 619 3823
rect 623 3819 624 3823
rect 618 3818 624 3819
rect 898 3823 904 3824
rect 898 3819 899 3823
rect 903 3819 904 3823
rect 898 3818 904 3819
rect 1194 3823 1200 3824
rect 1194 3819 1195 3823
rect 1199 3819 1200 3823
rect 1194 3818 1200 3819
rect 1498 3823 1504 3824
rect 1498 3819 1499 3823
rect 1503 3819 1504 3823
rect 1498 3818 1504 3819
rect 1786 3823 1792 3824
rect 1786 3819 1787 3823
rect 1791 3819 1792 3823
rect 1934 3820 1935 3824
rect 1939 3820 1940 3824
rect 1934 3819 1940 3820
rect 1786 3818 1792 3819
rect 158 3808 164 3809
rect 110 3807 116 3808
rect 110 3803 111 3807
rect 115 3803 116 3807
rect 158 3804 159 3808
rect 163 3804 164 3808
rect 158 3803 164 3804
rect 382 3808 388 3809
rect 382 3804 383 3808
rect 387 3804 388 3808
rect 382 3803 388 3804
rect 646 3808 652 3809
rect 646 3804 647 3808
rect 651 3804 652 3808
rect 646 3803 652 3804
rect 926 3808 932 3809
rect 926 3804 927 3808
rect 931 3804 932 3808
rect 926 3803 932 3804
rect 1222 3808 1228 3809
rect 1222 3804 1223 3808
rect 1227 3804 1228 3808
rect 1222 3803 1228 3804
rect 1526 3808 1532 3809
rect 1526 3804 1527 3808
rect 1531 3804 1532 3808
rect 1526 3803 1532 3804
rect 1814 3808 1820 3809
rect 1814 3804 1815 3808
rect 1819 3804 1820 3808
rect 1814 3803 1820 3804
rect 1934 3807 1940 3808
rect 1934 3803 1935 3807
rect 1939 3803 1940 3807
rect 110 3802 116 3803
rect 1934 3802 1940 3803
rect 1974 3793 1980 3794
rect 3798 3793 3804 3794
rect 1974 3789 1975 3793
rect 1979 3789 1980 3793
rect 1974 3788 1980 3789
rect 2022 3792 2028 3793
rect 2022 3788 2023 3792
rect 2027 3788 2028 3792
rect 2022 3787 2028 3788
rect 2174 3792 2180 3793
rect 2174 3788 2175 3792
rect 2179 3788 2180 3792
rect 2174 3787 2180 3788
rect 2350 3792 2356 3793
rect 2350 3788 2351 3792
rect 2355 3788 2356 3792
rect 2350 3787 2356 3788
rect 2534 3792 2540 3793
rect 2534 3788 2535 3792
rect 2539 3788 2540 3792
rect 2534 3787 2540 3788
rect 2718 3792 2724 3793
rect 2718 3788 2719 3792
rect 2723 3788 2724 3792
rect 2718 3787 2724 3788
rect 2894 3792 2900 3793
rect 2894 3788 2895 3792
rect 2899 3788 2900 3792
rect 2894 3787 2900 3788
rect 3070 3792 3076 3793
rect 3070 3788 3071 3792
rect 3075 3788 3076 3792
rect 3070 3787 3076 3788
rect 3246 3792 3252 3793
rect 3246 3788 3247 3792
rect 3251 3788 3252 3792
rect 3246 3787 3252 3788
rect 3422 3792 3428 3793
rect 3422 3788 3423 3792
rect 3427 3788 3428 3792
rect 3422 3787 3428 3788
rect 3606 3792 3612 3793
rect 3606 3788 3607 3792
rect 3611 3788 3612 3792
rect 3798 3789 3799 3793
rect 3803 3789 3804 3793
rect 3798 3788 3804 3789
rect 3838 3793 3844 3794
rect 5662 3793 5668 3794
rect 3838 3789 3839 3793
rect 3843 3789 3844 3793
rect 3838 3788 3844 3789
rect 4502 3792 4508 3793
rect 4502 3788 4503 3792
rect 4507 3788 4508 3792
rect 3606 3787 3612 3788
rect 4502 3787 4508 3788
rect 4638 3792 4644 3793
rect 4638 3788 4639 3792
rect 4643 3788 4644 3792
rect 4638 3787 4644 3788
rect 4774 3792 4780 3793
rect 4774 3788 4775 3792
rect 4779 3788 4780 3792
rect 4774 3787 4780 3788
rect 4910 3792 4916 3793
rect 4910 3788 4911 3792
rect 4915 3788 4916 3792
rect 4910 3787 4916 3788
rect 5046 3792 5052 3793
rect 5046 3788 5047 3792
rect 5051 3788 5052 3792
rect 5662 3789 5663 3793
rect 5667 3789 5668 3793
rect 5662 3788 5668 3789
rect 5046 3787 5052 3788
rect 1994 3777 2000 3778
rect 1974 3776 1980 3777
rect 1974 3772 1975 3776
rect 1979 3772 1980 3776
rect 1994 3773 1995 3777
rect 1999 3773 2000 3777
rect 1994 3772 2000 3773
rect 2146 3777 2152 3778
rect 2146 3773 2147 3777
rect 2151 3773 2152 3777
rect 2146 3772 2152 3773
rect 2322 3777 2328 3778
rect 2322 3773 2323 3777
rect 2327 3773 2328 3777
rect 2322 3772 2328 3773
rect 2506 3777 2512 3778
rect 2506 3773 2507 3777
rect 2511 3773 2512 3777
rect 2506 3772 2512 3773
rect 2690 3777 2696 3778
rect 2690 3773 2691 3777
rect 2695 3773 2696 3777
rect 2690 3772 2696 3773
rect 2866 3777 2872 3778
rect 2866 3773 2867 3777
rect 2871 3773 2872 3777
rect 2866 3772 2872 3773
rect 3042 3777 3048 3778
rect 3042 3773 3043 3777
rect 3047 3773 3048 3777
rect 3042 3772 3048 3773
rect 3218 3777 3224 3778
rect 3218 3773 3219 3777
rect 3223 3773 3224 3777
rect 3218 3772 3224 3773
rect 3394 3777 3400 3778
rect 3394 3773 3395 3777
rect 3399 3773 3400 3777
rect 3394 3772 3400 3773
rect 3578 3777 3584 3778
rect 4474 3777 4480 3778
rect 3578 3773 3579 3777
rect 3583 3773 3584 3777
rect 3578 3772 3584 3773
rect 3798 3776 3804 3777
rect 3798 3772 3799 3776
rect 3803 3772 3804 3776
rect 1974 3771 1980 3772
rect 3798 3771 3804 3772
rect 3838 3776 3844 3777
rect 3838 3772 3839 3776
rect 3843 3772 3844 3776
rect 4474 3773 4475 3777
rect 4479 3773 4480 3777
rect 4474 3772 4480 3773
rect 4610 3777 4616 3778
rect 4610 3773 4611 3777
rect 4615 3773 4616 3777
rect 4610 3772 4616 3773
rect 4746 3777 4752 3778
rect 4746 3773 4747 3777
rect 4751 3773 4752 3777
rect 4746 3772 4752 3773
rect 4882 3777 4888 3778
rect 4882 3773 4883 3777
rect 4887 3773 4888 3777
rect 4882 3772 4888 3773
rect 5018 3777 5024 3778
rect 5018 3773 5019 3777
rect 5023 3773 5024 3777
rect 5018 3772 5024 3773
rect 5662 3776 5668 3777
rect 5662 3772 5663 3776
rect 5667 3772 5668 3776
rect 3838 3771 3844 3772
rect 5662 3771 5668 3772
rect 2119 3767 2125 3768
rect 2119 3763 2120 3767
rect 2124 3766 2125 3767
rect 2162 3767 2168 3768
rect 2162 3766 2163 3767
rect 2124 3764 2163 3766
rect 2124 3763 2125 3764
rect 2119 3762 2125 3763
rect 2162 3763 2163 3764
rect 2167 3763 2168 3767
rect 2162 3762 2168 3763
rect 2271 3767 2277 3768
rect 2271 3763 2272 3767
rect 2276 3766 2277 3767
rect 2338 3767 2344 3768
rect 2338 3766 2339 3767
rect 2276 3764 2339 3766
rect 2276 3763 2277 3764
rect 2271 3762 2277 3763
rect 2338 3763 2339 3764
rect 2343 3763 2344 3767
rect 2338 3762 2344 3763
rect 2447 3767 2453 3768
rect 2447 3763 2448 3767
rect 2452 3766 2453 3767
rect 2522 3767 2528 3768
rect 2522 3766 2523 3767
rect 2452 3764 2523 3766
rect 2452 3763 2453 3764
rect 2447 3762 2453 3763
rect 2522 3763 2523 3764
rect 2527 3763 2528 3767
rect 2522 3762 2528 3763
rect 2631 3767 2637 3768
rect 2631 3763 2632 3767
rect 2636 3766 2637 3767
rect 2706 3767 2712 3768
rect 2706 3766 2707 3767
rect 2636 3764 2707 3766
rect 2636 3763 2637 3764
rect 2631 3762 2637 3763
rect 2706 3763 2707 3764
rect 2711 3763 2712 3767
rect 2815 3767 2821 3768
rect 2815 3766 2816 3767
rect 2706 3762 2712 3763
rect 2716 3764 2816 3766
rect 2135 3751 2141 3752
rect 2135 3747 2136 3751
rect 2140 3750 2141 3751
rect 2716 3750 2718 3764
rect 2815 3763 2816 3764
rect 2820 3763 2821 3767
rect 2815 3762 2821 3763
rect 2991 3767 2997 3768
rect 2991 3763 2992 3767
rect 2996 3766 2997 3767
rect 3058 3767 3064 3768
rect 3058 3766 3059 3767
rect 2996 3764 3059 3766
rect 2996 3763 2997 3764
rect 2991 3762 2997 3763
rect 3058 3763 3059 3764
rect 3063 3763 3064 3767
rect 3058 3762 3064 3763
rect 3167 3767 3173 3768
rect 3167 3763 3168 3767
rect 3172 3766 3173 3767
rect 3234 3767 3240 3768
rect 3234 3766 3235 3767
rect 3172 3764 3235 3766
rect 3172 3763 3173 3764
rect 3167 3762 3173 3763
rect 3234 3763 3235 3764
rect 3239 3763 3240 3767
rect 3234 3762 3240 3763
rect 3343 3767 3349 3768
rect 3343 3763 3344 3767
rect 3348 3766 3349 3767
rect 3410 3767 3416 3768
rect 3410 3766 3411 3767
rect 3348 3764 3411 3766
rect 3348 3763 3349 3764
rect 3343 3762 3349 3763
rect 3410 3763 3411 3764
rect 3415 3763 3416 3767
rect 3410 3762 3416 3763
rect 3519 3767 3525 3768
rect 3519 3763 3520 3767
rect 3524 3766 3525 3767
rect 3594 3767 3600 3768
rect 3594 3766 3595 3767
rect 3524 3764 3595 3766
rect 3524 3763 3525 3764
rect 3519 3762 3525 3763
rect 3594 3763 3595 3764
rect 3599 3763 3600 3767
rect 3594 3762 3600 3763
rect 3654 3767 3660 3768
rect 3654 3763 3655 3767
rect 3659 3766 3660 3767
rect 3703 3767 3709 3768
rect 3703 3766 3704 3767
rect 3659 3764 3704 3766
rect 3659 3763 3660 3764
rect 3654 3762 3660 3763
rect 3703 3763 3704 3764
rect 3708 3763 3709 3767
rect 3703 3762 3709 3763
rect 4599 3767 4605 3768
rect 4599 3763 4600 3767
rect 4604 3766 4605 3767
rect 4626 3767 4632 3768
rect 4626 3766 4627 3767
rect 4604 3764 4627 3766
rect 4604 3763 4605 3764
rect 4599 3762 4605 3763
rect 4626 3763 4627 3764
rect 4631 3763 4632 3767
rect 4626 3762 4632 3763
rect 4735 3767 4741 3768
rect 4735 3763 4736 3767
rect 4740 3766 4741 3767
rect 4762 3767 4768 3768
rect 4762 3766 4763 3767
rect 4740 3764 4763 3766
rect 4740 3763 4741 3764
rect 4735 3762 4741 3763
rect 4762 3763 4763 3764
rect 4767 3763 4768 3767
rect 4762 3762 4768 3763
rect 4871 3767 4877 3768
rect 4871 3763 4872 3767
rect 4876 3766 4877 3767
rect 4898 3767 4904 3768
rect 4898 3766 4899 3767
rect 4876 3764 4899 3766
rect 4876 3763 4877 3764
rect 4871 3762 4877 3763
rect 4898 3763 4899 3764
rect 4903 3763 4904 3767
rect 4898 3762 4904 3763
rect 5007 3767 5013 3768
rect 5007 3763 5008 3767
rect 5012 3766 5013 3767
rect 5034 3767 5040 3768
rect 5034 3766 5035 3767
rect 5012 3764 5035 3766
rect 5012 3763 5013 3764
rect 5007 3762 5013 3763
rect 5034 3763 5035 3764
rect 5039 3763 5040 3767
rect 5143 3767 5149 3768
rect 5143 3766 5144 3767
rect 5034 3762 5040 3763
rect 5044 3764 5144 3766
rect 4122 3759 4128 3760
rect 4122 3755 4123 3759
rect 4127 3758 4128 3759
rect 5044 3758 5046 3764
rect 5143 3763 5144 3764
rect 5148 3763 5149 3767
rect 5143 3762 5149 3763
rect 4127 3756 5046 3758
rect 4127 3755 4128 3756
rect 4122 3754 4128 3755
rect 4786 3751 4792 3752
rect 4786 3750 4787 3751
rect 2140 3748 2718 3750
rect 4616 3748 4787 3750
rect 2140 3747 2141 3748
rect 2135 3746 2141 3747
rect 110 3737 116 3738
rect 1934 3737 1940 3738
rect 110 3733 111 3737
rect 115 3733 116 3737
rect 110 3732 116 3733
rect 246 3736 252 3737
rect 246 3732 247 3736
rect 251 3732 252 3736
rect 246 3731 252 3732
rect 518 3736 524 3737
rect 518 3732 519 3736
rect 523 3732 524 3736
rect 518 3731 524 3732
rect 790 3736 796 3737
rect 790 3732 791 3736
rect 795 3732 796 3736
rect 790 3731 796 3732
rect 1062 3736 1068 3737
rect 1062 3732 1063 3736
rect 1067 3732 1068 3736
rect 1062 3731 1068 3732
rect 1342 3736 1348 3737
rect 1342 3732 1343 3736
rect 1347 3732 1348 3736
rect 1934 3733 1935 3737
rect 1939 3733 1940 3737
rect 1934 3732 1940 3733
rect 2082 3735 2088 3736
rect 1342 3731 1348 3732
rect 2082 3731 2083 3735
rect 2087 3731 2088 3735
rect 2082 3730 2088 3731
rect 2162 3735 2168 3736
rect 2162 3731 2163 3735
rect 2167 3731 2168 3735
rect 2162 3730 2168 3731
rect 2338 3735 2344 3736
rect 2338 3731 2339 3735
rect 2343 3731 2344 3735
rect 2338 3730 2344 3731
rect 2522 3735 2528 3736
rect 2522 3731 2523 3735
rect 2527 3731 2528 3735
rect 2522 3730 2528 3731
rect 2706 3735 2712 3736
rect 2706 3731 2707 3735
rect 2711 3731 2712 3735
rect 3058 3735 3064 3736
rect 2957 3732 3014 3734
rect 2706 3730 2712 3731
rect 218 3721 224 3722
rect 110 3720 116 3721
rect 110 3716 111 3720
rect 115 3716 116 3720
rect 218 3717 219 3721
rect 223 3717 224 3721
rect 218 3716 224 3717
rect 490 3721 496 3722
rect 490 3717 491 3721
rect 495 3717 496 3721
rect 490 3716 496 3717
rect 762 3721 768 3722
rect 762 3717 763 3721
rect 767 3717 768 3721
rect 762 3716 768 3717
rect 1034 3721 1040 3722
rect 1034 3717 1035 3721
rect 1039 3717 1040 3721
rect 1034 3716 1040 3717
rect 1314 3721 1320 3722
rect 1314 3717 1315 3721
rect 1319 3717 1320 3721
rect 1314 3716 1320 3717
rect 1934 3720 1940 3721
rect 1934 3716 1935 3720
rect 1939 3716 1940 3720
rect 3012 3718 3014 3732
rect 3058 3731 3059 3735
rect 3063 3731 3064 3735
rect 3058 3730 3064 3731
rect 3234 3735 3240 3736
rect 3234 3731 3235 3735
rect 3239 3731 3240 3735
rect 3234 3730 3240 3731
rect 3410 3735 3416 3736
rect 3410 3731 3411 3735
rect 3415 3731 3416 3735
rect 3410 3730 3416 3731
rect 3594 3735 3600 3736
rect 3594 3731 3595 3735
rect 3599 3731 3600 3735
rect 4616 3734 4618 3748
rect 4786 3747 4787 3748
rect 4791 3747 4792 3751
rect 4786 3746 4792 3747
rect 4565 3732 4618 3734
rect 4626 3735 4632 3736
rect 3594 3730 3600 3731
rect 4626 3731 4627 3735
rect 4631 3731 4632 3735
rect 4626 3730 4632 3731
rect 4762 3735 4768 3736
rect 4762 3731 4763 3735
rect 4767 3731 4768 3735
rect 4762 3730 4768 3731
rect 4898 3735 4904 3736
rect 4898 3731 4899 3735
rect 4903 3731 4904 3735
rect 4898 3730 4904 3731
rect 5034 3735 5040 3736
rect 5034 3731 5035 3735
rect 5039 3731 5040 3735
rect 5034 3730 5040 3731
rect 3422 3719 3428 3720
rect 3422 3718 3423 3719
rect 3012 3716 3423 3718
rect 110 3715 116 3716
rect 1934 3715 1940 3716
rect 3422 3715 3423 3716
rect 3427 3715 3428 3719
rect 3422 3714 3428 3715
rect 343 3711 349 3712
rect 343 3707 344 3711
rect 348 3710 349 3711
rect 506 3711 512 3712
rect 506 3710 507 3711
rect 348 3708 507 3710
rect 348 3707 349 3708
rect 343 3706 349 3707
rect 506 3707 507 3708
rect 511 3707 512 3711
rect 506 3706 512 3707
rect 594 3711 600 3712
rect 594 3707 595 3711
rect 599 3710 600 3711
rect 615 3711 621 3712
rect 615 3710 616 3711
rect 599 3708 616 3710
rect 599 3707 600 3708
rect 594 3706 600 3707
rect 615 3707 616 3708
rect 620 3707 621 3711
rect 887 3711 893 3712
rect 887 3710 888 3711
rect 615 3706 621 3707
rect 752 3708 888 3710
rect 306 3703 312 3704
rect 306 3699 307 3703
rect 311 3702 312 3703
rect 752 3702 754 3708
rect 887 3707 888 3708
rect 892 3707 893 3711
rect 887 3706 893 3707
rect 1159 3711 1165 3712
rect 1159 3707 1160 3711
rect 1164 3710 1165 3711
rect 1330 3711 1336 3712
rect 1330 3710 1331 3711
rect 1164 3708 1331 3710
rect 1164 3707 1165 3708
rect 1159 3706 1165 3707
rect 1330 3707 1331 3708
rect 1335 3707 1336 3711
rect 1330 3706 1336 3707
rect 1439 3711 1445 3712
rect 1439 3707 1440 3711
rect 1444 3710 1445 3711
rect 1447 3711 1453 3712
rect 1447 3710 1448 3711
rect 1444 3708 1448 3710
rect 1444 3707 1445 3708
rect 1439 3706 1445 3707
rect 1447 3707 1448 3708
rect 1452 3707 1453 3711
rect 1447 3706 1453 3707
rect 311 3700 754 3702
rect 311 3699 312 3700
rect 306 3698 312 3699
rect 306 3679 312 3680
rect 306 3675 307 3679
rect 311 3675 312 3679
rect 306 3674 312 3675
rect 506 3679 512 3680
rect 506 3675 507 3679
rect 511 3675 512 3679
rect 506 3674 512 3675
rect 850 3679 856 3680
rect 850 3675 851 3679
rect 855 3675 856 3679
rect 1202 3679 1208 3680
rect 1202 3678 1203 3679
rect 1125 3676 1203 3678
rect 850 3674 856 3675
rect 1202 3675 1203 3676
rect 1207 3675 1208 3679
rect 1202 3674 1208 3675
rect 1330 3679 1336 3680
rect 1330 3675 1331 3679
rect 1335 3675 1336 3679
rect 2135 3679 2141 3680
rect 2135 3678 2136 3679
rect 2101 3676 2136 3678
rect 1330 3674 1336 3675
rect 2135 3675 2136 3676
rect 2140 3675 2141 3679
rect 2135 3674 2141 3675
rect 2143 3679 2149 3680
rect 2143 3675 2144 3679
rect 2148 3678 2149 3679
rect 2274 3679 2280 3680
rect 2148 3676 2165 3678
rect 2148 3675 2149 3676
rect 2143 3674 2149 3675
rect 2274 3675 2275 3679
rect 2279 3678 2280 3679
rect 2418 3679 2424 3680
rect 2279 3676 2309 3678
rect 2279 3675 2280 3676
rect 2274 3674 2280 3675
rect 2418 3675 2419 3679
rect 2423 3678 2424 3679
rect 2562 3679 2568 3680
rect 2423 3676 2453 3678
rect 2423 3675 2424 3676
rect 2418 3674 2424 3675
rect 2562 3675 2563 3679
rect 2567 3678 2568 3679
rect 2850 3679 2856 3680
rect 2567 3676 2597 3678
rect 2567 3675 2568 3676
rect 2562 3674 2568 3675
rect 2850 3675 2851 3679
rect 2855 3678 2856 3679
rect 2994 3679 3000 3680
rect 2855 3676 2885 3678
rect 2855 3675 2856 3676
rect 2850 3674 2856 3675
rect 2994 3675 2995 3679
rect 2999 3678 3000 3679
rect 3151 3679 3157 3680
rect 2999 3676 3029 3678
rect 2999 3675 3000 3676
rect 2994 3674 3000 3675
rect 3151 3675 3152 3679
rect 3156 3678 3157 3679
rect 3282 3679 3288 3680
rect 3156 3676 3173 3678
rect 3156 3675 3157 3676
rect 3151 3674 3157 3675
rect 3282 3675 3283 3679
rect 3287 3678 3288 3679
rect 3287 3676 3317 3678
rect 3287 3675 3288 3676
rect 3282 3674 3288 3675
rect 2808 3662 2810 3673
rect 4122 3667 4128 3668
rect 4122 3666 4123 3667
rect 4109 3664 4123 3666
rect 2954 3663 2960 3664
rect 2954 3662 2955 3663
rect 2808 3660 2955 3662
rect 2954 3659 2955 3660
rect 2959 3659 2960 3663
rect 4122 3663 4123 3664
rect 4127 3663 4128 3667
rect 4122 3662 4128 3663
rect 4146 3667 4152 3668
rect 4146 3663 4147 3667
rect 4151 3666 4152 3667
rect 4282 3667 4288 3668
rect 4151 3664 4173 3666
rect 4151 3663 4152 3664
rect 4146 3662 4152 3663
rect 4282 3663 4283 3667
rect 4287 3666 4288 3667
rect 4418 3667 4424 3668
rect 4287 3664 4309 3666
rect 4287 3663 4288 3664
rect 4282 3662 4288 3663
rect 4418 3663 4419 3667
rect 4423 3666 4424 3667
rect 4554 3667 4560 3668
rect 4423 3664 4445 3666
rect 4423 3663 4424 3664
rect 4418 3662 4424 3663
rect 4554 3663 4555 3667
rect 4559 3666 4560 3667
rect 4690 3667 4696 3668
rect 4559 3664 4581 3666
rect 4559 3663 4560 3664
rect 4554 3662 4560 3663
rect 4690 3663 4691 3667
rect 4695 3666 4696 3667
rect 4826 3667 4832 3668
rect 4695 3664 4717 3666
rect 4695 3663 4696 3664
rect 4690 3662 4696 3663
rect 4826 3663 4827 3667
rect 4831 3666 4832 3667
rect 4967 3667 4973 3668
rect 4831 3664 4853 3666
rect 4831 3663 4832 3664
rect 4826 3662 4832 3663
rect 4967 3663 4968 3667
rect 4972 3666 4973 3667
rect 5103 3667 5109 3668
rect 4972 3664 4989 3666
rect 4972 3663 4973 3664
rect 4967 3662 4973 3663
rect 5103 3663 5104 3667
rect 5108 3666 5109 3667
rect 5239 3667 5245 3668
rect 5108 3664 5125 3666
rect 5108 3663 5109 3664
rect 5103 3662 5109 3663
rect 5239 3663 5240 3667
rect 5244 3666 5245 3667
rect 5375 3667 5381 3668
rect 5244 3664 5261 3666
rect 5244 3663 5245 3664
rect 5239 3662 5245 3663
rect 5375 3663 5376 3667
rect 5380 3666 5381 3667
rect 5511 3667 5517 3668
rect 5380 3664 5397 3666
rect 5380 3663 5381 3664
rect 5375 3662 5381 3663
rect 5511 3663 5512 3667
rect 5516 3666 5517 3667
rect 5516 3664 5533 3666
rect 5516 3663 5517 3664
rect 5511 3662 5517 3663
rect 2954 3658 2960 3659
rect 2135 3643 2141 3644
rect 2135 3639 2136 3643
rect 2140 3642 2141 3643
rect 2143 3643 2149 3644
rect 2143 3642 2144 3643
rect 2140 3640 2144 3642
rect 2140 3639 2141 3640
rect 2135 3638 2141 3639
rect 2143 3639 2144 3640
rect 2148 3639 2149 3643
rect 2143 3638 2149 3639
rect 2271 3643 2280 3644
rect 2271 3639 2272 3643
rect 2279 3639 2280 3643
rect 2271 3638 2280 3639
rect 2415 3643 2424 3644
rect 2415 3639 2416 3643
rect 2423 3639 2424 3643
rect 2415 3638 2424 3639
rect 2559 3643 2568 3644
rect 2559 3639 2560 3643
rect 2567 3639 2568 3643
rect 2559 3638 2568 3639
rect 2598 3643 2604 3644
rect 2598 3639 2599 3643
rect 2603 3642 2604 3643
rect 2703 3643 2709 3644
rect 2703 3642 2704 3643
rect 2603 3640 2704 3642
rect 2603 3639 2604 3640
rect 2598 3638 2604 3639
rect 2703 3639 2704 3640
rect 2708 3639 2709 3643
rect 2703 3638 2709 3639
rect 2847 3643 2856 3644
rect 2847 3639 2848 3643
rect 2855 3639 2856 3643
rect 2847 3638 2856 3639
rect 2991 3643 3000 3644
rect 2991 3639 2992 3643
rect 2999 3639 3000 3643
rect 2991 3638 3000 3639
rect 3135 3643 3141 3644
rect 3135 3639 3136 3643
rect 3140 3642 3141 3643
rect 3151 3643 3157 3644
rect 3151 3642 3152 3643
rect 3140 3640 3152 3642
rect 3140 3639 3141 3640
rect 3135 3638 3141 3639
rect 3151 3639 3152 3640
rect 3156 3639 3157 3643
rect 3151 3638 3157 3639
rect 3279 3643 3288 3644
rect 3279 3639 3280 3643
rect 3287 3639 3288 3643
rect 3279 3638 3288 3639
rect 3422 3643 3429 3644
rect 3422 3639 3423 3643
rect 3428 3639 3429 3643
rect 3422 3638 3429 3639
rect 1974 3636 1980 3637
rect 3798 3636 3804 3637
rect 1974 3632 1975 3636
rect 1979 3632 1980 3636
rect 1974 3631 1980 3632
rect 2010 3635 2016 3636
rect 2010 3631 2011 3635
rect 2015 3631 2016 3635
rect 2010 3630 2016 3631
rect 2146 3635 2152 3636
rect 2146 3631 2147 3635
rect 2151 3631 2152 3635
rect 2146 3630 2152 3631
rect 2290 3635 2296 3636
rect 2290 3631 2291 3635
rect 2295 3631 2296 3635
rect 2290 3630 2296 3631
rect 2434 3635 2440 3636
rect 2434 3631 2435 3635
rect 2439 3631 2440 3635
rect 2434 3630 2440 3631
rect 2578 3635 2584 3636
rect 2578 3631 2579 3635
rect 2583 3631 2584 3635
rect 2578 3630 2584 3631
rect 2722 3635 2728 3636
rect 2722 3631 2723 3635
rect 2727 3631 2728 3635
rect 2722 3630 2728 3631
rect 2866 3635 2872 3636
rect 2866 3631 2867 3635
rect 2871 3631 2872 3635
rect 2866 3630 2872 3631
rect 3010 3635 3016 3636
rect 3010 3631 3011 3635
rect 3015 3631 3016 3635
rect 3010 3630 3016 3631
rect 3154 3635 3160 3636
rect 3154 3631 3155 3635
rect 3159 3631 3160 3635
rect 3154 3630 3160 3631
rect 3298 3635 3304 3636
rect 3298 3631 3299 3635
rect 3303 3631 3304 3635
rect 3798 3632 3799 3636
rect 3803 3632 3804 3636
rect 3798 3631 3804 3632
rect 4143 3631 4152 3632
rect 3298 3630 3304 3631
rect 4143 3627 4144 3631
rect 4151 3627 4152 3631
rect 4143 3626 4152 3627
rect 4279 3631 4288 3632
rect 4279 3627 4280 3631
rect 4287 3627 4288 3631
rect 4279 3626 4288 3627
rect 4415 3631 4424 3632
rect 4415 3627 4416 3631
rect 4423 3627 4424 3631
rect 4415 3626 4424 3627
rect 4551 3631 4560 3632
rect 4551 3627 4552 3631
rect 4559 3627 4560 3631
rect 4551 3626 4560 3627
rect 4687 3631 4696 3632
rect 4687 3627 4688 3631
rect 4695 3627 4696 3631
rect 4687 3626 4696 3627
rect 4823 3631 4832 3632
rect 4823 3627 4824 3631
rect 4831 3627 4832 3631
rect 4823 3626 4832 3627
rect 4959 3631 4965 3632
rect 4959 3627 4960 3631
rect 4964 3630 4965 3631
rect 4967 3631 4973 3632
rect 4967 3630 4968 3631
rect 4964 3628 4968 3630
rect 4964 3627 4965 3628
rect 4959 3626 4965 3627
rect 4967 3627 4968 3628
rect 4972 3627 4973 3631
rect 4967 3626 4973 3627
rect 5095 3631 5101 3632
rect 5095 3627 5096 3631
rect 5100 3630 5101 3631
rect 5103 3631 5109 3632
rect 5103 3630 5104 3631
rect 5100 3628 5104 3630
rect 5100 3627 5101 3628
rect 5095 3626 5101 3627
rect 5103 3627 5104 3628
rect 5108 3627 5109 3631
rect 5103 3626 5109 3627
rect 5231 3631 5237 3632
rect 5231 3627 5232 3631
rect 5236 3630 5237 3631
rect 5239 3631 5245 3632
rect 5239 3630 5240 3631
rect 5236 3628 5240 3630
rect 5236 3627 5237 3628
rect 5231 3626 5237 3627
rect 5239 3627 5240 3628
rect 5244 3627 5245 3631
rect 5239 3626 5245 3627
rect 5367 3631 5373 3632
rect 5367 3627 5368 3631
rect 5372 3630 5373 3631
rect 5375 3631 5381 3632
rect 5375 3630 5376 3631
rect 5372 3628 5376 3630
rect 5372 3627 5373 3628
rect 5367 3626 5373 3627
rect 5375 3627 5376 3628
rect 5380 3627 5381 3631
rect 5375 3626 5381 3627
rect 5503 3631 5509 3632
rect 5503 3627 5504 3631
rect 5508 3630 5509 3631
rect 5511 3631 5517 3632
rect 5511 3630 5512 3631
rect 5508 3628 5512 3630
rect 5508 3627 5509 3628
rect 5503 3626 5509 3627
rect 5511 3627 5512 3628
rect 5516 3627 5517 3631
rect 5511 3626 5517 3627
rect 5550 3631 5556 3632
rect 5550 3627 5551 3631
rect 5555 3630 5556 3631
rect 5639 3631 5645 3632
rect 5639 3630 5640 3631
rect 5555 3628 5640 3630
rect 5555 3627 5556 3628
rect 5550 3626 5556 3627
rect 5639 3627 5640 3628
rect 5644 3627 5645 3631
rect 5639 3626 5645 3627
rect 3838 3624 3844 3625
rect 5662 3624 5668 3625
rect 2038 3620 2044 3621
rect 1974 3619 1980 3620
rect 594 3615 600 3616
rect 594 3614 595 3615
rect 581 3612 595 3614
rect 594 3611 595 3612
rect 599 3611 600 3615
rect 594 3610 600 3611
rect 631 3615 637 3616
rect 631 3611 632 3615
rect 636 3614 637 3615
rect 762 3615 768 3616
rect 636 3612 653 3614
rect 636 3611 637 3612
rect 631 3610 637 3611
rect 762 3611 763 3615
rect 767 3614 768 3615
rect 1050 3615 1056 3616
rect 767 3612 797 3614
rect 767 3611 768 3612
rect 762 3610 768 3611
rect 1010 3611 1016 3612
rect 1010 3607 1011 3611
rect 1015 3607 1016 3611
rect 1050 3611 1051 3615
rect 1055 3614 1056 3615
rect 1194 3615 1200 3616
rect 1055 3612 1085 3614
rect 1055 3611 1056 3612
rect 1050 3610 1056 3611
rect 1194 3611 1195 3615
rect 1199 3614 1200 3615
rect 1974 3615 1975 3619
rect 1979 3615 1980 3619
rect 2038 3616 2039 3620
rect 2043 3616 2044 3620
rect 2038 3615 2044 3616
rect 2174 3620 2180 3621
rect 2174 3616 2175 3620
rect 2179 3616 2180 3620
rect 2174 3615 2180 3616
rect 2318 3620 2324 3621
rect 2318 3616 2319 3620
rect 2323 3616 2324 3620
rect 2318 3615 2324 3616
rect 2462 3620 2468 3621
rect 2462 3616 2463 3620
rect 2467 3616 2468 3620
rect 2462 3615 2468 3616
rect 2606 3620 2612 3621
rect 2606 3616 2607 3620
rect 2611 3616 2612 3620
rect 2606 3615 2612 3616
rect 2750 3620 2756 3621
rect 2750 3616 2751 3620
rect 2755 3616 2756 3620
rect 2750 3615 2756 3616
rect 2894 3620 2900 3621
rect 2894 3616 2895 3620
rect 2899 3616 2900 3620
rect 2894 3615 2900 3616
rect 3038 3620 3044 3621
rect 3038 3616 3039 3620
rect 3043 3616 3044 3620
rect 3038 3615 3044 3616
rect 3182 3620 3188 3621
rect 3182 3616 3183 3620
rect 3187 3616 3188 3620
rect 3182 3615 3188 3616
rect 3326 3620 3332 3621
rect 3838 3620 3839 3624
rect 3843 3620 3844 3624
rect 3326 3616 3327 3620
rect 3331 3616 3332 3620
rect 3326 3615 3332 3616
rect 3798 3619 3804 3620
rect 3838 3619 3844 3620
rect 4018 3623 4024 3624
rect 4018 3619 4019 3623
rect 4023 3619 4024 3623
rect 3798 3615 3799 3619
rect 3803 3615 3804 3619
rect 4018 3618 4024 3619
rect 4154 3623 4160 3624
rect 4154 3619 4155 3623
rect 4159 3619 4160 3623
rect 4154 3618 4160 3619
rect 4290 3623 4296 3624
rect 4290 3619 4291 3623
rect 4295 3619 4296 3623
rect 4290 3618 4296 3619
rect 4426 3623 4432 3624
rect 4426 3619 4427 3623
rect 4431 3619 4432 3623
rect 4426 3618 4432 3619
rect 4562 3623 4568 3624
rect 4562 3619 4563 3623
rect 4567 3619 4568 3623
rect 4562 3618 4568 3619
rect 4698 3623 4704 3624
rect 4698 3619 4699 3623
rect 4703 3619 4704 3623
rect 4698 3618 4704 3619
rect 4834 3623 4840 3624
rect 4834 3619 4835 3623
rect 4839 3619 4840 3623
rect 4834 3618 4840 3619
rect 4970 3623 4976 3624
rect 4970 3619 4971 3623
rect 4975 3619 4976 3623
rect 4970 3618 4976 3619
rect 5106 3623 5112 3624
rect 5106 3619 5107 3623
rect 5111 3619 5112 3623
rect 5106 3618 5112 3619
rect 5242 3623 5248 3624
rect 5242 3619 5243 3623
rect 5247 3619 5248 3623
rect 5242 3618 5248 3619
rect 5378 3623 5384 3624
rect 5378 3619 5379 3623
rect 5383 3619 5384 3623
rect 5378 3618 5384 3619
rect 5514 3623 5520 3624
rect 5514 3619 5515 3623
rect 5519 3619 5520 3623
rect 5662 3620 5663 3624
rect 5667 3620 5668 3624
rect 5662 3619 5668 3620
rect 5514 3618 5520 3619
rect 1974 3614 1980 3615
rect 3798 3614 3804 3615
rect 1199 3612 1229 3614
rect 1199 3611 1200 3612
rect 1194 3610 1200 3611
rect 4046 3608 4052 3609
rect 1010 3606 1016 3607
rect 3838 3607 3844 3608
rect 3838 3603 3839 3607
rect 3843 3603 3844 3607
rect 4046 3604 4047 3608
rect 4051 3604 4052 3608
rect 4046 3603 4052 3604
rect 4182 3608 4188 3609
rect 4182 3604 4183 3608
rect 4187 3604 4188 3608
rect 4182 3603 4188 3604
rect 4318 3608 4324 3609
rect 4318 3604 4319 3608
rect 4323 3604 4324 3608
rect 4318 3603 4324 3604
rect 4454 3608 4460 3609
rect 4454 3604 4455 3608
rect 4459 3604 4460 3608
rect 4454 3603 4460 3604
rect 4590 3608 4596 3609
rect 4590 3604 4591 3608
rect 4595 3604 4596 3608
rect 4590 3603 4596 3604
rect 4726 3608 4732 3609
rect 4726 3604 4727 3608
rect 4731 3604 4732 3608
rect 4726 3603 4732 3604
rect 4862 3608 4868 3609
rect 4862 3604 4863 3608
rect 4867 3604 4868 3608
rect 4862 3603 4868 3604
rect 4998 3608 5004 3609
rect 4998 3604 4999 3608
rect 5003 3604 5004 3608
rect 4998 3603 5004 3604
rect 5134 3608 5140 3609
rect 5134 3604 5135 3608
rect 5139 3604 5140 3608
rect 5134 3603 5140 3604
rect 5270 3608 5276 3609
rect 5270 3604 5271 3608
rect 5275 3604 5276 3608
rect 5270 3603 5276 3604
rect 5406 3608 5412 3609
rect 5406 3604 5407 3608
rect 5411 3604 5412 3608
rect 5406 3603 5412 3604
rect 5542 3608 5548 3609
rect 5542 3604 5543 3608
rect 5547 3604 5548 3608
rect 5542 3603 5548 3604
rect 5662 3607 5668 3608
rect 5662 3603 5663 3607
rect 5667 3603 5668 3607
rect 3838 3602 3844 3603
rect 5662 3602 5668 3603
rect 615 3579 621 3580
rect 615 3575 616 3579
rect 620 3578 621 3579
rect 631 3579 637 3580
rect 631 3578 632 3579
rect 620 3576 632 3578
rect 620 3575 621 3576
rect 615 3574 621 3575
rect 631 3575 632 3576
rect 636 3575 637 3579
rect 631 3574 637 3575
rect 759 3579 768 3580
rect 759 3575 760 3579
rect 767 3575 768 3579
rect 759 3574 768 3575
rect 898 3579 909 3580
rect 898 3575 899 3579
rect 903 3575 904 3579
rect 908 3575 909 3579
rect 898 3574 909 3575
rect 1047 3579 1056 3580
rect 1047 3575 1048 3579
rect 1055 3575 1056 3579
rect 1047 3574 1056 3575
rect 1191 3579 1200 3580
rect 1191 3575 1192 3579
rect 1199 3575 1200 3579
rect 1191 3574 1200 3575
rect 1202 3579 1208 3580
rect 1202 3575 1203 3579
rect 1207 3578 1208 3579
rect 1335 3579 1341 3580
rect 1335 3578 1336 3579
rect 1207 3576 1336 3578
rect 1207 3575 1208 3576
rect 1202 3574 1208 3575
rect 1335 3575 1336 3576
rect 1340 3575 1341 3579
rect 1335 3574 1341 3575
rect 110 3572 116 3573
rect 1934 3572 1940 3573
rect 110 3568 111 3572
rect 115 3568 116 3572
rect 110 3567 116 3568
rect 490 3571 496 3572
rect 490 3567 491 3571
rect 495 3567 496 3571
rect 490 3566 496 3567
rect 634 3571 640 3572
rect 634 3567 635 3571
rect 639 3567 640 3571
rect 634 3566 640 3567
rect 778 3571 784 3572
rect 778 3567 779 3571
rect 783 3567 784 3571
rect 778 3566 784 3567
rect 922 3571 928 3572
rect 922 3567 923 3571
rect 927 3567 928 3571
rect 922 3566 928 3567
rect 1066 3571 1072 3572
rect 1066 3567 1067 3571
rect 1071 3567 1072 3571
rect 1066 3566 1072 3567
rect 1210 3571 1216 3572
rect 1210 3567 1211 3571
rect 1215 3567 1216 3571
rect 1934 3568 1935 3572
rect 1939 3568 1940 3572
rect 1934 3567 1940 3568
rect 1210 3566 1216 3567
rect 518 3556 524 3557
rect 110 3555 116 3556
rect 110 3551 111 3555
rect 115 3551 116 3555
rect 518 3552 519 3556
rect 523 3552 524 3556
rect 518 3551 524 3552
rect 662 3556 668 3557
rect 662 3552 663 3556
rect 667 3552 668 3556
rect 662 3551 668 3552
rect 806 3556 812 3557
rect 806 3552 807 3556
rect 811 3552 812 3556
rect 806 3551 812 3552
rect 950 3556 956 3557
rect 950 3552 951 3556
rect 955 3552 956 3556
rect 950 3551 956 3552
rect 1094 3556 1100 3557
rect 1094 3552 1095 3556
rect 1099 3552 1100 3556
rect 1094 3551 1100 3552
rect 1238 3556 1244 3557
rect 1238 3552 1239 3556
rect 1243 3552 1244 3556
rect 1238 3551 1244 3552
rect 1934 3555 1940 3556
rect 1934 3551 1935 3555
rect 1939 3551 1940 3555
rect 110 3550 116 3551
rect 1934 3550 1940 3551
rect 1974 3553 1980 3554
rect 3798 3553 3804 3554
rect 1974 3549 1975 3553
rect 1979 3549 1980 3553
rect 1974 3548 1980 3549
rect 2238 3552 2244 3553
rect 2238 3548 2239 3552
rect 2243 3548 2244 3552
rect 2238 3547 2244 3548
rect 2374 3552 2380 3553
rect 2374 3548 2375 3552
rect 2379 3548 2380 3552
rect 2374 3547 2380 3548
rect 2510 3552 2516 3553
rect 2510 3548 2511 3552
rect 2515 3548 2516 3552
rect 2510 3547 2516 3548
rect 2646 3552 2652 3553
rect 2646 3548 2647 3552
rect 2651 3548 2652 3552
rect 2646 3547 2652 3548
rect 2782 3552 2788 3553
rect 2782 3548 2783 3552
rect 2787 3548 2788 3552
rect 2782 3547 2788 3548
rect 2918 3552 2924 3553
rect 2918 3548 2919 3552
rect 2923 3548 2924 3552
rect 2918 3547 2924 3548
rect 3054 3552 3060 3553
rect 3054 3548 3055 3552
rect 3059 3548 3060 3552
rect 3054 3547 3060 3548
rect 3190 3552 3196 3553
rect 3190 3548 3191 3552
rect 3195 3548 3196 3552
rect 3190 3547 3196 3548
rect 3326 3552 3332 3553
rect 3326 3548 3327 3552
rect 3331 3548 3332 3552
rect 3326 3547 3332 3548
rect 3462 3552 3468 3553
rect 3462 3548 3463 3552
rect 3467 3548 3468 3552
rect 3798 3549 3799 3553
rect 3803 3549 3804 3553
rect 3798 3548 3804 3549
rect 3462 3547 3468 3548
rect 2210 3537 2216 3538
rect 1974 3536 1980 3537
rect 1974 3532 1975 3536
rect 1979 3532 1980 3536
rect 2210 3533 2211 3537
rect 2215 3533 2216 3537
rect 2210 3532 2216 3533
rect 2346 3537 2352 3538
rect 2346 3533 2347 3537
rect 2351 3533 2352 3537
rect 2346 3532 2352 3533
rect 2482 3537 2488 3538
rect 2482 3533 2483 3537
rect 2487 3533 2488 3537
rect 2482 3532 2488 3533
rect 2618 3537 2624 3538
rect 2618 3533 2619 3537
rect 2623 3533 2624 3537
rect 2618 3532 2624 3533
rect 2754 3537 2760 3538
rect 2754 3533 2755 3537
rect 2759 3533 2760 3537
rect 2754 3532 2760 3533
rect 2890 3537 2896 3538
rect 2890 3533 2891 3537
rect 2895 3533 2896 3537
rect 2890 3532 2896 3533
rect 3026 3537 3032 3538
rect 3026 3533 3027 3537
rect 3031 3533 3032 3537
rect 3026 3532 3032 3533
rect 3162 3537 3168 3538
rect 3162 3533 3163 3537
rect 3167 3533 3168 3537
rect 3162 3532 3168 3533
rect 3298 3537 3304 3538
rect 3298 3533 3299 3537
rect 3303 3533 3304 3537
rect 3298 3532 3304 3533
rect 3434 3537 3440 3538
rect 3434 3533 3435 3537
rect 3439 3533 3440 3537
rect 3434 3532 3440 3533
rect 3798 3536 3804 3537
rect 3798 3532 3799 3536
rect 3803 3532 3804 3536
rect 1974 3531 1980 3532
rect 3798 3531 3804 3532
rect 2335 3527 2341 3528
rect 2335 3523 2336 3527
rect 2340 3526 2341 3527
rect 2362 3527 2368 3528
rect 2362 3526 2363 3527
rect 2340 3524 2363 3526
rect 2340 3523 2341 3524
rect 2335 3522 2341 3523
rect 2362 3523 2363 3524
rect 2367 3523 2368 3527
rect 2362 3522 2368 3523
rect 2471 3527 2477 3528
rect 2471 3523 2472 3527
rect 2476 3526 2477 3527
rect 2498 3527 2504 3528
rect 2498 3526 2499 3527
rect 2476 3524 2499 3526
rect 2476 3523 2477 3524
rect 2471 3522 2477 3523
rect 2498 3523 2499 3524
rect 2503 3523 2504 3527
rect 2498 3522 2504 3523
rect 2607 3527 2613 3528
rect 2607 3523 2608 3527
rect 2612 3526 2613 3527
rect 2634 3527 2640 3528
rect 2634 3526 2635 3527
rect 2612 3524 2635 3526
rect 2612 3523 2613 3524
rect 2607 3522 2613 3523
rect 2634 3523 2635 3524
rect 2639 3523 2640 3527
rect 2634 3522 2640 3523
rect 2743 3527 2749 3528
rect 2743 3523 2744 3527
rect 2748 3526 2749 3527
rect 2770 3527 2776 3528
rect 2770 3526 2771 3527
rect 2748 3524 2771 3526
rect 2748 3523 2749 3524
rect 2743 3522 2749 3523
rect 2770 3523 2771 3524
rect 2775 3523 2776 3527
rect 2770 3522 2776 3523
rect 2802 3527 2808 3528
rect 2802 3523 2803 3527
rect 2807 3526 2808 3527
rect 2879 3527 2885 3528
rect 2879 3526 2880 3527
rect 2807 3524 2880 3526
rect 2807 3523 2808 3524
rect 2802 3522 2808 3523
rect 2879 3523 2880 3524
rect 2884 3523 2885 3527
rect 2879 3522 2885 3523
rect 2954 3527 2960 3528
rect 2954 3523 2955 3527
rect 2959 3526 2960 3527
rect 3015 3527 3021 3528
rect 3015 3526 3016 3527
rect 2959 3524 3016 3526
rect 2959 3523 2960 3524
rect 2954 3522 2960 3523
rect 3015 3523 3016 3524
rect 3020 3523 3021 3527
rect 3015 3522 3021 3523
rect 3023 3527 3029 3528
rect 3023 3523 3024 3527
rect 3028 3526 3029 3527
rect 3151 3527 3157 3528
rect 3151 3526 3152 3527
rect 3028 3524 3152 3526
rect 3028 3523 3029 3524
rect 3023 3522 3029 3523
rect 3151 3523 3152 3524
rect 3156 3523 3157 3527
rect 3151 3522 3157 3523
rect 3170 3527 3176 3528
rect 3170 3523 3171 3527
rect 3175 3526 3176 3527
rect 3287 3527 3293 3528
rect 3287 3526 3288 3527
rect 3175 3524 3288 3526
rect 3175 3523 3176 3524
rect 3170 3522 3176 3523
rect 3287 3523 3288 3524
rect 3292 3523 3293 3527
rect 3287 3522 3293 3523
rect 3423 3527 3429 3528
rect 3423 3523 3424 3527
rect 3428 3526 3429 3527
rect 3450 3527 3456 3528
rect 3450 3526 3451 3527
rect 3428 3524 3451 3526
rect 3428 3523 3429 3524
rect 3423 3522 3429 3523
rect 3450 3523 3451 3524
rect 3455 3523 3456 3527
rect 3559 3527 3565 3528
rect 3559 3526 3560 3527
rect 3450 3522 3456 3523
rect 3460 3524 3560 3526
rect 3250 3519 3256 3520
rect 3250 3515 3251 3519
rect 3255 3518 3256 3519
rect 3460 3518 3462 3524
rect 3559 3523 3560 3524
rect 3564 3523 3565 3527
rect 3559 3522 3565 3523
rect 3255 3516 3462 3518
rect 3255 3515 3256 3516
rect 3250 3514 3256 3515
rect 2598 3511 2604 3512
rect 2598 3510 2599 3511
rect 2300 3508 2599 3510
rect 2300 3493 2302 3508
rect 2598 3507 2599 3508
rect 2603 3507 2604 3511
rect 2598 3506 2604 3507
rect 3838 3501 3844 3502
rect 5662 3501 5668 3502
rect 3838 3497 3839 3501
rect 3843 3497 3844 3501
rect 3838 3496 3844 3497
rect 5406 3500 5412 3501
rect 5406 3496 5407 3500
rect 5411 3496 5412 3500
rect 2362 3495 2368 3496
rect 2362 3491 2363 3495
rect 2367 3491 2368 3495
rect 2362 3490 2368 3491
rect 2498 3495 2504 3496
rect 2498 3491 2499 3495
rect 2503 3491 2504 3495
rect 2498 3490 2504 3491
rect 2634 3495 2640 3496
rect 2634 3491 2635 3495
rect 2639 3491 2640 3495
rect 2634 3490 2640 3491
rect 2770 3495 2776 3496
rect 2770 3491 2771 3495
rect 2775 3491 2776 3495
rect 3023 3495 3029 3496
rect 3023 3494 3024 3495
rect 2981 3492 3024 3494
rect 2770 3490 2776 3491
rect 3023 3491 3024 3492
rect 3028 3491 3029 3495
rect 3170 3495 3176 3496
rect 3170 3494 3171 3495
rect 3117 3492 3171 3494
rect 3023 3490 3029 3491
rect 3170 3491 3171 3492
rect 3175 3491 3176 3495
rect 3170 3490 3176 3491
rect 3250 3495 3256 3496
rect 3250 3491 3251 3495
rect 3255 3491 3256 3495
rect 3250 3490 3256 3491
rect 3386 3495 3392 3496
rect 3386 3491 3387 3495
rect 3391 3491 3392 3495
rect 3386 3490 3392 3491
rect 3450 3495 3456 3496
rect 5406 3495 5412 3496
rect 5542 3500 5548 3501
rect 5542 3496 5543 3500
rect 5547 3496 5548 3500
rect 5662 3497 5663 3501
rect 5667 3497 5668 3501
rect 5662 3496 5668 3497
rect 5542 3495 5548 3496
rect 3450 3491 3451 3495
rect 3455 3491 3456 3495
rect 3450 3490 3456 3491
rect 5378 3485 5384 3486
rect 3838 3484 3844 3485
rect 3838 3480 3839 3484
rect 3843 3480 3844 3484
rect 5378 3481 5379 3485
rect 5383 3481 5384 3485
rect 5378 3480 5384 3481
rect 5514 3485 5520 3486
rect 5514 3481 5515 3485
rect 5519 3481 5520 3485
rect 5514 3480 5520 3481
rect 5662 3484 5668 3485
rect 5662 3480 5663 3484
rect 5667 3480 5668 3484
rect 3838 3479 3844 3480
rect 5662 3479 5668 3480
rect 110 3477 116 3478
rect 1934 3477 1940 3478
rect 110 3473 111 3477
rect 115 3473 116 3477
rect 110 3472 116 3473
rect 430 3476 436 3477
rect 430 3472 431 3476
rect 435 3472 436 3476
rect 430 3471 436 3472
rect 566 3476 572 3477
rect 566 3472 567 3476
rect 571 3472 572 3476
rect 566 3471 572 3472
rect 702 3476 708 3477
rect 702 3472 703 3476
rect 707 3472 708 3476
rect 702 3471 708 3472
rect 838 3476 844 3477
rect 838 3472 839 3476
rect 843 3472 844 3476
rect 838 3471 844 3472
rect 974 3476 980 3477
rect 974 3472 975 3476
rect 979 3472 980 3476
rect 1934 3473 1935 3477
rect 1939 3473 1940 3477
rect 1934 3472 1940 3473
rect 5503 3475 5509 3476
rect 974 3471 980 3472
rect 5503 3471 5504 3475
rect 5508 3474 5509 3475
rect 5530 3475 5536 3476
rect 5530 3474 5531 3475
rect 5508 3472 5531 3474
rect 5508 3471 5509 3472
rect 5503 3470 5509 3471
rect 5530 3471 5531 3472
rect 5535 3471 5536 3475
rect 5530 3470 5536 3471
rect 5602 3475 5608 3476
rect 5602 3471 5603 3475
rect 5607 3474 5608 3475
rect 5639 3475 5645 3476
rect 5639 3474 5640 3475
rect 5607 3472 5640 3474
rect 5607 3471 5608 3472
rect 5602 3470 5608 3471
rect 5639 3471 5640 3472
rect 5644 3471 5645 3475
rect 5639 3470 5645 3471
rect 402 3461 408 3462
rect 110 3460 116 3461
rect 110 3456 111 3460
rect 115 3456 116 3460
rect 402 3457 403 3461
rect 407 3457 408 3461
rect 402 3456 408 3457
rect 538 3461 544 3462
rect 538 3457 539 3461
rect 543 3457 544 3461
rect 538 3456 544 3457
rect 674 3461 680 3462
rect 674 3457 675 3461
rect 679 3457 680 3461
rect 674 3456 680 3457
rect 810 3461 816 3462
rect 810 3457 811 3461
rect 815 3457 816 3461
rect 810 3456 816 3457
rect 946 3461 952 3462
rect 946 3457 947 3461
rect 951 3457 952 3461
rect 946 3456 952 3457
rect 1934 3460 1940 3461
rect 1934 3456 1935 3460
rect 1939 3456 1940 3460
rect 5550 3459 5556 3460
rect 5550 3458 5551 3459
rect 110 3455 116 3456
rect 1934 3455 1940 3456
rect 5520 3456 5551 3458
rect 527 3451 533 3452
rect 527 3447 528 3451
rect 532 3450 533 3451
rect 618 3451 624 3452
rect 618 3450 619 3451
rect 532 3448 619 3450
rect 532 3447 533 3448
rect 527 3446 533 3447
rect 618 3447 619 3448
rect 623 3447 624 3451
rect 618 3446 624 3447
rect 663 3451 669 3452
rect 663 3447 664 3451
rect 668 3450 669 3451
rect 690 3451 696 3452
rect 690 3450 691 3451
rect 668 3448 691 3450
rect 668 3447 669 3448
rect 663 3446 669 3447
rect 690 3447 691 3448
rect 695 3447 696 3451
rect 690 3446 696 3447
rect 799 3451 805 3452
rect 799 3447 800 3451
rect 804 3450 805 3451
rect 818 3451 824 3452
rect 818 3450 819 3451
rect 804 3448 819 3450
rect 804 3447 805 3448
rect 799 3446 805 3447
rect 818 3447 819 3448
rect 823 3447 824 3451
rect 818 3446 824 3447
rect 935 3451 941 3452
rect 935 3447 936 3451
rect 940 3450 941 3451
rect 962 3451 968 3452
rect 962 3450 963 3451
rect 940 3448 963 3450
rect 940 3447 941 3448
rect 935 3446 941 3447
rect 962 3447 963 3448
rect 967 3447 968 3451
rect 962 3446 968 3447
rect 1010 3451 1016 3452
rect 1010 3447 1011 3451
rect 1015 3450 1016 3451
rect 1071 3451 1077 3452
rect 1071 3450 1072 3451
rect 1015 3448 1072 3450
rect 1015 3447 1016 3448
rect 1010 3446 1016 3447
rect 1071 3447 1072 3448
rect 1076 3447 1077 3451
rect 1071 3446 1077 3447
rect 2318 3443 2324 3444
rect 2318 3442 2319 3443
rect 2261 3440 2319 3442
rect 2318 3439 2319 3440
rect 2323 3439 2324 3443
rect 2318 3438 2324 3439
rect 2326 3443 2332 3444
rect 2326 3439 2327 3443
rect 2331 3442 2332 3443
rect 2474 3443 2480 3444
rect 2331 3440 2365 3442
rect 2331 3439 2332 3440
rect 2326 3438 2332 3439
rect 2474 3439 2475 3443
rect 2479 3442 2480 3443
rect 2818 3443 2824 3444
rect 2479 3440 2549 3442
rect 2479 3439 2480 3440
rect 2474 3438 2480 3439
rect 2802 3439 2808 3440
rect 2802 3435 2803 3439
rect 2807 3435 2808 3439
rect 2818 3439 2819 3443
rect 2823 3442 2824 3443
rect 3226 3443 3232 3444
rect 2823 3440 2925 3442
rect 2823 3439 2824 3440
rect 2818 3438 2824 3439
rect 3186 3439 3192 3440
rect 2802 3434 2808 3435
rect 3186 3435 3187 3439
rect 3191 3435 3192 3439
rect 3226 3439 3227 3443
rect 3231 3442 3232 3443
rect 3638 3443 3644 3444
rect 3638 3442 3639 3443
rect 3231 3440 3309 3442
rect 3573 3440 3639 3442
rect 3231 3439 3232 3440
rect 3226 3438 3232 3439
rect 3638 3439 3639 3440
rect 3643 3439 3644 3443
rect 5520 3442 5522 3456
rect 5550 3455 5551 3456
rect 5555 3455 5556 3459
rect 5550 3454 5556 3455
rect 5469 3440 5522 3442
rect 5530 3443 5536 3444
rect 3638 3438 3644 3439
rect 3738 3439 3744 3440
rect 3186 3434 3192 3435
rect 3738 3435 3739 3439
rect 3743 3435 3744 3439
rect 5530 3439 5531 3443
rect 5535 3439 5536 3443
rect 5530 3438 5536 3439
rect 3738 3434 3744 3435
rect 446 3419 452 3420
rect 446 3415 447 3419
rect 451 3415 452 3419
rect 446 3414 452 3415
rect 618 3419 624 3420
rect 618 3415 619 3419
rect 623 3415 624 3419
rect 618 3414 624 3415
rect 690 3419 696 3420
rect 690 3415 691 3419
rect 695 3415 696 3419
rect 690 3414 696 3415
rect 898 3419 904 3420
rect 898 3415 899 3419
rect 903 3415 904 3419
rect 898 3414 904 3415
rect 962 3419 968 3420
rect 962 3415 963 3419
rect 967 3415 968 3419
rect 962 3414 968 3415
rect 2318 3415 2324 3416
rect 2318 3411 2319 3415
rect 2323 3414 2324 3415
rect 3186 3415 3192 3416
rect 2323 3412 2830 3414
rect 2323 3411 2324 3412
rect 2318 3410 2324 3411
rect 2295 3407 2301 3408
rect 2295 3403 2296 3407
rect 2300 3406 2301 3407
rect 2326 3407 2332 3408
rect 2326 3406 2327 3407
rect 2300 3404 2327 3406
rect 2300 3403 2301 3404
rect 2295 3402 2301 3403
rect 2326 3403 2327 3404
rect 2331 3403 2332 3407
rect 2326 3402 2332 3403
rect 2471 3407 2480 3408
rect 2471 3403 2472 3407
rect 2479 3403 2480 3407
rect 2471 3402 2480 3403
rect 2655 3407 2661 3408
rect 2655 3403 2656 3407
rect 2660 3406 2661 3407
rect 2818 3407 2824 3408
rect 2818 3406 2819 3407
rect 2660 3404 2819 3406
rect 2660 3403 2661 3404
rect 2655 3402 2661 3403
rect 2818 3403 2819 3404
rect 2823 3403 2824 3407
rect 2828 3406 2830 3412
rect 3186 3411 3187 3415
rect 3191 3414 3192 3415
rect 3191 3412 3426 3414
rect 3191 3411 3192 3412
rect 3186 3410 3192 3411
rect 2839 3407 2845 3408
rect 2839 3406 2840 3407
rect 2828 3404 2840 3406
rect 2818 3402 2824 3403
rect 2839 3403 2840 3404
rect 2844 3403 2845 3407
rect 2839 3402 2845 3403
rect 3030 3407 3037 3408
rect 3030 3403 3031 3407
rect 3036 3403 3037 3407
rect 3030 3402 3037 3403
rect 3223 3407 3232 3408
rect 3223 3403 3224 3407
rect 3231 3403 3232 3407
rect 3223 3402 3232 3403
rect 3386 3407 3392 3408
rect 3386 3403 3387 3407
rect 3391 3406 3392 3407
rect 3415 3407 3421 3408
rect 3415 3406 3416 3407
rect 3391 3404 3416 3406
rect 3391 3403 3392 3404
rect 3386 3402 3392 3403
rect 3415 3403 3416 3404
rect 3420 3403 3421 3407
rect 3424 3406 3426 3412
rect 3607 3407 3613 3408
rect 3607 3406 3608 3407
rect 3424 3404 3608 3406
rect 3415 3402 3421 3403
rect 3607 3403 3608 3404
rect 3612 3403 3613 3407
rect 3607 3402 3613 3403
rect 3638 3407 3644 3408
rect 3638 3403 3639 3407
rect 3643 3406 3644 3407
rect 3775 3407 3781 3408
rect 3775 3406 3776 3407
rect 3643 3404 3776 3406
rect 3643 3403 3644 3404
rect 3638 3402 3644 3403
rect 3775 3403 3776 3404
rect 3780 3403 3781 3407
rect 3775 3402 3781 3403
rect 1974 3400 1980 3401
rect 3798 3400 3804 3401
rect 1974 3396 1975 3400
rect 1979 3396 1980 3400
rect 1974 3395 1980 3396
rect 2170 3399 2176 3400
rect 2170 3395 2171 3399
rect 2175 3395 2176 3399
rect 2170 3394 2176 3395
rect 2346 3399 2352 3400
rect 2346 3395 2347 3399
rect 2351 3395 2352 3399
rect 2346 3394 2352 3395
rect 2530 3399 2536 3400
rect 2530 3395 2531 3399
rect 2535 3395 2536 3399
rect 2530 3394 2536 3395
rect 2714 3399 2720 3400
rect 2714 3395 2715 3399
rect 2719 3395 2720 3399
rect 2714 3394 2720 3395
rect 2906 3399 2912 3400
rect 2906 3395 2907 3399
rect 2911 3395 2912 3399
rect 2906 3394 2912 3395
rect 3098 3399 3104 3400
rect 3098 3395 3099 3399
rect 3103 3395 3104 3399
rect 3098 3394 3104 3395
rect 3290 3399 3296 3400
rect 3290 3395 3291 3399
rect 3295 3395 3296 3399
rect 3290 3394 3296 3395
rect 3482 3399 3488 3400
rect 3482 3395 3483 3399
rect 3487 3395 3488 3399
rect 3482 3394 3488 3395
rect 3650 3399 3656 3400
rect 3650 3395 3651 3399
rect 3655 3395 3656 3399
rect 3798 3396 3799 3400
rect 3803 3396 3804 3400
rect 3798 3395 3804 3396
rect 3650 3394 3656 3395
rect 4095 3387 4101 3388
rect 4095 3386 4096 3387
rect 2198 3384 2204 3385
rect 1974 3383 1980 3384
rect 1974 3379 1975 3383
rect 1979 3379 1980 3383
rect 2198 3380 2199 3384
rect 2203 3380 2204 3384
rect 2198 3379 2204 3380
rect 2374 3384 2380 3385
rect 2374 3380 2375 3384
rect 2379 3380 2380 3384
rect 2374 3379 2380 3380
rect 2558 3384 2564 3385
rect 2558 3380 2559 3384
rect 2563 3380 2564 3384
rect 2558 3379 2564 3380
rect 2742 3384 2748 3385
rect 2742 3380 2743 3384
rect 2747 3380 2748 3384
rect 2742 3379 2748 3380
rect 2934 3384 2940 3385
rect 2934 3380 2935 3384
rect 2939 3380 2940 3384
rect 2934 3379 2940 3380
rect 3126 3384 3132 3385
rect 3126 3380 3127 3384
rect 3131 3380 3132 3384
rect 3126 3379 3132 3380
rect 3318 3384 3324 3385
rect 3318 3380 3319 3384
rect 3323 3380 3324 3384
rect 3318 3379 3324 3380
rect 3510 3384 3516 3385
rect 3510 3380 3511 3384
rect 3515 3380 3516 3384
rect 3510 3379 3516 3380
rect 3678 3384 3684 3385
rect 3949 3384 4096 3386
rect 3678 3380 3679 3384
rect 3683 3380 3684 3384
rect 3678 3379 3684 3380
rect 3798 3383 3804 3384
rect 3798 3379 3799 3383
rect 3803 3379 3804 3383
rect 4095 3383 4096 3384
rect 4100 3383 4101 3387
rect 4095 3382 4101 3383
rect 4226 3387 4232 3388
rect 4226 3383 4227 3387
rect 4231 3386 4232 3387
rect 4990 3387 4996 3388
rect 4990 3386 4991 3387
rect 4231 3384 4365 3386
rect 4901 3384 4991 3386
rect 4231 3383 4232 3384
rect 4226 3382 4232 3383
rect 4674 3383 4680 3384
rect 1974 3378 1980 3379
rect 3798 3378 3804 3379
rect 4184 3378 4186 3381
rect 4294 3379 4300 3380
rect 4294 3378 4295 3379
rect 4184 3376 4295 3378
rect 4294 3375 4295 3376
rect 4299 3375 4300 3379
rect 4674 3379 4675 3383
rect 4679 3379 4680 3383
rect 4990 3383 4991 3384
rect 4995 3383 4996 3387
rect 5199 3387 5205 3388
rect 5199 3386 5200 3387
rect 5117 3384 5200 3386
rect 4990 3382 4996 3383
rect 5199 3383 5200 3384
rect 5204 3383 5205 3387
rect 5414 3387 5420 3388
rect 5414 3386 5415 3387
rect 5325 3384 5415 3386
rect 5199 3382 5205 3383
rect 5414 3383 5415 3384
rect 5419 3383 5420 3387
rect 5414 3382 5420 3383
rect 5442 3387 5448 3388
rect 5442 3383 5443 3387
rect 5447 3386 5448 3387
rect 5447 3384 5469 3386
rect 5447 3383 5448 3384
rect 5442 3382 5448 3383
rect 4674 3378 4680 3379
rect 4294 3374 4300 3375
rect 455 3363 461 3364
rect 455 3362 456 3363
rect 413 3360 456 3362
rect 455 3359 456 3360
rect 460 3359 461 3363
rect 562 3363 568 3364
rect 562 3362 563 3363
rect 549 3360 563 3362
rect 455 3358 461 3359
rect 562 3359 563 3360
rect 567 3359 568 3363
rect 863 3363 869 3364
rect 562 3358 568 3359
rect 682 3359 688 3360
rect 682 3355 683 3359
rect 687 3355 688 3359
rect 682 3354 688 3355
rect 818 3359 824 3360
rect 818 3355 819 3359
rect 823 3355 824 3359
rect 863 3359 864 3363
rect 868 3362 869 3363
rect 868 3360 885 3362
rect 868 3359 869 3360
rect 863 3358 869 3359
rect 4674 3359 4680 3360
rect 818 3354 824 3355
rect 4674 3355 4675 3359
rect 4679 3358 4680 3359
rect 4679 3356 4821 3358
rect 4679 3355 4680 3356
rect 4674 3354 4680 3355
rect 3738 3351 3744 3352
rect 3738 3347 3739 3351
rect 3743 3350 3744 3351
rect 3983 3351 3989 3352
rect 3983 3350 3984 3351
rect 3743 3348 3984 3350
rect 3743 3347 3744 3348
rect 3738 3346 3744 3347
rect 3983 3347 3984 3348
rect 3988 3347 3989 3351
rect 3983 3346 3989 3347
rect 4095 3351 4101 3352
rect 4095 3347 4096 3351
rect 4100 3350 4101 3351
rect 4223 3351 4229 3352
rect 4223 3350 4224 3351
rect 4100 3348 4224 3350
rect 4100 3347 4101 3348
rect 4095 3346 4101 3347
rect 4223 3347 4224 3348
rect 4228 3347 4229 3351
rect 4223 3346 4229 3347
rect 4294 3351 4300 3352
rect 4294 3347 4295 3351
rect 4299 3350 4300 3351
rect 4471 3351 4477 3352
rect 4471 3350 4472 3351
rect 4299 3348 4472 3350
rect 4299 3347 4300 3348
rect 4294 3346 4300 3347
rect 4471 3347 4472 3348
rect 4476 3347 4477 3351
rect 4471 3346 4477 3347
rect 4711 3351 4717 3352
rect 4711 3347 4712 3351
rect 4716 3350 4717 3351
rect 4802 3351 4808 3352
rect 4802 3350 4803 3351
rect 4716 3348 4803 3350
rect 4716 3347 4717 3348
rect 4711 3346 4717 3347
rect 4802 3347 4803 3348
rect 4807 3347 4808 3351
rect 4819 3350 4821 3356
rect 4935 3351 4941 3352
rect 4935 3350 4936 3351
rect 4819 3348 4936 3350
rect 4802 3346 4808 3347
rect 4935 3347 4936 3348
rect 4940 3347 4941 3351
rect 4935 3346 4941 3347
rect 4990 3351 4996 3352
rect 4990 3347 4991 3351
rect 4995 3350 4996 3351
rect 5151 3351 5157 3352
rect 5151 3350 5152 3351
rect 4995 3348 5152 3350
rect 4995 3347 4996 3348
rect 4990 3346 4996 3347
rect 5151 3347 5152 3348
rect 5156 3347 5157 3351
rect 5151 3346 5157 3347
rect 5199 3351 5205 3352
rect 5199 3347 5200 3351
rect 5204 3350 5205 3351
rect 5359 3351 5365 3352
rect 5359 3350 5360 3351
rect 5204 3348 5360 3350
rect 5204 3347 5205 3348
rect 5199 3346 5205 3347
rect 5359 3347 5360 3348
rect 5364 3347 5365 3351
rect 5359 3346 5365 3347
rect 5414 3351 5420 3352
rect 5414 3347 5415 3351
rect 5419 3350 5420 3351
rect 5575 3351 5581 3352
rect 5575 3350 5576 3351
rect 5419 3348 5576 3350
rect 5419 3347 5420 3348
rect 5414 3346 5420 3347
rect 5575 3347 5576 3348
rect 5580 3347 5581 3351
rect 5575 3346 5581 3347
rect 3838 3344 3844 3345
rect 5662 3344 5668 3345
rect 3838 3340 3839 3344
rect 3843 3340 3844 3344
rect 3838 3339 3844 3340
rect 3858 3343 3864 3344
rect 3858 3339 3859 3343
rect 3863 3339 3864 3343
rect 3858 3338 3864 3339
rect 4098 3343 4104 3344
rect 4098 3339 4099 3343
rect 4103 3339 4104 3343
rect 4098 3338 4104 3339
rect 4346 3343 4352 3344
rect 4346 3339 4347 3343
rect 4351 3339 4352 3343
rect 4346 3338 4352 3339
rect 4586 3343 4592 3344
rect 4586 3339 4587 3343
rect 4591 3339 4592 3343
rect 4586 3338 4592 3339
rect 4810 3343 4816 3344
rect 4810 3339 4811 3343
rect 4815 3339 4816 3343
rect 4810 3338 4816 3339
rect 5026 3343 5032 3344
rect 5026 3339 5027 3343
rect 5031 3339 5032 3343
rect 5026 3338 5032 3339
rect 5234 3343 5240 3344
rect 5234 3339 5235 3343
rect 5239 3339 5240 3343
rect 5234 3338 5240 3339
rect 5450 3343 5456 3344
rect 5450 3339 5451 3343
rect 5455 3339 5456 3343
rect 5662 3340 5663 3344
rect 5667 3340 5668 3344
rect 5662 3339 5668 3340
rect 5450 3338 5456 3339
rect 682 3335 688 3336
rect 682 3331 683 3335
rect 687 3334 688 3335
rect 687 3332 874 3334
rect 687 3331 688 3332
rect 682 3330 688 3331
rect 446 3327 453 3328
rect 446 3323 447 3327
rect 452 3323 453 3327
rect 446 3322 453 3323
rect 455 3327 461 3328
rect 455 3323 456 3327
rect 460 3326 461 3327
rect 583 3327 589 3328
rect 583 3326 584 3327
rect 460 3324 584 3326
rect 460 3323 461 3324
rect 455 3322 461 3323
rect 583 3323 584 3324
rect 588 3323 589 3327
rect 583 3322 589 3323
rect 719 3327 725 3328
rect 719 3323 720 3327
rect 724 3326 725 3327
rect 738 3327 744 3328
rect 738 3326 739 3327
rect 724 3324 739 3326
rect 724 3323 725 3324
rect 719 3322 725 3323
rect 738 3323 739 3324
rect 743 3323 744 3327
rect 738 3322 744 3323
rect 855 3327 861 3328
rect 855 3323 856 3327
rect 860 3326 861 3327
rect 863 3327 869 3328
rect 863 3326 864 3327
rect 860 3324 864 3326
rect 860 3323 861 3324
rect 855 3322 861 3323
rect 863 3323 864 3324
rect 868 3323 869 3327
rect 872 3326 874 3332
rect 3886 3328 3892 3329
rect 991 3327 997 3328
rect 991 3326 992 3327
rect 872 3324 992 3326
rect 863 3322 869 3323
rect 991 3323 992 3324
rect 996 3323 997 3327
rect 991 3322 997 3323
rect 3838 3327 3844 3328
rect 3838 3323 3839 3327
rect 3843 3323 3844 3327
rect 3886 3324 3887 3328
rect 3891 3324 3892 3328
rect 3886 3323 3892 3324
rect 4126 3328 4132 3329
rect 4126 3324 4127 3328
rect 4131 3324 4132 3328
rect 4126 3323 4132 3324
rect 4374 3328 4380 3329
rect 4374 3324 4375 3328
rect 4379 3324 4380 3328
rect 4374 3323 4380 3324
rect 4614 3328 4620 3329
rect 4614 3324 4615 3328
rect 4619 3324 4620 3328
rect 4614 3323 4620 3324
rect 4838 3328 4844 3329
rect 4838 3324 4839 3328
rect 4843 3324 4844 3328
rect 4838 3323 4844 3324
rect 5054 3328 5060 3329
rect 5054 3324 5055 3328
rect 5059 3324 5060 3328
rect 5054 3323 5060 3324
rect 5262 3328 5268 3329
rect 5262 3324 5263 3328
rect 5267 3324 5268 3328
rect 5262 3323 5268 3324
rect 5478 3328 5484 3329
rect 5478 3324 5479 3328
rect 5483 3324 5484 3328
rect 5478 3323 5484 3324
rect 5662 3327 5668 3328
rect 5662 3323 5663 3327
rect 5667 3323 5668 3327
rect 3838 3322 3844 3323
rect 5662 3322 5668 3323
rect 110 3320 116 3321
rect 1934 3320 1940 3321
rect 110 3316 111 3320
rect 115 3316 116 3320
rect 110 3315 116 3316
rect 322 3319 328 3320
rect 322 3315 323 3319
rect 327 3315 328 3319
rect 322 3314 328 3315
rect 458 3319 464 3320
rect 458 3315 459 3319
rect 463 3315 464 3319
rect 458 3314 464 3315
rect 594 3319 600 3320
rect 594 3315 595 3319
rect 599 3315 600 3319
rect 594 3314 600 3315
rect 730 3319 736 3320
rect 730 3315 731 3319
rect 735 3315 736 3319
rect 730 3314 736 3315
rect 866 3319 872 3320
rect 866 3315 867 3319
rect 871 3315 872 3319
rect 1934 3316 1935 3320
rect 1939 3316 1940 3320
rect 1934 3315 1940 3316
rect 866 3314 872 3315
rect 350 3304 356 3305
rect 110 3303 116 3304
rect 110 3299 111 3303
rect 115 3299 116 3303
rect 350 3300 351 3304
rect 355 3300 356 3304
rect 350 3299 356 3300
rect 486 3304 492 3305
rect 486 3300 487 3304
rect 491 3300 492 3304
rect 486 3299 492 3300
rect 622 3304 628 3305
rect 622 3300 623 3304
rect 627 3300 628 3304
rect 622 3299 628 3300
rect 758 3304 764 3305
rect 758 3300 759 3304
rect 763 3300 764 3304
rect 758 3299 764 3300
rect 894 3304 900 3305
rect 894 3300 895 3304
rect 899 3300 900 3304
rect 894 3299 900 3300
rect 1934 3303 1940 3304
rect 1934 3299 1935 3303
rect 1939 3299 1940 3303
rect 110 3298 116 3299
rect 1934 3298 1940 3299
rect 1974 3301 1980 3302
rect 3798 3301 3804 3302
rect 1974 3297 1975 3301
rect 1979 3297 1980 3301
rect 1974 3296 1980 3297
rect 2150 3300 2156 3301
rect 2150 3296 2151 3300
rect 2155 3296 2156 3300
rect 2150 3295 2156 3296
rect 2398 3300 2404 3301
rect 2398 3296 2399 3300
rect 2403 3296 2404 3300
rect 2398 3295 2404 3296
rect 2686 3300 2692 3301
rect 2686 3296 2687 3300
rect 2691 3296 2692 3300
rect 2686 3295 2692 3296
rect 3014 3300 3020 3301
rect 3014 3296 3015 3300
rect 3019 3296 3020 3300
rect 3014 3295 3020 3296
rect 3358 3300 3364 3301
rect 3358 3296 3359 3300
rect 3363 3296 3364 3300
rect 3358 3295 3364 3296
rect 3678 3300 3684 3301
rect 3678 3296 3679 3300
rect 3683 3296 3684 3300
rect 3798 3297 3799 3301
rect 3803 3297 3804 3301
rect 3798 3296 3804 3297
rect 3678 3295 3684 3296
rect 2122 3285 2128 3286
rect 1974 3284 1980 3285
rect 1974 3280 1975 3284
rect 1979 3280 1980 3284
rect 2122 3281 2123 3285
rect 2127 3281 2128 3285
rect 2122 3280 2128 3281
rect 2370 3285 2376 3286
rect 2370 3281 2371 3285
rect 2375 3281 2376 3285
rect 2370 3280 2376 3281
rect 2658 3285 2664 3286
rect 2658 3281 2659 3285
rect 2663 3281 2664 3285
rect 2658 3280 2664 3281
rect 2986 3285 2992 3286
rect 2986 3281 2987 3285
rect 2991 3281 2992 3285
rect 2986 3280 2992 3281
rect 3330 3285 3336 3286
rect 3330 3281 3331 3285
rect 3335 3281 3336 3285
rect 3330 3280 3336 3281
rect 3650 3285 3656 3286
rect 3650 3281 3651 3285
rect 3655 3281 3656 3285
rect 3650 3280 3656 3281
rect 3798 3284 3804 3285
rect 3798 3280 3799 3284
rect 3803 3280 3804 3284
rect 1974 3279 1980 3280
rect 3798 3279 3804 3280
rect 2247 3275 2253 3276
rect 2247 3271 2248 3275
rect 2252 3274 2253 3275
rect 2386 3275 2392 3276
rect 2386 3274 2387 3275
rect 2252 3272 2387 3274
rect 2252 3271 2253 3272
rect 2247 3270 2253 3271
rect 2386 3271 2387 3272
rect 2391 3271 2392 3275
rect 2386 3270 2392 3271
rect 2495 3275 2501 3276
rect 2495 3271 2496 3275
rect 2500 3274 2501 3275
rect 2674 3275 2680 3276
rect 2674 3274 2675 3275
rect 2500 3272 2675 3274
rect 2500 3271 2501 3272
rect 2495 3270 2501 3271
rect 2674 3271 2675 3272
rect 2679 3271 2680 3275
rect 2674 3270 2680 3271
rect 2682 3275 2688 3276
rect 2682 3271 2683 3275
rect 2687 3274 2688 3275
rect 2783 3275 2789 3276
rect 2783 3274 2784 3275
rect 2687 3272 2784 3274
rect 2687 3271 2688 3272
rect 2682 3270 2688 3271
rect 2783 3271 2784 3272
rect 2788 3271 2789 3275
rect 2783 3270 2789 3271
rect 3111 3275 3117 3276
rect 3111 3271 3112 3275
rect 3116 3274 3117 3275
rect 3182 3275 3188 3276
rect 3182 3274 3183 3275
rect 3116 3272 3183 3274
rect 3116 3271 3117 3272
rect 3111 3270 3117 3271
rect 3182 3271 3183 3272
rect 3187 3271 3188 3275
rect 3455 3275 3461 3276
rect 3455 3274 3456 3275
rect 3182 3270 3188 3271
rect 3300 3272 3456 3274
rect 3087 3267 3093 3268
rect 3087 3263 3088 3267
rect 3092 3266 3093 3267
rect 3300 3266 3302 3272
rect 3455 3271 3456 3272
rect 3460 3271 3461 3275
rect 3455 3270 3461 3271
rect 3775 3275 3784 3276
rect 3775 3271 3776 3275
rect 3783 3271 3784 3275
rect 3775 3270 3784 3271
rect 3092 3264 3302 3266
rect 3838 3269 3844 3270
rect 5662 3269 5668 3270
rect 3838 3265 3839 3269
rect 3843 3265 3844 3269
rect 3838 3264 3844 3265
rect 3886 3268 3892 3269
rect 3886 3264 3887 3268
rect 3891 3264 3892 3268
rect 3092 3263 3093 3264
rect 3886 3263 3892 3264
rect 4126 3268 4132 3269
rect 4126 3264 4127 3268
rect 4131 3264 4132 3268
rect 4126 3263 4132 3264
rect 4374 3268 4380 3269
rect 4374 3264 4375 3268
rect 4379 3264 4380 3268
rect 4374 3263 4380 3264
rect 4606 3268 4612 3269
rect 4606 3264 4607 3268
rect 4611 3264 4612 3268
rect 4606 3263 4612 3264
rect 4814 3268 4820 3269
rect 4814 3264 4815 3268
rect 4819 3264 4820 3268
rect 4814 3263 4820 3264
rect 5014 3268 5020 3269
rect 5014 3264 5015 3268
rect 5019 3264 5020 3268
rect 5014 3263 5020 3264
rect 5198 3268 5204 3269
rect 5198 3264 5199 3268
rect 5203 3264 5204 3268
rect 5198 3263 5204 3264
rect 5382 3268 5388 3269
rect 5382 3264 5383 3268
rect 5387 3264 5388 3268
rect 5382 3263 5388 3264
rect 5542 3268 5548 3269
rect 5542 3264 5543 3268
rect 5547 3264 5548 3268
rect 5662 3265 5663 3269
rect 5667 3265 5668 3269
rect 5662 3264 5668 3265
rect 5542 3263 5548 3264
rect 3087 3262 3093 3263
rect 3858 3253 3864 3254
rect 3838 3252 3844 3253
rect 3838 3248 3839 3252
rect 3843 3248 3844 3252
rect 3858 3249 3859 3253
rect 3863 3249 3864 3253
rect 3858 3248 3864 3249
rect 4098 3253 4104 3254
rect 4098 3249 4099 3253
rect 4103 3249 4104 3253
rect 4098 3248 4104 3249
rect 4346 3253 4352 3254
rect 4346 3249 4347 3253
rect 4351 3249 4352 3253
rect 4346 3248 4352 3249
rect 4578 3253 4584 3254
rect 4578 3249 4579 3253
rect 4583 3249 4584 3253
rect 4578 3248 4584 3249
rect 4786 3253 4792 3254
rect 4786 3249 4787 3253
rect 4791 3249 4792 3253
rect 4786 3248 4792 3249
rect 4986 3253 4992 3254
rect 4986 3249 4987 3253
rect 4991 3249 4992 3253
rect 4986 3248 4992 3249
rect 5170 3253 5176 3254
rect 5170 3249 5171 3253
rect 5175 3249 5176 3253
rect 5170 3248 5176 3249
rect 5354 3253 5360 3254
rect 5354 3249 5355 3253
rect 5359 3249 5360 3253
rect 5354 3248 5360 3249
rect 5514 3253 5520 3254
rect 5514 3249 5515 3253
rect 5519 3249 5520 3253
rect 5514 3248 5520 3249
rect 5662 3252 5668 3253
rect 5662 3248 5663 3252
rect 5667 3248 5668 3252
rect 3838 3247 3844 3248
rect 5662 3247 5668 3248
rect 2290 3243 2296 3244
rect 2290 3242 2291 3243
rect 2213 3240 2291 3242
rect 2290 3239 2291 3240
rect 2295 3239 2296 3243
rect 2290 3238 2296 3239
rect 2386 3243 2392 3244
rect 2386 3239 2387 3243
rect 2391 3239 2392 3243
rect 2386 3238 2392 3239
rect 2674 3243 2680 3244
rect 2674 3239 2675 3243
rect 2679 3239 2680 3243
rect 2674 3238 2680 3239
rect 3030 3243 3036 3244
rect 3030 3239 3031 3243
rect 3035 3239 3036 3243
rect 3030 3238 3036 3239
rect 3182 3243 3188 3244
rect 3182 3239 3183 3243
rect 3187 3242 3188 3243
rect 3738 3243 3744 3244
rect 3187 3240 3349 3242
rect 3187 3239 3188 3240
rect 3182 3238 3188 3239
rect 3738 3239 3739 3243
rect 3743 3239 3744 3243
rect 3738 3238 3744 3239
rect 3983 3243 3989 3244
rect 3983 3239 3984 3243
rect 3988 3242 3989 3243
rect 4114 3243 4120 3244
rect 4114 3242 4115 3243
rect 3988 3240 4115 3242
rect 3988 3239 3989 3240
rect 3983 3238 3989 3239
rect 4114 3239 4115 3240
rect 4119 3239 4120 3243
rect 4114 3238 4120 3239
rect 4223 3243 4232 3244
rect 4223 3239 4224 3243
rect 4231 3239 4232 3243
rect 4223 3238 4232 3239
rect 4471 3243 4477 3244
rect 4471 3239 4472 3243
rect 4476 3242 4477 3243
rect 4594 3243 4600 3244
rect 4594 3242 4595 3243
rect 4476 3240 4595 3242
rect 4476 3239 4477 3240
rect 4471 3238 4477 3239
rect 4594 3239 4595 3240
rect 4599 3239 4600 3243
rect 4594 3238 4600 3239
rect 4703 3243 4709 3244
rect 4703 3239 4704 3243
rect 4708 3242 4709 3243
rect 4758 3243 4764 3244
rect 4758 3242 4759 3243
rect 4708 3240 4759 3242
rect 4708 3239 4709 3240
rect 4703 3238 4709 3239
rect 4758 3239 4759 3240
rect 4763 3239 4764 3243
rect 4758 3238 4764 3239
rect 4911 3243 4917 3244
rect 4911 3239 4912 3243
rect 4916 3242 4917 3243
rect 5002 3243 5008 3244
rect 5002 3242 5003 3243
rect 4916 3240 5003 3242
rect 4916 3239 4917 3240
rect 4911 3238 4917 3239
rect 5002 3239 5003 3240
rect 5007 3239 5008 3243
rect 5111 3243 5117 3244
rect 5111 3242 5112 3243
rect 5002 3238 5008 3239
rect 5012 3240 5112 3242
rect 110 3237 116 3238
rect 1934 3237 1940 3238
rect 110 3233 111 3237
rect 115 3233 116 3237
rect 110 3232 116 3233
rect 158 3236 164 3237
rect 158 3232 159 3236
rect 163 3232 164 3236
rect 158 3231 164 3232
rect 334 3236 340 3237
rect 334 3232 335 3236
rect 339 3232 340 3236
rect 334 3231 340 3232
rect 542 3236 548 3237
rect 542 3232 543 3236
rect 547 3232 548 3236
rect 542 3231 548 3232
rect 750 3236 756 3237
rect 750 3232 751 3236
rect 755 3232 756 3236
rect 750 3231 756 3232
rect 958 3236 964 3237
rect 958 3232 959 3236
rect 963 3232 964 3236
rect 1934 3233 1935 3237
rect 1939 3233 1940 3237
rect 1934 3232 1940 3233
rect 4434 3235 4440 3236
rect 958 3231 964 3232
rect 4434 3231 4435 3235
rect 4439 3234 4440 3235
rect 5012 3234 5014 3240
rect 5111 3239 5112 3240
rect 5116 3239 5117 3243
rect 5111 3238 5117 3239
rect 5295 3243 5301 3244
rect 5295 3239 5296 3243
rect 5300 3242 5301 3243
rect 5370 3243 5376 3244
rect 5370 3242 5371 3243
rect 5300 3240 5371 3242
rect 5300 3239 5301 3240
rect 5295 3238 5301 3239
rect 5370 3239 5371 3240
rect 5375 3239 5376 3243
rect 5370 3238 5376 3239
rect 5442 3243 5448 3244
rect 5442 3239 5443 3243
rect 5447 3242 5448 3243
rect 5479 3243 5485 3244
rect 5479 3242 5480 3243
rect 5447 3240 5480 3242
rect 5447 3239 5448 3240
rect 5442 3238 5448 3239
rect 5479 3239 5480 3240
rect 5484 3239 5485 3243
rect 5479 3238 5485 3239
rect 5618 3243 5624 3244
rect 5618 3239 5619 3243
rect 5623 3242 5624 3243
rect 5639 3243 5645 3244
rect 5639 3242 5640 3243
rect 5623 3240 5640 3242
rect 5623 3239 5624 3240
rect 5618 3238 5624 3239
rect 5639 3239 5640 3240
rect 5644 3239 5645 3243
rect 5639 3238 5645 3239
rect 4439 3232 5014 3234
rect 4439 3231 4440 3232
rect 4434 3230 4440 3231
rect 130 3221 136 3222
rect 110 3220 116 3221
rect 110 3216 111 3220
rect 115 3216 116 3220
rect 130 3217 131 3221
rect 135 3217 136 3221
rect 130 3216 136 3217
rect 306 3221 312 3222
rect 306 3217 307 3221
rect 311 3217 312 3221
rect 306 3216 312 3217
rect 514 3221 520 3222
rect 514 3217 515 3221
rect 519 3217 520 3221
rect 514 3216 520 3217
rect 722 3221 728 3222
rect 722 3217 723 3221
rect 727 3217 728 3221
rect 722 3216 728 3217
rect 930 3221 936 3222
rect 930 3217 931 3221
rect 935 3217 936 3221
rect 930 3216 936 3217
rect 1934 3220 1940 3221
rect 1934 3216 1935 3220
rect 1939 3216 1940 3220
rect 110 3215 116 3216
rect 1934 3215 1940 3216
rect 255 3211 261 3212
rect 255 3207 256 3211
rect 260 3210 261 3211
rect 322 3211 328 3212
rect 322 3210 323 3211
rect 260 3208 323 3210
rect 260 3207 261 3208
rect 255 3206 261 3207
rect 322 3207 323 3208
rect 327 3207 328 3211
rect 322 3206 328 3207
rect 431 3211 437 3212
rect 431 3207 432 3211
rect 436 3210 437 3211
rect 530 3211 536 3212
rect 530 3210 531 3211
rect 436 3208 531 3210
rect 436 3207 437 3208
rect 431 3206 437 3207
rect 530 3207 531 3208
rect 535 3207 536 3211
rect 530 3206 536 3207
rect 562 3211 568 3212
rect 562 3207 563 3211
rect 567 3210 568 3211
rect 639 3211 645 3212
rect 639 3210 640 3211
rect 567 3208 640 3210
rect 567 3207 568 3208
rect 562 3206 568 3207
rect 639 3207 640 3208
rect 644 3207 645 3211
rect 639 3206 645 3207
rect 847 3211 853 3212
rect 847 3207 848 3211
rect 852 3210 853 3211
rect 946 3211 952 3212
rect 946 3210 947 3211
rect 852 3208 947 3210
rect 852 3207 853 3208
rect 847 3206 853 3207
rect 946 3207 947 3208
rect 951 3207 952 3211
rect 946 3206 952 3207
rect 1055 3211 1064 3212
rect 1055 3207 1056 3211
rect 1063 3207 1064 3211
rect 1055 3206 1064 3207
rect 3778 3211 3784 3212
rect 3778 3207 3779 3211
rect 3783 3210 3784 3211
rect 4114 3211 4120 3212
rect 3783 3208 3877 3210
rect 3783 3207 3784 3208
rect 3778 3206 3784 3207
rect 4114 3207 4115 3211
rect 4119 3207 4120 3211
rect 4114 3206 4120 3207
rect 4434 3211 4440 3212
rect 4434 3207 4435 3211
rect 4439 3207 4440 3211
rect 4434 3206 4440 3207
rect 4594 3211 4600 3212
rect 4594 3207 4595 3211
rect 4599 3207 4600 3211
rect 4594 3206 4600 3207
rect 4802 3211 4808 3212
rect 4802 3207 4803 3211
rect 4807 3207 4808 3211
rect 4802 3206 4808 3207
rect 5002 3211 5008 3212
rect 5002 3207 5003 3211
rect 5007 3207 5008 3211
rect 5362 3211 5368 3212
rect 5362 3210 5363 3211
rect 5261 3208 5363 3210
rect 5002 3206 5008 3207
rect 5362 3207 5363 3208
rect 5367 3207 5368 3211
rect 5362 3206 5368 3207
rect 5370 3211 5376 3212
rect 5370 3207 5371 3211
rect 5375 3207 5376 3211
rect 5370 3206 5376 3207
rect 5602 3211 5608 3212
rect 5602 3207 5603 3211
rect 5607 3207 5608 3211
rect 5602 3206 5608 3207
rect 2682 3203 2688 3204
rect 2682 3202 2683 3203
rect 2676 3200 2683 3202
rect 1914 3195 1920 3196
rect 1914 3191 1915 3195
rect 1919 3194 1920 3195
rect 2122 3195 2128 3196
rect 1919 3192 2013 3194
rect 1919 3191 1920 3192
rect 1914 3190 1920 3191
rect 2122 3191 2123 3195
rect 2127 3194 2128 3195
rect 2274 3195 2280 3196
rect 2127 3192 2165 3194
rect 2127 3191 2128 3192
rect 2122 3190 2128 3191
rect 2274 3191 2275 3195
rect 2279 3194 2280 3195
rect 2676 3194 2678 3200
rect 2682 3199 2683 3200
rect 2687 3199 2688 3203
rect 2682 3198 2688 3199
rect 2279 3192 2365 3194
rect 2645 3192 2678 3194
rect 2682 3195 2688 3196
rect 2279 3191 2280 3192
rect 2274 3190 2280 3191
rect 2682 3191 2683 3195
rect 2687 3194 2688 3195
rect 3087 3195 3093 3196
rect 3087 3194 3088 3195
rect 2687 3192 2789 3194
rect 3077 3192 3088 3194
rect 2687 3191 2688 3192
rect 2682 3190 2688 3191
rect 3087 3191 3088 3192
rect 3092 3191 3093 3195
rect 3087 3190 3093 3191
rect 3414 3195 3420 3196
rect 3414 3191 3415 3195
rect 3419 3194 3420 3195
rect 3570 3195 3576 3196
rect 3419 3192 3461 3194
rect 3419 3191 3420 3192
rect 3414 3190 3420 3191
rect 3570 3191 3571 3195
rect 3575 3194 3576 3195
rect 3575 3192 3669 3194
rect 3575 3191 3576 3192
rect 3570 3190 3576 3191
rect 3296 3186 3298 3189
rect 3382 3187 3388 3188
rect 3382 3186 3383 3187
rect 3296 3184 3383 3186
rect 3382 3183 3383 3184
rect 3387 3183 3388 3187
rect 3382 3182 3388 3183
rect 226 3179 232 3180
rect 226 3178 227 3179
rect 221 3176 227 3178
rect 226 3175 227 3176
rect 231 3175 232 3179
rect 226 3174 232 3175
rect 322 3179 328 3180
rect 322 3175 323 3179
rect 327 3175 328 3179
rect 322 3174 328 3175
rect 530 3179 536 3180
rect 530 3175 531 3179
rect 535 3175 536 3179
rect 530 3174 536 3175
rect 738 3179 744 3180
rect 738 3175 739 3179
rect 743 3175 744 3179
rect 738 3174 744 3175
rect 946 3179 952 3180
rect 946 3175 947 3179
rect 951 3175 952 3179
rect 946 3174 952 3175
rect 2119 3159 2128 3160
rect 2119 3155 2120 3159
rect 2127 3155 2128 3159
rect 2119 3154 2128 3155
rect 2271 3159 2280 3160
rect 2271 3155 2272 3159
rect 2279 3155 2280 3159
rect 2271 3154 2280 3155
rect 2290 3159 2296 3160
rect 2290 3155 2291 3159
rect 2295 3158 2296 3159
rect 2471 3159 2477 3160
rect 2471 3158 2472 3159
rect 2295 3156 2472 3158
rect 2295 3155 2296 3156
rect 2290 3154 2296 3155
rect 2471 3155 2472 3156
rect 2476 3155 2477 3159
rect 2471 3154 2477 3155
rect 2679 3159 2688 3160
rect 2679 3155 2680 3159
rect 2687 3155 2688 3159
rect 2679 3154 2688 3155
rect 2895 3159 2901 3160
rect 2895 3155 2896 3159
rect 2900 3158 2901 3159
rect 2914 3159 2920 3160
rect 2914 3158 2915 3159
rect 2900 3156 2915 3158
rect 2900 3155 2901 3156
rect 2895 3154 2901 3155
rect 2914 3155 2915 3156
rect 2919 3155 2920 3159
rect 2914 3154 2920 3155
rect 3022 3159 3028 3160
rect 3022 3155 3023 3159
rect 3027 3158 3028 3159
rect 3111 3159 3117 3160
rect 3111 3158 3112 3159
rect 3027 3156 3112 3158
rect 3027 3155 3028 3156
rect 3022 3154 3028 3155
rect 3111 3155 3112 3156
rect 3116 3155 3117 3159
rect 3111 3154 3117 3155
rect 3335 3159 3341 3160
rect 3335 3155 3336 3159
rect 3340 3158 3341 3159
rect 3414 3159 3420 3160
rect 3414 3158 3415 3159
rect 3340 3156 3415 3158
rect 3340 3155 3341 3156
rect 3335 3154 3341 3155
rect 3414 3155 3415 3156
rect 3419 3155 3420 3159
rect 3414 3154 3420 3155
rect 3567 3159 3576 3160
rect 3567 3155 3568 3159
rect 3575 3155 3576 3159
rect 3567 3154 3576 3155
rect 3738 3159 3744 3160
rect 3738 3155 3739 3159
rect 3743 3158 3744 3159
rect 3775 3159 3781 3160
rect 3775 3158 3776 3159
rect 3743 3156 3776 3158
rect 3743 3155 3744 3156
rect 3738 3154 3744 3155
rect 3775 3155 3776 3156
rect 3780 3155 3781 3159
rect 3775 3154 3781 3155
rect 1974 3152 1980 3153
rect 3798 3152 3804 3153
rect 1974 3148 1975 3152
rect 1979 3148 1980 3152
rect 1974 3147 1980 3148
rect 1994 3151 2000 3152
rect 1994 3147 1995 3151
rect 1999 3147 2000 3151
rect 1994 3146 2000 3147
rect 2146 3151 2152 3152
rect 2146 3147 2147 3151
rect 2151 3147 2152 3151
rect 2146 3146 2152 3147
rect 2346 3151 2352 3152
rect 2346 3147 2347 3151
rect 2351 3147 2352 3151
rect 2346 3146 2352 3147
rect 2554 3151 2560 3152
rect 2554 3147 2555 3151
rect 2559 3147 2560 3151
rect 2554 3146 2560 3147
rect 2770 3151 2776 3152
rect 2770 3147 2771 3151
rect 2775 3147 2776 3151
rect 2770 3146 2776 3147
rect 2986 3151 2992 3152
rect 2986 3147 2987 3151
rect 2991 3147 2992 3151
rect 2986 3146 2992 3147
rect 3210 3151 3216 3152
rect 3210 3147 3211 3151
rect 3215 3147 3216 3151
rect 3210 3146 3216 3147
rect 3442 3151 3448 3152
rect 3442 3147 3443 3151
rect 3447 3147 3448 3151
rect 3442 3146 3448 3147
rect 3650 3151 3656 3152
rect 3650 3147 3651 3151
rect 3655 3147 3656 3151
rect 3798 3148 3799 3152
rect 3803 3148 3804 3152
rect 3798 3147 3804 3148
rect 4758 3147 4764 3148
rect 3650 3146 3656 3147
rect 4554 3143 4560 3144
rect 4554 3139 4555 3143
rect 4559 3139 4560 3143
rect 4758 3143 4759 3147
rect 4763 3146 4764 3147
rect 4986 3147 4992 3148
rect 4763 3144 4877 3146
rect 4763 3143 4764 3144
rect 4758 3142 4764 3143
rect 4986 3143 4987 3147
rect 4991 3146 4992 3147
rect 5202 3147 5208 3148
rect 4991 3144 5093 3146
rect 4991 3143 4992 3144
rect 4986 3142 4992 3143
rect 5202 3143 5203 3147
rect 5207 3146 5208 3147
rect 5618 3147 5624 3148
rect 5618 3146 5619 3147
rect 5207 3144 5325 3146
rect 5605 3144 5619 3146
rect 5207 3143 5208 3144
rect 5202 3142 5208 3143
rect 5618 3143 5619 3144
rect 5623 3143 5624 3147
rect 5618 3142 5624 3143
rect 4554 3138 4560 3139
rect 2022 3136 2028 3137
rect 1974 3135 1980 3136
rect 1974 3131 1975 3135
rect 1979 3131 1980 3135
rect 2022 3132 2023 3136
rect 2027 3132 2028 3136
rect 2022 3131 2028 3132
rect 2174 3136 2180 3137
rect 2174 3132 2175 3136
rect 2179 3132 2180 3136
rect 2174 3131 2180 3132
rect 2374 3136 2380 3137
rect 2374 3132 2375 3136
rect 2379 3132 2380 3136
rect 2374 3131 2380 3132
rect 2582 3136 2588 3137
rect 2582 3132 2583 3136
rect 2587 3132 2588 3136
rect 2582 3131 2588 3132
rect 2798 3136 2804 3137
rect 2798 3132 2799 3136
rect 2803 3132 2804 3136
rect 2798 3131 2804 3132
rect 3014 3136 3020 3137
rect 3014 3132 3015 3136
rect 3019 3132 3020 3136
rect 3014 3131 3020 3132
rect 3238 3136 3244 3137
rect 3238 3132 3239 3136
rect 3243 3132 3244 3136
rect 3238 3131 3244 3132
rect 3470 3136 3476 3137
rect 3470 3132 3471 3136
rect 3475 3132 3476 3136
rect 3470 3131 3476 3132
rect 3678 3136 3684 3137
rect 3678 3132 3679 3136
rect 3683 3132 3684 3136
rect 3678 3131 3684 3132
rect 3798 3135 3804 3136
rect 3798 3131 3799 3135
rect 3803 3131 3804 3135
rect 1974 3130 1980 3131
rect 3798 3130 3804 3131
rect 4736 3130 4738 3141
rect 5430 3131 5436 3132
rect 5430 3130 5431 3131
rect 4736 3128 5431 3130
rect 5430 3127 5431 3128
rect 5435 3127 5436 3131
rect 5430 3126 5436 3127
rect 4554 3119 4560 3120
rect 319 3115 325 3116
rect 319 3114 320 3115
rect 221 3112 320 3114
rect 319 3111 320 3112
rect 324 3111 325 3115
rect 319 3110 325 3111
rect 330 3115 336 3116
rect 330 3111 331 3115
rect 335 3114 336 3115
rect 822 3115 828 3116
rect 822 3114 823 3115
rect 335 3112 389 3114
rect 717 3112 823 3114
rect 335 3111 336 3112
rect 330 3110 336 3111
rect 822 3111 823 3112
rect 827 3111 828 3115
rect 1050 3115 1056 3116
rect 1050 3114 1051 3115
rect 965 3112 1051 3114
rect 822 3110 828 3111
rect 1050 3111 1051 3112
rect 1055 3111 1056 3115
rect 1050 3110 1056 3111
rect 1058 3115 1064 3116
rect 1058 3111 1059 3115
rect 1063 3114 1064 3115
rect 1450 3115 1456 3116
rect 1450 3114 1451 3115
rect 1063 3112 1133 3114
rect 1437 3112 1451 3114
rect 1063 3111 1064 3112
rect 1058 3110 1064 3111
rect 1450 3111 1451 3112
rect 1455 3111 1456 3115
rect 1450 3110 1456 3111
rect 1474 3115 1480 3116
rect 1474 3111 1475 3115
rect 1479 3114 1480 3115
rect 1706 3115 1712 3116
rect 1479 3112 1597 3114
rect 1479 3111 1480 3112
rect 1474 3110 1480 3111
rect 1706 3111 1707 3115
rect 1711 3114 1712 3115
rect 4554 3115 4555 3119
rect 4559 3118 4560 3119
rect 4559 3116 4670 3118
rect 4559 3115 4560 3116
rect 4554 3114 4560 3115
rect 1711 3112 1805 3114
rect 1711 3111 1712 3112
rect 1706 3110 1712 3111
rect 4591 3111 4597 3112
rect 4591 3107 4592 3111
rect 4596 3110 4597 3111
rect 4658 3111 4664 3112
rect 4658 3110 4659 3111
rect 4596 3108 4659 3110
rect 4596 3107 4597 3108
rect 4591 3106 4597 3107
rect 4658 3107 4659 3108
rect 4663 3107 4664 3111
rect 4668 3110 4670 3116
rect 4775 3111 4781 3112
rect 4775 3110 4776 3111
rect 4668 3108 4776 3110
rect 4658 3106 4664 3107
rect 4775 3107 4776 3108
rect 4780 3107 4781 3111
rect 4775 3106 4781 3107
rect 4983 3111 4992 3112
rect 4983 3107 4984 3111
rect 4991 3107 4992 3111
rect 4983 3106 4992 3107
rect 5199 3111 5208 3112
rect 5199 3107 5200 3111
rect 5207 3107 5208 3111
rect 5199 3106 5208 3107
rect 5430 3111 5437 3112
rect 5430 3107 5431 3111
rect 5436 3107 5437 3111
rect 5430 3106 5437 3107
rect 5618 3111 5624 3112
rect 5618 3107 5619 3111
rect 5623 3110 5624 3111
rect 5639 3111 5645 3112
rect 5639 3110 5640 3111
rect 5623 3108 5640 3110
rect 5623 3107 5624 3108
rect 5618 3106 5624 3107
rect 5639 3107 5640 3108
rect 5644 3107 5645 3111
rect 5639 3106 5645 3107
rect 3838 3104 3844 3105
rect 5662 3104 5668 3105
rect 3838 3100 3839 3104
rect 3843 3100 3844 3104
rect 3838 3099 3844 3100
rect 4466 3103 4472 3104
rect 4466 3099 4467 3103
rect 4471 3099 4472 3103
rect 4466 3098 4472 3099
rect 4650 3103 4656 3104
rect 4650 3099 4651 3103
rect 4655 3099 4656 3103
rect 4650 3098 4656 3099
rect 4858 3103 4864 3104
rect 4858 3099 4859 3103
rect 4863 3099 4864 3103
rect 4858 3098 4864 3099
rect 5074 3103 5080 3104
rect 5074 3099 5075 3103
rect 5079 3099 5080 3103
rect 5074 3098 5080 3099
rect 5306 3103 5312 3104
rect 5306 3099 5307 3103
rect 5311 3099 5312 3103
rect 5306 3098 5312 3099
rect 5514 3103 5520 3104
rect 5514 3099 5515 3103
rect 5519 3099 5520 3103
rect 5662 3100 5663 3104
rect 5667 3100 5668 3104
rect 5662 3099 5668 3100
rect 5514 3098 5520 3099
rect 4494 3088 4500 3089
rect 3838 3087 3844 3088
rect 3838 3083 3839 3087
rect 3843 3083 3844 3087
rect 4494 3084 4495 3088
rect 4499 3084 4500 3088
rect 4494 3083 4500 3084
rect 4678 3088 4684 3089
rect 4678 3084 4679 3088
rect 4683 3084 4684 3088
rect 4678 3083 4684 3084
rect 4886 3088 4892 3089
rect 4886 3084 4887 3088
rect 4891 3084 4892 3088
rect 4886 3083 4892 3084
rect 5102 3088 5108 3089
rect 5102 3084 5103 3088
rect 5107 3084 5108 3088
rect 5102 3083 5108 3084
rect 5334 3088 5340 3089
rect 5334 3084 5335 3088
rect 5339 3084 5340 3088
rect 5334 3083 5340 3084
rect 5542 3088 5548 3089
rect 5542 3084 5543 3088
rect 5547 3084 5548 3088
rect 5542 3083 5548 3084
rect 5662 3087 5668 3088
rect 5662 3083 5663 3087
rect 5667 3083 5668 3087
rect 3838 3082 3844 3083
rect 5662 3082 5668 3083
rect 226 3079 232 3080
rect 226 3075 227 3079
rect 231 3078 232 3079
rect 255 3079 261 3080
rect 255 3078 256 3079
rect 231 3076 256 3078
rect 231 3075 232 3076
rect 226 3074 232 3075
rect 255 3075 256 3076
rect 260 3075 261 3079
rect 255 3074 261 3075
rect 319 3079 325 3080
rect 319 3075 320 3079
rect 324 3078 325 3079
rect 495 3079 501 3080
rect 495 3078 496 3079
rect 324 3076 496 3078
rect 324 3075 325 3076
rect 319 3074 325 3075
rect 495 3075 496 3076
rect 500 3075 501 3079
rect 495 3074 501 3075
rect 682 3079 688 3080
rect 682 3075 683 3079
rect 687 3078 688 3079
rect 751 3079 757 3080
rect 751 3078 752 3079
rect 687 3076 752 3078
rect 687 3075 688 3076
rect 682 3074 688 3075
rect 751 3075 752 3076
rect 756 3075 757 3079
rect 751 3074 757 3075
rect 822 3079 828 3080
rect 822 3075 823 3079
rect 827 3078 828 3079
rect 999 3079 1005 3080
rect 999 3078 1000 3079
rect 827 3076 1000 3078
rect 827 3075 828 3076
rect 822 3074 828 3075
rect 999 3075 1000 3076
rect 1004 3075 1005 3079
rect 999 3074 1005 3075
rect 1050 3079 1056 3080
rect 1050 3075 1051 3079
rect 1055 3078 1056 3079
rect 1239 3079 1245 3080
rect 1239 3078 1240 3079
rect 1055 3076 1240 3078
rect 1055 3075 1056 3076
rect 1050 3074 1056 3075
rect 1239 3075 1240 3076
rect 1244 3075 1245 3079
rect 1239 3074 1245 3075
rect 1471 3079 1480 3080
rect 1471 3075 1472 3079
rect 1479 3075 1480 3079
rect 1471 3074 1480 3075
rect 1703 3079 1712 3080
rect 1703 3075 1704 3079
rect 1711 3075 1712 3079
rect 1703 3074 1712 3075
rect 1911 3079 1920 3080
rect 1911 3075 1912 3079
rect 1919 3075 1920 3079
rect 1911 3074 1920 3075
rect 1974 3077 1980 3078
rect 3798 3077 3804 3078
rect 1974 3073 1975 3077
rect 1979 3073 1980 3077
rect 110 3072 116 3073
rect 1934 3072 1940 3073
rect 1974 3072 1980 3073
rect 2646 3076 2652 3077
rect 2646 3072 2647 3076
rect 2651 3072 2652 3076
rect 110 3068 111 3072
rect 115 3068 116 3072
rect 110 3067 116 3068
rect 130 3071 136 3072
rect 130 3067 131 3071
rect 135 3067 136 3071
rect 130 3066 136 3067
rect 370 3071 376 3072
rect 370 3067 371 3071
rect 375 3067 376 3071
rect 370 3066 376 3067
rect 626 3071 632 3072
rect 626 3067 627 3071
rect 631 3067 632 3071
rect 626 3066 632 3067
rect 874 3071 880 3072
rect 874 3067 875 3071
rect 879 3067 880 3071
rect 874 3066 880 3067
rect 1114 3071 1120 3072
rect 1114 3067 1115 3071
rect 1119 3067 1120 3071
rect 1114 3066 1120 3067
rect 1346 3071 1352 3072
rect 1346 3067 1347 3071
rect 1351 3067 1352 3071
rect 1346 3066 1352 3067
rect 1578 3071 1584 3072
rect 1578 3067 1579 3071
rect 1583 3067 1584 3071
rect 1578 3066 1584 3067
rect 1786 3071 1792 3072
rect 1786 3067 1787 3071
rect 1791 3067 1792 3071
rect 1934 3068 1935 3072
rect 1939 3068 1940 3072
rect 2646 3071 2652 3072
rect 2782 3076 2788 3077
rect 2782 3072 2783 3076
rect 2787 3072 2788 3076
rect 2782 3071 2788 3072
rect 2926 3076 2932 3077
rect 2926 3072 2927 3076
rect 2931 3072 2932 3076
rect 2926 3071 2932 3072
rect 3078 3076 3084 3077
rect 3078 3072 3079 3076
rect 3083 3072 3084 3076
rect 3078 3071 3084 3072
rect 3238 3076 3244 3077
rect 3238 3072 3239 3076
rect 3243 3072 3244 3076
rect 3238 3071 3244 3072
rect 3398 3076 3404 3077
rect 3398 3072 3399 3076
rect 3403 3072 3404 3076
rect 3398 3071 3404 3072
rect 3566 3076 3572 3077
rect 3566 3072 3567 3076
rect 3571 3072 3572 3076
rect 3798 3073 3799 3077
rect 3803 3073 3804 3077
rect 3798 3072 3804 3073
rect 3566 3071 3572 3072
rect 1934 3067 1940 3068
rect 1786 3066 1792 3067
rect 2618 3061 2624 3062
rect 1974 3060 1980 3061
rect 158 3056 164 3057
rect 110 3055 116 3056
rect 110 3051 111 3055
rect 115 3051 116 3055
rect 158 3052 159 3056
rect 163 3052 164 3056
rect 158 3051 164 3052
rect 398 3056 404 3057
rect 398 3052 399 3056
rect 403 3052 404 3056
rect 398 3051 404 3052
rect 654 3056 660 3057
rect 654 3052 655 3056
rect 659 3052 660 3056
rect 654 3051 660 3052
rect 902 3056 908 3057
rect 902 3052 903 3056
rect 907 3052 908 3056
rect 902 3051 908 3052
rect 1142 3056 1148 3057
rect 1142 3052 1143 3056
rect 1147 3052 1148 3056
rect 1142 3051 1148 3052
rect 1374 3056 1380 3057
rect 1374 3052 1375 3056
rect 1379 3052 1380 3056
rect 1374 3051 1380 3052
rect 1606 3056 1612 3057
rect 1606 3052 1607 3056
rect 1611 3052 1612 3056
rect 1606 3051 1612 3052
rect 1814 3056 1820 3057
rect 1974 3056 1975 3060
rect 1979 3056 1980 3060
rect 2618 3057 2619 3061
rect 2623 3057 2624 3061
rect 2618 3056 2624 3057
rect 2754 3061 2760 3062
rect 2754 3057 2755 3061
rect 2759 3057 2760 3061
rect 2754 3056 2760 3057
rect 2898 3061 2904 3062
rect 2898 3057 2899 3061
rect 2903 3057 2904 3061
rect 2898 3056 2904 3057
rect 3050 3061 3056 3062
rect 3050 3057 3051 3061
rect 3055 3057 3056 3061
rect 3050 3056 3056 3057
rect 3210 3061 3216 3062
rect 3210 3057 3211 3061
rect 3215 3057 3216 3061
rect 3210 3056 3216 3057
rect 3370 3061 3376 3062
rect 3370 3057 3371 3061
rect 3375 3057 3376 3061
rect 3370 3056 3376 3057
rect 3538 3061 3544 3062
rect 3538 3057 3539 3061
rect 3543 3057 3544 3061
rect 3538 3056 3544 3057
rect 3798 3060 3804 3061
rect 3798 3056 3799 3060
rect 3803 3056 3804 3060
rect 1814 3052 1815 3056
rect 1819 3052 1820 3056
rect 1814 3051 1820 3052
rect 1934 3055 1940 3056
rect 1974 3055 1980 3056
rect 3798 3055 3804 3056
rect 1934 3051 1935 3055
rect 1939 3051 1940 3055
rect 110 3050 116 3051
rect 1934 3050 1940 3051
rect 2743 3051 2749 3052
rect 2743 3047 2744 3051
rect 2748 3050 2749 3051
rect 2770 3051 2776 3052
rect 2770 3050 2771 3051
rect 2748 3048 2771 3050
rect 2748 3047 2749 3048
rect 2743 3046 2749 3047
rect 2770 3047 2771 3048
rect 2775 3047 2776 3051
rect 2770 3046 2776 3047
rect 2879 3051 2885 3052
rect 2879 3047 2880 3051
rect 2884 3050 2885 3051
rect 2890 3051 2896 3052
rect 2890 3050 2891 3051
rect 2884 3048 2891 3050
rect 2884 3047 2885 3048
rect 2879 3046 2885 3047
rect 2890 3047 2891 3048
rect 2895 3047 2896 3051
rect 2890 3046 2896 3047
rect 3023 3051 3029 3052
rect 3023 3047 3024 3051
rect 3028 3050 3029 3051
rect 3066 3051 3072 3052
rect 3066 3050 3067 3051
rect 3028 3048 3067 3050
rect 3028 3047 3029 3048
rect 3023 3046 3029 3047
rect 3066 3047 3067 3048
rect 3071 3047 3072 3051
rect 3066 3046 3072 3047
rect 3175 3051 3181 3052
rect 3175 3047 3176 3051
rect 3180 3050 3181 3051
rect 3226 3051 3232 3052
rect 3226 3050 3227 3051
rect 3180 3048 3227 3050
rect 3180 3047 3181 3048
rect 3175 3046 3181 3047
rect 3226 3047 3227 3048
rect 3231 3047 3232 3051
rect 3335 3051 3341 3052
rect 3335 3050 3336 3051
rect 3226 3046 3232 3047
rect 3252 3048 3336 3050
rect 3199 3043 3205 3044
rect 3199 3039 3200 3043
rect 3204 3042 3205 3043
rect 3252 3042 3254 3048
rect 3335 3047 3336 3048
rect 3340 3047 3341 3051
rect 3335 3046 3341 3047
rect 3382 3051 3388 3052
rect 3382 3047 3383 3051
rect 3387 3050 3388 3051
rect 3495 3051 3501 3052
rect 3495 3050 3496 3051
rect 3387 3048 3496 3050
rect 3387 3047 3388 3048
rect 3382 3046 3388 3047
rect 3495 3047 3496 3048
rect 3500 3047 3501 3051
rect 3495 3046 3501 3047
rect 3526 3051 3532 3052
rect 3526 3047 3527 3051
rect 3531 3050 3532 3051
rect 3663 3051 3669 3052
rect 3663 3050 3664 3051
rect 3531 3048 3664 3050
rect 3531 3047 3532 3048
rect 3526 3046 3532 3047
rect 3663 3047 3664 3048
rect 3668 3047 3669 3051
rect 3663 3046 3669 3047
rect 3204 3040 3254 3042
rect 4358 3043 4364 3044
rect 3204 3039 3205 3040
rect 3199 3038 3205 3039
rect 4358 3039 4359 3043
rect 4363 3042 4364 3043
rect 5262 3043 5268 3044
rect 5262 3042 5263 3043
rect 4363 3040 5263 3042
rect 4363 3039 4364 3040
rect 4358 3038 4364 3039
rect 5262 3039 5263 3040
rect 5267 3039 5268 3043
rect 5262 3038 5268 3039
rect 3022 3035 3028 3036
rect 3022 3034 3023 3035
rect 2760 3032 3023 3034
rect 2760 3018 2762 3032
rect 3022 3031 3023 3032
rect 3027 3031 3028 3035
rect 3022 3030 3028 3031
rect 3838 3029 3844 3030
rect 5662 3029 5668 3030
rect 3838 3025 3839 3029
rect 3843 3025 3844 3029
rect 3838 3024 3844 3025
rect 4254 3028 4260 3029
rect 4254 3024 4255 3028
rect 4259 3024 4260 3028
rect 4254 3023 4260 3024
rect 4454 3028 4460 3029
rect 4454 3024 4455 3028
rect 4459 3024 4460 3028
rect 4454 3023 4460 3024
rect 4670 3028 4676 3029
rect 4670 3024 4671 3028
rect 4675 3024 4676 3028
rect 4670 3023 4676 3024
rect 4910 3028 4916 3029
rect 4910 3024 4911 3028
rect 4915 3024 4916 3028
rect 4910 3023 4916 3024
rect 5166 3028 5172 3029
rect 5166 3024 5167 3028
rect 5171 3024 5172 3028
rect 5166 3023 5172 3024
rect 5422 3028 5428 3029
rect 5422 3024 5423 3028
rect 5427 3024 5428 3028
rect 5662 3025 5663 3029
rect 5667 3025 5668 3029
rect 5662 3024 5668 3025
rect 5422 3023 5428 3024
rect 2709 3016 2762 3018
rect 2770 3019 2776 3020
rect 2770 3015 2771 3019
rect 2775 3015 2776 3019
rect 2770 3014 2776 3015
rect 2914 3019 2920 3020
rect 2914 3015 2915 3019
rect 2919 3015 2920 3019
rect 2914 3014 2920 3015
rect 3066 3019 3072 3020
rect 3066 3015 3067 3019
rect 3071 3015 3072 3019
rect 3066 3014 3072 3015
rect 3226 3019 3232 3020
rect 3226 3015 3227 3019
rect 3231 3015 3232 3019
rect 3526 3019 3532 3020
rect 3526 3018 3527 3019
rect 3461 3016 3527 3018
rect 3226 3014 3232 3015
rect 3526 3015 3527 3016
rect 3531 3015 3532 3019
rect 3526 3014 3532 3015
rect 3606 3019 3612 3020
rect 3606 3015 3607 3019
rect 3611 3015 3612 3019
rect 3606 3014 3612 3015
rect 4226 3013 4232 3014
rect 3838 3012 3844 3013
rect 1450 3011 1456 3012
rect 1450 3007 1451 3011
rect 1455 3010 1456 3011
rect 1910 3011 1916 3012
rect 1910 3010 1911 3011
rect 1455 3008 1911 3010
rect 1455 3007 1456 3008
rect 1450 3006 1456 3007
rect 1910 3007 1911 3008
rect 1915 3007 1916 3011
rect 3838 3008 3839 3012
rect 3843 3008 3844 3012
rect 4226 3009 4227 3013
rect 4231 3009 4232 3013
rect 4226 3008 4232 3009
rect 4426 3013 4432 3014
rect 4426 3009 4427 3013
rect 4431 3009 4432 3013
rect 4426 3008 4432 3009
rect 4642 3013 4648 3014
rect 4642 3009 4643 3013
rect 4647 3009 4648 3013
rect 4642 3008 4648 3009
rect 4882 3013 4888 3014
rect 4882 3009 4883 3013
rect 4887 3009 4888 3013
rect 4882 3008 4888 3009
rect 5138 3013 5144 3014
rect 5138 3009 5139 3013
rect 5143 3009 5144 3013
rect 5138 3008 5144 3009
rect 5394 3013 5400 3014
rect 5394 3009 5395 3013
rect 5399 3009 5400 3013
rect 5394 3008 5400 3009
rect 5662 3012 5668 3013
rect 5662 3008 5663 3012
rect 5667 3008 5668 3012
rect 3838 3007 3844 3008
rect 5662 3007 5668 3008
rect 1910 3006 1916 3007
rect 4351 3003 4357 3004
rect 4351 2999 4352 3003
rect 4356 3002 4357 3003
rect 4442 3003 4448 3004
rect 4442 3002 4443 3003
rect 4356 3000 4443 3002
rect 4356 2999 4357 3000
rect 4351 2998 4357 2999
rect 4442 2999 4443 3000
rect 4447 2999 4448 3003
rect 4442 2998 4448 2999
rect 4546 3003 4557 3004
rect 4546 2999 4547 3003
rect 4551 2999 4552 3003
rect 4556 2999 4557 3003
rect 4546 2998 4557 2999
rect 4767 3003 4773 3004
rect 4767 2999 4768 3003
rect 4772 3002 4773 3003
rect 4898 3003 4904 3004
rect 4898 3002 4899 3003
rect 4772 3000 4899 3002
rect 4772 2999 4773 3000
rect 4767 2998 4773 2999
rect 4898 2999 4899 3000
rect 4903 2999 4904 3003
rect 4898 2998 4904 2999
rect 5007 3003 5013 3004
rect 5007 2999 5008 3003
rect 5012 3002 5013 3003
rect 5154 3003 5160 3004
rect 5154 3002 5155 3003
rect 5012 3000 5155 3002
rect 5012 2999 5013 3000
rect 5007 2998 5013 2999
rect 5154 2999 5155 3000
rect 5159 2999 5160 3003
rect 5154 2998 5160 2999
rect 5262 3003 5269 3004
rect 5262 2999 5263 3003
rect 5268 2999 5269 3003
rect 5262 2998 5269 2999
rect 5362 3003 5368 3004
rect 5362 2999 5363 3003
rect 5367 3002 5368 3003
rect 5519 3003 5525 3004
rect 5519 3002 5520 3003
rect 5367 3000 5520 3002
rect 5367 2999 5368 3000
rect 5362 2998 5368 2999
rect 5519 2999 5520 3000
rect 5524 2999 5525 3003
rect 5519 2998 5525 2999
rect 110 2997 116 2998
rect 1934 2997 1940 2998
rect 110 2993 111 2997
rect 115 2993 116 2997
rect 110 2992 116 2993
rect 174 2996 180 2997
rect 174 2992 175 2996
rect 179 2992 180 2996
rect 174 2991 180 2992
rect 406 2996 412 2997
rect 406 2992 407 2996
rect 411 2992 412 2996
rect 406 2991 412 2992
rect 622 2996 628 2997
rect 622 2992 623 2996
rect 627 2992 628 2996
rect 622 2991 628 2992
rect 822 2996 828 2997
rect 822 2992 823 2996
rect 827 2992 828 2996
rect 822 2991 828 2992
rect 1006 2996 1012 2997
rect 1006 2992 1007 2996
rect 1011 2992 1012 2996
rect 1006 2991 1012 2992
rect 1182 2996 1188 2997
rect 1182 2992 1183 2996
rect 1187 2992 1188 2996
rect 1182 2991 1188 2992
rect 1350 2996 1356 2997
rect 1350 2992 1351 2996
rect 1355 2992 1356 2996
rect 1350 2991 1356 2992
rect 1510 2996 1516 2997
rect 1510 2992 1511 2996
rect 1515 2992 1516 2996
rect 1510 2991 1516 2992
rect 1670 2996 1676 2997
rect 1670 2992 1671 2996
rect 1675 2992 1676 2996
rect 1670 2991 1676 2992
rect 1814 2996 1820 2997
rect 1814 2992 1815 2996
rect 1819 2992 1820 2996
rect 1934 2993 1935 2997
rect 1939 2993 1940 2997
rect 1934 2992 1940 2993
rect 1814 2991 1820 2992
rect 146 2981 152 2982
rect 110 2980 116 2981
rect 110 2976 111 2980
rect 115 2976 116 2980
rect 146 2977 147 2981
rect 151 2977 152 2981
rect 146 2976 152 2977
rect 378 2981 384 2982
rect 378 2977 379 2981
rect 383 2977 384 2981
rect 378 2976 384 2977
rect 594 2981 600 2982
rect 594 2977 595 2981
rect 599 2977 600 2981
rect 594 2976 600 2977
rect 794 2981 800 2982
rect 794 2977 795 2981
rect 799 2977 800 2981
rect 794 2976 800 2977
rect 978 2981 984 2982
rect 978 2977 979 2981
rect 983 2977 984 2981
rect 978 2976 984 2977
rect 1154 2981 1160 2982
rect 1154 2977 1155 2981
rect 1159 2977 1160 2981
rect 1154 2976 1160 2977
rect 1322 2981 1328 2982
rect 1322 2977 1323 2981
rect 1327 2977 1328 2981
rect 1322 2976 1328 2977
rect 1482 2981 1488 2982
rect 1482 2977 1483 2981
rect 1487 2977 1488 2981
rect 1482 2976 1488 2977
rect 1642 2981 1648 2982
rect 1642 2977 1643 2981
rect 1647 2977 1648 2981
rect 1642 2976 1648 2977
rect 1786 2981 1792 2982
rect 1786 2977 1787 2981
rect 1791 2977 1792 2981
rect 1786 2976 1792 2977
rect 1934 2980 1940 2981
rect 1934 2976 1935 2980
rect 1939 2976 1940 2980
rect 110 2975 116 2976
rect 1934 2975 1940 2976
rect 271 2971 277 2972
rect 271 2967 272 2971
rect 276 2970 277 2971
rect 330 2971 336 2972
rect 330 2970 331 2971
rect 276 2968 331 2970
rect 276 2967 277 2968
rect 271 2966 277 2967
rect 330 2967 331 2968
rect 335 2967 336 2971
rect 330 2966 336 2967
rect 338 2971 344 2972
rect 338 2967 339 2971
rect 343 2970 344 2971
rect 503 2971 509 2972
rect 503 2970 504 2971
rect 343 2968 504 2970
rect 343 2967 344 2968
rect 338 2966 344 2967
rect 503 2967 504 2968
rect 508 2967 509 2971
rect 503 2966 509 2967
rect 719 2971 725 2972
rect 719 2967 720 2971
rect 724 2970 725 2971
rect 810 2971 816 2972
rect 810 2970 811 2971
rect 724 2968 811 2970
rect 724 2967 725 2968
rect 719 2966 725 2967
rect 810 2967 811 2968
rect 815 2967 816 2971
rect 810 2966 816 2967
rect 919 2971 925 2972
rect 919 2967 920 2971
rect 924 2970 925 2971
rect 994 2971 1000 2972
rect 994 2970 995 2971
rect 924 2968 995 2970
rect 924 2967 925 2968
rect 919 2966 925 2967
rect 994 2967 995 2968
rect 999 2967 1000 2971
rect 1103 2971 1109 2972
rect 1103 2970 1104 2971
rect 994 2966 1000 2967
rect 1004 2968 1104 2970
rect 906 2963 912 2964
rect 906 2959 907 2963
rect 911 2962 912 2963
rect 1004 2962 1006 2968
rect 1103 2967 1104 2968
rect 1108 2967 1109 2971
rect 1103 2966 1109 2967
rect 1279 2971 1285 2972
rect 1279 2967 1280 2971
rect 1284 2970 1285 2971
rect 1338 2971 1344 2972
rect 1338 2970 1339 2971
rect 1284 2968 1339 2970
rect 1284 2967 1285 2968
rect 1279 2966 1285 2967
rect 1338 2967 1339 2968
rect 1343 2967 1344 2971
rect 1338 2966 1344 2967
rect 1447 2971 1453 2972
rect 1447 2967 1448 2971
rect 1452 2970 1453 2971
rect 1498 2971 1504 2972
rect 1498 2970 1499 2971
rect 1452 2968 1499 2970
rect 1452 2967 1453 2968
rect 1447 2966 1453 2967
rect 1498 2967 1499 2968
rect 1503 2967 1504 2971
rect 1498 2966 1504 2967
rect 1607 2971 1613 2972
rect 1607 2967 1608 2971
rect 1612 2970 1613 2971
rect 1658 2971 1664 2972
rect 1658 2970 1659 2971
rect 1612 2968 1659 2970
rect 1612 2967 1613 2968
rect 1607 2966 1613 2967
rect 1658 2967 1659 2968
rect 1663 2967 1664 2971
rect 1658 2966 1664 2967
rect 1767 2971 1773 2972
rect 1767 2967 1768 2971
rect 1772 2970 1773 2971
rect 1802 2971 1808 2972
rect 1802 2970 1803 2971
rect 1772 2968 1803 2970
rect 1772 2967 1773 2968
rect 1767 2966 1773 2967
rect 1802 2967 1803 2968
rect 1807 2967 1808 2971
rect 1802 2966 1808 2967
rect 1910 2971 1917 2972
rect 1910 2967 1911 2971
rect 1916 2967 1917 2971
rect 2935 2971 2941 2972
rect 1910 2966 1917 2967
rect 2890 2967 2896 2968
rect 2890 2963 2891 2967
rect 2895 2963 2896 2967
rect 2935 2967 2936 2971
rect 2940 2970 2941 2971
rect 3199 2971 3205 2972
rect 3199 2970 3200 2971
rect 2940 2968 2957 2970
rect 3165 2968 3200 2970
rect 2940 2967 2941 2968
rect 2935 2966 2941 2967
rect 3199 2967 3200 2968
rect 3204 2967 3205 2971
rect 3199 2966 3205 2967
rect 3207 2971 3213 2972
rect 3207 2967 3208 2971
rect 3212 2970 3213 2971
rect 3343 2971 3349 2972
rect 3212 2968 3229 2970
rect 3212 2967 3213 2968
rect 3207 2966 3213 2967
rect 3343 2967 3344 2971
rect 3348 2970 3349 2971
rect 3479 2971 3485 2972
rect 3348 2968 3365 2970
rect 3348 2967 3349 2968
rect 3343 2966 3349 2967
rect 3479 2967 3480 2971
rect 3484 2970 3485 2971
rect 4358 2971 4364 2972
rect 4358 2970 4359 2971
rect 3484 2968 3501 2970
rect 4317 2968 4359 2970
rect 3484 2967 3485 2968
rect 3479 2966 3485 2967
rect 4358 2967 4359 2968
rect 4363 2967 4364 2971
rect 4358 2966 4364 2967
rect 4442 2971 4448 2972
rect 4442 2967 4443 2971
rect 4447 2967 4448 2971
rect 4442 2966 4448 2967
rect 4658 2971 4664 2972
rect 4658 2967 4659 2971
rect 4663 2967 4664 2971
rect 4658 2966 4664 2967
rect 4898 2971 4904 2972
rect 4898 2967 4899 2971
rect 4903 2967 4904 2971
rect 4898 2966 4904 2967
rect 5154 2971 5160 2972
rect 5154 2967 5155 2971
rect 5159 2967 5160 2971
rect 5154 2966 5160 2967
rect 5410 2971 5416 2972
rect 5410 2967 5411 2971
rect 5415 2967 5416 2971
rect 5410 2966 5416 2967
rect 2890 2962 2896 2963
rect 911 2960 1006 2962
rect 911 2959 912 2960
rect 906 2958 912 2959
rect 338 2939 344 2940
rect 338 2938 339 2939
rect 237 2936 339 2938
rect 338 2935 339 2936
rect 343 2935 344 2939
rect 338 2934 344 2935
rect 466 2939 472 2940
rect 466 2935 467 2939
rect 471 2935 472 2939
rect 466 2934 472 2935
rect 682 2939 688 2940
rect 682 2935 683 2939
rect 687 2935 688 2939
rect 682 2934 688 2935
rect 810 2939 816 2940
rect 810 2935 811 2939
rect 815 2935 816 2939
rect 810 2934 816 2935
rect 994 2939 1000 2940
rect 994 2935 995 2939
rect 999 2935 1000 2939
rect 1303 2939 1309 2940
rect 1303 2938 1304 2939
rect 1245 2936 1304 2938
rect 994 2934 1000 2935
rect 1303 2935 1304 2936
rect 1308 2935 1309 2939
rect 1303 2934 1309 2935
rect 1338 2939 1344 2940
rect 1338 2935 1339 2939
rect 1343 2935 1344 2939
rect 1338 2934 1344 2935
rect 1498 2939 1504 2940
rect 1498 2935 1499 2939
rect 1503 2935 1504 2939
rect 1498 2934 1504 2935
rect 1658 2939 1664 2940
rect 1658 2935 1659 2939
rect 1663 2935 1664 2939
rect 1658 2934 1664 2935
rect 1802 2939 1808 2940
rect 1802 2935 1803 2939
rect 1807 2935 1808 2939
rect 1802 2934 1808 2935
rect 2927 2935 2933 2936
rect 2927 2931 2928 2935
rect 2932 2934 2933 2935
rect 2935 2935 2941 2936
rect 2935 2934 2936 2935
rect 2932 2932 2936 2934
rect 2932 2931 2933 2932
rect 2927 2930 2933 2931
rect 2935 2931 2936 2932
rect 2940 2931 2941 2935
rect 2935 2930 2941 2931
rect 3058 2935 3069 2936
rect 3058 2931 3059 2935
rect 3063 2931 3064 2935
rect 3068 2931 3069 2935
rect 3058 2930 3069 2931
rect 3199 2935 3205 2936
rect 3199 2931 3200 2935
rect 3204 2934 3205 2935
rect 3207 2935 3213 2936
rect 3207 2934 3208 2935
rect 3204 2932 3208 2934
rect 3204 2931 3205 2932
rect 3199 2930 3205 2931
rect 3207 2931 3208 2932
rect 3212 2931 3213 2935
rect 3207 2930 3213 2931
rect 3335 2935 3341 2936
rect 3335 2931 3336 2935
rect 3340 2934 3341 2935
rect 3343 2935 3349 2936
rect 3343 2934 3344 2935
rect 3340 2932 3344 2934
rect 3340 2931 3341 2932
rect 3335 2930 3341 2931
rect 3343 2931 3344 2932
rect 3348 2931 3349 2935
rect 3343 2930 3349 2931
rect 3471 2935 3477 2936
rect 3471 2931 3472 2935
rect 3476 2934 3477 2935
rect 3479 2935 3485 2936
rect 3479 2934 3480 2935
rect 3476 2932 3480 2934
rect 3476 2931 3477 2932
rect 3471 2930 3477 2931
rect 3479 2931 3480 2932
rect 3484 2931 3485 2935
rect 3479 2930 3485 2931
rect 3606 2935 3613 2936
rect 3606 2931 3607 2935
rect 3612 2931 3613 2935
rect 3606 2930 3613 2931
rect 1974 2928 1980 2929
rect 3798 2928 3804 2929
rect 1974 2924 1975 2928
rect 1979 2924 1980 2928
rect 1974 2923 1980 2924
rect 2802 2927 2808 2928
rect 2802 2923 2803 2927
rect 2807 2923 2808 2927
rect 2802 2922 2808 2923
rect 2938 2927 2944 2928
rect 2938 2923 2939 2927
rect 2943 2923 2944 2927
rect 2938 2922 2944 2923
rect 3074 2927 3080 2928
rect 3074 2923 3075 2927
rect 3079 2923 3080 2927
rect 3074 2922 3080 2923
rect 3210 2927 3216 2928
rect 3210 2923 3211 2927
rect 3215 2923 3216 2927
rect 3210 2922 3216 2923
rect 3346 2927 3352 2928
rect 3346 2923 3347 2927
rect 3351 2923 3352 2927
rect 3346 2922 3352 2923
rect 3482 2927 3488 2928
rect 3482 2923 3483 2927
rect 3487 2923 3488 2927
rect 3798 2924 3799 2928
rect 3803 2924 3804 2928
rect 3798 2923 3804 2924
rect 3482 2922 3488 2923
rect 2830 2912 2836 2913
rect 1974 2911 1980 2912
rect 1974 2907 1975 2911
rect 1979 2907 1980 2911
rect 2830 2908 2831 2912
rect 2835 2908 2836 2912
rect 2830 2907 2836 2908
rect 2966 2912 2972 2913
rect 2966 2908 2967 2912
rect 2971 2908 2972 2912
rect 2966 2907 2972 2908
rect 3102 2912 3108 2913
rect 3102 2908 3103 2912
rect 3107 2908 3108 2912
rect 3102 2907 3108 2908
rect 3238 2912 3244 2913
rect 3238 2908 3239 2912
rect 3243 2908 3244 2912
rect 3238 2907 3244 2908
rect 3374 2912 3380 2913
rect 3374 2908 3375 2912
rect 3379 2908 3380 2912
rect 3374 2907 3380 2908
rect 3510 2912 3516 2913
rect 3510 2908 3511 2912
rect 3515 2908 3516 2912
rect 3510 2907 3516 2908
rect 3798 2911 3804 2912
rect 3798 2907 3799 2911
rect 3803 2907 3804 2911
rect 1974 2906 1980 2907
rect 3798 2906 3804 2907
rect 4174 2899 4180 2900
rect 4174 2898 4175 2899
rect 4085 2896 4175 2898
rect 4174 2895 4175 2896
rect 4179 2895 4180 2899
rect 4546 2899 4552 2900
rect 4546 2898 4547 2899
rect 4533 2896 4547 2898
rect 4174 2894 4180 2895
rect 4298 2895 4304 2896
rect 4298 2891 4299 2895
rect 4303 2891 4304 2895
rect 4546 2895 4547 2896
rect 4551 2895 4552 2899
rect 4546 2894 4552 2895
rect 4570 2899 4576 2900
rect 4570 2895 4571 2899
rect 4575 2898 4576 2899
rect 4826 2899 4832 2900
rect 4575 2896 4717 2898
rect 4575 2895 4576 2896
rect 4570 2894 4576 2895
rect 4826 2895 4827 2899
rect 4831 2898 4832 2899
rect 5618 2899 5624 2900
rect 5618 2898 5619 2899
rect 4831 2896 4989 2898
rect 5605 2896 5619 2898
rect 4831 2895 4832 2896
rect 4826 2894 4832 2895
rect 5338 2895 5344 2896
rect 4298 2890 4304 2891
rect 5338 2891 5339 2895
rect 5343 2891 5344 2895
rect 5618 2895 5619 2896
rect 5623 2895 5624 2899
rect 5618 2894 5624 2895
rect 5338 2890 5344 2891
rect 527 2887 533 2888
rect 527 2886 528 2887
rect 485 2884 528 2886
rect 527 2883 528 2884
rect 532 2883 533 2887
rect 906 2887 912 2888
rect 906 2886 907 2887
rect 877 2884 907 2886
rect 527 2882 533 2883
rect 682 2883 688 2884
rect 682 2879 683 2883
rect 687 2879 688 2883
rect 906 2883 907 2884
rect 911 2883 912 2887
rect 906 2882 912 2883
rect 914 2887 920 2888
rect 914 2883 915 2887
rect 919 2886 920 2887
rect 1098 2887 1104 2888
rect 919 2884 989 2886
rect 919 2883 920 2884
rect 914 2882 920 2883
rect 1098 2883 1099 2887
rect 1103 2886 1104 2887
rect 1479 2887 1485 2888
rect 1479 2886 1480 2887
rect 1103 2884 1165 2886
rect 1405 2884 1480 2886
rect 1103 2883 1104 2884
rect 1098 2882 1104 2883
rect 1479 2883 1480 2884
rect 1484 2883 1485 2887
rect 1631 2887 1637 2888
rect 1631 2886 1632 2887
rect 1573 2884 1632 2886
rect 1479 2882 1485 2883
rect 1631 2883 1632 2884
rect 1636 2883 1637 2887
rect 1783 2887 1789 2888
rect 1783 2886 1784 2887
rect 1733 2884 1784 2886
rect 1631 2882 1637 2883
rect 1783 2883 1784 2884
rect 1788 2883 1789 2887
rect 1783 2882 1789 2883
rect 1874 2883 1880 2884
rect 682 2878 688 2879
rect 1874 2879 1875 2883
rect 1879 2879 1880 2883
rect 1874 2878 1880 2879
rect 4298 2871 4304 2872
rect 4298 2867 4299 2871
rect 4303 2870 4304 2871
rect 4303 2868 4962 2870
rect 4303 2867 4304 2868
rect 4298 2866 4304 2867
rect 3978 2863 3984 2864
rect 3978 2859 3979 2863
rect 3983 2862 3984 2863
rect 4119 2863 4125 2864
rect 4119 2862 4120 2863
rect 3983 2860 4120 2862
rect 3983 2859 3984 2860
rect 3978 2858 3984 2859
rect 4119 2859 4120 2860
rect 4124 2859 4125 2863
rect 4119 2858 4125 2859
rect 4174 2863 4180 2864
rect 4174 2859 4175 2863
rect 4179 2862 4180 2863
rect 4335 2863 4341 2864
rect 4335 2862 4336 2863
rect 4179 2860 4336 2862
rect 4179 2859 4180 2860
rect 4174 2858 4180 2859
rect 4335 2859 4336 2860
rect 4340 2859 4341 2863
rect 4335 2858 4341 2859
rect 4567 2863 4576 2864
rect 4567 2859 4568 2863
rect 4575 2859 4576 2863
rect 4567 2858 4576 2859
rect 4823 2863 4832 2864
rect 4823 2859 4824 2863
rect 4831 2859 4832 2863
rect 4960 2862 4962 2868
rect 5095 2863 5101 2864
rect 5095 2862 5096 2863
rect 4960 2860 5096 2862
rect 4823 2858 4832 2859
rect 5095 2859 5096 2860
rect 5100 2859 5101 2863
rect 5095 2858 5101 2859
rect 5375 2863 5381 2864
rect 5375 2859 5376 2863
rect 5380 2862 5381 2863
rect 5410 2863 5416 2864
rect 5410 2862 5411 2863
rect 5380 2860 5411 2862
rect 5380 2859 5381 2860
rect 5375 2858 5381 2859
rect 5410 2859 5411 2860
rect 5415 2859 5416 2863
rect 5410 2858 5416 2859
rect 5618 2863 5624 2864
rect 5618 2859 5619 2863
rect 5623 2862 5624 2863
rect 5639 2863 5645 2864
rect 5639 2862 5640 2863
rect 5623 2860 5640 2862
rect 5623 2859 5624 2860
rect 5618 2858 5624 2859
rect 5639 2859 5640 2860
rect 5644 2859 5645 2863
rect 5639 2858 5645 2859
rect 3838 2856 3844 2857
rect 5662 2856 5668 2857
rect 3838 2852 3839 2856
rect 3843 2852 3844 2856
rect 466 2851 472 2852
rect 466 2847 467 2851
rect 471 2850 472 2851
rect 519 2851 525 2852
rect 519 2850 520 2851
rect 471 2848 520 2850
rect 471 2847 472 2848
rect 466 2846 472 2847
rect 519 2847 520 2848
rect 524 2847 525 2851
rect 519 2846 525 2847
rect 527 2851 533 2852
rect 527 2847 528 2851
rect 532 2850 533 2851
rect 719 2851 725 2852
rect 719 2850 720 2851
rect 532 2848 720 2850
rect 532 2847 533 2848
rect 527 2846 533 2847
rect 719 2847 720 2848
rect 724 2847 725 2851
rect 719 2846 725 2847
rect 911 2851 920 2852
rect 911 2847 912 2851
rect 919 2847 920 2851
rect 911 2846 920 2847
rect 1095 2851 1104 2852
rect 1095 2847 1096 2851
rect 1103 2847 1104 2851
rect 1095 2846 1104 2847
rect 1202 2851 1208 2852
rect 1202 2847 1203 2851
rect 1207 2850 1208 2851
rect 1271 2851 1277 2852
rect 1271 2850 1272 2851
rect 1207 2848 1272 2850
rect 1207 2847 1208 2848
rect 1202 2846 1208 2847
rect 1271 2847 1272 2848
rect 1276 2847 1277 2851
rect 1271 2846 1277 2847
rect 1303 2851 1309 2852
rect 1303 2847 1304 2851
rect 1308 2850 1309 2851
rect 1439 2851 1445 2852
rect 1439 2850 1440 2851
rect 1308 2848 1440 2850
rect 1308 2847 1309 2848
rect 1303 2846 1309 2847
rect 1439 2847 1440 2848
rect 1444 2847 1445 2851
rect 1439 2846 1445 2847
rect 1479 2851 1485 2852
rect 1479 2847 1480 2851
rect 1484 2850 1485 2851
rect 1607 2851 1613 2852
rect 1607 2850 1608 2851
rect 1484 2848 1608 2850
rect 1484 2847 1485 2848
rect 1479 2846 1485 2847
rect 1607 2847 1608 2848
rect 1612 2847 1613 2851
rect 1607 2846 1613 2847
rect 1631 2851 1637 2852
rect 1631 2847 1632 2851
rect 1636 2850 1637 2851
rect 1767 2851 1773 2852
rect 1767 2850 1768 2851
rect 1636 2848 1768 2850
rect 1636 2847 1637 2848
rect 1631 2846 1637 2847
rect 1767 2847 1768 2848
rect 1772 2847 1773 2851
rect 1767 2846 1773 2847
rect 1783 2851 1789 2852
rect 1783 2847 1784 2851
rect 1788 2850 1789 2851
rect 1911 2851 1917 2852
rect 3838 2851 3844 2852
rect 3994 2855 4000 2856
rect 3994 2851 3995 2855
rect 3999 2851 4000 2855
rect 1911 2850 1912 2851
rect 1788 2848 1912 2850
rect 1788 2847 1789 2848
rect 1783 2846 1789 2847
rect 1911 2847 1912 2848
rect 1916 2847 1917 2851
rect 3994 2850 4000 2851
rect 4210 2855 4216 2856
rect 4210 2851 4211 2855
rect 4215 2851 4216 2855
rect 4210 2850 4216 2851
rect 4442 2855 4448 2856
rect 4442 2851 4443 2855
rect 4447 2851 4448 2855
rect 4442 2850 4448 2851
rect 4698 2855 4704 2856
rect 4698 2851 4699 2855
rect 4703 2851 4704 2855
rect 4698 2850 4704 2851
rect 4970 2855 4976 2856
rect 4970 2851 4971 2855
rect 4975 2851 4976 2855
rect 4970 2850 4976 2851
rect 5250 2855 5256 2856
rect 5250 2851 5251 2855
rect 5255 2851 5256 2855
rect 5250 2850 5256 2851
rect 5514 2855 5520 2856
rect 5514 2851 5515 2855
rect 5519 2851 5520 2855
rect 5662 2852 5663 2856
rect 5667 2852 5668 2856
rect 5662 2851 5668 2852
rect 5514 2850 5520 2851
rect 1911 2846 1917 2847
rect 110 2844 116 2845
rect 1934 2844 1940 2845
rect 110 2840 111 2844
rect 115 2840 116 2844
rect 110 2839 116 2840
rect 394 2843 400 2844
rect 394 2839 395 2843
rect 399 2839 400 2843
rect 394 2838 400 2839
rect 594 2843 600 2844
rect 594 2839 595 2843
rect 599 2839 600 2843
rect 594 2838 600 2839
rect 786 2843 792 2844
rect 786 2839 787 2843
rect 791 2839 792 2843
rect 786 2838 792 2839
rect 970 2843 976 2844
rect 970 2839 971 2843
rect 975 2839 976 2843
rect 970 2838 976 2839
rect 1146 2843 1152 2844
rect 1146 2839 1147 2843
rect 1151 2839 1152 2843
rect 1146 2838 1152 2839
rect 1314 2843 1320 2844
rect 1314 2839 1315 2843
rect 1319 2839 1320 2843
rect 1314 2838 1320 2839
rect 1482 2843 1488 2844
rect 1482 2839 1483 2843
rect 1487 2839 1488 2843
rect 1482 2838 1488 2839
rect 1642 2843 1648 2844
rect 1642 2839 1643 2843
rect 1647 2839 1648 2843
rect 1642 2838 1648 2839
rect 1786 2843 1792 2844
rect 1786 2839 1787 2843
rect 1791 2839 1792 2843
rect 1934 2840 1935 2844
rect 1939 2840 1940 2844
rect 4022 2840 4028 2841
rect 1934 2839 1940 2840
rect 3838 2839 3844 2840
rect 1786 2838 1792 2839
rect 3838 2835 3839 2839
rect 3843 2835 3844 2839
rect 4022 2836 4023 2840
rect 4027 2836 4028 2840
rect 4022 2835 4028 2836
rect 4238 2840 4244 2841
rect 4238 2836 4239 2840
rect 4243 2836 4244 2840
rect 4238 2835 4244 2836
rect 4470 2840 4476 2841
rect 4470 2836 4471 2840
rect 4475 2836 4476 2840
rect 4470 2835 4476 2836
rect 4726 2840 4732 2841
rect 4726 2836 4727 2840
rect 4731 2836 4732 2840
rect 4726 2835 4732 2836
rect 4998 2840 5004 2841
rect 4998 2836 4999 2840
rect 5003 2836 5004 2840
rect 4998 2835 5004 2836
rect 5278 2840 5284 2841
rect 5278 2836 5279 2840
rect 5283 2836 5284 2840
rect 5278 2835 5284 2836
rect 5542 2840 5548 2841
rect 5542 2836 5543 2840
rect 5547 2836 5548 2840
rect 5542 2835 5548 2836
rect 5662 2839 5668 2840
rect 5662 2835 5663 2839
rect 5667 2835 5668 2839
rect 3838 2834 3844 2835
rect 5662 2834 5668 2835
rect 422 2828 428 2829
rect 110 2827 116 2828
rect 110 2823 111 2827
rect 115 2823 116 2827
rect 422 2824 423 2828
rect 427 2824 428 2828
rect 422 2823 428 2824
rect 622 2828 628 2829
rect 622 2824 623 2828
rect 627 2824 628 2828
rect 622 2823 628 2824
rect 814 2828 820 2829
rect 814 2824 815 2828
rect 819 2824 820 2828
rect 814 2823 820 2824
rect 998 2828 1004 2829
rect 998 2824 999 2828
rect 1003 2824 1004 2828
rect 998 2823 1004 2824
rect 1174 2828 1180 2829
rect 1174 2824 1175 2828
rect 1179 2824 1180 2828
rect 1174 2823 1180 2824
rect 1342 2828 1348 2829
rect 1342 2824 1343 2828
rect 1347 2824 1348 2828
rect 1342 2823 1348 2824
rect 1510 2828 1516 2829
rect 1510 2824 1511 2828
rect 1515 2824 1516 2828
rect 1510 2823 1516 2824
rect 1670 2828 1676 2829
rect 1670 2824 1671 2828
rect 1675 2824 1676 2828
rect 1670 2823 1676 2824
rect 1814 2828 1820 2829
rect 1814 2824 1815 2828
rect 1819 2824 1820 2828
rect 1814 2823 1820 2824
rect 1934 2827 1940 2828
rect 1934 2823 1935 2827
rect 1939 2823 1940 2827
rect 110 2822 116 2823
rect 1934 2822 1940 2823
rect 1974 2801 1980 2802
rect 3798 2801 3804 2802
rect 1974 2797 1975 2801
rect 1979 2797 1980 2801
rect 1974 2796 1980 2797
rect 2022 2800 2028 2801
rect 2022 2796 2023 2800
rect 2027 2796 2028 2800
rect 2022 2795 2028 2796
rect 2166 2800 2172 2801
rect 2166 2796 2167 2800
rect 2171 2796 2172 2800
rect 2166 2795 2172 2796
rect 2334 2800 2340 2801
rect 2334 2796 2335 2800
rect 2339 2796 2340 2800
rect 2334 2795 2340 2796
rect 2494 2800 2500 2801
rect 2494 2796 2495 2800
rect 2499 2796 2500 2800
rect 2494 2795 2500 2796
rect 2662 2800 2668 2801
rect 2662 2796 2663 2800
rect 2667 2796 2668 2800
rect 2662 2795 2668 2796
rect 2830 2800 2836 2801
rect 2830 2796 2831 2800
rect 2835 2796 2836 2800
rect 2830 2795 2836 2796
rect 2998 2800 3004 2801
rect 2998 2796 2999 2800
rect 3003 2796 3004 2800
rect 2998 2795 3004 2796
rect 3166 2800 3172 2801
rect 3166 2796 3167 2800
rect 3171 2796 3172 2800
rect 3798 2797 3799 2801
rect 3803 2797 3804 2801
rect 3798 2796 3804 2797
rect 3166 2795 3172 2796
rect 1994 2785 2000 2786
rect 1974 2784 1980 2785
rect 1974 2780 1975 2784
rect 1979 2780 1980 2784
rect 1994 2781 1995 2785
rect 1999 2781 2000 2785
rect 1994 2780 2000 2781
rect 2138 2785 2144 2786
rect 2138 2781 2139 2785
rect 2143 2781 2144 2785
rect 2138 2780 2144 2781
rect 2306 2785 2312 2786
rect 2306 2781 2307 2785
rect 2311 2781 2312 2785
rect 2306 2780 2312 2781
rect 2466 2785 2472 2786
rect 2466 2781 2467 2785
rect 2471 2781 2472 2785
rect 2466 2780 2472 2781
rect 2634 2785 2640 2786
rect 2634 2781 2635 2785
rect 2639 2781 2640 2785
rect 2634 2780 2640 2781
rect 2802 2785 2808 2786
rect 2802 2781 2803 2785
rect 2807 2781 2808 2785
rect 2802 2780 2808 2781
rect 2970 2785 2976 2786
rect 2970 2781 2971 2785
rect 2975 2781 2976 2785
rect 2970 2780 2976 2781
rect 3138 2785 3144 2786
rect 3138 2781 3139 2785
rect 3143 2781 3144 2785
rect 3138 2780 3144 2781
rect 3798 2784 3804 2785
rect 3798 2780 3799 2784
rect 3803 2780 3804 2784
rect 1974 2779 1980 2780
rect 3798 2779 3804 2780
rect 3838 2777 3844 2778
rect 5662 2777 5668 2778
rect 1874 2775 1880 2776
rect 1874 2771 1875 2775
rect 1879 2774 1880 2775
rect 2119 2775 2125 2776
rect 2119 2774 2120 2775
rect 1879 2772 2120 2774
rect 1879 2771 1880 2772
rect 1874 2770 1880 2771
rect 2119 2771 2120 2772
rect 2124 2771 2125 2775
rect 2119 2770 2125 2771
rect 2135 2775 2141 2776
rect 2135 2771 2136 2775
rect 2140 2774 2141 2775
rect 2263 2775 2269 2776
rect 2263 2774 2264 2775
rect 2140 2772 2264 2774
rect 2140 2771 2141 2772
rect 2135 2770 2141 2771
rect 2263 2771 2264 2772
rect 2268 2771 2269 2775
rect 2263 2770 2269 2771
rect 2271 2775 2277 2776
rect 2271 2771 2272 2775
rect 2276 2774 2277 2775
rect 2431 2775 2437 2776
rect 2431 2774 2432 2775
rect 2276 2772 2432 2774
rect 2276 2771 2277 2772
rect 2271 2770 2277 2771
rect 2431 2771 2432 2772
rect 2436 2771 2437 2775
rect 2431 2770 2437 2771
rect 2455 2775 2461 2776
rect 2455 2771 2456 2775
rect 2460 2774 2461 2775
rect 2591 2775 2597 2776
rect 2591 2774 2592 2775
rect 2460 2772 2592 2774
rect 2460 2771 2461 2772
rect 2455 2770 2461 2771
rect 2591 2771 2592 2772
rect 2596 2771 2597 2775
rect 2591 2770 2597 2771
rect 2746 2775 2752 2776
rect 2746 2771 2747 2775
rect 2751 2774 2752 2775
rect 2759 2775 2765 2776
rect 2759 2774 2760 2775
rect 2751 2772 2760 2774
rect 2751 2771 2752 2772
rect 2746 2770 2752 2771
rect 2759 2771 2760 2772
rect 2764 2771 2765 2775
rect 2759 2770 2765 2771
rect 2790 2775 2796 2776
rect 2790 2771 2791 2775
rect 2795 2774 2796 2775
rect 2927 2775 2933 2776
rect 2927 2774 2928 2775
rect 2795 2772 2928 2774
rect 2795 2771 2796 2772
rect 2790 2770 2796 2771
rect 2927 2771 2928 2772
rect 2932 2771 2933 2775
rect 2927 2770 2933 2771
rect 3095 2775 3101 2776
rect 3095 2771 3096 2775
rect 3100 2774 3101 2775
rect 3154 2775 3160 2776
rect 3154 2774 3155 2775
rect 3100 2772 3155 2774
rect 3100 2771 3101 2772
rect 3095 2770 3101 2771
rect 3154 2771 3155 2772
rect 3159 2771 3160 2775
rect 3263 2775 3269 2776
rect 3263 2774 3264 2775
rect 3154 2770 3160 2771
rect 3200 2772 3264 2774
rect 2890 2767 2896 2768
rect 2890 2763 2891 2767
rect 2895 2766 2896 2767
rect 3200 2766 3202 2772
rect 3263 2771 3264 2772
rect 3268 2771 3269 2775
rect 3838 2773 3839 2777
rect 3843 2773 3844 2777
rect 3838 2772 3844 2773
rect 3918 2776 3924 2777
rect 3918 2772 3919 2776
rect 3923 2772 3924 2776
rect 3918 2771 3924 2772
rect 4054 2776 4060 2777
rect 4054 2772 4055 2776
rect 4059 2772 4060 2776
rect 4054 2771 4060 2772
rect 4190 2776 4196 2777
rect 4190 2772 4191 2776
rect 4195 2772 4196 2776
rect 4190 2771 4196 2772
rect 4326 2776 4332 2777
rect 4326 2772 4327 2776
rect 4331 2772 4332 2776
rect 4326 2771 4332 2772
rect 4462 2776 4468 2777
rect 4462 2772 4463 2776
rect 4467 2772 4468 2776
rect 5662 2773 5663 2777
rect 5667 2773 5668 2777
rect 5662 2772 5668 2773
rect 4462 2771 4468 2772
rect 3263 2770 3269 2771
rect 2895 2764 3202 2766
rect 2895 2763 2896 2764
rect 2890 2762 2896 2763
rect 3890 2761 3896 2762
rect 3838 2760 3844 2761
rect 110 2757 116 2758
rect 1934 2757 1940 2758
rect 110 2753 111 2757
rect 115 2753 116 2757
rect 110 2752 116 2753
rect 654 2756 660 2757
rect 654 2752 655 2756
rect 659 2752 660 2756
rect 654 2751 660 2752
rect 814 2756 820 2757
rect 814 2752 815 2756
rect 819 2752 820 2756
rect 814 2751 820 2752
rect 974 2756 980 2757
rect 974 2752 975 2756
rect 979 2752 980 2756
rect 974 2751 980 2752
rect 1142 2756 1148 2757
rect 1142 2752 1143 2756
rect 1147 2752 1148 2756
rect 1142 2751 1148 2752
rect 1310 2756 1316 2757
rect 1310 2752 1311 2756
rect 1315 2752 1316 2756
rect 1310 2751 1316 2752
rect 1478 2756 1484 2757
rect 1478 2752 1479 2756
rect 1483 2752 1484 2756
rect 1934 2753 1935 2757
rect 1939 2753 1940 2757
rect 3838 2756 3839 2760
rect 3843 2756 3844 2760
rect 3890 2757 3891 2761
rect 3895 2757 3896 2761
rect 3890 2756 3896 2757
rect 4026 2761 4032 2762
rect 4026 2757 4027 2761
rect 4031 2757 4032 2761
rect 4026 2756 4032 2757
rect 4162 2761 4168 2762
rect 4162 2757 4163 2761
rect 4167 2757 4168 2761
rect 4162 2756 4168 2757
rect 4298 2761 4304 2762
rect 4298 2757 4299 2761
rect 4303 2757 4304 2761
rect 4298 2756 4304 2757
rect 4434 2761 4440 2762
rect 4434 2757 4435 2761
rect 4439 2757 4440 2761
rect 4434 2756 4440 2757
rect 5662 2760 5668 2761
rect 5662 2756 5663 2760
rect 5667 2756 5668 2760
rect 3838 2755 3844 2756
rect 5662 2755 5668 2756
rect 1934 2752 1940 2753
rect 1478 2751 1484 2752
rect 4015 2751 4021 2752
rect 4015 2747 4016 2751
rect 4020 2750 4021 2751
rect 4042 2751 4048 2752
rect 4042 2750 4043 2751
rect 4020 2748 4043 2750
rect 4020 2747 4021 2748
rect 4015 2746 4021 2747
rect 4042 2747 4043 2748
rect 4047 2747 4048 2751
rect 4042 2746 4048 2747
rect 4151 2751 4157 2752
rect 4151 2747 4152 2751
rect 4156 2750 4157 2751
rect 4178 2751 4184 2752
rect 4178 2750 4179 2751
rect 4156 2748 4179 2750
rect 4156 2747 4157 2748
rect 4151 2746 4157 2747
rect 4178 2747 4179 2748
rect 4183 2747 4184 2751
rect 4178 2746 4184 2747
rect 4287 2751 4293 2752
rect 4287 2747 4288 2751
rect 4292 2750 4293 2751
rect 4314 2751 4320 2752
rect 4314 2750 4315 2751
rect 4292 2748 4315 2750
rect 4292 2747 4293 2748
rect 4287 2746 4293 2747
rect 4314 2747 4315 2748
rect 4319 2747 4320 2751
rect 4314 2746 4320 2747
rect 4423 2751 4429 2752
rect 4423 2747 4424 2751
rect 4428 2750 4429 2751
rect 4450 2751 4456 2752
rect 4450 2750 4451 2751
rect 4428 2748 4451 2750
rect 4428 2747 4429 2748
rect 4423 2746 4429 2747
rect 4450 2747 4451 2748
rect 4455 2747 4456 2751
rect 4559 2751 4565 2752
rect 4559 2750 4560 2751
rect 4450 2746 4456 2747
rect 4460 2748 4560 2750
rect 2135 2743 2141 2744
rect 2135 2742 2136 2743
rect 626 2741 632 2742
rect 110 2740 116 2741
rect 110 2736 111 2740
rect 115 2736 116 2740
rect 626 2737 627 2741
rect 631 2737 632 2741
rect 626 2736 632 2737
rect 786 2741 792 2742
rect 786 2737 787 2741
rect 791 2737 792 2741
rect 786 2736 792 2737
rect 946 2741 952 2742
rect 946 2737 947 2741
rect 951 2737 952 2741
rect 946 2736 952 2737
rect 1114 2741 1120 2742
rect 1114 2737 1115 2741
rect 1119 2737 1120 2741
rect 1114 2736 1120 2737
rect 1282 2741 1288 2742
rect 1282 2737 1283 2741
rect 1287 2737 1288 2741
rect 1282 2736 1288 2737
rect 1450 2741 1456 2742
rect 1450 2737 1451 2741
rect 1455 2737 1456 2741
rect 1450 2736 1456 2737
rect 1934 2740 1940 2741
rect 2085 2740 2136 2742
rect 1934 2736 1935 2740
rect 1939 2736 1940 2740
rect 2135 2739 2136 2740
rect 2140 2739 2141 2743
rect 2271 2743 2277 2744
rect 2271 2742 2272 2743
rect 2229 2740 2272 2742
rect 2135 2738 2141 2739
rect 2271 2739 2272 2740
rect 2276 2739 2277 2743
rect 2455 2743 2461 2744
rect 2455 2742 2456 2743
rect 2397 2740 2456 2742
rect 2271 2738 2277 2739
rect 2455 2739 2456 2740
rect 2460 2739 2461 2743
rect 2455 2738 2461 2739
rect 2502 2743 2508 2744
rect 2502 2739 2503 2743
rect 2507 2739 2508 2743
rect 2790 2743 2796 2744
rect 2790 2742 2791 2743
rect 2725 2740 2791 2742
rect 2502 2738 2508 2739
rect 2790 2739 2791 2740
rect 2795 2739 2796 2743
rect 2790 2738 2796 2739
rect 2890 2743 2896 2744
rect 2890 2739 2891 2743
rect 2895 2739 2896 2743
rect 2890 2738 2896 2739
rect 3058 2743 3064 2744
rect 3058 2739 3059 2743
rect 3063 2739 3064 2743
rect 3058 2738 3064 2739
rect 3154 2743 3160 2744
rect 3154 2739 3155 2743
rect 3159 2739 3160 2743
rect 3154 2738 3160 2739
rect 4218 2743 4224 2744
rect 4218 2739 4219 2743
rect 4223 2742 4224 2743
rect 4460 2742 4462 2748
rect 4559 2747 4560 2748
rect 4564 2747 4565 2751
rect 4559 2746 4565 2747
rect 4223 2740 4462 2742
rect 4223 2739 4224 2740
rect 4218 2738 4224 2739
rect 110 2735 116 2736
rect 1934 2735 1940 2736
rect 682 2731 688 2732
rect 682 2727 683 2731
rect 687 2730 688 2731
rect 751 2731 757 2732
rect 751 2730 752 2731
rect 687 2728 752 2730
rect 687 2727 688 2728
rect 682 2726 688 2727
rect 751 2727 752 2728
rect 756 2727 757 2731
rect 751 2726 757 2727
rect 775 2731 781 2732
rect 775 2727 776 2731
rect 780 2730 781 2731
rect 911 2731 917 2732
rect 911 2730 912 2731
rect 780 2728 912 2730
rect 780 2727 781 2728
rect 775 2726 781 2727
rect 911 2727 912 2728
rect 916 2727 917 2731
rect 911 2726 917 2727
rect 935 2731 941 2732
rect 935 2727 936 2731
rect 940 2730 941 2731
rect 1071 2731 1077 2732
rect 1071 2730 1072 2731
rect 940 2728 1072 2730
rect 940 2727 941 2728
rect 935 2726 941 2727
rect 1071 2727 1072 2728
rect 1076 2727 1077 2731
rect 1071 2726 1077 2727
rect 1239 2731 1245 2732
rect 1239 2727 1240 2731
rect 1244 2730 1245 2731
rect 1298 2731 1304 2732
rect 1298 2730 1299 2731
rect 1244 2728 1299 2730
rect 1244 2727 1245 2728
rect 1239 2726 1245 2727
rect 1298 2727 1299 2728
rect 1303 2727 1304 2731
rect 1298 2726 1304 2727
rect 1407 2731 1413 2732
rect 1407 2727 1408 2731
rect 1412 2730 1413 2731
rect 1466 2731 1472 2732
rect 1466 2730 1467 2731
rect 1412 2728 1467 2730
rect 1412 2727 1413 2728
rect 1407 2726 1413 2727
rect 1466 2727 1467 2728
rect 1471 2727 1472 2731
rect 1466 2726 1472 2727
rect 1554 2731 1560 2732
rect 1554 2727 1555 2731
rect 1559 2730 1560 2731
rect 1575 2731 1581 2732
rect 1575 2730 1576 2731
rect 1559 2728 1576 2730
rect 1559 2727 1560 2728
rect 1554 2726 1560 2727
rect 1575 2727 1576 2728
rect 1580 2727 1581 2731
rect 1575 2726 1581 2727
rect 3978 2719 3984 2720
rect 3978 2715 3979 2719
rect 3983 2715 3984 2719
rect 3978 2714 3984 2715
rect 4042 2719 4048 2720
rect 4042 2715 4043 2719
rect 4047 2715 4048 2719
rect 4042 2714 4048 2715
rect 4178 2719 4184 2720
rect 4178 2715 4179 2719
rect 4183 2715 4184 2719
rect 4178 2714 4184 2715
rect 4314 2719 4320 2720
rect 4314 2715 4315 2719
rect 4319 2715 4320 2719
rect 4314 2714 4320 2715
rect 4450 2719 4456 2720
rect 4450 2715 4451 2719
rect 4455 2715 4456 2719
rect 4450 2714 4456 2715
rect 775 2699 781 2700
rect 775 2698 776 2699
rect 717 2696 776 2698
rect 775 2695 776 2696
rect 780 2695 781 2699
rect 935 2699 941 2700
rect 935 2698 936 2699
rect 877 2696 936 2698
rect 775 2694 781 2695
rect 935 2695 936 2696
rect 940 2695 941 2699
rect 935 2694 941 2695
rect 1030 2699 1036 2700
rect 1030 2695 1031 2699
rect 1035 2695 1036 2699
rect 1030 2694 1036 2695
rect 1202 2699 1208 2700
rect 1202 2695 1203 2699
rect 1207 2695 1208 2699
rect 1202 2694 1208 2695
rect 1298 2699 1304 2700
rect 1298 2695 1299 2699
rect 1303 2695 1304 2699
rect 1298 2694 1304 2695
rect 1466 2699 1472 2700
rect 1466 2695 1467 2699
rect 1471 2695 1472 2699
rect 1466 2694 1472 2695
rect 2511 2695 2517 2696
rect 2511 2694 2512 2695
rect 2469 2692 2512 2694
rect 2511 2691 2512 2692
rect 2516 2691 2517 2695
rect 2786 2695 2792 2696
rect 2511 2690 2517 2691
rect 2602 2691 2608 2692
rect 2602 2687 2603 2691
rect 2607 2687 2608 2691
rect 2602 2686 2608 2687
rect 2746 2691 2752 2692
rect 2746 2687 2747 2691
rect 2751 2687 2752 2691
rect 2786 2691 2787 2695
rect 2791 2694 2792 2695
rect 2930 2695 2936 2696
rect 2791 2692 2821 2694
rect 2791 2691 2792 2692
rect 2786 2690 2792 2691
rect 2930 2691 2931 2695
rect 2935 2694 2936 2695
rect 3074 2695 3080 2696
rect 2935 2692 2965 2694
rect 2935 2691 2936 2692
rect 2930 2690 2936 2691
rect 3074 2691 3075 2695
rect 3079 2694 3080 2695
rect 3218 2695 3224 2696
rect 3079 2692 3109 2694
rect 3079 2691 3080 2692
rect 3074 2690 3080 2691
rect 3218 2691 3219 2695
rect 3223 2694 3224 2695
rect 3223 2692 3253 2694
rect 3223 2691 3224 2692
rect 3218 2690 3224 2691
rect 2746 2686 2752 2687
rect 2502 2659 2509 2660
rect 2502 2655 2503 2659
rect 2508 2655 2509 2659
rect 2502 2654 2509 2655
rect 2511 2659 2517 2660
rect 2511 2655 2512 2659
rect 2516 2658 2517 2659
rect 2639 2659 2645 2660
rect 2639 2658 2640 2659
rect 2516 2656 2640 2658
rect 2516 2655 2517 2656
rect 2511 2654 2517 2655
rect 2639 2655 2640 2656
rect 2644 2655 2645 2659
rect 2639 2654 2645 2655
rect 2783 2659 2792 2660
rect 2783 2655 2784 2659
rect 2791 2655 2792 2659
rect 2783 2654 2792 2655
rect 2927 2659 2936 2660
rect 2927 2655 2928 2659
rect 2935 2655 2936 2659
rect 2927 2654 2936 2655
rect 3071 2659 3080 2660
rect 3071 2655 3072 2659
rect 3079 2655 3080 2659
rect 3071 2654 3080 2655
rect 3215 2659 3224 2660
rect 3215 2655 3216 2659
rect 3223 2655 3224 2659
rect 3215 2654 3224 2655
rect 3270 2659 3276 2660
rect 3270 2655 3271 2659
rect 3275 2658 3276 2659
rect 3359 2659 3365 2660
rect 3359 2658 3360 2659
rect 3275 2656 3360 2658
rect 3275 2655 3276 2656
rect 3270 2654 3276 2655
rect 3359 2655 3360 2656
rect 3364 2655 3365 2659
rect 4218 2659 4224 2660
rect 4218 2658 4219 2659
rect 4189 2656 4219 2658
rect 3359 2654 3365 2655
rect 4218 2655 4219 2656
rect 4223 2655 4224 2659
rect 4218 2654 4224 2655
rect 4226 2659 4232 2660
rect 4226 2655 4227 2659
rect 4231 2658 4232 2659
rect 4426 2659 4432 2660
rect 4231 2656 4317 2658
rect 4231 2655 4232 2656
rect 4226 2654 4232 2655
rect 4426 2655 4427 2659
rect 4431 2658 4432 2659
rect 4642 2659 4648 2660
rect 4431 2656 4533 2658
rect 4431 2655 4432 2656
rect 4426 2654 4432 2655
rect 4642 2655 4643 2659
rect 4647 2658 4648 2659
rect 4882 2659 4888 2660
rect 4647 2656 4773 2658
rect 4647 2655 4648 2656
rect 4642 2654 4648 2655
rect 4882 2655 4883 2659
rect 4887 2658 4888 2659
rect 5398 2659 5404 2660
rect 5398 2658 5399 2659
rect 4887 2656 5029 2658
rect 5365 2656 5399 2658
rect 4887 2655 4888 2656
rect 4882 2654 4888 2655
rect 5398 2655 5399 2656
rect 5403 2655 5404 2659
rect 5618 2659 5624 2660
rect 5618 2658 5619 2659
rect 5605 2656 5619 2658
rect 5398 2654 5404 2655
rect 5618 2655 5619 2656
rect 5623 2655 5624 2659
rect 5618 2654 5624 2655
rect 1974 2652 1980 2653
rect 3798 2652 3804 2653
rect 903 2651 909 2652
rect 858 2647 864 2648
rect 858 2643 859 2647
rect 863 2643 864 2647
rect 903 2647 904 2651
rect 908 2650 909 2651
rect 1175 2651 1181 2652
rect 1175 2650 1176 2651
rect 908 2648 925 2650
rect 1133 2648 1176 2650
rect 908 2647 909 2648
rect 903 2646 909 2647
rect 1175 2647 1176 2648
rect 1180 2647 1181 2651
rect 1311 2651 1317 2652
rect 1311 2650 1312 2651
rect 1269 2648 1312 2650
rect 1175 2646 1181 2647
rect 1311 2647 1312 2648
rect 1316 2647 1317 2651
rect 1554 2651 1560 2652
rect 1554 2650 1555 2651
rect 1541 2648 1555 2650
rect 1311 2646 1317 2647
rect 1402 2647 1408 2648
rect 858 2642 864 2643
rect 1402 2643 1403 2647
rect 1407 2643 1408 2647
rect 1554 2647 1555 2648
rect 1559 2647 1560 2651
rect 1554 2646 1560 2647
rect 1583 2651 1589 2652
rect 1583 2647 1584 2651
rect 1588 2650 1589 2651
rect 1719 2651 1725 2652
rect 1588 2648 1605 2650
rect 1588 2647 1589 2648
rect 1583 2646 1589 2647
rect 1719 2647 1720 2651
rect 1724 2650 1725 2651
rect 1724 2648 1741 2650
rect 1974 2648 1975 2652
rect 1979 2648 1980 2652
rect 1724 2647 1725 2648
rect 1974 2647 1980 2648
rect 2378 2651 2384 2652
rect 2378 2647 2379 2651
rect 2383 2647 2384 2651
rect 1719 2646 1725 2647
rect 2378 2646 2384 2647
rect 2514 2651 2520 2652
rect 2514 2647 2515 2651
rect 2519 2647 2520 2651
rect 2514 2646 2520 2647
rect 2658 2651 2664 2652
rect 2658 2647 2659 2651
rect 2663 2647 2664 2651
rect 2658 2646 2664 2647
rect 2802 2651 2808 2652
rect 2802 2647 2803 2651
rect 2807 2647 2808 2651
rect 2802 2646 2808 2647
rect 2946 2651 2952 2652
rect 2946 2647 2947 2651
rect 2951 2647 2952 2651
rect 2946 2646 2952 2647
rect 3090 2651 3096 2652
rect 3090 2647 3091 2651
rect 3095 2647 3096 2651
rect 3090 2646 3096 2647
rect 3234 2651 3240 2652
rect 3234 2647 3235 2651
rect 3239 2647 3240 2651
rect 3798 2648 3799 2652
rect 3803 2648 3804 2652
rect 3798 2647 3804 2648
rect 3234 2646 3240 2647
rect 1402 2642 1408 2643
rect 2406 2636 2412 2637
rect 1974 2635 1980 2636
rect 1974 2631 1975 2635
rect 1979 2631 1980 2635
rect 2406 2632 2407 2636
rect 2411 2632 2412 2636
rect 2406 2631 2412 2632
rect 2542 2636 2548 2637
rect 2542 2632 2543 2636
rect 2547 2632 2548 2636
rect 2542 2631 2548 2632
rect 2686 2636 2692 2637
rect 2686 2632 2687 2636
rect 2691 2632 2692 2636
rect 2686 2631 2692 2632
rect 2830 2636 2836 2637
rect 2830 2632 2831 2636
rect 2835 2632 2836 2636
rect 2830 2631 2836 2632
rect 2974 2636 2980 2637
rect 2974 2632 2975 2636
rect 2979 2632 2980 2636
rect 2974 2631 2980 2632
rect 3118 2636 3124 2637
rect 3118 2632 3119 2636
rect 3123 2632 3124 2636
rect 3118 2631 3124 2632
rect 3262 2636 3268 2637
rect 3262 2632 3263 2636
rect 3267 2632 3268 2636
rect 3262 2631 3268 2632
rect 3798 2635 3804 2636
rect 3798 2631 3799 2635
rect 3803 2631 3804 2635
rect 1974 2630 1980 2631
rect 3798 2630 3804 2631
rect 858 2623 864 2624
rect 858 2619 859 2623
rect 863 2622 864 2623
rect 4223 2623 4232 2624
rect 863 2620 1042 2622
rect 863 2619 864 2620
rect 858 2618 864 2619
rect 895 2615 901 2616
rect 895 2611 896 2615
rect 900 2614 901 2615
rect 903 2615 909 2616
rect 903 2614 904 2615
rect 900 2612 904 2614
rect 900 2611 901 2612
rect 895 2610 901 2611
rect 903 2611 904 2612
rect 908 2611 909 2615
rect 903 2610 909 2611
rect 1030 2615 1037 2616
rect 1030 2611 1031 2615
rect 1036 2611 1037 2615
rect 1040 2614 1042 2620
rect 4223 2619 4224 2623
rect 4231 2619 4232 2623
rect 4223 2618 4232 2619
rect 4423 2623 4432 2624
rect 4423 2619 4424 2623
rect 4431 2619 4432 2623
rect 4423 2618 4432 2619
rect 4639 2623 4648 2624
rect 4639 2619 4640 2623
rect 4647 2619 4648 2623
rect 4639 2618 4648 2619
rect 4879 2623 4888 2624
rect 4879 2619 4880 2623
rect 4887 2619 4888 2623
rect 4879 2618 4888 2619
rect 4998 2623 5004 2624
rect 4998 2619 4999 2623
rect 5003 2622 5004 2623
rect 5135 2623 5141 2624
rect 5135 2622 5136 2623
rect 5003 2620 5136 2622
rect 5003 2619 5004 2620
rect 4998 2618 5004 2619
rect 5135 2619 5136 2620
rect 5140 2619 5141 2623
rect 5135 2618 5141 2619
rect 5338 2623 5344 2624
rect 5338 2619 5339 2623
rect 5343 2622 5344 2623
rect 5399 2623 5405 2624
rect 5399 2622 5400 2623
rect 5343 2620 5400 2622
rect 5343 2619 5344 2620
rect 5338 2618 5344 2619
rect 5399 2619 5400 2620
rect 5404 2619 5405 2623
rect 5399 2618 5405 2619
rect 5618 2623 5624 2624
rect 5618 2619 5619 2623
rect 5623 2622 5624 2623
rect 5639 2623 5645 2624
rect 5639 2622 5640 2623
rect 5623 2620 5640 2622
rect 5623 2619 5624 2620
rect 5618 2618 5624 2619
rect 5639 2619 5640 2620
rect 5644 2619 5645 2623
rect 5639 2618 5645 2619
rect 3838 2616 3844 2617
rect 5662 2616 5668 2617
rect 1167 2615 1173 2616
rect 1167 2614 1168 2615
rect 1040 2612 1168 2614
rect 1030 2610 1037 2611
rect 1167 2611 1168 2612
rect 1172 2611 1173 2615
rect 1167 2610 1173 2611
rect 1175 2615 1181 2616
rect 1175 2611 1176 2615
rect 1180 2614 1181 2615
rect 1303 2615 1309 2616
rect 1303 2614 1304 2615
rect 1180 2612 1304 2614
rect 1180 2611 1181 2612
rect 1175 2610 1181 2611
rect 1303 2611 1304 2612
rect 1308 2611 1309 2615
rect 1303 2610 1309 2611
rect 1311 2615 1317 2616
rect 1311 2611 1312 2615
rect 1316 2614 1317 2615
rect 1439 2615 1445 2616
rect 1439 2614 1440 2615
rect 1316 2612 1440 2614
rect 1316 2611 1317 2612
rect 1311 2610 1317 2611
rect 1439 2611 1440 2612
rect 1444 2611 1445 2615
rect 1439 2610 1445 2611
rect 1575 2615 1581 2616
rect 1575 2611 1576 2615
rect 1580 2614 1581 2615
rect 1583 2615 1589 2616
rect 1583 2614 1584 2615
rect 1580 2612 1584 2614
rect 1580 2611 1581 2612
rect 1575 2610 1581 2611
rect 1583 2611 1584 2612
rect 1588 2611 1589 2615
rect 1583 2610 1589 2611
rect 1711 2615 1717 2616
rect 1711 2611 1712 2615
rect 1716 2614 1717 2615
rect 1719 2615 1725 2616
rect 1719 2614 1720 2615
rect 1716 2612 1720 2614
rect 1716 2611 1717 2612
rect 1711 2610 1717 2611
rect 1719 2611 1720 2612
rect 1724 2611 1725 2615
rect 1719 2610 1725 2611
rect 1842 2615 1853 2616
rect 1842 2611 1843 2615
rect 1847 2611 1848 2615
rect 1852 2611 1853 2615
rect 3838 2612 3839 2616
rect 3843 2612 3844 2616
rect 3838 2611 3844 2612
rect 4098 2615 4104 2616
rect 4098 2611 4099 2615
rect 4103 2611 4104 2615
rect 1842 2610 1853 2611
rect 4098 2610 4104 2611
rect 4298 2615 4304 2616
rect 4298 2611 4299 2615
rect 4303 2611 4304 2615
rect 4298 2610 4304 2611
rect 4514 2615 4520 2616
rect 4514 2611 4515 2615
rect 4519 2611 4520 2615
rect 4514 2610 4520 2611
rect 4754 2615 4760 2616
rect 4754 2611 4755 2615
rect 4759 2611 4760 2615
rect 4754 2610 4760 2611
rect 5010 2615 5016 2616
rect 5010 2611 5011 2615
rect 5015 2611 5016 2615
rect 5010 2610 5016 2611
rect 5274 2615 5280 2616
rect 5274 2611 5275 2615
rect 5279 2611 5280 2615
rect 5274 2610 5280 2611
rect 5514 2615 5520 2616
rect 5514 2611 5515 2615
rect 5519 2611 5520 2615
rect 5662 2612 5663 2616
rect 5667 2612 5668 2616
rect 5662 2611 5668 2612
rect 5514 2610 5520 2611
rect 110 2608 116 2609
rect 1934 2608 1940 2609
rect 110 2604 111 2608
rect 115 2604 116 2608
rect 110 2603 116 2604
rect 770 2607 776 2608
rect 770 2603 771 2607
rect 775 2603 776 2607
rect 770 2602 776 2603
rect 906 2607 912 2608
rect 906 2603 907 2607
rect 911 2603 912 2607
rect 906 2602 912 2603
rect 1042 2607 1048 2608
rect 1042 2603 1043 2607
rect 1047 2603 1048 2607
rect 1042 2602 1048 2603
rect 1178 2607 1184 2608
rect 1178 2603 1179 2607
rect 1183 2603 1184 2607
rect 1178 2602 1184 2603
rect 1314 2607 1320 2608
rect 1314 2603 1315 2607
rect 1319 2603 1320 2607
rect 1314 2602 1320 2603
rect 1450 2607 1456 2608
rect 1450 2603 1451 2607
rect 1455 2603 1456 2607
rect 1450 2602 1456 2603
rect 1586 2607 1592 2608
rect 1586 2603 1587 2607
rect 1591 2603 1592 2607
rect 1586 2602 1592 2603
rect 1722 2607 1728 2608
rect 1722 2603 1723 2607
rect 1727 2603 1728 2607
rect 1934 2604 1935 2608
rect 1939 2604 1940 2608
rect 1934 2603 1940 2604
rect 1722 2602 1728 2603
rect 4126 2600 4132 2601
rect 3838 2599 3844 2600
rect 3838 2595 3839 2599
rect 3843 2595 3844 2599
rect 4126 2596 4127 2600
rect 4131 2596 4132 2600
rect 4126 2595 4132 2596
rect 4326 2600 4332 2601
rect 4326 2596 4327 2600
rect 4331 2596 4332 2600
rect 4326 2595 4332 2596
rect 4542 2600 4548 2601
rect 4542 2596 4543 2600
rect 4547 2596 4548 2600
rect 4542 2595 4548 2596
rect 4782 2600 4788 2601
rect 4782 2596 4783 2600
rect 4787 2596 4788 2600
rect 4782 2595 4788 2596
rect 5038 2600 5044 2601
rect 5038 2596 5039 2600
rect 5043 2596 5044 2600
rect 5038 2595 5044 2596
rect 5302 2600 5308 2601
rect 5302 2596 5303 2600
rect 5307 2596 5308 2600
rect 5302 2595 5308 2596
rect 5542 2600 5548 2601
rect 5542 2596 5543 2600
rect 5547 2596 5548 2600
rect 5542 2595 5548 2596
rect 5662 2599 5668 2600
rect 5662 2595 5663 2599
rect 5667 2595 5668 2599
rect 3838 2594 3844 2595
rect 5662 2594 5668 2595
rect 798 2592 804 2593
rect 110 2591 116 2592
rect 110 2587 111 2591
rect 115 2587 116 2591
rect 798 2588 799 2592
rect 803 2588 804 2592
rect 798 2587 804 2588
rect 934 2592 940 2593
rect 934 2588 935 2592
rect 939 2588 940 2592
rect 934 2587 940 2588
rect 1070 2592 1076 2593
rect 1070 2588 1071 2592
rect 1075 2588 1076 2592
rect 1070 2587 1076 2588
rect 1206 2592 1212 2593
rect 1206 2588 1207 2592
rect 1211 2588 1212 2592
rect 1206 2587 1212 2588
rect 1342 2592 1348 2593
rect 1342 2588 1343 2592
rect 1347 2588 1348 2592
rect 1342 2587 1348 2588
rect 1478 2592 1484 2593
rect 1478 2588 1479 2592
rect 1483 2588 1484 2592
rect 1478 2587 1484 2588
rect 1614 2592 1620 2593
rect 1614 2588 1615 2592
rect 1619 2588 1620 2592
rect 1614 2587 1620 2588
rect 1750 2592 1756 2593
rect 1750 2588 1751 2592
rect 1755 2588 1756 2592
rect 1750 2587 1756 2588
rect 1934 2591 1940 2592
rect 1934 2587 1935 2591
rect 1939 2587 1940 2591
rect 110 2586 116 2587
rect 1934 2586 1940 2587
rect 1974 2573 1980 2574
rect 3798 2573 3804 2574
rect 1974 2569 1975 2573
rect 1979 2569 1980 2573
rect 1974 2568 1980 2569
rect 2510 2572 2516 2573
rect 2510 2568 2511 2572
rect 2515 2568 2516 2572
rect 2510 2567 2516 2568
rect 2646 2572 2652 2573
rect 2646 2568 2647 2572
rect 2651 2568 2652 2572
rect 2646 2567 2652 2568
rect 2782 2572 2788 2573
rect 2782 2568 2783 2572
rect 2787 2568 2788 2572
rect 2782 2567 2788 2568
rect 2918 2572 2924 2573
rect 2918 2568 2919 2572
rect 2923 2568 2924 2572
rect 2918 2567 2924 2568
rect 3054 2572 3060 2573
rect 3054 2568 3055 2572
rect 3059 2568 3060 2572
rect 3054 2567 3060 2568
rect 3190 2572 3196 2573
rect 3190 2568 3191 2572
rect 3195 2568 3196 2572
rect 3190 2567 3196 2568
rect 3326 2572 3332 2573
rect 3326 2568 3327 2572
rect 3331 2568 3332 2572
rect 3326 2567 3332 2568
rect 3462 2572 3468 2573
rect 3462 2568 3463 2572
rect 3467 2568 3468 2572
rect 3798 2569 3799 2573
rect 3803 2569 3804 2573
rect 3798 2568 3804 2569
rect 3462 2567 3468 2568
rect 2482 2557 2488 2558
rect 1974 2556 1980 2557
rect 1974 2552 1975 2556
rect 1979 2552 1980 2556
rect 2482 2553 2483 2557
rect 2487 2553 2488 2557
rect 2482 2552 2488 2553
rect 2618 2557 2624 2558
rect 2618 2553 2619 2557
rect 2623 2553 2624 2557
rect 2618 2552 2624 2553
rect 2754 2557 2760 2558
rect 2754 2553 2755 2557
rect 2759 2553 2760 2557
rect 2754 2552 2760 2553
rect 2890 2557 2896 2558
rect 2890 2553 2891 2557
rect 2895 2553 2896 2557
rect 2890 2552 2896 2553
rect 3026 2557 3032 2558
rect 3026 2553 3027 2557
rect 3031 2553 3032 2557
rect 3026 2552 3032 2553
rect 3162 2557 3168 2558
rect 3162 2553 3163 2557
rect 3167 2553 3168 2557
rect 3162 2552 3168 2553
rect 3298 2557 3304 2558
rect 3298 2553 3299 2557
rect 3303 2553 3304 2557
rect 3298 2552 3304 2553
rect 3434 2557 3440 2558
rect 3434 2553 3435 2557
rect 3439 2553 3440 2557
rect 3434 2552 3440 2553
rect 3798 2556 3804 2557
rect 3798 2552 3799 2556
rect 3803 2552 3804 2556
rect 1974 2551 1980 2552
rect 3798 2551 3804 2552
rect 2602 2547 2613 2548
rect 2602 2543 2603 2547
rect 2607 2543 2608 2547
rect 2612 2543 2613 2547
rect 2602 2542 2613 2543
rect 2615 2547 2621 2548
rect 2615 2543 2616 2547
rect 2620 2546 2621 2547
rect 2743 2547 2749 2548
rect 2743 2546 2744 2547
rect 2620 2544 2744 2546
rect 2620 2543 2621 2544
rect 2615 2542 2621 2543
rect 2743 2543 2744 2544
rect 2748 2543 2749 2547
rect 2743 2542 2749 2543
rect 2751 2547 2757 2548
rect 2751 2543 2752 2547
rect 2756 2546 2757 2547
rect 2879 2547 2885 2548
rect 2879 2546 2880 2547
rect 2756 2544 2880 2546
rect 2756 2543 2757 2544
rect 2751 2542 2757 2543
rect 2879 2543 2880 2544
rect 2884 2543 2885 2547
rect 2879 2542 2885 2543
rect 3015 2547 3021 2548
rect 3015 2543 3016 2547
rect 3020 2546 3021 2547
rect 3042 2547 3048 2548
rect 3042 2546 3043 2547
rect 3020 2544 3043 2546
rect 3020 2543 3021 2544
rect 3015 2542 3021 2543
rect 3042 2543 3043 2544
rect 3047 2543 3048 2547
rect 3042 2542 3048 2543
rect 3151 2547 3157 2548
rect 3151 2543 3152 2547
rect 3156 2546 3157 2547
rect 3178 2547 3184 2548
rect 3178 2546 3179 2547
rect 3156 2544 3179 2546
rect 3156 2543 3157 2544
rect 3151 2542 3157 2543
rect 3178 2543 3179 2544
rect 3183 2543 3184 2547
rect 3178 2542 3184 2543
rect 3287 2547 3293 2548
rect 3287 2543 3288 2547
rect 3292 2546 3293 2547
rect 3314 2547 3320 2548
rect 3314 2546 3315 2547
rect 3292 2544 3315 2546
rect 3292 2543 3293 2544
rect 3287 2542 3293 2543
rect 3314 2543 3315 2544
rect 3319 2543 3320 2547
rect 3314 2542 3320 2543
rect 3423 2547 3429 2548
rect 3423 2543 3424 2547
rect 3428 2546 3429 2547
rect 3450 2547 3456 2548
rect 3450 2546 3451 2547
rect 3428 2544 3451 2546
rect 3428 2543 3429 2544
rect 3423 2542 3429 2543
rect 3450 2543 3451 2544
rect 3455 2543 3456 2547
rect 3559 2547 3565 2548
rect 3559 2546 3560 2547
rect 3450 2542 3456 2543
rect 3460 2544 3560 2546
rect 2978 2539 2984 2540
rect 2978 2535 2979 2539
rect 2983 2538 2984 2539
rect 3270 2539 3276 2540
rect 3270 2538 3271 2539
rect 2983 2536 3271 2538
rect 2983 2535 2984 2536
rect 2978 2534 2984 2535
rect 3270 2535 3271 2536
rect 3275 2535 3276 2539
rect 3270 2534 3276 2535
rect 3014 2531 3020 2532
rect 3014 2527 3015 2531
rect 3019 2530 3020 2531
rect 3460 2530 3462 2544
rect 3559 2543 3560 2544
rect 3564 2543 3565 2547
rect 3559 2542 3565 2543
rect 3838 2537 3844 2538
rect 5662 2537 5668 2538
rect 3838 2533 3839 2537
rect 3843 2533 3844 2537
rect 3838 2532 3844 2533
rect 4494 2536 4500 2537
rect 4494 2532 4495 2536
rect 4499 2532 4500 2536
rect 4494 2531 4500 2532
rect 4630 2536 4636 2537
rect 4630 2532 4631 2536
rect 4635 2532 4636 2536
rect 4630 2531 4636 2532
rect 4766 2536 4772 2537
rect 4766 2532 4767 2536
rect 4771 2532 4772 2536
rect 4766 2531 4772 2532
rect 4902 2536 4908 2537
rect 4902 2532 4903 2536
rect 4907 2532 4908 2536
rect 4902 2531 4908 2532
rect 5038 2536 5044 2537
rect 5038 2532 5039 2536
rect 5043 2532 5044 2536
rect 5662 2533 5663 2537
rect 5667 2533 5668 2537
rect 5662 2532 5668 2533
rect 5038 2531 5044 2532
rect 3019 2528 3462 2530
rect 3019 2527 3020 2528
rect 3014 2526 3020 2527
rect 4466 2521 4472 2522
rect 3838 2520 3844 2521
rect 110 2517 116 2518
rect 1934 2517 1940 2518
rect 110 2513 111 2517
rect 115 2513 116 2517
rect 110 2512 116 2513
rect 550 2516 556 2517
rect 550 2512 551 2516
rect 555 2512 556 2516
rect 550 2511 556 2512
rect 686 2516 692 2517
rect 686 2512 687 2516
rect 691 2512 692 2516
rect 686 2511 692 2512
rect 830 2516 836 2517
rect 830 2512 831 2516
rect 835 2512 836 2516
rect 830 2511 836 2512
rect 982 2516 988 2517
rect 982 2512 983 2516
rect 987 2512 988 2516
rect 982 2511 988 2512
rect 1134 2516 1140 2517
rect 1134 2512 1135 2516
rect 1139 2512 1140 2516
rect 1134 2511 1140 2512
rect 1294 2516 1300 2517
rect 1294 2512 1295 2516
rect 1299 2512 1300 2516
rect 1294 2511 1300 2512
rect 1454 2516 1460 2517
rect 1454 2512 1455 2516
rect 1459 2512 1460 2516
rect 1454 2511 1460 2512
rect 1614 2516 1620 2517
rect 1614 2512 1615 2516
rect 1619 2512 1620 2516
rect 1614 2511 1620 2512
rect 1782 2516 1788 2517
rect 1782 2512 1783 2516
rect 1787 2512 1788 2516
rect 1934 2513 1935 2517
rect 1939 2513 1940 2517
rect 3838 2516 3839 2520
rect 3843 2516 3844 2520
rect 4466 2517 4467 2521
rect 4471 2517 4472 2521
rect 4466 2516 4472 2517
rect 4602 2521 4608 2522
rect 4602 2517 4603 2521
rect 4607 2517 4608 2521
rect 4602 2516 4608 2517
rect 4738 2521 4744 2522
rect 4738 2517 4739 2521
rect 4743 2517 4744 2521
rect 4738 2516 4744 2517
rect 4874 2521 4880 2522
rect 4874 2517 4875 2521
rect 4879 2517 4880 2521
rect 4874 2516 4880 2517
rect 5010 2521 5016 2522
rect 5010 2517 5011 2521
rect 5015 2517 5016 2521
rect 5010 2516 5016 2517
rect 5662 2520 5668 2521
rect 5662 2516 5663 2520
rect 5667 2516 5668 2520
rect 2615 2515 2621 2516
rect 2615 2514 2616 2515
rect 1934 2512 1940 2513
rect 2573 2512 2616 2514
rect 1782 2511 1788 2512
rect 2615 2511 2616 2512
rect 2620 2511 2621 2515
rect 2751 2515 2757 2516
rect 2751 2514 2752 2515
rect 2709 2512 2752 2514
rect 2615 2510 2621 2511
rect 2751 2511 2752 2512
rect 2756 2511 2757 2515
rect 2751 2510 2757 2511
rect 2838 2515 2844 2516
rect 2838 2511 2839 2515
rect 2843 2511 2844 2515
rect 2838 2510 2844 2511
rect 2978 2515 2984 2516
rect 2978 2511 2979 2515
rect 2983 2511 2984 2515
rect 2978 2510 2984 2511
rect 3042 2515 3048 2516
rect 3042 2511 3043 2515
rect 3047 2511 3048 2515
rect 3042 2510 3048 2511
rect 3178 2515 3184 2516
rect 3178 2511 3179 2515
rect 3183 2511 3184 2515
rect 3178 2510 3184 2511
rect 3314 2515 3320 2516
rect 3314 2511 3315 2515
rect 3319 2511 3320 2515
rect 3314 2510 3320 2511
rect 3450 2515 3456 2516
rect 3838 2515 3844 2516
rect 5662 2515 5668 2516
rect 3450 2511 3451 2515
rect 3455 2511 3456 2515
rect 3450 2510 3456 2511
rect 4591 2511 4597 2512
rect 4591 2507 4592 2511
rect 4596 2510 4597 2511
rect 4618 2511 4624 2512
rect 4618 2510 4619 2511
rect 4596 2508 4619 2510
rect 4596 2507 4597 2508
rect 4591 2506 4597 2507
rect 4618 2507 4619 2508
rect 4623 2507 4624 2511
rect 4618 2506 4624 2507
rect 4727 2511 4733 2512
rect 4727 2507 4728 2511
rect 4732 2510 4733 2511
rect 4754 2511 4760 2512
rect 4754 2510 4755 2511
rect 4732 2508 4755 2510
rect 4732 2507 4733 2508
rect 4727 2506 4733 2507
rect 4754 2507 4755 2508
rect 4759 2507 4760 2511
rect 4754 2506 4760 2507
rect 4863 2511 4869 2512
rect 4863 2507 4864 2511
rect 4868 2510 4869 2511
rect 4890 2511 4896 2512
rect 4890 2510 4891 2511
rect 4868 2508 4891 2510
rect 4868 2507 4869 2508
rect 4863 2506 4869 2507
rect 4890 2507 4891 2508
rect 4895 2507 4896 2511
rect 4890 2506 4896 2507
rect 4999 2511 5005 2512
rect 4999 2507 5000 2511
rect 5004 2510 5005 2511
rect 5026 2511 5032 2512
rect 5026 2510 5027 2511
rect 5004 2508 5027 2510
rect 5004 2507 5005 2508
rect 4999 2506 5005 2507
rect 5026 2507 5027 2508
rect 5031 2507 5032 2511
rect 5135 2511 5141 2512
rect 5135 2510 5136 2511
rect 5026 2506 5032 2507
rect 5036 2508 5136 2510
rect 4818 2503 4824 2504
rect 522 2501 528 2502
rect 110 2500 116 2501
rect 110 2496 111 2500
rect 115 2496 116 2500
rect 522 2497 523 2501
rect 527 2497 528 2501
rect 522 2496 528 2497
rect 658 2501 664 2502
rect 658 2497 659 2501
rect 663 2497 664 2501
rect 658 2496 664 2497
rect 802 2501 808 2502
rect 802 2497 803 2501
rect 807 2497 808 2501
rect 802 2496 808 2497
rect 954 2501 960 2502
rect 954 2497 955 2501
rect 959 2497 960 2501
rect 954 2496 960 2497
rect 1106 2501 1112 2502
rect 1106 2497 1107 2501
rect 1111 2497 1112 2501
rect 1106 2496 1112 2497
rect 1266 2501 1272 2502
rect 1266 2497 1267 2501
rect 1271 2497 1272 2501
rect 1266 2496 1272 2497
rect 1426 2501 1432 2502
rect 1426 2497 1427 2501
rect 1431 2497 1432 2501
rect 1426 2496 1432 2497
rect 1586 2501 1592 2502
rect 1586 2497 1587 2501
rect 1591 2497 1592 2501
rect 1586 2496 1592 2497
rect 1754 2501 1760 2502
rect 1754 2497 1755 2501
rect 1759 2497 1760 2501
rect 1754 2496 1760 2497
rect 1934 2500 1940 2501
rect 1934 2496 1935 2500
rect 1939 2496 1940 2500
rect 4818 2499 4819 2503
rect 4823 2502 4824 2503
rect 5036 2502 5038 2508
rect 5135 2507 5136 2508
rect 5140 2507 5141 2511
rect 5135 2506 5141 2507
rect 4823 2500 5038 2502
rect 4823 2499 4824 2500
rect 4818 2498 4824 2499
rect 110 2495 116 2496
rect 1934 2495 1940 2496
rect 4998 2495 5004 2496
rect 4998 2494 4999 2495
rect 4608 2492 4999 2494
rect 647 2491 653 2492
rect 647 2487 648 2491
rect 652 2490 653 2491
rect 674 2491 680 2492
rect 674 2490 675 2491
rect 652 2488 675 2490
rect 652 2487 653 2488
rect 647 2486 653 2487
rect 674 2487 675 2488
rect 679 2487 680 2491
rect 674 2486 680 2487
rect 783 2491 789 2492
rect 783 2487 784 2491
rect 788 2490 789 2491
rect 818 2491 824 2492
rect 818 2490 819 2491
rect 788 2488 819 2490
rect 788 2487 789 2488
rect 783 2486 789 2487
rect 818 2487 819 2488
rect 823 2487 824 2491
rect 818 2486 824 2487
rect 927 2491 933 2492
rect 927 2487 928 2491
rect 932 2490 933 2491
rect 970 2491 976 2492
rect 970 2490 971 2491
rect 932 2488 971 2490
rect 932 2487 933 2488
rect 927 2486 933 2487
rect 970 2487 971 2488
rect 975 2487 976 2491
rect 970 2486 976 2487
rect 1079 2491 1085 2492
rect 1079 2487 1080 2491
rect 1084 2490 1085 2491
rect 1122 2491 1128 2492
rect 1122 2490 1123 2491
rect 1084 2488 1123 2490
rect 1084 2487 1085 2488
rect 1079 2486 1085 2487
rect 1122 2487 1123 2488
rect 1127 2487 1128 2491
rect 1122 2486 1128 2487
rect 1231 2491 1237 2492
rect 1231 2487 1232 2491
rect 1236 2490 1237 2491
rect 1282 2491 1288 2492
rect 1282 2490 1283 2491
rect 1236 2488 1283 2490
rect 1236 2487 1237 2488
rect 1231 2486 1237 2487
rect 1282 2487 1283 2488
rect 1287 2487 1288 2491
rect 1282 2486 1288 2487
rect 1391 2491 1397 2492
rect 1391 2487 1392 2491
rect 1396 2490 1397 2491
rect 1402 2491 1408 2492
rect 1402 2490 1403 2491
rect 1396 2488 1403 2490
rect 1396 2487 1397 2488
rect 1391 2486 1397 2487
rect 1402 2487 1403 2488
rect 1407 2487 1408 2491
rect 1402 2486 1408 2487
rect 1410 2491 1416 2492
rect 1410 2487 1411 2491
rect 1415 2490 1416 2491
rect 1551 2491 1557 2492
rect 1551 2490 1552 2491
rect 1415 2488 1552 2490
rect 1415 2487 1416 2488
rect 1410 2486 1416 2487
rect 1551 2487 1552 2488
rect 1556 2487 1557 2491
rect 1551 2486 1557 2487
rect 1583 2491 1589 2492
rect 1583 2487 1584 2491
rect 1588 2490 1589 2491
rect 1711 2491 1717 2492
rect 1711 2490 1712 2491
rect 1588 2488 1712 2490
rect 1588 2487 1589 2488
rect 1583 2486 1589 2487
rect 1711 2487 1712 2488
rect 1716 2487 1717 2491
rect 1711 2486 1717 2487
rect 1742 2491 1748 2492
rect 1742 2487 1743 2491
rect 1747 2490 1748 2491
rect 1879 2491 1885 2492
rect 1879 2490 1880 2491
rect 1747 2488 1880 2490
rect 1747 2487 1748 2488
rect 1742 2486 1748 2487
rect 1879 2487 1880 2488
rect 1884 2487 1885 2491
rect 1879 2486 1885 2487
rect 4608 2478 4610 2492
rect 4998 2491 4999 2492
rect 5003 2491 5004 2495
rect 4998 2490 5004 2491
rect 4557 2476 4610 2478
rect 4618 2479 4624 2480
rect 4618 2475 4619 2479
rect 4623 2475 4624 2479
rect 4618 2474 4624 2475
rect 4754 2479 4760 2480
rect 4754 2475 4755 2479
rect 4759 2475 4760 2479
rect 4754 2474 4760 2475
rect 4890 2479 4896 2480
rect 4890 2475 4891 2479
rect 4895 2475 4896 2479
rect 4890 2474 4896 2475
rect 5026 2479 5032 2480
rect 5026 2475 5027 2479
rect 5031 2475 5032 2479
rect 5026 2474 5032 2475
rect 666 2459 672 2460
rect 666 2458 667 2459
rect 613 2456 667 2458
rect 666 2455 667 2456
rect 671 2455 672 2459
rect 666 2454 672 2455
rect 674 2459 680 2460
rect 674 2455 675 2459
rect 679 2455 680 2459
rect 674 2454 680 2455
rect 818 2459 824 2460
rect 818 2455 819 2459
rect 823 2455 824 2459
rect 818 2454 824 2455
rect 970 2459 976 2460
rect 970 2455 971 2459
rect 975 2455 976 2459
rect 970 2454 976 2455
rect 1122 2459 1128 2460
rect 1122 2455 1123 2459
rect 1127 2455 1128 2459
rect 1122 2454 1128 2455
rect 1282 2459 1288 2460
rect 1282 2455 1283 2459
rect 1287 2455 1288 2459
rect 1583 2459 1589 2460
rect 1583 2458 1584 2459
rect 1517 2456 1584 2458
rect 1282 2454 1288 2455
rect 1583 2455 1584 2456
rect 1588 2455 1589 2459
rect 1742 2459 1748 2460
rect 1742 2458 1743 2459
rect 1677 2456 1743 2458
rect 1583 2454 1589 2455
rect 1742 2455 1743 2456
rect 1747 2455 1748 2459
rect 1742 2454 1748 2455
rect 1842 2459 1848 2460
rect 1842 2455 1843 2459
rect 1847 2455 1848 2459
rect 1842 2454 1848 2455
rect 2298 2451 2304 2452
rect 2298 2447 2299 2451
rect 2303 2450 2304 2451
rect 2434 2451 2440 2452
rect 2303 2448 2325 2450
rect 2303 2447 2304 2448
rect 2298 2446 2304 2447
rect 2434 2447 2435 2451
rect 2439 2450 2440 2451
rect 2642 2451 2648 2452
rect 2439 2448 2533 2450
rect 2439 2447 2440 2448
rect 2434 2446 2440 2447
rect 2642 2447 2643 2451
rect 2647 2450 2648 2451
rect 3014 2451 3020 2452
rect 3014 2450 3015 2451
rect 2647 2448 2733 2450
rect 2997 2448 3015 2450
rect 2647 2447 2648 2448
rect 2642 2446 2648 2447
rect 3014 2447 3015 2448
rect 3019 2447 3020 2451
rect 3014 2446 3020 2447
rect 3034 2451 3040 2452
rect 3034 2447 3035 2451
rect 3039 2450 3040 2451
rect 3226 2451 3232 2452
rect 3039 2448 3117 2450
rect 3039 2447 3040 2448
rect 3034 2446 3040 2447
rect 3226 2447 3227 2451
rect 3231 2450 3232 2451
rect 3410 2451 3416 2452
rect 3231 2448 3301 2450
rect 3231 2447 3232 2448
rect 3226 2446 3232 2447
rect 3410 2447 3411 2451
rect 3415 2450 3416 2451
rect 3594 2451 3600 2452
rect 3415 2448 3485 2450
rect 3415 2447 3416 2448
rect 3410 2446 3416 2447
rect 3594 2447 3595 2451
rect 3599 2450 3600 2451
rect 3599 2448 3669 2450
rect 3599 2447 3600 2448
rect 3594 2446 3600 2447
rect 2431 2415 2440 2416
rect 2431 2411 2432 2415
rect 2439 2411 2440 2415
rect 2431 2410 2440 2411
rect 2639 2415 2648 2416
rect 2639 2411 2640 2415
rect 2647 2411 2648 2415
rect 2639 2410 2648 2411
rect 2838 2415 2845 2416
rect 2838 2411 2839 2415
rect 2844 2411 2845 2415
rect 2838 2410 2845 2411
rect 3031 2415 3040 2416
rect 3031 2411 3032 2415
rect 3039 2411 3040 2415
rect 3031 2410 3040 2411
rect 3223 2415 3232 2416
rect 3223 2411 3224 2415
rect 3231 2411 3232 2415
rect 3223 2410 3232 2411
rect 3407 2415 3416 2416
rect 3407 2411 3408 2415
rect 3415 2411 3416 2415
rect 3407 2410 3416 2411
rect 3591 2415 3600 2416
rect 3591 2411 3592 2415
rect 3599 2411 3600 2415
rect 3591 2410 3600 2411
rect 3738 2415 3744 2416
rect 3738 2411 3739 2415
rect 3743 2414 3744 2415
rect 3775 2415 3781 2416
rect 3775 2414 3776 2415
rect 3743 2412 3776 2414
rect 3743 2411 3744 2412
rect 3738 2410 3744 2411
rect 3775 2411 3776 2412
rect 3780 2411 3781 2415
rect 4818 2415 4824 2416
rect 4818 2414 4819 2415
rect 4789 2412 4819 2414
rect 3775 2410 3781 2411
rect 4818 2411 4819 2412
rect 4823 2411 4824 2415
rect 4818 2410 4824 2411
rect 4826 2415 4832 2416
rect 4826 2411 4827 2415
rect 4831 2414 4832 2415
rect 4967 2415 4973 2416
rect 4831 2412 4853 2414
rect 4831 2411 4832 2412
rect 4826 2410 4832 2411
rect 4967 2411 4968 2415
rect 4972 2414 4973 2415
rect 5103 2415 5109 2416
rect 4972 2412 4989 2414
rect 4972 2411 4973 2412
rect 4967 2410 4973 2411
rect 5103 2411 5104 2415
rect 5108 2414 5109 2415
rect 5239 2415 5245 2416
rect 5108 2412 5125 2414
rect 5108 2411 5109 2412
rect 5103 2410 5109 2411
rect 5239 2411 5240 2415
rect 5244 2414 5245 2415
rect 5618 2415 5624 2416
rect 5618 2414 5619 2415
rect 5244 2412 5261 2414
rect 5605 2412 5619 2414
rect 5244 2411 5245 2412
rect 5239 2410 5245 2411
rect 5466 2411 5472 2412
rect 1974 2408 1980 2409
rect 3798 2408 3804 2409
rect 1974 2404 1975 2408
rect 1979 2404 1980 2408
rect 1974 2403 1980 2404
rect 2306 2407 2312 2408
rect 2306 2403 2307 2407
rect 2311 2403 2312 2407
rect 2306 2402 2312 2403
rect 2514 2407 2520 2408
rect 2514 2403 2515 2407
rect 2519 2403 2520 2407
rect 2514 2402 2520 2403
rect 2714 2407 2720 2408
rect 2714 2403 2715 2407
rect 2719 2403 2720 2407
rect 2714 2402 2720 2403
rect 2906 2407 2912 2408
rect 2906 2403 2907 2407
rect 2911 2403 2912 2407
rect 2906 2402 2912 2403
rect 3098 2407 3104 2408
rect 3098 2403 3099 2407
rect 3103 2403 3104 2407
rect 3098 2402 3104 2403
rect 3282 2407 3288 2408
rect 3282 2403 3283 2407
rect 3287 2403 3288 2407
rect 3282 2402 3288 2403
rect 3466 2407 3472 2408
rect 3466 2403 3467 2407
rect 3471 2403 3472 2407
rect 3466 2402 3472 2403
rect 3650 2407 3656 2408
rect 3650 2403 3651 2407
rect 3655 2403 3656 2407
rect 3798 2404 3799 2408
rect 3803 2404 3804 2408
rect 5466 2407 5467 2411
rect 5471 2407 5472 2411
rect 5618 2411 5619 2412
rect 5623 2411 5624 2415
rect 5618 2410 5624 2411
rect 5466 2406 5472 2407
rect 3798 2403 3804 2404
rect 3650 2402 3656 2403
rect 306 2399 312 2400
rect 218 2395 224 2396
rect 218 2391 219 2395
rect 223 2391 224 2395
rect 306 2395 307 2399
rect 311 2398 312 2399
rect 466 2399 472 2400
rect 311 2396 357 2398
rect 311 2395 312 2396
rect 306 2394 312 2395
rect 466 2395 467 2399
rect 471 2398 472 2399
rect 690 2399 696 2400
rect 471 2396 581 2398
rect 471 2395 472 2396
rect 466 2394 472 2395
rect 690 2395 691 2399
rect 695 2398 696 2399
rect 930 2399 936 2400
rect 695 2396 821 2398
rect 695 2395 696 2396
rect 690 2394 696 2395
rect 930 2395 931 2399
rect 935 2398 936 2399
rect 1410 2399 1416 2400
rect 1410 2398 1411 2399
rect 935 2396 1061 2398
rect 1381 2396 1411 2398
rect 935 2395 936 2396
rect 930 2394 936 2395
rect 1410 2395 1411 2396
rect 1415 2395 1416 2399
rect 1410 2394 1416 2395
rect 1438 2399 1444 2400
rect 1438 2395 1439 2399
rect 1443 2398 1444 2399
rect 1674 2399 1680 2400
rect 1443 2396 1565 2398
rect 1443 2395 1444 2396
rect 1438 2394 1444 2395
rect 1674 2395 1675 2399
rect 1679 2398 1680 2399
rect 1679 2396 1805 2398
rect 1679 2395 1680 2396
rect 1674 2394 1680 2395
rect 2334 2392 2340 2393
rect 218 2390 224 2391
rect 1974 2391 1980 2392
rect 1974 2387 1975 2391
rect 1979 2387 1980 2391
rect 2334 2388 2335 2392
rect 2339 2388 2340 2392
rect 2334 2387 2340 2388
rect 2542 2392 2548 2393
rect 2542 2388 2543 2392
rect 2547 2388 2548 2392
rect 2542 2387 2548 2388
rect 2742 2392 2748 2393
rect 2742 2388 2743 2392
rect 2747 2388 2748 2392
rect 2742 2387 2748 2388
rect 2934 2392 2940 2393
rect 2934 2388 2935 2392
rect 2939 2388 2940 2392
rect 2934 2387 2940 2388
rect 3126 2392 3132 2393
rect 3126 2388 3127 2392
rect 3131 2388 3132 2392
rect 3126 2387 3132 2388
rect 3310 2392 3316 2393
rect 3310 2388 3311 2392
rect 3315 2388 3316 2392
rect 3310 2387 3316 2388
rect 3494 2392 3500 2393
rect 3494 2388 3495 2392
rect 3499 2388 3500 2392
rect 3494 2387 3500 2388
rect 3678 2392 3684 2393
rect 3678 2388 3679 2392
rect 3683 2388 3684 2392
rect 3678 2387 3684 2388
rect 3798 2391 3804 2392
rect 3798 2387 3799 2391
rect 3803 2387 3804 2391
rect 1974 2386 1980 2387
rect 3798 2386 3804 2387
rect 5466 2387 5472 2388
rect 5466 2383 5467 2387
rect 5471 2386 5472 2387
rect 5550 2387 5556 2388
rect 5550 2386 5551 2387
rect 5471 2384 5551 2386
rect 5471 2383 5472 2384
rect 5466 2382 5472 2383
rect 5550 2383 5551 2384
rect 5555 2383 5556 2387
rect 5550 2382 5556 2383
rect 4823 2379 4832 2380
rect 4823 2375 4824 2379
rect 4831 2375 4832 2379
rect 4823 2374 4832 2375
rect 4959 2379 4965 2380
rect 4959 2375 4960 2379
rect 4964 2378 4965 2379
rect 4967 2379 4973 2380
rect 4967 2378 4968 2379
rect 4964 2376 4968 2378
rect 4964 2375 4965 2376
rect 4959 2374 4965 2375
rect 4967 2375 4968 2376
rect 4972 2375 4973 2379
rect 4967 2374 4973 2375
rect 5095 2379 5101 2380
rect 5095 2375 5096 2379
rect 5100 2378 5101 2379
rect 5103 2379 5109 2380
rect 5103 2378 5104 2379
rect 5100 2376 5104 2378
rect 5100 2375 5101 2376
rect 5095 2374 5101 2375
rect 5103 2375 5104 2376
rect 5108 2375 5109 2379
rect 5103 2374 5109 2375
rect 5231 2379 5237 2380
rect 5231 2375 5232 2379
rect 5236 2378 5237 2379
rect 5239 2379 5245 2380
rect 5239 2378 5240 2379
rect 5236 2376 5240 2378
rect 5236 2375 5237 2376
rect 5231 2374 5237 2375
rect 5239 2375 5240 2376
rect 5244 2375 5245 2379
rect 5239 2374 5245 2375
rect 5367 2379 5376 2380
rect 5367 2375 5368 2379
rect 5375 2375 5376 2379
rect 5367 2374 5376 2375
rect 5398 2379 5404 2380
rect 5398 2375 5399 2379
rect 5403 2378 5404 2379
rect 5503 2379 5509 2380
rect 5503 2378 5504 2379
rect 5403 2376 5504 2378
rect 5403 2375 5404 2376
rect 5398 2374 5404 2375
rect 5503 2375 5504 2376
rect 5508 2375 5509 2379
rect 5503 2374 5509 2375
rect 5618 2379 5624 2380
rect 5618 2375 5619 2379
rect 5623 2378 5624 2379
rect 5639 2379 5645 2380
rect 5639 2378 5640 2379
rect 5623 2376 5640 2378
rect 5623 2375 5624 2376
rect 5618 2374 5624 2375
rect 5639 2375 5640 2376
rect 5644 2375 5645 2379
rect 5639 2374 5645 2375
rect 3838 2372 3844 2373
rect 5662 2372 5668 2373
rect 666 2371 672 2372
rect 666 2367 667 2371
rect 671 2370 672 2371
rect 671 2368 942 2370
rect 671 2367 672 2368
rect 666 2366 672 2367
rect 255 2363 261 2364
rect 255 2359 256 2363
rect 260 2362 261 2363
rect 306 2363 312 2364
rect 306 2362 307 2363
rect 260 2360 307 2362
rect 260 2359 261 2360
rect 255 2358 261 2359
rect 306 2359 307 2360
rect 311 2359 312 2363
rect 306 2358 312 2359
rect 463 2363 472 2364
rect 463 2359 464 2363
rect 471 2359 472 2363
rect 463 2358 472 2359
rect 687 2363 696 2364
rect 687 2359 688 2363
rect 695 2359 696 2363
rect 687 2358 696 2359
rect 927 2363 936 2364
rect 927 2359 928 2363
rect 935 2359 936 2363
rect 940 2362 942 2368
rect 3838 2368 3839 2372
rect 3843 2368 3844 2372
rect 3838 2367 3844 2368
rect 4698 2371 4704 2372
rect 4698 2367 4699 2371
rect 4703 2367 4704 2371
rect 4698 2366 4704 2367
rect 4834 2371 4840 2372
rect 4834 2367 4835 2371
rect 4839 2367 4840 2371
rect 4834 2366 4840 2367
rect 4970 2371 4976 2372
rect 4970 2367 4971 2371
rect 4975 2367 4976 2371
rect 4970 2366 4976 2367
rect 5106 2371 5112 2372
rect 5106 2367 5107 2371
rect 5111 2367 5112 2371
rect 5106 2366 5112 2367
rect 5242 2371 5248 2372
rect 5242 2367 5243 2371
rect 5247 2367 5248 2371
rect 5242 2366 5248 2367
rect 5378 2371 5384 2372
rect 5378 2367 5379 2371
rect 5383 2367 5384 2371
rect 5378 2366 5384 2367
rect 5514 2371 5520 2372
rect 5514 2367 5515 2371
rect 5519 2367 5520 2371
rect 5662 2368 5663 2372
rect 5667 2368 5668 2372
rect 5662 2367 5668 2368
rect 5514 2366 5520 2367
rect 1167 2363 1173 2364
rect 1167 2362 1168 2363
rect 940 2360 1168 2362
rect 927 2358 936 2359
rect 1167 2359 1168 2360
rect 1172 2359 1173 2363
rect 1167 2358 1173 2359
rect 1415 2363 1421 2364
rect 1415 2359 1416 2363
rect 1420 2362 1421 2363
rect 1438 2363 1444 2364
rect 1438 2362 1439 2363
rect 1420 2360 1439 2362
rect 1420 2359 1421 2360
rect 1415 2358 1421 2359
rect 1438 2359 1439 2360
rect 1443 2359 1444 2363
rect 1438 2358 1444 2359
rect 1671 2363 1680 2364
rect 1671 2359 1672 2363
rect 1679 2359 1680 2363
rect 1671 2358 1680 2359
rect 1874 2363 1880 2364
rect 1874 2359 1875 2363
rect 1879 2362 1880 2363
rect 1911 2363 1917 2364
rect 1911 2362 1912 2363
rect 1879 2360 1912 2362
rect 1879 2359 1880 2360
rect 1874 2358 1880 2359
rect 1911 2359 1912 2360
rect 1916 2359 1917 2363
rect 1911 2358 1917 2359
rect 110 2356 116 2357
rect 1934 2356 1940 2357
rect 4726 2356 4732 2357
rect 110 2352 111 2356
rect 115 2352 116 2356
rect 110 2351 116 2352
rect 130 2355 136 2356
rect 130 2351 131 2355
rect 135 2351 136 2355
rect 130 2350 136 2351
rect 338 2355 344 2356
rect 338 2351 339 2355
rect 343 2351 344 2355
rect 338 2350 344 2351
rect 562 2355 568 2356
rect 562 2351 563 2355
rect 567 2351 568 2355
rect 562 2350 568 2351
rect 802 2355 808 2356
rect 802 2351 803 2355
rect 807 2351 808 2355
rect 802 2350 808 2351
rect 1042 2355 1048 2356
rect 1042 2351 1043 2355
rect 1047 2351 1048 2355
rect 1042 2350 1048 2351
rect 1290 2355 1296 2356
rect 1290 2351 1291 2355
rect 1295 2351 1296 2355
rect 1290 2350 1296 2351
rect 1546 2355 1552 2356
rect 1546 2351 1547 2355
rect 1551 2351 1552 2355
rect 1546 2350 1552 2351
rect 1786 2355 1792 2356
rect 1786 2351 1787 2355
rect 1791 2351 1792 2355
rect 1934 2352 1935 2356
rect 1939 2352 1940 2356
rect 1934 2351 1940 2352
rect 3838 2355 3844 2356
rect 3838 2351 3839 2355
rect 3843 2351 3844 2355
rect 4726 2352 4727 2356
rect 4731 2352 4732 2356
rect 4726 2351 4732 2352
rect 4862 2356 4868 2357
rect 4862 2352 4863 2356
rect 4867 2352 4868 2356
rect 4862 2351 4868 2352
rect 4998 2356 5004 2357
rect 4998 2352 4999 2356
rect 5003 2352 5004 2356
rect 4998 2351 5004 2352
rect 5134 2356 5140 2357
rect 5134 2352 5135 2356
rect 5139 2352 5140 2356
rect 5134 2351 5140 2352
rect 5270 2356 5276 2357
rect 5270 2352 5271 2356
rect 5275 2352 5276 2356
rect 5270 2351 5276 2352
rect 5406 2356 5412 2357
rect 5406 2352 5407 2356
rect 5411 2352 5412 2356
rect 5406 2351 5412 2352
rect 5542 2356 5548 2357
rect 5542 2352 5543 2356
rect 5547 2352 5548 2356
rect 5542 2351 5548 2352
rect 5662 2355 5668 2356
rect 5662 2351 5663 2355
rect 5667 2351 5668 2355
rect 1786 2350 1792 2351
rect 3838 2350 3844 2351
rect 5662 2350 5668 2351
rect 158 2340 164 2341
rect 110 2339 116 2340
rect 110 2335 111 2339
rect 115 2335 116 2339
rect 158 2336 159 2340
rect 163 2336 164 2340
rect 158 2335 164 2336
rect 366 2340 372 2341
rect 366 2336 367 2340
rect 371 2336 372 2340
rect 366 2335 372 2336
rect 590 2340 596 2341
rect 590 2336 591 2340
rect 595 2336 596 2340
rect 590 2335 596 2336
rect 830 2340 836 2341
rect 830 2336 831 2340
rect 835 2336 836 2340
rect 830 2335 836 2336
rect 1070 2340 1076 2341
rect 1070 2336 1071 2340
rect 1075 2336 1076 2340
rect 1070 2335 1076 2336
rect 1318 2340 1324 2341
rect 1318 2336 1319 2340
rect 1323 2336 1324 2340
rect 1318 2335 1324 2336
rect 1574 2340 1580 2341
rect 1574 2336 1575 2340
rect 1579 2336 1580 2340
rect 1574 2335 1580 2336
rect 1814 2340 1820 2341
rect 1814 2336 1815 2340
rect 1819 2336 1820 2340
rect 1814 2335 1820 2336
rect 1934 2339 1940 2340
rect 1934 2335 1935 2339
rect 1939 2335 1940 2339
rect 110 2334 116 2335
rect 1934 2334 1940 2335
rect 1974 2325 1980 2326
rect 3798 2325 3804 2326
rect 1974 2321 1975 2325
rect 1979 2321 1980 2325
rect 1974 2320 1980 2321
rect 2222 2324 2228 2325
rect 2222 2320 2223 2324
rect 2227 2320 2228 2324
rect 2222 2319 2228 2320
rect 2502 2324 2508 2325
rect 2502 2320 2503 2324
rect 2507 2320 2508 2324
rect 2502 2319 2508 2320
rect 2766 2324 2772 2325
rect 2766 2320 2767 2324
rect 2771 2320 2772 2324
rect 2766 2319 2772 2320
rect 3006 2324 3012 2325
rect 3006 2320 3007 2324
rect 3011 2320 3012 2324
rect 3006 2319 3012 2320
rect 3238 2324 3244 2325
rect 3238 2320 3239 2324
rect 3243 2320 3244 2324
rect 3238 2319 3244 2320
rect 3470 2324 3476 2325
rect 3470 2320 3471 2324
rect 3475 2320 3476 2324
rect 3470 2319 3476 2320
rect 3678 2324 3684 2325
rect 3678 2320 3679 2324
rect 3683 2320 3684 2324
rect 3798 2321 3799 2325
rect 3803 2321 3804 2325
rect 3798 2320 3804 2321
rect 3678 2319 3684 2320
rect 2194 2309 2200 2310
rect 1974 2308 1980 2309
rect 1974 2304 1975 2308
rect 1979 2304 1980 2308
rect 2194 2305 2195 2309
rect 2199 2305 2200 2309
rect 2194 2304 2200 2305
rect 2474 2309 2480 2310
rect 2474 2305 2475 2309
rect 2479 2305 2480 2309
rect 2474 2304 2480 2305
rect 2738 2309 2744 2310
rect 2738 2305 2739 2309
rect 2743 2305 2744 2309
rect 2738 2304 2744 2305
rect 2978 2309 2984 2310
rect 2978 2305 2979 2309
rect 2983 2305 2984 2309
rect 2978 2304 2984 2305
rect 3210 2309 3216 2310
rect 3210 2305 3211 2309
rect 3215 2305 3216 2309
rect 3210 2304 3216 2305
rect 3442 2309 3448 2310
rect 3442 2305 3443 2309
rect 3447 2305 3448 2309
rect 3442 2304 3448 2305
rect 3650 2309 3656 2310
rect 3650 2305 3651 2309
rect 3655 2305 3656 2309
rect 3650 2304 3656 2305
rect 3798 2308 3804 2309
rect 3798 2304 3799 2308
rect 3803 2304 3804 2308
rect 1974 2303 1980 2304
rect 3798 2303 3804 2304
rect 2298 2299 2304 2300
rect 2298 2295 2299 2299
rect 2303 2298 2304 2299
rect 2319 2299 2325 2300
rect 2319 2298 2320 2299
rect 2303 2296 2320 2298
rect 2303 2295 2304 2296
rect 2298 2294 2304 2295
rect 2319 2295 2320 2296
rect 2324 2295 2325 2299
rect 2319 2294 2325 2295
rect 2334 2299 2340 2300
rect 2334 2295 2335 2299
rect 2339 2298 2340 2299
rect 2599 2299 2605 2300
rect 2599 2298 2600 2299
rect 2339 2296 2600 2298
rect 2339 2295 2340 2296
rect 2334 2294 2340 2295
rect 2599 2295 2600 2296
rect 2604 2295 2605 2299
rect 2599 2294 2605 2295
rect 2863 2299 2869 2300
rect 2863 2295 2864 2299
rect 2868 2298 2869 2299
rect 2994 2299 3000 2300
rect 2994 2298 2995 2299
rect 2868 2296 2995 2298
rect 2868 2295 2869 2296
rect 2863 2294 2869 2295
rect 2994 2295 2995 2296
rect 2999 2295 3000 2299
rect 2994 2294 3000 2295
rect 3103 2299 3109 2300
rect 3103 2295 3104 2299
rect 3108 2298 3109 2299
rect 3226 2299 3232 2300
rect 3226 2298 3227 2299
rect 3108 2296 3227 2298
rect 3108 2295 3109 2296
rect 3103 2294 3109 2295
rect 3226 2295 3227 2296
rect 3231 2295 3232 2299
rect 3226 2294 3232 2295
rect 3335 2299 3341 2300
rect 3335 2295 3336 2299
rect 3340 2298 3341 2299
rect 3458 2299 3464 2300
rect 3458 2298 3459 2299
rect 3340 2296 3459 2298
rect 3340 2295 3341 2296
rect 3335 2294 3341 2295
rect 3458 2295 3459 2296
rect 3463 2295 3464 2299
rect 3458 2294 3464 2295
rect 3567 2299 3573 2300
rect 3567 2295 3568 2299
rect 3572 2298 3573 2299
rect 3666 2299 3672 2300
rect 3666 2298 3667 2299
rect 3572 2296 3667 2298
rect 3572 2295 3573 2296
rect 3567 2294 3573 2295
rect 3666 2295 3667 2296
rect 3671 2295 3672 2299
rect 3666 2294 3672 2295
rect 3754 2299 3760 2300
rect 3754 2295 3755 2299
rect 3759 2298 3760 2299
rect 3775 2299 3781 2300
rect 3775 2298 3776 2299
rect 3759 2296 3776 2298
rect 3759 2295 3760 2296
rect 3754 2294 3760 2295
rect 3775 2295 3776 2296
rect 3780 2295 3781 2299
rect 3775 2294 3781 2295
rect 287 2291 293 2292
rect 287 2287 288 2291
rect 292 2290 293 2291
rect 1246 2291 1252 2292
rect 1246 2290 1247 2291
rect 292 2288 1247 2290
rect 292 2287 293 2288
rect 287 2286 293 2287
rect 1246 2287 1247 2288
rect 1251 2287 1252 2291
rect 1246 2286 1252 2287
rect 2826 2291 2832 2292
rect 2826 2287 2827 2291
rect 2831 2290 2832 2291
rect 3738 2291 3744 2292
rect 3738 2290 3739 2291
rect 2831 2288 3739 2290
rect 2831 2287 2832 2288
rect 2826 2286 2832 2287
rect 3738 2287 3739 2288
rect 3743 2287 3744 2291
rect 3738 2286 3744 2287
rect 3838 2285 3844 2286
rect 5662 2285 5668 2286
rect 3838 2281 3839 2285
rect 3843 2281 3844 2285
rect 3838 2280 3844 2281
rect 3886 2284 3892 2285
rect 3886 2280 3887 2284
rect 3891 2280 3892 2284
rect 3886 2279 3892 2280
rect 4182 2284 4188 2285
rect 4182 2280 4183 2284
rect 4187 2280 4188 2284
rect 4182 2279 4188 2280
rect 4494 2284 4500 2285
rect 4494 2280 4495 2284
rect 4499 2280 4500 2284
rect 4494 2279 4500 2280
rect 4790 2284 4796 2285
rect 4790 2280 4791 2284
rect 4795 2280 4796 2284
rect 4790 2279 4796 2280
rect 5086 2284 5092 2285
rect 5086 2280 5087 2284
rect 5091 2280 5092 2284
rect 5086 2279 5092 2280
rect 5382 2284 5388 2285
rect 5382 2280 5383 2284
rect 5387 2280 5388 2284
rect 5662 2281 5663 2285
rect 5667 2281 5668 2285
rect 5662 2280 5668 2281
rect 5382 2279 5388 2280
rect 110 2277 116 2278
rect 1934 2277 1940 2278
rect 110 2273 111 2277
rect 115 2273 116 2277
rect 110 2272 116 2273
rect 158 2276 164 2277
rect 158 2272 159 2276
rect 163 2272 164 2276
rect 158 2271 164 2272
rect 318 2276 324 2277
rect 318 2272 319 2276
rect 323 2272 324 2276
rect 318 2271 324 2272
rect 550 2276 556 2277
rect 550 2272 551 2276
rect 555 2272 556 2276
rect 550 2271 556 2272
rect 830 2276 836 2277
rect 830 2272 831 2276
rect 835 2272 836 2276
rect 830 2271 836 2272
rect 1150 2276 1156 2277
rect 1150 2272 1151 2276
rect 1155 2272 1156 2276
rect 1150 2271 1156 2272
rect 1494 2276 1500 2277
rect 1494 2272 1495 2276
rect 1499 2272 1500 2276
rect 1494 2271 1500 2272
rect 1814 2276 1820 2277
rect 1814 2272 1815 2276
rect 1819 2272 1820 2276
rect 1934 2273 1935 2277
rect 1939 2273 1940 2277
rect 1934 2272 1940 2273
rect 1814 2271 1820 2272
rect 3858 2269 3864 2270
rect 3838 2268 3844 2269
rect 2334 2267 2340 2268
rect 2334 2266 2335 2267
rect 2285 2264 2335 2266
rect 2334 2263 2335 2264
rect 2339 2263 2340 2267
rect 2334 2262 2340 2263
rect 2562 2267 2568 2268
rect 2562 2263 2563 2267
rect 2567 2263 2568 2267
rect 2562 2262 2568 2263
rect 2826 2267 2832 2268
rect 2826 2263 2827 2267
rect 2831 2263 2832 2267
rect 2826 2262 2832 2263
rect 2994 2267 3000 2268
rect 2994 2263 2995 2267
rect 2999 2263 3000 2267
rect 2994 2262 3000 2263
rect 3226 2267 3232 2268
rect 3226 2263 3227 2267
rect 3231 2263 3232 2267
rect 3226 2262 3232 2263
rect 3458 2267 3464 2268
rect 3458 2263 3459 2267
rect 3463 2263 3464 2267
rect 3458 2262 3464 2263
rect 3666 2267 3672 2268
rect 3666 2263 3667 2267
rect 3671 2263 3672 2267
rect 3838 2264 3839 2268
rect 3843 2264 3844 2268
rect 3858 2265 3859 2269
rect 3863 2265 3864 2269
rect 3858 2264 3864 2265
rect 4154 2269 4160 2270
rect 4154 2265 4155 2269
rect 4159 2265 4160 2269
rect 4154 2264 4160 2265
rect 4466 2269 4472 2270
rect 4466 2265 4467 2269
rect 4471 2265 4472 2269
rect 4466 2264 4472 2265
rect 4762 2269 4768 2270
rect 4762 2265 4763 2269
rect 4767 2265 4768 2269
rect 4762 2264 4768 2265
rect 5058 2269 5064 2270
rect 5058 2265 5059 2269
rect 5063 2265 5064 2269
rect 5058 2264 5064 2265
rect 5354 2269 5360 2270
rect 5354 2265 5355 2269
rect 5359 2265 5360 2269
rect 5354 2264 5360 2265
rect 5662 2268 5668 2269
rect 5662 2264 5663 2268
rect 5667 2264 5668 2268
rect 3838 2263 3844 2264
rect 5662 2263 5668 2264
rect 3666 2262 3672 2263
rect 130 2261 136 2262
rect 110 2260 116 2261
rect 110 2256 111 2260
rect 115 2256 116 2260
rect 130 2257 131 2261
rect 135 2257 136 2261
rect 130 2256 136 2257
rect 290 2261 296 2262
rect 290 2257 291 2261
rect 295 2257 296 2261
rect 290 2256 296 2257
rect 522 2261 528 2262
rect 522 2257 523 2261
rect 527 2257 528 2261
rect 522 2256 528 2257
rect 802 2261 808 2262
rect 802 2257 803 2261
rect 807 2257 808 2261
rect 802 2256 808 2257
rect 1122 2261 1128 2262
rect 1122 2257 1123 2261
rect 1127 2257 1128 2261
rect 1122 2256 1128 2257
rect 1466 2261 1472 2262
rect 1466 2257 1467 2261
rect 1471 2257 1472 2261
rect 1466 2256 1472 2257
rect 1786 2261 1792 2262
rect 1786 2257 1787 2261
rect 1791 2257 1792 2261
rect 1786 2256 1792 2257
rect 1934 2260 1940 2261
rect 1934 2256 1935 2260
rect 1939 2256 1940 2260
rect 110 2255 116 2256
rect 1934 2255 1940 2256
rect 3962 2259 3968 2260
rect 3962 2255 3963 2259
rect 3967 2258 3968 2259
rect 3983 2259 3989 2260
rect 3983 2258 3984 2259
rect 3967 2256 3984 2258
rect 3967 2255 3968 2256
rect 3962 2254 3968 2255
rect 3983 2255 3984 2256
rect 3988 2255 3989 2259
rect 3983 2254 3989 2255
rect 4279 2259 4285 2260
rect 4279 2255 4280 2259
rect 4284 2258 4285 2259
rect 4482 2259 4488 2260
rect 4482 2258 4483 2259
rect 4284 2256 4483 2258
rect 4284 2255 4285 2256
rect 4279 2254 4285 2255
rect 4482 2255 4483 2256
rect 4487 2255 4488 2259
rect 4482 2254 4488 2255
rect 4591 2259 4597 2260
rect 4591 2255 4592 2259
rect 4596 2258 4597 2259
rect 4626 2259 4632 2260
rect 4626 2258 4627 2259
rect 4596 2256 4627 2258
rect 4596 2255 4597 2256
rect 4591 2254 4597 2255
rect 4626 2255 4627 2256
rect 4631 2255 4632 2259
rect 4887 2259 4893 2260
rect 4887 2258 4888 2259
rect 4626 2254 4632 2255
rect 4819 2256 4888 2258
rect 255 2251 261 2252
rect 255 2247 256 2251
rect 260 2250 261 2251
rect 306 2251 312 2252
rect 306 2250 307 2251
rect 260 2248 307 2250
rect 260 2247 261 2248
rect 255 2246 261 2247
rect 306 2247 307 2248
rect 311 2247 312 2251
rect 306 2246 312 2247
rect 415 2251 421 2252
rect 415 2247 416 2251
rect 420 2250 421 2251
rect 538 2251 544 2252
rect 538 2250 539 2251
rect 420 2248 539 2250
rect 420 2247 421 2248
rect 415 2246 421 2247
rect 538 2247 539 2248
rect 543 2247 544 2251
rect 538 2246 544 2247
rect 647 2251 653 2252
rect 647 2247 648 2251
rect 652 2250 653 2251
rect 818 2251 824 2252
rect 818 2250 819 2251
rect 652 2248 819 2250
rect 652 2247 653 2248
rect 647 2246 653 2247
rect 818 2247 819 2248
rect 823 2247 824 2251
rect 818 2246 824 2247
rect 927 2251 933 2252
rect 927 2247 928 2251
rect 932 2247 933 2251
rect 927 2246 933 2247
rect 1246 2251 1253 2252
rect 1246 2247 1247 2251
rect 1252 2247 1253 2251
rect 1246 2246 1253 2247
rect 1266 2251 1272 2252
rect 1266 2247 1267 2251
rect 1271 2250 1272 2251
rect 1591 2251 1597 2252
rect 1591 2250 1592 2251
rect 1271 2248 1592 2250
rect 1271 2247 1272 2248
rect 1266 2246 1272 2247
rect 1591 2247 1592 2248
rect 1596 2247 1597 2251
rect 1591 2246 1597 2247
rect 1911 2251 1920 2252
rect 1911 2247 1912 2251
rect 1919 2247 1920 2251
rect 1911 2246 1920 2247
rect 4242 2251 4248 2252
rect 4242 2247 4243 2251
rect 4247 2250 4248 2251
rect 4819 2250 4821 2256
rect 4887 2255 4888 2256
rect 4892 2255 4893 2259
rect 4887 2254 4893 2255
rect 5002 2259 5008 2260
rect 5002 2255 5003 2259
rect 5007 2258 5008 2259
rect 5183 2259 5189 2260
rect 5183 2258 5184 2259
rect 5007 2256 5184 2258
rect 5007 2255 5008 2256
rect 5002 2254 5008 2255
rect 5183 2255 5184 2256
rect 5188 2255 5189 2259
rect 5183 2254 5189 2255
rect 5278 2259 5284 2260
rect 5278 2255 5279 2259
rect 5283 2258 5284 2259
rect 5479 2259 5485 2260
rect 5479 2258 5480 2259
rect 5283 2256 5480 2258
rect 5283 2255 5284 2256
rect 5278 2254 5284 2255
rect 5479 2255 5480 2256
rect 5484 2255 5485 2259
rect 5479 2254 5485 2255
rect 4247 2248 4821 2250
rect 4247 2247 4248 2248
rect 4242 2246 4248 2247
rect 218 2243 224 2244
rect 218 2239 219 2243
rect 223 2242 224 2243
rect 929 2242 931 2246
rect 223 2240 931 2242
rect 223 2239 224 2240
rect 218 2238 224 2239
rect 3778 2227 3784 2228
rect 3778 2223 3779 2227
rect 3783 2226 3784 2227
rect 4242 2227 4248 2228
rect 3783 2224 3877 2226
rect 3783 2223 3784 2224
rect 3778 2222 3784 2223
rect 4242 2223 4243 2227
rect 4247 2223 4248 2227
rect 4242 2222 4248 2223
rect 4482 2227 4488 2228
rect 4482 2223 4483 2227
rect 4487 2223 4488 2227
rect 5002 2227 5008 2228
rect 5002 2226 5003 2227
rect 4853 2224 5003 2226
rect 4482 2222 4488 2223
rect 5002 2223 5003 2224
rect 5007 2223 5008 2227
rect 5278 2227 5284 2228
rect 5278 2226 5279 2227
rect 5149 2224 5279 2226
rect 5002 2222 5008 2223
rect 5278 2223 5279 2224
rect 5283 2223 5284 2227
rect 5278 2222 5284 2223
rect 5370 2227 5376 2228
rect 5370 2223 5371 2227
rect 5375 2223 5376 2227
rect 5370 2222 5376 2223
rect 287 2219 293 2220
rect 287 2218 288 2219
rect 221 2216 288 2218
rect 287 2215 288 2216
rect 292 2215 293 2219
rect 287 2214 293 2215
rect 306 2219 312 2220
rect 306 2215 307 2219
rect 311 2215 312 2219
rect 306 2214 312 2215
rect 538 2219 544 2220
rect 538 2215 539 2219
rect 543 2215 544 2219
rect 538 2214 544 2215
rect 818 2219 824 2220
rect 818 2215 819 2219
rect 823 2215 824 2219
rect 1266 2219 1272 2220
rect 1266 2218 1267 2219
rect 1213 2216 1267 2218
rect 818 2214 824 2215
rect 1266 2215 1267 2216
rect 1271 2215 1272 2219
rect 1266 2214 1272 2215
rect 1274 2219 1280 2220
rect 1274 2215 1275 2219
rect 1279 2218 1280 2219
rect 1874 2219 1880 2220
rect 1279 2216 1485 2218
rect 1279 2215 1280 2216
rect 1274 2214 1280 2215
rect 1874 2215 1875 2219
rect 1879 2215 1880 2219
rect 1874 2214 1880 2215
rect 1914 2219 1920 2220
rect 1914 2215 1915 2219
rect 1919 2218 1920 2219
rect 2122 2219 2128 2220
rect 1919 2216 2013 2218
rect 1919 2215 1920 2216
rect 1914 2214 1920 2215
rect 2122 2215 2123 2219
rect 2127 2218 2128 2219
rect 2287 2219 2293 2220
rect 2127 2216 2173 2218
rect 2127 2215 2128 2216
rect 2122 2214 2128 2215
rect 2287 2215 2288 2219
rect 2292 2218 2293 2219
rect 2514 2219 2520 2220
rect 2292 2216 2405 2218
rect 2292 2215 2293 2216
rect 2287 2214 2293 2215
rect 2514 2215 2515 2219
rect 2519 2218 2520 2219
rect 2794 2219 2800 2220
rect 2519 2216 2685 2218
rect 2519 2215 2520 2216
rect 2514 2214 2520 2215
rect 2794 2215 2795 2219
rect 2799 2218 2800 2219
rect 3114 2219 3120 2220
rect 2799 2216 3005 2218
rect 2799 2215 2800 2216
rect 2794 2214 2800 2215
rect 3114 2215 3115 2219
rect 3119 2218 3120 2219
rect 3754 2219 3760 2220
rect 3754 2218 3755 2219
rect 3119 2216 3349 2218
rect 3741 2216 3755 2218
rect 3119 2215 3120 2216
rect 3114 2214 3120 2215
rect 3754 2215 3755 2216
rect 3759 2215 3760 2219
rect 3754 2214 3760 2215
rect 2562 2191 2568 2192
rect 2562 2187 2563 2191
rect 2567 2190 2568 2191
rect 2567 2188 3141 2190
rect 2567 2187 2568 2188
rect 2562 2186 2568 2187
rect 2119 2183 2128 2184
rect 2119 2179 2120 2183
rect 2127 2179 2128 2183
rect 2119 2178 2128 2179
rect 2279 2183 2285 2184
rect 2279 2179 2280 2183
rect 2284 2182 2285 2183
rect 2287 2183 2293 2184
rect 2287 2182 2288 2183
rect 2284 2180 2288 2182
rect 2284 2179 2285 2180
rect 2279 2178 2285 2179
rect 2287 2179 2288 2180
rect 2292 2179 2293 2183
rect 2287 2178 2293 2179
rect 2511 2183 2520 2184
rect 2511 2179 2512 2183
rect 2519 2179 2520 2183
rect 2511 2178 2520 2179
rect 2791 2183 2800 2184
rect 2791 2179 2792 2183
rect 2799 2179 2800 2183
rect 2791 2178 2800 2179
rect 3111 2183 3120 2184
rect 3111 2179 3112 2183
rect 3119 2179 3120 2183
rect 3139 2182 3141 2188
rect 3455 2183 3461 2184
rect 3455 2182 3456 2183
rect 3139 2180 3456 2182
rect 3111 2178 3120 2179
rect 3455 2179 3456 2180
rect 3460 2179 3461 2183
rect 3455 2178 3461 2179
rect 3775 2183 3784 2184
rect 3775 2179 3776 2183
rect 3783 2179 3784 2183
rect 3775 2178 3784 2179
rect 1974 2176 1980 2177
rect 3798 2176 3804 2177
rect 1974 2172 1975 2176
rect 1979 2172 1980 2176
rect 1974 2171 1980 2172
rect 1994 2175 2000 2176
rect 1994 2171 1995 2175
rect 1999 2171 2000 2175
rect 1994 2170 2000 2171
rect 2154 2175 2160 2176
rect 2154 2171 2155 2175
rect 2159 2171 2160 2175
rect 2154 2170 2160 2171
rect 2386 2175 2392 2176
rect 2386 2171 2387 2175
rect 2391 2171 2392 2175
rect 2386 2170 2392 2171
rect 2666 2175 2672 2176
rect 2666 2171 2667 2175
rect 2671 2171 2672 2175
rect 2666 2170 2672 2171
rect 2986 2175 2992 2176
rect 2986 2171 2987 2175
rect 2991 2171 2992 2175
rect 2986 2170 2992 2171
rect 3330 2175 3336 2176
rect 3330 2171 3331 2175
rect 3335 2171 3336 2175
rect 3330 2170 3336 2171
rect 3650 2175 3656 2176
rect 3650 2171 3651 2175
rect 3655 2171 3656 2175
rect 3798 2172 3799 2176
rect 3803 2172 3804 2176
rect 3962 2175 3968 2176
rect 3962 2174 3963 2175
rect 3949 2172 3963 2174
rect 3798 2171 3804 2172
rect 3962 2171 3963 2172
rect 3967 2171 3968 2175
rect 3650 2170 3656 2171
rect 3962 2170 3968 2171
rect 3986 2175 3992 2176
rect 3986 2171 3987 2175
rect 3991 2174 3992 2175
rect 4127 2175 4133 2176
rect 3991 2172 4013 2174
rect 3991 2171 3992 2172
rect 3986 2170 3992 2171
rect 4127 2171 4128 2175
rect 4132 2174 4133 2175
rect 4263 2175 4269 2176
rect 4132 2172 4149 2174
rect 4132 2171 4133 2172
rect 4127 2170 4133 2171
rect 4263 2171 4264 2175
rect 4268 2174 4269 2175
rect 4399 2175 4405 2176
rect 4268 2172 4285 2174
rect 4268 2171 4269 2172
rect 4263 2170 4269 2171
rect 4399 2171 4400 2175
rect 4404 2174 4405 2175
rect 4666 2175 4672 2176
rect 4404 2172 4421 2174
rect 4404 2171 4405 2172
rect 4399 2170 4405 2171
rect 4626 2171 4632 2172
rect 4626 2167 4627 2171
rect 4631 2167 4632 2171
rect 4666 2171 4667 2175
rect 4671 2174 4672 2175
rect 4826 2175 4832 2176
rect 4671 2172 4717 2174
rect 4671 2171 4672 2172
rect 4666 2170 4672 2171
rect 4826 2171 4827 2175
rect 4831 2174 4832 2175
rect 5018 2175 5024 2176
rect 4831 2172 4909 2174
rect 4831 2171 4832 2172
rect 4826 2170 4832 2171
rect 5018 2171 5019 2175
rect 5023 2174 5024 2175
rect 5231 2175 5237 2176
rect 5023 2172 5117 2174
rect 5023 2171 5024 2172
rect 5018 2170 5024 2171
rect 5231 2171 5232 2175
rect 5236 2174 5237 2175
rect 5618 2175 5624 2176
rect 5618 2174 5619 2175
rect 5236 2172 5333 2174
rect 5605 2172 5619 2174
rect 5236 2171 5237 2172
rect 5231 2170 5237 2171
rect 5618 2171 5619 2172
rect 5623 2171 5624 2175
rect 5618 2170 5624 2171
rect 4626 2166 4632 2167
rect 2022 2160 2028 2161
rect 1974 2159 1980 2160
rect 1974 2155 1975 2159
rect 1979 2155 1980 2159
rect 2022 2156 2023 2160
rect 2027 2156 2028 2160
rect 2022 2155 2028 2156
rect 2182 2160 2188 2161
rect 2182 2156 2183 2160
rect 2187 2156 2188 2160
rect 2182 2155 2188 2156
rect 2414 2160 2420 2161
rect 2414 2156 2415 2160
rect 2419 2156 2420 2160
rect 2414 2155 2420 2156
rect 2694 2160 2700 2161
rect 2694 2156 2695 2160
rect 2699 2156 2700 2160
rect 2694 2155 2700 2156
rect 3014 2160 3020 2161
rect 3014 2156 3015 2160
rect 3019 2156 3020 2160
rect 3014 2155 3020 2156
rect 3358 2160 3364 2161
rect 3358 2156 3359 2160
rect 3363 2156 3364 2160
rect 3358 2155 3364 2156
rect 3678 2160 3684 2161
rect 3678 2156 3679 2160
rect 3683 2156 3684 2160
rect 3678 2155 3684 2156
rect 3798 2159 3804 2160
rect 3798 2155 3799 2159
rect 3803 2155 3804 2159
rect 1974 2154 1980 2155
rect 3798 2154 3804 2155
rect 418 2147 424 2148
rect 418 2143 419 2147
rect 423 2146 424 2147
rect 871 2147 877 2148
rect 871 2146 872 2147
rect 423 2144 501 2146
rect 781 2144 872 2146
rect 423 2143 424 2144
rect 418 2142 424 2143
rect 871 2143 872 2144
rect 876 2143 877 2147
rect 1018 2147 1024 2148
rect 871 2142 877 2143
rect 1002 2143 1008 2144
rect 376 2130 378 2141
rect 1002 2139 1003 2143
rect 1007 2139 1008 2143
rect 1018 2143 1019 2147
rect 1023 2146 1024 2147
rect 1614 2147 1620 2148
rect 1614 2146 1615 2147
rect 1023 2144 1165 2146
rect 1477 2144 1615 2146
rect 1023 2143 1024 2144
rect 1018 2142 1024 2143
rect 1614 2143 1615 2144
rect 1619 2143 1620 2147
rect 1614 2142 1620 2143
rect 1626 2147 1632 2148
rect 1626 2143 1627 2147
rect 1631 2146 1632 2147
rect 1631 2144 1653 2146
rect 1631 2143 1632 2144
rect 1626 2142 1632 2143
rect 1002 2138 1008 2139
rect 3983 2139 3992 2140
rect 3983 2135 3984 2139
rect 3991 2135 3992 2139
rect 3983 2134 3992 2135
rect 4119 2139 4125 2140
rect 4119 2135 4120 2139
rect 4124 2138 4125 2139
rect 4127 2139 4133 2140
rect 4127 2138 4128 2139
rect 4124 2136 4128 2138
rect 4124 2135 4125 2136
rect 4119 2134 4125 2135
rect 4127 2135 4128 2136
rect 4132 2135 4133 2139
rect 4127 2134 4133 2135
rect 4255 2139 4261 2140
rect 4255 2135 4256 2139
rect 4260 2138 4261 2139
rect 4263 2139 4269 2140
rect 4263 2138 4264 2139
rect 4260 2136 4264 2138
rect 4260 2135 4261 2136
rect 4255 2134 4261 2135
rect 4263 2135 4264 2136
rect 4268 2135 4269 2139
rect 4263 2134 4269 2135
rect 4391 2139 4397 2140
rect 4391 2135 4392 2139
rect 4396 2138 4397 2139
rect 4399 2139 4405 2140
rect 4399 2138 4400 2139
rect 4396 2136 4400 2138
rect 4396 2135 4397 2136
rect 4391 2134 4397 2135
rect 4399 2135 4400 2136
rect 4404 2135 4405 2139
rect 4399 2134 4405 2135
rect 4490 2139 4496 2140
rect 4490 2135 4491 2139
rect 4495 2138 4496 2139
rect 4527 2139 4533 2140
rect 4527 2138 4528 2139
rect 4495 2136 4528 2138
rect 4495 2135 4496 2136
rect 4490 2134 4496 2135
rect 4527 2135 4528 2136
rect 4532 2135 4533 2139
rect 4527 2134 4533 2135
rect 4663 2139 4672 2140
rect 4663 2135 4664 2139
rect 4671 2135 4672 2139
rect 4663 2134 4672 2135
rect 4823 2139 4832 2140
rect 4823 2135 4824 2139
rect 4831 2135 4832 2139
rect 4823 2134 4832 2135
rect 5015 2139 5024 2140
rect 5015 2135 5016 2139
rect 5023 2135 5024 2139
rect 5015 2134 5024 2135
rect 5223 2139 5229 2140
rect 5223 2135 5224 2139
rect 5228 2138 5229 2139
rect 5231 2139 5237 2140
rect 5231 2138 5232 2139
rect 5228 2136 5232 2138
rect 5228 2135 5229 2136
rect 5223 2134 5229 2135
rect 5231 2135 5232 2136
rect 5236 2135 5237 2139
rect 5231 2134 5237 2135
rect 5354 2139 5360 2140
rect 5354 2135 5355 2139
rect 5359 2138 5360 2139
rect 5439 2139 5445 2140
rect 5439 2138 5440 2139
rect 5359 2136 5440 2138
rect 5359 2135 5360 2136
rect 5354 2134 5360 2135
rect 5439 2135 5440 2136
rect 5444 2135 5445 2139
rect 5439 2134 5445 2135
rect 5618 2139 5624 2140
rect 5618 2135 5619 2139
rect 5623 2138 5624 2139
rect 5639 2139 5645 2140
rect 5639 2138 5640 2139
rect 5623 2136 5640 2138
rect 5623 2135 5624 2136
rect 5618 2134 5624 2135
rect 5639 2135 5640 2136
rect 5644 2135 5645 2139
rect 5639 2134 5645 2135
rect 3838 2132 3844 2133
rect 5662 2132 5668 2133
rect 814 2131 820 2132
rect 814 2130 815 2131
rect 376 2128 815 2130
rect 814 2127 815 2128
rect 819 2127 820 2131
rect 3838 2128 3839 2132
rect 3843 2128 3844 2132
rect 3838 2127 3844 2128
rect 3858 2131 3864 2132
rect 3858 2127 3859 2131
rect 3863 2127 3864 2131
rect 814 2126 820 2127
rect 3858 2126 3864 2127
rect 3994 2131 4000 2132
rect 3994 2127 3995 2131
rect 3999 2127 4000 2131
rect 3994 2126 4000 2127
rect 4130 2131 4136 2132
rect 4130 2127 4131 2131
rect 4135 2127 4136 2131
rect 4130 2126 4136 2127
rect 4266 2131 4272 2132
rect 4266 2127 4267 2131
rect 4271 2127 4272 2131
rect 4266 2126 4272 2127
rect 4402 2131 4408 2132
rect 4402 2127 4403 2131
rect 4407 2127 4408 2131
rect 4402 2126 4408 2127
rect 4538 2131 4544 2132
rect 4538 2127 4539 2131
rect 4543 2127 4544 2131
rect 4538 2126 4544 2127
rect 4698 2131 4704 2132
rect 4698 2127 4699 2131
rect 4703 2127 4704 2131
rect 4698 2126 4704 2127
rect 4890 2131 4896 2132
rect 4890 2127 4891 2131
rect 4895 2127 4896 2131
rect 4890 2126 4896 2127
rect 5098 2131 5104 2132
rect 5098 2127 5099 2131
rect 5103 2127 5104 2131
rect 5098 2126 5104 2127
rect 5314 2131 5320 2132
rect 5314 2127 5315 2131
rect 5319 2127 5320 2131
rect 5314 2126 5320 2127
rect 5514 2131 5520 2132
rect 5514 2127 5515 2131
rect 5519 2127 5520 2131
rect 5662 2128 5663 2132
rect 5667 2128 5668 2132
rect 5662 2127 5668 2128
rect 5514 2126 5520 2127
rect 1018 2119 1024 2120
rect 1018 2118 1019 2119
rect 619 2116 1019 2118
rect 415 2111 424 2112
rect 415 2107 416 2111
rect 423 2107 424 2111
rect 415 2106 424 2107
rect 607 2111 613 2112
rect 607 2107 608 2111
rect 612 2110 613 2111
rect 619 2110 621 2116
rect 1018 2115 1019 2116
rect 1023 2115 1024 2119
rect 3886 2116 3892 2117
rect 1018 2114 1024 2115
rect 3838 2115 3844 2116
rect 612 2108 621 2110
rect 814 2111 821 2112
rect 612 2107 613 2108
rect 607 2106 613 2107
rect 814 2107 815 2111
rect 820 2107 821 2111
rect 814 2106 821 2107
rect 871 2111 877 2112
rect 871 2107 872 2111
rect 876 2110 877 2111
rect 1039 2111 1045 2112
rect 1039 2110 1040 2111
rect 876 2108 1040 2110
rect 876 2107 877 2108
rect 871 2106 877 2107
rect 1039 2107 1040 2108
rect 1044 2107 1045 2111
rect 1039 2106 1045 2107
rect 1271 2111 1280 2112
rect 1271 2107 1272 2111
rect 1279 2107 1280 2111
rect 1271 2106 1280 2107
rect 1458 2111 1464 2112
rect 1458 2107 1459 2111
rect 1463 2110 1464 2111
rect 1511 2111 1517 2112
rect 1511 2110 1512 2111
rect 1463 2108 1512 2110
rect 1463 2107 1464 2108
rect 1458 2106 1464 2107
rect 1511 2107 1512 2108
rect 1516 2107 1517 2111
rect 1511 2106 1517 2107
rect 1614 2111 1620 2112
rect 1614 2107 1615 2111
rect 1619 2110 1620 2111
rect 1759 2111 1765 2112
rect 1759 2110 1760 2111
rect 1619 2108 1760 2110
rect 1619 2107 1620 2108
rect 1614 2106 1620 2107
rect 1759 2107 1760 2108
rect 1764 2107 1765 2111
rect 3838 2111 3839 2115
rect 3843 2111 3844 2115
rect 3886 2112 3887 2116
rect 3891 2112 3892 2116
rect 3886 2111 3892 2112
rect 4022 2116 4028 2117
rect 4022 2112 4023 2116
rect 4027 2112 4028 2116
rect 4022 2111 4028 2112
rect 4158 2116 4164 2117
rect 4158 2112 4159 2116
rect 4163 2112 4164 2116
rect 4158 2111 4164 2112
rect 4294 2116 4300 2117
rect 4294 2112 4295 2116
rect 4299 2112 4300 2116
rect 4294 2111 4300 2112
rect 4430 2116 4436 2117
rect 4430 2112 4431 2116
rect 4435 2112 4436 2116
rect 4430 2111 4436 2112
rect 4566 2116 4572 2117
rect 4566 2112 4567 2116
rect 4571 2112 4572 2116
rect 4566 2111 4572 2112
rect 4726 2116 4732 2117
rect 4726 2112 4727 2116
rect 4731 2112 4732 2116
rect 4726 2111 4732 2112
rect 4918 2116 4924 2117
rect 4918 2112 4919 2116
rect 4923 2112 4924 2116
rect 4918 2111 4924 2112
rect 5126 2116 5132 2117
rect 5126 2112 5127 2116
rect 5131 2112 5132 2116
rect 5126 2111 5132 2112
rect 5342 2116 5348 2117
rect 5342 2112 5343 2116
rect 5347 2112 5348 2116
rect 5342 2111 5348 2112
rect 5542 2116 5548 2117
rect 5542 2112 5543 2116
rect 5547 2112 5548 2116
rect 5542 2111 5548 2112
rect 5662 2115 5668 2116
rect 5662 2111 5663 2115
rect 5667 2111 5668 2115
rect 3838 2110 3844 2111
rect 5662 2110 5668 2111
rect 1759 2106 1765 2107
rect 110 2104 116 2105
rect 1934 2104 1940 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 290 2103 296 2104
rect 290 2099 291 2103
rect 295 2099 296 2103
rect 290 2098 296 2099
rect 482 2103 488 2104
rect 482 2099 483 2103
rect 487 2099 488 2103
rect 482 2098 488 2099
rect 690 2103 696 2104
rect 690 2099 691 2103
rect 695 2099 696 2103
rect 690 2098 696 2099
rect 914 2103 920 2104
rect 914 2099 915 2103
rect 919 2099 920 2103
rect 914 2098 920 2099
rect 1146 2103 1152 2104
rect 1146 2099 1147 2103
rect 1151 2099 1152 2103
rect 1146 2098 1152 2099
rect 1386 2103 1392 2104
rect 1386 2099 1387 2103
rect 1391 2099 1392 2103
rect 1386 2098 1392 2099
rect 1634 2103 1640 2104
rect 1634 2099 1635 2103
rect 1639 2099 1640 2103
rect 1934 2100 1935 2104
rect 1939 2100 1940 2104
rect 1934 2099 1940 2100
rect 1634 2098 1640 2099
rect 318 2088 324 2089
rect 110 2087 116 2088
rect 110 2083 111 2087
rect 115 2083 116 2087
rect 318 2084 319 2088
rect 323 2084 324 2088
rect 318 2083 324 2084
rect 510 2088 516 2089
rect 510 2084 511 2088
rect 515 2084 516 2088
rect 510 2083 516 2084
rect 718 2088 724 2089
rect 718 2084 719 2088
rect 723 2084 724 2088
rect 718 2083 724 2084
rect 942 2088 948 2089
rect 942 2084 943 2088
rect 947 2084 948 2088
rect 942 2083 948 2084
rect 1174 2088 1180 2089
rect 1174 2084 1175 2088
rect 1179 2084 1180 2088
rect 1174 2083 1180 2084
rect 1414 2088 1420 2089
rect 1414 2084 1415 2088
rect 1419 2084 1420 2088
rect 1414 2083 1420 2084
rect 1662 2088 1668 2089
rect 1662 2084 1663 2088
rect 1667 2084 1668 2088
rect 1662 2083 1668 2084
rect 1934 2087 1940 2088
rect 1934 2083 1935 2087
rect 1939 2083 1940 2087
rect 110 2082 116 2083
rect 1934 2082 1940 2083
rect 3838 2037 3844 2038
rect 5662 2037 5668 2038
rect 3838 2033 3839 2037
rect 3843 2033 3844 2037
rect 3838 2032 3844 2033
rect 3886 2036 3892 2037
rect 3886 2032 3887 2036
rect 3891 2032 3892 2036
rect 3886 2031 3892 2032
rect 4022 2036 4028 2037
rect 4022 2032 4023 2036
rect 4027 2032 4028 2036
rect 4022 2031 4028 2032
rect 4158 2036 4164 2037
rect 4158 2032 4159 2036
rect 4163 2032 4164 2036
rect 4158 2031 4164 2032
rect 4294 2036 4300 2037
rect 4294 2032 4295 2036
rect 4299 2032 4300 2036
rect 4294 2031 4300 2032
rect 4430 2036 4436 2037
rect 4430 2032 4431 2036
rect 4435 2032 4436 2036
rect 4430 2031 4436 2032
rect 4566 2036 4572 2037
rect 4566 2032 4567 2036
rect 4571 2032 4572 2036
rect 4566 2031 4572 2032
rect 4718 2036 4724 2037
rect 4718 2032 4719 2036
rect 4723 2032 4724 2036
rect 4718 2031 4724 2032
rect 4894 2036 4900 2037
rect 4894 2032 4895 2036
rect 4899 2032 4900 2036
rect 4894 2031 4900 2032
rect 5086 2036 5092 2037
rect 5086 2032 5087 2036
rect 5091 2032 5092 2036
rect 5086 2031 5092 2032
rect 5278 2036 5284 2037
rect 5278 2032 5279 2036
rect 5283 2032 5284 2036
rect 5278 2031 5284 2032
rect 5478 2036 5484 2037
rect 5478 2032 5479 2036
rect 5483 2032 5484 2036
rect 5662 2033 5663 2037
rect 5667 2033 5668 2037
rect 5662 2032 5668 2033
rect 5478 2031 5484 2032
rect 110 2025 116 2026
rect 1934 2025 1940 2026
rect 110 2021 111 2025
rect 115 2021 116 2025
rect 110 2020 116 2021
rect 262 2024 268 2025
rect 262 2020 263 2024
rect 267 2020 268 2024
rect 262 2019 268 2020
rect 398 2024 404 2025
rect 398 2020 399 2024
rect 403 2020 404 2024
rect 398 2019 404 2020
rect 534 2024 540 2025
rect 534 2020 535 2024
rect 539 2020 540 2024
rect 534 2019 540 2020
rect 678 2024 684 2025
rect 678 2020 679 2024
rect 683 2020 684 2024
rect 678 2019 684 2020
rect 822 2024 828 2025
rect 822 2020 823 2024
rect 827 2020 828 2024
rect 822 2019 828 2020
rect 966 2024 972 2025
rect 966 2020 967 2024
rect 971 2020 972 2024
rect 966 2019 972 2020
rect 1110 2024 1116 2025
rect 1110 2020 1111 2024
rect 1115 2020 1116 2024
rect 1110 2019 1116 2020
rect 1254 2024 1260 2025
rect 1254 2020 1255 2024
rect 1259 2020 1260 2024
rect 1254 2019 1260 2020
rect 1398 2024 1404 2025
rect 1398 2020 1399 2024
rect 1403 2020 1404 2024
rect 1398 2019 1404 2020
rect 1542 2024 1548 2025
rect 1542 2020 1543 2024
rect 1547 2020 1548 2024
rect 1542 2019 1548 2020
rect 1678 2024 1684 2025
rect 1678 2020 1679 2024
rect 1683 2020 1684 2024
rect 1678 2019 1684 2020
rect 1814 2024 1820 2025
rect 1814 2020 1815 2024
rect 1819 2020 1820 2024
rect 1934 2021 1935 2025
rect 1939 2021 1940 2025
rect 3858 2021 3864 2022
rect 1934 2020 1940 2021
rect 3838 2020 3844 2021
rect 1814 2019 1820 2020
rect 3838 2016 3839 2020
rect 3843 2016 3844 2020
rect 3858 2017 3859 2021
rect 3863 2017 3864 2021
rect 3858 2016 3864 2017
rect 3994 2021 4000 2022
rect 3994 2017 3995 2021
rect 3999 2017 4000 2021
rect 3994 2016 4000 2017
rect 4130 2021 4136 2022
rect 4130 2017 4131 2021
rect 4135 2017 4136 2021
rect 4130 2016 4136 2017
rect 4266 2021 4272 2022
rect 4266 2017 4267 2021
rect 4271 2017 4272 2021
rect 4266 2016 4272 2017
rect 4402 2021 4408 2022
rect 4402 2017 4403 2021
rect 4407 2017 4408 2021
rect 4402 2016 4408 2017
rect 4538 2021 4544 2022
rect 4538 2017 4539 2021
rect 4543 2017 4544 2021
rect 4538 2016 4544 2017
rect 4690 2021 4696 2022
rect 4690 2017 4691 2021
rect 4695 2017 4696 2021
rect 4690 2016 4696 2017
rect 4866 2021 4872 2022
rect 4866 2017 4867 2021
rect 4871 2017 4872 2021
rect 4866 2016 4872 2017
rect 5058 2021 5064 2022
rect 5058 2017 5059 2021
rect 5063 2017 5064 2021
rect 5058 2016 5064 2017
rect 5250 2021 5256 2022
rect 5250 2017 5251 2021
rect 5255 2017 5256 2021
rect 5250 2016 5256 2017
rect 5450 2021 5456 2022
rect 5450 2017 5451 2021
rect 5455 2017 5456 2021
rect 5450 2016 5456 2017
rect 5662 2020 5668 2021
rect 5662 2016 5663 2020
rect 5667 2016 5668 2020
rect 3838 2015 3844 2016
rect 5662 2015 5668 2016
rect 3962 2011 3968 2012
rect 234 2009 240 2010
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 234 2005 235 2009
rect 239 2005 240 2009
rect 234 2004 240 2005
rect 370 2009 376 2010
rect 370 2005 371 2009
rect 375 2005 376 2009
rect 370 2004 376 2005
rect 506 2009 512 2010
rect 506 2005 507 2009
rect 511 2005 512 2009
rect 506 2004 512 2005
rect 650 2009 656 2010
rect 650 2005 651 2009
rect 655 2005 656 2009
rect 650 2004 656 2005
rect 794 2009 800 2010
rect 794 2005 795 2009
rect 799 2005 800 2009
rect 794 2004 800 2005
rect 938 2009 944 2010
rect 938 2005 939 2009
rect 943 2005 944 2009
rect 938 2004 944 2005
rect 1082 2009 1088 2010
rect 1082 2005 1083 2009
rect 1087 2005 1088 2009
rect 1082 2004 1088 2005
rect 1226 2009 1232 2010
rect 1226 2005 1227 2009
rect 1231 2005 1232 2009
rect 1226 2004 1232 2005
rect 1370 2009 1376 2010
rect 1370 2005 1371 2009
rect 1375 2005 1376 2009
rect 1370 2004 1376 2005
rect 1514 2009 1520 2010
rect 1514 2005 1515 2009
rect 1519 2005 1520 2009
rect 1514 2004 1520 2005
rect 1650 2009 1656 2010
rect 1650 2005 1651 2009
rect 1655 2005 1656 2009
rect 1650 2004 1656 2005
rect 1786 2009 1792 2010
rect 1786 2005 1787 2009
rect 1791 2005 1792 2009
rect 1786 2004 1792 2005
rect 1934 2008 1940 2009
rect 1934 2004 1935 2008
rect 1939 2004 1940 2008
rect 3962 2007 3963 2011
rect 3967 2010 3968 2011
rect 3983 2011 3989 2012
rect 3983 2010 3984 2011
rect 3967 2008 3984 2010
rect 3967 2007 3968 2008
rect 3962 2006 3968 2007
rect 3983 2007 3984 2008
rect 3988 2007 3989 2011
rect 3983 2006 3989 2007
rect 3991 2011 3997 2012
rect 3991 2007 3992 2011
rect 3996 2010 3997 2011
rect 4119 2011 4125 2012
rect 4119 2010 4120 2011
rect 3996 2008 4120 2010
rect 3996 2007 3997 2008
rect 3991 2006 3997 2007
rect 4119 2007 4120 2008
rect 4124 2007 4125 2011
rect 4119 2006 4125 2007
rect 4127 2011 4133 2012
rect 4127 2007 4128 2011
rect 4132 2010 4133 2011
rect 4255 2011 4261 2012
rect 4255 2010 4256 2011
rect 4132 2008 4256 2010
rect 4132 2007 4133 2008
rect 4127 2006 4133 2007
rect 4255 2007 4256 2008
rect 4260 2007 4261 2011
rect 4255 2006 4261 2007
rect 4263 2011 4269 2012
rect 4263 2007 4264 2011
rect 4268 2010 4269 2011
rect 4391 2011 4397 2012
rect 4391 2010 4392 2011
rect 4268 2008 4392 2010
rect 4268 2007 4269 2008
rect 4263 2006 4269 2007
rect 4391 2007 4392 2008
rect 4396 2007 4397 2011
rect 4391 2006 4397 2007
rect 4399 2011 4405 2012
rect 4399 2007 4400 2011
rect 4404 2010 4405 2011
rect 4527 2011 4533 2012
rect 4527 2010 4528 2011
rect 4404 2008 4528 2010
rect 4404 2007 4405 2008
rect 4399 2006 4405 2007
rect 4527 2007 4528 2008
rect 4532 2007 4533 2011
rect 4527 2006 4533 2007
rect 4535 2011 4541 2012
rect 4535 2007 4536 2011
rect 4540 2010 4541 2011
rect 4663 2011 4669 2012
rect 4663 2010 4664 2011
rect 4540 2008 4664 2010
rect 4540 2007 4541 2008
rect 4535 2006 4541 2007
rect 4663 2007 4664 2008
rect 4668 2007 4669 2011
rect 4663 2006 4669 2007
rect 4682 2011 4688 2012
rect 4682 2007 4683 2011
rect 4687 2010 4688 2011
rect 4815 2011 4821 2012
rect 4815 2010 4816 2011
rect 4687 2008 4816 2010
rect 4687 2007 4688 2008
rect 4682 2006 4688 2007
rect 4815 2007 4816 2008
rect 4820 2007 4821 2011
rect 4815 2006 4821 2007
rect 4834 2011 4840 2012
rect 4834 2007 4835 2011
rect 4839 2010 4840 2011
rect 4991 2011 4997 2012
rect 4991 2010 4992 2011
rect 4839 2008 4992 2010
rect 4839 2007 4840 2008
rect 4834 2006 4840 2007
rect 4991 2007 4992 2008
rect 4996 2007 4997 2011
rect 4991 2006 4997 2007
rect 5031 2011 5037 2012
rect 5031 2007 5032 2011
rect 5036 2010 5037 2011
rect 5183 2011 5189 2012
rect 5183 2010 5184 2011
rect 5036 2008 5184 2010
rect 5036 2007 5037 2008
rect 5031 2006 5037 2007
rect 5183 2007 5184 2008
rect 5188 2007 5189 2011
rect 5183 2006 5189 2007
rect 5223 2011 5229 2012
rect 5223 2007 5224 2011
rect 5228 2010 5229 2011
rect 5375 2011 5381 2012
rect 5375 2010 5376 2011
rect 5228 2008 5376 2010
rect 5228 2007 5229 2008
rect 5223 2006 5229 2007
rect 5375 2007 5376 2008
rect 5380 2007 5381 2011
rect 5375 2006 5381 2007
rect 5550 2011 5556 2012
rect 5550 2007 5551 2011
rect 5555 2010 5556 2011
rect 5575 2011 5581 2012
rect 5575 2010 5576 2011
rect 5555 2008 5576 2010
rect 5555 2007 5556 2008
rect 5550 2006 5556 2007
rect 5575 2007 5576 2008
rect 5580 2007 5581 2011
rect 5575 2006 5581 2007
rect 110 2003 116 2004
rect 1934 2003 1940 2004
rect 359 1999 365 2000
rect 359 1995 360 1999
rect 364 1998 365 1999
rect 386 1999 392 2000
rect 386 1998 387 1999
rect 364 1996 387 1998
rect 364 1995 365 1996
rect 359 1994 365 1995
rect 386 1995 387 1996
rect 391 1995 392 1999
rect 386 1994 392 1995
rect 495 1999 501 2000
rect 495 1995 496 1999
rect 500 1998 501 1999
rect 522 1999 528 2000
rect 522 1998 523 1999
rect 500 1996 523 1998
rect 500 1995 501 1996
rect 495 1994 501 1995
rect 522 1995 523 1996
rect 527 1995 528 1999
rect 522 1994 528 1995
rect 631 1999 637 2000
rect 631 1995 632 1999
rect 636 1998 637 1999
rect 666 1999 672 2000
rect 666 1998 667 1999
rect 636 1996 667 1998
rect 636 1995 637 1996
rect 631 1994 637 1995
rect 666 1995 667 1996
rect 671 1995 672 1999
rect 666 1994 672 1995
rect 775 1999 781 2000
rect 775 1995 776 1999
rect 780 1998 781 1999
rect 810 1999 816 2000
rect 810 1998 811 1999
rect 780 1996 811 1998
rect 780 1995 781 1996
rect 775 1994 781 1995
rect 810 1995 811 1996
rect 815 1995 816 1999
rect 810 1994 816 1995
rect 919 1999 925 2000
rect 919 1995 920 1999
rect 924 1998 925 1999
rect 954 1999 960 2000
rect 954 1998 955 1999
rect 924 1996 955 1998
rect 924 1995 925 1996
rect 919 1994 925 1995
rect 954 1995 955 1996
rect 959 1995 960 1999
rect 954 1994 960 1995
rect 1002 1999 1008 2000
rect 1002 1995 1003 1999
rect 1007 1998 1008 1999
rect 1063 1999 1069 2000
rect 1063 1998 1064 1999
rect 1007 1996 1064 1998
rect 1007 1995 1008 1996
rect 1002 1994 1008 1995
rect 1063 1995 1064 1996
rect 1068 1995 1069 1999
rect 1207 1999 1213 2000
rect 1207 1998 1208 1999
rect 1063 1994 1069 1995
rect 1100 1996 1208 1998
rect 930 1991 936 1992
rect 930 1987 931 1991
rect 935 1990 936 1991
rect 1100 1990 1102 1996
rect 1207 1995 1208 1996
rect 1212 1995 1213 1999
rect 1207 1994 1213 1995
rect 1215 1999 1221 2000
rect 1215 1995 1216 1999
rect 1220 1998 1221 1999
rect 1351 1999 1357 2000
rect 1351 1998 1352 1999
rect 1220 1996 1352 1998
rect 1220 1995 1221 1996
rect 1215 1994 1221 1995
rect 1351 1995 1352 1996
rect 1356 1995 1357 1999
rect 1351 1994 1357 1995
rect 1359 1999 1365 2000
rect 1359 1995 1360 1999
rect 1364 1998 1365 1999
rect 1495 1999 1501 2000
rect 1495 1998 1496 1999
rect 1364 1996 1496 1998
rect 1364 1995 1365 1996
rect 1359 1994 1365 1995
rect 1495 1995 1496 1996
rect 1500 1995 1501 1999
rect 1495 1994 1501 1995
rect 1626 1999 1632 2000
rect 1626 1995 1627 1999
rect 1631 1998 1632 1999
rect 1639 1999 1645 2000
rect 1639 1998 1640 1999
rect 1631 1996 1640 1998
rect 1631 1995 1632 1996
rect 1626 1994 1632 1995
rect 1639 1995 1640 1996
rect 1644 1995 1645 1999
rect 1639 1994 1645 1995
rect 1775 1999 1781 2000
rect 1775 1995 1776 1999
rect 1780 1998 1781 1999
rect 1802 1999 1808 2000
rect 1802 1998 1803 1999
rect 1780 1996 1803 1998
rect 1780 1995 1781 1996
rect 1775 1994 1781 1995
rect 1802 1995 1803 1996
rect 1807 1995 1808 1999
rect 1802 1994 1808 1995
rect 1911 1999 1917 2000
rect 1911 1995 1912 1999
rect 1916 1995 1917 1999
rect 1911 1994 1917 1995
rect 935 1988 1102 1990
rect 1602 1991 1608 1992
rect 935 1987 936 1988
rect 930 1986 936 1987
rect 1602 1987 1603 1991
rect 1607 1990 1608 1991
rect 1913 1990 1915 1994
rect 1607 1988 1915 1990
rect 1607 1987 1608 1988
rect 1602 1986 1608 1987
rect 3991 1979 3997 1980
rect 3991 1978 3992 1979
rect 3949 1976 3992 1978
rect 3991 1975 3992 1976
rect 3996 1975 3997 1979
rect 4127 1979 4133 1980
rect 4127 1978 4128 1979
rect 4085 1976 4128 1978
rect 3991 1974 3997 1975
rect 4127 1975 4128 1976
rect 4132 1975 4133 1979
rect 4263 1979 4269 1980
rect 4263 1978 4264 1979
rect 4221 1976 4264 1978
rect 4127 1974 4133 1975
rect 4263 1975 4264 1976
rect 4268 1975 4269 1979
rect 4399 1979 4405 1980
rect 4399 1978 4400 1979
rect 4357 1976 4400 1978
rect 4263 1974 4269 1975
rect 4399 1975 4400 1976
rect 4404 1975 4405 1979
rect 4399 1974 4405 1975
rect 4490 1979 4496 1980
rect 4490 1975 4491 1979
rect 4495 1975 4496 1979
rect 4682 1979 4688 1980
rect 4682 1978 4683 1979
rect 4629 1976 4683 1978
rect 4490 1974 4496 1975
rect 4682 1975 4683 1976
rect 4687 1975 4688 1979
rect 4834 1979 4840 1980
rect 4834 1978 4835 1979
rect 4781 1976 4835 1978
rect 4682 1974 4688 1975
rect 4834 1975 4835 1976
rect 4839 1975 4840 1979
rect 5031 1979 5037 1980
rect 5031 1978 5032 1979
rect 4957 1976 5032 1978
rect 4834 1974 4840 1975
rect 5031 1975 5032 1976
rect 5036 1975 5037 1979
rect 5223 1979 5229 1980
rect 5223 1978 5224 1979
rect 5149 1976 5224 1978
rect 5031 1974 5037 1975
rect 5223 1975 5224 1976
rect 5228 1975 5229 1979
rect 5354 1979 5360 1980
rect 5354 1978 5355 1979
rect 5341 1976 5355 1978
rect 5223 1974 5229 1975
rect 5354 1975 5355 1976
rect 5359 1975 5360 1979
rect 5354 1974 5360 1975
rect 5502 1979 5508 1980
rect 5502 1975 5503 1979
rect 5507 1975 5508 1979
rect 5502 1974 5508 1975
rect 386 1967 392 1968
rect 325 1964 374 1966
rect 372 1950 374 1964
rect 386 1963 387 1967
rect 391 1963 392 1967
rect 386 1962 392 1963
rect 522 1967 528 1968
rect 522 1963 523 1967
rect 527 1963 528 1967
rect 522 1962 528 1963
rect 666 1967 672 1968
rect 666 1963 667 1967
rect 671 1963 672 1967
rect 666 1962 672 1963
rect 810 1967 816 1968
rect 810 1963 811 1967
rect 815 1963 816 1967
rect 810 1962 816 1963
rect 954 1967 960 1968
rect 954 1963 955 1967
rect 959 1963 960 1967
rect 1215 1967 1221 1968
rect 1215 1966 1216 1967
rect 1173 1964 1216 1966
rect 954 1962 960 1963
rect 1215 1963 1216 1964
rect 1220 1963 1221 1967
rect 1359 1967 1365 1968
rect 1359 1966 1360 1967
rect 1317 1964 1360 1966
rect 1215 1962 1221 1963
rect 1359 1963 1360 1964
rect 1364 1963 1365 1967
rect 1359 1962 1365 1963
rect 1458 1967 1464 1968
rect 1458 1963 1459 1967
rect 1463 1963 1464 1967
rect 1458 1962 1464 1963
rect 1602 1967 1608 1968
rect 1602 1963 1603 1967
rect 1607 1963 1608 1967
rect 1602 1962 1608 1963
rect 1738 1967 1744 1968
rect 1738 1963 1739 1967
rect 1743 1963 1744 1967
rect 1738 1962 1744 1963
rect 1802 1967 1808 1968
rect 1802 1963 1803 1967
rect 1807 1963 1808 1967
rect 1802 1962 1808 1963
rect 750 1951 756 1952
rect 750 1950 751 1951
rect 372 1948 751 1950
rect 750 1947 751 1948
rect 755 1947 756 1951
rect 750 1946 756 1947
rect 4535 1943 4541 1944
rect 4535 1942 4536 1943
rect 4164 1940 4536 1942
rect 3962 1931 3968 1932
rect 3962 1930 3963 1931
rect 3949 1928 3963 1930
rect 3962 1927 3963 1928
rect 3967 1927 3968 1931
rect 4164 1930 4166 1940
rect 4535 1939 4536 1940
rect 4540 1939 4541 1943
rect 4535 1938 4541 1939
rect 4666 1943 4672 1944
rect 4666 1939 4667 1943
rect 4671 1942 4672 1943
rect 5326 1943 5332 1944
rect 5326 1942 5327 1943
rect 4671 1940 5327 1942
rect 4671 1939 4672 1940
rect 4666 1938 4672 1939
rect 5326 1939 5327 1940
rect 5331 1939 5332 1943
rect 5326 1938 5332 1939
rect 4133 1928 4166 1930
rect 4170 1931 4176 1932
rect 3962 1926 3968 1927
rect 4170 1927 4171 1931
rect 4175 1930 4176 1931
rect 4410 1931 4416 1932
rect 4175 1928 4301 1930
rect 4175 1927 4176 1928
rect 4170 1926 4176 1927
rect 4410 1927 4411 1931
rect 4415 1930 4416 1931
rect 4690 1931 4696 1932
rect 4415 1928 4581 1930
rect 4415 1927 4416 1928
rect 4410 1926 4416 1927
rect 4690 1927 4691 1931
rect 4695 1930 4696 1931
rect 5002 1931 5008 1932
rect 4695 1928 4893 1930
rect 4695 1927 4696 1928
rect 4690 1926 4696 1927
rect 5002 1927 5003 1931
rect 5007 1930 5008 1931
rect 5618 1931 5624 1932
rect 5618 1930 5619 1931
rect 5007 1928 5221 1930
rect 5605 1928 5619 1930
rect 5007 1927 5008 1928
rect 5002 1926 5008 1927
rect 5618 1927 5619 1928
rect 5623 1927 5624 1931
rect 5618 1926 5624 1927
rect 362 1907 368 1908
rect 322 1903 328 1904
rect 322 1899 323 1903
rect 327 1899 328 1903
rect 362 1903 363 1907
rect 367 1906 368 1907
rect 562 1907 568 1908
rect 367 1904 453 1906
rect 367 1903 368 1904
rect 362 1902 368 1903
rect 562 1903 563 1907
rect 567 1906 568 1907
rect 930 1907 936 1908
rect 930 1906 931 1907
rect 567 1904 645 1906
rect 901 1904 931 1906
rect 567 1903 568 1904
rect 562 1902 568 1903
rect 930 1903 931 1904
rect 935 1903 936 1907
rect 930 1902 936 1903
rect 938 1907 944 1908
rect 938 1903 939 1907
rect 943 1906 944 1907
rect 1114 1907 1120 1908
rect 943 1904 1005 1906
rect 943 1903 944 1904
rect 938 1902 944 1903
rect 1114 1903 1115 1907
rect 1119 1906 1120 1907
rect 1450 1907 1456 1908
rect 1119 1904 1173 1906
rect 1119 1903 1120 1904
rect 1114 1902 1120 1903
rect 1410 1903 1416 1904
rect 322 1898 328 1899
rect 1410 1899 1411 1903
rect 1415 1899 1416 1903
rect 1450 1903 1451 1907
rect 1455 1906 1456 1907
rect 1610 1907 1616 1908
rect 1455 1904 1501 1906
rect 1455 1903 1456 1904
rect 1450 1902 1456 1903
rect 1610 1903 1611 1907
rect 1615 1906 1616 1907
rect 2002 1907 2008 1908
rect 2002 1906 2003 1907
rect 1615 1904 1661 1906
rect 1877 1904 2003 1906
rect 1615 1903 1616 1904
rect 1610 1902 1616 1903
rect 2002 1903 2003 1904
rect 2007 1903 2008 1907
rect 2002 1902 2008 1903
rect 1410 1898 1416 1899
rect 1974 1901 1980 1902
rect 3798 1901 3804 1902
rect 1974 1897 1975 1901
rect 1979 1897 1980 1901
rect 1974 1896 1980 1897
rect 3134 1900 3140 1901
rect 3134 1896 3135 1900
rect 3139 1896 3140 1900
rect 3134 1895 3140 1896
rect 3270 1900 3276 1901
rect 3270 1896 3271 1900
rect 3275 1896 3276 1900
rect 3270 1895 3276 1896
rect 3406 1900 3412 1901
rect 3406 1896 3407 1900
rect 3411 1896 3412 1900
rect 3406 1895 3412 1896
rect 3542 1900 3548 1901
rect 3542 1896 3543 1900
rect 3547 1896 3548 1900
rect 3542 1895 3548 1896
rect 3678 1900 3684 1901
rect 3678 1896 3679 1900
rect 3683 1896 3684 1900
rect 3798 1897 3799 1901
rect 3803 1897 3804 1901
rect 3798 1896 3804 1897
rect 3678 1895 3684 1896
rect 3822 1895 3828 1896
rect 3822 1891 3823 1895
rect 3827 1894 3828 1895
rect 3983 1895 3989 1896
rect 3983 1894 3984 1895
rect 3827 1892 3984 1894
rect 3827 1891 3828 1892
rect 3822 1890 3828 1891
rect 3983 1891 3984 1892
rect 3988 1891 3989 1895
rect 3983 1890 3989 1891
rect 4167 1895 4176 1896
rect 4167 1891 4168 1895
rect 4175 1891 4176 1895
rect 4167 1890 4176 1891
rect 4407 1895 4416 1896
rect 4407 1891 4408 1895
rect 4415 1891 4416 1895
rect 4407 1890 4416 1891
rect 4466 1895 4472 1896
rect 4466 1891 4467 1895
rect 4471 1894 4472 1895
rect 4666 1895 4672 1896
rect 4666 1894 4667 1895
rect 4471 1892 4667 1894
rect 4471 1891 4472 1892
rect 4466 1890 4472 1891
rect 4666 1891 4667 1892
rect 4671 1891 4672 1895
rect 4666 1890 4672 1891
rect 4687 1895 4696 1896
rect 4687 1891 4688 1895
rect 4695 1891 4696 1895
rect 4687 1890 4696 1891
rect 4999 1895 5008 1896
rect 4999 1891 5000 1895
rect 5007 1891 5008 1895
rect 4999 1890 5008 1891
rect 5326 1895 5333 1896
rect 5326 1891 5327 1895
rect 5332 1891 5333 1895
rect 5326 1890 5333 1891
rect 5618 1895 5624 1896
rect 5618 1891 5619 1895
rect 5623 1894 5624 1895
rect 5639 1895 5645 1896
rect 5639 1894 5640 1895
rect 5623 1892 5640 1894
rect 5623 1891 5624 1892
rect 5618 1890 5624 1891
rect 5639 1891 5640 1892
rect 5644 1891 5645 1895
rect 5639 1890 5645 1891
rect 3838 1888 3844 1889
rect 5662 1888 5668 1889
rect 3106 1885 3112 1886
rect 1974 1884 1980 1885
rect 1974 1880 1975 1884
rect 1979 1880 1980 1884
rect 3106 1881 3107 1885
rect 3111 1881 3112 1885
rect 3106 1880 3112 1881
rect 3242 1885 3248 1886
rect 3242 1881 3243 1885
rect 3247 1881 3248 1885
rect 3242 1880 3248 1881
rect 3378 1885 3384 1886
rect 3378 1881 3379 1885
rect 3383 1881 3384 1885
rect 3378 1880 3384 1881
rect 3514 1885 3520 1886
rect 3514 1881 3515 1885
rect 3519 1881 3520 1885
rect 3514 1880 3520 1881
rect 3650 1885 3656 1886
rect 3650 1881 3651 1885
rect 3655 1881 3656 1885
rect 3650 1880 3656 1881
rect 3798 1884 3804 1885
rect 3798 1880 3799 1884
rect 3803 1880 3804 1884
rect 3838 1884 3839 1888
rect 3843 1884 3844 1888
rect 3838 1883 3844 1884
rect 3858 1887 3864 1888
rect 3858 1883 3859 1887
rect 3863 1883 3864 1887
rect 3858 1882 3864 1883
rect 4042 1887 4048 1888
rect 4042 1883 4043 1887
rect 4047 1883 4048 1887
rect 4042 1882 4048 1883
rect 4282 1887 4288 1888
rect 4282 1883 4283 1887
rect 4287 1883 4288 1887
rect 4282 1882 4288 1883
rect 4562 1887 4568 1888
rect 4562 1883 4563 1887
rect 4567 1883 4568 1887
rect 4562 1882 4568 1883
rect 4874 1887 4880 1888
rect 4874 1883 4875 1887
rect 4879 1883 4880 1887
rect 4874 1882 4880 1883
rect 5202 1887 5208 1888
rect 5202 1883 5203 1887
rect 5207 1883 5208 1887
rect 5202 1882 5208 1883
rect 5514 1887 5520 1888
rect 5514 1883 5515 1887
rect 5519 1883 5520 1887
rect 5662 1884 5663 1888
rect 5667 1884 5668 1888
rect 5662 1883 5668 1884
rect 5514 1882 5520 1883
rect 1410 1879 1416 1880
rect 1974 1879 1980 1880
rect 3798 1879 3804 1880
rect 1410 1875 1411 1879
rect 1415 1878 1416 1879
rect 1415 1876 1915 1878
rect 1415 1875 1416 1876
rect 1410 1874 1416 1875
rect 1913 1872 1915 1876
rect 3231 1875 3237 1876
rect 359 1871 368 1872
rect 359 1867 360 1871
rect 367 1867 368 1871
rect 359 1866 368 1867
rect 559 1871 568 1872
rect 559 1867 560 1871
rect 567 1867 568 1871
rect 559 1866 568 1867
rect 750 1871 757 1872
rect 750 1867 751 1871
rect 756 1867 757 1871
rect 750 1866 757 1867
rect 935 1871 944 1872
rect 935 1867 936 1871
rect 943 1867 944 1871
rect 935 1866 944 1867
rect 1111 1871 1120 1872
rect 1111 1867 1112 1871
rect 1119 1867 1120 1871
rect 1111 1866 1120 1867
rect 1279 1871 1285 1872
rect 1279 1867 1280 1871
rect 1284 1870 1285 1871
rect 1378 1871 1384 1872
rect 1378 1870 1379 1871
rect 1284 1868 1379 1870
rect 1284 1867 1285 1868
rect 1279 1866 1285 1867
rect 1378 1867 1379 1868
rect 1383 1867 1384 1871
rect 1378 1866 1384 1867
rect 1447 1871 1456 1872
rect 1447 1867 1448 1871
rect 1455 1867 1456 1871
rect 1447 1866 1456 1867
rect 1607 1871 1616 1872
rect 1607 1867 1608 1871
rect 1615 1867 1616 1871
rect 1607 1866 1616 1867
rect 1738 1871 1744 1872
rect 1738 1867 1739 1871
rect 1743 1870 1744 1871
rect 1767 1871 1773 1872
rect 1767 1870 1768 1871
rect 1743 1868 1768 1870
rect 1743 1867 1744 1868
rect 1738 1866 1744 1867
rect 1767 1867 1768 1868
rect 1772 1867 1773 1871
rect 1767 1866 1773 1867
rect 1911 1871 1917 1872
rect 1911 1867 1912 1871
rect 1916 1867 1917 1871
rect 3231 1871 3232 1875
rect 3236 1874 3237 1875
rect 3258 1875 3264 1876
rect 3258 1874 3259 1875
rect 3236 1872 3259 1874
rect 3236 1871 3237 1872
rect 3231 1870 3237 1871
rect 3258 1871 3259 1872
rect 3263 1871 3264 1875
rect 3258 1870 3264 1871
rect 3346 1875 3352 1876
rect 3346 1871 3347 1875
rect 3351 1874 3352 1875
rect 3367 1875 3373 1876
rect 3367 1874 3368 1875
rect 3351 1872 3368 1874
rect 3351 1871 3352 1872
rect 3346 1870 3352 1871
rect 3367 1871 3368 1872
rect 3372 1871 3373 1875
rect 3503 1875 3509 1876
rect 3503 1874 3504 1875
rect 3367 1870 3373 1871
rect 3376 1872 3504 1874
rect 1911 1866 1917 1867
rect 3194 1867 3200 1868
rect 110 1864 116 1865
rect 1934 1864 1940 1865
rect 110 1860 111 1864
rect 115 1860 116 1864
rect 110 1859 116 1860
rect 234 1863 240 1864
rect 234 1859 235 1863
rect 239 1859 240 1863
rect 234 1858 240 1859
rect 434 1863 440 1864
rect 434 1859 435 1863
rect 439 1859 440 1863
rect 434 1858 440 1859
rect 626 1863 632 1864
rect 626 1859 627 1863
rect 631 1859 632 1863
rect 626 1858 632 1859
rect 810 1863 816 1864
rect 810 1859 811 1863
rect 815 1859 816 1863
rect 810 1858 816 1859
rect 986 1863 992 1864
rect 986 1859 987 1863
rect 991 1859 992 1863
rect 986 1858 992 1859
rect 1154 1863 1160 1864
rect 1154 1859 1155 1863
rect 1159 1859 1160 1863
rect 1154 1858 1160 1859
rect 1322 1863 1328 1864
rect 1322 1859 1323 1863
rect 1327 1859 1328 1863
rect 1322 1858 1328 1859
rect 1482 1863 1488 1864
rect 1482 1859 1483 1863
rect 1487 1859 1488 1863
rect 1482 1858 1488 1859
rect 1642 1863 1648 1864
rect 1642 1859 1643 1863
rect 1647 1859 1648 1863
rect 1642 1858 1648 1859
rect 1786 1863 1792 1864
rect 1786 1859 1787 1863
rect 1791 1859 1792 1863
rect 1934 1860 1935 1864
rect 1939 1860 1940 1864
rect 3194 1863 3195 1867
rect 3199 1866 3200 1867
rect 3376 1866 3378 1872
rect 3503 1871 3504 1872
rect 3508 1871 3509 1875
rect 3503 1870 3509 1871
rect 3511 1875 3517 1876
rect 3511 1871 3512 1875
rect 3516 1874 3517 1875
rect 3639 1875 3645 1876
rect 3639 1874 3640 1875
rect 3516 1872 3640 1874
rect 3516 1871 3517 1872
rect 3511 1870 3517 1871
rect 3639 1871 3640 1872
rect 3644 1871 3645 1875
rect 3639 1870 3645 1871
rect 3647 1875 3653 1876
rect 3647 1871 3648 1875
rect 3652 1874 3653 1875
rect 3775 1875 3781 1876
rect 3775 1874 3776 1875
rect 3652 1872 3776 1874
rect 3652 1871 3653 1872
rect 3647 1870 3653 1871
rect 3775 1871 3776 1872
rect 3780 1871 3781 1875
rect 3886 1872 3892 1873
rect 3775 1870 3781 1871
rect 3838 1871 3844 1872
rect 3838 1867 3839 1871
rect 3843 1867 3844 1871
rect 3886 1868 3887 1872
rect 3891 1868 3892 1872
rect 3886 1867 3892 1868
rect 4070 1872 4076 1873
rect 4070 1868 4071 1872
rect 4075 1868 4076 1872
rect 4070 1867 4076 1868
rect 4310 1872 4316 1873
rect 4310 1868 4311 1872
rect 4315 1868 4316 1872
rect 4310 1867 4316 1868
rect 4590 1872 4596 1873
rect 4590 1868 4591 1872
rect 4595 1868 4596 1872
rect 4590 1867 4596 1868
rect 4902 1872 4908 1873
rect 4902 1868 4903 1872
rect 4907 1868 4908 1872
rect 4902 1867 4908 1868
rect 5230 1872 5236 1873
rect 5230 1868 5231 1872
rect 5235 1868 5236 1872
rect 5230 1867 5236 1868
rect 5542 1872 5548 1873
rect 5542 1868 5543 1872
rect 5547 1868 5548 1872
rect 5542 1867 5548 1868
rect 5662 1871 5668 1872
rect 5662 1867 5663 1871
rect 5667 1867 5668 1871
rect 3838 1866 3844 1867
rect 5662 1866 5668 1867
rect 3199 1864 3378 1866
rect 3199 1863 3200 1864
rect 3194 1862 3200 1863
rect 1934 1859 1940 1860
rect 1786 1858 1792 1859
rect 262 1848 268 1849
rect 110 1847 116 1848
rect 110 1843 111 1847
rect 115 1843 116 1847
rect 262 1844 263 1848
rect 267 1844 268 1848
rect 262 1843 268 1844
rect 462 1848 468 1849
rect 462 1844 463 1848
rect 467 1844 468 1848
rect 462 1843 468 1844
rect 654 1848 660 1849
rect 654 1844 655 1848
rect 659 1844 660 1848
rect 654 1843 660 1844
rect 838 1848 844 1849
rect 838 1844 839 1848
rect 843 1844 844 1848
rect 838 1843 844 1844
rect 1014 1848 1020 1849
rect 1014 1844 1015 1848
rect 1019 1844 1020 1848
rect 1014 1843 1020 1844
rect 1182 1848 1188 1849
rect 1182 1844 1183 1848
rect 1187 1844 1188 1848
rect 1182 1843 1188 1844
rect 1350 1848 1356 1849
rect 1350 1844 1351 1848
rect 1355 1844 1356 1848
rect 1350 1843 1356 1844
rect 1510 1848 1516 1849
rect 1510 1844 1511 1848
rect 1515 1844 1516 1848
rect 1510 1843 1516 1844
rect 1670 1848 1676 1849
rect 1670 1844 1671 1848
rect 1675 1844 1676 1848
rect 1670 1843 1676 1844
rect 1814 1848 1820 1849
rect 1814 1844 1815 1848
rect 1819 1844 1820 1848
rect 1814 1843 1820 1844
rect 1934 1847 1940 1848
rect 1934 1843 1935 1847
rect 1939 1843 1940 1847
rect 110 1842 116 1843
rect 1934 1842 1940 1843
rect 3194 1843 3200 1844
rect 3194 1839 3195 1843
rect 3199 1839 3200 1843
rect 3194 1838 3200 1839
rect 3258 1843 3264 1844
rect 3258 1839 3259 1843
rect 3263 1839 3264 1843
rect 3511 1843 3517 1844
rect 3511 1842 3512 1843
rect 3469 1840 3512 1842
rect 3258 1838 3264 1839
rect 3511 1839 3512 1840
rect 3516 1839 3517 1843
rect 3647 1843 3653 1844
rect 3647 1842 3648 1843
rect 3605 1840 3648 1842
rect 3511 1838 3517 1839
rect 3647 1839 3648 1840
rect 3652 1839 3653 1843
rect 3822 1843 3828 1844
rect 3822 1842 3823 1843
rect 3741 1840 3823 1842
rect 3647 1838 3653 1839
rect 3822 1839 3823 1840
rect 3827 1839 3828 1843
rect 3822 1838 3828 1839
rect 3838 1813 3844 1814
rect 5662 1813 5668 1814
rect 3838 1809 3839 1813
rect 3843 1809 3844 1813
rect 3838 1808 3844 1809
rect 4406 1812 4412 1813
rect 4406 1808 4407 1812
rect 4411 1808 4412 1812
rect 4406 1807 4412 1808
rect 4542 1812 4548 1813
rect 4542 1808 4543 1812
rect 4547 1808 4548 1812
rect 4542 1807 4548 1808
rect 4678 1812 4684 1813
rect 4678 1808 4679 1812
rect 4683 1808 4684 1812
rect 4678 1807 4684 1808
rect 4814 1812 4820 1813
rect 4814 1808 4815 1812
rect 4819 1808 4820 1812
rect 4814 1807 4820 1808
rect 4950 1812 4956 1813
rect 4950 1808 4951 1812
rect 4955 1808 4956 1812
rect 5662 1809 5663 1813
rect 5667 1809 5668 1813
rect 5662 1808 5668 1809
rect 4950 1807 4956 1808
rect 4378 1797 4384 1798
rect 3838 1796 3844 1797
rect 3838 1792 3839 1796
rect 3843 1792 3844 1796
rect 4378 1793 4379 1797
rect 4383 1793 4384 1797
rect 4378 1792 4384 1793
rect 4514 1797 4520 1798
rect 4514 1793 4515 1797
rect 4519 1793 4520 1797
rect 4514 1792 4520 1793
rect 4650 1797 4656 1798
rect 4650 1793 4651 1797
rect 4655 1793 4656 1797
rect 4650 1792 4656 1793
rect 4786 1797 4792 1798
rect 4786 1793 4787 1797
rect 4791 1793 4792 1797
rect 4786 1792 4792 1793
rect 4922 1797 4928 1798
rect 4922 1793 4923 1797
rect 4927 1793 4928 1797
rect 4922 1792 4928 1793
rect 5662 1796 5668 1797
rect 5662 1792 5663 1796
rect 5667 1792 5668 1796
rect 3838 1791 3844 1792
rect 5662 1791 5668 1792
rect 4503 1787 4509 1788
rect 2127 1783 2133 1784
rect 2127 1782 2128 1783
rect 2085 1780 2128 1782
rect 2127 1779 2128 1780
rect 2132 1779 2133 1783
rect 2263 1783 2269 1784
rect 2263 1782 2264 1783
rect 2221 1780 2264 1782
rect 2127 1778 2133 1779
rect 2263 1779 2264 1780
rect 2268 1779 2269 1783
rect 2415 1783 2421 1784
rect 2415 1782 2416 1783
rect 2357 1780 2416 1782
rect 2263 1778 2269 1779
rect 2415 1779 2416 1780
rect 2420 1779 2421 1783
rect 2567 1783 2573 1784
rect 2567 1782 2568 1783
rect 2509 1780 2568 1782
rect 2415 1778 2421 1779
rect 2567 1779 2568 1780
rect 2572 1779 2573 1783
rect 2722 1783 2728 1784
rect 2722 1782 2723 1783
rect 2669 1780 2723 1782
rect 2567 1778 2573 1779
rect 2722 1779 2723 1780
rect 2727 1779 2728 1783
rect 2722 1778 2728 1779
rect 2730 1783 2736 1784
rect 2730 1779 2731 1783
rect 2735 1782 2736 1783
rect 3022 1783 3028 1784
rect 3022 1782 3023 1783
rect 2735 1780 2757 1782
rect 2989 1780 3023 1782
rect 2735 1779 2736 1780
rect 2730 1778 2736 1779
rect 3022 1779 3023 1780
rect 3027 1779 3028 1783
rect 3022 1778 3028 1779
rect 3031 1783 3037 1784
rect 3031 1779 3032 1783
rect 3036 1782 3037 1783
rect 3178 1783 3184 1784
rect 3036 1780 3069 1782
rect 3036 1779 3037 1780
rect 3031 1778 3037 1779
rect 3178 1779 3179 1783
rect 3183 1782 3184 1783
rect 3346 1783 3352 1784
rect 3183 1780 3221 1782
rect 3183 1779 3184 1780
rect 3178 1778 3184 1779
rect 3346 1779 3347 1783
rect 3351 1782 3352 1783
rect 3482 1783 3488 1784
rect 3351 1780 3373 1782
rect 3351 1779 3352 1780
rect 3346 1778 3352 1779
rect 3482 1779 3483 1783
rect 3487 1782 3488 1783
rect 3647 1783 3653 1784
rect 3487 1780 3533 1782
rect 3487 1779 3488 1780
rect 3482 1778 3488 1779
rect 3647 1779 3648 1783
rect 3652 1782 3653 1783
rect 4503 1783 4504 1787
rect 4508 1786 4509 1787
rect 4530 1787 4536 1788
rect 4530 1786 4531 1787
rect 4508 1784 4531 1786
rect 4508 1783 4509 1784
rect 4503 1782 4509 1783
rect 4530 1783 4531 1784
rect 4535 1783 4536 1787
rect 4530 1782 4536 1783
rect 4639 1787 4645 1788
rect 4639 1783 4640 1787
rect 4644 1786 4645 1787
rect 4666 1787 4672 1788
rect 4666 1786 4667 1787
rect 4644 1784 4667 1786
rect 4644 1783 4645 1784
rect 4639 1782 4645 1783
rect 4666 1783 4667 1784
rect 4671 1783 4672 1787
rect 4666 1782 4672 1783
rect 4775 1787 4781 1788
rect 4775 1783 4776 1787
rect 4780 1786 4781 1787
rect 4802 1787 4808 1788
rect 4802 1786 4803 1787
rect 4780 1784 4803 1786
rect 4780 1783 4781 1784
rect 4775 1782 4781 1783
rect 4802 1783 4803 1784
rect 4807 1783 4808 1787
rect 4802 1782 4808 1783
rect 4911 1787 4917 1788
rect 4911 1783 4912 1787
rect 4916 1786 4917 1787
rect 4938 1787 4944 1788
rect 4938 1786 4939 1787
rect 4916 1784 4939 1786
rect 4916 1783 4917 1784
rect 4911 1782 4917 1783
rect 4938 1783 4939 1784
rect 4943 1783 4944 1787
rect 4938 1782 4944 1783
rect 4950 1787 4956 1788
rect 4950 1783 4951 1787
rect 4955 1786 4956 1787
rect 5047 1787 5053 1788
rect 5047 1786 5048 1787
rect 4955 1784 5048 1786
rect 4955 1783 4956 1784
rect 4950 1782 4956 1783
rect 5047 1783 5048 1784
rect 5052 1783 5053 1787
rect 5047 1782 5053 1783
rect 3652 1780 3669 1782
rect 3652 1779 3653 1780
rect 3647 1778 3653 1779
rect 110 1777 116 1778
rect 1934 1777 1940 1778
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 110 1772 116 1773
rect 222 1776 228 1777
rect 222 1772 223 1776
rect 227 1772 228 1776
rect 222 1771 228 1772
rect 462 1776 468 1777
rect 462 1772 463 1776
rect 467 1772 468 1776
rect 462 1771 468 1772
rect 694 1776 700 1777
rect 694 1772 695 1776
rect 699 1772 700 1776
rect 694 1771 700 1772
rect 926 1776 932 1777
rect 926 1772 927 1776
rect 931 1772 932 1776
rect 926 1771 932 1772
rect 1158 1776 1164 1777
rect 1158 1772 1159 1776
rect 1163 1772 1164 1776
rect 1158 1771 1164 1772
rect 1390 1776 1396 1777
rect 1390 1772 1391 1776
rect 1395 1772 1396 1776
rect 1934 1773 1935 1777
rect 1939 1773 1940 1777
rect 1934 1772 1940 1773
rect 1390 1771 1396 1772
rect 194 1761 200 1762
rect 110 1760 116 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 194 1757 195 1761
rect 199 1757 200 1761
rect 194 1756 200 1757
rect 434 1761 440 1762
rect 434 1757 435 1761
rect 439 1757 440 1761
rect 434 1756 440 1757
rect 666 1761 672 1762
rect 666 1757 667 1761
rect 671 1757 672 1761
rect 666 1756 672 1757
rect 898 1761 904 1762
rect 898 1757 899 1761
rect 903 1757 904 1761
rect 898 1756 904 1757
rect 1130 1761 1136 1762
rect 1130 1757 1131 1761
rect 1135 1757 1136 1761
rect 1130 1756 1136 1757
rect 1362 1761 1368 1762
rect 1362 1757 1363 1761
rect 1367 1757 1368 1761
rect 1362 1756 1368 1757
rect 1934 1760 1940 1761
rect 1934 1756 1935 1760
rect 1939 1756 1940 1760
rect 110 1755 116 1756
rect 1934 1755 1940 1756
rect 4466 1755 4472 1756
rect 319 1751 328 1752
rect 319 1747 320 1751
rect 327 1747 328 1751
rect 319 1746 328 1747
rect 383 1751 389 1752
rect 383 1747 384 1751
rect 388 1750 389 1751
rect 559 1751 565 1752
rect 559 1750 560 1751
rect 388 1748 560 1750
rect 388 1747 389 1748
rect 383 1746 389 1747
rect 559 1747 560 1748
rect 564 1747 565 1751
rect 559 1746 565 1747
rect 791 1751 797 1752
rect 791 1747 792 1751
rect 796 1750 797 1751
rect 914 1751 920 1752
rect 914 1750 915 1751
rect 796 1748 915 1750
rect 796 1747 797 1748
rect 791 1746 797 1747
rect 914 1747 915 1748
rect 919 1747 920 1751
rect 914 1746 920 1747
rect 1023 1751 1029 1752
rect 1023 1747 1024 1751
rect 1028 1750 1029 1751
rect 1146 1751 1152 1752
rect 1146 1750 1147 1751
rect 1028 1748 1147 1750
rect 1028 1747 1029 1748
rect 1023 1746 1029 1747
rect 1146 1747 1147 1748
rect 1151 1747 1152 1751
rect 1146 1746 1152 1747
rect 1242 1751 1248 1752
rect 1242 1747 1243 1751
rect 1247 1750 1248 1751
rect 1255 1751 1261 1752
rect 1255 1750 1256 1751
rect 1247 1748 1256 1750
rect 1247 1747 1248 1748
rect 1242 1746 1248 1747
rect 1255 1747 1256 1748
rect 1260 1747 1261 1751
rect 1487 1751 1493 1752
rect 1487 1750 1488 1751
rect 1255 1746 1261 1747
rect 1459 1748 1488 1750
rect 754 1743 760 1744
rect 754 1739 755 1743
rect 759 1742 760 1743
rect 1459 1742 1461 1748
rect 1487 1747 1488 1748
rect 1492 1747 1493 1751
rect 4466 1751 4467 1755
rect 4471 1751 4472 1755
rect 4466 1750 4472 1751
rect 4530 1755 4536 1756
rect 4530 1751 4531 1755
rect 4535 1751 4536 1755
rect 4530 1750 4536 1751
rect 4666 1755 4672 1756
rect 4666 1751 4667 1755
rect 4671 1751 4672 1755
rect 4666 1750 4672 1751
rect 4802 1755 4808 1756
rect 4802 1751 4803 1755
rect 4807 1751 4808 1755
rect 4802 1750 4808 1751
rect 4938 1755 4944 1756
rect 4938 1751 4939 1755
rect 4943 1751 4944 1755
rect 4938 1750 4944 1751
rect 1487 1746 1493 1747
rect 2002 1747 2008 1748
rect 2002 1743 2003 1747
rect 2007 1746 2008 1747
rect 2119 1747 2125 1748
rect 2119 1746 2120 1747
rect 2007 1744 2120 1746
rect 2007 1743 2008 1744
rect 2002 1742 2008 1743
rect 2119 1743 2120 1744
rect 2124 1743 2125 1747
rect 2119 1742 2125 1743
rect 2127 1747 2133 1748
rect 2127 1743 2128 1747
rect 2132 1746 2133 1747
rect 2255 1747 2261 1748
rect 2255 1746 2256 1747
rect 2132 1744 2256 1746
rect 2132 1743 2133 1744
rect 2127 1742 2133 1743
rect 2255 1743 2256 1744
rect 2260 1743 2261 1747
rect 2255 1742 2261 1743
rect 2263 1747 2269 1748
rect 2263 1743 2264 1747
rect 2268 1746 2269 1747
rect 2391 1747 2397 1748
rect 2391 1746 2392 1747
rect 2268 1744 2392 1746
rect 2268 1743 2269 1744
rect 2263 1742 2269 1743
rect 2391 1743 2392 1744
rect 2396 1743 2397 1747
rect 2391 1742 2397 1743
rect 2415 1747 2421 1748
rect 2415 1743 2416 1747
rect 2420 1746 2421 1747
rect 2543 1747 2549 1748
rect 2543 1746 2544 1747
rect 2420 1744 2544 1746
rect 2420 1743 2421 1744
rect 2415 1742 2421 1743
rect 2543 1743 2544 1744
rect 2548 1743 2549 1747
rect 2543 1742 2549 1743
rect 2567 1747 2573 1748
rect 2567 1743 2568 1747
rect 2572 1746 2573 1747
rect 2703 1747 2709 1748
rect 2703 1746 2704 1747
rect 2572 1744 2704 1746
rect 2572 1743 2573 1744
rect 2567 1742 2573 1743
rect 2703 1743 2704 1744
rect 2708 1743 2709 1747
rect 2703 1742 2709 1743
rect 2722 1747 2728 1748
rect 2722 1743 2723 1747
rect 2727 1746 2728 1747
rect 2863 1747 2869 1748
rect 2863 1746 2864 1747
rect 2727 1744 2864 1746
rect 2727 1743 2728 1744
rect 2722 1742 2728 1743
rect 2863 1743 2864 1744
rect 2868 1743 2869 1747
rect 2863 1742 2869 1743
rect 3023 1747 3029 1748
rect 3023 1743 3024 1747
rect 3028 1746 3029 1747
rect 3031 1747 3037 1748
rect 3031 1746 3032 1747
rect 3028 1744 3032 1746
rect 3028 1743 3029 1744
rect 3023 1742 3029 1743
rect 3031 1743 3032 1744
rect 3036 1743 3037 1747
rect 3031 1742 3037 1743
rect 3175 1747 3184 1748
rect 3175 1743 3176 1747
rect 3183 1743 3184 1747
rect 3175 1742 3184 1743
rect 3322 1747 3333 1748
rect 3322 1743 3323 1747
rect 3327 1743 3328 1747
rect 3332 1743 3333 1747
rect 3322 1742 3333 1743
rect 3479 1747 3488 1748
rect 3479 1743 3480 1747
rect 3487 1743 3488 1747
rect 3479 1742 3488 1743
rect 3639 1747 3645 1748
rect 3639 1743 3640 1747
rect 3644 1746 3645 1747
rect 3647 1747 3653 1748
rect 3647 1746 3648 1747
rect 3644 1744 3648 1746
rect 3644 1743 3645 1744
rect 3639 1742 3645 1743
rect 3647 1743 3648 1744
rect 3652 1743 3653 1747
rect 3647 1742 3653 1743
rect 3770 1747 3781 1748
rect 3770 1743 3771 1747
rect 3775 1743 3776 1747
rect 3780 1743 3781 1747
rect 3770 1742 3781 1743
rect 759 1740 1461 1742
rect 1974 1740 1980 1741
rect 3798 1740 3804 1741
rect 759 1739 760 1740
rect 754 1738 760 1739
rect 1974 1736 1975 1740
rect 1979 1736 1980 1740
rect 1974 1735 1980 1736
rect 1994 1739 2000 1740
rect 1994 1735 1995 1739
rect 1999 1735 2000 1739
rect 1994 1734 2000 1735
rect 2130 1739 2136 1740
rect 2130 1735 2131 1739
rect 2135 1735 2136 1739
rect 2130 1734 2136 1735
rect 2266 1739 2272 1740
rect 2266 1735 2267 1739
rect 2271 1735 2272 1739
rect 2266 1734 2272 1735
rect 2418 1739 2424 1740
rect 2418 1735 2419 1739
rect 2423 1735 2424 1739
rect 2418 1734 2424 1735
rect 2578 1739 2584 1740
rect 2578 1735 2579 1739
rect 2583 1735 2584 1739
rect 2578 1734 2584 1735
rect 2738 1739 2744 1740
rect 2738 1735 2739 1739
rect 2743 1735 2744 1739
rect 2738 1734 2744 1735
rect 2898 1739 2904 1740
rect 2898 1735 2899 1739
rect 2903 1735 2904 1739
rect 2898 1734 2904 1735
rect 3050 1739 3056 1740
rect 3050 1735 3051 1739
rect 3055 1735 3056 1739
rect 3050 1734 3056 1735
rect 3202 1739 3208 1740
rect 3202 1735 3203 1739
rect 3207 1735 3208 1739
rect 3202 1734 3208 1735
rect 3354 1739 3360 1740
rect 3354 1735 3355 1739
rect 3359 1735 3360 1739
rect 3354 1734 3360 1735
rect 3514 1739 3520 1740
rect 3514 1735 3515 1739
rect 3519 1735 3520 1739
rect 3514 1734 3520 1735
rect 3650 1739 3656 1740
rect 3650 1735 3651 1739
rect 3655 1735 3656 1739
rect 3798 1736 3799 1740
rect 3803 1736 3804 1740
rect 3798 1735 3804 1736
rect 3650 1734 3656 1735
rect 2022 1724 2028 1725
rect 1974 1723 1980 1724
rect 383 1719 389 1720
rect 383 1718 384 1719
rect 285 1716 384 1718
rect 383 1715 384 1716
rect 388 1715 389 1719
rect 383 1714 389 1715
rect 486 1719 492 1720
rect 486 1715 487 1719
rect 491 1715 492 1719
rect 486 1714 492 1715
rect 754 1719 760 1720
rect 754 1715 755 1719
rect 759 1715 760 1719
rect 754 1714 760 1715
rect 914 1719 920 1720
rect 914 1715 915 1719
rect 919 1715 920 1719
rect 914 1714 920 1715
rect 1146 1719 1152 1720
rect 1146 1715 1147 1719
rect 1151 1715 1152 1719
rect 1146 1714 1152 1715
rect 1378 1719 1384 1720
rect 1378 1715 1379 1719
rect 1383 1715 1384 1719
rect 1974 1719 1975 1723
rect 1979 1719 1980 1723
rect 2022 1720 2023 1724
rect 2027 1720 2028 1724
rect 2022 1719 2028 1720
rect 2158 1724 2164 1725
rect 2158 1720 2159 1724
rect 2163 1720 2164 1724
rect 2158 1719 2164 1720
rect 2294 1724 2300 1725
rect 2294 1720 2295 1724
rect 2299 1720 2300 1724
rect 2294 1719 2300 1720
rect 2446 1724 2452 1725
rect 2446 1720 2447 1724
rect 2451 1720 2452 1724
rect 2446 1719 2452 1720
rect 2606 1724 2612 1725
rect 2606 1720 2607 1724
rect 2611 1720 2612 1724
rect 2606 1719 2612 1720
rect 2766 1724 2772 1725
rect 2766 1720 2767 1724
rect 2771 1720 2772 1724
rect 2766 1719 2772 1720
rect 2926 1724 2932 1725
rect 2926 1720 2927 1724
rect 2931 1720 2932 1724
rect 2926 1719 2932 1720
rect 3078 1724 3084 1725
rect 3078 1720 3079 1724
rect 3083 1720 3084 1724
rect 3078 1719 3084 1720
rect 3230 1724 3236 1725
rect 3230 1720 3231 1724
rect 3235 1720 3236 1724
rect 3230 1719 3236 1720
rect 3382 1724 3388 1725
rect 3382 1720 3383 1724
rect 3387 1720 3388 1724
rect 3382 1719 3388 1720
rect 3542 1724 3548 1725
rect 3542 1720 3543 1724
rect 3547 1720 3548 1724
rect 3542 1719 3548 1720
rect 3678 1724 3684 1725
rect 3678 1720 3679 1724
rect 3683 1720 3684 1724
rect 3678 1719 3684 1720
rect 3798 1723 3804 1724
rect 3798 1719 3799 1723
rect 3803 1719 3804 1723
rect 1974 1718 1980 1719
rect 3798 1718 3804 1719
rect 1378 1714 1384 1715
rect 4695 1691 4701 1692
rect 4695 1690 4696 1691
rect 4653 1688 4696 1690
rect 4695 1687 4696 1688
rect 4700 1687 4701 1691
rect 4950 1691 4956 1692
rect 4950 1690 4951 1691
rect 4925 1688 4951 1690
rect 4695 1686 4701 1687
rect 4950 1687 4951 1688
rect 4955 1687 4956 1691
rect 4950 1686 4956 1687
rect 5098 1691 5104 1692
rect 5098 1687 5099 1691
rect 5103 1690 5104 1691
rect 5370 1691 5376 1692
rect 5103 1688 5125 1690
rect 5103 1687 5104 1688
rect 5098 1686 5104 1687
rect 5330 1687 5336 1688
rect 4784 1682 4786 1685
rect 4831 1683 4837 1684
rect 4831 1682 4832 1683
rect 4784 1680 4832 1682
rect 4831 1679 4832 1680
rect 4836 1679 4837 1683
rect 4831 1678 4837 1679
rect 5056 1674 5058 1685
rect 5330 1683 5331 1687
rect 5335 1683 5336 1687
rect 5370 1687 5371 1691
rect 5375 1690 5376 1691
rect 5618 1691 5624 1692
rect 5618 1690 5619 1691
rect 5375 1688 5397 1690
rect 5605 1688 5619 1690
rect 5375 1687 5376 1688
rect 5370 1686 5376 1687
rect 5618 1687 5619 1688
rect 5623 1687 5624 1691
rect 5618 1686 5624 1687
rect 5330 1682 5336 1683
rect 5327 1675 5333 1676
rect 5327 1674 5328 1675
rect 5056 1672 5328 1674
rect 5327 1671 5328 1672
rect 5332 1671 5333 1675
rect 5327 1670 5333 1671
rect 5330 1663 5336 1664
rect 258 1659 264 1660
rect 218 1655 224 1656
rect 218 1651 219 1655
rect 223 1651 224 1655
rect 258 1655 259 1659
rect 263 1658 264 1659
rect 815 1659 821 1660
rect 815 1658 816 1659
rect 263 1656 381 1658
rect 709 1656 816 1658
rect 263 1655 264 1656
rect 258 1654 264 1655
rect 815 1655 816 1656
rect 820 1655 821 1659
rect 1242 1659 1248 1660
rect 1242 1658 1243 1659
rect 1229 1656 1243 1658
rect 815 1654 821 1655
rect 962 1655 968 1656
rect 218 1650 224 1651
rect 962 1651 963 1655
rect 967 1651 968 1655
rect 1242 1655 1243 1656
rect 1247 1655 1248 1659
rect 5330 1659 5331 1663
rect 5335 1662 5336 1663
rect 5335 1660 5643 1662
rect 5335 1659 5336 1660
rect 5330 1658 5336 1659
rect 5641 1656 5643 1660
rect 1242 1654 1248 1655
rect 4650 1655 4656 1656
rect 962 1650 968 1651
rect 1974 1653 1980 1654
rect 3798 1653 3804 1654
rect 1974 1649 1975 1653
rect 1979 1649 1980 1653
rect 1974 1648 1980 1649
rect 2022 1652 2028 1653
rect 2022 1648 2023 1652
rect 2027 1648 2028 1652
rect 2022 1647 2028 1648
rect 2166 1652 2172 1653
rect 2166 1648 2167 1652
rect 2171 1648 2172 1652
rect 2166 1647 2172 1648
rect 2318 1652 2324 1653
rect 2318 1648 2319 1652
rect 2323 1648 2324 1652
rect 2318 1647 2324 1648
rect 2478 1652 2484 1653
rect 2478 1648 2479 1652
rect 2483 1648 2484 1652
rect 2478 1647 2484 1648
rect 2638 1652 2644 1653
rect 2638 1648 2639 1652
rect 2643 1648 2644 1652
rect 2638 1647 2644 1648
rect 2790 1652 2796 1653
rect 2790 1648 2791 1652
rect 2795 1648 2796 1652
rect 2790 1647 2796 1648
rect 2942 1652 2948 1653
rect 2942 1648 2943 1652
rect 2947 1648 2948 1652
rect 2942 1647 2948 1648
rect 3102 1652 3108 1653
rect 3102 1648 3103 1652
rect 3107 1648 3108 1652
rect 3102 1647 3108 1648
rect 3262 1652 3268 1653
rect 3262 1648 3263 1652
rect 3267 1648 3268 1652
rect 3262 1647 3268 1648
rect 3422 1652 3428 1653
rect 3422 1648 3423 1652
rect 3427 1648 3428 1652
rect 3798 1649 3799 1653
rect 3803 1649 3804 1653
rect 4650 1651 4651 1655
rect 4655 1654 4656 1655
rect 4687 1655 4693 1656
rect 4687 1654 4688 1655
rect 4655 1652 4688 1654
rect 4655 1651 4656 1652
rect 4650 1650 4656 1651
rect 4687 1651 4688 1652
rect 4692 1651 4693 1655
rect 4687 1650 4693 1651
rect 4695 1655 4701 1656
rect 4695 1651 4696 1655
rect 4700 1654 4701 1655
rect 4823 1655 4829 1656
rect 4823 1654 4824 1655
rect 4700 1652 4824 1654
rect 4700 1651 4701 1652
rect 4695 1650 4701 1651
rect 4823 1651 4824 1652
rect 4828 1651 4829 1655
rect 4823 1650 4829 1651
rect 4831 1655 4837 1656
rect 4831 1651 4832 1655
rect 4836 1654 4837 1655
rect 4959 1655 4965 1656
rect 4959 1654 4960 1655
rect 4836 1652 4960 1654
rect 4836 1651 4837 1652
rect 4831 1650 4837 1651
rect 4959 1651 4960 1652
rect 4964 1651 4965 1655
rect 4959 1650 4965 1651
rect 5095 1655 5104 1656
rect 5095 1651 5096 1655
rect 5103 1651 5104 1655
rect 5095 1650 5104 1651
rect 5231 1655 5237 1656
rect 5231 1651 5232 1655
rect 5236 1654 5237 1655
rect 5338 1655 5344 1656
rect 5338 1654 5339 1655
rect 5236 1652 5339 1654
rect 5236 1651 5237 1652
rect 5231 1650 5237 1651
rect 5338 1651 5339 1652
rect 5343 1651 5344 1655
rect 5338 1650 5344 1651
rect 5367 1655 5376 1656
rect 5367 1651 5368 1655
rect 5375 1651 5376 1655
rect 5367 1650 5376 1651
rect 5502 1655 5509 1656
rect 5502 1651 5503 1655
rect 5508 1651 5509 1655
rect 5502 1650 5509 1651
rect 5639 1655 5645 1656
rect 5639 1651 5640 1655
rect 5644 1651 5645 1655
rect 5639 1650 5645 1651
rect 3798 1648 3804 1649
rect 3838 1648 3844 1649
rect 5662 1648 5668 1649
rect 3422 1647 3428 1648
rect 3838 1644 3839 1648
rect 3843 1644 3844 1648
rect 3838 1643 3844 1644
rect 4562 1647 4568 1648
rect 4562 1643 4563 1647
rect 4567 1643 4568 1647
rect 4562 1642 4568 1643
rect 4698 1647 4704 1648
rect 4698 1643 4699 1647
rect 4703 1643 4704 1647
rect 4698 1642 4704 1643
rect 4834 1647 4840 1648
rect 4834 1643 4835 1647
rect 4839 1643 4840 1647
rect 4834 1642 4840 1643
rect 4970 1647 4976 1648
rect 4970 1643 4971 1647
rect 4975 1643 4976 1647
rect 4970 1642 4976 1643
rect 5106 1647 5112 1648
rect 5106 1643 5107 1647
rect 5111 1643 5112 1647
rect 5106 1642 5112 1643
rect 5242 1647 5248 1648
rect 5242 1643 5243 1647
rect 5247 1643 5248 1647
rect 5242 1642 5248 1643
rect 5378 1647 5384 1648
rect 5378 1643 5379 1647
rect 5383 1643 5384 1647
rect 5378 1642 5384 1643
rect 5514 1647 5520 1648
rect 5514 1643 5515 1647
rect 5519 1643 5520 1647
rect 5662 1644 5663 1648
rect 5667 1644 5668 1648
rect 5662 1643 5668 1644
rect 5514 1642 5520 1643
rect 1994 1637 2000 1638
rect 1974 1636 1980 1637
rect 962 1635 968 1636
rect 962 1631 963 1635
rect 967 1634 968 1635
rect 967 1632 1162 1634
rect 967 1631 968 1632
rect 962 1630 968 1631
rect 255 1623 264 1624
rect 255 1619 256 1623
rect 263 1619 264 1623
rect 255 1618 264 1619
rect 486 1623 493 1624
rect 486 1619 487 1623
rect 492 1619 493 1623
rect 486 1618 493 1619
rect 570 1623 576 1624
rect 570 1619 571 1623
rect 575 1622 576 1623
rect 743 1623 749 1624
rect 743 1622 744 1623
rect 575 1620 744 1622
rect 575 1619 576 1620
rect 570 1618 576 1619
rect 743 1619 744 1620
rect 748 1619 749 1623
rect 743 1618 749 1619
rect 815 1623 821 1624
rect 815 1619 816 1623
rect 820 1622 821 1623
rect 999 1623 1005 1624
rect 999 1622 1000 1623
rect 820 1620 1000 1622
rect 820 1619 821 1620
rect 815 1618 821 1619
rect 999 1619 1000 1620
rect 1004 1619 1005 1623
rect 1160 1622 1162 1632
rect 1974 1632 1975 1636
rect 1979 1632 1980 1636
rect 1994 1633 1995 1637
rect 1999 1633 2000 1637
rect 1994 1632 2000 1633
rect 2138 1637 2144 1638
rect 2138 1633 2139 1637
rect 2143 1633 2144 1637
rect 2138 1632 2144 1633
rect 2290 1637 2296 1638
rect 2290 1633 2291 1637
rect 2295 1633 2296 1637
rect 2290 1632 2296 1633
rect 2450 1637 2456 1638
rect 2450 1633 2451 1637
rect 2455 1633 2456 1637
rect 2450 1632 2456 1633
rect 2610 1637 2616 1638
rect 2610 1633 2611 1637
rect 2615 1633 2616 1637
rect 2610 1632 2616 1633
rect 2762 1637 2768 1638
rect 2762 1633 2763 1637
rect 2767 1633 2768 1637
rect 2762 1632 2768 1633
rect 2914 1637 2920 1638
rect 2914 1633 2915 1637
rect 2919 1633 2920 1637
rect 2914 1632 2920 1633
rect 3074 1637 3080 1638
rect 3074 1633 3075 1637
rect 3079 1633 3080 1637
rect 3074 1632 3080 1633
rect 3234 1637 3240 1638
rect 3234 1633 3235 1637
rect 3239 1633 3240 1637
rect 3234 1632 3240 1633
rect 3394 1637 3400 1638
rect 3394 1633 3395 1637
rect 3399 1633 3400 1637
rect 3394 1632 3400 1633
rect 3798 1636 3804 1637
rect 3798 1632 3799 1636
rect 3803 1632 3804 1636
rect 4590 1632 4596 1633
rect 1974 1631 1980 1632
rect 3798 1631 3804 1632
rect 3838 1631 3844 1632
rect 2119 1627 2125 1628
rect 1263 1623 1269 1624
rect 1263 1622 1264 1623
rect 1160 1620 1264 1622
rect 999 1618 1005 1619
rect 1263 1619 1264 1620
rect 1268 1619 1269 1623
rect 2119 1623 2120 1627
rect 2124 1626 2125 1627
rect 2154 1627 2160 1628
rect 2154 1626 2155 1627
rect 2124 1624 2155 1626
rect 2124 1623 2125 1624
rect 2119 1622 2125 1623
rect 2154 1623 2155 1624
rect 2159 1623 2160 1627
rect 2154 1622 2160 1623
rect 2263 1627 2269 1628
rect 2263 1623 2264 1627
rect 2268 1626 2269 1627
rect 2306 1627 2312 1628
rect 2306 1626 2307 1627
rect 2268 1624 2307 1626
rect 2268 1623 2269 1624
rect 2263 1622 2269 1623
rect 2306 1623 2307 1624
rect 2311 1623 2312 1627
rect 2306 1622 2312 1623
rect 2415 1627 2421 1628
rect 2415 1623 2416 1627
rect 2420 1626 2421 1627
rect 2466 1627 2472 1628
rect 2466 1626 2467 1627
rect 2420 1624 2467 1626
rect 2420 1623 2421 1624
rect 2415 1622 2421 1623
rect 2466 1623 2467 1624
rect 2471 1623 2472 1627
rect 2466 1622 2472 1623
rect 2575 1627 2581 1628
rect 2575 1623 2576 1627
rect 2580 1626 2581 1627
rect 2626 1627 2632 1628
rect 2626 1626 2627 1627
rect 2580 1624 2627 1626
rect 2580 1623 2581 1624
rect 2575 1622 2581 1623
rect 2626 1623 2627 1624
rect 2631 1623 2632 1627
rect 2626 1622 2632 1623
rect 2730 1627 2741 1628
rect 2730 1623 2731 1627
rect 2735 1623 2736 1627
rect 2740 1623 2741 1627
rect 2730 1622 2741 1623
rect 2887 1627 2893 1628
rect 2887 1623 2888 1627
rect 2892 1626 2893 1627
rect 2930 1627 2936 1628
rect 2930 1626 2931 1627
rect 2892 1624 2931 1626
rect 2892 1623 2893 1624
rect 2887 1622 2893 1623
rect 2930 1623 2931 1624
rect 2935 1623 2936 1627
rect 2930 1622 2936 1623
rect 3039 1627 3045 1628
rect 3039 1623 3040 1627
rect 3044 1626 3045 1627
rect 3090 1627 3096 1628
rect 3090 1626 3091 1627
rect 3044 1624 3091 1626
rect 3044 1623 3045 1624
rect 3039 1622 3045 1623
rect 3090 1623 3091 1624
rect 3095 1623 3096 1627
rect 3090 1622 3096 1623
rect 3199 1627 3205 1628
rect 3199 1623 3200 1627
rect 3204 1626 3205 1627
rect 3215 1627 3221 1628
rect 3215 1626 3216 1627
rect 3204 1624 3216 1626
rect 3204 1623 3205 1624
rect 3199 1622 3205 1623
rect 3215 1623 3216 1624
rect 3220 1623 3221 1627
rect 3215 1622 3221 1623
rect 3359 1627 3365 1628
rect 3359 1623 3360 1627
rect 3364 1626 3365 1627
rect 3410 1627 3416 1628
rect 3410 1626 3411 1627
rect 3364 1624 3411 1626
rect 3364 1623 3365 1624
rect 3359 1622 3365 1623
rect 3410 1623 3411 1624
rect 3415 1623 3416 1627
rect 3519 1627 3525 1628
rect 3519 1626 3520 1627
rect 3410 1622 3416 1623
rect 3420 1624 3520 1626
rect 1263 1618 1269 1619
rect 2850 1619 2856 1620
rect 110 1616 116 1617
rect 1934 1616 1940 1617
rect 110 1612 111 1616
rect 115 1612 116 1616
rect 110 1611 116 1612
rect 130 1615 136 1616
rect 130 1611 131 1615
rect 135 1611 136 1615
rect 130 1610 136 1611
rect 362 1615 368 1616
rect 362 1611 363 1615
rect 367 1611 368 1615
rect 362 1610 368 1611
rect 618 1615 624 1616
rect 618 1611 619 1615
rect 623 1611 624 1615
rect 618 1610 624 1611
rect 874 1615 880 1616
rect 874 1611 875 1615
rect 879 1611 880 1615
rect 874 1610 880 1611
rect 1138 1615 1144 1616
rect 1138 1611 1139 1615
rect 1143 1611 1144 1615
rect 1934 1612 1935 1616
rect 1939 1612 1940 1616
rect 2850 1615 2851 1619
rect 2855 1618 2856 1619
rect 3420 1618 3422 1624
rect 3519 1623 3520 1624
rect 3524 1623 3525 1627
rect 3838 1627 3839 1631
rect 3843 1627 3844 1631
rect 4590 1628 4591 1632
rect 4595 1628 4596 1632
rect 4590 1627 4596 1628
rect 4726 1632 4732 1633
rect 4726 1628 4727 1632
rect 4731 1628 4732 1632
rect 4726 1627 4732 1628
rect 4862 1632 4868 1633
rect 4862 1628 4863 1632
rect 4867 1628 4868 1632
rect 4862 1627 4868 1628
rect 4998 1632 5004 1633
rect 4998 1628 4999 1632
rect 5003 1628 5004 1632
rect 4998 1627 5004 1628
rect 5134 1632 5140 1633
rect 5134 1628 5135 1632
rect 5139 1628 5140 1632
rect 5134 1627 5140 1628
rect 5270 1632 5276 1633
rect 5270 1628 5271 1632
rect 5275 1628 5276 1632
rect 5270 1627 5276 1628
rect 5406 1632 5412 1633
rect 5406 1628 5407 1632
rect 5411 1628 5412 1632
rect 5406 1627 5412 1628
rect 5542 1632 5548 1633
rect 5542 1628 5543 1632
rect 5547 1628 5548 1632
rect 5542 1627 5548 1628
rect 5662 1631 5668 1632
rect 5662 1627 5663 1631
rect 5667 1627 5668 1631
rect 3838 1626 3844 1627
rect 5662 1626 5668 1627
rect 3519 1622 3525 1623
rect 2855 1616 3422 1618
rect 2855 1615 2856 1616
rect 2850 1614 2856 1615
rect 1934 1611 1940 1612
rect 1138 1610 1144 1611
rect 158 1600 164 1601
rect 110 1599 116 1600
rect 110 1595 111 1599
rect 115 1595 116 1599
rect 158 1596 159 1600
rect 163 1596 164 1600
rect 158 1595 164 1596
rect 390 1600 396 1601
rect 390 1596 391 1600
rect 395 1596 396 1600
rect 390 1595 396 1596
rect 646 1600 652 1601
rect 646 1596 647 1600
rect 651 1596 652 1600
rect 646 1595 652 1596
rect 902 1600 908 1601
rect 902 1596 903 1600
rect 907 1596 908 1600
rect 902 1595 908 1596
rect 1166 1600 1172 1601
rect 1166 1596 1167 1600
rect 1171 1596 1172 1600
rect 1166 1595 1172 1596
rect 1934 1599 1940 1600
rect 1934 1595 1935 1599
rect 1939 1595 1940 1599
rect 110 1594 116 1595
rect 1934 1594 1940 1595
rect 2090 1595 2096 1596
rect 2090 1594 2091 1595
rect 2085 1592 2091 1594
rect 2090 1591 2091 1592
rect 2095 1591 2096 1595
rect 2090 1590 2096 1591
rect 2154 1595 2160 1596
rect 2154 1591 2155 1595
rect 2159 1591 2160 1595
rect 2154 1590 2160 1591
rect 2306 1595 2312 1596
rect 2306 1591 2307 1595
rect 2311 1591 2312 1595
rect 2306 1590 2312 1591
rect 2466 1595 2472 1596
rect 2466 1591 2467 1595
rect 2471 1591 2472 1595
rect 2466 1590 2472 1591
rect 2626 1595 2632 1596
rect 2626 1591 2627 1595
rect 2631 1591 2632 1595
rect 2626 1590 2632 1591
rect 2850 1595 2856 1596
rect 2850 1591 2851 1595
rect 2855 1591 2856 1595
rect 2850 1590 2856 1591
rect 2930 1595 2936 1596
rect 2930 1591 2931 1595
rect 2935 1591 2936 1595
rect 2930 1590 2936 1591
rect 3090 1595 3096 1596
rect 3090 1591 3091 1595
rect 3095 1591 3096 1595
rect 3090 1590 3096 1591
rect 3322 1595 3328 1596
rect 3322 1591 3323 1595
rect 3327 1591 3328 1595
rect 3322 1590 3328 1591
rect 3410 1595 3416 1596
rect 3410 1591 3411 1595
rect 3415 1591 3416 1595
rect 3410 1590 3416 1591
rect 3838 1557 3844 1558
rect 5662 1557 5668 1558
rect 3838 1553 3839 1557
rect 3843 1553 3844 1557
rect 3838 1552 3844 1553
rect 4590 1556 4596 1557
rect 4590 1552 4591 1556
rect 4595 1552 4596 1556
rect 4590 1551 4596 1552
rect 4726 1556 4732 1557
rect 4726 1552 4727 1556
rect 4731 1552 4732 1556
rect 4726 1551 4732 1552
rect 4862 1556 4868 1557
rect 4862 1552 4863 1556
rect 4867 1552 4868 1556
rect 4862 1551 4868 1552
rect 4998 1556 5004 1557
rect 4998 1552 4999 1556
rect 5003 1552 5004 1556
rect 4998 1551 5004 1552
rect 5134 1556 5140 1557
rect 5134 1552 5135 1556
rect 5139 1552 5140 1556
rect 5134 1551 5140 1552
rect 5270 1556 5276 1557
rect 5270 1552 5271 1556
rect 5275 1552 5276 1556
rect 5270 1551 5276 1552
rect 5406 1556 5412 1557
rect 5406 1552 5407 1556
rect 5411 1552 5412 1556
rect 5406 1551 5412 1552
rect 5542 1556 5548 1557
rect 5542 1552 5543 1556
rect 5547 1552 5548 1556
rect 5662 1553 5663 1557
rect 5667 1553 5668 1557
rect 5662 1552 5668 1553
rect 5542 1551 5548 1552
rect 4562 1541 4568 1542
rect 3838 1540 3844 1541
rect 3838 1536 3839 1540
rect 3843 1536 3844 1540
rect 4562 1537 4563 1541
rect 4567 1537 4568 1541
rect 4562 1536 4568 1537
rect 4698 1541 4704 1542
rect 4698 1537 4699 1541
rect 4703 1537 4704 1541
rect 4698 1536 4704 1537
rect 4834 1541 4840 1542
rect 4834 1537 4835 1541
rect 4839 1537 4840 1541
rect 4834 1536 4840 1537
rect 4970 1541 4976 1542
rect 4970 1537 4971 1541
rect 4975 1537 4976 1541
rect 4970 1536 4976 1537
rect 5106 1541 5112 1542
rect 5106 1537 5107 1541
rect 5111 1537 5112 1541
rect 5106 1536 5112 1537
rect 5242 1541 5248 1542
rect 5242 1537 5243 1541
rect 5247 1537 5248 1541
rect 5242 1536 5248 1537
rect 5378 1541 5384 1542
rect 5378 1537 5379 1541
rect 5383 1537 5384 1541
rect 5378 1536 5384 1537
rect 5514 1541 5520 1542
rect 5514 1537 5515 1541
rect 5519 1537 5520 1541
rect 5514 1536 5520 1537
rect 5662 1540 5668 1541
rect 5662 1536 5663 1540
rect 5667 1536 5668 1540
rect 2127 1535 2133 1536
rect 2127 1534 2128 1535
rect 2085 1532 2128 1534
rect 2127 1531 2128 1532
rect 2132 1531 2133 1535
rect 2127 1530 2133 1531
rect 2258 1535 2264 1536
rect 2258 1531 2259 1535
rect 2263 1534 2264 1535
rect 2807 1535 2813 1536
rect 2807 1534 2808 1535
rect 2263 1532 2285 1534
rect 2765 1532 2808 1534
rect 2263 1531 2264 1532
rect 2258 1530 2264 1531
rect 2626 1531 2632 1532
rect 110 1529 116 1530
rect 1934 1529 1940 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 158 1528 164 1529
rect 158 1524 159 1528
rect 163 1524 164 1528
rect 158 1523 164 1524
rect 326 1528 332 1529
rect 326 1524 327 1528
rect 331 1524 332 1528
rect 326 1523 332 1524
rect 510 1528 516 1529
rect 510 1524 511 1528
rect 515 1524 516 1528
rect 510 1523 516 1524
rect 694 1528 700 1529
rect 694 1524 695 1528
rect 699 1524 700 1528
rect 694 1523 700 1524
rect 886 1528 892 1529
rect 886 1524 887 1528
rect 891 1524 892 1528
rect 886 1523 892 1524
rect 1078 1528 1084 1529
rect 1078 1524 1079 1528
rect 1083 1524 1084 1528
rect 1934 1525 1935 1529
rect 1939 1525 1940 1529
rect 1934 1524 1940 1525
rect 2216 1526 2218 1529
rect 2263 1527 2269 1528
rect 2263 1526 2264 1527
rect 2216 1524 2264 1526
rect 1078 1523 1084 1524
rect 2263 1523 2264 1524
rect 2268 1523 2269 1527
rect 2263 1522 2269 1523
rect 2488 1518 2490 1529
rect 2626 1527 2627 1531
rect 2631 1527 2632 1531
rect 2807 1531 2808 1532
rect 2812 1531 2813 1535
rect 2943 1535 2949 1536
rect 2943 1534 2944 1535
rect 2901 1532 2944 1534
rect 2807 1530 2813 1531
rect 2943 1531 2944 1532
rect 2948 1531 2949 1535
rect 3079 1535 3085 1536
rect 3079 1534 3080 1535
rect 3037 1532 3080 1534
rect 2943 1530 2949 1531
rect 3079 1531 3080 1532
rect 3084 1531 3085 1535
rect 3079 1530 3085 1531
rect 3215 1535 3221 1536
rect 3215 1531 3216 1535
rect 3220 1534 3221 1535
rect 3351 1535 3357 1536
rect 3220 1532 3237 1534
rect 3220 1531 3221 1532
rect 3215 1530 3221 1531
rect 3351 1531 3352 1535
rect 3356 1534 3357 1535
rect 3487 1535 3493 1536
rect 3838 1535 3844 1536
rect 5662 1535 5668 1536
rect 3356 1532 3373 1534
rect 3356 1531 3357 1532
rect 3351 1530 3357 1531
rect 3487 1531 3488 1535
rect 3492 1534 3493 1535
rect 3492 1532 3509 1534
rect 3492 1531 3493 1532
rect 3487 1530 3493 1531
rect 4687 1531 4693 1532
rect 2626 1526 2632 1527
rect 2798 1519 2804 1520
rect 2798 1518 2799 1519
rect 2488 1516 2799 1518
rect 2798 1515 2799 1516
rect 2803 1515 2804 1519
rect 3168 1518 3170 1529
rect 4687 1527 4688 1531
rect 4692 1530 4693 1531
rect 4714 1531 4720 1532
rect 4714 1530 4715 1531
rect 4692 1528 4715 1530
rect 4692 1527 4693 1528
rect 4687 1526 4693 1527
rect 4714 1527 4715 1528
rect 4719 1527 4720 1531
rect 4714 1526 4720 1527
rect 4823 1531 4829 1532
rect 4823 1527 4824 1531
rect 4828 1530 4829 1531
rect 4850 1531 4856 1532
rect 4850 1530 4851 1531
rect 4828 1528 4851 1530
rect 4828 1527 4829 1528
rect 4823 1526 4829 1527
rect 4850 1527 4851 1528
rect 4855 1527 4856 1531
rect 4850 1526 4856 1527
rect 4959 1531 4965 1532
rect 4959 1527 4960 1531
rect 4964 1530 4965 1531
rect 4986 1531 4992 1532
rect 4986 1530 4987 1531
rect 4964 1528 4987 1530
rect 4964 1527 4965 1528
rect 4959 1526 4965 1527
rect 4986 1527 4987 1528
rect 4991 1527 4992 1531
rect 4986 1526 4992 1527
rect 5095 1531 5101 1532
rect 5095 1527 5096 1531
rect 5100 1530 5101 1531
rect 5122 1531 5128 1532
rect 5122 1530 5123 1531
rect 5100 1528 5123 1530
rect 5100 1527 5101 1528
rect 5095 1526 5101 1527
rect 5122 1527 5123 1528
rect 5127 1527 5128 1531
rect 5122 1526 5128 1527
rect 5231 1531 5237 1532
rect 5231 1527 5232 1531
rect 5236 1530 5237 1531
rect 5258 1531 5264 1532
rect 5258 1530 5259 1531
rect 5236 1528 5259 1530
rect 5236 1527 5237 1528
rect 5231 1526 5237 1527
rect 5258 1527 5259 1528
rect 5263 1527 5264 1531
rect 5258 1526 5264 1527
rect 5327 1531 5333 1532
rect 5327 1527 5328 1531
rect 5332 1530 5333 1531
rect 5367 1531 5373 1532
rect 5367 1530 5368 1531
rect 5332 1528 5368 1530
rect 5332 1527 5333 1528
rect 5327 1526 5333 1527
rect 5367 1527 5368 1528
rect 5372 1527 5373 1531
rect 5367 1526 5373 1527
rect 5503 1531 5509 1532
rect 5503 1527 5504 1531
rect 5508 1530 5509 1531
rect 5530 1531 5536 1532
rect 5530 1530 5531 1531
rect 5508 1528 5531 1530
rect 5508 1527 5509 1528
rect 5503 1526 5509 1527
rect 5530 1527 5531 1528
rect 5535 1527 5536 1531
rect 5530 1526 5536 1527
rect 5639 1531 5645 1532
rect 5639 1527 5640 1531
rect 5644 1527 5645 1531
rect 5639 1526 5645 1527
rect 5479 1523 5485 1524
rect 3614 1519 3620 1520
rect 3614 1518 3615 1519
rect 3168 1516 3615 1518
rect 2798 1514 2804 1515
rect 3614 1515 3615 1516
rect 3619 1515 3620 1519
rect 5479 1519 5480 1523
rect 5484 1522 5485 1523
rect 5641 1522 5643 1526
rect 5484 1520 5643 1522
rect 5484 1519 5485 1520
rect 5479 1518 5485 1519
rect 3614 1514 3620 1515
rect 130 1513 136 1514
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 130 1509 131 1513
rect 135 1509 136 1513
rect 130 1508 136 1509
rect 298 1513 304 1514
rect 298 1509 299 1513
rect 303 1509 304 1513
rect 298 1508 304 1509
rect 482 1513 488 1514
rect 482 1509 483 1513
rect 487 1509 488 1513
rect 482 1508 488 1509
rect 666 1513 672 1514
rect 666 1509 667 1513
rect 671 1509 672 1513
rect 666 1508 672 1509
rect 858 1513 864 1514
rect 858 1509 859 1513
rect 863 1509 864 1513
rect 858 1508 864 1509
rect 1050 1513 1056 1514
rect 1050 1509 1051 1513
rect 1055 1509 1056 1513
rect 1050 1508 1056 1509
rect 1934 1512 1940 1513
rect 1934 1508 1935 1512
rect 1939 1508 1940 1512
rect 110 1507 116 1508
rect 1934 1507 1940 1508
rect 218 1503 224 1504
rect 218 1499 219 1503
rect 223 1502 224 1503
rect 255 1503 261 1504
rect 255 1502 256 1503
rect 223 1500 256 1502
rect 223 1499 224 1500
rect 218 1498 224 1499
rect 255 1499 256 1500
rect 260 1499 261 1503
rect 255 1498 261 1499
rect 286 1503 292 1504
rect 286 1499 287 1503
rect 291 1502 292 1503
rect 423 1503 429 1504
rect 423 1502 424 1503
rect 291 1500 424 1502
rect 291 1499 292 1500
rect 286 1498 292 1499
rect 423 1499 424 1500
rect 428 1499 429 1503
rect 423 1498 429 1499
rect 607 1503 613 1504
rect 607 1499 608 1503
rect 612 1502 613 1503
rect 682 1503 688 1504
rect 682 1502 683 1503
rect 612 1500 683 1502
rect 612 1499 613 1500
rect 607 1498 613 1499
rect 682 1499 683 1500
rect 687 1499 688 1503
rect 682 1498 688 1499
rect 791 1503 797 1504
rect 791 1499 792 1503
rect 796 1502 797 1503
rect 874 1503 880 1504
rect 874 1502 875 1503
rect 796 1500 875 1502
rect 796 1499 797 1500
rect 791 1498 797 1499
rect 874 1499 875 1500
rect 879 1499 880 1503
rect 874 1498 880 1499
rect 983 1503 989 1504
rect 983 1499 984 1503
rect 988 1502 989 1503
rect 1066 1503 1072 1504
rect 1066 1502 1067 1503
rect 988 1500 1067 1502
rect 988 1499 989 1500
rect 983 1498 989 1499
rect 1066 1499 1067 1500
rect 1071 1499 1072 1503
rect 1175 1503 1181 1504
rect 1175 1502 1176 1503
rect 1066 1498 1072 1499
rect 1076 1500 1176 1502
rect 802 1495 808 1496
rect 802 1491 803 1495
rect 807 1494 808 1495
rect 1076 1494 1078 1500
rect 1175 1499 1176 1500
rect 1180 1499 1181 1503
rect 1175 1498 1181 1499
rect 2090 1499 2096 1500
rect 2090 1495 2091 1499
rect 2095 1498 2096 1499
rect 2119 1499 2125 1500
rect 2119 1498 2120 1499
rect 2095 1496 2120 1498
rect 2095 1495 2096 1496
rect 2090 1494 2096 1495
rect 2119 1495 2120 1496
rect 2124 1495 2125 1499
rect 2119 1494 2125 1495
rect 2127 1499 2133 1500
rect 2127 1495 2128 1499
rect 2132 1498 2133 1499
rect 2255 1499 2261 1500
rect 2255 1498 2256 1499
rect 2132 1496 2256 1498
rect 2132 1495 2133 1496
rect 2127 1494 2133 1495
rect 2255 1495 2256 1496
rect 2260 1495 2261 1499
rect 2255 1494 2261 1495
rect 2263 1499 2269 1500
rect 2263 1495 2264 1499
rect 2268 1498 2269 1499
rect 2391 1499 2397 1500
rect 2391 1498 2392 1499
rect 2268 1496 2392 1498
rect 2268 1495 2269 1496
rect 2263 1494 2269 1495
rect 2391 1495 2392 1496
rect 2396 1495 2397 1499
rect 2391 1494 2397 1495
rect 2527 1499 2533 1500
rect 2527 1495 2528 1499
rect 2532 1498 2533 1499
rect 2626 1499 2632 1500
rect 2626 1498 2627 1499
rect 2532 1496 2627 1498
rect 2532 1495 2533 1496
rect 2527 1494 2533 1495
rect 2626 1495 2627 1496
rect 2631 1495 2632 1499
rect 2626 1494 2632 1495
rect 2634 1499 2640 1500
rect 2634 1495 2635 1499
rect 2639 1498 2640 1499
rect 2663 1499 2669 1500
rect 2663 1498 2664 1499
rect 2639 1496 2664 1498
rect 2639 1495 2640 1496
rect 2634 1494 2640 1495
rect 2663 1495 2664 1496
rect 2668 1495 2669 1499
rect 2663 1494 2669 1495
rect 2798 1499 2805 1500
rect 2798 1495 2799 1499
rect 2804 1495 2805 1499
rect 2798 1494 2805 1495
rect 2807 1499 2813 1500
rect 2807 1495 2808 1499
rect 2812 1498 2813 1499
rect 2935 1499 2941 1500
rect 2935 1498 2936 1499
rect 2812 1496 2936 1498
rect 2812 1495 2813 1496
rect 2807 1494 2813 1495
rect 2935 1495 2936 1496
rect 2940 1495 2941 1499
rect 2935 1494 2941 1495
rect 2943 1499 2949 1500
rect 2943 1495 2944 1499
rect 2948 1498 2949 1499
rect 3071 1499 3077 1500
rect 3071 1498 3072 1499
rect 2948 1496 3072 1498
rect 2948 1495 2949 1496
rect 2943 1494 2949 1495
rect 3071 1495 3072 1496
rect 3076 1495 3077 1499
rect 3071 1494 3077 1495
rect 3079 1499 3085 1500
rect 3079 1495 3080 1499
rect 3084 1498 3085 1499
rect 3207 1499 3213 1500
rect 3207 1498 3208 1499
rect 3084 1496 3208 1498
rect 3084 1495 3085 1496
rect 3079 1494 3085 1495
rect 3207 1495 3208 1496
rect 3212 1495 3213 1499
rect 3207 1494 3213 1495
rect 3343 1499 3349 1500
rect 3343 1495 3344 1499
rect 3348 1498 3349 1499
rect 3351 1499 3357 1500
rect 3351 1498 3352 1499
rect 3348 1496 3352 1498
rect 3348 1495 3349 1496
rect 3343 1494 3349 1495
rect 3351 1495 3352 1496
rect 3356 1495 3357 1499
rect 3351 1494 3357 1495
rect 3479 1499 3485 1500
rect 3479 1495 3480 1499
rect 3484 1498 3485 1499
rect 3487 1499 3493 1500
rect 3487 1498 3488 1499
rect 3484 1496 3488 1498
rect 3484 1495 3485 1496
rect 3479 1494 3485 1495
rect 3487 1495 3488 1496
rect 3492 1495 3493 1499
rect 3487 1494 3493 1495
rect 3614 1499 3621 1500
rect 3614 1495 3615 1499
rect 3620 1495 3621 1499
rect 3614 1494 3621 1495
rect 4650 1499 4656 1500
rect 4650 1495 4651 1499
rect 4655 1495 4656 1499
rect 4650 1494 4656 1495
rect 4714 1499 4720 1500
rect 4714 1495 4715 1499
rect 4719 1495 4720 1499
rect 4714 1494 4720 1495
rect 4850 1499 4856 1500
rect 4850 1495 4851 1499
rect 4855 1495 4856 1499
rect 4850 1494 4856 1495
rect 4986 1499 4992 1500
rect 4986 1495 4987 1499
rect 4991 1495 4992 1499
rect 4986 1494 4992 1495
rect 5122 1499 5128 1500
rect 5122 1495 5123 1499
rect 5127 1495 5128 1499
rect 5122 1494 5128 1495
rect 5258 1499 5264 1500
rect 5258 1495 5259 1499
rect 5263 1495 5264 1499
rect 5258 1494 5264 1495
rect 5338 1499 5344 1500
rect 5338 1495 5339 1499
rect 5343 1498 5344 1499
rect 5530 1499 5536 1500
rect 5343 1496 5397 1498
rect 5343 1495 5344 1496
rect 5338 1494 5344 1495
rect 5530 1495 5531 1499
rect 5535 1495 5536 1499
rect 5530 1494 5536 1495
rect 807 1492 1078 1494
rect 1974 1492 1980 1493
rect 3798 1492 3804 1493
rect 807 1491 808 1492
rect 802 1490 808 1491
rect 1974 1488 1975 1492
rect 1979 1488 1980 1492
rect 1974 1487 1980 1488
rect 1994 1491 2000 1492
rect 1994 1487 1995 1491
rect 1999 1487 2000 1491
rect 1994 1486 2000 1487
rect 2130 1491 2136 1492
rect 2130 1487 2131 1491
rect 2135 1487 2136 1491
rect 2130 1486 2136 1487
rect 2266 1491 2272 1492
rect 2266 1487 2267 1491
rect 2271 1487 2272 1491
rect 2266 1486 2272 1487
rect 2402 1491 2408 1492
rect 2402 1487 2403 1491
rect 2407 1487 2408 1491
rect 2402 1486 2408 1487
rect 2538 1491 2544 1492
rect 2538 1487 2539 1491
rect 2543 1487 2544 1491
rect 2538 1486 2544 1487
rect 2674 1491 2680 1492
rect 2674 1487 2675 1491
rect 2679 1487 2680 1491
rect 2674 1486 2680 1487
rect 2810 1491 2816 1492
rect 2810 1487 2811 1491
rect 2815 1487 2816 1491
rect 2810 1486 2816 1487
rect 2946 1491 2952 1492
rect 2946 1487 2947 1491
rect 2951 1487 2952 1491
rect 2946 1486 2952 1487
rect 3082 1491 3088 1492
rect 3082 1487 3083 1491
rect 3087 1487 3088 1491
rect 3082 1486 3088 1487
rect 3218 1491 3224 1492
rect 3218 1487 3219 1491
rect 3223 1487 3224 1491
rect 3218 1486 3224 1487
rect 3354 1491 3360 1492
rect 3354 1487 3355 1491
rect 3359 1487 3360 1491
rect 3354 1486 3360 1487
rect 3490 1491 3496 1492
rect 3490 1487 3491 1491
rect 3495 1487 3496 1491
rect 3798 1488 3799 1492
rect 3803 1488 3804 1492
rect 3798 1487 3804 1488
rect 3490 1486 3496 1487
rect 2022 1476 2028 1477
rect 1974 1475 1980 1476
rect 286 1471 292 1472
rect 286 1470 287 1471
rect 221 1468 287 1470
rect 286 1467 287 1468
rect 291 1467 292 1471
rect 286 1466 292 1467
rect 386 1471 392 1472
rect 386 1467 387 1471
rect 391 1467 392 1471
rect 386 1466 392 1467
rect 570 1471 576 1472
rect 570 1467 571 1471
rect 575 1467 576 1471
rect 570 1466 576 1467
rect 682 1471 688 1472
rect 682 1467 683 1471
rect 687 1467 688 1471
rect 682 1466 688 1467
rect 874 1471 880 1472
rect 874 1467 875 1471
rect 879 1467 880 1471
rect 874 1466 880 1467
rect 1066 1471 1072 1472
rect 1066 1467 1067 1471
rect 1071 1467 1072 1471
rect 1974 1471 1975 1475
rect 1979 1471 1980 1475
rect 2022 1472 2023 1476
rect 2027 1472 2028 1476
rect 2022 1471 2028 1472
rect 2158 1476 2164 1477
rect 2158 1472 2159 1476
rect 2163 1472 2164 1476
rect 2158 1471 2164 1472
rect 2294 1476 2300 1477
rect 2294 1472 2295 1476
rect 2299 1472 2300 1476
rect 2294 1471 2300 1472
rect 2430 1476 2436 1477
rect 2430 1472 2431 1476
rect 2435 1472 2436 1476
rect 2430 1471 2436 1472
rect 2566 1476 2572 1477
rect 2566 1472 2567 1476
rect 2571 1472 2572 1476
rect 2566 1471 2572 1472
rect 2702 1476 2708 1477
rect 2702 1472 2703 1476
rect 2707 1472 2708 1476
rect 2702 1471 2708 1472
rect 2838 1476 2844 1477
rect 2838 1472 2839 1476
rect 2843 1472 2844 1476
rect 2838 1471 2844 1472
rect 2974 1476 2980 1477
rect 2974 1472 2975 1476
rect 2979 1472 2980 1476
rect 2974 1471 2980 1472
rect 3110 1476 3116 1477
rect 3110 1472 3111 1476
rect 3115 1472 3116 1476
rect 3110 1471 3116 1472
rect 3246 1476 3252 1477
rect 3246 1472 3247 1476
rect 3251 1472 3252 1476
rect 3246 1471 3252 1472
rect 3382 1476 3388 1477
rect 3382 1472 3383 1476
rect 3387 1472 3388 1476
rect 3382 1471 3388 1472
rect 3518 1476 3524 1477
rect 3518 1472 3519 1476
rect 3523 1472 3524 1476
rect 3518 1471 3524 1472
rect 3798 1475 3804 1476
rect 3798 1471 3799 1475
rect 3803 1471 3804 1475
rect 1974 1470 1980 1471
rect 3798 1470 3804 1471
rect 1066 1466 1072 1467
rect 258 1411 264 1412
rect 218 1407 224 1408
rect 218 1403 219 1407
rect 223 1403 224 1407
rect 258 1407 259 1411
rect 263 1410 264 1411
rect 802 1411 808 1412
rect 802 1410 803 1411
rect 263 1408 413 1410
rect 773 1408 803 1410
rect 263 1407 264 1408
rect 258 1406 264 1407
rect 802 1407 803 1408
rect 807 1407 808 1411
rect 802 1406 808 1407
rect 810 1411 816 1412
rect 810 1407 811 1411
rect 815 1410 816 1411
rect 1098 1411 1104 1412
rect 815 1408 989 1410
rect 815 1407 816 1408
rect 810 1406 816 1407
rect 1098 1407 1099 1411
rect 1103 1410 1104 1411
rect 1103 1408 1277 1410
rect 1103 1407 1104 1408
rect 1098 1406 1104 1407
rect 218 1402 224 1403
rect 1974 1405 1980 1406
rect 3798 1405 3804 1406
rect 1974 1401 1975 1405
rect 1979 1401 1980 1405
rect 1974 1400 1980 1401
rect 2166 1404 2172 1405
rect 2166 1400 2167 1404
rect 2171 1400 2172 1404
rect 2166 1399 2172 1400
rect 2302 1404 2308 1405
rect 2302 1400 2303 1404
rect 2307 1400 2308 1404
rect 2302 1399 2308 1400
rect 2438 1404 2444 1405
rect 2438 1400 2439 1404
rect 2443 1400 2444 1404
rect 2438 1399 2444 1400
rect 2574 1404 2580 1405
rect 2574 1400 2575 1404
rect 2579 1400 2580 1404
rect 2574 1399 2580 1400
rect 2710 1404 2716 1405
rect 2710 1400 2711 1404
rect 2715 1400 2716 1404
rect 2710 1399 2716 1400
rect 2846 1404 2852 1405
rect 2846 1400 2847 1404
rect 2851 1400 2852 1404
rect 2846 1399 2852 1400
rect 2982 1404 2988 1405
rect 2982 1400 2983 1404
rect 2987 1400 2988 1404
rect 2982 1399 2988 1400
rect 3118 1404 3124 1405
rect 3118 1400 3119 1404
rect 3123 1400 3124 1404
rect 3118 1399 3124 1400
rect 3254 1404 3260 1405
rect 3254 1400 3255 1404
rect 3259 1400 3260 1404
rect 3798 1401 3799 1405
rect 3803 1401 3804 1405
rect 3798 1400 3804 1401
rect 3254 1399 3260 1400
rect 2138 1389 2144 1390
rect 1974 1388 1980 1389
rect 1974 1384 1975 1388
rect 1979 1384 1980 1388
rect 2138 1385 2139 1389
rect 2143 1385 2144 1389
rect 2138 1384 2144 1385
rect 2274 1389 2280 1390
rect 2274 1385 2275 1389
rect 2279 1385 2280 1389
rect 2274 1384 2280 1385
rect 2410 1389 2416 1390
rect 2410 1385 2411 1389
rect 2415 1385 2416 1389
rect 2410 1384 2416 1385
rect 2546 1389 2552 1390
rect 2546 1385 2547 1389
rect 2551 1385 2552 1389
rect 2546 1384 2552 1385
rect 2682 1389 2688 1390
rect 2682 1385 2683 1389
rect 2687 1385 2688 1389
rect 2682 1384 2688 1385
rect 2818 1389 2824 1390
rect 2818 1385 2819 1389
rect 2823 1385 2824 1389
rect 2818 1384 2824 1385
rect 2954 1389 2960 1390
rect 2954 1385 2955 1389
rect 2959 1385 2960 1389
rect 2954 1384 2960 1385
rect 3090 1389 3096 1390
rect 3090 1385 3091 1389
rect 3095 1385 3096 1389
rect 3090 1384 3096 1385
rect 3226 1389 3232 1390
rect 3226 1385 3227 1389
rect 3231 1385 3232 1389
rect 3226 1384 3232 1385
rect 3798 1388 3804 1389
rect 3798 1384 3799 1388
rect 3803 1384 3804 1388
rect 1974 1383 1980 1384
rect 3798 1383 3804 1384
rect 2258 1379 2269 1380
rect 255 1375 264 1376
rect 255 1371 256 1375
rect 263 1371 264 1375
rect 255 1370 264 1371
rect 386 1375 392 1376
rect 386 1371 387 1375
rect 391 1374 392 1375
rect 519 1375 525 1376
rect 519 1374 520 1375
rect 391 1372 520 1374
rect 391 1371 392 1372
rect 386 1370 392 1371
rect 519 1371 520 1372
rect 524 1371 525 1375
rect 519 1370 525 1371
rect 807 1375 816 1376
rect 807 1371 808 1375
rect 815 1371 816 1375
rect 807 1370 816 1371
rect 1095 1375 1104 1376
rect 1095 1371 1096 1375
rect 1103 1371 1104 1375
rect 1095 1370 1104 1371
rect 1383 1375 1389 1376
rect 1383 1371 1384 1375
rect 1388 1374 1389 1375
rect 1410 1375 1416 1376
rect 1410 1374 1411 1375
rect 1388 1372 1411 1374
rect 1388 1371 1389 1372
rect 1383 1370 1389 1371
rect 1410 1371 1411 1372
rect 1415 1371 1416 1375
rect 2258 1375 2259 1379
rect 2263 1375 2264 1379
rect 2268 1375 2269 1379
rect 2258 1374 2269 1375
rect 2271 1379 2277 1380
rect 2271 1375 2272 1379
rect 2276 1378 2277 1379
rect 2399 1379 2405 1380
rect 2399 1378 2400 1379
rect 2276 1376 2400 1378
rect 2276 1375 2277 1376
rect 2271 1374 2277 1375
rect 2399 1375 2400 1376
rect 2404 1375 2405 1379
rect 2399 1374 2405 1375
rect 2418 1379 2424 1380
rect 2418 1375 2419 1379
rect 2423 1378 2424 1379
rect 2535 1379 2541 1380
rect 2535 1378 2536 1379
rect 2423 1376 2536 1378
rect 2423 1375 2424 1376
rect 2418 1374 2424 1375
rect 2535 1375 2536 1376
rect 2540 1375 2541 1379
rect 2535 1374 2541 1375
rect 2671 1379 2677 1380
rect 2671 1375 2672 1379
rect 2676 1378 2677 1379
rect 2698 1379 2704 1380
rect 2698 1378 2699 1379
rect 2676 1376 2699 1378
rect 2676 1375 2677 1376
rect 2671 1374 2677 1375
rect 2698 1375 2699 1376
rect 2703 1375 2704 1379
rect 2698 1374 2704 1375
rect 2807 1379 2813 1380
rect 2807 1375 2808 1379
rect 2812 1378 2813 1379
rect 2834 1379 2840 1380
rect 2834 1378 2835 1379
rect 2812 1376 2835 1378
rect 2812 1375 2813 1376
rect 2807 1374 2813 1375
rect 2834 1375 2835 1376
rect 2839 1375 2840 1379
rect 2834 1374 2840 1375
rect 2943 1379 2949 1380
rect 2943 1375 2944 1379
rect 2948 1378 2949 1379
rect 2970 1379 2976 1380
rect 2970 1378 2971 1379
rect 2948 1376 2971 1378
rect 2948 1375 2949 1376
rect 2943 1374 2949 1375
rect 2970 1375 2971 1376
rect 2975 1375 2976 1379
rect 2970 1374 2976 1375
rect 3079 1379 3085 1380
rect 3079 1375 3080 1379
rect 3084 1378 3085 1379
rect 3106 1379 3112 1380
rect 3106 1378 3107 1379
rect 3084 1376 3107 1378
rect 3084 1375 3085 1376
rect 3079 1374 3085 1375
rect 3106 1375 3107 1376
rect 3111 1375 3112 1379
rect 3106 1374 3112 1375
rect 3215 1379 3221 1380
rect 3215 1375 3216 1379
rect 3220 1378 3221 1379
rect 3242 1379 3248 1380
rect 3242 1378 3243 1379
rect 3220 1376 3243 1378
rect 3220 1375 3221 1376
rect 3215 1374 3221 1375
rect 3242 1375 3243 1376
rect 3247 1375 3248 1379
rect 3242 1374 3248 1375
rect 3351 1379 3360 1380
rect 3351 1375 3352 1379
rect 3359 1375 3360 1379
rect 4943 1379 4949 1380
rect 4943 1378 4944 1379
rect 4901 1376 4944 1378
rect 3351 1374 3360 1375
rect 4943 1375 4944 1376
rect 4948 1375 4949 1379
rect 5079 1379 5085 1380
rect 5079 1378 5080 1379
rect 5037 1376 5080 1378
rect 4943 1374 4949 1375
rect 5079 1375 5080 1376
rect 5084 1375 5085 1379
rect 5215 1379 5221 1380
rect 5215 1378 5216 1379
rect 5173 1376 5216 1378
rect 5079 1374 5085 1375
rect 5215 1375 5216 1376
rect 5220 1375 5221 1379
rect 5471 1379 5477 1380
rect 5471 1378 5472 1379
rect 5445 1376 5472 1378
rect 5215 1374 5221 1375
rect 5306 1375 5312 1376
rect 1410 1370 1416 1371
rect 5306 1371 5307 1375
rect 5311 1371 5312 1375
rect 5471 1375 5472 1376
rect 5476 1375 5477 1379
rect 5471 1374 5477 1375
rect 5482 1379 5488 1380
rect 5482 1375 5483 1379
rect 5487 1378 5488 1379
rect 5487 1376 5509 1378
rect 5487 1375 5488 1376
rect 5482 1374 5488 1375
rect 5306 1370 5312 1371
rect 110 1368 116 1369
rect 1934 1368 1940 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 130 1367 136 1368
rect 130 1363 131 1367
rect 135 1363 136 1367
rect 130 1362 136 1363
rect 394 1367 400 1368
rect 394 1363 395 1367
rect 399 1363 400 1367
rect 394 1362 400 1363
rect 682 1367 688 1368
rect 682 1363 683 1367
rect 687 1363 688 1367
rect 682 1362 688 1363
rect 970 1367 976 1368
rect 970 1363 971 1367
rect 975 1363 976 1367
rect 970 1362 976 1363
rect 1258 1367 1264 1368
rect 1258 1363 1259 1367
rect 1263 1363 1264 1367
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 1934 1363 1940 1364
rect 1258 1362 1264 1363
rect 158 1352 164 1353
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 158 1348 159 1352
rect 163 1348 164 1352
rect 158 1347 164 1348
rect 422 1352 428 1353
rect 422 1348 423 1352
rect 427 1348 428 1352
rect 422 1347 428 1348
rect 710 1352 716 1353
rect 710 1348 711 1352
rect 715 1348 716 1352
rect 710 1347 716 1348
rect 998 1352 1004 1353
rect 998 1348 999 1352
rect 1003 1348 1004 1352
rect 998 1347 1004 1348
rect 1286 1352 1292 1353
rect 1286 1348 1287 1352
rect 1291 1348 1292 1352
rect 1286 1347 1292 1348
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 110 1346 116 1347
rect 1934 1346 1940 1347
rect 2271 1347 2277 1348
rect 2271 1346 2272 1347
rect 2229 1344 2272 1346
rect 2271 1343 2272 1344
rect 2276 1343 2277 1347
rect 2418 1347 2424 1348
rect 2418 1346 2419 1347
rect 2365 1344 2419 1346
rect 2271 1342 2277 1343
rect 2418 1343 2419 1344
rect 2423 1343 2424 1347
rect 2418 1342 2424 1343
rect 2498 1347 2504 1348
rect 2498 1343 2499 1347
rect 2503 1343 2504 1347
rect 2498 1342 2504 1343
rect 2634 1347 2640 1348
rect 2634 1343 2635 1347
rect 2639 1343 2640 1347
rect 2634 1342 2640 1343
rect 2698 1347 2704 1348
rect 2698 1343 2699 1347
rect 2703 1343 2704 1347
rect 2698 1342 2704 1343
rect 2834 1347 2840 1348
rect 2834 1343 2835 1347
rect 2839 1343 2840 1347
rect 2834 1342 2840 1343
rect 2970 1347 2976 1348
rect 2970 1343 2971 1347
rect 2975 1343 2976 1347
rect 2970 1342 2976 1343
rect 3106 1347 3112 1348
rect 3106 1343 3107 1347
rect 3111 1343 3112 1347
rect 3106 1342 3112 1343
rect 3242 1347 3248 1348
rect 3242 1343 3243 1347
rect 3247 1343 3248 1347
rect 3242 1342 3248 1343
rect 4934 1343 4941 1344
rect 4934 1339 4935 1343
rect 4940 1339 4941 1343
rect 4934 1338 4941 1339
rect 4943 1343 4949 1344
rect 4943 1339 4944 1343
rect 4948 1342 4949 1343
rect 5071 1343 5077 1344
rect 5071 1342 5072 1343
rect 4948 1340 5072 1342
rect 4948 1339 4949 1340
rect 4943 1338 4949 1339
rect 5071 1339 5072 1340
rect 5076 1339 5077 1343
rect 5071 1338 5077 1339
rect 5079 1343 5085 1344
rect 5079 1339 5080 1343
rect 5084 1342 5085 1343
rect 5207 1343 5213 1344
rect 5207 1342 5208 1343
rect 5084 1340 5208 1342
rect 5084 1339 5085 1340
rect 5079 1338 5085 1339
rect 5207 1339 5208 1340
rect 5212 1339 5213 1343
rect 5207 1338 5213 1339
rect 5215 1343 5221 1344
rect 5215 1339 5216 1343
rect 5220 1342 5221 1343
rect 5343 1343 5349 1344
rect 5343 1342 5344 1343
rect 5220 1340 5344 1342
rect 5220 1339 5221 1340
rect 5215 1338 5221 1339
rect 5343 1339 5344 1340
rect 5348 1339 5349 1343
rect 5343 1338 5349 1339
rect 5479 1343 5488 1344
rect 5479 1339 5480 1343
rect 5487 1339 5488 1343
rect 5479 1338 5488 1339
rect 5586 1343 5592 1344
rect 5586 1339 5587 1343
rect 5591 1342 5592 1343
rect 5615 1343 5621 1344
rect 5615 1342 5616 1343
rect 5591 1340 5616 1342
rect 5591 1339 5592 1340
rect 5586 1338 5592 1339
rect 5615 1339 5616 1340
rect 5620 1339 5621 1343
rect 5615 1338 5621 1339
rect 3838 1336 3844 1337
rect 5662 1336 5668 1337
rect 3838 1332 3839 1336
rect 3843 1332 3844 1336
rect 3838 1331 3844 1332
rect 4810 1335 4816 1336
rect 4810 1331 4811 1335
rect 4815 1331 4816 1335
rect 4810 1330 4816 1331
rect 4946 1335 4952 1336
rect 4946 1331 4947 1335
rect 4951 1331 4952 1335
rect 4946 1330 4952 1331
rect 5082 1335 5088 1336
rect 5082 1331 5083 1335
rect 5087 1331 5088 1335
rect 5082 1330 5088 1331
rect 5218 1335 5224 1336
rect 5218 1331 5219 1335
rect 5223 1331 5224 1335
rect 5218 1330 5224 1331
rect 5354 1335 5360 1336
rect 5354 1331 5355 1335
rect 5359 1331 5360 1335
rect 5354 1330 5360 1331
rect 5490 1335 5496 1336
rect 5490 1331 5491 1335
rect 5495 1331 5496 1335
rect 5662 1332 5663 1336
rect 5667 1332 5668 1336
rect 5662 1331 5668 1332
rect 5490 1330 5496 1331
rect 4838 1320 4844 1321
rect 3838 1319 3844 1320
rect 3838 1315 3839 1319
rect 3843 1315 3844 1319
rect 4838 1316 4839 1320
rect 4843 1316 4844 1320
rect 4838 1315 4844 1316
rect 4974 1320 4980 1321
rect 4974 1316 4975 1320
rect 4979 1316 4980 1320
rect 4974 1315 4980 1316
rect 5110 1320 5116 1321
rect 5110 1316 5111 1320
rect 5115 1316 5116 1320
rect 5110 1315 5116 1316
rect 5246 1320 5252 1321
rect 5246 1316 5247 1320
rect 5251 1316 5252 1320
rect 5246 1315 5252 1316
rect 5382 1320 5388 1321
rect 5382 1316 5383 1320
rect 5387 1316 5388 1320
rect 5382 1315 5388 1316
rect 5518 1320 5524 1321
rect 5518 1316 5519 1320
rect 5523 1316 5524 1320
rect 5518 1315 5524 1316
rect 5662 1319 5668 1320
rect 5662 1315 5663 1319
rect 5667 1315 5668 1319
rect 3838 1314 3844 1315
rect 5662 1314 5668 1315
rect 2246 1299 2252 1300
rect 2246 1298 2247 1299
rect 2221 1296 2247 1298
rect 2246 1295 2247 1296
rect 2251 1295 2252 1299
rect 2246 1294 2252 1295
rect 2258 1299 2264 1300
rect 2258 1295 2259 1299
rect 2263 1298 2264 1299
rect 2399 1299 2405 1300
rect 2263 1296 2285 1298
rect 2263 1295 2264 1296
rect 2258 1294 2264 1295
rect 2399 1295 2400 1299
rect 2404 1298 2405 1299
rect 2530 1299 2536 1300
rect 2404 1296 2421 1298
rect 2404 1295 2405 1296
rect 2399 1294 2405 1295
rect 2530 1295 2531 1299
rect 2535 1298 2536 1299
rect 2706 1299 2712 1300
rect 2535 1296 2573 1298
rect 2535 1295 2536 1296
rect 2530 1294 2536 1295
rect 2706 1295 2707 1299
rect 2711 1298 2712 1299
rect 3023 1299 3029 1300
rect 3023 1298 3024 1299
rect 2711 1296 2733 1298
rect 2981 1296 3024 1298
rect 2711 1295 2712 1296
rect 2706 1294 2712 1295
rect 3023 1295 3024 1296
rect 3028 1295 3029 1299
rect 3263 1299 3269 1300
rect 3263 1298 3264 1299
rect 3165 1296 3264 1298
rect 3023 1294 3029 1295
rect 3263 1295 3264 1296
rect 3268 1295 3269 1299
rect 3594 1299 3600 1300
rect 3263 1294 3269 1295
rect 3354 1295 3360 1296
rect 110 1293 116 1294
rect 1934 1293 1940 1294
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 158 1292 164 1293
rect 158 1288 159 1292
rect 163 1288 164 1292
rect 158 1287 164 1288
rect 454 1292 460 1293
rect 454 1288 455 1292
rect 459 1288 460 1292
rect 454 1287 460 1288
rect 774 1292 780 1293
rect 774 1288 775 1292
rect 779 1288 780 1292
rect 774 1287 780 1288
rect 1094 1292 1100 1293
rect 1094 1288 1095 1292
rect 1099 1288 1100 1292
rect 1094 1287 1100 1288
rect 1422 1292 1428 1293
rect 1422 1288 1423 1292
rect 1427 1288 1428 1292
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 3354 1291 3355 1295
rect 3359 1291 3360 1295
rect 3354 1290 3360 1291
rect 3554 1295 3560 1296
rect 3554 1291 3555 1295
rect 3559 1291 3560 1295
rect 3594 1295 3595 1299
rect 3599 1298 3600 1299
rect 3599 1296 3669 1298
rect 3599 1295 3600 1296
rect 3594 1294 3600 1295
rect 3554 1290 3560 1291
rect 1934 1288 1940 1289
rect 1422 1287 1428 1288
rect 130 1277 136 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 130 1273 131 1277
rect 135 1273 136 1277
rect 130 1272 136 1273
rect 426 1277 432 1278
rect 426 1273 427 1277
rect 431 1273 432 1277
rect 426 1272 432 1273
rect 746 1277 752 1278
rect 746 1273 747 1277
rect 751 1273 752 1277
rect 746 1272 752 1273
rect 1066 1277 1072 1278
rect 1066 1273 1067 1277
rect 1071 1273 1072 1277
rect 1066 1272 1072 1273
rect 1394 1277 1400 1278
rect 1394 1273 1395 1277
rect 1399 1273 1400 1277
rect 1394 1272 1400 1273
rect 1934 1276 1940 1277
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 110 1271 116 1272
rect 1934 1271 1940 1272
rect 218 1267 224 1268
rect 218 1263 219 1267
rect 223 1266 224 1267
rect 255 1267 261 1268
rect 255 1266 256 1267
rect 223 1264 256 1266
rect 223 1263 224 1264
rect 218 1262 224 1263
rect 255 1263 256 1264
rect 260 1263 261 1267
rect 255 1262 261 1263
rect 298 1267 304 1268
rect 298 1263 299 1267
rect 303 1266 304 1267
rect 551 1267 557 1268
rect 551 1266 552 1267
rect 303 1264 552 1266
rect 303 1263 304 1264
rect 298 1262 304 1263
rect 551 1263 552 1264
rect 556 1263 557 1267
rect 551 1262 557 1263
rect 871 1267 877 1268
rect 871 1263 872 1267
rect 876 1266 877 1267
rect 1082 1267 1088 1268
rect 1082 1266 1083 1267
rect 876 1264 1083 1266
rect 876 1263 877 1264
rect 871 1262 877 1263
rect 1082 1263 1083 1264
rect 1087 1263 1088 1267
rect 1082 1262 1088 1263
rect 1191 1267 1197 1268
rect 1191 1263 1192 1267
rect 1196 1266 1197 1267
rect 1199 1267 1205 1268
rect 1199 1266 1200 1267
rect 1196 1264 1200 1266
rect 1196 1263 1197 1264
rect 1191 1262 1197 1263
rect 1199 1263 1200 1264
rect 1204 1263 1205 1267
rect 1519 1267 1525 1268
rect 1519 1266 1520 1267
rect 1199 1262 1205 1263
rect 1459 1264 1520 1266
rect 834 1259 840 1260
rect 834 1255 835 1259
rect 839 1258 840 1259
rect 1459 1258 1461 1264
rect 1519 1263 1520 1264
rect 1524 1263 1525 1267
rect 1519 1262 1525 1263
rect 2255 1263 2264 1264
rect 2255 1259 2256 1263
rect 2263 1259 2264 1263
rect 2255 1258 2264 1259
rect 2391 1263 2397 1264
rect 2391 1259 2392 1263
rect 2396 1262 2397 1263
rect 2399 1263 2405 1264
rect 2399 1262 2400 1263
rect 2396 1260 2400 1262
rect 2396 1259 2397 1260
rect 2391 1258 2397 1259
rect 2399 1259 2400 1260
rect 2404 1259 2405 1263
rect 2399 1258 2405 1259
rect 2527 1263 2536 1264
rect 2527 1259 2528 1263
rect 2535 1259 2536 1263
rect 2527 1258 2536 1259
rect 2679 1263 2685 1264
rect 2679 1259 2680 1263
rect 2684 1262 2685 1263
rect 2706 1263 2712 1264
rect 2706 1262 2707 1263
rect 2684 1260 2707 1262
rect 2684 1259 2685 1260
rect 2679 1258 2685 1259
rect 2706 1259 2707 1260
rect 2711 1259 2712 1263
rect 2706 1258 2712 1259
rect 2722 1263 2728 1264
rect 2722 1259 2723 1263
rect 2727 1262 2728 1263
rect 2839 1263 2845 1264
rect 2839 1262 2840 1263
rect 2727 1260 2840 1262
rect 2727 1259 2728 1260
rect 2722 1258 2728 1259
rect 2839 1259 2840 1260
rect 2844 1259 2845 1263
rect 2839 1258 2845 1259
rect 3014 1263 3021 1264
rect 3014 1259 3015 1263
rect 3020 1259 3021 1263
rect 3014 1258 3021 1259
rect 3023 1263 3029 1264
rect 3023 1259 3024 1263
rect 3028 1262 3029 1263
rect 3199 1263 3205 1264
rect 3199 1262 3200 1263
rect 3028 1260 3200 1262
rect 3028 1259 3029 1260
rect 3023 1258 3029 1259
rect 3199 1259 3200 1260
rect 3204 1259 3205 1263
rect 3199 1258 3205 1259
rect 3263 1263 3269 1264
rect 3263 1259 3264 1263
rect 3268 1262 3269 1263
rect 3391 1263 3397 1264
rect 3391 1262 3392 1263
rect 3268 1260 3392 1262
rect 3268 1259 3269 1260
rect 3263 1258 3269 1259
rect 3391 1259 3392 1260
rect 3396 1259 3397 1263
rect 3391 1258 3397 1259
rect 3591 1263 3600 1264
rect 3591 1259 3592 1263
rect 3599 1259 3600 1263
rect 3591 1258 3600 1259
rect 3738 1263 3744 1264
rect 3738 1259 3739 1263
rect 3743 1262 3744 1263
rect 3775 1263 3781 1264
rect 3775 1262 3776 1263
rect 3743 1260 3776 1262
rect 3743 1259 3744 1260
rect 3738 1258 3744 1259
rect 3775 1259 3776 1260
rect 3780 1259 3781 1263
rect 3775 1258 3781 1259
rect 839 1256 1461 1258
rect 3838 1257 3844 1258
rect 5662 1257 5668 1258
rect 1974 1256 1980 1257
rect 3798 1256 3804 1257
rect 839 1255 840 1256
rect 834 1254 840 1255
rect 1974 1252 1975 1256
rect 1979 1252 1980 1256
rect 1974 1251 1980 1252
rect 2130 1255 2136 1256
rect 2130 1251 2131 1255
rect 2135 1251 2136 1255
rect 2130 1250 2136 1251
rect 2266 1255 2272 1256
rect 2266 1251 2267 1255
rect 2271 1251 2272 1255
rect 2266 1250 2272 1251
rect 2402 1255 2408 1256
rect 2402 1251 2403 1255
rect 2407 1251 2408 1255
rect 2402 1250 2408 1251
rect 2554 1255 2560 1256
rect 2554 1251 2555 1255
rect 2559 1251 2560 1255
rect 2554 1250 2560 1251
rect 2714 1255 2720 1256
rect 2714 1251 2715 1255
rect 2719 1251 2720 1255
rect 2714 1250 2720 1251
rect 2890 1255 2896 1256
rect 2890 1251 2891 1255
rect 2895 1251 2896 1255
rect 2890 1250 2896 1251
rect 3074 1255 3080 1256
rect 3074 1251 3075 1255
rect 3079 1251 3080 1255
rect 3074 1250 3080 1251
rect 3266 1255 3272 1256
rect 3266 1251 3267 1255
rect 3271 1251 3272 1255
rect 3266 1250 3272 1251
rect 3466 1255 3472 1256
rect 3466 1251 3467 1255
rect 3471 1251 3472 1255
rect 3466 1250 3472 1251
rect 3650 1255 3656 1256
rect 3650 1251 3651 1255
rect 3655 1251 3656 1255
rect 3798 1252 3799 1256
rect 3803 1252 3804 1256
rect 3838 1253 3839 1257
rect 3843 1253 3844 1257
rect 3838 1252 3844 1253
rect 4734 1256 4740 1257
rect 4734 1252 4735 1256
rect 4739 1252 4740 1256
rect 3798 1251 3804 1252
rect 4734 1251 4740 1252
rect 4878 1256 4884 1257
rect 4878 1252 4879 1256
rect 4883 1252 4884 1256
rect 4878 1251 4884 1252
rect 5030 1256 5036 1257
rect 5030 1252 5031 1256
rect 5035 1252 5036 1256
rect 5030 1251 5036 1252
rect 5190 1256 5196 1257
rect 5190 1252 5191 1256
rect 5195 1252 5196 1256
rect 5190 1251 5196 1252
rect 5358 1256 5364 1257
rect 5358 1252 5359 1256
rect 5363 1252 5364 1256
rect 5358 1251 5364 1252
rect 5526 1256 5532 1257
rect 5526 1252 5527 1256
rect 5531 1252 5532 1256
rect 5662 1253 5663 1257
rect 5667 1253 5668 1257
rect 5662 1252 5668 1253
rect 5526 1251 5532 1252
rect 3650 1250 3656 1251
rect 4706 1241 4712 1242
rect 2158 1240 2164 1241
rect 1974 1239 1980 1240
rect 298 1235 304 1236
rect 298 1234 299 1235
rect 221 1232 299 1234
rect 298 1231 299 1232
rect 303 1231 304 1235
rect 298 1230 304 1231
rect 514 1235 520 1236
rect 514 1231 515 1235
rect 519 1231 520 1235
rect 514 1230 520 1231
rect 834 1235 840 1236
rect 834 1231 835 1235
rect 839 1231 840 1235
rect 834 1230 840 1231
rect 1082 1235 1088 1236
rect 1082 1231 1083 1235
rect 1087 1231 1088 1235
rect 1082 1230 1088 1231
rect 1410 1235 1416 1236
rect 1410 1231 1411 1235
rect 1415 1231 1416 1235
rect 1974 1235 1975 1239
rect 1979 1235 1980 1239
rect 2158 1236 2159 1240
rect 2163 1236 2164 1240
rect 2158 1235 2164 1236
rect 2294 1240 2300 1241
rect 2294 1236 2295 1240
rect 2299 1236 2300 1240
rect 2294 1235 2300 1236
rect 2430 1240 2436 1241
rect 2430 1236 2431 1240
rect 2435 1236 2436 1240
rect 2430 1235 2436 1236
rect 2582 1240 2588 1241
rect 2582 1236 2583 1240
rect 2587 1236 2588 1240
rect 2582 1235 2588 1236
rect 2742 1240 2748 1241
rect 2742 1236 2743 1240
rect 2747 1236 2748 1240
rect 2742 1235 2748 1236
rect 2918 1240 2924 1241
rect 2918 1236 2919 1240
rect 2923 1236 2924 1240
rect 2918 1235 2924 1236
rect 3102 1240 3108 1241
rect 3102 1236 3103 1240
rect 3107 1236 3108 1240
rect 3102 1235 3108 1236
rect 3294 1240 3300 1241
rect 3294 1236 3295 1240
rect 3299 1236 3300 1240
rect 3294 1235 3300 1236
rect 3494 1240 3500 1241
rect 3494 1236 3495 1240
rect 3499 1236 3500 1240
rect 3494 1235 3500 1236
rect 3678 1240 3684 1241
rect 3838 1240 3844 1241
rect 3678 1236 3679 1240
rect 3683 1236 3684 1240
rect 3678 1235 3684 1236
rect 3798 1239 3804 1240
rect 3798 1235 3799 1239
rect 3803 1235 3804 1239
rect 3838 1236 3839 1240
rect 3843 1236 3844 1240
rect 4706 1237 4707 1241
rect 4711 1237 4712 1241
rect 4706 1236 4712 1237
rect 4850 1241 4856 1242
rect 4850 1237 4851 1241
rect 4855 1237 4856 1241
rect 4850 1236 4856 1237
rect 5002 1241 5008 1242
rect 5002 1237 5003 1241
rect 5007 1237 5008 1241
rect 5002 1236 5008 1237
rect 5162 1241 5168 1242
rect 5162 1237 5163 1241
rect 5167 1237 5168 1241
rect 5162 1236 5168 1237
rect 5330 1241 5336 1242
rect 5330 1237 5331 1241
rect 5335 1237 5336 1241
rect 5330 1236 5336 1237
rect 5498 1241 5504 1242
rect 5498 1237 5499 1241
rect 5503 1237 5504 1241
rect 5498 1236 5504 1237
rect 5662 1240 5668 1241
rect 5662 1236 5663 1240
rect 5667 1236 5668 1240
rect 3838 1235 3844 1236
rect 5662 1235 5668 1236
rect 1974 1234 1980 1235
rect 3798 1234 3804 1235
rect 1410 1230 1416 1231
rect 4831 1231 4837 1232
rect 4831 1227 4832 1231
rect 4836 1230 4837 1231
rect 4858 1231 4864 1232
rect 4858 1230 4859 1231
rect 4836 1228 4859 1230
rect 4836 1227 4837 1228
rect 4831 1226 4837 1227
rect 4858 1227 4859 1228
rect 4863 1227 4864 1231
rect 4858 1226 4864 1227
rect 4975 1231 4981 1232
rect 4975 1227 4976 1231
rect 4980 1230 4981 1231
rect 5018 1231 5024 1232
rect 5018 1230 5019 1231
rect 4980 1228 5019 1230
rect 4980 1227 4981 1228
rect 4975 1226 4981 1227
rect 5018 1227 5019 1228
rect 5023 1227 5024 1231
rect 5127 1231 5133 1232
rect 5127 1230 5128 1231
rect 5018 1226 5024 1227
rect 5028 1228 5128 1230
rect 4794 1223 4800 1224
rect 4794 1219 4795 1223
rect 4799 1222 4800 1223
rect 5028 1222 5030 1228
rect 5127 1227 5128 1228
rect 5132 1227 5133 1231
rect 5127 1226 5133 1227
rect 5287 1231 5293 1232
rect 5287 1227 5288 1231
rect 5292 1230 5293 1231
rect 5306 1231 5312 1232
rect 5306 1230 5307 1231
rect 5292 1228 5307 1230
rect 5292 1227 5293 1228
rect 5287 1226 5293 1227
rect 5306 1227 5307 1228
rect 5311 1227 5312 1231
rect 5306 1226 5312 1227
rect 5318 1231 5324 1232
rect 5318 1227 5319 1231
rect 5323 1230 5324 1231
rect 5455 1231 5461 1232
rect 5455 1230 5456 1231
rect 5323 1228 5456 1230
rect 5323 1227 5324 1228
rect 5318 1226 5324 1227
rect 5455 1227 5456 1228
rect 5460 1227 5461 1231
rect 5455 1226 5461 1227
rect 5618 1231 5629 1232
rect 5618 1227 5619 1231
rect 5623 1227 5624 1231
rect 5628 1227 5629 1231
rect 5618 1226 5629 1227
rect 4799 1220 5030 1222
rect 4799 1219 4800 1220
rect 4794 1218 4800 1219
rect 2246 1215 2252 1216
rect 2246 1211 2247 1215
rect 2251 1211 2252 1215
rect 2246 1210 2252 1211
rect 2248 1208 2814 1210
rect 2810 1207 2816 1208
rect 2810 1203 2811 1207
rect 2815 1203 2816 1207
rect 2810 1202 2816 1203
rect 4794 1199 4800 1200
rect 4794 1195 4795 1199
rect 4799 1195 4800 1199
rect 4794 1194 4800 1195
rect 4934 1199 4940 1200
rect 4934 1195 4935 1199
rect 4939 1195 4940 1199
rect 4934 1194 4940 1195
rect 5018 1199 5024 1200
rect 5018 1195 5019 1199
rect 5023 1195 5024 1199
rect 5318 1199 5324 1200
rect 5318 1198 5319 1199
rect 5253 1196 5319 1198
rect 5018 1194 5024 1195
rect 5318 1195 5319 1196
rect 5323 1195 5324 1199
rect 5318 1194 5324 1195
rect 5406 1199 5412 1200
rect 5406 1195 5407 1199
rect 5411 1195 5412 1199
rect 5406 1194 5412 1195
rect 5586 1199 5592 1200
rect 5586 1195 5587 1199
rect 5591 1195 5592 1199
rect 5586 1194 5592 1195
rect 1974 1181 1980 1182
rect 3798 1181 3804 1182
rect 1974 1177 1975 1181
rect 1979 1177 1980 1181
rect 1974 1176 1980 1177
rect 2022 1180 2028 1181
rect 2022 1176 2023 1180
rect 2027 1176 2028 1180
rect 2022 1175 2028 1176
rect 2238 1180 2244 1181
rect 2238 1176 2239 1180
rect 2243 1176 2244 1180
rect 2238 1175 2244 1176
rect 2478 1180 2484 1181
rect 2478 1176 2479 1180
rect 2483 1176 2484 1180
rect 2478 1175 2484 1176
rect 2718 1180 2724 1181
rect 2718 1176 2719 1180
rect 2723 1176 2724 1180
rect 2718 1175 2724 1176
rect 2958 1180 2964 1181
rect 2958 1176 2959 1180
rect 2963 1176 2964 1180
rect 2958 1175 2964 1176
rect 3206 1180 3212 1181
rect 3206 1176 3207 1180
rect 3211 1176 3212 1180
rect 3206 1175 3212 1176
rect 3454 1180 3460 1181
rect 3454 1176 3455 1180
rect 3459 1176 3460 1180
rect 3454 1175 3460 1176
rect 3678 1180 3684 1181
rect 3678 1176 3679 1180
rect 3683 1176 3684 1180
rect 3798 1177 3799 1181
rect 3803 1177 3804 1181
rect 3798 1176 3804 1177
rect 3678 1175 3684 1176
rect 1994 1165 2000 1166
rect 1974 1164 1980 1165
rect 258 1163 264 1164
rect 258 1159 259 1163
rect 263 1162 264 1163
rect 458 1163 464 1164
rect 263 1160 349 1162
rect 263 1159 264 1160
rect 258 1158 264 1159
rect 458 1159 459 1163
rect 463 1162 464 1163
rect 991 1163 997 1164
rect 991 1162 992 1163
rect 463 1160 581 1162
rect 893 1160 992 1162
rect 463 1159 464 1160
rect 458 1158 464 1159
rect 991 1159 992 1160
rect 996 1159 997 1163
rect 1191 1163 1197 1164
rect 1191 1162 1192 1163
rect 1133 1160 1192 1162
rect 991 1158 997 1159
rect 1191 1159 1192 1160
rect 1196 1159 1197 1163
rect 1191 1158 1197 1159
rect 1199 1163 1205 1164
rect 1199 1159 1200 1163
rect 1204 1162 1205 1163
rect 1650 1163 1656 1164
rect 1204 1160 1301 1162
rect 1204 1159 1205 1160
rect 1199 1158 1205 1159
rect 1650 1159 1651 1163
rect 1655 1162 1656 1163
rect 1655 1160 1789 1162
rect 1974 1160 1975 1164
rect 1979 1160 1980 1164
rect 1994 1161 1995 1165
rect 1999 1161 2000 1165
rect 1994 1160 2000 1161
rect 2210 1165 2216 1166
rect 2210 1161 2211 1165
rect 2215 1161 2216 1165
rect 2210 1160 2216 1161
rect 2450 1165 2456 1166
rect 2450 1161 2451 1165
rect 2455 1161 2456 1165
rect 2450 1160 2456 1161
rect 2690 1165 2696 1166
rect 2690 1161 2691 1165
rect 2695 1161 2696 1165
rect 2690 1160 2696 1161
rect 2930 1165 2936 1166
rect 2930 1161 2931 1165
rect 2935 1161 2936 1165
rect 2930 1160 2936 1161
rect 3178 1165 3184 1166
rect 3178 1161 3179 1165
rect 3183 1161 3184 1165
rect 3178 1160 3184 1161
rect 3426 1165 3432 1166
rect 3426 1161 3427 1165
rect 3431 1161 3432 1165
rect 3426 1160 3432 1161
rect 3650 1165 3656 1166
rect 3650 1161 3651 1165
rect 3655 1161 3656 1165
rect 3650 1160 3656 1161
rect 3798 1164 3804 1165
rect 3798 1160 3799 1164
rect 3803 1160 3804 1164
rect 1655 1159 1656 1160
rect 1974 1159 1980 1160
rect 3798 1159 3804 1160
rect 1650 1158 1656 1159
rect 216 1154 218 1157
rect 270 1155 276 1156
rect 270 1154 271 1155
rect 216 1152 271 1154
rect 270 1151 271 1152
rect 275 1151 276 1155
rect 1608 1154 1610 1157
rect 1758 1155 1764 1156
rect 1758 1154 1759 1155
rect 1608 1152 1759 1154
rect 270 1150 276 1151
rect 1758 1151 1759 1152
rect 1763 1151 1764 1155
rect 1758 1150 1764 1151
rect 2119 1155 2125 1156
rect 2119 1151 2120 1155
rect 2124 1154 2125 1155
rect 2226 1155 2232 1156
rect 2226 1154 2227 1155
rect 2124 1152 2227 1154
rect 2124 1151 2125 1152
rect 2119 1150 2125 1151
rect 2226 1151 2227 1152
rect 2231 1151 2232 1155
rect 2226 1150 2232 1151
rect 2335 1155 2341 1156
rect 2335 1151 2336 1155
rect 2340 1154 2341 1155
rect 2466 1155 2472 1156
rect 2466 1154 2467 1155
rect 2340 1152 2467 1154
rect 2340 1151 2341 1152
rect 2335 1150 2341 1151
rect 2466 1151 2467 1152
rect 2471 1151 2472 1155
rect 2466 1150 2472 1151
rect 2575 1155 2581 1156
rect 2575 1151 2576 1155
rect 2580 1154 2581 1155
rect 2706 1155 2712 1156
rect 2706 1154 2707 1155
rect 2580 1152 2707 1154
rect 2580 1151 2581 1152
rect 2575 1150 2581 1151
rect 2706 1151 2707 1152
rect 2711 1151 2712 1155
rect 2706 1150 2712 1151
rect 2810 1155 2821 1156
rect 2810 1151 2811 1155
rect 2815 1151 2816 1155
rect 2820 1151 2821 1155
rect 2810 1150 2821 1151
rect 3055 1155 3061 1156
rect 3055 1151 3056 1155
rect 3060 1154 3061 1155
rect 3082 1155 3088 1156
rect 3082 1154 3083 1155
rect 3060 1152 3083 1154
rect 3060 1151 3061 1152
rect 3055 1150 3061 1151
rect 3082 1151 3083 1152
rect 3087 1151 3088 1155
rect 3082 1150 3088 1151
rect 3303 1155 3309 1156
rect 3303 1151 3304 1155
rect 3308 1154 3309 1155
rect 3442 1155 3448 1156
rect 3442 1154 3443 1155
rect 3308 1152 3443 1154
rect 3308 1151 3309 1152
rect 3303 1150 3309 1151
rect 3442 1151 3443 1152
rect 3447 1151 3448 1155
rect 3442 1150 3448 1151
rect 3551 1155 3560 1156
rect 3551 1151 3552 1155
rect 3559 1151 3560 1155
rect 3551 1150 3560 1151
rect 3775 1155 3781 1156
rect 3775 1151 3776 1155
rect 3780 1154 3781 1155
rect 3780 1152 3830 1154
rect 3780 1151 3781 1152
rect 3775 1150 3781 1151
rect 3828 1142 3830 1152
rect 4034 1143 4040 1144
rect 3828 1140 3877 1142
rect 4034 1139 4035 1143
rect 4039 1142 4040 1143
rect 4426 1143 4432 1144
rect 4039 1140 4085 1142
rect 4039 1139 4040 1140
rect 4034 1138 4040 1139
rect 4386 1139 4392 1140
rect 4386 1135 4387 1139
rect 4391 1135 4392 1139
rect 4426 1139 4427 1143
rect 4431 1142 4432 1143
rect 4906 1143 4912 1144
rect 4431 1140 4557 1142
rect 4431 1139 4432 1140
rect 4426 1138 4432 1139
rect 4866 1139 4872 1140
rect 4386 1134 4392 1135
rect 4866 1135 4867 1139
rect 4871 1135 4872 1139
rect 4906 1139 4907 1143
rect 4911 1142 4912 1143
rect 5618 1143 5624 1144
rect 5618 1142 5619 1143
rect 4911 1140 5045 1142
rect 5605 1140 5619 1142
rect 4911 1139 4912 1140
rect 4906 1138 4912 1139
rect 5370 1139 5376 1140
rect 4866 1134 4872 1135
rect 5370 1135 5371 1139
rect 5375 1135 5376 1139
rect 5618 1139 5619 1140
rect 5623 1139 5624 1143
rect 5618 1138 5624 1139
rect 5370 1134 5376 1135
rect 255 1127 264 1128
rect 255 1123 256 1127
rect 263 1123 264 1127
rect 255 1122 264 1123
rect 455 1127 464 1128
rect 455 1123 456 1127
rect 463 1123 464 1127
rect 455 1122 464 1123
rect 514 1127 520 1128
rect 514 1123 515 1127
rect 519 1126 520 1127
rect 687 1127 693 1128
rect 687 1126 688 1127
rect 519 1124 688 1126
rect 519 1123 520 1124
rect 514 1122 520 1123
rect 687 1123 688 1124
rect 692 1123 693 1127
rect 687 1122 693 1123
rect 927 1127 933 1128
rect 927 1123 928 1127
rect 932 1126 933 1127
rect 938 1127 944 1128
rect 938 1126 939 1127
rect 932 1124 939 1126
rect 932 1123 933 1124
rect 927 1122 933 1123
rect 938 1123 939 1124
rect 943 1123 944 1127
rect 938 1122 944 1123
rect 991 1127 997 1128
rect 991 1123 992 1127
rect 996 1126 997 1127
rect 1167 1127 1173 1128
rect 1167 1126 1168 1127
rect 996 1124 1168 1126
rect 996 1123 997 1124
rect 991 1122 997 1123
rect 1167 1123 1168 1124
rect 1172 1123 1173 1127
rect 1167 1122 1173 1123
rect 1191 1127 1197 1128
rect 1191 1123 1192 1127
rect 1196 1126 1197 1127
rect 1407 1127 1413 1128
rect 1407 1126 1408 1127
rect 1196 1124 1408 1126
rect 1196 1123 1197 1124
rect 1191 1122 1197 1123
rect 1407 1123 1408 1124
rect 1412 1123 1413 1127
rect 1407 1122 1413 1123
rect 1647 1127 1656 1128
rect 1647 1123 1648 1127
rect 1655 1123 1656 1127
rect 1647 1122 1656 1123
rect 1895 1127 1901 1128
rect 1895 1123 1896 1127
rect 1900 1126 1901 1127
rect 1900 1124 1958 1126
rect 1900 1123 1901 1124
rect 1895 1122 1901 1123
rect 1956 1122 1958 1124
rect 2226 1123 2232 1124
rect 110 1120 116 1121
rect 1934 1120 1940 1121
rect 1956 1120 2013 1122
rect 110 1116 111 1120
rect 115 1116 116 1120
rect 110 1115 116 1116
rect 130 1119 136 1120
rect 130 1115 131 1119
rect 135 1115 136 1119
rect 130 1114 136 1115
rect 330 1119 336 1120
rect 330 1115 331 1119
rect 335 1115 336 1119
rect 330 1114 336 1115
rect 562 1119 568 1120
rect 562 1115 563 1119
rect 567 1115 568 1119
rect 562 1114 568 1115
rect 802 1119 808 1120
rect 802 1115 803 1119
rect 807 1115 808 1119
rect 802 1114 808 1115
rect 1042 1119 1048 1120
rect 1042 1115 1043 1119
rect 1047 1115 1048 1119
rect 1042 1114 1048 1115
rect 1282 1119 1288 1120
rect 1282 1115 1283 1119
rect 1287 1115 1288 1119
rect 1282 1114 1288 1115
rect 1522 1119 1528 1120
rect 1522 1115 1523 1119
rect 1527 1115 1528 1119
rect 1522 1114 1528 1115
rect 1770 1119 1776 1120
rect 1770 1115 1771 1119
rect 1775 1115 1776 1119
rect 1934 1116 1935 1120
rect 1939 1116 1940 1120
rect 2226 1119 2227 1123
rect 2231 1119 2232 1123
rect 2226 1118 2232 1119
rect 2466 1123 2472 1124
rect 2466 1119 2467 1123
rect 2471 1119 2472 1123
rect 2466 1118 2472 1119
rect 2706 1123 2712 1124
rect 2706 1119 2707 1123
rect 2711 1119 2712 1123
rect 2706 1118 2712 1119
rect 3014 1123 3020 1124
rect 3014 1119 3015 1123
rect 3019 1119 3020 1123
rect 3378 1123 3384 1124
rect 3378 1122 3379 1123
rect 3269 1120 3379 1122
rect 3014 1118 3020 1119
rect 3378 1119 3379 1120
rect 3383 1119 3384 1123
rect 3378 1118 3384 1119
rect 3442 1123 3448 1124
rect 3442 1119 3443 1123
rect 3447 1119 3448 1123
rect 3442 1118 3448 1119
rect 3738 1123 3744 1124
rect 3738 1119 3739 1123
rect 3743 1119 3744 1123
rect 3738 1118 3744 1119
rect 1934 1115 1940 1116
rect 4386 1115 4392 1116
rect 1770 1114 1776 1115
rect 4386 1111 4387 1115
rect 4391 1114 4392 1115
rect 4391 1112 4990 1114
rect 4391 1111 4392 1112
rect 4386 1110 4392 1111
rect 3983 1107 3989 1108
rect 158 1104 164 1105
rect 110 1103 116 1104
rect 110 1099 111 1103
rect 115 1099 116 1103
rect 158 1100 159 1104
rect 163 1100 164 1104
rect 158 1099 164 1100
rect 358 1104 364 1105
rect 358 1100 359 1104
rect 363 1100 364 1104
rect 358 1099 364 1100
rect 590 1104 596 1105
rect 590 1100 591 1104
rect 595 1100 596 1104
rect 590 1099 596 1100
rect 830 1104 836 1105
rect 830 1100 831 1104
rect 835 1100 836 1104
rect 830 1099 836 1100
rect 1070 1104 1076 1105
rect 1070 1100 1071 1104
rect 1075 1100 1076 1104
rect 1070 1099 1076 1100
rect 1310 1104 1316 1105
rect 1310 1100 1311 1104
rect 1315 1100 1316 1104
rect 1310 1099 1316 1100
rect 1550 1104 1556 1105
rect 1550 1100 1551 1104
rect 1555 1100 1556 1104
rect 1550 1099 1556 1100
rect 1798 1104 1804 1105
rect 1798 1100 1799 1104
rect 1803 1100 1804 1104
rect 1798 1099 1804 1100
rect 1934 1103 1940 1104
rect 1934 1099 1935 1103
rect 1939 1099 1940 1103
rect 3983 1103 3984 1107
rect 3988 1106 3989 1107
rect 4034 1107 4040 1108
rect 4034 1106 4035 1107
rect 3988 1104 4035 1106
rect 3988 1103 3989 1104
rect 3983 1102 3989 1103
rect 4034 1103 4035 1104
rect 4039 1103 4040 1107
rect 4034 1102 4040 1103
rect 4130 1107 4136 1108
rect 4130 1103 4131 1107
rect 4135 1106 4136 1107
rect 4191 1107 4197 1108
rect 4191 1106 4192 1107
rect 4135 1104 4192 1106
rect 4135 1103 4136 1104
rect 4130 1102 4136 1103
rect 4191 1103 4192 1104
rect 4196 1103 4197 1107
rect 4191 1102 4197 1103
rect 4423 1107 4432 1108
rect 4423 1103 4424 1107
rect 4431 1103 4432 1107
rect 4423 1102 4432 1103
rect 4663 1107 4669 1108
rect 4663 1103 4664 1107
rect 4668 1106 4669 1107
rect 4746 1107 4752 1108
rect 4746 1106 4747 1107
rect 4668 1104 4747 1106
rect 4668 1103 4669 1104
rect 4663 1102 4669 1103
rect 4746 1103 4747 1104
rect 4751 1103 4752 1107
rect 4746 1102 4752 1103
rect 4903 1107 4912 1108
rect 4903 1103 4904 1107
rect 4911 1103 4912 1107
rect 4988 1106 4990 1112
rect 5151 1107 5157 1108
rect 5151 1106 5152 1107
rect 4988 1104 5152 1106
rect 4903 1102 4912 1103
rect 5151 1103 5152 1104
rect 5156 1103 5157 1107
rect 5151 1102 5157 1103
rect 5406 1107 5413 1108
rect 5406 1103 5407 1107
rect 5412 1103 5413 1107
rect 5406 1102 5413 1103
rect 5602 1107 5608 1108
rect 5602 1103 5603 1107
rect 5607 1106 5608 1107
rect 5639 1107 5645 1108
rect 5639 1106 5640 1107
rect 5607 1104 5640 1106
rect 5607 1103 5608 1104
rect 5602 1102 5608 1103
rect 5639 1103 5640 1104
rect 5644 1103 5645 1107
rect 5639 1102 5645 1103
rect 110 1098 116 1099
rect 1934 1098 1940 1099
rect 3838 1100 3844 1101
rect 5662 1100 5668 1101
rect 3838 1096 3839 1100
rect 3843 1096 3844 1100
rect 3838 1095 3844 1096
rect 3858 1099 3864 1100
rect 3858 1095 3859 1099
rect 3863 1095 3864 1099
rect 3858 1094 3864 1095
rect 4066 1099 4072 1100
rect 4066 1095 4067 1099
rect 4071 1095 4072 1099
rect 4066 1094 4072 1095
rect 4298 1099 4304 1100
rect 4298 1095 4299 1099
rect 4303 1095 4304 1099
rect 4298 1094 4304 1095
rect 4538 1099 4544 1100
rect 4538 1095 4539 1099
rect 4543 1095 4544 1099
rect 4538 1094 4544 1095
rect 4778 1099 4784 1100
rect 4778 1095 4779 1099
rect 4783 1095 4784 1099
rect 4778 1094 4784 1095
rect 5026 1099 5032 1100
rect 5026 1095 5027 1099
rect 5031 1095 5032 1099
rect 5026 1094 5032 1095
rect 5282 1099 5288 1100
rect 5282 1095 5283 1099
rect 5287 1095 5288 1099
rect 5282 1094 5288 1095
rect 5514 1099 5520 1100
rect 5514 1095 5515 1099
rect 5519 1095 5520 1099
rect 5662 1096 5663 1100
rect 5667 1096 5668 1100
rect 5662 1095 5668 1096
rect 5514 1094 5520 1095
rect 3886 1084 3892 1085
rect 3838 1083 3844 1084
rect 3838 1079 3839 1083
rect 3843 1079 3844 1083
rect 3886 1080 3887 1084
rect 3891 1080 3892 1084
rect 3886 1079 3892 1080
rect 4094 1084 4100 1085
rect 4094 1080 4095 1084
rect 4099 1080 4100 1084
rect 4094 1079 4100 1080
rect 4326 1084 4332 1085
rect 4326 1080 4327 1084
rect 4331 1080 4332 1084
rect 4326 1079 4332 1080
rect 4566 1084 4572 1085
rect 4566 1080 4567 1084
rect 4571 1080 4572 1084
rect 4566 1079 4572 1080
rect 4806 1084 4812 1085
rect 4806 1080 4807 1084
rect 4811 1080 4812 1084
rect 4806 1079 4812 1080
rect 5054 1084 5060 1085
rect 5054 1080 5055 1084
rect 5059 1080 5060 1084
rect 5054 1079 5060 1080
rect 5310 1084 5316 1085
rect 5310 1080 5311 1084
rect 5315 1080 5316 1084
rect 5310 1079 5316 1080
rect 5542 1084 5548 1085
rect 5542 1080 5543 1084
rect 5547 1080 5548 1084
rect 5542 1079 5548 1080
rect 5662 1083 5668 1084
rect 5662 1079 5663 1083
rect 5667 1079 5668 1083
rect 3838 1078 3844 1079
rect 5662 1078 5668 1079
rect 3082 1051 3088 1052
rect 3082 1047 3083 1051
rect 3087 1050 3088 1051
rect 3370 1051 3376 1052
rect 3087 1048 3109 1050
rect 3087 1047 3088 1048
rect 3082 1046 3088 1047
rect 3330 1047 3336 1048
rect 110 1045 116 1046
rect 1934 1045 1940 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 262 1044 268 1045
rect 262 1040 263 1044
rect 267 1040 268 1044
rect 262 1039 268 1040
rect 438 1044 444 1045
rect 438 1040 439 1044
rect 443 1040 444 1044
rect 438 1039 444 1040
rect 614 1044 620 1045
rect 614 1040 615 1044
rect 619 1040 620 1044
rect 614 1039 620 1040
rect 782 1044 788 1045
rect 782 1040 783 1044
rect 787 1040 788 1044
rect 782 1039 788 1040
rect 950 1044 956 1045
rect 950 1040 951 1044
rect 955 1040 956 1044
rect 950 1039 956 1040
rect 1110 1044 1116 1045
rect 1110 1040 1111 1044
rect 1115 1040 1116 1044
rect 1110 1039 1116 1040
rect 1270 1044 1276 1045
rect 1270 1040 1271 1044
rect 1275 1040 1276 1044
rect 1270 1039 1276 1040
rect 1430 1044 1436 1045
rect 1430 1040 1431 1044
rect 1435 1040 1436 1044
rect 1430 1039 1436 1040
rect 1590 1044 1596 1045
rect 1590 1040 1591 1044
rect 1595 1040 1596 1044
rect 1590 1039 1596 1040
rect 1750 1044 1756 1045
rect 1750 1040 1751 1044
rect 1755 1040 1756 1044
rect 1934 1041 1935 1045
rect 1939 1041 1940 1045
rect 3330 1043 3331 1047
rect 3335 1043 3336 1047
rect 3370 1047 3371 1051
rect 3375 1050 3376 1051
rect 3375 1048 3413 1050
rect 3375 1047 3376 1048
rect 3370 1046 3376 1047
rect 3330 1042 3336 1043
rect 1934 1040 1940 1041
rect 1750 1039 1756 1040
rect 234 1029 240 1030
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 234 1025 235 1029
rect 239 1025 240 1029
rect 234 1024 240 1025
rect 410 1029 416 1030
rect 410 1025 411 1029
rect 415 1025 416 1029
rect 410 1024 416 1025
rect 586 1029 592 1030
rect 586 1025 587 1029
rect 591 1025 592 1029
rect 586 1024 592 1025
rect 754 1029 760 1030
rect 754 1025 755 1029
rect 759 1025 760 1029
rect 754 1024 760 1025
rect 922 1029 928 1030
rect 922 1025 923 1029
rect 927 1025 928 1029
rect 922 1024 928 1025
rect 1082 1029 1088 1030
rect 1082 1025 1083 1029
rect 1087 1025 1088 1029
rect 1082 1024 1088 1025
rect 1242 1029 1248 1030
rect 1242 1025 1243 1029
rect 1247 1025 1248 1029
rect 1242 1024 1248 1025
rect 1402 1029 1408 1030
rect 1402 1025 1403 1029
rect 1407 1025 1408 1029
rect 1402 1024 1408 1025
rect 1562 1029 1568 1030
rect 1562 1025 1563 1029
rect 1567 1025 1568 1029
rect 1562 1024 1568 1025
rect 1722 1029 1728 1030
rect 1722 1025 1723 1029
rect 1727 1025 1728 1029
rect 1722 1024 1728 1025
rect 1934 1028 1940 1029
rect 1934 1024 1935 1028
rect 1939 1024 1940 1028
rect 110 1023 116 1024
rect 1934 1023 1940 1024
rect 3838 1025 3844 1026
rect 5662 1025 5668 1026
rect 3838 1021 3839 1025
rect 3843 1021 3844 1025
rect 3838 1020 3844 1021
rect 3886 1024 3892 1025
rect 3886 1020 3887 1024
rect 3891 1020 3892 1024
rect 270 1019 276 1020
rect 270 1015 271 1019
rect 275 1018 276 1019
rect 359 1019 365 1020
rect 359 1018 360 1019
rect 275 1016 360 1018
rect 275 1015 276 1016
rect 270 1014 276 1015
rect 359 1015 360 1016
rect 364 1015 365 1019
rect 359 1014 365 1015
rect 391 1019 397 1020
rect 391 1015 392 1019
rect 396 1018 397 1019
rect 535 1019 541 1020
rect 535 1018 536 1019
rect 396 1016 536 1018
rect 396 1015 397 1016
rect 391 1014 397 1015
rect 535 1015 536 1016
rect 540 1015 541 1019
rect 535 1014 541 1015
rect 658 1019 664 1020
rect 658 1015 659 1019
rect 663 1018 664 1019
rect 711 1019 717 1020
rect 711 1018 712 1019
rect 663 1016 712 1018
rect 663 1015 664 1016
rect 658 1014 664 1015
rect 711 1015 712 1016
rect 716 1015 717 1019
rect 711 1014 717 1015
rect 746 1019 752 1020
rect 746 1015 747 1019
rect 751 1018 752 1019
rect 879 1019 885 1020
rect 879 1018 880 1019
rect 751 1016 880 1018
rect 751 1015 752 1016
rect 746 1014 752 1015
rect 879 1015 880 1016
rect 884 1015 885 1019
rect 879 1014 885 1015
rect 910 1019 916 1020
rect 910 1015 911 1019
rect 915 1018 916 1019
rect 1047 1019 1053 1020
rect 1047 1018 1048 1019
rect 915 1016 1048 1018
rect 915 1015 916 1016
rect 910 1014 916 1015
rect 1047 1015 1048 1016
rect 1052 1015 1053 1019
rect 1047 1014 1053 1015
rect 1207 1019 1213 1020
rect 1207 1015 1208 1019
rect 1212 1018 1213 1019
rect 1258 1019 1264 1020
rect 1258 1018 1259 1019
rect 1212 1016 1259 1018
rect 1212 1015 1213 1016
rect 1207 1014 1213 1015
rect 1258 1015 1259 1016
rect 1263 1015 1264 1019
rect 1258 1014 1264 1015
rect 1367 1019 1373 1020
rect 1367 1015 1368 1019
rect 1372 1018 1373 1019
rect 1418 1019 1424 1020
rect 1418 1018 1419 1019
rect 1372 1016 1419 1018
rect 1372 1015 1373 1016
rect 1367 1014 1373 1015
rect 1418 1015 1419 1016
rect 1423 1015 1424 1019
rect 1418 1014 1424 1015
rect 1527 1019 1533 1020
rect 1527 1015 1528 1019
rect 1532 1018 1533 1019
rect 1578 1019 1584 1020
rect 1578 1018 1579 1019
rect 1532 1016 1579 1018
rect 1532 1015 1533 1016
rect 1527 1014 1533 1015
rect 1578 1015 1579 1016
rect 1583 1015 1584 1019
rect 1578 1014 1584 1015
rect 1687 1019 1693 1020
rect 1687 1015 1688 1019
rect 1692 1018 1693 1019
rect 1738 1019 1744 1020
rect 1738 1018 1739 1019
rect 1692 1016 1739 1018
rect 1692 1015 1693 1016
rect 1687 1014 1693 1015
rect 1738 1015 1739 1016
rect 1743 1015 1744 1019
rect 1738 1014 1744 1015
rect 1758 1019 1764 1020
rect 1758 1015 1759 1019
rect 1763 1018 1764 1019
rect 1847 1019 1853 1020
rect 3886 1019 3892 1020
rect 4070 1024 4076 1025
rect 4070 1020 4071 1024
rect 4075 1020 4076 1024
rect 4070 1019 4076 1020
rect 4278 1024 4284 1025
rect 4278 1020 4279 1024
rect 4283 1020 4284 1024
rect 4278 1019 4284 1020
rect 4510 1024 4516 1025
rect 4510 1020 4511 1024
rect 4515 1020 4516 1024
rect 4510 1019 4516 1020
rect 4758 1024 4764 1025
rect 4758 1020 4759 1024
rect 4763 1020 4764 1024
rect 4758 1019 4764 1020
rect 5022 1024 5028 1025
rect 5022 1020 5023 1024
rect 5027 1020 5028 1024
rect 5022 1019 5028 1020
rect 5294 1024 5300 1025
rect 5294 1020 5295 1024
rect 5299 1020 5300 1024
rect 5294 1019 5300 1020
rect 5542 1024 5548 1025
rect 5542 1020 5543 1024
rect 5547 1020 5548 1024
rect 5662 1021 5663 1025
rect 5667 1021 5668 1025
rect 5662 1020 5668 1021
rect 5542 1019 5548 1020
rect 1847 1018 1848 1019
rect 1763 1016 1848 1018
rect 1763 1015 1764 1016
rect 1758 1014 1764 1015
rect 1847 1015 1848 1016
rect 1852 1015 1853 1019
rect 1847 1014 1853 1015
rect 2986 1015 2992 1016
rect 2986 1011 2987 1015
rect 2991 1014 2992 1015
rect 3215 1015 3221 1016
rect 3215 1014 3216 1015
rect 2991 1012 3216 1014
rect 2991 1011 2992 1012
rect 2986 1010 2992 1011
rect 3215 1011 3216 1012
rect 3220 1011 3221 1015
rect 3215 1010 3221 1011
rect 3367 1015 3376 1016
rect 3367 1011 3368 1015
rect 3375 1011 3376 1015
rect 3367 1010 3376 1011
rect 3378 1015 3384 1016
rect 3378 1011 3379 1015
rect 3383 1014 3384 1015
rect 3519 1015 3525 1016
rect 3519 1014 3520 1015
rect 3383 1012 3520 1014
rect 3383 1011 3384 1012
rect 3378 1010 3384 1011
rect 3519 1011 3520 1012
rect 3524 1011 3525 1015
rect 3519 1010 3525 1011
rect 3858 1009 3864 1010
rect 1974 1008 1980 1009
rect 3798 1008 3804 1009
rect 1974 1004 1975 1008
rect 1979 1004 1980 1008
rect 1974 1003 1980 1004
rect 3090 1007 3096 1008
rect 3090 1003 3091 1007
rect 3095 1003 3096 1007
rect 3090 1002 3096 1003
rect 3242 1007 3248 1008
rect 3242 1003 3243 1007
rect 3247 1003 3248 1007
rect 3242 1002 3248 1003
rect 3394 1007 3400 1008
rect 3394 1003 3395 1007
rect 3399 1003 3400 1007
rect 3798 1004 3799 1008
rect 3803 1004 3804 1008
rect 3798 1003 3804 1004
rect 3838 1008 3844 1009
rect 3838 1004 3839 1008
rect 3843 1004 3844 1008
rect 3858 1005 3859 1009
rect 3863 1005 3864 1009
rect 3858 1004 3864 1005
rect 4042 1009 4048 1010
rect 4042 1005 4043 1009
rect 4047 1005 4048 1009
rect 4042 1004 4048 1005
rect 4250 1009 4256 1010
rect 4250 1005 4251 1009
rect 4255 1005 4256 1009
rect 4250 1004 4256 1005
rect 4482 1009 4488 1010
rect 4482 1005 4483 1009
rect 4487 1005 4488 1009
rect 4482 1004 4488 1005
rect 4730 1009 4736 1010
rect 4730 1005 4731 1009
rect 4735 1005 4736 1009
rect 4730 1004 4736 1005
rect 4994 1009 5000 1010
rect 4994 1005 4995 1009
rect 4999 1005 5000 1009
rect 4994 1004 5000 1005
rect 5266 1009 5272 1010
rect 5266 1005 5267 1009
rect 5271 1005 5272 1009
rect 5266 1004 5272 1005
rect 5514 1009 5520 1010
rect 5514 1005 5515 1009
rect 5519 1005 5520 1009
rect 5514 1004 5520 1005
rect 5662 1008 5668 1009
rect 5662 1004 5663 1008
rect 5667 1004 5668 1008
rect 3838 1003 3844 1004
rect 5662 1003 5668 1004
rect 3394 1002 3400 1003
rect 3962 999 3968 1000
rect 3962 995 3963 999
rect 3967 998 3968 999
rect 3983 999 3989 1000
rect 3983 998 3984 999
rect 3967 996 3984 998
rect 3967 995 3968 996
rect 3962 994 3968 995
rect 3983 995 3984 996
rect 3988 995 3989 999
rect 3983 994 3989 995
rect 4018 999 4024 1000
rect 4018 995 4019 999
rect 4023 998 4024 999
rect 4167 999 4173 1000
rect 4167 998 4168 999
rect 4023 996 4168 998
rect 4023 995 4024 996
rect 4018 994 4024 995
rect 4167 995 4168 996
rect 4172 995 4173 999
rect 4167 994 4173 995
rect 4375 999 4381 1000
rect 4375 995 4376 999
rect 4380 998 4381 999
rect 4498 999 4504 1000
rect 4498 998 4499 999
rect 4380 996 4499 998
rect 4380 995 4381 996
rect 4375 994 4381 995
rect 4498 995 4499 996
rect 4503 995 4504 999
rect 4498 994 4504 995
rect 4607 999 4616 1000
rect 4607 995 4608 999
rect 4615 995 4616 999
rect 4607 994 4616 995
rect 4855 999 4861 1000
rect 4855 995 4856 999
rect 4860 998 4861 999
rect 5010 999 5016 1000
rect 5010 998 5011 999
rect 4860 996 5011 998
rect 4860 995 4861 996
rect 4855 994 4861 995
rect 5010 995 5011 996
rect 5015 995 5016 999
rect 5010 994 5016 995
rect 5119 999 5125 1000
rect 5119 995 5120 999
rect 5124 995 5125 999
rect 5119 994 5125 995
rect 5370 999 5376 1000
rect 5370 995 5371 999
rect 5375 998 5376 999
rect 5391 999 5397 1000
rect 5391 998 5392 999
rect 5375 996 5392 998
rect 5375 995 5376 996
rect 5370 994 5376 995
rect 5391 995 5392 996
rect 5396 995 5397 999
rect 5391 994 5397 995
rect 5610 999 5616 1000
rect 5610 995 5611 999
rect 5615 998 5616 999
rect 5639 999 5645 1000
rect 5639 998 5640 999
rect 5615 996 5640 998
rect 5615 995 5616 996
rect 5610 994 5616 995
rect 5639 995 5640 996
rect 5644 995 5645 999
rect 5639 994 5645 995
rect 3118 992 3124 993
rect 1974 991 1980 992
rect 391 987 397 988
rect 391 986 392 987
rect 325 984 392 986
rect 391 983 392 984
rect 396 983 397 987
rect 391 982 397 983
rect 498 987 504 988
rect 498 983 499 987
rect 503 983 504 987
rect 746 987 752 988
rect 746 986 747 987
rect 677 984 747 986
rect 498 982 504 983
rect 746 983 747 984
rect 751 983 752 987
rect 910 987 916 988
rect 910 986 911 987
rect 845 984 911 986
rect 746 982 752 983
rect 910 983 911 984
rect 915 983 916 987
rect 910 982 916 983
rect 938 987 944 988
rect 938 983 939 987
rect 943 983 944 987
rect 1239 987 1245 988
rect 1239 986 1240 987
rect 1173 984 1240 986
rect 938 982 944 983
rect 1239 983 1240 984
rect 1244 983 1245 987
rect 1239 982 1245 983
rect 1258 987 1264 988
rect 1258 983 1259 987
rect 1263 983 1264 987
rect 1258 982 1264 983
rect 1418 987 1424 988
rect 1418 983 1419 987
rect 1423 983 1424 987
rect 1418 982 1424 983
rect 1578 987 1584 988
rect 1578 983 1579 987
rect 1583 983 1584 987
rect 1578 982 1584 983
rect 1738 987 1744 988
rect 1738 983 1739 987
rect 1743 983 1744 987
rect 1974 987 1975 991
rect 1979 987 1980 991
rect 3118 988 3119 992
rect 3123 988 3124 992
rect 3118 987 3124 988
rect 3270 992 3276 993
rect 3270 988 3271 992
rect 3275 988 3276 992
rect 3270 987 3276 988
rect 3422 992 3428 993
rect 3422 988 3423 992
rect 3427 988 3428 992
rect 3422 987 3428 988
rect 3798 991 3804 992
rect 3798 987 3799 991
rect 3803 987 3804 991
rect 1974 986 1980 987
rect 3798 986 3804 987
rect 4338 991 4344 992
rect 4338 987 4339 991
rect 4343 990 4344 991
rect 5121 990 5123 994
rect 4343 988 5123 990
rect 4343 987 4344 988
rect 4338 986 4344 987
rect 1738 982 1744 983
rect 4018 967 4024 968
rect 4018 966 4019 967
rect 3949 964 4019 966
rect 4018 963 4019 964
rect 4023 963 4024 967
rect 4018 962 4024 963
rect 4130 967 4136 968
rect 4130 963 4131 967
rect 4135 963 4136 967
rect 4130 962 4136 963
rect 4338 967 4344 968
rect 4338 963 4339 967
rect 4343 963 4344 967
rect 4338 962 4344 963
rect 4498 967 4504 968
rect 4498 963 4499 967
rect 4503 963 4504 967
rect 4498 962 4504 963
rect 4746 967 4752 968
rect 4746 963 4747 967
rect 4751 963 4752 967
rect 4746 962 4752 963
rect 5010 967 5016 968
rect 5010 963 5011 967
rect 5015 963 5016 967
rect 5010 962 5016 963
rect 5294 967 5300 968
rect 5294 963 5295 967
rect 5299 963 5300 967
rect 5294 962 5300 963
rect 5602 967 5608 968
rect 5602 963 5603 967
rect 5607 963 5608 967
rect 5602 962 5608 963
rect 354 935 360 936
rect 314 931 320 932
rect 314 927 315 931
rect 319 927 320 931
rect 354 931 355 935
rect 359 934 360 935
rect 658 935 664 936
rect 658 934 659 935
rect 359 932 397 934
rect 629 932 659 934
rect 359 931 360 932
rect 354 930 360 931
rect 658 931 659 932
rect 663 931 664 935
rect 658 930 664 931
rect 666 935 672 936
rect 666 931 667 935
rect 671 934 672 935
rect 842 935 848 936
rect 671 932 733 934
rect 671 931 672 932
rect 666 930 672 931
rect 842 931 843 935
rect 847 934 848 935
rect 1018 935 1024 936
rect 847 932 909 934
rect 847 931 848 932
rect 842 930 848 931
rect 1018 931 1019 935
rect 1023 934 1024 935
rect 1391 935 1397 936
rect 1391 934 1392 935
rect 1023 932 1093 934
rect 1349 932 1392 934
rect 1023 931 1024 932
rect 1018 930 1024 931
rect 1391 931 1392 932
rect 1396 931 1397 935
rect 1606 935 1612 936
rect 1606 934 1607 935
rect 1533 932 1607 934
rect 1391 930 1397 931
rect 1606 931 1607 932
rect 1611 931 1612 935
rect 1775 935 1781 936
rect 1775 934 1776 935
rect 1717 932 1776 934
rect 1606 930 1612 931
rect 1775 931 1776 932
rect 1780 931 1781 935
rect 1967 935 1973 936
rect 1967 934 1968 935
rect 1877 932 1968 934
rect 1775 930 1781 931
rect 1967 931 1968 932
rect 1972 931 1973 935
rect 1967 930 1973 931
rect 314 926 320 927
rect 3962 919 3968 920
rect 3962 915 3963 919
rect 3967 918 3968 919
rect 4306 919 4312 920
rect 3967 916 3989 918
rect 3967 915 3968 916
rect 3962 914 3968 915
rect 4266 915 4272 916
rect 4266 911 4267 915
rect 4271 911 4272 915
rect 4306 915 4307 919
rect 4311 918 4312 919
rect 4610 919 4616 920
rect 4311 916 4421 918
rect 4311 915 4312 916
rect 4306 914 4312 915
rect 4610 915 4611 919
rect 4615 918 4616 919
rect 4866 919 4872 920
rect 4615 916 4661 918
rect 4615 915 4616 916
rect 4610 914 4616 915
rect 4866 915 4867 919
rect 4871 918 4872 919
rect 5375 919 5381 920
rect 5375 918 5376 919
rect 4871 916 4917 918
rect 5261 916 5376 918
rect 4871 915 4872 916
rect 4866 914 4872 915
rect 5375 915 5376 916
rect 5380 915 5381 919
rect 5375 914 5381 915
rect 5530 915 5536 916
rect 4266 910 4272 911
rect 5530 911 5531 915
rect 5535 911 5536 915
rect 5530 910 5536 911
rect 1974 905 1980 906
rect 3798 905 3804 906
rect 1974 901 1975 905
rect 1979 901 1980 905
rect 1974 900 1980 901
rect 2046 904 2052 905
rect 2046 900 2047 904
rect 2051 900 2052 904
rect 351 899 360 900
rect 351 895 352 899
rect 359 895 360 899
rect 351 894 360 895
rect 498 899 509 900
rect 498 895 499 899
rect 503 895 504 899
rect 508 895 509 899
rect 498 894 509 895
rect 663 899 672 900
rect 663 895 664 899
rect 671 895 672 899
rect 663 894 672 895
rect 839 899 848 900
rect 839 895 840 899
rect 847 895 848 899
rect 839 894 848 895
rect 1015 899 1024 900
rect 1015 895 1016 899
rect 1023 895 1024 899
rect 1015 894 1024 895
rect 1199 899 1205 900
rect 1199 895 1200 899
rect 1204 898 1205 899
rect 1226 899 1232 900
rect 1226 898 1227 899
rect 1204 896 1227 898
rect 1204 895 1205 896
rect 1199 894 1205 895
rect 1226 895 1227 896
rect 1231 895 1232 899
rect 1226 894 1232 895
rect 1239 899 1245 900
rect 1239 895 1240 899
rect 1244 898 1245 899
rect 1383 899 1389 900
rect 1383 898 1384 899
rect 1244 896 1384 898
rect 1244 895 1245 896
rect 1239 894 1245 895
rect 1383 895 1384 896
rect 1388 895 1389 899
rect 1383 894 1389 895
rect 1391 899 1397 900
rect 1391 895 1392 899
rect 1396 898 1397 899
rect 1567 899 1573 900
rect 1567 898 1568 899
rect 1396 896 1568 898
rect 1396 895 1397 896
rect 1391 894 1397 895
rect 1567 895 1568 896
rect 1572 895 1573 899
rect 1567 894 1573 895
rect 1606 899 1612 900
rect 1606 895 1607 899
rect 1611 898 1612 899
rect 1751 899 1757 900
rect 1751 898 1752 899
rect 1611 896 1752 898
rect 1611 895 1612 896
rect 1606 894 1612 895
rect 1751 895 1752 896
rect 1756 895 1757 899
rect 1751 894 1757 895
rect 1775 899 1781 900
rect 1775 895 1776 899
rect 1780 898 1781 899
rect 1911 899 1917 900
rect 2046 899 2052 900
rect 2350 904 2356 905
rect 2350 900 2351 904
rect 2355 900 2356 904
rect 2350 899 2356 900
rect 2646 904 2652 905
rect 2646 900 2647 904
rect 2651 900 2652 904
rect 2646 899 2652 900
rect 2926 904 2932 905
rect 2926 900 2927 904
rect 2931 900 2932 904
rect 2926 899 2932 900
rect 3206 904 3212 905
rect 3206 900 3207 904
rect 3211 900 3212 904
rect 3206 899 3212 900
rect 3494 904 3500 905
rect 3494 900 3495 904
rect 3499 900 3500 904
rect 3798 901 3799 905
rect 3803 901 3804 905
rect 3798 900 3804 901
rect 3494 899 3500 900
rect 1911 898 1912 899
rect 1780 896 1912 898
rect 1780 895 1781 896
rect 1775 894 1781 895
rect 1911 895 1912 896
rect 1916 895 1917 899
rect 1911 894 1917 895
rect 110 892 116 893
rect 1934 892 1940 893
rect 110 888 111 892
rect 115 888 116 892
rect 110 887 116 888
rect 226 891 232 892
rect 226 887 227 891
rect 231 887 232 891
rect 226 886 232 887
rect 378 891 384 892
rect 378 887 379 891
rect 383 887 384 891
rect 378 886 384 887
rect 538 891 544 892
rect 538 887 539 891
rect 543 887 544 891
rect 538 886 544 887
rect 714 891 720 892
rect 714 887 715 891
rect 719 887 720 891
rect 714 886 720 887
rect 890 891 896 892
rect 890 887 891 891
rect 895 887 896 891
rect 890 886 896 887
rect 1074 891 1080 892
rect 1074 887 1075 891
rect 1079 887 1080 891
rect 1074 886 1080 887
rect 1258 891 1264 892
rect 1258 887 1259 891
rect 1263 887 1264 891
rect 1258 886 1264 887
rect 1442 891 1448 892
rect 1442 887 1443 891
rect 1447 887 1448 891
rect 1442 886 1448 887
rect 1626 891 1632 892
rect 1626 887 1627 891
rect 1631 887 1632 891
rect 1626 886 1632 887
rect 1786 891 1792 892
rect 1786 887 1787 891
rect 1791 887 1792 891
rect 1934 888 1935 892
rect 1939 888 1940 892
rect 4266 891 4272 892
rect 2018 889 2024 890
rect 1934 887 1940 888
rect 1974 888 1980 889
rect 1786 886 1792 887
rect 1974 884 1975 888
rect 1979 884 1980 888
rect 2018 885 2019 889
rect 2023 885 2024 889
rect 2018 884 2024 885
rect 2322 889 2328 890
rect 2322 885 2323 889
rect 2327 885 2328 889
rect 2322 884 2328 885
rect 2618 889 2624 890
rect 2618 885 2619 889
rect 2623 885 2624 889
rect 2618 884 2624 885
rect 2898 889 2904 890
rect 2898 885 2899 889
rect 2903 885 2904 889
rect 2898 884 2904 885
rect 3178 889 3184 890
rect 3178 885 3179 889
rect 3183 885 3184 889
rect 3178 884 3184 885
rect 3466 889 3472 890
rect 3466 885 3467 889
rect 3471 885 3472 889
rect 3466 884 3472 885
rect 3798 888 3804 889
rect 3798 884 3799 888
rect 3803 884 3804 888
rect 4266 887 4267 891
rect 4271 890 4272 891
rect 4271 888 4821 890
rect 4271 887 4272 888
rect 4266 886 4272 887
rect 4819 886 4821 888
rect 4819 884 4926 886
rect 1974 883 1980 884
rect 3798 883 3804 884
rect 4095 883 4101 884
rect 1967 879 1973 880
rect 254 876 260 877
rect 110 875 116 876
rect 110 871 111 875
rect 115 871 116 875
rect 254 872 255 876
rect 259 872 260 876
rect 254 871 260 872
rect 406 876 412 877
rect 406 872 407 876
rect 411 872 412 876
rect 406 871 412 872
rect 566 876 572 877
rect 566 872 567 876
rect 571 872 572 876
rect 566 871 572 872
rect 742 876 748 877
rect 742 872 743 876
rect 747 872 748 876
rect 742 871 748 872
rect 918 876 924 877
rect 918 872 919 876
rect 923 872 924 876
rect 918 871 924 872
rect 1102 876 1108 877
rect 1102 872 1103 876
rect 1107 872 1108 876
rect 1102 871 1108 872
rect 1286 876 1292 877
rect 1286 872 1287 876
rect 1291 872 1292 876
rect 1286 871 1292 872
rect 1470 876 1476 877
rect 1470 872 1471 876
rect 1475 872 1476 876
rect 1470 871 1476 872
rect 1654 876 1660 877
rect 1654 872 1655 876
rect 1659 872 1660 876
rect 1654 871 1660 872
rect 1814 876 1820 877
rect 1814 872 1815 876
rect 1819 872 1820 876
rect 1814 871 1820 872
rect 1934 875 1940 876
rect 1934 871 1935 875
rect 1939 871 1940 875
rect 1967 875 1968 879
rect 1972 878 1973 879
rect 2143 879 2149 880
rect 2143 878 2144 879
rect 1972 876 2144 878
rect 1972 875 1973 876
rect 1967 874 1973 875
rect 2143 875 2144 876
rect 2148 875 2149 879
rect 2143 874 2149 875
rect 2166 879 2172 880
rect 2166 875 2167 879
rect 2171 878 2172 879
rect 2447 879 2453 880
rect 2447 878 2448 879
rect 2171 876 2448 878
rect 2171 875 2172 876
rect 2166 874 2172 875
rect 2447 875 2448 876
rect 2452 875 2453 879
rect 2447 874 2453 875
rect 2743 879 2752 880
rect 2743 875 2744 879
rect 2751 875 2752 879
rect 2743 874 2752 875
rect 2830 879 2836 880
rect 2830 875 2831 879
rect 2835 878 2836 879
rect 3023 879 3029 880
rect 3023 878 3024 879
rect 2835 876 3024 878
rect 2835 875 2836 876
rect 2830 874 2836 875
rect 3023 875 3024 876
rect 3028 875 3029 879
rect 3023 874 3029 875
rect 3303 879 3309 880
rect 3303 875 3304 879
rect 3308 878 3309 879
rect 3330 879 3336 880
rect 3330 878 3331 879
rect 3308 876 3331 878
rect 3308 875 3309 876
rect 3303 874 3309 875
rect 3330 875 3331 876
rect 3335 875 3336 879
rect 3330 874 3336 875
rect 3378 879 3384 880
rect 3378 875 3379 879
rect 3383 878 3384 879
rect 3591 879 3597 880
rect 3591 878 3592 879
rect 3383 876 3592 878
rect 3383 875 3384 876
rect 3378 874 3384 875
rect 3591 875 3592 876
rect 3596 875 3597 879
rect 4095 879 4096 883
rect 4100 882 4101 883
rect 4266 883 4272 884
rect 4266 882 4267 883
rect 4100 880 4267 882
rect 4100 879 4101 880
rect 4095 878 4101 879
rect 4266 879 4267 880
rect 4271 879 4272 883
rect 4266 878 4272 879
rect 4303 883 4312 884
rect 4303 879 4304 883
rect 4311 879 4312 883
rect 4303 878 4312 879
rect 4527 883 4533 884
rect 4527 879 4528 883
rect 4532 882 4533 883
rect 4546 883 4552 884
rect 4546 882 4547 883
rect 4532 880 4547 882
rect 4532 879 4533 880
rect 4527 878 4533 879
rect 4546 879 4547 880
rect 4551 879 4552 883
rect 4546 878 4552 879
rect 4767 883 4773 884
rect 4767 879 4768 883
rect 4772 882 4773 883
rect 4924 882 4926 884
rect 5023 883 5029 884
rect 5023 882 5024 883
rect 4772 880 4821 882
rect 4924 880 5024 882
rect 4772 879 4773 880
rect 4767 878 4773 879
rect 4819 878 4821 880
rect 4866 879 4872 880
rect 4866 878 4867 879
rect 3591 874 3597 875
rect 3838 876 3844 877
rect 4819 876 4867 878
rect 3838 872 3839 876
rect 3843 872 3844 876
rect 3838 871 3844 872
rect 3970 875 3976 876
rect 3970 871 3971 875
rect 3975 871 3976 875
rect 110 870 116 871
rect 1934 870 1940 871
rect 3970 870 3976 871
rect 4178 875 4184 876
rect 4178 871 4179 875
rect 4183 871 4184 875
rect 4178 870 4184 871
rect 4402 875 4408 876
rect 4402 871 4403 875
rect 4407 871 4408 875
rect 4402 870 4408 871
rect 4642 875 4648 876
rect 4642 871 4643 875
rect 4647 871 4648 875
rect 4866 875 4867 876
rect 4871 875 4872 879
rect 5023 879 5024 880
rect 5028 879 5029 883
rect 5023 878 5029 879
rect 5294 883 5301 884
rect 5294 879 5295 883
rect 5300 879 5301 883
rect 5294 878 5301 879
rect 5375 883 5381 884
rect 5375 879 5376 883
rect 5380 882 5381 883
rect 5567 883 5573 884
rect 5567 882 5568 883
rect 5380 880 5568 882
rect 5380 879 5381 880
rect 5375 878 5381 879
rect 5567 879 5568 880
rect 5572 879 5573 883
rect 5567 878 5573 879
rect 5662 876 5668 877
rect 4866 874 4872 875
rect 4898 875 4904 876
rect 4642 870 4648 871
rect 4898 871 4899 875
rect 4903 871 4904 875
rect 4898 870 4904 871
rect 5170 875 5176 876
rect 5170 871 5171 875
rect 5175 871 5176 875
rect 5170 870 5176 871
rect 5442 875 5448 876
rect 5442 871 5443 875
rect 5447 871 5448 875
rect 5662 872 5663 876
rect 5667 872 5668 876
rect 5662 871 5668 872
rect 5442 870 5448 871
rect 3998 860 4004 861
rect 3838 859 3844 860
rect 3838 855 3839 859
rect 3843 855 3844 859
rect 3998 856 3999 860
rect 4003 856 4004 860
rect 3998 855 4004 856
rect 4206 860 4212 861
rect 4206 856 4207 860
rect 4211 856 4212 860
rect 4206 855 4212 856
rect 4430 860 4436 861
rect 4430 856 4431 860
rect 4435 856 4436 860
rect 4430 855 4436 856
rect 4670 860 4676 861
rect 4670 856 4671 860
rect 4675 856 4676 860
rect 4670 855 4676 856
rect 4926 860 4932 861
rect 4926 856 4927 860
rect 4931 856 4932 860
rect 4926 855 4932 856
rect 5198 860 5204 861
rect 5198 856 5199 860
rect 5203 856 5204 860
rect 5198 855 5204 856
rect 5470 860 5476 861
rect 5470 856 5471 860
rect 5475 856 5476 860
rect 5470 855 5476 856
rect 5662 859 5668 860
rect 5662 855 5663 859
rect 5667 855 5668 859
rect 3838 854 3844 855
rect 5662 854 5668 855
rect 2166 847 2172 848
rect 2166 846 2167 847
rect 2109 844 2167 846
rect 2166 843 2167 844
rect 2171 843 2172 847
rect 2166 842 2172 843
rect 2410 847 2416 848
rect 2410 843 2411 847
rect 2415 843 2416 847
rect 2830 847 2836 848
rect 2830 846 2831 847
rect 2709 844 2831 846
rect 2410 842 2416 843
rect 2830 843 2831 844
rect 2835 843 2836 847
rect 2830 842 2836 843
rect 2986 847 2992 848
rect 2986 843 2987 847
rect 2991 843 2992 847
rect 3378 847 3384 848
rect 3378 846 3379 847
rect 3269 844 3379 846
rect 2986 842 2992 843
rect 3378 843 3379 844
rect 3383 843 3384 847
rect 3378 842 3384 843
rect 3554 847 3560 848
rect 3554 843 3555 847
rect 3559 843 3560 847
rect 3554 842 3560 843
rect 110 801 116 802
rect 1934 801 1940 802
rect 110 797 111 801
rect 115 797 116 801
rect 110 796 116 797
rect 374 800 380 801
rect 374 796 375 800
rect 379 796 380 800
rect 374 795 380 796
rect 654 800 660 801
rect 654 796 655 800
rect 659 796 660 800
rect 654 795 660 796
rect 942 800 948 801
rect 942 796 943 800
rect 947 796 948 800
rect 942 795 948 796
rect 1238 800 1244 801
rect 1238 796 1239 800
rect 1243 796 1244 800
rect 1238 795 1244 796
rect 1534 800 1540 801
rect 1534 796 1535 800
rect 1539 796 1540 800
rect 1534 795 1540 796
rect 1814 800 1820 801
rect 1814 796 1815 800
rect 1819 796 1820 800
rect 1934 797 1935 801
rect 1939 797 1940 801
rect 3838 801 3844 802
rect 5662 801 5668 802
rect 1934 796 1940 797
rect 1942 799 1948 800
rect 1814 795 1820 796
rect 1942 795 1943 799
rect 1947 798 1948 799
rect 2122 799 2128 800
rect 1947 796 2013 798
rect 1947 795 1948 796
rect 1942 794 1948 795
rect 2122 795 2123 799
rect 2127 798 2128 799
rect 2378 799 2384 800
rect 2127 796 2269 798
rect 2127 795 2128 796
rect 2122 794 2128 795
rect 2378 795 2379 799
rect 2383 798 2384 799
rect 2746 799 2752 800
rect 2383 796 2541 798
rect 2383 795 2384 796
rect 2378 794 2384 795
rect 2746 795 2747 799
rect 2751 798 2752 799
rect 2898 799 2904 800
rect 2751 796 2789 798
rect 2751 795 2752 796
rect 2746 794 2752 795
rect 2898 795 2899 799
rect 2903 798 2904 799
rect 3354 799 3360 800
rect 2903 796 3021 798
rect 2903 795 2904 796
rect 2898 794 2904 795
rect 3314 795 3320 796
rect 3314 791 3315 795
rect 3319 791 3320 795
rect 3354 795 3355 799
rect 3359 798 3360 799
rect 3359 796 3469 798
rect 3741 796 3834 798
rect 3838 797 3839 801
rect 3843 797 3844 801
rect 3838 796 3844 797
rect 3886 800 3892 801
rect 3886 796 3887 800
rect 3891 796 3892 800
rect 3359 795 3360 796
rect 3354 794 3360 795
rect 3832 794 3834 796
rect 3866 795 3872 796
rect 3886 795 3892 796
rect 4046 800 4052 801
rect 4046 796 4047 800
rect 4051 796 4052 800
rect 4046 795 4052 796
rect 4278 800 4284 801
rect 4278 796 4279 800
rect 4283 796 4284 800
rect 4278 795 4284 796
rect 4558 800 4564 801
rect 4558 796 4559 800
rect 4563 796 4564 800
rect 4558 795 4564 796
rect 4878 800 4884 801
rect 4878 796 4879 800
rect 4883 796 4884 800
rect 4878 795 4884 796
rect 5222 800 5228 801
rect 5222 796 5223 800
rect 5227 796 5228 800
rect 5222 795 5228 796
rect 5542 800 5548 801
rect 5542 796 5543 800
rect 5547 796 5548 800
rect 5662 797 5663 801
rect 5667 797 5668 801
rect 5662 796 5668 797
rect 5542 795 5548 796
rect 3866 794 3867 795
rect 3832 792 3867 794
rect 3314 790 3320 791
rect 3866 791 3867 792
rect 3871 791 3872 795
rect 3866 790 3872 791
rect 346 785 352 786
rect 110 784 116 785
rect 110 780 111 784
rect 115 780 116 784
rect 346 781 347 785
rect 351 781 352 785
rect 346 780 352 781
rect 626 785 632 786
rect 626 781 627 785
rect 631 781 632 785
rect 626 780 632 781
rect 914 785 920 786
rect 914 781 915 785
rect 919 781 920 785
rect 914 780 920 781
rect 1210 785 1216 786
rect 1210 781 1211 785
rect 1215 781 1216 785
rect 1210 780 1216 781
rect 1506 785 1512 786
rect 1506 781 1507 785
rect 1511 781 1512 785
rect 1506 780 1512 781
rect 1786 785 1792 786
rect 3858 785 3864 786
rect 1786 781 1787 785
rect 1791 781 1792 785
rect 1786 780 1792 781
rect 1934 784 1940 785
rect 1934 780 1935 784
rect 1939 780 1940 784
rect 110 779 116 780
rect 1934 779 1940 780
rect 3838 784 3844 785
rect 3838 780 3839 784
rect 3843 780 3844 784
rect 3858 781 3859 785
rect 3863 781 3864 785
rect 3858 780 3864 781
rect 4018 785 4024 786
rect 4018 781 4019 785
rect 4023 781 4024 785
rect 4018 780 4024 781
rect 4250 785 4256 786
rect 4250 781 4251 785
rect 4255 781 4256 785
rect 4250 780 4256 781
rect 4530 785 4536 786
rect 4530 781 4531 785
rect 4535 781 4536 785
rect 4530 780 4536 781
rect 4850 785 4856 786
rect 4850 781 4851 785
rect 4855 781 4856 785
rect 4850 780 4856 781
rect 5194 785 5200 786
rect 5194 781 5195 785
rect 5199 781 5200 785
rect 5194 780 5200 781
rect 5514 785 5520 786
rect 5514 781 5515 785
rect 5519 781 5520 785
rect 5514 780 5520 781
rect 5662 784 5668 785
rect 5662 780 5663 784
rect 5667 780 5668 784
rect 3838 779 3844 780
rect 5662 779 5668 780
rect 471 775 477 776
rect 471 771 472 775
rect 476 774 477 775
rect 642 775 648 776
rect 642 774 643 775
rect 476 772 643 774
rect 476 771 477 772
rect 471 770 477 771
rect 642 771 643 772
rect 647 771 648 775
rect 751 775 757 776
rect 751 774 752 775
rect 642 770 648 771
rect 684 772 752 774
rect 314 767 320 768
rect 314 763 315 767
rect 319 766 320 767
rect 684 766 686 772
rect 751 771 752 772
rect 756 771 757 775
rect 751 770 757 771
rect 1018 775 1024 776
rect 1018 771 1019 775
rect 1023 774 1024 775
rect 1039 775 1045 776
rect 1039 774 1040 775
rect 1023 772 1040 774
rect 1023 771 1024 772
rect 1018 770 1024 771
rect 1039 771 1040 772
rect 1044 771 1045 775
rect 1039 770 1045 771
rect 1134 775 1140 776
rect 1134 771 1135 775
rect 1139 774 1140 775
rect 1335 775 1341 776
rect 1335 774 1336 775
rect 1139 772 1336 774
rect 1139 771 1140 772
rect 1134 770 1140 771
rect 1335 771 1336 772
rect 1340 771 1341 775
rect 1335 770 1341 771
rect 1631 775 1637 776
rect 1631 771 1632 775
rect 1636 774 1637 775
rect 1802 775 1808 776
rect 1802 774 1803 775
rect 1636 772 1803 774
rect 1636 771 1637 772
rect 1631 770 1637 771
rect 1802 771 1803 772
rect 1807 771 1808 775
rect 1802 770 1808 771
rect 1911 775 1917 776
rect 1911 771 1912 775
rect 1916 774 1917 775
rect 1942 775 1948 776
rect 1942 774 1943 775
rect 1916 772 1943 774
rect 1916 771 1917 772
rect 1911 770 1917 771
rect 1942 771 1943 772
rect 1947 771 1948 775
rect 3983 775 3992 776
rect 1942 770 1948 771
rect 3314 771 3320 772
rect 3314 767 3315 771
rect 3319 770 3320 771
rect 3983 771 3984 775
rect 3991 771 3992 775
rect 3983 770 3992 771
rect 4026 775 4032 776
rect 4026 771 4027 775
rect 4031 774 4032 775
rect 4143 775 4149 776
rect 4143 774 4144 775
rect 4031 772 4144 774
rect 4031 771 4032 772
rect 4026 770 4032 771
rect 4143 771 4144 772
rect 4148 771 4149 775
rect 4143 770 4149 771
rect 4375 775 4381 776
rect 4375 771 4376 775
rect 4380 774 4381 775
rect 4503 775 4509 776
rect 4503 774 4504 775
rect 4380 772 4504 774
rect 4380 771 4381 772
rect 4375 770 4381 771
rect 4503 771 4504 772
rect 4508 771 4509 775
rect 4503 770 4509 771
rect 4655 775 4661 776
rect 4655 771 4656 775
rect 4660 774 4661 775
rect 4866 775 4872 776
rect 4866 774 4867 775
rect 4660 772 4867 774
rect 4660 771 4661 772
rect 4655 770 4661 771
rect 4866 771 4867 772
rect 4871 771 4872 775
rect 4866 770 4872 771
rect 4975 775 4981 776
rect 4975 771 4976 775
rect 4980 774 4981 775
rect 5210 775 5216 776
rect 5210 774 5211 775
rect 4980 772 5211 774
rect 4980 771 4981 772
rect 4975 770 4981 771
rect 5210 771 5211 772
rect 5215 771 5216 775
rect 5319 775 5325 776
rect 5319 774 5320 775
rect 5210 770 5216 771
rect 5220 772 5320 774
rect 3319 768 3586 770
rect 3319 767 3320 768
rect 3314 766 3320 767
rect 319 764 686 766
rect 319 763 320 764
rect 314 762 320 763
rect 2119 763 2128 764
rect 1910 759 1916 760
rect 1910 758 1911 759
rect 1596 756 1911 758
rect 430 743 436 744
rect 430 739 431 743
rect 435 739 436 743
rect 430 738 436 739
rect 642 743 648 744
rect 642 739 643 743
rect 647 739 648 743
rect 1134 743 1140 744
rect 1134 742 1135 743
rect 1005 740 1135 742
rect 642 738 648 739
rect 1134 739 1135 740
rect 1139 739 1140 743
rect 1134 738 1140 739
rect 1226 743 1232 744
rect 1226 739 1227 743
rect 1231 739 1232 743
rect 1596 741 1598 756
rect 1910 755 1911 756
rect 1915 755 1916 759
rect 2119 759 2120 763
rect 2127 759 2128 763
rect 2119 758 2128 759
rect 2375 763 2384 764
rect 2375 759 2376 763
rect 2383 759 2384 763
rect 2375 758 2384 759
rect 2410 763 2416 764
rect 2410 759 2411 763
rect 2415 762 2416 763
rect 2647 763 2653 764
rect 2647 762 2648 763
rect 2415 760 2648 762
rect 2415 759 2416 760
rect 2410 758 2416 759
rect 2647 759 2648 760
rect 2652 759 2653 763
rect 2647 758 2653 759
rect 2895 763 2904 764
rect 2895 759 2896 763
rect 2903 759 2904 763
rect 2895 758 2904 759
rect 3127 763 3133 764
rect 3127 759 3128 763
rect 3132 762 3133 763
rect 3298 763 3304 764
rect 3298 762 3299 763
rect 3132 760 3299 762
rect 3132 759 3133 760
rect 3127 758 3133 759
rect 3298 759 3299 760
rect 3303 759 3304 763
rect 3298 758 3304 759
rect 3351 763 3360 764
rect 3351 759 3352 763
rect 3359 759 3360 763
rect 3351 758 3360 759
rect 3554 763 3560 764
rect 3554 759 3555 763
rect 3559 762 3560 763
rect 3575 763 3581 764
rect 3575 762 3576 763
rect 3559 760 3576 762
rect 3559 759 3560 760
rect 3554 758 3560 759
rect 3575 759 3576 760
rect 3580 759 3581 763
rect 3584 762 3586 768
rect 3775 763 3781 764
rect 3775 762 3776 763
rect 3584 760 3776 762
rect 3575 758 3581 759
rect 3775 759 3776 760
rect 3780 759 3781 763
rect 3775 758 3781 759
rect 5220 758 5222 772
rect 5319 771 5320 772
rect 5324 771 5325 775
rect 5319 770 5325 771
rect 5530 775 5536 776
rect 5530 771 5531 775
rect 5535 774 5536 775
rect 5639 775 5645 776
rect 5639 774 5640 775
rect 5535 772 5640 774
rect 5535 771 5536 772
rect 5530 770 5536 771
rect 5639 771 5640 772
rect 5644 771 5645 775
rect 5639 770 5645 771
rect 1910 754 1916 755
rect 1974 756 1980 757
rect 3798 756 3804 757
rect 1974 752 1975 756
rect 1979 752 1980 756
rect 1974 751 1980 752
rect 1994 755 2000 756
rect 1994 751 1995 755
rect 1999 751 2000 755
rect 1994 750 2000 751
rect 2250 755 2256 756
rect 2250 751 2251 755
rect 2255 751 2256 755
rect 2250 750 2256 751
rect 2522 755 2528 756
rect 2522 751 2523 755
rect 2527 751 2528 755
rect 2522 750 2528 751
rect 2770 755 2776 756
rect 2770 751 2771 755
rect 2775 751 2776 755
rect 2770 750 2776 751
rect 3002 755 3008 756
rect 3002 751 3003 755
rect 3007 751 3008 755
rect 3002 750 3008 751
rect 3226 755 3232 756
rect 3226 751 3227 755
rect 3231 751 3232 755
rect 3226 750 3232 751
rect 3450 755 3456 756
rect 3450 751 3451 755
rect 3455 751 3456 755
rect 3450 750 3456 751
rect 3650 755 3656 756
rect 3650 751 3651 755
rect 3655 751 3656 755
rect 3798 752 3799 756
rect 3803 752 3804 756
rect 3798 751 3804 752
rect 4257 756 5222 758
rect 3650 750 3656 751
rect 1802 743 1808 744
rect 1226 738 1232 739
rect 1802 739 1803 743
rect 1807 739 1808 743
rect 4026 743 4032 744
rect 4026 742 4027 743
rect 2022 740 2028 741
rect 1802 738 1808 739
rect 1974 739 1980 740
rect 1974 735 1975 739
rect 1979 735 1980 739
rect 2022 736 2023 740
rect 2027 736 2028 740
rect 2022 735 2028 736
rect 2278 740 2284 741
rect 2278 736 2279 740
rect 2283 736 2284 740
rect 2278 735 2284 736
rect 2550 740 2556 741
rect 2550 736 2551 740
rect 2555 736 2556 740
rect 2550 735 2556 736
rect 2798 740 2804 741
rect 2798 736 2799 740
rect 2803 736 2804 740
rect 2798 735 2804 736
rect 3030 740 3036 741
rect 3030 736 3031 740
rect 3035 736 3036 740
rect 3030 735 3036 736
rect 3254 740 3260 741
rect 3254 736 3255 740
rect 3259 736 3260 740
rect 3254 735 3260 736
rect 3478 740 3484 741
rect 3478 736 3479 740
rect 3483 736 3484 740
rect 3478 735 3484 736
rect 3678 740 3684 741
rect 3949 740 4027 742
rect 3678 736 3679 740
rect 3683 736 3684 740
rect 3678 735 3684 736
rect 3798 739 3804 740
rect 3798 735 3799 739
rect 3803 735 3804 739
rect 4026 739 4027 740
rect 4031 739 4032 743
rect 4257 742 4259 756
rect 4109 740 4259 742
rect 4266 743 4272 744
rect 4026 738 4032 739
rect 4266 739 4267 743
rect 4271 739 4272 743
rect 4266 738 4272 739
rect 4546 743 4552 744
rect 4546 739 4547 743
rect 4551 739 4552 743
rect 4546 738 4552 739
rect 4866 743 4872 744
rect 4866 739 4867 743
rect 4871 739 4872 743
rect 4866 738 4872 739
rect 5210 743 5216 744
rect 5210 739 5211 743
rect 5215 739 5216 743
rect 5610 743 5616 744
rect 5610 742 5611 743
rect 5605 740 5611 742
rect 5210 738 5216 739
rect 5610 739 5611 740
rect 5615 739 5616 743
rect 5610 738 5616 739
rect 1974 734 1980 735
rect 3798 734 3804 735
rect 258 695 264 696
rect 258 691 259 695
rect 263 694 264 695
rect 474 695 480 696
rect 263 692 325 694
rect 263 691 264 692
rect 258 690 264 691
rect 474 691 475 695
rect 479 694 480 695
rect 810 695 816 696
rect 479 692 517 694
rect 479 691 480 692
rect 474 690 480 691
rect 810 691 811 695
rect 815 694 816 695
rect 1018 695 1024 696
rect 815 692 877 694
rect 815 691 816 692
rect 810 690 816 691
rect 1018 691 1019 695
rect 1023 694 1024 695
rect 1319 695 1325 696
rect 1023 692 1045 694
rect 1023 691 1024 692
rect 1018 690 1024 691
rect 1274 691 1280 692
rect 216 678 218 689
rect 583 679 589 680
rect 583 678 584 679
rect 216 676 584 678
rect 583 675 584 676
rect 588 675 589 679
rect 768 678 770 689
rect 1274 687 1275 691
rect 1279 687 1280 691
rect 1319 691 1320 695
rect 1324 694 1325 695
rect 1471 695 1477 696
rect 1324 692 1357 694
rect 1324 691 1325 692
rect 1319 690 1325 691
rect 1471 691 1472 695
rect 1476 694 1477 695
rect 1639 695 1645 696
rect 1476 692 1509 694
rect 1476 691 1477 692
rect 1471 690 1477 691
rect 1639 691 1640 695
rect 1644 694 1645 695
rect 1783 695 1789 696
rect 1644 692 1669 694
rect 1644 691 1645 692
rect 1639 690 1645 691
rect 1783 691 1784 695
rect 1788 694 1789 695
rect 1788 692 1805 694
rect 1788 691 1789 692
rect 1783 690 1789 691
rect 1274 686 1280 687
rect 3986 687 3992 688
rect 3946 683 3952 684
rect 1150 679 1156 680
rect 1150 678 1151 679
rect 768 676 1151 678
rect 583 674 589 675
rect 1150 675 1151 676
rect 1155 675 1156 679
rect 3946 679 3947 683
rect 3951 679 3952 683
rect 3986 683 3987 687
rect 3991 686 3992 687
rect 4127 687 4133 688
rect 3991 684 4013 686
rect 3991 683 3992 684
rect 3986 682 3992 683
rect 4127 683 4128 687
rect 4132 686 4133 687
rect 4263 687 4269 688
rect 4132 684 4149 686
rect 4132 683 4133 684
rect 4127 682 4133 683
rect 4263 683 4264 687
rect 4268 686 4269 687
rect 4399 687 4405 688
rect 4268 684 4285 686
rect 4268 683 4269 684
rect 4263 682 4269 683
rect 4399 683 4400 687
rect 4404 686 4405 687
rect 4503 687 4509 688
rect 4404 684 4421 686
rect 4404 683 4405 684
rect 4399 682 4405 683
rect 4503 683 4504 687
rect 4508 686 4509 687
rect 4698 687 4704 688
rect 4508 684 4589 686
rect 4508 683 4509 684
rect 4503 682 4509 683
rect 4698 683 4699 687
rect 4703 686 4704 687
rect 4898 687 4904 688
rect 4703 684 4789 686
rect 4703 683 4704 684
rect 4698 682 4704 683
rect 4898 683 4899 687
rect 4903 686 4904 687
rect 5122 687 5128 688
rect 4903 684 5013 686
rect 4903 683 4904 684
rect 4898 682 4904 683
rect 5122 683 5123 687
rect 5127 686 5128 687
rect 5127 684 5245 686
rect 5127 683 5128 684
rect 5122 682 5128 683
rect 5546 683 5552 684
rect 3946 678 3952 679
rect 5546 679 5547 683
rect 5551 679 5552 683
rect 5546 678 5552 679
rect 1150 674 1156 675
rect 255 659 264 660
rect 255 655 256 659
rect 263 655 264 659
rect 255 654 264 655
rect 430 659 437 660
rect 430 655 431 659
rect 436 655 437 659
rect 430 654 437 655
rect 583 659 589 660
rect 583 655 584 659
rect 588 658 589 659
rect 623 659 629 660
rect 623 658 624 659
rect 588 656 624 658
rect 588 655 589 656
rect 583 654 589 655
rect 623 655 624 656
rect 628 655 629 659
rect 623 654 629 655
rect 807 659 816 660
rect 807 655 808 659
rect 815 655 816 659
rect 807 654 816 655
rect 983 659 992 660
rect 983 655 984 659
rect 991 655 992 659
rect 983 654 992 655
rect 1150 659 1157 660
rect 1150 655 1151 659
rect 1156 655 1157 659
rect 1150 654 1157 655
rect 1311 659 1317 660
rect 1311 655 1312 659
rect 1316 658 1317 659
rect 1319 659 1325 660
rect 1319 658 1320 659
rect 1316 656 1320 658
rect 1316 655 1317 656
rect 1311 654 1317 655
rect 1319 655 1320 656
rect 1324 655 1325 659
rect 1319 654 1325 655
rect 1463 659 1469 660
rect 1463 655 1464 659
rect 1468 658 1469 659
rect 1471 659 1477 660
rect 1471 658 1472 659
rect 1468 656 1472 658
rect 1468 655 1469 656
rect 1463 654 1469 655
rect 1471 655 1472 656
rect 1476 655 1477 659
rect 1471 654 1477 655
rect 1615 659 1621 660
rect 1615 655 1616 659
rect 1620 658 1621 659
rect 1639 659 1645 660
rect 1639 658 1640 659
rect 1620 656 1640 658
rect 1620 655 1621 656
rect 1615 654 1621 655
rect 1639 655 1640 656
rect 1644 655 1645 659
rect 1639 654 1645 655
rect 1775 659 1781 660
rect 1775 655 1776 659
rect 1780 658 1781 659
rect 1783 659 1789 660
rect 1783 658 1784 659
rect 1780 656 1784 658
rect 1780 655 1781 656
rect 1775 654 1781 655
rect 1783 655 1784 656
rect 1788 655 1789 659
rect 1783 654 1789 655
rect 1910 659 1917 660
rect 1910 655 1911 659
rect 1916 655 1917 659
rect 1910 654 1917 655
rect 4218 659 4224 660
rect 4218 655 4219 659
rect 4223 658 4224 659
rect 4223 656 4410 658
rect 4223 655 4224 656
rect 4218 654 4224 655
rect 110 652 116 653
rect 1934 652 1940 653
rect 110 648 111 652
rect 115 648 116 652
rect 110 647 116 648
rect 130 651 136 652
rect 130 647 131 651
rect 135 647 136 651
rect 130 646 136 647
rect 306 651 312 652
rect 306 647 307 651
rect 311 647 312 651
rect 306 646 312 647
rect 498 651 504 652
rect 498 647 499 651
rect 503 647 504 651
rect 498 646 504 647
rect 682 651 688 652
rect 682 647 683 651
rect 687 647 688 651
rect 682 646 688 647
rect 858 651 864 652
rect 858 647 859 651
rect 863 647 864 651
rect 858 646 864 647
rect 1026 651 1032 652
rect 1026 647 1027 651
rect 1031 647 1032 651
rect 1026 646 1032 647
rect 1186 651 1192 652
rect 1186 647 1187 651
rect 1191 647 1192 651
rect 1186 646 1192 647
rect 1338 651 1344 652
rect 1338 647 1339 651
rect 1343 647 1344 651
rect 1338 646 1344 647
rect 1490 651 1496 652
rect 1490 647 1491 651
rect 1495 647 1496 651
rect 1490 646 1496 647
rect 1650 651 1656 652
rect 1650 647 1651 651
rect 1655 647 1656 651
rect 1650 646 1656 647
rect 1786 651 1792 652
rect 1786 647 1787 651
rect 1791 647 1792 651
rect 1934 648 1935 652
rect 1939 648 1940 652
rect 1934 647 1940 648
rect 3866 651 3872 652
rect 3866 647 3867 651
rect 3871 650 3872 651
rect 3983 651 3989 652
rect 3983 650 3984 651
rect 3871 648 3984 650
rect 3871 647 3872 648
rect 1786 646 1792 647
rect 3866 646 3872 647
rect 3983 647 3984 648
rect 3988 647 3989 651
rect 3983 646 3989 647
rect 4119 651 4125 652
rect 4119 647 4120 651
rect 4124 650 4125 651
rect 4127 651 4133 652
rect 4127 650 4128 651
rect 4124 648 4128 650
rect 4124 647 4125 648
rect 4119 646 4125 647
rect 4127 647 4128 648
rect 4132 647 4133 651
rect 4127 646 4133 647
rect 4255 651 4261 652
rect 4255 647 4256 651
rect 4260 650 4261 651
rect 4263 651 4269 652
rect 4263 650 4264 651
rect 4260 648 4264 650
rect 4260 647 4261 648
rect 4255 646 4261 647
rect 4263 647 4264 648
rect 4268 647 4269 651
rect 4263 646 4269 647
rect 4391 651 4397 652
rect 4391 647 4392 651
rect 4396 650 4397 651
rect 4399 651 4405 652
rect 4399 650 4400 651
rect 4396 648 4400 650
rect 4396 647 4397 648
rect 4391 646 4397 647
rect 4399 647 4400 648
rect 4404 647 4405 651
rect 4408 650 4410 656
rect 4527 651 4533 652
rect 4527 650 4528 651
rect 4408 648 4528 650
rect 4399 646 4405 647
rect 4527 647 4528 648
rect 4532 647 4533 651
rect 4527 646 4533 647
rect 4695 651 4704 652
rect 4695 647 4696 651
rect 4703 647 4704 651
rect 4695 646 4704 647
rect 4895 651 4904 652
rect 4895 647 4896 651
rect 4903 647 4904 651
rect 4895 646 4904 647
rect 5119 651 5128 652
rect 5119 647 5120 651
rect 5127 647 5128 651
rect 5119 646 5128 647
rect 5334 651 5340 652
rect 5334 647 5335 651
rect 5339 650 5340 651
rect 5351 651 5357 652
rect 5351 650 5352 651
rect 5339 648 5352 650
rect 5339 647 5340 648
rect 5334 646 5340 647
rect 5351 647 5352 648
rect 5356 647 5357 651
rect 5351 646 5357 647
rect 5583 651 5589 652
rect 5583 647 5584 651
rect 5588 650 5589 651
rect 5594 651 5600 652
rect 5594 650 5595 651
rect 5588 648 5595 650
rect 5588 647 5589 648
rect 5583 646 5589 647
rect 5594 647 5595 648
rect 5599 647 5600 651
rect 5594 646 5600 647
rect 3838 644 3844 645
rect 5662 644 5668 645
rect 3838 640 3839 644
rect 3843 640 3844 644
rect 3838 639 3844 640
rect 3858 643 3864 644
rect 3858 639 3859 643
rect 3863 639 3864 643
rect 3858 638 3864 639
rect 3994 643 4000 644
rect 3994 639 3995 643
rect 3999 639 4000 643
rect 3994 638 4000 639
rect 4130 643 4136 644
rect 4130 639 4131 643
rect 4135 639 4136 643
rect 4130 638 4136 639
rect 4266 643 4272 644
rect 4266 639 4267 643
rect 4271 639 4272 643
rect 4266 638 4272 639
rect 4402 643 4408 644
rect 4402 639 4403 643
rect 4407 639 4408 643
rect 4402 638 4408 639
rect 4570 643 4576 644
rect 4570 639 4571 643
rect 4575 639 4576 643
rect 4570 638 4576 639
rect 4770 643 4776 644
rect 4770 639 4771 643
rect 4775 639 4776 643
rect 4770 638 4776 639
rect 4994 643 5000 644
rect 4994 639 4995 643
rect 4999 639 5000 643
rect 4994 638 5000 639
rect 5226 643 5232 644
rect 5226 639 5227 643
rect 5231 639 5232 643
rect 5226 638 5232 639
rect 5458 643 5464 644
rect 5458 639 5459 643
rect 5463 639 5464 643
rect 5662 640 5663 644
rect 5667 640 5668 644
rect 5662 639 5668 640
rect 5458 638 5464 639
rect 158 636 164 637
rect 110 635 116 636
rect 110 631 111 635
rect 115 631 116 635
rect 158 632 159 636
rect 163 632 164 636
rect 158 631 164 632
rect 334 636 340 637
rect 334 632 335 636
rect 339 632 340 636
rect 334 631 340 632
rect 526 636 532 637
rect 526 632 527 636
rect 531 632 532 636
rect 526 631 532 632
rect 710 636 716 637
rect 710 632 711 636
rect 715 632 716 636
rect 710 631 716 632
rect 886 636 892 637
rect 886 632 887 636
rect 891 632 892 636
rect 886 631 892 632
rect 1054 636 1060 637
rect 1054 632 1055 636
rect 1059 632 1060 636
rect 1054 631 1060 632
rect 1214 636 1220 637
rect 1214 632 1215 636
rect 1219 632 1220 636
rect 1214 631 1220 632
rect 1366 636 1372 637
rect 1366 632 1367 636
rect 1371 632 1372 636
rect 1366 631 1372 632
rect 1518 636 1524 637
rect 1518 632 1519 636
rect 1523 632 1524 636
rect 1518 631 1524 632
rect 1678 636 1684 637
rect 1678 632 1679 636
rect 1683 632 1684 636
rect 1678 631 1684 632
rect 1814 636 1820 637
rect 1814 632 1815 636
rect 1819 632 1820 636
rect 1814 631 1820 632
rect 1934 635 1940 636
rect 1934 631 1935 635
rect 1939 631 1940 635
rect 110 630 116 631
rect 1934 630 1940 631
rect 3886 628 3892 629
rect 3838 627 3844 628
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3886 624 3887 628
rect 3891 624 3892 628
rect 3886 623 3892 624
rect 4022 628 4028 629
rect 4022 624 4023 628
rect 4027 624 4028 628
rect 4022 623 4028 624
rect 4158 628 4164 629
rect 4158 624 4159 628
rect 4163 624 4164 628
rect 4158 623 4164 624
rect 4294 628 4300 629
rect 4294 624 4295 628
rect 4299 624 4300 628
rect 4294 623 4300 624
rect 4430 628 4436 629
rect 4430 624 4431 628
rect 4435 624 4436 628
rect 4430 623 4436 624
rect 4598 628 4604 629
rect 4598 624 4599 628
rect 4603 624 4604 628
rect 4598 623 4604 624
rect 4798 628 4804 629
rect 4798 624 4799 628
rect 4803 624 4804 628
rect 4798 623 4804 624
rect 5022 628 5028 629
rect 5022 624 5023 628
rect 5027 624 5028 628
rect 5022 623 5028 624
rect 5254 628 5260 629
rect 5254 624 5255 628
rect 5259 624 5260 628
rect 5254 623 5260 624
rect 5486 628 5492 629
rect 5486 624 5487 628
rect 5491 624 5492 628
rect 5486 623 5492 624
rect 5662 627 5668 628
rect 5662 623 5663 627
rect 5667 623 5668 627
rect 3838 622 3844 623
rect 5662 622 5668 623
rect 4407 611 4413 612
rect 4407 607 4408 611
rect 4412 610 4413 611
rect 5334 611 5340 612
rect 5334 610 5335 611
rect 4412 608 5335 610
rect 4412 607 4413 608
rect 4407 606 4413 607
rect 5334 607 5335 608
rect 5339 607 5340 611
rect 5334 606 5340 607
rect 110 577 116 578
rect 1934 577 1940 578
rect 110 573 111 577
rect 115 573 116 577
rect 110 572 116 573
rect 158 576 164 577
rect 158 572 159 576
rect 163 572 164 576
rect 158 571 164 572
rect 374 576 380 577
rect 374 572 375 576
rect 379 572 380 576
rect 374 571 380 572
rect 598 576 604 577
rect 598 572 599 576
rect 603 572 604 576
rect 598 571 604 572
rect 806 576 812 577
rect 806 572 807 576
rect 811 572 812 576
rect 806 571 812 572
rect 998 576 1004 577
rect 998 572 999 576
rect 1003 572 1004 576
rect 998 571 1004 572
rect 1174 576 1180 577
rect 1174 572 1175 576
rect 1179 572 1180 576
rect 1174 571 1180 572
rect 1342 576 1348 577
rect 1342 572 1343 576
rect 1347 572 1348 576
rect 1342 571 1348 572
rect 1510 576 1516 577
rect 1510 572 1511 576
rect 1515 572 1516 576
rect 1510 571 1516 572
rect 1670 576 1676 577
rect 1670 572 1671 576
rect 1675 572 1676 576
rect 1670 571 1676 572
rect 1814 576 1820 577
rect 1814 572 1815 576
rect 1819 572 1820 576
rect 1934 573 1935 577
rect 1939 573 1940 577
rect 1934 572 1940 573
rect 1814 571 1820 572
rect 3838 569 3844 570
rect 5662 569 5668 570
rect 3838 565 3839 569
rect 3843 565 3844 569
rect 3838 564 3844 565
rect 3886 568 3892 569
rect 3886 564 3887 568
rect 3891 564 3892 568
rect 3886 563 3892 564
rect 4022 568 4028 569
rect 4022 564 4023 568
rect 4027 564 4028 568
rect 4022 563 4028 564
rect 4158 568 4164 569
rect 4158 564 4159 568
rect 4163 564 4164 568
rect 4158 563 4164 564
rect 4294 568 4300 569
rect 4294 564 4295 568
rect 4299 564 4300 568
rect 4294 563 4300 564
rect 4478 568 4484 569
rect 4478 564 4479 568
rect 4483 564 4484 568
rect 4478 563 4484 564
rect 4694 568 4700 569
rect 4694 564 4695 568
rect 4699 564 4700 568
rect 4694 563 4700 564
rect 4934 568 4940 569
rect 4934 564 4935 568
rect 4939 564 4940 568
rect 4934 563 4940 564
rect 5190 568 5196 569
rect 5190 564 5191 568
rect 5195 564 5196 568
rect 5190 563 5196 564
rect 5446 568 5452 569
rect 5446 564 5447 568
rect 5451 564 5452 568
rect 5662 565 5663 569
rect 5667 565 5668 569
rect 5662 564 5668 565
rect 5446 563 5452 564
rect 130 561 136 562
rect 110 560 116 561
rect 110 556 111 560
rect 115 556 116 560
rect 130 557 131 561
rect 135 557 136 561
rect 130 556 136 557
rect 346 561 352 562
rect 346 557 347 561
rect 351 557 352 561
rect 346 556 352 557
rect 570 561 576 562
rect 570 557 571 561
rect 575 557 576 561
rect 570 556 576 557
rect 778 561 784 562
rect 778 557 779 561
rect 783 557 784 561
rect 778 556 784 557
rect 970 561 976 562
rect 970 557 971 561
rect 975 557 976 561
rect 970 556 976 557
rect 1146 561 1152 562
rect 1146 557 1147 561
rect 1151 557 1152 561
rect 1146 556 1152 557
rect 1314 561 1320 562
rect 1314 557 1315 561
rect 1319 557 1320 561
rect 1314 556 1320 557
rect 1482 561 1488 562
rect 1482 557 1483 561
rect 1487 557 1488 561
rect 1482 556 1488 557
rect 1642 561 1648 562
rect 1642 557 1643 561
rect 1647 557 1648 561
rect 1642 556 1648 557
rect 1786 561 1792 562
rect 1786 557 1787 561
rect 1791 557 1792 561
rect 1786 556 1792 557
rect 1934 560 1940 561
rect 1934 556 1935 560
rect 1939 556 1940 560
rect 110 555 116 556
rect 1934 555 1940 556
rect 3858 553 3864 554
rect 3838 552 3844 553
rect 255 551 261 552
rect 255 547 256 551
rect 260 550 261 551
rect 362 551 368 552
rect 362 550 363 551
rect 260 548 363 550
rect 260 547 261 548
rect 255 546 261 547
rect 362 547 363 548
rect 367 547 368 551
rect 362 546 368 547
rect 471 551 480 552
rect 471 547 472 551
rect 479 547 480 551
rect 471 546 480 547
rect 695 551 704 552
rect 695 547 696 551
rect 703 547 704 551
rect 695 546 704 547
rect 759 551 765 552
rect 759 547 760 551
rect 764 550 765 551
rect 903 551 909 552
rect 903 550 904 551
rect 764 548 904 550
rect 764 547 765 548
rect 759 546 765 547
rect 903 547 904 548
rect 908 547 909 551
rect 903 546 909 547
rect 943 551 949 552
rect 943 547 944 551
rect 948 550 949 551
rect 1095 551 1101 552
rect 1095 550 1096 551
rect 948 548 1096 550
rect 948 547 949 548
rect 943 546 949 547
rect 1095 547 1096 548
rect 1100 547 1101 551
rect 1095 546 1101 547
rect 1271 551 1280 552
rect 1271 547 1272 551
rect 1279 547 1280 551
rect 1271 546 1280 547
rect 1302 551 1308 552
rect 1302 547 1303 551
rect 1307 550 1308 551
rect 1439 551 1445 552
rect 1439 550 1440 551
rect 1307 548 1440 550
rect 1307 547 1308 548
rect 1302 546 1308 547
rect 1439 547 1440 548
rect 1444 547 1445 551
rect 1439 546 1445 547
rect 1490 551 1496 552
rect 1490 547 1491 551
rect 1495 550 1496 551
rect 1607 551 1613 552
rect 1607 550 1608 551
rect 1495 548 1608 550
rect 1495 547 1496 548
rect 1490 546 1496 547
rect 1607 547 1608 548
rect 1612 547 1613 551
rect 1607 546 1613 547
rect 1631 551 1637 552
rect 1631 547 1632 551
rect 1636 550 1637 551
rect 1767 551 1773 552
rect 1767 550 1768 551
rect 1636 548 1768 550
rect 1636 547 1637 548
rect 1631 546 1637 547
rect 1767 547 1768 548
rect 1772 547 1773 551
rect 1767 546 1773 547
rect 1778 551 1784 552
rect 1778 547 1779 551
rect 1783 550 1784 551
rect 1911 551 1917 552
rect 1911 550 1912 551
rect 1783 548 1912 550
rect 1783 547 1784 548
rect 1778 546 1784 547
rect 1911 547 1912 548
rect 1916 547 1917 551
rect 1911 546 1917 547
rect 1974 549 1980 550
rect 3798 549 3804 550
rect 1974 545 1975 549
rect 1979 545 1980 549
rect 1974 544 1980 545
rect 3310 548 3316 549
rect 3310 544 3311 548
rect 3315 544 3316 548
rect 3310 543 3316 544
rect 3446 548 3452 549
rect 3446 544 3447 548
rect 3451 544 3452 548
rect 3446 543 3452 544
rect 3582 548 3588 549
rect 3582 544 3583 548
rect 3587 544 3588 548
rect 3798 545 3799 549
rect 3803 545 3804 549
rect 3838 548 3839 552
rect 3843 548 3844 552
rect 3858 549 3859 553
rect 3863 549 3864 553
rect 3858 548 3864 549
rect 3994 553 4000 554
rect 3994 549 3995 553
rect 3999 549 4000 553
rect 3994 548 4000 549
rect 4130 553 4136 554
rect 4130 549 4131 553
rect 4135 549 4136 553
rect 4130 548 4136 549
rect 4266 553 4272 554
rect 4266 549 4267 553
rect 4271 549 4272 553
rect 4266 548 4272 549
rect 4450 553 4456 554
rect 4450 549 4451 553
rect 4455 549 4456 553
rect 4450 548 4456 549
rect 4666 553 4672 554
rect 4666 549 4667 553
rect 4671 549 4672 553
rect 4666 548 4672 549
rect 4906 553 4912 554
rect 4906 549 4907 553
rect 4911 549 4912 553
rect 4906 548 4912 549
rect 5162 553 5168 554
rect 5162 549 5163 553
rect 5167 549 5168 553
rect 5162 548 5168 549
rect 5418 553 5424 554
rect 5418 549 5419 553
rect 5423 549 5424 553
rect 5418 548 5424 549
rect 5662 552 5668 553
rect 5662 548 5663 552
rect 5667 548 5668 552
rect 3838 547 3844 548
rect 5662 547 5668 548
rect 3798 544 3804 545
rect 3582 543 3588 544
rect 3946 543 3952 544
rect 3946 539 3947 543
rect 3951 542 3952 543
rect 3983 543 3989 544
rect 3983 542 3984 543
rect 3951 540 3984 542
rect 3951 539 3952 540
rect 3946 538 3952 539
rect 3983 539 3984 540
rect 3988 539 3989 543
rect 3983 538 3989 539
rect 4002 543 4008 544
rect 4002 539 4003 543
rect 4007 542 4008 543
rect 4119 543 4125 544
rect 4119 542 4120 543
rect 4007 540 4120 542
rect 4007 539 4008 540
rect 4002 538 4008 539
rect 4119 539 4120 540
rect 4124 539 4125 543
rect 4119 538 4125 539
rect 4127 543 4133 544
rect 4127 539 4128 543
rect 4132 542 4133 543
rect 4255 543 4261 544
rect 4255 542 4256 543
rect 4132 540 4256 542
rect 4132 539 4133 540
rect 4127 538 4133 539
rect 4255 539 4256 540
rect 4260 539 4261 543
rect 4255 538 4261 539
rect 4391 543 4397 544
rect 4391 539 4392 543
rect 4396 542 4397 543
rect 4466 543 4472 544
rect 4466 542 4467 543
rect 4396 540 4467 542
rect 4396 539 4397 540
rect 4391 538 4397 539
rect 4466 539 4467 540
rect 4471 539 4472 543
rect 4466 538 4472 539
rect 4575 543 4581 544
rect 4575 539 4576 543
rect 4580 542 4581 543
rect 4682 543 4688 544
rect 4682 542 4683 543
rect 4580 540 4683 542
rect 4580 539 4581 540
rect 4575 538 4581 539
rect 4682 539 4683 540
rect 4687 539 4688 543
rect 4682 538 4688 539
rect 4791 543 4797 544
rect 4791 539 4792 543
rect 4796 542 4797 543
rect 4922 543 4928 544
rect 4922 542 4923 543
rect 4796 540 4923 542
rect 4796 539 4797 540
rect 4791 538 4797 539
rect 4922 539 4923 540
rect 4927 539 4928 543
rect 4922 538 4928 539
rect 5031 543 5037 544
rect 5031 539 5032 543
rect 5036 542 5037 543
rect 5178 543 5184 544
rect 5178 542 5179 543
rect 5036 540 5179 542
rect 5036 539 5037 540
rect 5031 538 5037 539
rect 5178 539 5179 540
rect 5183 539 5184 543
rect 5178 538 5184 539
rect 5186 543 5192 544
rect 5186 539 5187 543
rect 5191 542 5192 543
rect 5287 543 5293 544
rect 5287 542 5288 543
rect 5191 540 5288 542
rect 5191 539 5192 540
rect 5186 538 5192 539
rect 5287 539 5288 540
rect 5292 539 5293 543
rect 5287 538 5293 539
rect 5543 543 5552 544
rect 5543 539 5544 543
rect 5551 539 5552 543
rect 5543 538 5552 539
rect 3282 533 3288 534
rect 1974 532 1980 533
rect 1974 528 1975 532
rect 1979 528 1980 532
rect 3282 529 3283 533
rect 3287 529 3288 533
rect 3282 528 3288 529
rect 3418 533 3424 534
rect 3418 529 3419 533
rect 3423 529 3424 533
rect 3418 528 3424 529
rect 3554 533 3560 534
rect 3554 529 3555 533
rect 3559 529 3560 533
rect 3554 528 3560 529
rect 3798 532 3804 533
rect 3798 528 3799 532
rect 3803 528 3804 532
rect 1974 527 1980 528
rect 3798 527 3804 528
rect 3407 523 3413 524
rect 226 519 232 520
rect 226 518 227 519
rect 221 516 227 518
rect 226 515 227 516
rect 231 515 232 519
rect 226 514 232 515
rect 362 519 368 520
rect 362 515 363 519
rect 367 515 368 519
rect 759 519 765 520
rect 759 518 760 519
rect 661 516 760 518
rect 362 514 368 515
rect 759 515 760 516
rect 764 515 765 519
rect 943 519 949 520
rect 943 518 944 519
rect 869 516 944 518
rect 759 514 765 515
rect 943 515 944 516
rect 948 515 949 519
rect 943 514 949 515
rect 986 519 992 520
rect 986 515 987 519
rect 991 515 992 519
rect 1302 519 1308 520
rect 1302 518 1303 519
rect 1237 516 1303 518
rect 986 514 992 515
rect 1302 515 1303 516
rect 1307 515 1308 519
rect 1490 519 1496 520
rect 1490 518 1491 519
rect 1405 516 1491 518
rect 1302 514 1308 515
rect 1490 515 1491 516
rect 1495 515 1496 519
rect 1631 519 1637 520
rect 1631 518 1632 519
rect 1573 516 1632 518
rect 1490 514 1496 515
rect 1631 515 1632 516
rect 1636 515 1637 519
rect 1778 519 1784 520
rect 1778 518 1779 519
rect 1733 516 1779 518
rect 1631 514 1637 515
rect 1778 515 1779 516
rect 1783 515 1784 519
rect 1882 519 1888 520
rect 1882 518 1883 519
rect 1877 516 1883 518
rect 1778 514 1784 515
rect 1882 515 1883 516
rect 1887 515 1888 519
rect 3407 519 3408 523
rect 3412 522 3413 523
rect 3434 523 3440 524
rect 3434 522 3435 523
rect 3412 520 3435 522
rect 3412 519 3413 520
rect 3407 518 3413 519
rect 3434 519 3435 520
rect 3439 519 3440 523
rect 3434 518 3440 519
rect 3543 523 3549 524
rect 3543 519 3544 523
rect 3548 522 3549 523
rect 3570 523 3576 524
rect 3570 522 3571 523
rect 3548 520 3571 522
rect 3548 519 3549 520
rect 3543 518 3549 519
rect 3570 519 3571 520
rect 3575 519 3576 523
rect 3570 518 3576 519
rect 3642 523 3648 524
rect 3642 519 3643 523
rect 3647 522 3648 523
rect 3679 523 3685 524
rect 3679 522 3680 523
rect 3647 520 3680 522
rect 3647 519 3648 520
rect 3642 518 3648 519
rect 3679 519 3680 520
rect 3684 519 3685 523
rect 3679 518 3685 519
rect 1882 514 1888 515
rect 4002 511 4008 512
rect 4002 510 4003 511
rect 3949 508 4003 510
rect 4002 507 4003 508
rect 4007 507 4008 511
rect 4127 511 4133 512
rect 4127 510 4128 511
rect 4085 508 4128 510
rect 4002 506 4008 507
rect 4127 507 4128 508
rect 4132 507 4133 511
rect 4127 506 4133 507
rect 4218 511 4224 512
rect 4218 507 4219 511
rect 4223 507 4224 511
rect 4407 511 4413 512
rect 4407 510 4408 511
rect 4357 508 4408 510
rect 4218 506 4224 507
rect 4407 507 4408 508
rect 4412 507 4413 511
rect 4407 506 4413 507
rect 4466 511 4472 512
rect 4466 507 4467 511
rect 4471 507 4472 511
rect 4466 506 4472 507
rect 4682 511 4688 512
rect 4682 507 4683 511
rect 4687 507 4688 511
rect 4682 506 4688 507
rect 4922 511 4928 512
rect 4922 507 4923 511
rect 4927 507 4928 511
rect 4922 506 4928 507
rect 5178 511 5184 512
rect 5178 507 5179 511
rect 5183 507 5184 511
rect 5178 506 5184 507
rect 5434 511 5440 512
rect 5434 507 5435 511
rect 5439 507 5440 511
rect 5434 506 5440 507
rect 4570 495 4576 496
rect 3298 491 3304 492
rect 3298 487 3299 491
rect 3303 487 3304 491
rect 3298 486 3304 487
rect 3434 491 3440 492
rect 3434 487 3435 491
rect 3439 487 3440 491
rect 3434 486 3440 487
rect 3570 491 3576 492
rect 3570 487 3571 491
rect 3575 487 3576 491
rect 4570 491 4571 495
rect 4575 494 4576 495
rect 5186 495 5192 496
rect 5186 494 5187 495
rect 4575 492 5187 494
rect 4575 491 4576 492
rect 4570 490 4576 491
rect 5186 491 5187 492
rect 5191 491 5192 495
rect 5186 490 5192 491
rect 3570 486 3576 487
rect 350 471 356 472
rect 350 470 351 471
rect 221 468 351 470
rect 350 467 351 468
rect 355 467 356 471
rect 558 471 564 472
rect 558 470 559 471
rect 517 468 559 470
rect 350 466 356 467
rect 558 467 559 468
rect 563 467 564 471
rect 558 466 564 467
rect 698 471 704 472
rect 698 467 699 471
rect 703 470 704 471
rect 890 471 896 472
rect 703 468 781 470
rect 703 467 704 468
rect 698 466 704 467
rect 890 467 891 471
rect 895 470 896 471
rect 1234 471 1240 472
rect 895 468 1125 470
rect 895 467 896 468
rect 890 466 896 467
rect 1234 467 1235 471
rect 1239 470 1240 471
rect 1959 471 1965 472
rect 1959 470 1960 471
rect 1239 468 1477 470
rect 1877 468 1960 470
rect 1239 467 1240 468
rect 1234 466 1240 467
rect 1959 467 1960 468
rect 1964 467 1965 471
rect 1959 466 1965 467
rect 4570 451 4576 452
rect 4570 450 4571 451
rect 4541 448 4571 450
rect 4570 447 4571 448
rect 4575 447 4576 451
rect 4570 446 4576 447
rect 4578 451 4584 452
rect 4578 447 4579 451
rect 4583 450 4584 451
rect 4778 451 4784 452
rect 4583 448 4669 450
rect 4583 447 4584 448
rect 4578 446 4584 447
rect 4778 447 4779 451
rect 4783 450 4784 451
rect 4986 451 4992 452
rect 4783 448 4877 450
rect 4783 447 4784 448
rect 4778 446 4784 447
rect 4986 447 4987 451
rect 4991 450 4992 451
rect 4991 448 5085 450
rect 4991 447 4992 448
rect 4986 446 4992 447
rect 5594 447 5600 448
rect 2143 443 2149 444
rect 2143 442 2144 443
rect 2085 440 2144 442
rect 2143 439 2144 440
rect 2148 439 2149 443
rect 2143 438 2149 439
rect 2258 443 2264 444
rect 2258 439 2259 443
rect 2263 442 2264 443
rect 2474 443 2480 444
rect 2263 440 2365 442
rect 2263 439 2264 440
rect 2258 438 2264 439
rect 2474 439 2475 443
rect 2479 442 2480 443
rect 2666 443 2672 444
rect 2479 440 2557 442
rect 2479 439 2480 440
rect 2474 438 2480 439
rect 2666 439 2667 443
rect 2671 442 2672 443
rect 3050 443 3056 444
rect 2671 440 2749 442
rect 2671 439 2672 440
rect 2666 438 2672 439
rect 3010 439 3016 440
rect 226 435 232 436
rect 226 431 227 435
rect 231 434 232 435
rect 255 435 261 436
rect 255 434 256 435
rect 231 432 256 434
rect 231 431 232 432
rect 226 430 232 431
rect 255 431 256 432
rect 260 431 261 435
rect 255 430 261 431
rect 350 435 356 436
rect 350 431 351 435
rect 355 434 356 435
rect 551 435 557 436
rect 551 434 552 435
rect 355 432 552 434
rect 355 431 356 432
rect 350 430 356 431
rect 551 431 552 432
rect 556 431 557 435
rect 551 430 557 431
rect 887 435 896 436
rect 887 431 888 435
rect 895 431 896 435
rect 887 430 896 431
rect 1231 435 1240 436
rect 1231 431 1232 435
rect 1239 431 1240 435
rect 1231 430 1240 431
rect 1518 435 1524 436
rect 1518 431 1519 435
rect 1523 434 1524 435
rect 1583 435 1589 436
rect 1583 434 1584 435
rect 1523 432 1584 434
rect 1523 431 1524 432
rect 1518 430 1524 431
rect 1583 431 1584 432
rect 1588 431 1589 435
rect 1583 430 1589 431
rect 1882 435 1888 436
rect 1882 431 1883 435
rect 1887 434 1888 435
rect 1911 435 1917 436
rect 1911 434 1912 435
rect 1887 432 1912 434
rect 1887 431 1888 432
rect 1882 430 1888 431
rect 1911 431 1912 432
rect 1916 431 1917 435
rect 2240 434 2242 437
rect 3010 435 3011 439
rect 3015 435 3016 439
rect 3050 439 3051 443
rect 3055 442 3056 443
rect 3242 443 3248 444
rect 3055 440 3133 442
rect 3055 439 3056 440
rect 3050 438 3056 439
rect 3242 439 3243 443
rect 3247 442 3248 443
rect 3634 443 3640 444
rect 3634 442 3635 443
rect 3247 440 3317 442
rect 3573 440 3635 442
rect 3247 439 3248 440
rect 3242 438 3248 439
rect 3634 439 3635 440
rect 3639 439 3640 443
rect 3634 438 3640 439
rect 3642 443 3648 444
rect 3642 439 3643 443
rect 3647 442 3648 443
rect 3647 440 3669 442
rect 5368 440 5370 445
rect 5594 443 5595 447
rect 5599 443 5600 447
rect 5594 442 5600 443
rect 3647 439 3648 440
rect 3642 438 3648 439
rect 5367 439 5373 440
rect 3010 434 3016 435
rect 5367 435 5368 439
rect 5372 435 5373 439
rect 5367 434 5373 435
rect 2240 432 2301 434
rect 1911 430 1917 431
rect 110 428 116 429
rect 1934 428 1940 429
rect 110 424 111 428
rect 115 424 116 428
rect 110 423 116 424
rect 130 427 136 428
rect 130 423 131 427
rect 135 423 136 427
rect 130 422 136 423
rect 426 427 432 428
rect 426 423 427 427
rect 431 423 432 427
rect 426 422 432 423
rect 762 427 768 428
rect 762 423 763 427
rect 767 423 768 427
rect 762 422 768 423
rect 1106 427 1112 428
rect 1106 423 1107 427
rect 1111 423 1112 427
rect 1106 422 1112 423
rect 1458 427 1464 428
rect 1458 423 1459 427
rect 1463 423 1464 427
rect 1458 422 1464 423
rect 1786 427 1792 428
rect 1786 423 1787 427
rect 1791 423 1792 427
rect 1934 424 1935 428
rect 1939 424 1940 428
rect 2299 426 2301 432
rect 2854 427 2860 428
rect 2854 426 2855 427
rect 2299 424 2855 426
rect 1934 423 1940 424
rect 2854 423 2855 424
rect 2859 423 2860 427
rect 1786 422 1792 423
rect 2854 422 2860 423
rect 3010 415 3016 416
rect 158 412 164 413
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 158 408 159 412
rect 163 408 164 412
rect 158 407 164 408
rect 454 412 460 413
rect 454 408 455 412
rect 459 408 460 412
rect 454 407 460 408
rect 790 412 796 413
rect 790 408 791 412
rect 795 408 796 412
rect 790 407 796 408
rect 1134 412 1140 413
rect 1134 408 1135 412
rect 1139 408 1140 412
rect 1134 407 1140 408
rect 1486 412 1492 413
rect 1486 408 1487 412
rect 1491 408 1492 412
rect 1486 407 1492 408
rect 1814 412 1820 413
rect 1814 408 1815 412
rect 1819 408 1820 412
rect 1814 407 1820 408
rect 1934 411 1940 412
rect 1934 407 1935 411
rect 1939 407 1940 411
rect 3010 411 3011 415
rect 3015 414 3016 415
rect 4575 415 4584 416
rect 3015 412 3434 414
rect 3015 411 3016 412
rect 3010 410 3016 411
rect 110 406 116 407
rect 1934 406 1940 407
rect 1959 407 1965 408
rect 1959 403 1960 407
rect 1964 406 1965 407
rect 2119 407 2125 408
rect 2119 406 2120 407
rect 1964 404 2120 406
rect 1964 403 1965 404
rect 1959 402 1965 403
rect 2119 403 2120 404
rect 2124 403 2125 407
rect 2119 402 2125 403
rect 2143 407 2149 408
rect 2143 403 2144 407
rect 2148 406 2149 407
rect 2279 407 2285 408
rect 2279 406 2280 407
rect 2148 404 2280 406
rect 2148 403 2149 404
rect 2143 402 2149 403
rect 2279 403 2280 404
rect 2284 403 2285 407
rect 2279 402 2285 403
rect 2471 407 2480 408
rect 2471 403 2472 407
rect 2479 403 2480 407
rect 2471 402 2480 403
rect 2663 407 2672 408
rect 2663 403 2664 407
rect 2671 403 2672 407
rect 2663 402 2672 403
rect 2854 407 2861 408
rect 2854 403 2855 407
rect 2860 403 2861 407
rect 2854 402 2861 403
rect 3047 407 3056 408
rect 3047 403 3048 407
rect 3055 403 3056 407
rect 3047 402 3056 403
rect 3239 407 3248 408
rect 3239 403 3240 407
rect 3247 403 3248 407
rect 3239 402 3248 403
rect 3422 407 3429 408
rect 3422 403 3423 407
rect 3428 403 3429 407
rect 3432 406 3434 412
rect 4575 411 4576 415
rect 4583 411 4584 415
rect 4575 410 4584 411
rect 4775 415 4784 416
rect 4775 411 4776 415
rect 4783 411 4784 415
rect 4775 410 4784 411
rect 4983 415 4992 416
rect 4983 411 4984 415
rect 4991 411 4992 415
rect 4983 410 4992 411
rect 5034 415 5040 416
rect 5034 411 5035 415
rect 5039 414 5040 415
rect 5191 415 5197 416
rect 5191 414 5192 415
rect 5039 412 5192 414
rect 5039 411 5040 412
rect 5034 410 5040 411
rect 5191 411 5192 412
rect 5196 411 5197 415
rect 5191 410 5197 411
rect 5407 415 5413 416
rect 5407 411 5408 415
rect 5412 414 5413 415
rect 5434 415 5440 416
rect 5434 414 5435 415
rect 5412 412 5435 414
rect 5412 411 5413 412
rect 5407 410 5413 411
rect 5434 411 5435 412
rect 5439 411 5440 415
rect 5434 410 5440 411
rect 5602 415 5608 416
rect 5602 411 5603 415
rect 5607 414 5608 415
rect 5631 415 5637 416
rect 5631 414 5632 415
rect 5607 412 5632 414
rect 5607 411 5608 412
rect 5602 410 5608 411
rect 5631 411 5632 412
rect 5636 411 5637 415
rect 5631 410 5637 411
rect 3838 408 3844 409
rect 5662 408 5668 409
rect 3607 407 3613 408
rect 3607 406 3608 407
rect 3432 404 3608 406
rect 3422 402 3429 403
rect 3607 403 3608 404
rect 3612 403 3613 407
rect 3607 402 3613 403
rect 3634 407 3640 408
rect 3634 403 3635 407
rect 3639 406 3640 407
rect 3775 407 3781 408
rect 3775 406 3776 407
rect 3639 404 3776 406
rect 3639 403 3640 404
rect 3634 402 3640 403
rect 3775 403 3776 404
rect 3780 403 3781 407
rect 3838 404 3839 408
rect 3843 404 3844 408
rect 3838 403 3844 404
rect 4450 407 4456 408
rect 4450 403 4451 407
rect 4455 403 4456 407
rect 3775 402 3781 403
rect 4450 402 4456 403
rect 4650 407 4656 408
rect 4650 403 4651 407
rect 4655 403 4656 407
rect 4650 402 4656 403
rect 4858 407 4864 408
rect 4858 403 4859 407
rect 4863 403 4864 407
rect 4858 402 4864 403
rect 5066 407 5072 408
rect 5066 403 5067 407
rect 5071 403 5072 407
rect 5066 402 5072 403
rect 5282 407 5288 408
rect 5282 403 5283 407
rect 5287 403 5288 407
rect 5282 402 5288 403
rect 5506 407 5512 408
rect 5506 403 5507 407
rect 5511 403 5512 407
rect 5662 404 5663 408
rect 5667 404 5668 408
rect 5662 403 5668 404
rect 5506 402 5512 403
rect 1974 400 1980 401
rect 3798 400 3804 401
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 1994 399 2000 400
rect 1994 395 1995 399
rect 1999 395 2000 399
rect 1994 394 2000 395
rect 2154 399 2160 400
rect 2154 395 2155 399
rect 2159 395 2160 399
rect 2154 394 2160 395
rect 2346 399 2352 400
rect 2346 395 2347 399
rect 2351 395 2352 399
rect 2346 394 2352 395
rect 2538 399 2544 400
rect 2538 395 2539 399
rect 2543 395 2544 399
rect 2538 394 2544 395
rect 2730 399 2736 400
rect 2730 395 2731 399
rect 2735 395 2736 399
rect 2730 394 2736 395
rect 2922 399 2928 400
rect 2922 395 2923 399
rect 2927 395 2928 399
rect 2922 394 2928 395
rect 3114 399 3120 400
rect 3114 395 3115 399
rect 3119 395 3120 399
rect 3114 394 3120 395
rect 3298 399 3304 400
rect 3298 395 3299 399
rect 3303 395 3304 399
rect 3298 394 3304 395
rect 3482 399 3488 400
rect 3482 395 3483 399
rect 3487 395 3488 399
rect 3482 394 3488 395
rect 3650 399 3656 400
rect 3650 395 3651 399
rect 3655 395 3656 399
rect 3798 396 3799 400
rect 3803 396 3804 400
rect 3798 395 3804 396
rect 3650 394 3656 395
rect 4478 392 4484 393
rect 3838 391 3844 392
rect 3838 387 3839 391
rect 3843 387 3844 391
rect 4478 388 4479 392
rect 4483 388 4484 392
rect 4478 387 4484 388
rect 4678 392 4684 393
rect 4678 388 4679 392
rect 4683 388 4684 392
rect 4678 387 4684 388
rect 4886 392 4892 393
rect 4886 388 4887 392
rect 4891 388 4892 392
rect 4886 387 4892 388
rect 5094 392 5100 393
rect 5094 388 5095 392
rect 5099 388 5100 392
rect 5094 387 5100 388
rect 5310 392 5316 393
rect 5310 388 5311 392
rect 5315 388 5316 392
rect 5310 387 5316 388
rect 5534 392 5540 393
rect 5534 388 5535 392
rect 5539 388 5540 392
rect 5534 387 5540 388
rect 5662 391 5668 392
rect 5662 387 5663 391
rect 5667 387 5668 391
rect 3838 386 3844 387
rect 5662 386 5668 387
rect 2022 384 2028 385
rect 1974 383 1980 384
rect 1974 379 1975 383
rect 1979 379 1980 383
rect 2022 380 2023 384
rect 2027 380 2028 384
rect 2022 379 2028 380
rect 2182 384 2188 385
rect 2182 380 2183 384
rect 2187 380 2188 384
rect 2182 379 2188 380
rect 2374 384 2380 385
rect 2374 380 2375 384
rect 2379 380 2380 384
rect 2374 379 2380 380
rect 2566 384 2572 385
rect 2566 380 2567 384
rect 2571 380 2572 384
rect 2566 379 2572 380
rect 2758 384 2764 385
rect 2758 380 2759 384
rect 2763 380 2764 384
rect 2758 379 2764 380
rect 2950 384 2956 385
rect 2950 380 2951 384
rect 2955 380 2956 384
rect 2950 379 2956 380
rect 3142 384 3148 385
rect 3142 380 3143 384
rect 3147 380 3148 384
rect 3142 379 3148 380
rect 3326 384 3332 385
rect 3326 380 3327 384
rect 3331 380 3332 384
rect 3326 379 3332 380
rect 3510 384 3516 385
rect 3510 380 3511 384
rect 3515 380 3516 384
rect 3510 379 3516 380
rect 3678 384 3684 385
rect 3678 380 3679 384
rect 3683 380 3684 384
rect 3678 379 3684 380
rect 3798 383 3804 384
rect 3798 379 3799 383
rect 3803 379 3804 383
rect 1974 378 1980 379
rect 3798 378 3804 379
rect 110 337 116 338
rect 1934 337 1940 338
rect 110 333 111 337
rect 115 333 116 337
rect 110 332 116 333
rect 238 336 244 337
rect 238 332 239 336
rect 243 332 244 336
rect 238 331 244 332
rect 390 336 396 337
rect 390 332 391 336
rect 395 332 396 336
rect 390 331 396 332
rect 550 336 556 337
rect 550 332 551 336
rect 555 332 556 336
rect 550 331 556 332
rect 710 336 716 337
rect 710 332 711 336
rect 715 332 716 336
rect 710 331 716 332
rect 870 336 876 337
rect 870 332 871 336
rect 875 332 876 336
rect 870 331 876 332
rect 1030 336 1036 337
rect 1030 332 1031 336
rect 1035 332 1036 336
rect 1934 333 1935 337
rect 1939 333 1940 337
rect 1934 332 1940 333
rect 1030 331 1036 332
rect 3838 329 3844 330
rect 5662 329 5668 330
rect 3838 325 3839 329
rect 3843 325 3844 329
rect 3838 324 3844 325
rect 4750 328 4756 329
rect 4750 324 4751 328
rect 4755 324 4756 328
rect 4750 323 4756 324
rect 4910 328 4916 329
rect 4910 324 4911 328
rect 4915 324 4916 328
rect 4910 323 4916 324
rect 5070 328 5076 329
rect 5070 324 5071 328
rect 5075 324 5076 328
rect 5070 323 5076 324
rect 5230 328 5236 329
rect 5230 324 5231 328
rect 5235 324 5236 328
rect 5230 323 5236 324
rect 5398 328 5404 329
rect 5398 324 5399 328
rect 5403 324 5404 328
rect 5398 323 5404 324
rect 5542 328 5548 329
rect 5542 324 5543 328
rect 5547 324 5548 328
rect 5662 325 5663 329
rect 5667 325 5668 329
rect 5662 324 5668 325
rect 5542 323 5548 324
rect 210 321 216 322
rect 110 320 116 321
rect 110 316 111 320
rect 115 316 116 320
rect 210 317 211 321
rect 215 317 216 321
rect 210 316 216 317
rect 362 321 368 322
rect 362 317 363 321
rect 367 317 368 321
rect 362 316 368 317
rect 522 321 528 322
rect 522 317 523 321
rect 527 317 528 321
rect 522 316 528 317
rect 682 321 688 322
rect 682 317 683 321
rect 687 317 688 321
rect 682 316 688 317
rect 842 321 848 322
rect 842 317 843 321
rect 847 317 848 321
rect 842 316 848 317
rect 1002 321 1008 322
rect 1002 317 1003 321
rect 1007 317 1008 321
rect 1002 316 1008 317
rect 1934 320 1940 321
rect 1934 316 1935 320
rect 1939 316 1940 320
rect 110 315 116 316
rect 1934 315 1940 316
rect 4722 313 4728 314
rect 3838 312 3844 313
rect 335 311 341 312
rect 335 307 336 311
rect 340 310 341 311
rect 378 311 384 312
rect 378 310 379 311
rect 340 308 379 310
rect 340 307 341 308
rect 335 306 341 307
rect 378 307 379 308
rect 383 307 384 311
rect 378 306 384 307
rect 487 311 493 312
rect 487 307 488 311
rect 492 310 493 311
rect 538 311 544 312
rect 538 310 539 311
rect 492 308 539 310
rect 492 307 493 308
rect 487 306 493 307
rect 538 307 539 308
rect 543 307 544 311
rect 538 306 544 307
rect 558 311 564 312
rect 558 307 559 311
rect 563 310 564 311
rect 647 311 653 312
rect 647 310 648 311
rect 563 308 648 310
rect 563 307 564 308
rect 558 306 564 307
rect 647 307 648 308
rect 652 307 653 311
rect 647 306 653 307
rect 807 311 816 312
rect 807 307 808 311
rect 815 307 816 311
rect 807 306 816 307
rect 831 311 837 312
rect 831 307 832 311
rect 836 310 837 311
rect 967 311 973 312
rect 967 310 968 311
rect 836 308 968 310
rect 836 307 837 308
rect 831 306 837 307
rect 967 307 968 308
rect 972 307 973 311
rect 967 306 973 307
rect 991 311 997 312
rect 991 307 992 311
rect 996 310 997 311
rect 1127 311 1133 312
rect 1127 310 1128 311
rect 996 308 1128 310
rect 996 307 997 308
rect 991 306 997 307
rect 1127 307 1128 308
rect 1132 307 1133 311
rect 3838 308 3839 312
rect 3843 308 3844 312
rect 4722 309 4723 313
rect 4727 309 4728 313
rect 4722 308 4728 309
rect 4882 313 4888 314
rect 4882 309 4883 313
rect 4887 309 4888 313
rect 4882 308 4888 309
rect 5042 313 5048 314
rect 5042 309 5043 313
rect 5047 309 5048 313
rect 5042 308 5048 309
rect 5202 313 5208 314
rect 5202 309 5203 313
rect 5207 309 5208 313
rect 5202 308 5208 309
rect 5370 313 5376 314
rect 5370 309 5371 313
rect 5375 309 5376 313
rect 5370 308 5376 309
rect 5514 313 5520 314
rect 5514 309 5515 313
rect 5519 309 5520 313
rect 5514 308 5520 309
rect 5662 312 5668 313
rect 5662 308 5663 312
rect 5667 308 5668 312
rect 3838 307 3844 308
rect 5662 307 5668 308
rect 1127 306 1133 307
rect 4415 303 4421 304
rect 1974 301 1980 302
rect 3798 301 3804 302
rect 1974 297 1975 301
rect 1979 297 1980 301
rect 1974 296 1980 297
rect 2046 300 2052 301
rect 2046 296 2047 300
rect 2051 296 2052 300
rect 2046 295 2052 296
rect 2182 300 2188 301
rect 2182 296 2183 300
rect 2187 296 2188 300
rect 2182 295 2188 296
rect 2318 300 2324 301
rect 2318 296 2319 300
rect 2323 296 2324 300
rect 2318 295 2324 296
rect 2454 300 2460 301
rect 2454 296 2455 300
rect 2459 296 2460 300
rect 2454 295 2460 296
rect 2590 300 2596 301
rect 2590 296 2591 300
rect 2595 296 2596 300
rect 2590 295 2596 296
rect 2726 300 2732 301
rect 2726 296 2727 300
rect 2731 296 2732 300
rect 2726 295 2732 296
rect 2862 300 2868 301
rect 2862 296 2863 300
rect 2867 296 2868 300
rect 2862 295 2868 296
rect 2998 300 3004 301
rect 2998 296 2999 300
rect 3003 296 3004 300
rect 2998 295 3004 296
rect 3134 300 3140 301
rect 3134 296 3135 300
rect 3139 296 3140 300
rect 3134 295 3140 296
rect 3270 300 3276 301
rect 3270 296 3271 300
rect 3275 296 3276 300
rect 3270 295 3276 296
rect 3406 300 3412 301
rect 3406 296 3407 300
rect 3411 296 3412 300
rect 3406 295 3412 296
rect 3542 300 3548 301
rect 3542 296 3543 300
rect 3547 296 3548 300
rect 3542 295 3548 296
rect 3678 300 3684 301
rect 3678 296 3679 300
rect 3683 296 3684 300
rect 3798 297 3799 301
rect 3803 297 3804 301
rect 4415 299 4416 303
rect 4420 302 4421 303
rect 4847 303 4853 304
rect 4847 302 4848 303
rect 4420 300 4848 302
rect 4420 299 4421 300
rect 4415 298 4421 299
rect 4847 299 4848 300
rect 4852 299 4853 303
rect 4847 298 4853 299
rect 4858 303 4864 304
rect 4858 299 4859 303
rect 4863 302 4864 303
rect 5007 303 5013 304
rect 5007 302 5008 303
rect 4863 300 5008 302
rect 4863 299 4864 300
rect 4858 298 4864 299
rect 5007 299 5008 300
rect 5012 299 5013 303
rect 5007 298 5013 299
rect 5167 303 5173 304
rect 5167 299 5168 303
rect 5172 302 5173 303
rect 5218 303 5224 304
rect 5218 302 5219 303
rect 5172 300 5219 302
rect 5172 299 5173 300
rect 5167 298 5173 299
rect 5218 299 5219 300
rect 5223 299 5224 303
rect 5218 298 5224 299
rect 5327 303 5333 304
rect 5327 299 5328 303
rect 5332 302 5333 303
rect 5367 303 5373 304
rect 5367 302 5368 303
rect 5332 300 5368 302
rect 5332 299 5333 300
rect 5327 298 5333 299
rect 5367 299 5368 300
rect 5372 299 5373 303
rect 5495 303 5501 304
rect 5495 302 5496 303
rect 5367 298 5373 299
rect 5376 300 5496 302
rect 3798 296 3804 297
rect 3678 295 3684 296
rect 5130 295 5136 296
rect 5130 291 5131 295
rect 5135 294 5136 295
rect 5376 294 5378 300
rect 5495 299 5496 300
rect 5500 299 5501 303
rect 5495 298 5501 299
rect 5618 303 5624 304
rect 5618 299 5619 303
rect 5623 302 5624 303
rect 5639 303 5645 304
rect 5639 302 5640 303
rect 5623 300 5640 302
rect 5623 299 5624 300
rect 5618 298 5624 299
rect 5639 299 5640 300
rect 5644 299 5645 303
rect 5639 298 5645 299
rect 5135 292 5378 294
rect 5135 291 5136 292
rect 5130 290 5136 291
rect 2018 285 2024 286
rect 1974 284 1980 285
rect 1974 280 1975 284
rect 1979 280 1980 284
rect 2018 281 2019 285
rect 2023 281 2024 285
rect 2018 280 2024 281
rect 2154 285 2160 286
rect 2154 281 2155 285
rect 2159 281 2160 285
rect 2154 280 2160 281
rect 2290 285 2296 286
rect 2290 281 2291 285
rect 2295 281 2296 285
rect 2290 280 2296 281
rect 2426 285 2432 286
rect 2426 281 2427 285
rect 2431 281 2432 285
rect 2426 280 2432 281
rect 2562 285 2568 286
rect 2562 281 2563 285
rect 2567 281 2568 285
rect 2562 280 2568 281
rect 2698 285 2704 286
rect 2698 281 2699 285
rect 2703 281 2704 285
rect 2698 280 2704 281
rect 2834 285 2840 286
rect 2834 281 2835 285
rect 2839 281 2840 285
rect 2834 280 2840 281
rect 2970 285 2976 286
rect 2970 281 2971 285
rect 2975 281 2976 285
rect 2970 280 2976 281
rect 3106 285 3112 286
rect 3106 281 3107 285
rect 3111 281 3112 285
rect 3106 280 3112 281
rect 3242 285 3248 286
rect 3242 281 3243 285
rect 3247 281 3248 285
rect 3242 280 3248 281
rect 3378 285 3384 286
rect 3378 281 3379 285
rect 3383 281 3384 285
rect 3378 280 3384 281
rect 3514 285 3520 286
rect 3514 281 3515 285
rect 3519 281 3520 285
rect 3514 280 3520 281
rect 3650 285 3656 286
rect 3650 281 3651 285
rect 3655 281 3656 285
rect 3650 280 3656 281
rect 3798 284 3804 285
rect 3798 280 3799 284
rect 3803 280 3804 284
rect 270 279 276 280
rect 270 275 271 279
rect 275 275 276 279
rect 270 274 276 275
rect 378 279 384 280
rect 378 275 379 279
rect 383 275 384 279
rect 378 274 384 275
rect 538 279 544 280
rect 538 275 539 279
rect 543 275 544 279
rect 831 279 837 280
rect 831 278 832 279
rect 773 276 832 278
rect 538 274 544 275
rect 831 275 832 276
rect 836 275 837 279
rect 991 279 997 280
rect 991 278 992 279
rect 933 276 992 278
rect 831 274 837 275
rect 991 275 992 276
rect 996 275 997 279
rect 1518 279 1524 280
rect 1974 279 1980 280
rect 3798 279 3804 280
rect 1518 278 1519 279
rect 1093 276 1519 278
rect 991 274 997 275
rect 1518 275 1519 276
rect 1523 275 1524 279
rect 1518 274 1524 275
rect 2143 275 2149 276
rect 2143 271 2144 275
rect 2148 274 2149 275
rect 2258 275 2264 276
rect 2258 274 2259 275
rect 2148 272 2259 274
rect 2148 271 2149 272
rect 2143 270 2149 271
rect 2258 271 2259 272
rect 2263 271 2264 275
rect 2258 270 2264 271
rect 2279 275 2285 276
rect 2279 271 2280 275
rect 2284 274 2285 275
rect 2306 275 2312 276
rect 2306 274 2307 275
rect 2284 272 2307 274
rect 2284 271 2285 272
rect 2279 270 2285 271
rect 2306 271 2307 272
rect 2311 271 2312 275
rect 2306 270 2312 271
rect 2415 275 2421 276
rect 2415 271 2416 275
rect 2420 274 2421 275
rect 2442 275 2448 276
rect 2442 274 2443 275
rect 2420 272 2443 274
rect 2420 271 2421 272
rect 2415 270 2421 271
rect 2442 271 2443 272
rect 2447 271 2448 275
rect 2442 270 2448 271
rect 2530 275 2536 276
rect 2530 271 2531 275
rect 2535 274 2536 275
rect 2551 275 2557 276
rect 2551 274 2552 275
rect 2535 272 2552 274
rect 2535 271 2536 272
rect 2530 270 2536 271
rect 2551 271 2552 272
rect 2556 271 2557 275
rect 2687 275 2693 276
rect 2687 274 2688 275
rect 2551 270 2557 271
rect 2560 272 2688 274
rect 2560 258 2562 272
rect 2687 271 2688 272
rect 2692 271 2693 275
rect 2687 270 2693 271
rect 2695 275 2701 276
rect 2695 271 2696 275
rect 2700 274 2701 275
rect 2823 275 2829 276
rect 2823 274 2824 275
rect 2700 272 2824 274
rect 2700 271 2701 272
rect 2695 270 2701 271
rect 2823 271 2824 272
rect 2828 271 2829 275
rect 2823 270 2829 271
rect 2959 275 2965 276
rect 2959 271 2960 275
rect 2964 274 2965 275
rect 2986 275 2992 276
rect 2986 274 2987 275
rect 2964 272 2987 274
rect 2964 271 2965 272
rect 2959 270 2965 271
rect 2986 271 2987 272
rect 2991 271 2992 275
rect 2986 270 2992 271
rect 3095 275 3101 276
rect 3095 271 3096 275
rect 3100 274 3101 275
rect 3122 275 3128 276
rect 3122 274 3123 275
rect 3100 272 3123 274
rect 3100 271 3101 272
rect 3095 270 3101 271
rect 3122 271 3123 272
rect 3127 271 3128 275
rect 3122 270 3128 271
rect 3231 275 3240 276
rect 3231 271 3232 275
rect 3239 271 3240 275
rect 3367 275 3373 276
rect 3367 274 3368 275
rect 3231 270 3240 271
rect 3252 272 3368 274
rect 2922 267 2928 268
rect 2922 263 2923 267
rect 2927 266 2928 267
rect 3252 266 3254 272
rect 3367 271 3368 272
rect 3372 271 3373 275
rect 3367 270 3373 271
rect 3503 275 3509 276
rect 3503 271 3504 275
rect 3508 274 3509 275
rect 3530 275 3536 276
rect 3530 274 3531 275
rect 3508 272 3531 274
rect 3508 271 3509 272
rect 3503 270 3509 271
rect 3530 271 3531 272
rect 3535 271 3536 275
rect 3530 270 3536 271
rect 3639 275 3645 276
rect 3639 271 3640 275
rect 3644 274 3645 275
rect 3666 275 3672 276
rect 3666 274 3667 275
rect 3644 272 3667 274
rect 3644 271 3645 272
rect 3639 270 3645 271
rect 3666 271 3667 272
rect 3671 271 3672 275
rect 3775 275 3781 276
rect 3775 274 3776 275
rect 3666 270 3672 271
rect 3676 272 3776 274
rect 2927 264 3254 266
rect 3330 267 3336 268
rect 2927 263 2928 264
rect 2922 262 2928 263
rect 3330 263 3331 267
rect 3335 266 3336 267
rect 3676 266 3678 272
rect 3775 271 3776 272
rect 3780 271 3781 275
rect 3775 270 3781 271
rect 4858 271 4864 272
rect 4858 270 4859 271
rect 4813 268 4859 270
rect 4858 267 4859 268
rect 4863 267 4864 271
rect 5034 271 5040 272
rect 5034 270 5035 271
rect 4973 268 5035 270
rect 4858 266 4864 267
rect 5034 267 5035 268
rect 5039 267 5040 271
rect 5034 266 5040 267
rect 5130 271 5136 272
rect 5130 267 5131 271
rect 5135 267 5136 271
rect 5130 266 5136 267
rect 5218 271 5224 272
rect 5218 267 5219 271
rect 5223 267 5224 271
rect 5218 266 5224 267
rect 5386 271 5392 272
rect 5386 267 5387 271
rect 5391 267 5392 271
rect 5386 266 5392 267
rect 5602 271 5608 272
rect 5602 267 5603 271
rect 5607 267 5608 271
rect 5602 266 5608 267
rect 3335 264 3678 266
rect 3335 263 3336 264
rect 3330 262 3336 263
rect 2248 256 2562 258
rect 2106 243 2112 244
rect 2106 239 2107 243
rect 2111 239 2112 243
rect 2248 242 2250 256
rect 2245 240 2250 242
rect 2306 243 2312 244
rect 2106 238 2112 239
rect 2306 239 2307 243
rect 2311 239 2312 243
rect 2306 238 2312 239
rect 2442 243 2448 244
rect 2442 239 2443 243
rect 2447 239 2448 243
rect 2695 243 2701 244
rect 2695 242 2696 243
rect 2653 240 2696 242
rect 2442 238 2448 239
rect 2695 239 2696 240
rect 2700 239 2701 243
rect 2842 243 2848 244
rect 2842 242 2843 243
rect 2789 240 2843 242
rect 2695 238 2701 239
rect 2842 239 2843 240
rect 2847 239 2848 243
rect 2842 238 2848 239
rect 2922 243 2928 244
rect 2922 239 2923 243
rect 2927 239 2928 243
rect 2922 238 2928 239
rect 2986 243 2992 244
rect 2986 239 2987 243
rect 2991 239 2992 243
rect 2986 238 2992 239
rect 3122 243 3128 244
rect 3122 239 3123 243
rect 3127 239 3128 243
rect 3122 238 3128 239
rect 3330 243 3336 244
rect 3330 239 3331 243
rect 3335 239 3336 243
rect 3330 238 3336 239
rect 3422 243 3428 244
rect 3422 239 3423 243
rect 3427 239 3428 243
rect 3422 238 3428 239
rect 3530 243 3536 244
rect 3530 239 3531 243
rect 3535 239 3536 243
rect 3530 238 3536 239
rect 3666 243 3672 244
rect 3666 239 3667 243
rect 3671 239 3672 243
rect 3666 238 3672 239
rect 1202 211 1208 212
rect 1202 210 1203 211
rect 804 208 1203 210
rect 279 199 285 200
rect 279 198 280 199
rect 237 196 280 198
rect 279 195 280 196
rect 284 195 285 199
rect 415 199 421 200
rect 415 198 416 199
rect 373 196 416 198
rect 279 194 285 195
rect 415 195 416 196
rect 420 195 421 199
rect 551 199 557 200
rect 551 198 552 199
rect 509 196 552 198
rect 415 194 421 195
rect 551 195 552 196
rect 556 195 557 199
rect 687 199 693 200
rect 687 198 688 199
rect 645 196 688 198
rect 551 194 557 195
rect 687 195 688 196
rect 692 195 693 199
rect 804 198 806 208
rect 1202 207 1203 208
rect 1207 207 1208 211
rect 1202 206 1208 207
rect 781 196 806 198
rect 810 199 816 200
rect 687 194 693 195
rect 810 195 811 199
rect 815 198 816 199
rect 959 199 965 200
rect 815 196 845 198
rect 815 195 816 196
rect 810 194 816 195
rect 959 195 960 199
rect 964 198 965 199
rect 1095 199 1101 200
rect 964 196 981 198
rect 964 195 965 196
rect 959 194 965 195
rect 1095 195 1096 199
rect 1100 198 1101 199
rect 1100 196 1117 198
rect 1100 195 1101 196
rect 1095 194 1101 195
rect 3234 195 3240 196
rect 3234 191 3235 195
rect 3239 194 3240 195
rect 3239 192 3322 194
rect 3239 191 3240 192
rect 3234 190 3240 191
rect 2127 179 2133 180
rect 2127 178 2128 179
rect 2085 176 2128 178
rect 2127 175 2128 176
rect 2132 175 2133 179
rect 2263 179 2269 180
rect 2263 178 2264 179
rect 2221 176 2264 178
rect 2127 174 2133 175
rect 2263 175 2264 176
rect 2268 175 2269 179
rect 2399 179 2405 180
rect 2399 178 2400 179
rect 2357 176 2400 178
rect 2263 174 2269 175
rect 2399 175 2400 176
rect 2404 175 2405 179
rect 2530 179 2536 180
rect 2399 174 2405 175
rect 2490 175 2496 176
rect 2490 171 2491 175
rect 2495 171 2496 175
rect 2530 175 2531 179
rect 2535 178 2536 179
rect 2671 179 2677 180
rect 2535 176 2557 178
rect 2535 175 2536 176
rect 2530 174 2536 175
rect 2671 175 2672 179
rect 2676 178 2677 179
rect 2807 179 2813 180
rect 2676 176 2693 178
rect 2676 175 2677 176
rect 2671 174 2677 175
rect 2807 175 2808 179
rect 2812 178 2813 179
rect 3079 179 3085 180
rect 3079 178 3080 179
rect 2812 176 2829 178
rect 3037 176 3080 178
rect 2812 175 2813 176
rect 2807 174 2813 175
rect 3079 175 3080 176
rect 3084 175 3085 179
rect 3215 179 3221 180
rect 3215 178 3216 179
rect 3173 176 3216 178
rect 3079 174 3085 175
rect 3215 175 3216 176
rect 3220 175 3221 179
rect 3320 178 3322 192
rect 4415 183 4421 184
rect 4415 182 4416 183
rect 4381 180 4416 182
rect 3487 179 3493 180
rect 3320 176 3373 178
rect 3215 174 3221 175
rect 3306 175 3312 176
rect 2490 170 2496 171
rect 3306 171 3307 175
rect 3311 171 3312 175
rect 3487 175 3488 179
rect 3492 178 3493 179
rect 3623 179 3629 180
rect 3492 176 3509 178
rect 3492 175 3493 176
rect 3487 174 3493 175
rect 3623 175 3624 179
rect 3628 178 3629 179
rect 4415 179 4416 180
rect 4420 179 4421 183
rect 4415 178 4421 179
rect 4423 183 4429 184
rect 4423 179 4424 183
rect 4428 182 4429 183
rect 4559 183 4565 184
rect 4428 180 4445 182
rect 4428 179 4429 180
rect 4423 178 4429 179
rect 4559 179 4560 183
rect 4564 182 4565 183
rect 4695 183 4701 184
rect 4564 180 4581 182
rect 4564 179 4565 180
rect 4559 178 4565 179
rect 4695 179 4696 183
rect 4700 182 4701 183
rect 4826 183 4832 184
rect 4700 180 4717 182
rect 4700 179 4701 180
rect 4695 178 4701 179
rect 4826 179 4827 183
rect 4831 182 4832 183
rect 4967 183 4973 184
rect 4831 180 4853 182
rect 4831 179 4832 180
rect 4826 178 4832 179
rect 4967 179 4968 183
rect 4972 182 4973 183
rect 5103 183 5109 184
rect 4972 180 4989 182
rect 4972 179 4973 180
rect 4967 178 4973 179
rect 5103 179 5104 183
rect 5108 182 5109 183
rect 5239 183 5245 184
rect 5108 180 5125 182
rect 5108 179 5109 180
rect 5103 178 5109 179
rect 5239 179 5240 183
rect 5244 182 5245 183
rect 5618 183 5624 184
rect 5618 182 5619 183
rect 5244 180 5261 182
rect 5605 180 5619 182
rect 5244 179 5245 180
rect 5239 178 5245 179
rect 5466 179 5472 180
rect 3628 176 3645 178
rect 3628 175 3629 176
rect 3623 174 3629 175
rect 5466 175 5467 179
rect 5471 175 5472 179
rect 5618 179 5619 180
rect 5623 179 5624 183
rect 5618 178 5624 179
rect 5466 174 5472 175
rect 3306 170 3312 171
rect 270 163 277 164
rect 270 159 271 163
rect 276 159 277 163
rect 270 158 277 159
rect 279 163 285 164
rect 279 159 280 163
rect 284 162 285 163
rect 407 163 413 164
rect 407 162 408 163
rect 284 160 408 162
rect 284 159 285 160
rect 279 158 285 159
rect 407 159 408 160
rect 412 159 413 163
rect 407 158 413 159
rect 415 163 421 164
rect 415 159 416 163
rect 420 162 421 163
rect 543 163 549 164
rect 543 162 544 163
rect 420 160 544 162
rect 420 159 421 160
rect 415 158 421 159
rect 543 159 544 160
rect 548 159 549 163
rect 543 158 549 159
rect 551 163 557 164
rect 551 159 552 163
rect 556 162 557 163
rect 679 163 685 164
rect 679 162 680 163
rect 556 160 680 162
rect 556 159 557 160
rect 551 158 557 159
rect 679 159 680 160
rect 684 159 685 163
rect 679 158 685 159
rect 687 163 693 164
rect 687 159 688 163
rect 692 162 693 163
rect 815 163 821 164
rect 815 162 816 163
rect 692 160 816 162
rect 692 159 693 160
rect 687 158 693 159
rect 815 159 816 160
rect 820 159 821 163
rect 815 158 821 159
rect 951 163 957 164
rect 951 159 952 163
rect 956 162 957 163
rect 959 163 965 164
rect 959 162 960 163
rect 956 160 960 162
rect 956 159 957 160
rect 951 158 957 159
rect 959 159 960 160
rect 964 159 965 163
rect 959 158 965 159
rect 1087 163 1093 164
rect 1087 159 1088 163
rect 1092 162 1093 163
rect 1095 163 1101 164
rect 1095 162 1096 163
rect 1092 160 1096 162
rect 1092 159 1093 160
rect 1087 158 1093 159
rect 1095 159 1096 160
rect 1100 159 1101 163
rect 1095 158 1101 159
rect 1202 163 1208 164
rect 1202 159 1203 163
rect 1207 162 1208 163
rect 1223 163 1229 164
rect 1223 162 1224 163
rect 1207 160 1224 162
rect 1207 159 1208 160
rect 1202 158 1208 159
rect 1223 159 1224 160
rect 1228 159 1229 163
rect 1223 158 1229 159
rect 110 156 116 157
rect 1934 156 1940 157
rect 110 152 111 156
rect 115 152 116 156
rect 110 151 116 152
rect 146 155 152 156
rect 146 151 147 155
rect 151 151 152 155
rect 146 150 152 151
rect 282 155 288 156
rect 282 151 283 155
rect 287 151 288 155
rect 282 150 288 151
rect 418 155 424 156
rect 418 151 419 155
rect 423 151 424 155
rect 418 150 424 151
rect 554 155 560 156
rect 554 151 555 155
rect 559 151 560 155
rect 554 150 560 151
rect 690 155 696 156
rect 690 151 691 155
rect 695 151 696 155
rect 690 150 696 151
rect 826 155 832 156
rect 826 151 827 155
rect 831 151 832 155
rect 826 150 832 151
rect 962 155 968 156
rect 962 151 963 155
rect 967 151 968 155
rect 962 150 968 151
rect 1098 155 1104 156
rect 1098 151 1099 155
rect 1103 151 1104 155
rect 1934 152 1935 156
rect 1939 152 1940 156
rect 1934 151 1940 152
rect 2490 151 2496 152
rect 1098 150 1104 151
rect 2490 147 2491 151
rect 2495 150 2496 151
rect 2842 151 2848 152
rect 2495 148 2818 150
rect 2495 147 2496 148
rect 2490 146 2496 147
rect 2106 143 2112 144
rect 174 140 180 141
rect 110 139 116 140
rect 110 135 111 139
rect 115 135 116 139
rect 174 136 175 140
rect 179 136 180 140
rect 174 135 180 136
rect 310 140 316 141
rect 310 136 311 140
rect 315 136 316 140
rect 310 135 316 136
rect 446 140 452 141
rect 446 136 447 140
rect 451 136 452 140
rect 446 135 452 136
rect 582 140 588 141
rect 582 136 583 140
rect 587 136 588 140
rect 582 135 588 136
rect 718 140 724 141
rect 718 136 719 140
rect 723 136 724 140
rect 718 135 724 136
rect 854 140 860 141
rect 854 136 855 140
rect 859 136 860 140
rect 854 135 860 136
rect 990 140 996 141
rect 990 136 991 140
rect 995 136 996 140
rect 990 135 996 136
rect 1126 140 1132 141
rect 1126 136 1127 140
rect 1131 136 1132 140
rect 1126 135 1132 136
rect 1934 139 1940 140
rect 1934 135 1935 139
rect 1939 135 1940 139
rect 2106 139 2107 143
rect 2111 142 2112 143
rect 2119 143 2125 144
rect 2119 142 2120 143
rect 2111 140 2120 142
rect 2111 139 2112 140
rect 2106 138 2112 139
rect 2119 139 2120 140
rect 2124 139 2125 143
rect 2119 138 2125 139
rect 2127 143 2133 144
rect 2127 139 2128 143
rect 2132 142 2133 143
rect 2255 143 2261 144
rect 2255 142 2256 143
rect 2132 140 2256 142
rect 2132 139 2133 140
rect 2127 138 2133 139
rect 2255 139 2256 140
rect 2260 139 2261 143
rect 2255 138 2261 139
rect 2263 143 2269 144
rect 2263 139 2264 143
rect 2268 142 2269 143
rect 2391 143 2397 144
rect 2391 142 2392 143
rect 2268 140 2392 142
rect 2268 139 2269 140
rect 2263 138 2269 139
rect 2391 139 2392 140
rect 2396 139 2397 143
rect 2391 138 2397 139
rect 2399 143 2405 144
rect 2399 139 2400 143
rect 2404 142 2405 143
rect 2527 143 2533 144
rect 2527 142 2528 143
rect 2404 140 2528 142
rect 2404 139 2405 140
rect 2399 138 2405 139
rect 2527 139 2528 140
rect 2532 139 2533 143
rect 2527 138 2533 139
rect 2663 143 2669 144
rect 2663 139 2664 143
rect 2668 142 2669 143
rect 2671 143 2677 144
rect 2671 142 2672 143
rect 2668 140 2672 142
rect 2668 139 2669 140
rect 2663 138 2669 139
rect 2671 139 2672 140
rect 2676 139 2677 143
rect 2671 138 2677 139
rect 2799 143 2805 144
rect 2799 139 2800 143
rect 2804 142 2805 143
rect 2807 143 2813 144
rect 2807 142 2808 143
rect 2804 140 2808 142
rect 2804 139 2805 140
rect 2799 138 2805 139
rect 2807 139 2808 140
rect 2812 139 2813 143
rect 2816 142 2818 148
rect 2842 147 2843 151
rect 2847 150 2848 151
rect 3306 151 3312 152
rect 2847 148 2946 150
rect 2847 147 2848 148
rect 2842 146 2848 147
rect 2935 143 2941 144
rect 2935 142 2936 143
rect 2816 140 2936 142
rect 2807 138 2813 139
rect 2935 139 2936 140
rect 2940 139 2941 143
rect 2944 142 2946 148
rect 3306 147 3307 151
rect 3311 150 3312 151
rect 3311 148 3634 150
rect 3311 147 3312 148
rect 3306 146 3312 147
rect 3071 143 3077 144
rect 3071 142 3072 143
rect 2944 140 3072 142
rect 2935 138 2941 139
rect 3071 139 3072 140
rect 3076 139 3077 143
rect 3071 138 3077 139
rect 3079 143 3085 144
rect 3079 139 3080 143
rect 3084 142 3085 143
rect 3207 143 3213 144
rect 3207 142 3208 143
rect 3084 140 3208 142
rect 3084 139 3085 140
rect 3079 138 3085 139
rect 3207 139 3208 140
rect 3212 139 3213 143
rect 3207 138 3213 139
rect 3215 143 3221 144
rect 3215 139 3216 143
rect 3220 142 3221 143
rect 3343 143 3349 144
rect 3343 142 3344 143
rect 3220 140 3344 142
rect 3220 139 3221 140
rect 3215 138 3221 139
rect 3343 139 3344 140
rect 3348 139 3349 143
rect 3343 138 3349 139
rect 3479 143 3485 144
rect 3479 139 3480 143
rect 3484 142 3485 143
rect 3487 143 3493 144
rect 3487 142 3488 143
rect 3484 140 3488 142
rect 3484 139 3485 140
rect 3479 138 3485 139
rect 3487 139 3488 140
rect 3492 139 3493 143
rect 3487 138 3493 139
rect 3615 143 3621 144
rect 3615 139 3616 143
rect 3620 142 3621 143
rect 3623 143 3629 144
rect 3623 142 3624 143
rect 3620 140 3624 142
rect 3620 139 3621 140
rect 3615 138 3621 139
rect 3623 139 3624 140
rect 3628 139 3629 143
rect 3632 142 3634 148
rect 4415 147 4421 148
rect 3751 143 3757 144
rect 3751 142 3752 143
rect 3632 140 3752 142
rect 3623 138 3629 139
rect 3751 139 3752 140
rect 3756 139 3757 143
rect 4415 143 4416 147
rect 4420 146 4421 147
rect 4423 147 4429 148
rect 4423 146 4424 147
rect 4420 144 4424 146
rect 4420 143 4421 144
rect 4415 142 4421 143
rect 4423 143 4424 144
rect 4428 143 4429 147
rect 4423 142 4429 143
rect 4551 147 4557 148
rect 4551 143 4552 147
rect 4556 146 4557 147
rect 4559 147 4565 148
rect 4559 146 4560 147
rect 4556 144 4560 146
rect 4556 143 4557 144
rect 4551 142 4557 143
rect 4559 143 4560 144
rect 4564 143 4565 147
rect 4559 142 4565 143
rect 4687 147 4693 148
rect 4687 143 4688 147
rect 4692 146 4693 147
rect 4695 147 4701 148
rect 4695 146 4696 147
rect 4692 144 4696 146
rect 4692 143 4693 144
rect 4687 142 4693 143
rect 4695 143 4696 144
rect 4700 143 4701 147
rect 4695 142 4701 143
rect 4823 147 4832 148
rect 4823 143 4824 147
rect 4831 143 4832 147
rect 4823 142 4832 143
rect 4959 147 4965 148
rect 4959 143 4960 147
rect 4964 146 4965 147
rect 4967 147 4973 148
rect 4967 146 4968 147
rect 4964 144 4968 146
rect 4964 143 4965 144
rect 4959 142 4965 143
rect 4967 143 4968 144
rect 4972 143 4973 147
rect 4967 142 4973 143
rect 5095 147 5101 148
rect 5095 143 5096 147
rect 5100 146 5101 147
rect 5103 147 5109 148
rect 5103 146 5104 147
rect 5100 144 5104 146
rect 5100 143 5101 144
rect 5095 142 5101 143
rect 5103 143 5104 144
rect 5108 143 5109 147
rect 5103 142 5109 143
rect 5231 147 5237 148
rect 5231 143 5232 147
rect 5236 146 5237 147
rect 5239 147 5245 148
rect 5239 146 5240 147
rect 5236 144 5240 146
rect 5236 143 5237 144
rect 5231 142 5237 143
rect 5239 143 5240 144
rect 5244 143 5245 147
rect 5239 142 5245 143
rect 5367 147 5373 148
rect 5367 143 5368 147
rect 5372 146 5373 147
rect 5386 147 5392 148
rect 5386 146 5387 147
rect 5372 144 5387 146
rect 5372 143 5373 144
rect 5367 142 5373 143
rect 5386 143 5387 144
rect 5391 143 5392 147
rect 5386 142 5392 143
rect 5466 147 5472 148
rect 5466 143 5467 147
rect 5471 146 5472 147
rect 5639 147 5645 148
rect 5639 146 5640 147
rect 5471 144 5640 146
rect 5471 143 5472 144
rect 5466 142 5472 143
rect 5639 143 5640 144
rect 5644 143 5645 147
rect 5639 142 5645 143
rect 3751 138 3757 139
rect 3838 140 3844 141
rect 5662 140 5668 141
rect 110 134 116 135
rect 1934 134 1940 135
rect 1974 136 1980 137
rect 3798 136 3804 137
rect 1974 132 1975 136
rect 1979 132 1980 136
rect 1974 131 1980 132
rect 1994 135 2000 136
rect 1994 131 1995 135
rect 1999 131 2000 135
rect 1994 130 2000 131
rect 2130 135 2136 136
rect 2130 131 2131 135
rect 2135 131 2136 135
rect 2130 130 2136 131
rect 2266 135 2272 136
rect 2266 131 2267 135
rect 2271 131 2272 135
rect 2266 130 2272 131
rect 2402 135 2408 136
rect 2402 131 2403 135
rect 2407 131 2408 135
rect 2402 130 2408 131
rect 2538 135 2544 136
rect 2538 131 2539 135
rect 2543 131 2544 135
rect 2538 130 2544 131
rect 2674 135 2680 136
rect 2674 131 2675 135
rect 2679 131 2680 135
rect 2674 130 2680 131
rect 2810 135 2816 136
rect 2810 131 2811 135
rect 2815 131 2816 135
rect 2810 130 2816 131
rect 2946 135 2952 136
rect 2946 131 2947 135
rect 2951 131 2952 135
rect 2946 130 2952 131
rect 3082 135 3088 136
rect 3082 131 3083 135
rect 3087 131 3088 135
rect 3082 130 3088 131
rect 3218 135 3224 136
rect 3218 131 3219 135
rect 3223 131 3224 135
rect 3218 130 3224 131
rect 3354 135 3360 136
rect 3354 131 3355 135
rect 3359 131 3360 135
rect 3354 130 3360 131
rect 3490 135 3496 136
rect 3490 131 3491 135
rect 3495 131 3496 135
rect 3490 130 3496 131
rect 3626 135 3632 136
rect 3626 131 3627 135
rect 3631 131 3632 135
rect 3798 132 3799 136
rect 3803 132 3804 136
rect 3838 136 3839 140
rect 3843 136 3844 140
rect 3838 135 3844 136
rect 4290 139 4296 140
rect 4290 135 4291 139
rect 4295 135 4296 139
rect 4290 134 4296 135
rect 4426 139 4432 140
rect 4426 135 4427 139
rect 4431 135 4432 139
rect 4426 134 4432 135
rect 4562 139 4568 140
rect 4562 135 4563 139
rect 4567 135 4568 139
rect 4562 134 4568 135
rect 4698 139 4704 140
rect 4698 135 4699 139
rect 4703 135 4704 139
rect 4698 134 4704 135
rect 4834 139 4840 140
rect 4834 135 4835 139
rect 4839 135 4840 139
rect 4834 134 4840 135
rect 4970 139 4976 140
rect 4970 135 4971 139
rect 4975 135 4976 139
rect 4970 134 4976 135
rect 5106 139 5112 140
rect 5106 135 5107 139
rect 5111 135 5112 139
rect 5106 134 5112 135
rect 5242 139 5248 140
rect 5242 135 5243 139
rect 5247 135 5248 139
rect 5242 134 5248 135
rect 5378 139 5384 140
rect 5378 135 5379 139
rect 5383 135 5384 139
rect 5378 134 5384 135
rect 5514 139 5520 140
rect 5514 135 5515 139
rect 5519 135 5520 139
rect 5662 136 5663 140
rect 5667 136 5668 140
rect 5662 135 5668 136
rect 5514 134 5520 135
rect 3798 131 3804 132
rect 3626 130 3632 131
rect 4318 124 4324 125
rect 3838 123 3844 124
rect 2022 120 2028 121
rect 1974 119 1980 120
rect 1974 115 1975 119
rect 1979 115 1980 119
rect 2022 116 2023 120
rect 2027 116 2028 120
rect 2022 115 2028 116
rect 2158 120 2164 121
rect 2158 116 2159 120
rect 2163 116 2164 120
rect 2158 115 2164 116
rect 2294 120 2300 121
rect 2294 116 2295 120
rect 2299 116 2300 120
rect 2294 115 2300 116
rect 2430 120 2436 121
rect 2430 116 2431 120
rect 2435 116 2436 120
rect 2430 115 2436 116
rect 2566 120 2572 121
rect 2566 116 2567 120
rect 2571 116 2572 120
rect 2566 115 2572 116
rect 2702 120 2708 121
rect 2702 116 2703 120
rect 2707 116 2708 120
rect 2702 115 2708 116
rect 2838 120 2844 121
rect 2838 116 2839 120
rect 2843 116 2844 120
rect 2838 115 2844 116
rect 2974 120 2980 121
rect 2974 116 2975 120
rect 2979 116 2980 120
rect 2974 115 2980 116
rect 3110 120 3116 121
rect 3110 116 3111 120
rect 3115 116 3116 120
rect 3110 115 3116 116
rect 3246 120 3252 121
rect 3246 116 3247 120
rect 3251 116 3252 120
rect 3246 115 3252 116
rect 3382 120 3388 121
rect 3382 116 3383 120
rect 3387 116 3388 120
rect 3382 115 3388 116
rect 3518 120 3524 121
rect 3518 116 3519 120
rect 3523 116 3524 120
rect 3518 115 3524 116
rect 3654 120 3660 121
rect 3654 116 3655 120
rect 3659 116 3660 120
rect 3654 115 3660 116
rect 3798 119 3804 120
rect 3798 115 3799 119
rect 3803 115 3804 119
rect 3838 119 3839 123
rect 3843 119 3844 123
rect 4318 120 4319 124
rect 4323 120 4324 124
rect 4318 119 4324 120
rect 4454 124 4460 125
rect 4454 120 4455 124
rect 4459 120 4460 124
rect 4454 119 4460 120
rect 4590 124 4596 125
rect 4590 120 4591 124
rect 4595 120 4596 124
rect 4590 119 4596 120
rect 4726 124 4732 125
rect 4726 120 4727 124
rect 4731 120 4732 124
rect 4726 119 4732 120
rect 4862 124 4868 125
rect 4862 120 4863 124
rect 4867 120 4868 124
rect 4862 119 4868 120
rect 4998 124 5004 125
rect 4998 120 4999 124
rect 5003 120 5004 124
rect 4998 119 5004 120
rect 5134 124 5140 125
rect 5134 120 5135 124
rect 5139 120 5140 124
rect 5134 119 5140 120
rect 5270 124 5276 125
rect 5270 120 5271 124
rect 5275 120 5276 124
rect 5270 119 5276 120
rect 5406 124 5412 125
rect 5406 120 5407 124
rect 5411 120 5412 124
rect 5406 119 5412 120
rect 5542 124 5548 125
rect 5542 120 5543 124
rect 5547 120 5548 124
rect 5542 119 5548 120
rect 5662 123 5668 124
rect 5662 119 5663 123
rect 5667 119 5668 123
rect 3838 118 3844 119
rect 5662 118 5668 119
rect 1974 114 1980 115
rect 3798 114 3804 115
<< m3c >>
rect 259 5731 263 5735
rect 259 5695 260 5699
rect 260 5695 263 5699
rect 423 5695 427 5699
rect 111 5688 115 5692
rect 131 5687 135 5691
rect 267 5687 271 5691
rect 403 5687 407 5691
rect 1935 5688 1939 5692
rect 111 5671 115 5675
rect 159 5672 163 5676
rect 295 5672 299 5676
rect 431 5672 435 5676
rect 1935 5671 1939 5675
rect 2651 5659 2655 5663
rect 2875 5663 2879 5667
rect 3059 5663 3063 5667
rect 3235 5663 3239 5667
rect 3403 5663 3407 5667
rect 3571 5663 3575 5667
rect 4555 5663 4559 5667
rect 3067 5647 3071 5651
rect 1943 5627 1947 5631
rect 2875 5627 2876 5631
rect 2876 5627 2879 5631
rect 3059 5627 3060 5631
rect 3060 5627 3063 5631
rect 3235 5627 3236 5631
rect 3236 5627 3239 5631
rect 3403 5627 3404 5631
rect 3404 5627 3407 5631
rect 3571 5627 3572 5631
rect 3572 5627 3575 5631
rect 3739 5627 3743 5631
rect 4911 5631 4915 5635
rect 1975 5620 1979 5624
rect 1995 5619 1999 5623
rect 2171 5619 2175 5623
rect 2371 5619 2375 5623
rect 2563 5619 2567 5623
rect 2747 5619 2751 5623
rect 2931 5619 2935 5623
rect 3107 5619 3111 5623
rect 3275 5619 3279 5623
rect 3443 5619 3447 5623
rect 3619 5619 3623 5623
rect 3799 5620 3803 5624
rect 3839 5624 3843 5628
rect 4467 5623 4471 5627
rect 4603 5623 4607 5627
rect 4739 5623 4743 5627
rect 4875 5623 4879 5627
rect 5663 5624 5667 5628
rect 111 5613 115 5617
rect 343 5612 347 5616
rect 535 5612 539 5616
rect 735 5612 739 5616
rect 943 5612 947 5616
rect 1159 5612 1163 5616
rect 1383 5612 1387 5616
rect 1607 5612 1611 5616
rect 1815 5612 1819 5616
rect 1935 5613 1939 5617
rect 1975 5603 1979 5607
rect 2023 5604 2027 5608
rect 2199 5604 2203 5608
rect 2399 5604 2403 5608
rect 2591 5604 2595 5608
rect 2775 5604 2779 5608
rect 2959 5604 2963 5608
rect 3135 5604 3139 5608
rect 3303 5604 3307 5608
rect 3471 5604 3475 5608
rect 3647 5604 3651 5608
rect 3799 5603 3803 5607
rect 3839 5607 3843 5611
rect 4495 5608 4499 5612
rect 4631 5608 4635 5612
rect 4767 5608 4771 5612
rect 4903 5608 4907 5612
rect 5663 5607 5667 5611
rect 111 5596 115 5600
rect 315 5597 319 5601
rect 507 5597 511 5601
rect 707 5597 711 5601
rect 915 5597 919 5601
rect 1131 5597 1135 5601
rect 1355 5597 1359 5601
rect 1579 5597 1583 5601
rect 1787 5597 1791 5601
rect 1935 5596 1939 5600
rect 523 5587 527 5591
rect 723 5587 727 5591
rect 931 5587 935 5591
rect 1147 5587 1151 5591
rect 999 5579 1003 5583
rect 423 5555 427 5559
rect 523 5555 527 5559
rect 723 5555 727 5559
rect 931 5555 935 5559
rect 1147 5555 1151 5559
rect 1943 5555 1947 5559
rect 1975 5545 1979 5549
rect 2375 5544 2379 5548
rect 2607 5544 2611 5548
rect 2831 5544 2835 5548
rect 3047 5544 3051 5548
rect 3263 5544 3267 5548
rect 3479 5544 3483 5548
rect 3679 5544 3683 5548
rect 3799 5545 3803 5549
rect 3839 5549 3843 5553
rect 4431 5548 4435 5552
rect 4567 5548 4571 5552
rect 4703 5548 4707 5552
rect 4839 5548 4843 5552
rect 4975 5548 4979 5552
rect 5111 5548 5115 5552
rect 5663 5549 5667 5553
rect 1847 5527 1851 5531
rect 1975 5528 1979 5532
rect 2347 5529 2351 5533
rect 2579 5529 2583 5533
rect 2803 5529 2807 5533
rect 3019 5529 3023 5533
rect 3235 5529 3239 5533
rect 3451 5529 3455 5533
rect 3651 5529 3655 5533
rect 3799 5528 3803 5532
rect 3839 5532 3843 5536
rect 4403 5533 4407 5537
rect 4539 5533 4543 5537
rect 4675 5533 4679 5537
rect 4811 5533 4815 5537
rect 4947 5533 4951 5537
rect 5083 5533 5087 5537
rect 5663 5532 5667 5536
rect 2595 5519 2599 5523
rect 2651 5519 2655 5523
rect 3035 5519 3039 5523
rect 3067 5519 3071 5523
rect 3467 5519 3471 5523
rect 3579 5519 3580 5523
rect 3580 5519 3583 5523
rect 999 5507 1003 5511
rect 1419 5507 1423 5511
rect 1707 5507 1711 5511
rect 3323 5511 3327 5515
rect 4555 5523 4559 5527
rect 4491 5515 4495 5519
rect 4827 5523 4831 5527
rect 4963 5523 4967 5527
rect 5099 5523 5103 5527
rect 4887 5515 4891 5519
rect 2435 5487 2439 5491
rect 2595 5487 2599 5491
rect 2823 5487 2827 5491
rect 3035 5487 3039 5491
rect 3323 5487 3327 5491
rect 3467 5487 3471 5491
rect 3739 5487 3743 5491
rect 4491 5491 4495 5495
rect 4627 5491 4631 5495
rect 4911 5507 4915 5511
rect 4827 5491 4831 5495
rect 4963 5491 4967 5495
rect 5099 5491 5103 5495
rect 1271 5471 1272 5475
rect 1272 5471 1275 5475
rect 1419 5471 1420 5475
rect 1420 5471 1423 5475
rect 1559 5471 1560 5475
rect 1560 5471 1563 5475
rect 1707 5471 1708 5475
rect 1708 5471 1711 5475
rect 1847 5471 1848 5475
rect 1848 5471 1851 5475
rect 111 5464 115 5468
rect 875 5463 879 5467
rect 1011 5463 1015 5467
rect 1147 5463 1151 5467
rect 1291 5463 1295 5467
rect 1435 5463 1439 5467
rect 1579 5463 1583 5467
rect 1723 5463 1727 5467
rect 1935 5464 1939 5468
rect 111 5447 115 5451
rect 903 5448 907 5452
rect 1039 5448 1043 5452
rect 1175 5448 1179 5452
rect 1319 5448 1323 5452
rect 1463 5448 1467 5452
rect 1607 5448 1611 5452
rect 1751 5448 1755 5452
rect 1935 5447 1939 5451
rect 2419 5435 2423 5439
rect 2895 5435 2899 5439
rect 3035 5431 3039 5435
rect 3275 5431 3279 5435
rect 3315 5435 3319 5439
rect 3579 5435 3583 5439
rect 4515 5439 4519 5443
rect 4887 5443 4891 5447
rect 3275 5411 3279 5415
rect 2435 5399 2439 5403
rect 2823 5399 2824 5403
rect 2824 5399 2827 5403
rect 2895 5399 2899 5403
rect 3315 5399 3316 5403
rect 3316 5399 3319 5403
rect 3551 5399 3552 5403
rect 3552 5399 3555 5403
rect 4627 5407 4631 5411
rect 5199 5407 5200 5411
rect 5200 5407 5203 5411
rect 3839 5400 3843 5404
rect 4427 5399 4431 5403
rect 4587 5399 4591 5403
rect 4747 5399 4751 5403
rect 4907 5399 4911 5403
rect 5075 5399 5079 5403
rect 5663 5400 5667 5404
rect 111 5389 115 5393
rect 719 5388 723 5392
rect 855 5388 859 5392
rect 991 5388 995 5392
rect 1127 5388 1131 5392
rect 1263 5388 1267 5392
rect 1399 5388 1403 5392
rect 1535 5388 1539 5392
rect 1671 5388 1675 5392
rect 1807 5388 1811 5392
rect 1935 5389 1939 5393
rect 1975 5392 1979 5396
rect 2451 5391 2455 5395
rect 2699 5391 2703 5395
rect 2947 5391 2951 5395
rect 3187 5391 3191 5395
rect 3427 5391 3431 5395
rect 3651 5391 3655 5395
rect 3799 5392 3803 5396
rect 3839 5383 3843 5387
rect 4455 5384 4459 5388
rect 4615 5384 4619 5388
rect 4775 5384 4779 5388
rect 4935 5384 4939 5388
rect 5103 5384 5107 5388
rect 5663 5383 5667 5387
rect 111 5372 115 5376
rect 691 5373 695 5377
rect 827 5373 831 5377
rect 963 5373 967 5377
rect 1099 5373 1103 5377
rect 1235 5373 1239 5377
rect 1371 5373 1375 5377
rect 1507 5373 1511 5377
rect 1643 5373 1647 5377
rect 1779 5373 1783 5377
rect 1935 5372 1939 5376
rect 1975 5375 1979 5379
rect 2479 5376 2483 5380
rect 2727 5376 2731 5380
rect 2975 5376 2979 5380
rect 3215 5376 3219 5380
rect 3455 5376 3459 5380
rect 3679 5376 3683 5380
rect 3799 5375 3803 5379
rect 811 5363 815 5367
rect 1387 5363 1391 5367
rect 1475 5363 1479 5367
rect 1659 5363 1663 5367
rect 1795 5363 1799 5367
rect 1187 5351 1191 5355
rect 1187 5331 1191 5335
rect 1271 5331 1275 5335
rect 1387 5331 1391 5335
rect 1559 5331 1563 5335
rect 1659 5331 1663 5335
rect 1795 5331 1799 5335
rect 1975 5317 1979 5321
rect 2319 5316 2323 5320
rect 2519 5316 2523 5320
rect 2719 5316 2723 5320
rect 2919 5316 2923 5320
rect 3119 5316 3123 5320
rect 3327 5316 3331 5320
rect 3535 5316 3539 5320
rect 3799 5317 3803 5321
rect 3839 5317 3843 5321
rect 4431 5316 4435 5320
rect 4615 5316 4619 5320
rect 4799 5316 4803 5320
rect 4983 5316 4987 5320
rect 5175 5316 5179 5320
rect 5663 5317 5667 5321
rect 1975 5300 1979 5304
rect 2291 5301 2295 5305
rect 2491 5301 2495 5305
rect 2691 5301 2695 5305
rect 2891 5301 2895 5305
rect 3091 5301 3095 5305
rect 3299 5301 3303 5305
rect 3507 5301 3511 5305
rect 3799 5300 3803 5304
rect 3839 5300 3843 5304
rect 4403 5301 4407 5305
rect 4587 5301 4591 5305
rect 4771 5301 4775 5305
rect 4955 5301 4959 5305
rect 5147 5301 5151 5305
rect 5663 5300 5667 5304
rect 2419 5291 2420 5295
rect 2420 5291 2423 5295
rect 2707 5291 2711 5295
rect 811 5279 815 5283
rect 851 5283 855 5287
rect 1003 5283 1007 5287
rect 1155 5283 1159 5287
rect 1475 5283 1479 5287
rect 2379 5283 2383 5287
rect 3035 5291 3039 5295
rect 3315 5291 3319 5295
rect 3411 5291 3415 5295
rect 3179 5283 3183 5287
rect 4515 5291 4519 5295
rect 4567 5291 4571 5295
rect 4947 5291 4951 5295
rect 2379 5259 2383 5263
rect 2579 5259 2583 5263
rect 2707 5259 2711 5263
rect 2979 5259 2983 5263
rect 3179 5259 3183 5263
rect 3315 5259 3319 5263
rect 3551 5259 3555 5263
rect 4567 5259 4571 5263
rect 4603 5259 4607 5263
rect 4947 5259 4951 5263
rect 5199 5259 5203 5263
rect 851 5247 852 5251
rect 852 5247 855 5251
rect 1003 5247 1004 5251
rect 1004 5247 1007 5251
rect 1155 5247 1156 5251
rect 1156 5247 1159 5251
rect 1259 5247 1263 5251
rect 1647 5247 1648 5251
rect 1648 5247 1651 5251
rect 111 5240 115 5244
rect 723 5239 727 5243
rect 875 5239 879 5243
rect 1027 5239 1031 5243
rect 1187 5239 1191 5243
rect 1355 5239 1359 5243
rect 1523 5239 1527 5243
rect 1935 5240 1939 5244
rect 111 5223 115 5227
rect 751 5224 755 5228
rect 903 5224 907 5228
rect 1055 5224 1059 5228
rect 1215 5224 1219 5228
rect 1383 5224 1387 5228
rect 1551 5224 1555 5228
rect 1935 5223 1939 5227
rect 2363 5203 2367 5207
rect 2403 5207 2407 5211
rect 2771 5203 2775 5207
rect 2811 5207 2815 5211
rect 3411 5207 3415 5211
rect 4427 5195 4431 5199
rect 2403 5171 2404 5175
rect 2404 5171 2407 5175
rect 2579 5171 2583 5175
rect 2811 5171 2812 5175
rect 2812 5171 2815 5175
rect 2979 5171 2983 5175
rect 3079 5171 3083 5175
rect 111 5165 115 5169
rect 447 5164 451 5168
rect 623 5164 627 5168
rect 807 5164 811 5168
rect 999 5164 1003 5168
rect 1199 5164 1203 5168
rect 1399 5164 1403 5168
rect 1607 5164 1611 5168
rect 1815 5164 1819 5168
rect 1935 5165 1939 5169
rect 1975 5164 1979 5168
rect 2275 5163 2279 5167
rect 2475 5163 2479 5167
rect 2683 5163 2687 5167
rect 2891 5163 2895 5167
rect 3099 5163 3103 5167
rect 3307 5163 3311 5167
rect 3799 5164 3803 5168
rect 4603 5159 4607 5163
rect 5603 5159 5607 5163
rect 111 5148 115 5152
rect 419 5149 423 5153
rect 595 5149 599 5153
rect 779 5149 783 5153
rect 971 5149 975 5153
rect 1171 5149 1175 5153
rect 1371 5149 1375 5153
rect 1579 5149 1583 5153
rect 1787 5149 1791 5153
rect 1935 5148 1939 5152
rect 1975 5147 1979 5151
rect 2303 5148 2307 5152
rect 2503 5148 2507 5152
rect 2711 5148 2715 5152
rect 2919 5148 2923 5152
rect 3127 5148 3131 5152
rect 3839 5152 3843 5156
rect 3335 5148 3339 5152
rect 4435 5151 4439 5155
rect 3799 5147 3803 5151
rect 4595 5151 4599 5155
rect 4755 5151 4759 5155
rect 4915 5151 4919 5155
rect 5067 5151 5071 5155
rect 5219 5151 5223 5155
rect 5379 5151 5383 5155
rect 5515 5151 5519 5155
rect 5663 5152 5667 5156
rect 611 5139 615 5143
rect 715 5139 719 5143
rect 735 5139 739 5143
rect 1143 5139 1147 5143
rect 1491 5139 1495 5143
rect 1803 5139 1807 5143
rect 1459 5131 1463 5135
rect 3839 5135 3843 5139
rect 4463 5136 4467 5140
rect 4623 5136 4627 5140
rect 4783 5136 4787 5140
rect 4943 5136 4947 5140
rect 5095 5136 5099 5140
rect 5247 5136 5251 5140
rect 5407 5136 5411 5140
rect 5543 5136 5547 5140
rect 5663 5135 5667 5139
rect 611 5107 615 5111
rect 1143 5107 1147 5111
rect 1259 5107 1263 5111
rect 1459 5107 1463 5111
rect 1647 5107 1651 5111
rect 1803 5107 1807 5111
rect 735 5091 739 5095
rect 275 5075 279 5079
rect 1319 5075 1323 5079
rect 1975 5073 1979 5077
rect 2119 5072 2123 5076
rect 2327 5072 2331 5076
rect 2535 5072 2539 5076
rect 2751 5072 2755 5076
rect 2975 5072 2979 5076
rect 3207 5072 3211 5076
rect 3799 5073 3803 5077
rect 3839 5069 3843 5073
rect 3887 5068 3891 5072
rect 4087 5068 4091 5072
rect 4327 5068 4331 5072
rect 4567 5068 4571 5072
rect 4815 5068 4819 5072
rect 5063 5068 5067 5072
rect 5311 5068 5315 5072
rect 5543 5068 5547 5072
rect 5663 5069 5667 5073
rect 1975 5056 1979 5060
rect 2091 5057 2095 5061
rect 2299 5057 2303 5061
rect 2507 5057 2511 5061
rect 2723 5057 2727 5061
rect 2947 5057 2951 5061
rect 3179 5057 3183 5061
rect 3799 5056 3803 5060
rect 275 5051 279 5055
rect 283 5051 287 5055
rect 715 5047 719 5051
rect 755 5051 759 5055
rect 1119 5051 1123 5055
rect 1491 5051 1495 5055
rect 1627 5051 1631 5055
rect 3839 5052 3843 5056
rect 3859 5053 3863 5057
rect 4059 5053 4063 5057
rect 4299 5053 4303 5057
rect 4539 5053 4543 5057
rect 4787 5053 4791 5057
rect 5035 5053 5039 5057
rect 5283 5053 5287 5057
rect 5515 5053 5519 5057
rect 5663 5052 5667 5056
rect 2355 5047 2359 5051
rect 2179 5039 2183 5043
rect 2771 5047 2775 5051
rect 3195 5047 3199 5051
rect 4075 5043 4079 5047
rect 4219 5043 4223 5047
rect 4427 5043 4428 5047
rect 4428 5043 4431 5047
rect 4459 5043 4463 5047
rect 4683 5043 4687 5047
rect 5299 5043 5303 5047
rect 5371 5043 5375 5047
rect 5123 5035 5127 5039
rect 283 5015 284 5019
rect 284 5015 287 5019
rect 491 5015 495 5019
rect 755 5015 756 5019
rect 756 5015 759 5019
rect 1119 5015 1123 5019
rect 1319 5015 1320 5019
rect 1320 5015 1323 5019
rect 1627 5015 1628 5019
rect 1628 5015 1631 5019
rect 2179 5015 2183 5019
rect 111 5008 115 5012
rect 155 5007 159 5011
rect 379 5007 383 5011
rect 627 5007 631 5011
rect 899 5007 903 5011
rect 1195 5007 1199 5011
rect 1499 5007 1503 5011
rect 1787 5007 1791 5011
rect 1935 5008 1939 5012
rect 2839 4999 2843 5003
rect 3079 5015 3083 5019
rect 3195 5015 3199 5019
rect 4067 5011 4071 5015
rect 4075 5011 4079 5015
rect 4459 5011 4463 5015
rect 4683 5011 4687 5015
rect 4875 5011 4879 5015
rect 5123 5011 5127 5015
rect 5299 5011 5303 5015
rect 5603 5011 5607 5015
rect 3247 4999 3251 5003
rect 111 4991 115 4995
rect 183 4992 187 4996
rect 407 4992 411 4996
rect 655 4992 659 4996
rect 927 4992 931 4996
rect 1223 4992 1227 4996
rect 1527 4992 1531 4996
rect 1815 4992 1819 4996
rect 1935 4991 1939 4995
rect 2395 4959 2399 4963
rect 2547 4959 2551 4963
rect 2747 4959 2751 4963
rect 2963 4959 2967 4963
rect 3791 4963 3795 4967
rect 3987 4963 3991 4967
rect 3739 4955 3743 4959
rect 4219 4959 4223 4963
rect 4803 4963 4807 4967
rect 5211 4963 5215 4967
rect 5371 4963 5375 4967
rect 2395 4923 2396 4927
rect 2396 4923 2399 4927
rect 2547 4923 2548 4927
rect 2548 4923 2551 4927
rect 2747 4923 2748 4927
rect 2748 4923 2751 4927
rect 2839 4923 2843 4927
rect 3247 4923 3248 4927
rect 3248 4923 3251 4927
rect 3459 4923 3463 4927
rect 3791 4923 3795 4927
rect 3987 4927 3988 4931
rect 3988 4927 3991 4931
rect 4067 4927 4071 4931
rect 4803 4927 4804 4931
rect 4804 4927 4807 4931
rect 5211 4927 5212 4931
rect 5212 4927 5215 4931
rect 5239 4927 5243 4931
rect 5603 4927 5607 4931
rect 1975 4916 1979 4920
rect 1995 4915 1999 4919
rect 2131 4915 2135 4919
rect 2267 4915 2271 4919
rect 2419 4915 2423 4919
rect 2619 4915 2623 4919
rect 2859 4915 2863 4919
rect 3123 4915 3127 4919
rect 3395 4915 3399 4919
rect 3651 4915 3655 4919
rect 3799 4916 3803 4920
rect 3839 4920 3843 4924
rect 3859 4919 3863 4923
rect 3995 4919 3999 4923
rect 4131 4919 4135 4923
rect 4267 4919 4271 4923
rect 4403 4919 4407 4923
rect 4539 4919 4543 4923
rect 4675 4919 4679 4923
rect 4811 4919 4815 4923
rect 4947 4919 4951 4923
rect 5083 4919 5087 4923
rect 5227 4919 5231 4923
rect 5379 4919 5383 4923
rect 5515 4919 5519 4923
rect 5663 4920 5667 4924
rect 111 4905 115 4909
rect 159 4904 163 4908
rect 295 4904 299 4908
rect 431 4904 435 4908
rect 567 4904 571 4908
rect 703 4904 707 4908
rect 1935 4905 1939 4909
rect 1975 4899 1979 4903
rect 2023 4900 2027 4904
rect 2159 4900 2163 4904
rect 2295 4900 2299 4904
rect 2447 4900 2451 4904
rect 2647 4900 2651 4904
rect 2887 4900 2891 4904
rect 3151 4900 3155 4904
rect 3423 4900 3427 4904
rect 3679 4900 3683 4904
rect 3799 4899 3803 4903
rect 3839 4903 3843 4907
rect 3887 4904 3891 4908
rect 4023 4904 4027 4908
rect 4159 4904 4163 4908
rect 4295 4904 4299 4908
rect 4431 4904 4435 4908
rect 4567 4904 4571 4908
rect 4703 4904 4707 4908
rect 4839 4904 4843 4908
rect 4975 4904 4979 4908
rect 5111 4904 5115 4908
rect 5255 4904 5259 4908
rect 5407 4904 5411 4908
rect 5543 4904 5547 4908
rect 5663 4903 5667 4907
rect 111 4888 115 4892
rect 131 4889 135 4893
rect 267 4889 271 4893
rect 403 4889 407 4893
rect 539 4889 543 4893
rect 675 4889 679 4893
rect 1935 4888 1939 4892
rect 235 4879 239 4883
rect 555 4879 559 4883
rect 691 4879 695 4883
rect 355 4871 359 4875
rect 355 4847 359 4851
rect 491 4847 495 4851
rect 555 4847 559 4851
rect 691 4847 695 4851
rect 1975 4833 1979 4837
rect 2327 4832 2331 4836
rect 2559 4832 2563 4836
rect 2823 4832 2827 4836
rect 3103 4832 3107 4836
rect 3399 4832 3403 4836
rect 3679 4832 3683 4836
rect 3799 4833 3803 4837
rect 1975 4816 1979 4820
rect 2299 4817 2303 4821
rect 2531 4817 2535 4821
rect 2795 4817 2799 4821
rect 3075 4817 3079 4821
rect 3371 4817 3375 4821
rect 3651 4817 3655 4821
rect 3799 4816 3803 4820
rect 2547 4807 2551 4811
rect 2811 4807 2815 4811
rect 2963 4807 2967 4811
rect 2667 4799 2671 4803
rect 3739 4807 3743 4811
rect 235 4787 239 4791
rect 259 4787 263 4791
rect 395 4787 399 4791
rect 531 4787 535 4791
rect 667 4787 671 4791
rect 2387 4775 2391 4779
rect 2547 4775 2551 4779
rect 2811 4775 2815 4779
rect 3459 4775 3463 4779
rect 3739 4775 3743 4779
rect 3839 4769 3843 4773
rect 3887 4768 3891 4772
rect 4071 4768 4075 4772
rect 4295 4768 4299 4772
rect 4535 4768 4539 4772
rect 4783 4768 4787 4772
rect 5039 4768 5043 4772
rect 5303 4768 5307 4772
rect 5543 4768 5547 4772
rect 5663 4769 5667 4773
rect 219 4759 223 4763
rect 259 4751 260 4755
rect 260 4751 263 4755
rect 395 4751 396 4755
rect 396 4751 399 4755
rect 531 4751 532 4755
rect 532 4751 535 4755
rect 667 4751 668 4755
rect 668 4751 671 4755
rect 3839 4752 3843 4756
rect 3859 4753 3863 4757
rect 4043 4753 4047 4757
rect 4267 4753 4271 4757
rect 4507 4753 4511 4757
rect 4755 4753 4759 4757
rect 5011 4753 5015 4757
rect 5275 4753 5279 4757
rect 5515 4753 5519 4757
rect 5663 4752 5667 4756
rect 111 4744 115 4748
rect 131 4743 135 4747
rect 267 4743 271 4747
rect 403 4743 407 4747
rect 539 4743 543 4747
rect 675 4743 679 4747
rect 1935 4744 1939 4748
rect 3739 4743 3743 4747
rect 4003 4743 4007 4747
rect 4523 4743 4527 4747
rect 4771 4743 4775 4747
rect 4131 4735 4135 4739
rect 5291 4743 5295 4747
rect 5371 4743 5375 4747
rect 5099 4735 5103 4739
rect 111 4727 115 4731
rect 159 4728 163 4732
rect 295 4728 299 4732
rect 431 4728 435 4732
rect 567 4728 571 4732
rect 703 4728 707 4732
rect 1935 4727 1939 4731
rect 2107 4711 2111 4715
rect 2147 4715 2151 4719
rect 2323 4715 2327 4719
rect 2667 4715 2671 4719
rect 2675 4715 2679 4719
rect 4003 4711 4007 4715
rect 4131 4711 4135 4715
rect 4139 4711 4143 4715
rect 4523 4711 4527 4715
rect 4771 4711 4775 4715
rect 5099 4711 5103 4715
rect 5291 4711 5295 4715
rect 5603 4711 5607 4715
rect 2147 4679 2148 4683
rect 2148 4679 2151 4683
rect 2323 4679 2324 4683
rect 2324 4679 2327 4683
rect 2387 4679 2391 4683
rect 2675 4679 2676 4683
rect 2676 4679 2679 4683
rect 2835 4679 2839 4683
rect 1975 4672 1979 4676
rect 2019 4671 2023 4675
rect 2195 4671 2199 4675
rect 2371 4671 2375 4675
rect 2547 4671 2551 4675
rect 2723 4671 2727 4675
rect 3799 4672 3803 4676
rect 111 4665 115 4669
rect 159 4664 163 4668
rect 295 4664 299 4668
rect 431 4664 435 4668
rect 567 4664 571 4668
rect 703 4664 707 4668
rect 1935 4665 1939 4669
rect 3779 4663 3783 4667
rect 3987 4663 3991 4667
rect 1975 4655 1979 4659
rect 2047 4656 2051 4660
rect 2223 4656 2227 4660
rect 2399 4656 2403 4660
rect 2575 4656 2579 4660
rect 2751 4656 2755 4660
rect 3799 4655 3803 4659
rect 4219 4659 4223 4663
rect 4259 4663 4263 4667
rect 4395 4663 4399 4667
rect 5331 4659 5335 4663
rect 5371 4663 5375 4667
rect 111 4648 115 4652
rect 131 4649 135 4653
rect 267 4649 271 4653
rect 403 4649 407 4653
rect 539 4649 543 4653
rect 675 4649 679 4653
rect 1935 4648 1939 4652
rect 283 4639 287 4643
rect 419 4639 423 4643
rect 555 4639 559 4643
rect 691 4639 695 4643
rect 755 4639 759 4643
rect 4219 4635 4223 4639
rect 5331 4635 5335 4639
rect 3987 4627 3988 4631
rect 3988 4627 3991 4631
rect 4139 4627 4143 4631
rect 4259 4627 4260 4631
rect 4260 4627 4263 4631
rect 4395 4627 4396 4631
rect 4396 4627 4399 4631
rect 4595 4627 4599 4631
rect 3839 4620 3843 4624
rect 3859 4619 3863 4623
rect 3995 4619 3999 4623
rect 4131 4619 4135 4623
rect 4267 4619 4271 4623
rect 4403 4619 4407 4623
rect 4539 4619 4543 4623
rect 4675 4619 4679 4623
rect 4819 4619 4823 4623
rect 4963 4619 4967 4623
rect 5107 4619 5111 4623
rect 5243 4619 5247 4623
rect 5379 4619 5383 4623
rect 5515 4619 5519 4623
rect 5663 4620 5667 4624
rect 219 4607 223 4611
rect 283 4607 287 4611
rect 419 4607 423 4611
rect 555 4607 559 4611
rect 691 4607 695 4611
rect 3839 4603 3843 4607
rect 3887 4604 3891 4608
rect 4023 4604 4027 4608
rect 4159 4604 4163 4608
rect 4295 4604 4299 4608
rect 4431 4604 4435 4608
rect 4567 4604 4571 4608
rect 4703 4604 4707 4608
rect 4847 4604 4851 4608
rect 4991 4604 4995 4608
rect 5135 4604 5139 4608
rect 5271 4604 5275 4608
rect 5407 4604 5411 4608
rect 5543 4604 5547 4608
rect 5663 4603 5667 4607
rect 1975 4593 1979 4597
rect 2023 4592 2027 4596
rect 2263 4592 2267 4596
rect 2527 4592 2531 4596
rect 2775 4592 2779 4596
rect 3015 4592 3019 4596
rect 3247 4592 3251 4596
rect 3471 4592 3475 4596
rect 3679 4592 3683 4596
rect 3799 4593 3803 4597
rect 1975 4576 1979 4580
rect 1995 4577 1999 4581
rect 2235 4577 2239 4581
rect 2499 4577 2503 4581
rect 2747 4577 2751 4581
rect 2987 4577 2991 4581
rect 3219 4577 3223 4581
rect 3443 4577 3447 4581
rect 3651 4577 3655 4581
rect 3799 4576 3803 4580
rect 579 4567 583 4571
rect 1223 4567 1227 4571
rect 2107 4567 2111 4571
rect 2515 4567 2519 4571
rect 2619 4567 2623 4571
rect 755 4559 759 4563
rect 2323 4559 2327 4563
rect 3235 4567 3239 4571
rect 3459 4567 3463 4571
rect 3667 4567 3671 4571
rect 3779 4567 3780 4571
rect 3780 4567 3783 4571
rect 379 4547 383 4551
rect 567 4547 571 4551
rect 779 4547 783 4551
rect 1003 4547 1007 4551
rect 1523 4547 1527 4551
rect 3839 4545 3843 4549
rect 4671 4544 4675 4548
rect 4807 4544 4811 4548
rect 4943 4544 4947 4548
rect 5079 4544 5083 4548
rect 5663 4545 5667 4549
rect 1563 4539 1567 4543
rect 2011 4535 2015 4539
rect 2323 4535 2327 4539
rect 2515 4535 2519 4539
rect 2835 4535 2839 4539
rect 3075 4535 3079 4539
rect 3235 4535 3239 4539
rect 3459 4535 3463 4539
rect 3667 4535 3671 4539
rect 3839 4528 3843 4532
rect 4643 4529 4647 4533
rect 4779 4529 4783 4533
rect 4915 4529 4919 4533
rect 5051 4529 5055 4533
rect 5663 4528 5667 4532
rect 4795 4519 4799 4523
rect 4931 4519 4935 4523
rect 5067 4519 5071 4523
rect 5075 4519 5079 4523
rect 379 4511 380 4515
rect 380 4511 383 4515
rect 567 4511 568 4515
rect 568 4511 571 4515
rect 779 4511 780 4515
rect 780 4511 783 4515
rect 1003 4511 1004 4515
rect 1004 4511 1007 4515
rect 1223 4511 1224 4515
rect 1224 4511 1227 4515
rect 1523 4511 1527 4515
rect 2011 4511 2015 4515
rect 111 4504 115 4508
rect 251 4503 255 4507
rect 443 4503 447 4507
rect 651 4503 655 4507
rect 875 4503 879 4507
rect 1099 4503 1103 4507
rect 1331 4503 1335 4507
rect 1571 4503 1575 4507
rect 1787 4503 1791 4507
rect 1935 4504 1939 4508
rect 111 4487 115 4491
rect 279 4488 283 4492
rect 471 4488 475 4492
rect 679 4488 683 4492
rect 903 4488 907 4492
rect 1127 4488 1131 4492
rect 1359 4488 1363 4492
rect 1599 4488 1603 4492
rect 1815 4488 1819 4492
rect 1935 4487 1939 4491
rect 4595 4487 4599 4491
rect 4795 4487 4799 4491
rect 4931 4487 4935 4491
rect 5067 4487 5071 4491
rect 2495 4475 2499 4479
rect 2619 4475 2623 4479
rect 2835 4471 2839 4475
rect 2875 4475 2879 4479
rect 3099 4475 3103 4479
rect 3315 4475 3319 4479
rect 3523 4475 3527 4479
rect 2391 4439 2392 4443
rect 2392 4439 2395 4443
rect 2495 4439 2499 4443
rect 2875 4439 2876 4443
rect 2876 4439 2879 4443
rect 3099 4439 3100 4443
rect 3100 4439 3103 4443
rect 3315 4439 3316 4443
rect 3316 4439 3319 4443
rect 3523 4439 3524 4443
rect 3524 4439 3527 4443
rect 3735 4439 3736 4443
rect 3736 4439 3739 4443
rect 111 4429 115 4433
rect 511 4428 515 4432
rect 687 4428 691 4432
rect 871 4428 875 4432
rect 1071 4428 1075 4432
rect 1279 4428 1283 4432
rect 1495 4428 1499 4432
rect 1719 4428 1723 4432
rect 1935 4429 1939 4433
rect 1975 4432 1979 4436
rect 2267 4431 2271 4435
rect 2515 4431 2519 4435
rect 2747 4431 2751 4435
rect 2971 4431 2975 4435
rect 3187 4431 3191 4435
rect 3395 4431 3399 4435
rect 3611 4431 3615 4435
rect 3799 4432 3803 4436
rect 5075 4435 5079 4439
rect 111 4412 115 4416
rect 483 4413 487 4417
rect 659 4413 663 4417
rect 843 4413 847 4417
rect 1043 4413 1047 4417
rect 1251 4413 1255 4417
rect 1467 4413 1471 4417
rect 1691 4413 1695 4417
rect 1935 4412 1939 4416
rect 1975 4415 1979 4419
rect 2295 4416 2299 4420
rect 2543 4416 2547 4420
rect 2775 4416 2779 4420
rect 2999 4416 3003 4420
rect 3215 4416 3219 4420
rect 3423 4416 3427 4420
rect 3639 4416 3643 4420
rect 3799 4415 3803 4419
rect 675 4403 679 4407
rect 859 4403 863 4407
rect 1059 4403 1063 4407
rect 1267 4403 1271 4407
rect 1363 4403 1367 4407
rect 1563 4403 1567 4407
rect 1611 4403 1615 4407
rect 4467 4399 4471 4403
rect 3839 4392 3843 4396
rect 4347 4391 4351 4395
rect 4483 4391 4487 4395
rect 4619 4391 4623 4395
rect 4755 4391 4759 4395
rect 4891 4391 4895 4395
rect 5663 4392 5667 4396
rect 579 4371 583 4375
rect 675 4371 679 4375
rect 859 4371 863 4375
rect 1059 4371 1063 4375
rect 1267 4371 1271 4375
rect 1611 4371 1615 4375
rect 1779 4371 1783 4375
rect 3839 4375 3843 4379
rect 4375 4376 4379 4380
rect 4511 4376 4515 4380
rect 4647 4376 4651 4380
rect 4783 4376 4787 4380
rect 4919 4376 4923 4380
rect 5663 4375 5667 4379
rect 1975 4345 1979 4349
rect 2023 4344 2027 4348
rect 2199 4344 2203 4348
rect 2399 4344 2403 4348
rect 2591 4344 2595 4348
rect 2775 4344 2779 4348
rect 2951 4344 2955 4348
rect 3135 4344 3139 4348
rect 3319 4344 3323 4348
rect 3799 4345 3803 4349
rect 1363 4331 1367 4335
rect 1975 4328 1979 4332
rect 1995 4329 1999 4333
rect 2171 4329 2175 4333
rect 2371 4329 2375 4333
rect 2563 4329 2567 4333
rect 2747 4329 2751 4333
rect 2923 4329 2927 4333
rect 3107 4329 3111 4333
rect 3291 4329 3295 4333
rect 3799 4328 3803 4332
rect 1523 4319 1527 4323
rect 1659 4319 1663 4323
rect 2099 4319 2103 4323
rect 2311 4319 2315 4323
rect 2763 4319 2767 4323
rect 2939 4319 2943 4323
rect 3123 4319 3127 4323
rect 3307 4319 3311 4323
rect 2835 4311 2839 4315
rect 1619 4303 1623 4307
rect 3839 4301 3843 4305
rect 4135 4300 4139 4304
rect 4271 4300 4275 4304
rect 4407 4300 4411 4304
rect 4543 4300 4547 4304
rect 4679 4300 4683 4304
rect 5663 4301 5667 4305
rect 1331 4283 1335 4287
rect 1523 4283 1524 4287
rect 1524 4283 1527 4287
rect 1659 4283 1660 4287
rect 1660 4283 1663 4287
rect 1779 4283 1783 4287
rect 2311 4287 2315 4291
rect 2391 4287 2395 4291
rect 2631 4287 2635 4291
rect 2763 4287 2767 4291
rect 2939 4287 2943 4291
rect 3123 4287 3127 4291
rect 3307 4287 3311 4291
rect 3839 4284 3843 4288
rect 4107 4285 4111 4289
rect 4243 4285 4247 4289
rect 4379 4285 4383 4289
rect 4515 4285 4519 4289
rect 4651 4285 4655 4289
rect 5663 4284 5667 4288
rect 111 4276 115 4280
rect 715 4275 719 4279
rect 851 4275 855 4279
rect 987 4275 991 4279
rect 1123 4275 1127 4279
rect 1259 4275 1263 4279
rect 1395 4275 1399 4279
rect 1531 4275 1535 4279
rect 1667 4275 1671 4279
rect 1935 4276 1939 4280
rect 4235 4275 4236 4279
rect 4236 4275 4239 4279
rect 4251 4275 4255 4279
rect 4531 4275 4535 4279
rect 4667 4275 4671 4279
rect 4331 4267 4335 4271
rect 111 4259 115 4263
rect 743 4260 747 4264
rect 879 4260 883 4264
rect 1015 4260 1019 4264
rect 1151 4260 1155 4264
rect 1287 4260 1291 4264
rect 1423 4260 1427 4264
rect 1559 4260 1563 4264
rect 1695 4260 1699 4264
rect 1935 4259 1939 4263
rect 4251 4243 4255 4247
rect 4331 4243 4335 4247
rect 4467 4243 4471 4247
rect 4531 4243 4535 4247
rect 4667 4243 4671 4247
rect 2099 4235 2103 4239
rect 2331 4231 2335 4235
rect 2959 4235 2963 4239
rect 3371 4231 3375 4235
rect 2331 4207 2335 4211
rect 1947 4199 1951 4203
rect 2631 4199 2632 4203
rect 2632 4199 2635 4203
rect 2959 4199 2963 4203
rect 111 4193 115 4197
rect 727 4192 731 4196
rect 863 4192 867 4196
rect 999 4192 1003 4196
rect 1135 4192 1139 4196
rect 1271 4192 1275 4196
rect 1407 4192 1411 4196
rect 1543 4192 1547 4196
rect 1679 4192 1683 4196
rect 1815 4192 1819 4196
rect 1935 4193 1939 4197
rect 1975 4192 1979 4196
rect 1995 4191 1999 4195
rect 2243 4191 2247 4195
rect 2507 4191 2511 4195
rect 2763 4191 2767 4195
rect 3019 4191 3023 4195
rect 3283 4191 3287 4195
rect 3799 4192 3803 4196
rect 111 4176 115 4180
rect 699 4177 703 4181
rect 835 4177 839 4181
rect 971 4177 975 4181
rect 1107 4177 1111 4181
rect 1243 4177 1247 4181
rect 1379 4177 1383 4181
rect 1515 4177 1519 4181
rect 1651 4177 1655 4181
rect 1787 4177 1791 4181
rect 1935 4176 1939 4180
rect 1975 4175 1979 4179
rect 2023 4176 2027 4180
rect 2271 4176 2275 4180
rect 2535 4176 2539 4180
rect 2791 4176 2795 4180
rect 3047 4176 3051 4180
rect 3311 4176 3315 4180
rect 3799 4175 3803 4179
rect 4059 4179 4063 4183
rect 4235 4183 4239 4187
rect 851 4167 855 4171
rect 963 4167 964 4171
rect 964 4167 967 4171
rect 787 4159 791 4163
rect 1531 4167 1535 4171
rect 1619 4167 1623 4171
rect 1779 4167 1780 4171
rect 1780 4167 1783 4171
rect 1795 4167 1799 4171
rect 4283 4147 4287 4151
rect 4523 4147 4527 4151
rect 3839 4140 3843 4144
rect 787 4135 791 4139
rect 851 4135 855 4139
rect 1331 4135 1335 4139
rect 1467 4135 1471 4139
rect 1531 4135 1535 4139
rect 1795 4135 1799 4139
rect 3971 4139 3975 4143
rect 1947 4135 1951 4139
rect 4107 4139 4111 4143
rect 4243 4139 4247 4143
rect 4379 4139 4383 4143
rect 4515 4139 4519 4143
rect 5663 4140 5667 4144
rect 3839 4123 3843 4127
rect 3999 4124 4003 4128
rect 4135 4124 4139 4128
rect 4271 4124 4275 4128
rect 4407 4124 4411 4128
rect 4543 4124 4547 4128
rect 5663 4123 5667 4127
rect 1975 4105 1979 4109
rect 3135 4104 3139 4108
rect 3271 4104 3275 4108
rect 3407 4104 3411 4108
rect 3543 4104 3547 4108
rect 3679 4104 3683 4108
rect 3799 4105 3803 4109
rect 651 4083 655 4087
rect 963 4087 967 4091
rect 1779 4087 1783 4091
rect 1975 4088 1979 4092
rect 3107 4089 3111 4093
rect 3243 4089 3247 4093
rect 3379 4089 3383 4093
rect 3515 4089 3519 4093
rect 3651 4089 3655 4093
rect 3799 4088 3803 4092
rect 3259 4079 3263 4083
rect 3371 4079 3372 4083
rect 3372 4079 3375 4083
rect 1475 4071 1479 4075
rect 3195 4071 3199 4075
rect 651 4059 655 4063
rect 959 4051 960 4055
rect 960 4051 963 4055
rect 1467 4051 1471 4055
rect 1639 4051 1640 4055
rect 1640 4051 1643 4055
rect 111 4044 115 4048
rect 563 4043 567 4047
rect 699 4043 703 4047
rect 835 4043 839 4047
rect 971 4043 975 4047
rect 1107 4043 1111 4047
rect 1243 4043 1247 4047
rect 1379 4043 1383 4047
rect 1515 4043 1519 4047
rect 1651 4043 1655 4047
rect 1787 4043 1791 4047
rect 1935 4044 1939 4048
rect 3195 4047 3199 4051
rect 3259 4047 3263 4051
rect 3739 4047 3743 4051
rect 3839 4041 3843 4045
rect 3887 4040 3891 4044
rect 4023 4040 4027 4044
rect 4159 4040 4163 4044
rect 4295 4040 4299 4044
rect 4431 4040 4435 4044
rect 4567 4040 4571 4044
rect 4703 4040 4707 4044
rect 4839 4040 4843 4044
rect 5663 4041 5667 4045
rect 111 4027 115 4031
rect 591 4028 595 4032
rect 727 4028 731 4032
rect 863 4028 867 4032
rect 999 4028 1003 4032
rect 1135 4028 1139 4032
rect 1271 4028 1275 4032
rect 1407 4028 1411 4032
rect 1543 4028 1547 4032
rect 1679 4028 1683 4032
rect 1815 4028 1819 4032
rect 1935 4027 1939 4031
rect 3839 4024 3843 4028
rect 3859 4025 3863 4029
rect 3995 4025 3999 4029
rect 4131 4025 4135 4029
rect 4267 4025 4271 4029
rect 4403 4025 4407 4029
rect 4539 4025 4543 4029
rect 4675 4025 4679 4029
rect 4811 4025 4815 4029
rect 5663 4024 5667 4028
rect 3739 4015 3743 4019
rect 4003 4015 4007 4019
rect 4083 4007 4087 4011
rect 4419 4015 4423 4019
rect 4555 4015 4559 4019
rect 4691 4015 4695 4019
rect 4827 4015 4831 4019
rect 4003 3983 4007 3987
rect 4083 3983 4087 3987
rect 4123 3983 4127 3987
rect 4283 3983 4287 3987
rect 4419 3983 4423 3987
rect 4555 3983 4559 3987
rect 4691 3983 4695 3987
rect 4827 3983 4831 3987
rect 111 3969 115 3973
rect 159 3968 163 3972
rect 327 3968 331 3972
rect 535 3968 539 3972
rect 751 3968 755 3972
rect 967 3968 971 3972
rect 1183 3968 1187 3972
rect 1399 3968 1403 3972
rect 1615 3968 1619 3972
rect 1815 3968 1819 3972
rect 1935 3969 1939 3973
rect 111 3952 115 3956
rect 131 3953 135 3957
rect 299 3953 303 3957
rect 507 3953 511 3957
rect 723 3953 727 3957
rect 939 3953 943 3957
rect 1155 3953 1159 3957
rect 1371 3953 1375 3957
rect 1587 3953 1591 3957
rect 1787 3953 1791 3957
rect 1935 3952 1939 3956
rect 235 3943 239 3947
rect 287 3943 291 3947
rect 451 3943 455 3947
rect 703 3943 707 3947
rect 879 3943 883 3947
rect 1387 3943 1391 3947
rect 1475 3943 1479 3947
rect 1803 3943 1807 3947
rect 1891 3943 1895 3947
rect 3779 3935 3783 3939
rect 3987 3935 3991 3939
rect 4275 3935 4279 3939
rect 4451 3935 4455 3939
rect 4611 3935 4615 3939
rect 4771 3935 4775 3939
rect 287 3911 291 3915
rect 451 3911 455 3915
rect 703 3911 707 3915
rect 879 3911 883 3915
rect 959 3911 963 3915
rect 1243 3911 1247 3915
rect 1387 3911 1391 3915
rect 1639 3911 1643 3915
rect 1803 3911 1807 3915
rect 1915 3907 1919 3911
rect 2523 3907 2527 3911
rect 2531 3907 2535 3911
rect 2955 3907 2959 3911
rect 3379 3907 3383 3911
rect 3987 3899 3988 3903
rect 3988 3899 3991 3903
rect 4123 3899 4124 3903
rect 4124 3899 4127 3903
rect 4275 3899 4276 3903
rect 4276 3899 4279 3903
rect 4451 3899 4455 3903
rect 4611 3899 4615 3903
rect 4771 3899 4775 3903
rect 4787 3899 4791 3903
rect 3839 3892 3843 3896
rect 3859 3891 3863 3895
rect 3995 3891 3999 3895
rect 4147 3891 4151 3895
rect 4299 3891 4303 3895
rect 4459 3891 4463 3895
rect 4619 3891 4623 3895
rect 4779 3891 4783 3895
rect 5663 3892 5667 3896
rect 2083 3871 2087 3875
rect 2531 3871 2532 3875
rect 2532 3871 2535 3875
rect 2955 3871 2956 3875
rect 2956 3871 2959 3875
rect 3379 3871 3380 3875
rect 3380 3871 3383 3875
rect 3779 3871 3780 3875
rect 3780 3871 3783 3875
rect 3839 3875 3843 3879
rect 3887 3876 3891 3880
rect 4023 3876 4027 3880
rect 4175 3876 4179 3880
rect 4327 3876 4331 3880
rect 4487 3876 4491 3880
rect 4647 3876 4651 3880
rect 4807 3876 4811 3880
rect 5663 3875 5667 3879
rect 235 3863 239 3867
rect 259 3863 263 3867
rect 483 3863 487 3867
rect 747 3863 751 3867
rect 1335 3863 1339 3867
rect 1891 3863 1895 3867
rect 1975 3864 1979 3868
rect 1995 3863 1999 3867
rect 2403 3863 2407 3867
rect 2827 3863 2831 3867
rect 3251 3863 3255 3867
rect 3651 3863 3655 3867
rect 3799 3864 3803 3868
rect 1975 3847 1979 3851
rect 2023 3848 2027 3852
rect 2431 3848 2435 3852
rect 2855 3848 2859 3852
rect 3279 3848 3283 3852
rect 3679 3848 3683 3852
rect 3799 3847 3803 3851
rect 259 3827 260 3831
rect 260 3827 263 3831
rect 483 3827 484 3831
rect 484 3827 487 3831
rect 747 3827 748 3831
rect 748 3827 751 3831
rect 851 3827 855 3831
rect 1243 3827 1247 3831
rect 1335 3827 1339 3831
rect 1915 3827 1916 3831
rect 1916 3827 1919 3831
rect 2523 3831 2527 3835
rect 3655 3831 3659 3835
rect 111 3820 115 3824
rect 131 3819 135 3823
rect 355 3819 359 3823
rect 619 3819 623 3823
rect 899 3819 903 3823
rect 1195 3819 1199 3823
rect 1499 3819 1503 3823
rect 1787 3819 1791 3823
rect 1935 3820 1939 3824
rect 111 3803 115 3807
rect 159 3804 163 3808
rect 383 3804 387 3808
rect 647 3804 651 3808
rect 927 3804 931 3808
rect 1223 3804 1227 3808
rect 1527 3804 1531 3808
rect 1815 3804 1819 3808
rect 1935 3803 1939 3807
rect 1975 3789 1979 3793
rect 2023 3788 2027 3792
rect 2175 3788 2179 3792
rect 2351 3788 2355 3792
rect 2535 3788 2539 3792
rect 2719 3788 2723 3792
rect 2895 3788 2899 3792
rect 3071 3788 3075 3792
rect 3247 3788 3251 3792
rect 3423 3788 3427 3792
rect 3607 3788 3611 3792
rect 3799 3789 3803 3793
rect 3839 3789 3843 3793
rect 4503 3788 4507 3792
rect 4639 3788 4643 3792
rect 4775 3788 4779 3792
rect 4911 3788 4915 3792
rect 5047 3788 5051 3792
rect 5663 3789 5667 3793
rect 1975 3772 1979 3776
rect 1995 3773 1999 3777
rect 2147 3773 2151 3777
rect 2323 3773 2327 3777
rect 2507 3773 2511 3777
rect 2691 3773 2695 3777
rect 2867 3773 2871 3777
rect 3043 3773 3047 3777
rect 3219 3773 3223 3777
rect 3395 3773 3399 3777
rect 3579 3773 3583 3777
rect 3799 3772 3803 3776
rect 3839 3772 3843 3776
rect 4475 3773 4479 3777
rect 4611 3773 4615 3777
rect 4747 3773 4751 3777
rect 4883 3773 4887 3777
rect 5019 3773 5023 3777
rect 5663 3772 5667 3776
rect 2163 3763 2167 3767
rect 2339 3763 2343 3767
rect 2523 3763 2527 3767
rect 2707 3763 2711 3767
rect 3059 3763 3063 3767
rect 3235 3763 3239 3767
rect 3411 3763 3415 3767
rect 3595 3763 3599 3767
rect 3655 3763 3659 3767
rect 4627 3763 4631 3767
rect 4763 3763 4767 3767
rect 4899 3763 4903 3767
rect 5035 3763 5039 3767
rect 4123 3755 4127 3759
rect 111 3733 115 3737
rect 247 3732 251 3736
rect 519 3732 523 3736
rect 791 3732 795 3736
rect 1063 3732 1067 3736
rect 1343 3732 1347 3736
rect 1935 3733 1939 3737
rect 2083 3731 2087 3735
rect 2163 3731 2167 3735
rect 2339 3731 2343 3735
rect 2523 3731 2527 3735
rect 2707 3731 2711 3735
rect 111 3716 115 3720
rect 219 3717 223 3721
rect 491 3717 495 3721
rect 763 3717 767 3721
rect 1035 3717 1039 3721
rect 1315 3717 1319 3721
rect 1935 3716 1939 3720
rect 3059 3731 3063 3735
rect 3235 3731 3239 3735
rect 3411 3731 3415 3735
rect 3595 3731 3599 3735
rect 4787 3747 4791 3751
rect 4627 3731 4631 3735
rect 4763 3731 4767 3735
rect 4899 3731 4903 3735
rect 5035 3731 5039 3735
rect 3423 3715 3427 3719
rect 507 3707 511 3711
rect 595 3707 599 3711
rect 307 3699 311 3703
rect 1331 3707 1335 3711
rect 307 3675 311 3679
rect 507 3675 511 3679
rect 851 3675 855 3679
rect 1203 3675 1207 3679
rect 1331 3675 1335 3679
rect 2275 3675 2279 3679
rect 2419 3675 2423 3679
rect 2563 3675 2567 3679
rect 2851 3675 2855 3679
rect 2995 3675 2999 3679
rect 3283 3675 3287 3679
rect 2955 3659 2959 3663
rect 4123 3663 4127 3667
rect 4147 3663 4151 3667
rect 4283 3663 4287 3667
rect 4419 3663 4423 3667
rect 4555 3663 4559 3667
rect 4691 3663 4695 3667
rect 4827 3663 4831 3667
rect 2275 3639 2276 3643
rect 2276 3639 2279 3643
rect 2419 3639 2420 3643
rect 2420 3639 2423 3643
rect 2563 3639 2564 3643
rect 2564 3639 2567 3643
rect 2599 3639 2603 3643
rect 2851 3639 2852 3643
rect 2852 3639 2855 3643
rect 2995 3639 2996 3643
rect 2996 3639 2999 3643
rect 3283 3639 3284 3643
rect 3284 3639 3287 3643
rect 3423 3639 3424 3643
rect 3424 3639 3427 3643
rect 1975 3632 1979 3636
rect 2011 3631 2015 3635
rect 2147 3631 2151 3635
rect 2291 3631 2295 3635
rect 2435 3631 2439 3635
rect 2579 3631 2583 3635
rect 2723 3631 2727 3635
rect 2867 3631 2871 3635
rect 3011 3631 3015 3635
rect 3155 3631 3159 3635
rect 3299 3631 3303 3635
rect 3799 3632 3803 3636
rect 4147 3627 4148 3631
rect 4148 3627 4151 3631
rect 4283 3627 4284 3631
rect 4284 3627 4287 3631
rect 4419 3627 4420 3631
rect 4420 3627 4423 3631
rect 4555 3627 4556 3631
rect 4556 3627 4559 3631
rect 4691 3627 4692 3631
rect 4692 3627 4695 3631
rect 4827 3627 4828 3631
rect 4828 3627 4831 3631
rect 5551 3627 5555 3631
rect 595 3611 599 3615
rect 763 3611 767 3615
rect 1011 3607 1015 3611
rect 1051 3611 1055 3615
rect 1195 3611 1199 3615
rect 1975 3615 1979 3619
rect 2039 3616 2043 3620
rect 2175 3616 2179 3620
rect 2319 3616 2323 3620
rect 2463 3616 2467 3620
rect 2607 3616 2611 3620
rect 2751 3616 2755 3620
rect 2895 3616 2899 3620
rect 3039 3616 3043 3620
rect 3183 3616 3187 3620
rect 3839 3620 3843 3624
rect 3327 3616 3331 3620
rect 4019 3619 4023 3623
rect 3799 3615 3803 3619
rect 4155 3619 4159 3623
rect 4291 3619 4295 3623
rect 4427 3619 4431 3623
rect 4563 3619 4567 3623
rect 4699 3619 4703 3623
rect 4835 3619 4839 3623
rect 4971 3619 4975 3623
rect 5107 3619 5111 3623
rect 5243 3619 5247 3623
rect 5379 3619 5383 3623
rect 5515 3619 5519 3623
rect 5663 3620 5667 3624
rect 3839 3603 3843 3607
rect 4047 3604 4051 3608
rect 4183 3604 4187 3608
rect 4319 3604 4323 3608
rect 4455 3604 4459 3608
rect 4591 3604 4595 3608
rect 4727 3604 4731 3608
rect 4863 3604 4867 3608
rect 4999 3604 5003 3608
rect 5135 3604 5139 3608
rect 5271 3604 5275 3608
rect 5407 3604 5411 3608
rect 5543 3604 5547 3608
rect 5663 3603 5667 3607
rect 763 3575 764 3579
rect 764 3575 767 3579
rect 899 3575 903 3579
rect 1051 3575 1052 3579
rect 1052 3575 1055 3579
rect 1195 3575 1196 3579
rect 1196 3575 1199 3579
rect 1203 3575 1207 3579
rect 111 3568 115 3572
rect 491 3567 495 3571
rect 635 3567 639 3571
rect 779 3567 783 3571
rect 923 3567 927 3571
rect 1067 3567 1071 3571
rect 1211 3567 1215 3571
rect 1935 3568 1939 3572
rect 111 3551 115 3555
rect 519 3552 523 3556
rect 663 3552 667 3556
rect 807 3552 811 3556
rect 951 3552 955 3556
rect 1095 3552 1099 3556
rect 1239 3552 1243 3556
rect 1935 3551 1939 3555
rect 1975 3549 1979 3553
rect 2239 3548 2243 3552
rect 2375 3548 2379 3552
rect 2511 3548 2515 3552
rect 2647 3548 2651 3552
rect 2783 3548 2787 3552
rect 2919 3548 2923 3552
rect 3055 3548 3059 3552
rect 3191 3548 3195 3552
rect 3327 3548 3331 3552
rect 3463 3548 3467 3552
rect 3799 3549 3803 3553
rect 1975 3532 1979 3536
rect 2211 3533 2215 3537
rect 2347 3533 2351 3537
rect 2483 3533 2487 3537
rect 2619 3533 2623 3537
rect 2755 3533 2759 3537
rect 2891 3533 2895 3537
rect 3027 3533 3031 3537
rect 3163 3533 3167 3537
rect 3299 3533 3303 3537
rect 3435 3533 3439 3537
rect 3799 3532 3803 3536
rect 2363 3523 2367 3527
rect 2499 3523 2503 3527
rect 2635 3523 2639 3527
rect 2771 3523 2775 3527
rect 2803 3523 2807 3527
rect 2955 3523 2959 3527
rect 3171 3523 3175 3527
rect 3451 3523 3455 3527
rect 3251 3515 3255 3519
rect 2599 3507 2603 3511
rect 3839 3497 3843 3501
rect 5407 3496 5411 3500
rect 2363 3491 2367 3495
rect 2499 3491 2503 3495
rect 2635 3491 2639 3495
rect 2771 3491 2775 3495
rect 3171 3491 3175 3495
rect 3251 3491 3255 3495
rect 3387 3491 3391 3495
rect 5543 3496 5547 3500
rect 5663 3497 5667 3501
rect 3451 3491 3455 3495
rect 3839 3480 3843 3484
rect 5379 3481 5383 3485
rect 5515 3481 5519 3485
rect 5663 3480 5667 3484
rect 111 3473 115 3477
rect 431 3472 435 3476
rect 567 3472 571 3476
rect 703 3472 707 3476
rect 839 3472 843 3476
rect 975 3472 979 3476
rect 1935 3473 1939 3477
rect 5531 3471 5535 3475
rect 5603 3471 5607 3475
rect 111 3456 115 3460
rect 403 3457 407 3461
rect 539 3457 543 3461
rect 675 3457 679 3461
rect 811 3457 815 3461
rect 947 3457 951 3461
rect 1935 3456 1939 3460
rect 619 3447 623 3451
rect 691 3447 695 3451
rect 819 3447 823 3451
rect 963 3447 967 3451
rect 1011 3447 1015 3451
rect 2319 3439 2323 3443
rect 2327 3439 2331 3443
rect 2475 3439 2479 3443
rect 2803 3435 2807 3439
rect 2819 3439 2823 3443
rect 3187 3435 3191 3439
rect 3227 3439 3231 3443
rect 3639 3439 3643 3443
rect 5551 3455 5555 3459
rect 3739 3435 3743 3439
rect 5531 3439 5535 3443
rect 447 3415 451 3419
rect 619 3415 623 3419
rect 691 3415 695 3419
rect 899 3415 903 3419
rect 963 3415 967 3419
rect 2319 3411 2323 3415
rect 2327 3403 2331 3407
rect 2475 3403 2476 3407
rect 2476 3403 2479 3407
rect 2819 3403 2823 3407
rect 3187 3411 3191 3415
rect 3031 3403 3032 3407
rect 3032 3403 3035 3407
rect 3227 3403 3228 3407
rect 3228 3403 3231 3407
rect 3387 3403 3391 3407
rect 3639 3403 3643 3407
rect 1975 3396 1979 3400
rect 2171 3395 2175 3399
rect 2347 3395 2351 3399
rect 2531 3395 2535 3399
rect 2715 3395 2719 3399
rect 2907 3395 2911 3399
rect 3099 3395 3103 3399
rect 3291 3395 3295 3399
rect 3483 3395 3487 3399
rect 3651 3395 3655 3399
rect 3799 3396 3803 3400
rect 1975 3379 1979 3383
rect 2199 3380 2203 3384
rect 2375 3380 2379 3384
rect 2559 3380 2563 3384
rect 2743 3380 2747 3384
rect 2935 3380 2939 3384
rect 3127 3380 3131 3384
rect 3319 3380 3323 3384
rect 3511 3380 3515 3384
rect 3679 3380 3683 3384
rect 3799 3379 3803 3383
rect 4227 3383 4231 3387
rect 4295 3375 4299 3379
rect 4675 3379 4679 3383
rect 4991 3383 4995 3387
rect 5415 3383 5419 3387
rect 5443 3383 5447 3387
rect 563 3359 567 3363
rect 683 3355 687 3359
rect 819 3355 823 3359
rect 4675 3355 4679 3359
rect 3739 3347 3743 3351
rect 4295 3347 4299 3351
rect 4803 3347 4807 3351
rect 4991 3347 4995 3351
rect 5415 3347 5419 3351
rect 3839 3340 3843 3344
rect 3859 3339 3863 3343
rect 4099 3339 4103 3343
rect 4347 3339 4351 3343
rect 4587 3339 4591 3343
rect 4811 3339 4815 3343
rect 5027 3339 5031 3343
rect 5235 3339 5239 3343
rect 5451 3339 5455 3343
rect 5663 3340 5667 3344
rect 683 3331 687 3335
rect 447 3323 448 3327
rect 448 3323 451 3327
rect 739 3323 743 3327
rect 3839 3323 3843 3327
rect 3887 3324 3891 3328
rect 4127 3324 4131 3328
rect 4375 3324 4379 3328
rect 4615 3324 4619 3328
rect 4839 3324 4843 3328
rect 5055 3324 5059 3328
rect 5263 3324 5267 3328
rect 5479 3324 5483 3328
rect 5663 3323 5667 3327
rect 111 3316 115 3320
rect 323 3315 327 3319
rect 459 3315 463 3319
rect 595 3315 599 3319
rect 731 3315 735 3319
rect 867 3315 871 3319
rect 1935 3316 1939 3320
rect 111 3299 115 3303
rect 351 3300 355 3304
rect 487 3300 491 3304
rect 623 3300 627 3304
rect 759 3300 763 3304
rect 895 3300 899 3304
rect 1935 3299 1939 3303
rect 1975 3297 1979 3301
rect 2151 3296 2155 3300
rect 2399 3296 2403 3300
rect 2687 3296 2691 3300
rect 3015 3296 3019 3300
rect 3359 3296 3363 3300
rect 3679 3296 3683 3300
rect 3799 3297 3803 3301
rect 1975 3280 1979 3284
rect 2123 3281 2127 3285
rect 2371 3281 2375 3285
rect 2659 3281 2663 3285
rect 2987 3281 2991 3285
rect 3331 3281 3335 3285
rect 3651 3281 3655 3285
rect 3799 3280 3803 3284
rect 2387 3271 2391 3275
rect 2675 3271 2679 3275
rect 2683 3271 2687 3275
rect 3183 3271 3187 3275
rect 3779 3271 3780 3275
rect 3780 3271 3783 3275
rect 3839 3265 3843 3269
rect 3887 3264 3891 3268
rect 4127 3264 4131 3268
rect 4375 3264 4379 3268
rect 4607 3264 4611 3268
rect 4815 3264 4819 3268
rect 5015 3264 5019 3268
rect 5199 3264 5203 3268
rect 5383 3264 5387 3268
rect 5543 3264 5547 3268
rect 5663 3265 5667 3269
rect 3839 3248 3843 3252
rect 3859 3249 3863 3253
rect 4099 3249 4103 3253
rect 4347 3249 4351 3253
rect 4579 3249 4583 3253
rect 4787 3249 4791 3253
rect 4987 3249 4991 3253
rect 5171 3249 5175 3253
rect 5355 3249 5359 3253
rect 5515 3249 5519 3253
rect 5663 3248 5667 3252
rect 2291 3239 2295 3243
rect 2387 3239 2391 3243
rect 2675 3239 2679 3243
rect 3031 3239 3035 3243
rect 3183 3239 3187 3243
rect 3739 3239 3743 3243
rect 4115 3239 4119 3243
rect 4227 3239 4228 3243
rect 4228 3239 4231 3243
rect 4595 3239 4599 3243
rect 4759 3239 4763 3243
rect 5003 3239 5007 3243
rect 111 3233 115 3237
rect 159 3232 163 3236
rect 335 3232 339 3236
rect 543 3232 547 3236
rect 751 3232 755 3236
rect 959 3232 963 3236
rect 1935 3233 1939 3237
rect 4435 3231 4439 3235
rect 5371 3239 5375 3243
rect 5443 3239 5447 3243
rect 5619 3239 5623 3243
rect 111 3216 115 3220
rect 131 3217 135 3221
rect 307 3217 311 3221
rect 515 3217 519 3221
rect 723 3217 727 3221
rect 931 3217 935 3221
rect 1935 3216 1939 3220
rect 323 3207 327 3211
rect 531 3207 535 3211
rect 563 3207 567 3211
rect 947 3207 951 3211
rect 1059 3207 1060 3211
rect 1060 3207 1063 3211
rect 3779 3207 3783 3211
rect 4115 3207 4119 3211
rect 4435 3207 4439 3211
rect 4595 3207 4599 3211
rect 4803 3207 4807 3211
rect 5003 3207 5007 3211
rect 5363 3207 5367 3211
rect 5371 3207 5375 3211
rect 5603 3207 5607 3211
rect 1915 3191 1919 3195
rect 2123 3191 2127 3195
rect 2275 3191 2279 3195
rect 2683 3199 2687 3203
rect 2683 3191 2687 3195
rect 3415 3191 3419 3195
rect 3571 3191 3575 3195
rect 3383 3183 3387 3187
rect 227 3175 231 3179
rect 323 3175 327 3179
rect 531 3175 535 3179
rect 739 3175 743 3179
rect 947 3175 951 3179
rect 2123 3155 2124 3159
rect 2124 3155 2127 3159
rect 2275 3155 2276 3159
rect 2276 3155 2279 3159
rect 2291 3155 2295 3159
rect 2683 3155 2684 3159
rect 2684 3155 2687 3159
rect 2915 3155 2919 3159
rect 3023 3155 3027 3159
rect 3415 3155 3419 3159
rect 3571 3155 3572 3159
rect 3572 3155 3575 3159
rect 3739 3155 3743 3159
rect 1975 3148 1979 3152
rect 1995 3147 1999 3151
rect 2147 3147 2151 3151
rect 2347 3147 2351 3151
rect 2555 3147 2559 3151
rect 2771 3147 2775 3151
rect 2987 3147 2991 3151
rect 3211 3147 3215 3151
rect 3443 3147 3447 3151
rect 3651 3147 3655 3151
rect 3799 3148 3803 3152
rect 4555 3139 4559 3143
rect 4759 3143 4763 3147
rect 4987 3143 4991 3147
rect 5203 3143 5207 3147
rect 5619 3143 5623 3147
rect 1975 3131 1979 3135
rect 2023 3132 2027 3136
rect 2175 3132 2179 3136
rect 2375 3132 2379 3136
rect 2583 3132 2587 3136
rect 2799 3132 2803 3136
rect 3015 3132 3019 3136
rect 3239 3132 3243 3136
rect 3471 3132 3475 3136
rect 3679 3132 3683 3136
rect 3799 3131 3803 3135
rect 5431 3127 5435 3131
rect 331 3111 335 3115
rect 823 3111 827 3115
rect 1051 3111 1055 3115
rect 1059 3111 1063 3115
rect 1451 3111 1455 3115
rect 1475 3111 1479 3115
rect 1707 3111 1711 3115
rect 4555 3115 4559 3119
rect 4659 3107 4663 3111
rect 4987 3107 4988 3111
rect 4988 3107 4991 3111
rect 5203 3107 5204 3111
rect 5204 3107 5207 3111
rect 5431 3107 5432 3111
rect 5432 3107 5435 3111
rect 5619 3107 5623 3111
rect 3839 3100 3843 3104
rect 4467 3099 4471 3103
rect 4651 3099 4655 3103
rect 4859 3099 4863 3103
rect 5075 3099 5079 3103
rect 5307 3099 5311 3103
rect 5515 3099 5519 3103
rect 5663 3100 5667 3104
rect 3839 3083 3843 3087
rect 4495 3084 4499 3088
rect 4679 3084 4683 3088
rect 4887 3084 4891 3088
rect 5103 3084 5107 3088
rect 5335 3084 5339 3088
rect 5543 3084 5547 3088
rect 5663 3083 5667 3087
rect 227 3075 231 3079
rect 683 3075 687 3079
rect 823 3075 827 3079
rect 1051 3075 1055 3079
rect 1475 3075 1476 3079
rect 1476 3075 1479 3079
rect 1707 3075 1708 3079
rect 1708 3075 1711 3079
rect 1915 3075 1916 3079
rect 1916 3075 1919 3079
rect 1975 3073 1979 3077
rect 2647 3072 2651 3076
rect 111 3068 115 3072
rect 131 3067 135 3071
rect 371 3067 375 3071
rect 627 3067 631 3071
rect 875 3067 879 3071
rect 1115 3067 1119 3071
rect 1347 3067 1351 3071
rect 1579 3067 1583 3071
rect 1787 3067 1791 3071
rect 1935 3068 1939 3072
rect 2783 3072 2787 3076
rect 2927 3072 2931 3076
rect 3079 3072 3083 3076
rect 3239 3072 3243 3076
rect 3399 3072 3403 3076
rect 3567 3072 3571 3076
rect 3799 3073 3803 3077
rect 111 3051 115 3055
rect 159 3052 163 3056
rect 399 3052 403 3056
rect 655 3052 659 3056
rect 903 3052 907 3056
rect 1143 3052 1147 3056
rect 1375 3052 1379 3056
rect 1607 3052 1611 3056
rect 1975 3056 1979 3060
rect 2619 3057 2623 3061
rect 2755 3057 2759 3061
rect 2899 3057 2903 3061
rect 3051 3057 3055 3061
rect 3211 3057 3215 3061
rect 3371 3057 3375 3061
rect 3539 3057 3543 3061
rect 3799 3056 3803 3060
rect 1815 3052 1819 3056
rect 1935 3051 1939 3055
rect 2771 3047 2775 3051
rect 2891 3047 2895 3051
rect 3067 3047 3071 3051
rect 3227 3047 3231 3051
rect 3383 3047 3387 3051
rect 3527 3047 3531 3051
rect 4359 3039 4363 3043
rect 5263 3039 5267 3043
rect 3023 3031 3027 3035
rect 3839 3025 3843 3029
rect 4255 3024 4259 3028
rect 4455 3024 4459 3028
rect 4671 3024 4675 3028
rect 4911 3024 4915 3028
rect 5167 3024 5171 3028
rect 5423 3024 5427 3028
rect 5663 3025 5667 3029
rect 2771 3015 2775 3019
rect 2915 3015 2919 3019
rect 3067 3015 3071 3019
rect 3227 3015 3231 3019
rect 3527 3015 3531 3019
rect 3607 3015 3611 3019
rect 1451 3007 1455 3011
rect 1911 3007 1915 3011
rect 3839 3008 3843 3012
rect 4227 3009 4231 3013
rect 4427 3009 4431 3013
rect 4643 3009 4647 3013
rect 4883 3009 4887 3013
rect 5139 3009 5143 3013
rect 5395 3009 5399 3013
rect 5663 3008 5667 3012
rect 4443 2999 4447 3003
rect 4547 2999 4551 3003
rect 4899 2999 4903 3003
rect 5155 2999 5159 3003
rect 5263 2999 5264 3003
rect 5264 2999 5267 3003
rect 5363 2999 5367 3003
rect 111 2993 115 2997
rect 175 2992 179 2996
rect 407 2992 411 2996
rect 623 2992 627 2996
rect 823 2992 827 2996
rect 1007 2992 1011 2996
rect 1183 2992 1187 2996
rect 1351 2992 1355 2996
rect 1511 2992 1515 2996
rect 1671 2992 1675 2996
rect 1815 2992 1819 2996
rect 1935 2993 1939 2997
rect 111 2976 115 2980
rect 147 2977 151 2981
rect 379 2977 383 2981
rect 595 2977 599 2981
rect 795 2977 799 2981
rect 979 2977 983 2981
rect 1155 2977 1159 2981
rect 1323 2977 1327 2981
rect 1483 2977 1487 2981
rect 1643 2977 1647 2981
rect 1787 2977 1791 2981
rect 1935 2976 1939 2980
rect 331 2967 335 2971
rect 339 2967 343 2971
rect 811 2967 815 2971
rect 995 2967 999 2971
rect 907 2959 911 2963
rect 1339 2967 1343 2971
rect 1499 2967 1503 2971
rect 1659 2967 1663 2971
rect 1803 2967 1807 2971
rect 1911 2967 1912 2971
rect 1912 2967 1915 2971
rect 2891 2963 2895 2967
rect 4359 2967 4363 2971
rect 4443 2967 4447 2971
rect 4659 2967 4663 2971
rect 4899 2967 4903 2971
rect 5155 2967 5159 2971
rect 5411 2967 5415 2971
rect 339 2935 343 2939
rect 467 2935 471 2939
rect 683 2935 687 2939
rect 811 2935 815 2939
rect 995 2935 999 2939
rect 1339 2935 1343 2939
rect 1499 2935 1503 2939
rect 1659 2935 1663 2939
rect 1803 2935 1807 2939
rect 3059 2931 3063 2935
rect 3607 2931 3608 2935
rect 3608 2931 3611 2935
rect 1975 2924 1979 2928
rect 2803 2923 2807 2927
rect 2939 2923 2943 2927
rect 3075 2923 3079 2927
rect 3211 2923 3215 2927
rect 3347 2923 3351 2927
rect 3483 2923 3487 2927
rect 3799 2924 3803 2928
rect 1975 2907 1979 2911
rect 2831 2908 2835 2912
rect 2967 2908 2971 2912
rect 3103 2908 3107 2912
rect 3239 2908 3243 2912
rect 3375 2908 3379 2912
rect 3511 2908 3515 2912
rect 3799 2907 3803 2911
rect 4175 2895 4179 2899
rect 4299 2891 4303 2895
rect 4547 2895 4551 2899
rect 4571 2895 4575 2899
rect 4827 2895 4831 2899
rect 5339 2891 5343 2895
rect 5619 2895 5623 2899
rect 683 2879 687 2883
rect 907 2883 911 2887
rect 915 2883 919 2887
rect 1099 2883 1103 2887
rect 1875 2879 1879 2883
rect 4299 2867 4303 2871
rect 3979 2859 3983 2863
rect 4175 2859 4179 2863
rect 4571 2859 4572 2863
rect 4572 2859 4575 2863
rect 4827 2859 4828 2863
rect 4828 2859 4831 2863
rect 5411 2859 5415 2863
rect 5619 2859 5623 2863
rect 3839 2852 3843 2856
rect 467 2847 471 2851
rect 915 2847 916 2851
rect 916 2847 919 2851
rect 1099 2847 1100 2851
rect 1100 2847 1103 2851
rect 1203 2847 1207 2851
rect 3995 2851 3999 2855
rect 4211 2851 4215 2855
rect 4443 2851 4447 2855
rect 4699 2851 4703 2855
rect 4971 2851 4975 2855
rect 5251 2851 5255 2855
rect 5515 2851 5519 2855
rect 5663 2852 5667 2856
rect 111 2840 115 2844
rect 395 2839 399 2843
rect 595 2839 599 2843
rect 787 2839 791 2843
rect 971 2839 975 2843
rect 1147 2839 1151 2843
rect 1315 2839 1319 2843
rect 1483 2839 1487 2843
rect 1643 2839 1647 2843
rect 1787 2839 1791 2843
rect 1935 2840 1939 2844
rect 3839 2835 3843 2839
rect 4023 2836 4027 2840
rect 4239 2836 4243 2840
rect 4471 2836 4475 2840
rect 4727 2836 4731 2840
rect 4999 2836 5003 2840
rect 5279 2836 5283 2840
rect 5543 2836 5547 2840
rect 5663 2835 5667 2839
rect 111 2823 115 2827
rect 423 2824 427 2828
rect 623 2824 627 2828
rect 815 2824 819 2828
rect 999 2824 1003 2828
rect 1175 2824 1179 2828
rect 1343 2824 1347 2828
rect 1511 2824 1515 2828
rect 1671 2824 1675 2828
rect 1815 2824 1819 2828
rect 1935 2823 1939 2827
rect 1975 2797 1979 2801
rect 2023 2796 2027 2800
rect 2167 2796 2171 2800
rect 2335 2796 2339 2800
rect 2495 2796 2499 2800
rect 2663 2796 2667 2800
rect 2831 2796 2835 2800
rect 2999 2796 3003 2800
rect 3167 2796 3171 2800
rect 3799 2797 3803 2801
rect 1975 2780 1979 2784
rect 1995 2781 1999 2785
rect 2139 2781 2143 2785
rect 2307 2781 2311 2785
rect 2467 2781 2471 2785
rect 2635 2781 2639 2785
rect 2803 2781 2807 2785
rect 2971 2781 2975 2785
rect 3139 2781 3143 2785
rect 3799 2780 3803 2784
rect 1875 2771 1879 2775
rect 2747 2771 2751 2775
rect 2791 2771 2795 2775
rect 3155 2771 3159 2775
rect 2891 2763 2895 2767
rect 3839 2773 3843 2777
rect 3919 2772 3923 2776
rect 4055 2772 4059 2776
rect 4191 2772 4195 2776
rect 4327 2772 4331 2776
rect 4463 2772 4467 2776
rect 5663 2773 5667 2777
rect 111 2753 115 2757
rect 655 2752 659 2756
rect 815 2752 819 2756
rect 975 2752 979 2756
rect 1143 2752 1147 2756
rect 1311 2752 1315 2756
rect 1479 2752 1483 2756
rect 1935 2753 1939 2757
rect 3839 2756 3843 2760
rect 3891 2757 3895 2761
rect 4027 2757 4031 2761
rect 4163 2757 4167 2761
rect 4299 2757 4303 2761
rect 4435 2757 4439 2761
rect 5663 2756 5667 2760
rect 4043 2747 4047 2751
rect 4179 2747 4183 2751
rect 4315 2747 4319 2751
rect 4451 2747 4455 2751
rect 111 2736 115 2740
rect 627 2737 631 2741
rect 787 2737 791 2741
rect 947 2737 951 2741
rect 1115 2737 1119 2741
rect 1283 2737 1287 2741
rect 1451 2737 1455 2741
rect 1935 2736 1939 2740
rect 2503 2739 2507 2743
rect 2791 2739 2795 2743
rect 2891 2739 2895 2743
rect 3059 2739 3063 2743
rect 3155 2739 3159 2743
rect 4219 2739 4223 2743
rect 683 2727 687 2731
rect 1299 2727 1303 2731
rect 1467 2727 1471 2731
rect 1555 2727 1559 2731
rect 3979 2715 3983 2719
rect 4043 2715 4047 2719
rect 4179 2715 4183 2719
rect 4315 2715 4319 2719
rect 4451 2715 4455 2719
rect 1031 2695 1035 2699
rect 1203 2695 1207 2699
rect 1299 2695 1303 2699
rect 1467 2695 1471 2699
rect 2603 2687 2607 2691
rect 2747 2687 2751 2691
rect 2787 2691 2791 2695
rect 2931 2691 2935 2695
rect 3075 2691 3079 2695
rect 3219 2691 3223 2695
rect 2503 2655 2504 2659
rect 2504 2655 2507 2659
rect 2787 2655 2788 2659
rect 2788 2655 2791 2659
rect 2931 2655 2932 2659
rect 2932 2655 2935 2659
rect 3075 2655 3076 2659
rect 3076 2655 3079 2659
rect 3219 2655 3220 2659
rect 3220 2655 3223 2659
rect 3271 2655 3275 2659
rect 4219 2655 4223 2659
rect 4227 2655 4231 2659
rect 4427 2655 4431 2659
rect 4643 2655 4647 2659
rect 4883 2655 4887 2659
rect 5399 2655 5403 2659
rect 5619 2655 5623 2659
rect 859 2643 863 2647
rect 1403 2643 1407 2647
rect 1555 2647 1559 2651
rect 1975 2648 1979 2652
rect 2379 2647 2383 2651
rect 2515 2647 2519 2651
rect 2659 2647 2663 2651
rect 2803 2647 2807 2651
rect 2947 2647 2951 2651
rect 3091 2647 3095 2651
rect 3235 2647 3239 2651
rect 3799 2648 3803 2652
rect 1975 2631 1979 2635
rect 2407 2632 2411 2636
rect 2543 2632 2547 2636
rect 2687 2632 2691 2636
rect 2831 2632 2835 2636
rect 2975 2632 2979 2636
rect 3119 2632 3123 2636
rect 3263 2632 3267 2636
rect 3799 2631 3803 2635
rect 859 2619 863 2623
rect 1031 2611 1032 2615
rect 1032 2611 1035 2615
rect 4227 2619 4228 2623
rect 4228 2619 4231 2623
rect 4427 2619 4428 2623
rect 4428 2619 4431 2623
rect 4643 2619 4644 2623
rect 4644 2619 4647 2623
rect 4883 2619 4884 2623
rect 4884 2619 4887 2623
rect 4999 2619 5003 2623
rect 5339 2619 5343 2623
rect 5619 2619 5623 2623
rect 1843 2611 1847 2615
rect 3839 2612 3843 2616
rect 4099 2611 4103 2615
rect 4299 2611 4303 2615
rect 4515 2611 4519 2615
rect 4755 2611 4759 2615
rect 5011 2611 5015 2615
rect 5275 2611 5279 2615
rect 5515 2611 5519 2615
rect 5663 2612 5667 2616
rect 111 2604 115 2608
rect 771 2603 775 2607
rect 907 2603 911 2607
rect 1043 2603 1047 2607
rect 1179 2603 1183 2607
rect 1315 2603 1319 2607
rect 1451 2603 1455 2607
rect 1587 2603 1591 2607
rect 1723 2603 1727 2607
rect 1935 2604 1939 2608
rect 3839 2595 3843 2599
rect 4127 2596 4131 2600
rect 4327 2596 4331 2600
rect 4543 2596 4547 2600
rect 4783 2596 4787 2600
rect 5039 2596 5043 2600
rect 5303 2596 5307 2600
rect 5543 2596 5547 2600
rect 5663 2595 5667 2599
rect 111 2587 115 2591
rect 799 2588 803 2592
rect 935 2588 939 2592
rect 1071 2588 1075 2592
rect 1207 2588 1211 2592
rect 1343 2588 1347 2592
rect 1479 2588 1483 2592
rect 1615 2588 1619 2592
rect 1751 2588 1755 2592
rect 1935 2587 1939 2591
rect 1975 2569 1979 2573
rect 2511 2568 2515 2572
rect 2647 2568 2651 2572
rect 2783 2568 2787 2572
rect 2919 2568 2923 2572
rect 3055 2568 3059 2572
rect 3191 2568 3195 2572
rect 3327 2568 3331 2572
rect 3463 2568 3467 2572
rect 3799 2569 3803 2573
rect 1975 2552 1979 2556
rect 2483 2553 2487 2557
rect 2619 2553 2623 2557
rect 2755 2553 2759 2557
rect 2891 2553 2895 2557
rect 3027 2553 3031 2557
rect 3163 2553 3167 2557
rect 3299 2553 3303 2557
rect 3435 2553 3439 2557
rect 3799 2552 3803 2556
rect 2603 2543 2607 2547
rect 3043 2543 3047 2547
rect 3179 2543 3183 2547
rect 3315 2543 3319 2547
rect 3451 2543 3455 2547
rect 2979 2535 2983 2539
rect 3271 2535 3275 2539
rect 3015 2527 3019 2531
rect 3839 2533 3843 2537
rect 4495 2532 4499 2536
rect 4631 2532 4635 2536
rect 4767 2532 4771 2536
rect 4903 2532 4907 2536
rect 5039 2532 5043 2536
rect 5663 2533 5667 2537
rect 111 2513 115 2517
rect 551 2512 555 2516
rect 687 2512 691 2516
rect 831 2512 835 2516
rect 983 2512 987 2516
rect 1135 2512 1139 2516
rect 1295 2512 1299 2516
rect 1455 2512 1459 2516
rect 1615 2512 1619 2516
rect 1783 2512 1787 2516
rect 1935 2513 1939 2517
rect 3839 2516 3843 2520
rect 4467 2517 4471 2521
rect 4603 2517 4607 2521
rect 4739 2517 4743 2521
rect 4875 2517 4879 2521
rect 5011 2517 5015 2521
rect 5663 2516 5667 2520
rect 2839 2511 2843 2515
rect 2979 2511 2983 2515
rect 3043 2511 3047 2515
rect 3179 2511 3183 2515
rect 3315 2511 3319 2515
rect 3451 2511 3455 2515
rect 4619 2507 4623 2511
rect 4755 2507 4759 2511
rect 4891 2507 4895 2511
rect 5027 2507 5031 2511
rect 111 2496 115 2500
rect 523 2497 527 2501
rect 659 2497 663 2501
rect 803 2497 807 2501
rect 955 2497 959 2501
rect 1107 2497 1111 2501
rect 1267 2497 1271 2501
rect 1427 2497 1431 2501
rect 1587 2497 1591 2501
rect 1755 2497 1759 2501
rect 1935 2496 1939 2500
rect 4819 2499 4823 2503
rect 675 2487 679 2491
rect 819 2487 823 2491
rect 971 2487 975 2491
rect 1123 2487 1127 2491
rect 1283 2487 1287 2491
rect 1403 2487 1407 2491
rect 1411 2487 1415 2491
rect 1743 2487 1747 2491
rect 4999 2491 5003 2495
rect 4619 2475 4623 2479
rect 4755 2475 4759 2479
rect 4891 2475 4895 2479
rect 5027 2475 5031 2479
rect 667 2455 671 2459
rect 675 2455 679 2459
rect 819 2455 823 2459
rect 971 2455 975 2459
rect 1123 2455 1127 2459
rect 1283 2455 1287 2459
rect 1743 2455 1747 2459
rect 1843 2455 1847 2459
rect 2299 2447 2303 2451
rect 2435 2447 2439 2451
rect 2643 2447 2647 2451
rect 3015 2447 3019 2451
rect 3035 2447 3039 2451
rect 3227 2447 3231 2451
rect 3411 2447 3415 2451
rect 3595 2447 3599 2451
rect 2435 2411 2436 2415
rect 2436 2411 2439 2415
rect 2643 2411 2644 2415
rect 2644 2411 2647 2415
rect 2839 2411 2840 2415
rect 2840 2411 2843 2415
rect 3035 2411 3036 2415
rect 3036 2411 3039 2415
rect 3227 2411 3228 2415
rect 3228 2411 3231 2415
rect 3411 2411 3412 2415
rect 3412 2411 3415 2415
rect 3595 2411 3596 2415
rect 3596 2411 3599 2415
rect 3739 2411 3743 2415
rect 4819 2411 4823 2415
rect 4827 2411 4831 2415
rect 1975 2404 1979 2408
rect 2307 2403 2311 2407
rect 2515 2403 2519 2407
rect 2715 2403 2719 2407
rect 2907 2403 2911 2407
rect 3099 2403 3103 2407
rect 3283 2403 3287 2407
rect 3467 2403 3471 2407
rect 3651 2403 3655 2407
rect 3799 2404 3803 2408
rect 5467 2407 5471 2411
rect 5619 2411 5623 2415
rect 219 2391 223 2395
rect 307 2395 311 2399
rect 467 2395 471 2399
rect 691 2395 695 2399
rect 931 2395 935 2399
rect 1411 2395 1415 2399
rect 1439 2395 1443 2399
rect 1675 2395 1679 2399
rect 1975 2387 1979 2391
rect 2335 2388 2339 2392
rect 2543 2388 2547 2392
rect 2743 2388 2747 2392
rect 2935 2388 2939 2392
rect 3127 2388 3131 2392
rect 3311 2388 3315 2392
rect 3495 2388 3499 2392
rect 3679 2388 3683 2392
rect 3799 2387 3803 2391
rect 5467 2383 5471 2387
rect 5551 2383 5555 2387
rect 4827 2375 4828 2379
rect 4828 2375 4831 2379
rect 5371 2375 5372 2379
rect 5372 2375 5375 2379
rect 5399 2375 5403 2379
rect 5619 2375 5623 2379
rect 667 2367 671 2371
rect 307 2359 311 2363
rect 467 2359 468 2363
rect 468 2359 471 2363
rect 691 2359 692 2363
rect 692 2359 695 2363
rect 931 2359 932 2363
rect 932 2359 935 2363
rect 3839 2368 3843 2372
rect 4699 2367 4703 2371
rect 4835 2367 4839 2371
rect 4971 2367 4975 2371
rect 5107 2367 5111 2371
rect 5243 2367 5247 2371
rect 5379 2367 5383 2371
rect 5515 2367 5519 2371
rect 5663 2368 5667 2372
rect 1439 2359 1443 2363
rect 1675 2359 1676 2363
rect 1676 2359 1679 2363
rect 1875 2359 1879 2363
rect 111 2352 115 2356
rect 131 2351 135 2355
rect 339 2351 343 2355
rect 563 2351 567 2355
rect 803 2351 807 2355
rect 1043 2351 1047 2355
rect 1291 2351 1295 2355
rect 1547 2351 1551 2355
rect 1787 2351 1791 2355
rect 1935 2352 1939 2356
rect 3839 2351 3843 2355
rect 4727 2352 4731 2356
rect 4863 2352 4867 2356
rect 4999 2352 5003 2356
rect 5135 2352 5139 2356
rect 5271 2352 5275 2356
rect 5407 2352 5411 2356
rect 5543 2352 5547 2356
rect 5663 2351 5667 2355
rect 111 2335 115 2339
rect 159 2336 163 2340
rect 367 2336 371 2340
rect 591 2336 595 2340
rect 831 2336 835 2340
rect 1071 2336 1075 2340
rect 1319 2336 1323 2340
rect 1575 2336 1579 2340
rect 1815 2336 1819 2340
rect 1935 2335 1939 2339
rect 1975 2321 1979 2325
rect 2223 2320 2227 2324
rect 2503 2320 2507 2324
rect 2767 2320 2771 2324
rect 3007 2320 3011 2324
rect 3239 2320 3243 2324
rect 3471 2320 3475 2324
rect 3679 2320 3683 2324
rect 3799 2321 3803 2325
rect 1975 2304 1979 2308
rect 2195 2305 2199 2309
rect 2475 2305 2479 2309
rect 2739 2305 2743 2309
rect 2979 2305 2983 2309
rect 3211 2305 3215 2309
rect 3443 2305 3447 2309
rect 3651 2305 3655 2309
rect 3799 2304 3803 2308
rect 2299 2295 2303 2299
rect 2335 2295 2339 2299
rect 2995 2295 2999 2299
rect 3227 2295 3231 2299
rect 3459 2295 3463 2299
rect 3667 2295 3671 2299
rect 3755 2295 3759 2299
rect 1247 2287 1251 2291
rect 2827 2287 2831 2291
rect 3739 2287 3743 2291
rect 3839 2281 3843 2285
rect 3887 2280 3891 2284
rect 4183 2280 4187 2284
rect 4495 2280 4499 2284
rect 4791 2280 4795 2284
rect 5087 2280 5091 2284
rect 5383 2280 5387 2284
rect 5663 2281 5667 2285
rect 111 2273 115 2277
rect 159 2272 163 2276
rect 319 2272 323 2276
rect 551 2272 555 2276
rect 831 2272 835 2276
rect 1151 2272 1155 2276
rect 1495 2272 1499 2276
rect 1815 2272 1819 2276
rect 1935 2273 1939 2277
rect 2335 2263 2339 2267
rect 2563 2263 2567 2267
rect 2827 2263 2831 2267
rect 2995 2263 2999 2267
rect 3227 2263 3231 2267
rect 3459 2263 3463 2267
rect 3667 2263 3671 2267
rect 3839 2264 3843 2268
rect 3859 2265 3863 2269
rect 4155 2265 4159 2269
rect 4467 2265 4471 2269
rect 4763 2265 4767 2269
rect 5059 2265 5063 2269
rect 5355 2265 5359 2269
rect 5663 2264 5667 2268
rect 111 2256 115 2260
rect 131 2257 135 2261
rect 291 2257 295 2261
rect 523 2257 527 2261
rect 803 2257 807 2261
rect 1123 2257 1127 2261
rect 1467 2257 1471 2261
rect 1787 2257 1791 2261
rect 1935 2256 1939 2260
rect 3963 2255 3967 2259
rect 4483 2255 4487 2259
rect 4627 2255 4631 2259
rect 307 2247 311 2251
rect 539 2247 543 2251
rect 819 2247 823 2251
rect 1247 2247 1248 2251
rect 1248 2247 1251 2251
rect 1267 2247 1271 2251
rect 1915 2247 1916 2251
rect 1916 2247 1919 2251
rect 4243 2247 4247 2251
rect 5003 2255 5007 2259
rect 5279 2255 5283 2259
rect 219 2239 223 2243
rect 3779 2223 3783 2227
rect 4243 2223 4247 2227
rect 4483 2223 4487 2227
rect 5003 2223 5007 2227
rect 5279 2223 5283 2227
rect 5371 2223 5375 2227
rect 307 2215 311 2219
rect 539 2215 543 2219
rect 819 2215 823 2219
rect 1267 2215 1271 2219
rect 1275 2215 1279 2219
rect 1875 2215 1879 2219
rect 1915 2215 1919 2219
rect 2123 2215 2127 2219
rect 2515 2215 2519 2219
rect 2795 2215 2799 2219
rect 3115 2215 3119 2219
rect 3755 2215 3759 2219
rect 2563 2187 2567 2191
rect 2123 2179 2124 2183
rect 2124 2179 2127 2183
rect 2515 2179 2516 2183
rect 2516 2179 2519 2183
rect 2795 2179 2796 2183
rect 2796 2179 2799 2183
rect 3115 2179 3116 2183
rect 3116 2179 3119 2183
rect 3779 2179 3780 2183
rect 3780 2179 3783 2183
rect 1975 2172 1979 2176
rect 1995 2171 1999 2175
rect 2155 2171 2159 2175
rect 2387 2171 2391 2175
rect 2667 2171 2671 2175
rect 2987 2171 2991 2175
rect 3331 2171 3335 2175
rect 3651 2171 3655 2175
rect 3799 2172 3803 2176
rect 3963 2171 3967 2175
rect 3987 2171 3991 2175
rect 4627 2167 4631 2171
rect 4667 2171 4671 2175
rect 4827 2171 4831 2175
rect 5019 2171 5023 2175
rect 5619 2171 5623 2175
rect 1975 2155 1979 2159
rect 2023 2156 2027 2160
rect 2183 2156 2187 2160
rect 2415 2156 2419 2160
rect 2695 2156 2699 2160
rect 3015 2156 3019 2160
rect 3359 2156 3363 2160
rect 3679 2156 3683 2160
rect 3799 2155 3803 2159
rect 419 2143 423 2147
rect 1003 2139 1007 2143
rect 1019 2143 1023 2147
rect 1615 2143 1619 2147
rect 1627 2143 1631 2147
rect 3987 2135 3988 2139
rect 3988 2135 3991 2139
rect 4491 2135 4495 2139
rect 4667 2135 4668 2139
rect 4668 2135 4671 2139
rect 4827 2135 4828 2139
rect 4828 2135 4831 2139
rect 5019 2135 5020 2139
rect 5020 2135 5023 2139
rect 5355 2135 5359 2139
rect 5619 2135 5623 2139
rect 815 2127 819 2131
rect 3839 2128 3843 2132
rect 3859 2127 3863 2131
rect 3995 2127 3999 2131
rect 4131 2127 4135 2131
rect 4267 2127 4271 2131
rect 4403 2127 4407 2131
rect 4539 2127 4543 2131
rect 4699 2127 4703 2131
rect 4891 2127 4895 2131
rect 5099 2127 5103 2131
rect 5315 2127 5319 2131
rect 5515 2127 5519 2131
rect 5663 2128 5667 2132
rect 419 2107 420 2111
rect 420 2107 423 2111
rect 1019 2115 1023 2119
rect 815 2107 816 2111
rect 816 2107 819 2111
rect 1275 2107 1276 2111
rect 1276 2107 1279 2111
rect 1459 2107 1463 2111
rect 1615 2107 1619 2111
rect 3839 2111 3843 2115
rect 3887 2112 3891 2116
rect 4023 2112 4027 2116
rect 4159 2112 4163 2116
rect 4295 2112 4299 2116
rect 4431 2112 4435 2116
rect 4567 2112 4571 2116
rect 4727 2112 4731 2116
rect 4919 2112 4923 2116
rect 5127 2112 5131 2116
rect 5343 2112 5347 2116
rect 5543 2112 5547 2116
rect 5663 2111 5667 2115
rect 111 2100 115 2104
rect 291 2099 295 2103
rect 483 2099 487 2103
rect 691 2099 695 2103
rect 915 2099 919 2103
rect 1147 2099 1151 2103
rect 1387 2099 1391 2103
rect 1635 2099 1639 2103
rect 1935 2100 1939 2104
rect 111 2083 115 2087
rect 319 2084 323 2088
rect 511 2084 515 2088
rect 719 2084 723 2088
rect 943 2084 947 2088
rect 1175 2084 1179 2088
rect 1415 2084 1419 2088
rect 1663 2084 1667 2088
rect 1935 2083 1939 2087
rect 3839 2033 3843 2037
rect 3887 2032 3891 2036
rect 4023 2032 4027 2036
rect 4159 2032 4163 2036
rect 4295 2032 4299 2036
rect 4431 2032 4435 2036
rect 4567 2032 4571 2036
rect 4719 2032 4723 2036
rect 4895 2032 4899 2036
rect 5087 2032 5091 2036
rect 5279 2032 5283 2036
rect 5479 2032 5483 2036
rect 5663 2033 5667 2037
rect 111 2021 115 2025
rect 263 2020 267 2024
rect 399 2020 403 2024
rect 535 2020 539 2024
rect 679 2020 683 2024
rect 823 2020 827 2024
rect 967 2020 971 2024
rect 1111 2020 1115 2024
rect 1255 2020 1259 2024
rect 1399 2020 1403 2024
rect 1543 2020 1547 2024
rect 1679 2020 1683 2024
rect 1815 2020 1819 2024
rect 1935 2021 1939 2025
rect 3839 2016 3843 2020
rect 3859 2017 3863 2021
rect 3995 2017 3999 2021
rect 4131 2017 4135 2021
rect 4267 2017 4271 2021
rect 4403 2017 4407 2021
rect 4539 2017 4543 2021
rect 4691 2017 4695 2021
rect 4867 2017 4871 2021
rect 5059 2017 5063 2021
rect 5251 2017 5255 2021
rect 5451 2017 5455 2021
rect 5663 2016 5667 2020
rect 111 2004 115 2008
rect 235 2005 239 2009
rect 371 2005 375 2009
rect 507 2005 511 2009
rect 651 2005 655 2009
rect 795 2005 799 2009
rect 939 2005 943 2009
rect 1083 2005 1087 2009
rect 1227 2005 1231 2009
rect 1371 2005 1375 2009
rect 1515 2005 1519 2009
rect 1651 2005 1655 2009
rect 1787 2005 1791 2009
rect 1935 2004 1939 2008
rect 3963 2007 3967 2011
rect 4683 2007 4687 2011
rect 4835 2007 4839 2011
rect 5551 2007 5555 2011
rect 387 1995 391 1999
rect 523 1995 527 1999
rect 667 1995 671 1999
rect 811 1995 815 1999
rect 955 1995 959 1999
rect 1003 1995 1007 1999
rect 931 1987 935 1991
rect 1627 1995 1631 1999
rect 1803 1995 1807 1999
rect 1603 1987 1607 1991
rect 4491 1975 4495 1979
rect 4683 1975 4687 1979
rect 4835 1975 4839 1979
rect 5355 1975 5359 1979
rect 5503 1975 5507 1979
rect 387 1963 391 1967
rect 523 1963 527 1967
rect 667 1963 671 1967
rect 811 1963 815 1967
rect 955 1963 959 1967
rect 1459 1963 1463 1967
rect 1603 1963 1607 1967
rect 1739 1963 1743 1967
rect 1803 1963 1807 1967
rect 751 1947 755 1951
rect 3963 1927 3967 1931
rect 4667 1939 4671 1943
rect 5327 1939 5331 1943
rect 4171 1927 4175 1931
rect 4411 1927 4415 1931
rect 4691 1927 4695 1931
rect 5003 1927 5007 1931
rect 5619 1927 5623 1931
rect 323 1899 327 1903
rect 363 1903 367 1907
rect 563 1903 567 1907
rect 931 1903 935 1907
rect 939 1903 943 1907
rect 1115 1903 1119 1907
rect 1411 1899 1415 1903
rect 1451 1903 1455 1907
rect 1611 1903 1615 1907
rect 2003 1903 2007 1907
rect 1975 1897 1979 1901
rect 3135 1896 3139 1900
rect 3271 1896 3275 1900
rect 3407 1896 3411 1900
rect 3543 1896 3547 1900
rect 3679 1896 3683 1900
rect 3799 1897 3803 1901
rect 3823 1891 3827 1895
rect 4171 1891 4172 1895
rect 4172 1891 4175 1895
rect 4411 1891 4412 1895
rect 4412 1891 4415 1895
rect 4467 1891 4471 1895
rect 4667 1891 4671 1895
rect 4691 1891 4692 1895
rect 4692 1891 4695 1895
rect 5003 1891 5004 1895
rect 5004 1891 5007 1895
rect 5327 1891 5328 1895
rect 5328 1891 5331 1895
rect 5619 1891 5623 1895
rect 1975 1880 1979 1884
rect 3107 1881 3111 1885
rect 3243 1881 3247 1885
rect 3379 1881 3383 1885
rect 3515 1881 3519 1885
rect 3651 1881 3655 1885
rect 3799 1880 3803 1884
rect 3839 1884 3843 1888
rect 3859 1883 3863 1887
rect 4043 1883 4047 1887
rect 4283 1883 4287 1887
rect 4563 1883 4567 1887
rect 4875 1883 4879 1887
rect 5203 1883 5207 1887
rect 5515 1883 5519 1887
rect 5663 1884 5667 1888
rect 1411 1875 1415 1879
rect 363 1867 364 1871
rect 364 1867 367 1871
rect 563 1867 564 1871
rect 564 1867 567 1871
rect 751 1867 752 1871
rect 752 1867 755 1871
rect 939 1867 940 1871
rect 940 1867 943 1871
rect 1115 1867 1116 1871
rect 1116 1867 1119 1871
rect 1379 1867 1383 1871
rect 1451 1867 1452 1871
rect 1452 1867 1455 1871
rect 1611 1867 1612 1871
rect 1612 1867 1615 1871
rect 1739 1867 1743 1871
rect 3259 1871 3263 1875
rect 3347 1871 3351 1875
rect 111 1860 115 1864
rect 235 1859 239 1863
rect 435 1859 439 1863
rect 627 1859 631 1863
rect 811 1859 815 1863
rect 987 1859 991 1863
rect 1155 1859 1159 1863
rect 1323 1859 1327 1863
rect 1483 1859 1487 1863
rect 1643 1859 1647 1863
rect 1787 1859 1791 1863
rect 1935 1860 1939 1864
rect 3195 1863 3199 1867
rect 3839 1867 3843 1871
rect 3887 1868 3891 1872
rect 4071 1868 4075 1872
rect 4311 1868 4315 1872
rect 4591 1868 4595 1872
rect 4903 1868 4907 1872
rect 5231 1868 5235 1872
rect 5543 1868 5547 1872
rect 5663 1867 5667 1871
rect 111 1843 115 1847
rect 263 1844 267 1848
rect 463 1844 467 1848
rect 655 1844 659 1848
rect 839 1844 843 1848
rect 1015 1844 1019 1848
rect 1183 1844 1187 1848
rect 1351 1844 1355 1848
rect 1511 1844 1515 1848
rect 1671 1844 1675 1848
rect 1815 1844 1819 1848
rect 1935 1843 1939 1847
rect 3195 1839 3199 1843
rect 3259 1839 3263 1843
rect 3823 1839 3827 1843
rect 3839 1809 3843 1813
rect 4407 1808 4411 1812
rect 4543 1808 4547 1812
rect 4679 1808 4683 1812
rect 4815 1808 4819 1812
rect 4951 1808 4955 1812
rect 5663 1809 5667 1813
rect 3839 1792 3843 1796
rect 4379 1793 4383 1797
rect 4515 1793 4519 1797
rect 4651 1793 4655 1797
rect 4787 1793 4791 1797
rect 4923 1793 4927 1797
rect 5663 1792 5667 1796
rect 2723 1779 2727 1783
rect 2731 1779 2735 1783
rect 3023 1779 3027 1783
rect 3179 1779 3183 1783
rect 3347 1779 3351 1783
rect 3483 1779 3487 1783
rect 4531 1783 4535 1787
rect 4667 1783 4671 1787
rect 4803 1783 4807 1787
rect 4939 1783 4943 1787
rect 4951 1783 4955 1787
rect 111 1773 115 1777
rect 223 1772 227 1776
rect 463 1772 467 1776
rect 695 1772 699 1776
rect 927 1772 931 1776
rect 1159 1772 1163 1776
rect 1391 1772 1395 1776
rect 1935 1773 1939 1777
rect 111 1756 115 1760
rect 195 1757 199 1761
rect 435 1757 439 1761
rect 667 1757 671 1761
rect 899 1757 903 1761
rect 1131 1757 1135 1761
rect 1363 1757 1367 1761
rect 1935 1756 1939 1760
rect 323 1747 324 1751
rect 324 1747 327 1751
rect 915 1747 919 1751
rect 1147 1747 1151 1751
rect 1243 1747 1247 1751
rect 755 1739 759 1743
rect 4467 1751 4471 1755
rect 4531 1751 4535 1755
rect 4667 1751 4671 1755
rect 4803 1751 4807 1755
rect 4939 1751 4943 1755
rect 2003 1743 2007 1747
rect 2723 1743 2727 1747
rect 3179 1743 3180 1747
rect 3180 1743 3183 1747
rect 3323 1743 3327 1747
rect 3483 1743 3484 1747
rect 3484 1743 3487 1747
rect 3771 1743 3775 1747
rect 1975 1736 1979 1740
rect 1995 1735 1999 1739
rect 2131 1735 2135 1739
rect 2267 1735 2271 1739
rect 2419 1735 2423 1739
rect 2579 1735 2583 1739
rect 2739 1735 2743 1739
rect 2899 1735 2903 1739
rect 3051 1735 3055 1739
rect 3203 1735 3207 1739
rect 3355 1735 3359 1739
rect 3515 1735 3519 1739
rect 3651 1735 3655 1739
rect 3799 1736 3803 1740
rect 487 1715 491 1719
rect 755 1715 759 1719
rect 915 1715 919 1719
rect 1147 1715 1151 1719
rect 1379 1715 1383 1719
rect 1975 1719 1979 1723
rect 2023 1720 2027 1724
rect 2159 1720 2163 1724
rect 2295 1720 2299 1724
rect 2447 1720 2451 1724
rect 2607 1720 2611 1724
rect 2767 1720 2771 1724
rect 2927 1720 2931 1724
rect 3079 1720 3083 1724
rect 3231 1720 3235 1724
rect 3383 1720 3387 1724
rect 3543 1720 3547 1724
rect 3679 1720 3683 1724
rect 3799 1719 3803 1723
rect 4951 1687 4955 1691
rect 5099 1687 5103 1691
rect 5331 1683 5335 1687
rect 5371 1687 5375 1691
rect 5619 1687 5623 1691
rect 219 1651 223 1655
rect 259 1655 263 1659
rect 963 1651 967 1655
rect 1243 1655 1247 1659
rect 5331 1659 5335 1663
rect 1975 1649 1979 1653
rect 2023 1648 2027 1652
rect 2167 1648 2171 1652
rect 2319 1648 2323 1652
rect 2479 1648 2483 1652
rect 2639 1648 2643 1652
rect 2791 1648 2795 1652
rect 2943 1648 2947 1652
rect 3103 1648 3107 1652
rect 3263 1648 3267 1652
rect 3423 1648 3427 1652
rect 3799 1649 3803 1653
rect 4651 1651 4655 1655
rect 5099 1651 5100 1655
rect 5100 1651 5103 1655
rect 5339 1651 5343 1655
rect 5371 1651 5372 1655
rect 5372 1651 5375 1655
rect 5503 1651 5504 1655
rect 5504 1651 5507 1655
rect 3839 1644 3843 1648
rect 4563 1643 4567 1647
rect 4699 1643 4703 1647
rect 4835 1643 4839 1647
rect 4971 1643 4975 1647
rect 5107 1643 5111 1647
rect 5243 1643 5247 1647
rect 5379 1643 5383 1647
rect 5515 1643 5519 1647
rect 5663 1644 5667 1648
rect 963 1631 967 1635
rect 259 1619 260 1623
rect 260 1619 263 1623
rect 487 1619 488 1623
rect 488 1619 491 1623
rect 571 1619 575 1623
rect 1975 1632 1979 1636
rect 1995 1633 1999 1637
rect 2139 1633 2143 1637
rect 2291 1633 2295 1637
rect 2451 1633 2455 1637
rect 2611 1633 2615 1637
rect 2763 1633 2767 1637
rect 2915 1633 2919 1637
rect 3075 1633 3079 1637
rect 3235 1633 3239 1637
rect 3395 1633 3399 1637
rect 3799 1632 3803 1636
rect 2155 1623 2159 1627
rect 2307 1623 2311 1627
rect 2467 1623 2471 1627
rect 2627 1623 2631 1627
rect 2731 1623 2735 1627
rect 2931 1623 2935 1627
rect 3091 1623 3095 1627
rect 3411 1623 3415 1627
rect 111 1612 115 1616
rect 131 1611 135 1615
rect 363 1611 367 1615
rect 619 1611 623 1615
rect 875 1611 879 1615
rect 1139 1611 1143 1615
rect 1935 1612 1939 1616
rect 2851 1615 2855 1619
rect 3839 1627 3843 1631
rect 4591 1628 4595 1632
rect 4727 1628 4731 1632
rect 4863 1628 4867 1632
rect 4999 1628 5003 1632
rect 5135 1628 5139 1632
rect 5271 1628 5275 1632
rect 5407 1628 5411 1632
rect 5543 1628 5547 1632
rect 5663 1627 5667 1631
rect 111 1595 115 1599
rect 159 1596 163 1600
rect 391 1596 395 1600
rect 647 1596 651 1600
rect 903 1596 907 1600
rect 1167 1596 1171 1600
rect 1935 1595 1939 1599
rect 2091 1591 2095 1595
rect 2155 1591 2159 1595
rect 2307 1591 2311 1595
rect 2467 1591 2471 1595
rect 2627 1591 2631 1595
rect 2851 1591 2855 1595
rect 2931 1591 2935 1595
rect 3091 1591 3095 1595
rect 3323 1591 3327 1595
rect 3411 1591 3415 1595
rect 3839 1553 3843 1557
rect 4591 1552 4595 1556
rect 4727 1552 4731 1556
rect 4863 1552 4867 1556
rect 4999 1552 5003 1556
rect 5135 1552 5139 1556
rect 5271 1552 5275 1556
rect 5407 1552 5411 1556
rect 5543 1552 5547 1556
rect 5663 1553 5667 1557
rect 3839 1536 3843 1540
rect 4563 1537 4567 1541
rect 4699 1537 4703 1541
rect 4835 1537 4839 1541
rect 4971 1537 4975 1541
rect 5107 1537 5111 1541
rect 5243 1537 5247 1541
rect 5379 1537 5383 1541
rect 5515 1537 5519 1541
rect 5663 1536 5667 1540
rect 2259 1531 2263 1535
rect 111 1525 115 1529
rect 159 1524 163 1528
rect 327 1524 331 1528
rect 511 1524 515 1528
rect 695 1524 699 1528
rect 887 1524 891 1528
rect 1079 1524 1083 1528
rect 1935 1525 1939 1529
rect 2627 1527 2631 1531
rect 2799 1515 2803 1519
rect 4715 1527 4719 1531
rect 4851 1527 4855 1531
rect 4987 1527 4991 1531
rect 5123 1527 5127 1531
rect 5259 1527 5263 1531
rect 5531 1527 5535 1531
rect 3615 1515 3619 1519
rect 111 1508 115 1512
rect 131 1509 135 1513
rect 299 1509 303 1513
rect 483 1509 487 1513
rect 667 1509 671 1513
rect 859 1509 863 1513
rect 1051 1509 1055 1513
rect 1935 1508 1939 1512
rect 219 1499 223 1503
rect 287 1499 291 1503
rect 683 1499 687 1503
rect 875 1499 879 1503
rect 1067 1499 1071 1503
rect 803 1491 807 1495
rect 2091 1495 2095 1499
rect 2627 1495 2631 1499
rect 2635 1495 2639 1499
rect 2799 1495 2800 1499
rect 2800 1495 2803 1499
rect 3615 1495 3616 1499
rect 3616 1495 3619 1499
rect 4651 1495 4655 1499
rect 4715 1495 4719 1499
rect 4851 1495 4855 1499
rect 4987 1495 4991 1499
rect 5123 1495 5127 1499
rect 5259 1495 5263 1499
rect 5339 1495 5343 1499
rect 5531 1495 5535 1499
rect 1975 1488 1979 1492
rect 1995 1487 1999 1491
rect 2131 1487 2135 1491
rect 2267 1487 2271 1491
rect 2403 1487 2407 1491
rect 2539 1487 2543 1491
rect 2675 1487 2679 1491
rect 2811 1487 2815 1491
rect 2947 1487 2951 1491
rect 3083 1487 3087 1491
rect 3219 1487 3223 1491
rect 3355 1487 3359 1491
rect 3491 1487 3495 1491
rect 3799 1488 3803 1492
rect 287 1467 291 1471
rect 387 1467 391 1471
rect 571 1467 575 1471
rect 683 1467 687 1471
rect 875 1467 879 1471
rect 1067 1467 1071 1471
rect 1975 1471 1979 1475
rect 2023 1472 2027 1476
rect 2159 1472 2163 1476
rect 2295 1472 2299 1476
rect 2431 1472 2435 1476
rect 2567 1472 2571 1476
rect 2703 1472 2707 1476
rect 2839 1472 2843 1476
rect 2975 1472 2979 1476
rect 3111 1472 3115 1476
rect 3247 1472 3251 1476
rect 3383 1472 3387 1476
rect 3519 1472 3523 1476
rect 3799 1471 3803 1475
rect 219 1403 223 1407
rect 259 1407 263 1411
rect 803 1407 807 1411
rect 811 1407 815 1411
rect 1099 1407 1103 1411
rect 1975 1401 1979 1405
rect 2167 1400 2171 1404
rect 2303 1400 2307 1404
rect 2439 1400 2443 1404
rect 2575 1400 2579 1404
rect 2711 1400 2715 1404
rect 2847 1400 2851 1404
rect 2983 1400 2987 1404
rect 3119 1400 3123 1404
rect 3255 1400 3259 1404
rect 3799 1401 3803 1405
rect 1975 1384 1979 1388
rect 2139 1385 2143 1389
rect 2275 1385 2279 1389
rect 2411 1385 2415 1389
rect 2547 1385 2551 1389
rect 2683 1385 2687 1389
rect 2819 1385 2823 1389
rect 2955 1385 2959 1389
rect 3091 1385 3095 1389
rect 3227 1385 3231 1389
rect 3799 1384 3803 1388
rect 259 1371 260 1375
rect 260 1371 263 1375
rect 387 1371 391 1375
rect 811 1371 812 1375
rect 812 1371 815 1375
rect 1099 1371 1100 1375
rect 1100 1371 1103 1375
rect 1411 1371 1415 1375
rect 2259 1375 2263 1379
rect 2419 1375 2423 1379
rect 2699 1375 2703 1379
rect 2835 1375 2839 1379
rect 2971 1375 2975 1379
rect 3107 1375 3111 1379
rect 3243 1375 3247 1379
rect 3355 1375 3356 1379
rect 3356 1375 3359 1379
rect 5307 1371 5311 1375
rect 5483 1375 5487 1379
rect 111 1364 115 1368
rect 131 1363 135 1367
rect 395 1363 399 1367
rect 683 1363 687 1367
rect 971 1363 975 1367
rect 1259 1363 1263 1367
rect 1935 1364 1939 1368
rect 111 1347 115 1351
rect 159 1348 163 1352
rect 423 1348 427 1352
rect 711 1348 715 1352
rect 999 1348 1003 1352
rect 1287 1348 1291 1352
rect 1935 1347 1939 1351
rect 2419 1343 2423 1347
rect 2499 1343 2503 1347
rect 2635 1343 2639 1347
rect 2699 1343 2703 1347
rect 2835 1343 2839 1347
rect 2971 1343 2975 1347
rect 3107 1343 3111 1347
rect 3243 1343 3247 1347
rect 4935 1339 4936 1343
rect 4936 1339 4939 1343
rect 5483 1339 5484 1343
rect 5484 1339 5487 1343
rect 5587 1339 5591 1343
rect 3839 1332 3843 1336
rect 4811 1331 4815 1335
rect 4947 1331 4951 1335
rect 5083 1331 5087 1335
rect 5219 1331 5223 1335
rect 5355 1331 5359 1335
rect 5491 1331 5495 1335
rect 5663 1332 5667 1336
rect 3839 1315 3843 1319
rect 4839 1316 4843 1320
rect 4975 1316 4979 1320
rect 5111 1316 5115 1320
rect 5247 1316 5251 1320
rect 5383 1316 5387 1320
rect 5519 1316 5523 1320
rect 5663 1315 5667 1319
rect 2247 1295 2251 1299
rect 2259 1295 2263 1299
rect 2531 1295 2535 1299
rect 2707 1295 2711 1299
rect 111 1289 115 1293
rect 159 1288 163 1292
rect 455 1288 459 1292
rect 775 1288 779 1292
rect 1095 1288 1099 1292
rect 1423 1288 1427 1292
rect 1935 1289 1939 1293
rect 3355 1291 3359 1295
rect 3555 1291 3559 1295
rect 3595 1295 3599 1299
rect 111 1272 115 1276
rect 131 1273 135 1277
rect 427 1273 431 1277
rect 747 1273 751 1277
rect 1067 1273 1071 1277
rect 1395 1273 1399 1277
rect 1935 1272 1939 1276
rect 219 1263 223 1267
rect 299 1263 303 1267
rect 1083 1263 1087 1267
rect 835 1255 839 1259
rect 2259 1259 2260 1263
rect 2260 1259 2263 1263
rect 2531 1259 2532 1263
rect 2532 1259 2535 1263
rect 2707 1259 2711 1263
rect 2723 1259 2727 1263
rect 3015 1259 3016 1263
rect 3016 1259 3019 1263
rect 3595 1259 3596 1263
rect 3596 1259 3599 1263
rect 3739 1259 3743 1263
rect 1975 1252 1979 1256
rect 2131 1251 2135 1255
rect 2267 1251 2271 1255
rect 2403 1251 2407 1255
rect 2555 1251 2559 1255
rect 2715 1251 2719 1255
rect 2891 1251 2895 1255
rect 3075 1251 3079 1255
rect 3267 1251 3271 1255
rect 3467 1251 3471 1255
rect 3651 1251 3655 1255
rect 3799 1252 3803 1256
rect 3839 1253 3843 1257
rect 4735 1252 4739 1256
rect 4879 1252 4883 1256
rect 5031 1252 5035 1256
rect 5191 1252 5195 1256
rect 5359 1252 5363 1256
rect 5527 1252 5531 1256
rect 5663 1253 5667 1257
rect 299 1231 303 1235
rect 515 1231 519 1235
rect 835 1231 839 1235
rect 1083 1231 1087 1235
rect 1411 1231 1415 1235
rect 1975 1235 1979 1239
rect 2159 1236 2163 1240
rect 2295 1236 2299 1240
rect 2431 1236 2435 1240
rect 2583 1236 2587 1240
rect 2743 1236 2747 1240
rect 2919 1236 2923 1240
rect 3103 1236 3107 1240
rect 3295 1236 3299 1240
rect 3495 1236 3499 1240
rect 3679 1236 3683 1240
rect 3799 1235 3803 1239
rect 3839 1236 3843 1240
rect 4707 1237 4711 1241
rect 4851 1237 4855 1241
rect 5003 1237 5007 1241
rect 5163 1237 5167 1241
rect 5331 1237 5335 1241
rect 5499 1237 5503 1241
rect 5663 1236 5667 1240
rect 4859 1227 4863 1231
rect 5019 1227 5023 1231
rect 4795 1219 4799 1223
rect 5307 1227 5311 1231
rect 5319 1227 5323 1231
rect 5619 1227 5623 1231
rect 2247 1211 2251 1215
rect 2811 1203 2815 1207
rect 4795 1195 4799 1199
rect 4935 1195 4939 1199
rect 5019 1195 5023 1199
rect 5319 1195 5323 1199
rect 5407 1195 5411 1199
rect 5587 1195 5591 1199
rect 1975 1177 1979 1181
rect 2023 1176 2027 1180
rect 2239 1176 2243 1180
rect 2479 1176 2483 1180
rect 2719 1176 2723 1180
rect 2959 1176 2963 1180
rect 3207 1176 3211 1180
rect 3455 1176 3459 1180
rect 3679 1176 3683 1180
rect 3799 1177 3803 1181
rect 259 1159 263 1163
rect 459 1159 463 1163
rect 1651 1159 1655 1163
rect 1975 1160 1979 1164
rect 1995 1161 1999 1165
rect 2211 1161 2215 1165
rect 2451 1161 2455 1165
rect 2691 1161 2695 1165
rect 2931 1161 2935 1165
rect 3179 1161 3183 1165
rect 3427 1161 3431 1165
rect 3651 1161 3655 1165
rect 3799 1160 3803 1164
rect 271 1151 275 1155
rect 1759 1151 1763 1155
rect 2227 1151 2231 1155
rect 2467 1151 2471 1155
rect 2707 1151 2711 1155
rect 2811 1151 2815 1155
rect 3083 1151 3087 1155
rect 3443 1151 3447 1155
rect 3555 1151 3556 1155
rect 3556 1151 3559 1155
rect 4035 1139 4039 1143
rect 4387 1135 4391 1139
rect 4427 1139 4431 1143
rect 4867 1135 4871 1139
rect 4907 1139 4911 1143
rect 5371 1135 5375 1139
rect 5619 1139 5623 1143
rect 259 1123 260 1127
rect 260 1123 263 1127
rect 459 1123 460 1127
rect 460 1123 463 1127
rect 515 1123 519 1127
rect 939 1123 943 1127
rect 1651 1123 1652 1127
rect 1652 1123 1655 1127
rect 111 1116 115 1120
rect 131 1115 135 1119
rect 331 1115 335 1119
rect 563 1115 567 1119
rect 803 1115 807 1119
rect 1043 1115 1047 1119
rect 1283 1115 1287 1119
rect 1523 1115 1527 1119
rect 1771 1115 1775 1119
rect 1935 1116 1939 1120
rect 2227 1119 2231 1123
rect 2467 1119 2471 1123
rect 2707 1119 2711 1123
rect 3015 1119 3019 1123
rect 3379 1119 3383 1123
rect 3443 1119 3447 1123
rect 3739 1119 3743 1123
rect 4387 1111 4391 1115
rect 111 1099 115 1103
rect 159 1100 163 1104
rect 359 1100 363 1104
rect 591 1100 595 1104
rect 831 1100 835 1104
rect 1071 1100 1075 1104
rect 1311 1100 1315 1104
rect 1551 1100 1555 1104
rect 1799 1100 1803 1104
rect 1935 1099 1939 1103
rect 4035 1103 4039 1107
rect 4131 1103 4135 1107
rect 4427 1103 4428 1107
rect 4428 1103 4431 1107
rect 4747 1103 4751 1107
rect 4907 1103 4908 1107
rect 4908 1103 4911 1107
rect 5407 1103 5408 1107
rect 5408 1103 5411 1107
rect 5603 1103 5607 1107
rect 3839 1096 3843 1100
rect 3859 1095 3863 1099
rect 4067 1095 4071 1099
rect 4299 1095 4303 1099
rect 4539 1095 4543 1099
rect 4779 1095 4783 1099
rect 5027 1095 5031 1099
rect 5283 1095 5287 1099
rect 5515 1095 5519 1099
rect 5663 1096 5667 1100
rect 3839 1079 3843 1083
rect 3887 1080 3891 1084
rect 4095 1080 4099 1084
rect 4327 1080 4331 1084
rect 4567 1080 4571 1084
rect 4807 1080 4811 1084
rect 5055 1080 5059 1084
rect 5311 1080 5315 1084
rect 5543 1080 5547 1084
rect 5663 1079 5667 1083
rect 3083 1047 3087 1051
rect 111 1041 115 1045
rect 263 1040 267 1044
rect 439 1040 443 1044
rect 615 1040 619 1044
rect 783 1040 787 1044
rect 951 1040 955 1044
rect 1111 1040 1115 1044
rect 1271 1040 1275 1044
rect 1431 1040 1435 1044
rect 1591 1040 1595 1044
rect 1751 1040 1755 1044
rect 1935 1041 1939 1045
rect 3331 1043 3335 1047
rect 3371 1047 3375 1051
rect 111 1024 115 1028
rect 235 1025 239 1029
rect 411 1025 415 1029
rect 587 1025 591 1029
rect 755 1025 759 1029
rect 923 1025 927 1029
rect 1083 1025 1087 1029
rect 1243 1025 1247 1029
rect 1403 1025 1407 1029
rect 1563 1025 1567 1029
rect 1723 1025 1727 1029
rect 1935 1024 1939 1028
rect 3839 1021 3843 1025
rect 3887 1020 3891 1024
rect 271 1015 275 1019
rect 659 1015 663 1019
rect 747 1015 751 1019
rect 911 1015 915 1019
rect 1259 1015 1263 1019
rect 1419 1015 1423 1019
rect 1579 1015 1583 1019
rect 1739 1015 1743 1019
rect 1759 1015 1763 1019
rect 4071 1020 4075 1024
rect 4279 1020 4283 1024
rect 4511 1020 4515 1024
rect 4759 1020 4763 1024
rect 5023 1020 5027 1024
rect 5295 1020 5299 1024
rect 5543 1020 5547 1024
rect 5663 1021 5667 1025
rect 2987 1011 2991 1015
rect 3371 1011 3372 1015
rect 3372 1011 3375 1015
rect 3379 1011 3383 1015
rect 1975 1004 1979 1008
rect 3091 1003 3095 1007
rect 3243 1003 3247 1007
rect 3395 1003 3399 1007
rect 3799 1004 3803 1008
rect 3839 1004 3843 1008
rect 3859 1005 3863 1009
rect 4043 1005 4047 1009
rect 4251 1005 4255 1009
rect 4483 1005 4487 1009
rect 4731 1005 4735 1009
rect 4995 1005 4999 1009
rect 5267 1005 5271 1009
rect 5515 1005 5519 1009
rect 5663 1004 5667 1008
rect 3963 995 3967 999
rect 4019 995 4023 999
rect 4499 995 4503 999
rect 4611 995 4612 999
rect 4612 995 4615 999
rect 5011 995 5015 999
rect 5371 995 5375 999
rect 5611 995 5615 999
rect 499 983 503 987
rect 747 983 751 987
rect 911 983 915 987
rect 939 983 943 987
rect 1259 983 1263 987
rect 1419 983 1423 987
rect 1579 983 1583 987
rect 1739 983 1743 987
rect 1975 987 1979 991
rect 3119 988 3123 992
rect 3271 988 3275 992
rect 3423 988 3427 992
rect 3799 987 3803 991
rect 4339 987 4343 991
rect 4019 963 4023 967
rect 4131 963 4135 967
rect 4339 963 4343 967
rect 4499 963 4503 967
rect 4747 963 4751 967
rect 5011 963 5015 967
rect 5295 963 5299 967
rect 5603 963 5607 967
rect 315 927 319 931
rect 355 931 359 935
rect 659 931 663 935
rect 667 931 671 935
rect 843 931 847 935
rect 1019 931 1023 935
rect 1607 931 1611 935
rect 3963 915 3967 919
rect 4267 911 4271 915
rect 4307 915 4311 919
rect 4611 915 4615 919
rect 4867 915 4871 919
rect 5531 911 5535 915
rect 1975 901 1979 905
rect 2047 900 2051 904
rect 355 895 356 899
rect 356 895 359 899
rect 499 895 503 899
rect 667 895 668 899
rect 668 895 671 899
rect 843 895 844 899
rect 844 895 847 899
rect 1019 895 1020 899
rect 1020 895 1023 899
rect 1227 895 1231 899
rect 1607 895 1611 899
rect 2351 900 2355 904
rect 2647 900 2651 904
rect 2927 900 2931 904
rect 3207 900 3211 904
rect 3495 900 3499 904
rect 3799 901 3803 905
rect 111 888 115 892
rect 227 887 231 891
rect 379 887 383 891
rect 539 887 543 891
rect 715 887 719 891
rect 891 887 895 891
rect 1075 887 1079 891
rect 1259 887 1263 891
rect 1443 887 1447 891
rect 1627 887 1631 891
rect 1787 887 1791 891
rect 1935 888 1939 892
rect 1975 884 1979 888
rect 2019 885 2023 889
rect 2323 885 2327 889
rect 2619 885 2623 889
rect 2899 885 2903 889
rect 3179 885 3183 889
rect 3467 885 3471 889
rect 3799 884 3803 888
rect 4267 887 4271 891
rect 111 871 115 875
rect 255 872 259 876
rect 407 872 411 876
rect 567 872 571 876
rect 743 872 747 876
rect 919 872 923 876
rect 1103 872 1107 876
rect 1287 872 1291 876
rect 1471 872 1475 876
rect 1655 872 1659 876
rect 1815 872 1819 876
rect 1935 871 1939 875
rect 2167 875 2171 879
rect 2747 875 2748 879
rect 2748 875 2751 879
rect 2831 875 2835 879
rect 3331 875 3335 879
rect 3379 875 3383 879
rect 4267 879 4271 883
rect 4307 879 4308 883
rect 4308 879 4311 883
rect 4547 879 4551 883
rect 3839 872 3843 876
rect 3971 871 3975 875
rect 4179 871 4183 875
rect 4403 871 4407 875
rect 4643 871 4647 875
rect 4867 875 4871 879
rect 5295 879 5296 883
rect 5296 879 5299 883
rect 4899 871 4903 875
rect 5171 871 5175 875
rect 5443 871 5447 875
rect 5663 872 5667 876
rect 3839 855 3843 859
rect 3999 856 4003 860
rect 4207 856 4211 860
rect 4431 856 4435 860
rect 4671 856 4675 860
rect 4927 856 4931 860
rect 5199 856 5203 860
rect 5471 856 5475 860
rect 5663 855 5667 859
rect 2167 843 2171 847
rect 2411 843 2415 847
rect 2831 843 2835 847
rect 2987 843 2991 847
rect 3379 843 3383 847
rect 3555 843 3559 847
rect 111 797 115 801
rect 375 796 379 800
rect 655 796 659 800
rect 943 796 947 800
rect 1239 796 1243 800
rect 1535 796 1539 800
rect 1815 796 1819 800
rect 1935 797 1939 801
rect 1943 795 1947 799
rect 2123 795 2127 799
rect 2379 795 2383 799
rect 2747 795 2751 799
rect 2899 795 2903 799
rect 3315 791 3319 795
rect 3355 795 3359 799
rect 3839 797 3843 801
rect 3887 796 3891 800
rect 4047 796 4051 800
rect 4279 796 4283 800
rect 4559 796 4563 800
rect 4879 796 4883 800
rect 5223 796 5227 800
rect 5543 796 5547 800
rect 5663 797 5667 801
rect 3867 791 3871 795
rect 111 780 115 784
rect 347 781 351 785
rect 627 781 631 785
rect 915 781 919 785
rect 1211 781 1215 785
rect 1507 781 1511 785
rect 1787 781 1791 785
rect 1935 780 1939 784
rect 3839 780 3843 784
rect 3859 781 3863 785
rect 4019 781 4023 785
rect 4251 781 4255 785
rect 4531 781 4535 785
rect 4851 781 4855 785
rect 5195 781 5199 785
rect 5515 781 5519 785
rect 5663 780 5667 784
rect 643 771 647 775
rect 315 763 319 767
rect 1019 771 1023 775
rect 1135 771 1139 775
rect 1803 771 1807 775
rect 1943 771 1947 775
rect 3315 767 3319 771
rect 3987 771 3988 775
rect 3988 771 3991 775
rect 4027 771 4031 775
rect 4867 771 4871 775
rect 5211 771 5215 775
rect 431 739 435 743
rect 643 739 647 743
rect 1135 739 1139 743
rect 1227 739 1231 743
rect 1911 755 1915 759
rect 2123 759 2124 763
rect 2124 759 2127 763
rect 2379 759 2380 763
rect 2380 759 2383 763
rect 2411 759 2415 763
rect 2899 759 2900 763
rect 2900 759 2903 763
rect 3299 759 3303 763
rect 3355 759 3356 763
rect 3356 759 3359 763
rect 3555 759 3559 763
rect 5531 771 5535 775
rect 1975 752 1979 756
rect 1995 751 1999 755
rect 2251 751 2255 755
rect 2523 751 2527 755
rect 2771 751 2775 755
rect 3003 751 3007 755
rect 3227 751 3231 755
rect 3451 751 3455 755
rect 3651 751 3655 755
rect 3799 752 3803 756
rect 1803 739 1807 743
rect 1975 735 1979 739
rect 2023 736 2027 740
rect 2279 736 2283 740
rect 2551 736 2555 740
rect 2799 736 2803 740
rect 3031 736 3035 740
rect 3255 736 3259 740
rect 3479 736 3483 740
rect 3679 736 3683 740
rect 3799 735 3803 739
rect 4027 739 4031 743
rect 4267 739 4271 743
rect 4547 739 4551 743
rect 4867 739 4871 743
rect 5211 739 5215 743
rect 5611 739 5615 743
rect 259 691 263 695
rect 475 691 479 695
rect 811 691 815 695
rect 1019 691 1023 695
rect 1275 687 1279 691
rect 1151 675 1155 679
rect 3947 679 3951 683
rect 3987 683 3991 687
rect 4699 683 4703 687
rect 4899 683 4903 687
rect 5123 683 5127 687
rect 5547 679 5551 683
rect 259 655 260 659
rect 260 655 263 659
rect 431 655 432 659
rect 432 655 435 659
rect 811 655 812 659
rect 812 655 815 659
rect 987 655 988 659
rect 988 655 991 659
rect 1151 655 1152 659
rect 1152 655 1155 659
rect 1911 655 1912 659
rect 1912 655 1915 659
rect 4219 655 4223 659
rect 111 648 115 652
rect 131 647 135 651
rect 307 647 311 651
rect 499 647 503 651
rect 683 647 687 651
rect 859 647 863 651
rect 1027 647 1031 651
rect 1187 647 1191 651
rect 1339 647 1343 651
rect 1491 647 1495 651
rect 1651 647 1655 651
rect 1787 647 1791 651
rect 1935 648 1939 652
rect 3867 647 3871 651
rect 4699 647 4700 651
rect 4700 647 4703 651
rect 4899 647 4900 651
rect 4900 647 4903 651
rect 5123 647 5124 651
rect 5124 647 5127 651
rect 5335 647 5339 651
rect 5595 647 5599 651
rect 3839 640 3843 644
rect 3859 639 3863 643
rect 3995 639 3999 643
rect 4131 639 4135 643
rect 4267 639 4271 643
rect 4403 639 4407 643
rect 4571 639 4575 643
rect 4771 639 4775 643
rect 4995 639 4999 643
rect 5227 639 5231 643
rect 5459 639 5463 643
rect 5663 640 5667 644
rect 111 631 115 635
rect 159 632 163 636
rect 335 632 339 636
rect 527 632 531 636
rect 711 632 715 636
rect 887 632 891 636
rect 1055 632 1059 636
rect 1215 632 1219 636
rect 1367 632 1371 636
rect 1519 632 1523 636
rect 1679 632 1683 636
rect 1815 632 1819 636
rect 1935 631 1939 635
rect 3839 623 3843 627
rect 3887 624 3891 628
rect 4023 624 4027 628
rect 4159 624 4163 628
rect 4295 624 4299 628
rect 4431 624 4435 628
rect 4599 624 4603 628
rect 4799 624 4803 628
rect 5023 624 5027 628
rect 5255 624 5259 628
rect 5487 624 5491 628
rect 5663 623 5667 627
rect 5335 607 5339 611
rect 111 573 115 577
rect 159 572 163 576
rect 375 572 379 576
rect 599 572 603 576
rect 807 572 811 576
rect 999 572 1003 576
rect 1175 572 1179 576
rect 1343 572 1347 576
rect 1511 572 1515 576
rect 1671 572 1675 576
rect 1815 572 1819 576
rect 1935 573 1939 577
rect 3839 565 3843 569
rect 3887 564 3891 568
rect 4023 564 4027 568
rect 4159 564 4163 568
rect 4295 564 4299 568
rect 4479 564 4483 568
rect 4695 564 4699 568
rect 4935 564 4939 568
rect 5191 564 5195 568
rect 5447 564 5451 568
rect 5663 565 5667 569
rect 111 556 115 560
rect 131 557 135 561
rect 347 557 351 561
rect 571 557 575 561
rect 779 557 783 561
rect 971 557 975 561
rect 1147 557 1151 561
rect 1315 557 1319 561
rect 1483 557 1487 561
rect 1643 557 1647 561
rect 1787 557 1791 561
rect 1935 556 1939 560
rect 363 547 367 551
rect 475 547 476 551
rect 476 547 479 551
rect 699 547 700 551
rect 700 547 703 551
rect 1275 547 1276 551
rect 1276 547 1279 551
rect 1303 547 1307 551
rect 1491 547 1495 551
rect 1779 547 1783 551
rect 1975 545 1979 549
rect 3311 544 3315 548
rect 3447 544 3451 548
rect 3583 544 3587 548
rect 3799 545 3803 549
rect 3839 548 3843 552
rect 3859 549 3863 553
rect 3995 549 3999 553
rect 4131 549 4135 553
rect 4267 549 4271 553
rect 4451 549 4455 553
rect 4667 549 4671 553
rect 4907 549 4911 553
rect 5163 549 5167 553
rect 5419 549 5423 553
rect 5663 548 5667 552
rect 3947 539 3951 543
rect 4003 539 4007 543
rect 4467 539 4471 543
rect 4683 539 4687 543
rect 4923 539 4927 543
rect 5179 539 5183 543
rect 5187 539 5191 543
rect 5547 539 5548 543
rect 5548 539 5551 543
rect 1975 528 1979 532
rect 3283 529 3287 533
rect 3419 529 3423 533
rect 3555 529 3559 533
rect 3799 528 3803 532
rect 227 515 231 519
rect 363 515 367 519
rect 987 515 991 519
rect 1303 515 1307 519
rect 1491 515 1495 519
rect 1779 515 1783 519
rect 1883 515 1887 519
rect 3435 519 3439 523
rect 3571 519 3575 523
rect 3643 519 3647 523
rect 4003 507 4007 511
rect 4219 507 4223 511
rect 4467 507 4471 511
rect 4683 507 4687 511
rect 4923 507 4927 511
rect 5179 507 5183 511
rect 5435 507 5439 511
rect 3299 487 3303 491
rect 3435 487 3439 491
rect 3571 487 3575 491
rect 4571 491 4575 495
rect 5187 491 5191 495
rect 351 467 355 471
rect 559 467 563 471
rect 699 467 703 471
rect 891 467 895 471
rect 1235 467 1239 471
rect 4571 447 4575 451
rect 4579 447 4583 451
rect 4779 447 4783 451
rect 4987 447 4991 451
rect 2259 439 2263 443
rect 2475 439 2479 443
rect 2667 439 2671 443
rect 227 431 231 435
rect 351 431 355 435
rect 891 431 892 435
rect 892 431 895 435
rect 1235 431 1236 435
rect 1236 431 1239 435
rect 1519 431 1523 435
rect 1883 431 1887 435
rect 3011 435 3015 439
rect 3051 439 3055 443
rect 3243 439 3247 443
rect 3635 439 3639 443
rect 3643 439 3647 443
rect 5595 443 5599 447
rect 111 424 115 428
rect 131 423 135 427
rect 427 423 431 427
rect 763 423 767 427
rect 1107 423 1111 427
rect 1459 423 1463 427
rect 1787 423 1791 427
rect 1935 424 1939 428
rect 2855 423 2859 427
rect 111 407 115 411
rect 159 408 163 412
rect 455 408 459 412
rect 791 408 795 412
rect 1135 408 1139 412
rect 1487 408 1491 412
rect 1815 408 1819 412
rect 1935 407 1939 411
rect 3011 411 3015 415
rect 2475 403 2476 407
rect 2476 403 2479 407
rect 2667 403 2668 407
rect 2668 403 2671 407
rect 2855 403 2856 407
rect 2856 403 2859 407
rect 3051 403 3052 407
rect 3052 403 3055 407
rect 3243 403 3244 407
rect 3244 403 3247 407
rect 3423 403 3424 407
rect 3424 403 3427 407
rect 4579 411 4580 415
rect 4580 411 4583 415
rect 4779 411 4780 415
rect 4780 411 4783 415
rect 4987 411 4988 415
rect 4988 411 4991 415
rect 5035 411 5039 415
rect 5435 411 5439 415
rect 5603 411 5607 415
rect 3635 403 3639 407
rect 3839 404 3843 408
rect 4451 403 4455 407
rect 4651 403 4655 407
rect 4859 403 4863 407
rect 5067 403 5071 407
rect 5283 403 5287 407
rect 5507 403 5511 407
rect 5663 404 5667 408
rect 1975 396 1979 400
rect 1995 395 1999 399
rect 2155 395 2159 399
rect 2347 395 2351 399
rect 2539 395 2543 399
rect 2731 395 2735 399
rect 2923 395 2927 399
rect 3115 395 3119 399
rect 3299 395 3303 399
rect 3483 395 3487 399
rect 3651 395 3655 399
rect 3799 396 3803 400
rect 3839 387 3843 391
rect 4479 388 4483 392
rect 4679 388 4683 392
rect 4887 388 4891 392
rect 5095 388 5099 392
rect 5311 388 5315 392
rect 5535 388 5539 392
rect 5663 387 5667 391
rect 1975 379 1979 383
rect 2023 380 2027 384
rect 2183 380 2187 384
rect 2375 380 2379 384
rect 2567 380 2571 384
rect 2759 380 2763 384
rect 2951 380 2955 384
rect 3143 380 3147 384
rect 3327 380 3331 384
rect 3511 380 3515 384
rect 3679 380 3683 384
rect 3799 379 3803 383
rect 111 333 115 337
rect 239 332 243 336
rect 391 332 395 336
rect 551 332 555 336
rect 711 332 715 336
rect 871 332 875 336
rect 1031 332 1035 336
rect 1935 333 1939 337
rect 3839 325 3843 329
rect 4751 324 4755 328
rect 4911 324 4915 328
rect 5071 324 5075 328
rect 5231 324 5235 328
rect 5399 324 5403 328
rect 5543 324 5547 328
rect 5663 325 5667 329
rect 111 316 115 320
rect 211 317 215 321
rect 363 317 367 321
rect 523 317 527 321
rect 683 317 687 321
rect 843 317 847 321
rect 1003 317 1007 321
rect 1935 316 1939 320
rect 379 307 383 311
rect 539 307 543 311
rect 559 307 563 311
rect 811 307 812 311
rect 812 307 815 311
rect 3839 308 3843 312
rect 4723 309 4727 313
rect 4883 309 4887 313
rect 5043 309 5047 313
rect 5203 309 5207 313
rect 5371 309 5375 313
rect 5515 309 5519 313
rect 5663 308 5667 312
rect 1975 297 1979 301
rect 2047 296 2051 300
rect 2183 296 2187 300
rect 2319 296 2323 300
rect 2455 296 2459 300
rect 2591 296 2595 300
rect 2727 296 2731 300
rect 2863 296 2867 300
rect 2999 296 3003 300
rect 3135 296 3139 300
rect 3271 296 3275 300
rect 3407 296 3411 300
rect 3543 296 3547 300
rect 3679 296 3683 300
rect 3799 297 3803 301
rect 4859 299 4863 303
rect 5219 299 5223 303
rect 5131 291 5135 295
rect 5619 299 5623 303
rect 1975 280 1979 284
rect 2019 281 2023 285
rect 2155 281 2159 285
rect 2291 281 2295 285
rect 2427 281 2431 285
rect 2563 281 2567 285
rect 2699 281 2703 285
rect 2835 281 2839 285
rect 2971 281 2975 285
rect 3107 281 3111 285
rect 3243 281 3247 285
rect 3379 281 3383 285
rect 3515 281 3519 285
rect 3651 281 3655 285
rect 3799 280 3803 284
rect 271 275 275 279
rect 379 275 383 279
rect 539 275 543 279
rect 1519 275 1523 279
rect 2259 271 2263 275
rect 2307 271 2311 275
rect 2443 271 2447 275
rect 2531 271 2535 275
rect 2987 271 2991 275
rect 3123 271 3127 275
rect 3235 271 3236 275
rect 3236 271 3239 275
rect 2923 263 2927 267
rect 3531 271 3535 275
rect 3667 271 3671 275
rect 3331 263 3335 267
rect 4859 267 4863 271
rect 5035 267 5039 271
rect 5131 267 5135 271
rect 5219 267 5223 271
rect 5387 267 5391 271
rect 5603 267 5607 271
rect 2107 239 2111 243
rect 2307 239 2311 243
rect 2443 239 2447 243
rect 2843 239 2847 243
rect 2923 239 2927 243
rect 2987 239 2991 243
rect 3123 239 3127 243
rect 3331 239 3335 243
rect 3423 239 3427 243
rect 3531 239 3535 243
rect 3667 239 3671 243
rect 1203 207 1207 211
rect 811 195 815 199
rect 3235 191 3239 195
rect 2491 171 2495 175
rect 2531 175 2535 179
rect 3307 171 3311 175
rect 4827 179 4831 183
rect 5467 175 5471 179
rect 5619 179 5623 183
rect 271 159 272 163
rect 272 159 275 163
rect 1203 159 1207 163
rect 111 152 115 156
rect 147 151 151 155
rect 283 151 287 155
rect 419 151 423 155
rect 555 151 559 155
rect 691 151 695 155
rect 827 151 831 155
rect 963 151 967 155
rect 1099 151 1103 155
rect 1935 152 1939 156
rect 2491 147 2495 151
rect 111 135 115 139
rect 175 136 179 140
rect 311 136 315 140
rect 447 136 451 140
rect 583 136 587 140
rect 719 136 723 140
rect 855 136 859 140
rect 991 136 995 140
rect 1127 136 1131 140
rect 1935 135 1939 139
rect 2107 139 2111 143
rect 2843 147 2847 151
rect 3307 147 3311 151
rect 4827 143 4828 147
rect 4828 143 4831 147
rect 5387 143 5391 147
rect 5467 143 5471 147
rect 1975 132 1979 136
rect 1995 131 1999 135
rect 2131 131 2135 135
rect 2267 131 2271 135
rect 2403 131 2407 135
rect 2539 131 2543 135
rect 2675 131 2679 135
rect 2811 131 2815 135
rect 2947 131 2951 135
rect 3083 131 3087 135
rect 3219 131 3223 135
rect 3355 131 3359 135
rect 3491 131 3495 135
rect 3627 131 3631 135
rect 3799 132 3803 136
rect 3839 136 3843 140
rect 4291 135 4295 139
rect 4427 135 4431 139
rect 4563 135 4567 139
rect 4699 135 4703 139
rect 4835 135 4839 139
rect 4971 135 4975 139
rect 5107 135 5111 139
rect 5243 135 5247 139
rect 5379 135 5383 139
rect 5515 135 5519 139
rect 5663 136 5667 140
rect 1975 115 1979 119
rect 2023 116 2027 120
rect 2159 116 2163 120
rect 2295 116 2299 120
rect 2431 116 2435 120
rect 2567 116 2571 120
rect 2703 116 2707 120
rect 2839 116 2843 120
rect 2975 116 2979 120
rect 3111 116 3115 120
rect 3247 116 3251 120
rect 3383 116 3387 120
rect 3519 116 3523 120
rect 3655 116 3659 120
rect 3799 115 3803 119
rect 3839 119 3843 123
rect 4319 120 4323 124
rect 4455 120 4459 124
rect 4591 120 4595 124
rect 4727 120 4731 124
rect 4863 120 4867 124
rect 4999 120 5003 124
rect 5135 120 5139 124
rect 5271 120 5275 124
rect 5407 120 5411 124
rect 5543 120 5547 124
rect 5663 119 5667 123
<< m3 >>
rect 111 5758 115 5759
rect 111 5753 115 5754
rect 131 5758 135 5759
rect 131 5753 135 5754
rect 267 5758 271 5759
rect 267 5753 271 5754
rect 403 5758 407 5759
rect 403 5753 407 5754
rect 1935 5758 1939 5759
rect 1935 5753 1939 5754
rect 112 5693 114 5753
rect 110 5692 116 5693
rect 132 5692 134 5753
rect 258 5735 264 5736
rect 258 5731 259 5735
rect 263 5731 264 5735
rect 258 5730 264 5731
rect 260 5700 262 5730
rect 258 5699 264 5700
rect 258 5695 259 5699
rect 263 5695 264 5699
rect 258 5694 264 5695
rect 268 5692 270 5753
rect 404 5692 406 5753
rect 422 5699 428 5700
rect 422 5695 423 5699
rect 427 5695 428 5699
rect 422 5694 428 5695
rect 110 5688 111 5692
rect 115 5688 116 5692
rect 110 5687 116 5688
rect 130 5691 136 5692
rect 130 5687 131 5691
rect 135 5687 136 5691
rect 130 5686 136 5687
rect 266 5691 272 5692
rect 266 5687 267 5691
rect 271 5687 272 5691
rect 266 5686 272 5687
rect 402 5691 408 5692
rect 402 5687 403 5691
rect 407 5687 408 5691
rect 402 5686 408 5687
rect 158 5676 164 5677
rect 110 5675 116 5676
rect 110 5671 111 5675
rect 115 5671 116 5675
rect 158 5672 159 5676
rect 163 5672 164 5676
rect 158 5671 164 5672
rect 294 5676 300 5677
rect 294 5672 295 5676
rect 299 5672 300 5676
rect 294 5671 300 5672
rect 110 5670 116 5671
rect 112 5647 114 5670
rect 160 5647 162 5671
rect 296 5647 298 5671
rect 111 5646 115 5647
rect 111 5641 115 5642
rect 159 5646 163 5647
rect 159 5641 163 5642
rect 295 5646 299 5647
rect 295 5641 299 5642
rect 343 5646 347 5647
rect 343 5641 347 5642
rect 112 5618 114 5641
rect 110 5617 116 5618
rect 344 5617 346 5641
rect 110 5613 111 5617
rect 115 5613 116 5617
rect 110 5612 116 5613
rect 342 5616 348 5617
rect 342 5612 343 5616
rect 347 5612 348 5616
rect 342 5611 348 5612
rect 314 5601 320 5602
rect 110 5600 116 5601
rect 110 5596 111 5600
rect 115 5596 116 5600
rect 314 5597 315 5601
rect 319 5597 320 5601
rect 314 5596 320 5597
rect 110 5595 116 5596
rect 112 5535 114 5595
rect 316 5535 318 5596
rect 424 5560 426 5694
rect 1936 5693 1938 5753
rect 3839 5694 3843 5695
rect 1934 5692 1940 5693
rect 1934 5688 1935 5692
rect 1939 5688 1940 5692
rect 1934 5687 1940 5688
rect 1975 5690 1979 5691
rect 1975 5685 1979 5686
rect 1995 5690 1999 5691
rect 1995 5685 1999 5686
rect 2171 5690 2175 5691
rect 2171 5685 2175 5686
rect 2371 5690 2375 5691
rect 2371 5685 2375 5686
rect 2563 5690 2567 5691
rect 2563 5685 2567 5686
rect 2747 5690 2751 5691
rect 2747 5685 2751 5686
rect 2931 5690 2935 5691
rect 2931 5685 2935 5686
rect 3107 5690 3111 5691
rect 3107 5685 3111 5686
rect 3275 5690 3279 5691
rect 3275 5685 3279 5686
rect 3443 5690 3447 5691
rect 3443 5685 3447 5686
rect 3619 5690 3623 5691
rect 3619 5685 3623 5686
rect 3799 5690 3803 5691
rect 3839 5689 3843 5690
rect 4467 5694 4471 5695
rect 4467 5689 4471 5690
rect 4603 5694 4607 5695
rect 4603 5689 4607 5690
rect 4739 5694 4743 5695
rect 4739 5689 4743 5690
rect 4875 5694 4879 5695
rect 4875 5689 4879 5690
rect 5663 5694 5667 5695
rect 5663 5689 5667 5690
rect 3799 5685 3803 5686
rect 430 5676 436 5677
rect 430 5672 431 5676
rect 435 5672 436 5676
rect 430 5671 436 5672
rect 1934 5675 1940 5676
rect 1934 5671 1935 5675
rect 1939 5671 1940 5675
rect 432 5647 434 5671
rect 1934 5670 1940 5671
rect 1936 5647 1938 5670
rect 431 5646 435 5647
rect 431 5641 435 5642
rect 535 5646 539 5647
rect 535 5641 539 5642
rect 735 5646 739 5647
rect 735 5641 739 5642
rect 943 5646 947 5647
rect 943 5641 947 5642
rect 1159 5646 1163 5647
rect 1159 5641 1163 5642
rect 1383 5646 1387 5647
rect 1383 5641 1387 5642
rect 1607 5646 1611 5647
rect 1607 5641 1611 5642
rect 1815 5646 1819 5647
rect 1815 5641 1819 5642
rect 1935 5646 1939 5647
rect 1935 5641 1939 5642
rect 536 5617 538 5641
rect 736 5617 738 5641
rect 944 5617 946 5641
rect 1160 5617 1162 5641
rect 1384 5617 1386 5641
rect 1608 5617 1610 5641
rect 1816 5617 1818 5641
rect 1936 5618 1938 5641
rect 1942 5631 1948 5632
rect 1942 5627 1943 5631
rect 1947 5627 1948 5631
rect 1942 5626 1948 5627
rect 1934 5617 1940 5618
rect 534 5616 540 5617
rect 534 5612 535 5616
rect 539 5612 540 5616
rect 534 5611 540 5612
rect 734 5616 740 5617
rect 734 5612 735 5616
rect 739 5612 740 5616
rect 734 5611 740 5612
rect 942 5616 948 5617
rect 942 5612 943 5616
rect 947 5612 948 5616
rect 942 5611 948 5612
rect 1158 5616 1164 5617
rect 1158 5612 1159 5616
rect 1163 5612 1164 5616
rect 1158 5611 1164 5612
rect 1382 5616 1388 5617
rect 1382 5612 1383 5616
rect 1387 5612 1388 5616
rect 1382 5611 1388 5612
rect 1606 5616 1612 5617
rect 1606 5612 1607 5616
rect 1611 5612 1612 5616
rect 1606 5611 1612 5612
rect 1814 5616 1820 5617
rect 1814 5612 1815 5616
rect 1819 5612 1820 5616
rect 1934 5613 1935 5617
rect 1939 5613 1940 5617
rect 1934 5612 1940 5613
rect 1814 5611 1820 5612
rect 506 5601 512 5602
rect 506 5597 507 5601
rect 511 5597 512 5601
rect 506 5596 512 5597
rect 706 5601 712 5602
rect 706 5597 707 5601
rect 711 5597 712 5601
rect 706 5596 712 5597
rect 914 5601 920 5602
rect 914 5597 915 5601
rect 919 5597 920 5601
rect 914 5596 920 5597
rect 1130 5601 1136 5602
rect 1130 5597 1131 5601
rect 1135 5597 1136 5601
rect 1130 5596 1136 5597
rect 1354 5601 1360 5602
rect 1354 5597 1355 5601
rect 1359 5597 1360 5601
rect 1354 5596 1360 5597
rect 1578 5601 1584 5602
rect 1578 5597 1579 5601
rect 1583 5597 1584 5601
rect 1578 5596 1584 5597
rect 1786 5601 1792 5602
rect 1786 5597 1787 5601
rect 1791 5597 1792 5601
rect 1786 5596 1792 5597
rect 1934 5600 1940 5601
rect 1934 5596 1935 5600
rect 1939 5596 1940 5600
rect 422 5559 428 5560
rect 422 5555 423 5559
rect 427 5555 428 5559
rect 422 5554 428 5555
rect 508 5535 510 5596
rect 522 5591 528 5592
rect 522 5587 523 5591
rect 527 5587 528 5591
rect 522 5586 528 5587
rect 524 5560 526 5586
rect 522 5559 528 5560
rect 522 5555 523 5559
rect 527 5555 528 5559
rect 522 5554 528 5555
rect 708 5535 710 5596
rect 722 5591 728 5592
rect 722 5587 723 5591
rect 727 5587 728 5591
rect 722 5586 728 5587
rect 724 5560 726 5586
rect 722 5559 728 5560
rect 722 5555 723 5559
rect 727 5555 728 5559
rect 722 5554 728 5555
rect 916 5535 918 5596
rect 930 5591 936 5592
rect 930 5587 931 5591
rect 935 5587 936 5591
rect 930 5586 936 5587
rect 932 5560 934 5586
rect 998 5583 1004 5584
rect 998 5579 999 5583
rect 1003 5579 1004 5583
rect 998 5578 1004 5579
rect 930 5559 936 5560
rect 930 5555 931 5559
rect 935 5555 936 5559
rect 930 5554 936 5555
rect 111 5534 115 5535
rect 111 5529 115 5530
rect 315 5534 319 5535
rect 315 5529 319 5530
rect 507 5534 511 5535
rect 507 5529 511 5530
rect 707 5534 711 5535
rect 707 5529 711 5530
rect 875 5534 879 5535
rect 875 5529 879 5530
rect 915 5534 919 5535
rect 915 5529 919 5530
rect 112 5469 114 5529
rect 110 5468 116 5469
rect 876 5468 878 5529
rect 1000 5512 1002 5578
rect 1132 5535 1134 5596
rect 1146 5591 1152 5592
rect 1146 5587 1147 5591
rect 1151 5587 1152 5591
rect 1146 5586 1152 5587
rect 1148 5560 1150 5586
rect 1146 5559 1152 5560
rect 1146 5555 1147 5559
rect 1151 5555 1152 5559
rect 1146 5554 1152 5555
rect 1356 5535 1358 5596
rect 1580 5535 1582 5596
rect 1788 5535 1790 5596
rect 1934 5595 1940 5596
rect 1936 5535 1938 5595
rect 1944 5560 1946 5626
rect 1976 5625 1978 5685
rect 1974 5624 1980 5625
rect 1996 5624 1998 5685
rect 2172 5624 2174 5685
rect 2372 5624 2374 5685
rect 2564 5624 2566 5685
rect 2650 5663 2656 5664
rect 2650 5659 2651 5663
rect 2655 5659 2656 5663
rect 2650 5658 2656 5659
rect 1974 5620 1975 5624
rect 1979 5620 1980 5624
rect 1974 5619 1980 5620
rect 1994 5623 2000 5624
rect 1994 5619 1995 5623
rect 1999 5619 2000 5623
rect 1994 5618 2000 5619
rect 2170 5623 2176 5624
rect 2170 5619 2171 5623
rect 2175 5619 2176 5623
rect 2170 5618 2176 5619
rect 2370 5623 2376 5624
rect 2370 5619 2371 5623
rect 2375 5619 2376 5623
rect 2370 5618 2376 5619
rect 2562 5623 2568 5624
rect 2562 5619 2563 5623
rect 2567 5619 2568 5623
rect 2562 5618 2568 5619
rect 2022 5608 2028 5609
rect 1974 5607 1980 5608
rect 1974 5603 1975 5607
rect 1979 5603 1980 5607
rect 2022 5604 2023 5608
rect 2027 5604 2028 5608
rect 2022 5603 2028 5604
rect 2198 5608 2204 5609
rect 2198 5604 2199 5608
rect 2203 5604 2204 5608
rect 2198 5603 2204 5604
rect 2398 5608 2404 5609
rect 2398 5604 2399 5608
rect 2403 5604 2404 5608
rect 2398 5603 2404 5604
rect 2590 5608 2596 5609
rect 2590 5604 2591 5608
rect 2595 5604 2596 5608
rect 2590 5603 2596 5604
rect 1974 5602 1980 5603
rect 1976 5579 1978 5602
rect 2024 5579 2026 5603
rect 2200 5579 2202 5603
rect 2400 5579 2402 5603
rect 2592 5579 2594 5603
rect 1975 5578 1979 5579
rect 1975 5573 1979 5574
rect 2023 5578 2027 5579
rect 2023 5573 2027 5574
rect 2199 5578 2203 5579
rect 2199 5573 2203 5574
rect 2375 5578 2379 5579
rect 2375 5573 2379 5574
rect 2399 5578 2403 5579
rect 2399 5573 2403 5574
rect 2591 5578 2595 5579
rect 2591 5573 2595 5574
rect 2607 5578 2611 5579
rect 2607 5573 2611 5574
rect 1942 5559 1948 5560
rect 1942 5555 1943 5559
rect 1947 5555 1948 5559
rect 1942 5554 1948 5555
rect 1976 5550 1978 5573
rect 1974 5549 1980 5550
rect 2376 5549 2378 5573
rect 2608 5549 2610 5573
rect 1974 5545 1975 5549
rect 1979 5545 1980 5549
rect 1974 5544 1980 5545
rect 2374 5548 2380 5549
rect 2374 5544 2375 5548
rect 2379 5544 2380 5548
rect 2374 5543 2380 5544
rect 2606 5548 2612 5549
rect 2606 5544 2607 5548
rect 2611 5544 2612 5548
rect 2606 5543 2612 5544
rect 1011 5534 1015 5535
rect 1011 5529 1015 5530
rect 1131 5534 1135 5535
rect 1131 5529 1135 5530
rect 1147 5534 1151 5535
rect 1147 5529 1151 5530
rect 1291 5534 1295 5535
rect 1291 5529 1295 5530
rect 1355 5534 1359 5535
rect 1355 5529 1359 5530
rect 1435 5534 1439 5535
rect 1435 5529 1439 5530
rect 1579 5534 1583 5535
rect 1579 5529 1583 5530
rect 1723 5534 1727 5535
rect 1723 5529 1727 5530
rect 1787 5534 1791 5535
rect 1935 5534 1939 5535
rect 1787 5529 1791 5530
rect 1846 5531 1852 5532
rect 998 5511 1004 5512
rect 998 5507 999 5511
rect 1003 5507 1004 5511
rect 998 5506 1004 5507
rect 1012 5468 1014 5529
rect 1148 5468 1150 5529
rect 1270 5475 1276 5476
rect 1270 5471 1271 5475
rect 1275 5471 1276 5475
rect 1270 5470 1276 5471
rect 110 5464 111 5468
rect 115 5464 116 5468
rect 110 5463 116 5464
rect 874 5467 880 5468
rect 874 5463 875 5467
rect 879 5463 880 5467
rect 874 5462 880 5463
rect 1010 5467 1016 5468
rect 1010 5463 1011 5467
rect 1015 5463 1016 5467
rect 1010 5462 1016 5463
rect 1146 5467 1152 5468
rect 1146 5463 1147 5467
rect 1151 5463 1152 5467
rect 1146 5462 1152 5463
rect 902 5452 908 5453
rect 110 5451 116 5452
rect 110 5447 111 5451
rect 115 5447 116 5451
rect 902 5448 903 5452
rect 907 5448 908 5452
rect 902 5447 908 5448
rect 1038 5452 1044 5453
rect 1038 5448 1039 5452
rect 1043 5448 1044 5452
rect 1038 5447 1044 5448
rect 1174 5452 1180 5453
rect 1174 5448 1175 5452
rect 1179 5448 1180 5452
rect 1174 5447 1180 5448
rect 110 5446 116 5447
rect 112 5423 114 5446
rect 904 5423 906 5447
rect 1040 5423 1042 5447
rect 1176 5423 1178 5447
rect 111 5422 115 5423
rect 111 5417 115 5418
rect 719 5422 723 5423
rect 719 5417 723 5418
rect 855 5422 859 5423
rect 855 5417 859 5418
rect 903 5422 907 5423
rect 903 5417 907 5418
rect 991 5422 995 5423
rect 991 5417 995 5418
rect 1039 5422 1043 5423
rect 1039 5417 1043 5418
rect 1127 5422 1131 5423
rect 1127 5417 1131 5418
rect 1175 5422 1179 5423
rect 1175 5417 1179 5418
rect 1263 5422 1267 5423
rect 1263 5417 1267 5418
rect 112 5394 114 5417
rect 110 5393 116 5394
rect 720 5393 722 5417
rect 856 5393 858 5417
rect 992 5393 994 5417
rect 1128 5393 1130 5417
rect 1264 5393 1266 5417
rect 110 5389 111 5393
rect 115 5389 116 5393
rect 110 5388 116 5389
rect 718 5392 724 5393
rect 718 5388 719 5392
rect 723 5388 724 5392
rect 718 5387 724 5388
rect 854 5392 860 5393
rect 854 5388 855 5392
rect 859 5388 860 5392
rect 854 5387 860 5388
rect 990 5392 996 5393
rect 990 5388 991 5392
rect 995 5388 996 5392
rect 990 5387 996 5388
rect 1126 5392 1132 5393
rect 1126 5388 1127 5392
rect 1131 5388 1132 5392
rect 1126 5387 1132 5388
rect 1262 5392 1268 5393
rect 1262 5388 1263 5392
rect 1267 5388 1268 5392
rect 1262 5387 1268 5388
rect 690 5377 696 5378
rect 110 5376 116 5377
rect 110 5372 111 5376
rect 115 5372 116 5376
rect 690 5373 691 5377
rect 695 5373 696 5377
rect 690 5372 696 5373
rect 826 5377 832 5378
rect 826 5373 827 5377
rect 831 5373 832 5377
rect 826 5372 832 5373
rect 962 5377 968 5378
rect 962 5373 963 5377
rect 967 5373 968 5377
rect 962 5372 968 5373
rect 1098 5377 1104 5378
rect 1098 5373 1099 5377
rect 1103 5373 1104 5377
rect 1098 5372 1104 5373
rect 1234 5377 1240 5378
rect 1234 5373 1235 5377
rect 1239 5373 1240 5377
rect 1234 5372 1240 5373
rect 110 5371 116 5372
rect 112 5311 114 5371
rect 692 5311 694 5372
rect 810 5367 816 5368
rect 810 5363 811 5367
rect 815 5363 816 5367
rect 810 5362 816 5363
rect 111 5310 115 5311
rect 111 5305 115 5306
rect 691 5310 695 5311
rect 691 5305 695 5306
rect 723 5310 727 5311
rect 723 5305 727 5306
rect 112 5245 114 5305
rect 110 5244 116 5245
rect 724 5244 726 5305
rect 812 5284 814 5362
rect 828 5311 830 5372
rect 964 5311 966 5372
rect 1100 5311 1102 5372
rect 1186 5355 1192 5356
rect 1186 5351 1187 5355
rect 1191 5351 1192 5355
rect 1186 5350 1192 5351
rect 1188 5336 1190 5350
rect 1186 5335 1192 5336
rect 1186 5331 1187 5335
rect 1191 5331 1192 5335
rect 1186 5330 1192 5331
rect 1236 5311 1238 5372
rect 1272 5336 1274 5470
rect 1292 5468 1294 5529
rect 1418 5511 1424 5512
rect 1418 5507 1419 5511
rect 1423 5507 1424 5511
rect 1418 5506 1424 5507
rect 1420 5476 1422 5506
rect 1418 5475 1424 5476
rect 1418 5471 1419 5475
rect 1423 5471 1424 5475
rect 1418 5470 1424 5471
rect 1436 5468 1438 5529
rect 1558 5475 1564 5476
rect 1558 5471 1559 5475
rect 1563 5471 1564 5475
rect 1558 5470 1564 5471
rect 1290 5467 1296 5468
rect 1290 5463 1291 5467
rect 1295 5463 1296 5467
rect 1290 5462 1296 5463
rect 1434 5467 1440 5468
rect 1434 5463 1435 5467
rect 1439 5463 1440 5467
rect 1434 5462 1440 5463
rect 1318 5452 1324 5453
rect 1318 5448 1319 5452
rect 1323 5448 1324 5452
rect 1318 5447 1324 5448
rect 1462 5452 1468 5453
rect 1462 5448 1463 5452
rect 1467 5448 1468 5452
rect 1462 5447 1468 5448
rect 1320 5423 1322 5447
rect 1464 5423 1466 5447
rect 1319 5422 1323 5423
rect 1319 5417 1323 5418
rect 1399 5422 1403 5423
rect 1399 5417 1403 5418
rect 1463 5422 1467 5423
rect 1463 5417 1467 5418
rect 1535 5422 1539 5423
rect 1535 5417 1539 5418
rect 1400 5393 1402 5417
rect 1536 5393 1538 5417
rect 1398 5392 1404 5393
rect 1398 5388 1399 5392
rect 1403 5388 1404 5392
rect 1398 5387 1404 5388
rect 1534 5392 1540 5393
rect 1534 5388 1535 5392
rect 1539 5388 1540 5392
rect 1534 5387 1540 5388
rect 1370 5377 1376 5378
rect 1370 5373 1371 5377
rect 1375 5373 1376 5377
rect 1370 5372 1376 5373
rect 1506 5377 1512 5378
rect 1506 5373 1507 5377
rect 1511 5373 1512 5377
rect 1506 5372 1512 5373
rect 1270 5335 1276 5336
rect 1270 5331 1271 5335
rect 1275 5331 1276 5335
rect 1270 5330 1276 5331
rect 1372 5311 1374 5372
rect 1386 5367 1392 5368
rect 1386 5363 1387 5367
rect 1391 5363 1392 5367
rect 1386 5362 1392 5363
rect 1474 5367 1480 5368
rect 1474 5363 1475 5367
rect 1479 5363 1480 5367
rect 1474 5362 1480 5363
rect 1388 5336 1390 5362
rect 1386 5335 1392 5336
rect 1386 5331 1387 5335
rect 1391 5331 1392 5335
rect 1386 5330 1392 5331
rect 827 5310 831 5311
rect 827 5305 831 5306
rect 875 5310 879 5311
rect 875 5305 879 5306
rect 963 5310 967 5311
rect 963 5305 967 5306
rect 1027 5310 1031 5311
rect 1027 5305 1031 5306
rect 1099 5310 1103 5311
rect 1099 5305 1103 5306
rect 1187 5310 1191 5311
rect 1187 5305 1191 5306
rect 1235 5310 1239 5311
rect 1235 5305 1239 5306
rect 1355 5310 1359 5311
rect 1355 5305 1359 5306
rect 1371 5310 1375 5311
rect 1371 5305 1375 5306
rect 850 5287 856 5288
rect 810 5283 816 5284
rect 810 5279 811 5283
rect 815 5279 816 5283
rect 850 5283 851 5287
rect 855 5283 856 5287
rect 850 5282 856 5283
rect 810 5278 816 5279
rect 852 5252 854 5282
rect 850 5251 856 5252
rect 850 5247 851 5251
rect 855 5247 856 5251
rect 850 5246 856 5247
rect 876 5244 878 5305
rect 1002 5287 1008 5288
rect 1002 5283 1003 5287
rect 1007 5283 1008 5287
rect 1002 5282 1008 5283
rect 1004 5252 1006 5282
rect 1002 5251 1008 5252
rect 1002 5247 1003 5251
rect 1007 5247 1008 5251
rect 1002 5246 1008 5247
rect 1028 5244 1030 5305
rect 1154 5287 1160 5288
rect 1154 5283 1155 5287
rect 1159 5283 1160 5287
rect 1154 5282 1160 5283
rect 1156 5252 1158 5282
rect 1154 5251 1160 5252
rect 1154 5247 1155 5251
rect 1159 5247 1160 5251
rect 1154 5246 1160 5247
rect 1188 5244 1190 5305
rect 1258 5251 1264 5252
rect 1258 5247 1259 5251
rect 1263 5247 1264 5251
rect 1258 5246 1264 5247
rect 110 5240 111 5244
rect 115 5240 116 5244
rect 110 5239 116 5240
rect 722 5243 728 5244
rect 722 5239 723 5243
rect 727 5239 728 5243
rect 722 5238 728 5239
rect 874 5243 880 5244
rect 874 5239 875 5243
rect 879 5239 880 5243
rect 874 5238 880 5239
rect 1026 5243 1032 5244
rect 1026 5239 1027 5243
rect 1031 5239 1032 5243
rect 1026 5238 1032 5239
rect 1186 5243 1192 5244
rect 1186 5239 1187 5243
rect 1191 5239 1192 5243
rect 1186 5238 1192 5239
rect 750 5228 756 5229
rect 110 5227 116 5228
rect 110 5223 111 5227
rect 115 5223 116 5227
rect 750 5224 751 5228
rect 755 5224 756 5228
rect 750 5223 756 5224
rect 902 5228 908 5229
rect 902 5224 903 5228
rect 907 5224 908 5228
rect 902 5223 908 5224
rect 1054 5228 1060 5229
rect 1054 5224 1055 5228
rect 1059 5224 1060 5228
rect 1054 5223 1060 5224
rect 1214 5228 1220 5229
rect 1214 5224 1215 5228
rect 1219 5224 1220 5228
rect 1214 5223 1220 5224
rect 110 5222 116 5223
rect 112 5199 114 5222
rect 752 5199 754 5223
rect 904 5199 906 5223
rect 1056 5199 1058 5223
rect 1216 5199 1218 5223
rect 111 5198 115 5199
rect 111 5193 115 5194
rect 447 5198 451 5199
rect 447 5193 451 5194
rect 623 5198 627 5199
rect 623 5193 627 5194
rect 751 5198 755 5199
rect 751 5193 755 5194
rect 807 5198 811 5199
rect 807 5193 811 5194
rect 903 5198 907 5199
rect 903 5193 907 5194
rect 999 5198 1003 5199
rect 999 5193 1003 5194
rect 1055 5198 1059 5199
rect 1055 5193 1059 5194
rect 1199 5198 1203 5199
rect 1199 5193 1203 5194
rect 1215 5198 1219 5199
rect 1215 5193 1219 5194
rect 112 5170 114 5193
rect 110 5169 116 5170
rect 448 5169 450 5193
rect 624 5169 626 5193
rect 808 5169 810 5193
rect 1000 5169 1002 5193
rect 1200 5169 1202 5193
rect 110 5165 111 5169
rect 115 5165 116 5169
rect 110 5164 116 5165
rect 446 5168 452 5169
rect 446 5164 447 5168
rect 451 5164 452 5168
rect 446 5163 452 5164
rect 622 5168 628 5169
rect 622 5164 623 5168
rect 627 5164 628 5168
rect 622 5163 628 5164
rect 806 5168 812 5169
rect 806 5164 807 5168
rect 811 5164 812 5168
rect 806 5163 812 5164
rect 998 5168 1004 5169
rect 998 5164 999 5168
rect 1003 5164 1004 5168
rect 998 5163 1004 5164
rect 1198 5168 1204 5169
rect 1198 5164 1199 5168
rect 1203 5164 1204 5168
rect 1198 5163 1204 5164
rect 418 5153 424 5154
rect 110 5152 116 5153
rect 110 5148 111 5152
rect 115 5148 116 5152
rect 418 5149 419 5153
rect 423 5149 424 5153
rect 418 5148 424 5149
rect 594 5153 600 5154
rect 594 5149 595 5153
rect 599 5149 600 5153
rect 594 5148 600 5149
rect 778 5153 784 5154
rect 778 5149 779 5153
rect 783 5149 784 5153
rect 778 5148 784 5149
rect 970 5153 976 5154
rect 970 5149 971 5153
rect 975 5149 976 5153
rect 970 5148 976 5149
rect 1170 5153 1176 5154
rect 1170 5149 1171 5153
rect 1175 5149 1176 5153
rect 1170 5148 1176 5149
rect 110 5147 116 5148
rect 112 5079 114 5147
rect 274 5079 280 5080
rect 420 5079 422 5148
rect 596 5079 598 5148
rect 610 5143 616 5144
rect 610 5139 611 5143
rect 615 5139 616 5143
rect 610 5138 616 5139
rect 714 5143 720 5144
rect 714 5139 715 5143
rect 719 5139 720 5143
rect 714 5138 720 5139
rect 734 5143 740 5144
rect 734 5139 735 5143
rect 739 5139 740 5143
rect 734 5138 740 5139
rect 612 5112 614 5138
rect 610 5111 616 5112
rect 610 5107 611 5111
rect 615 5107 616 5111
rect 610 5106 616 5107
rect 111 5078 115 5079
rect 111 5073 115 5074
rect 155 5078 159 5079
rect 274 5075 275 5079
rect 279 5075 280 5079
rect 274 5074 280 5075
rect 379 5078 383 5079
rect 155 5073 159 5074
rect 112 5013 114 5073
rect 110 5012 116 5013
rect 156 5012 158 5073
rect 276 5056 278 5074
rect 379 5073 383 5074
rect 419 5078 423 5079
rect 419 5073 423 5074
rect 595 5078 599 5079
rect 595 5073 599 5074
rect 627 5078 631 5079
rect 627 5073 631 5074
rect 274 5055 280 5056
rect 274 5051 275 5055
rect 279 5051 280 5055
rect 274 5050 280 5051
rect 282 5055 288 5056
rect 282 5051 283 5055
rect 287 5051 288 5055
rect 282 5050 288 5051
rect 284 5020 286 5050
rect 282 5019 288 5020
rect 282 5015 283 5019
rect 287 5015 288 5019
rect 282 5014 288 5015
rect 380 5012 382 5073
rect 490 5019 496 5020
rect 490 5015 491 5019
rect 495 5015 496 5019
rect 490 5014 496 5015
rect 110 5008 111 5012
rect 115 5008 116 5012
rect 110 5007 116 5008
rect 154 5011 160 5012
rect 154 5007 155 5011
rect 159 5007 160 5011
rect 154 5006 160 5007
rect 378 5011 384 5012
rect 378 5007 379 5011
rect 383 5007 384 5011
rect 378 5006 384 5007
rect 182 4996 188 4997
rect 110 4995 116 4996
rect 110 4991 111 4995
rect 115 4991 116 4995
rect 182 4992 183 4996
rect 187 4992 188 4996
rect 182 4991 188 4992
rect 406 4996 412 4997
rect 406 4992 407 4996
rect 411 4992 412 4996
rect 406 4991 412 4992
rect 110 4990 116 4991
rect 112 4939 114 4990
rect 184 4939 186 4991
rect 408 4939 410 4991
rect 111 4938 115 4939
rect 111 4933 115 4934
rect 159 4938 163 4939
rect 159 4933 163 4934
rect 183 4938 187 4939
rect 183 4933 187 4934
rect 295 4938 299 4939
rect 295 4933 299 4934
rect 407 4938 411 4939
rect 407 4933 411 4934
rect 431 4938 435 4939
rect 431 4933 435 4934
rect 112 4910 114 4933
rect 110 4909 116 4910
rect 160 4909 162 4933
rect 296 4909 298 4933
rect 432 4909 434 4933
rect 110 4905 111 4909
rect 115 4905 116 4909
rect 110 4904 116 4905
rect 158 4908 164 4909
rect 158 4904 159 4908
rect 163 4904 164 4908
rect 158 4903 164 4904
rect 294 4908 300 4909
rect 294 4904 295 4908
rect 299 4904 300 4908
rect 294 4903 300 4904
rect 430 4908 436 4909
rect 430 4904 431 4908
rect 435 4904 436 4908
rect 430 4903 436 4904
rect 130 4893 136 4894
rect 110 4892 116 4893
rect 110 4888 111 4892
rect 115 4888 116 4892
rect 130 4889 131 4893
rect 135 4889 136 4893
rect 130 4888 136 4889
rect 266 4893 272 4894
rect 266 4889 267 4893
rect 271 4889 272 4893
rect 266 4888 272 4889
rect 402 4893 408 4894
rect 402 4889 403 4893
rect 407 4889 408 4893
rect 402 4888 408 4889
rect 110 4887 116 4888
rect 112 4815 114 4887
rect 132 4815 134 4888
rect 234 4883 240 4884
rect 234 4879 235 4883
rect 239 4879 240 4883
rect 234 4878 240 4879
rect 111 4814 115 4815
rect 111 4809 115 4810
rect 131 4814 135 4815
rect 131 4809 135 4810
rect 112 4749 114 4809
rect 110 4748 116 4749
rect 132 4748 134 4809
rect 236 4792 238 4878
rect 268 4815 270 4888
rect 354 4875 360 4876
rect 354 4871 355 4875
rect 359 4871 360 4875
rect 354 4870 360 4871
rect 356 4852 358 4870
rect 354 4851 360 4852
rect 354 4847 355 4851
rect 359 4847 360 4851
rect 354 4846 360 4847
rect 404 4815 406 4888
rect 492 4852 494 5014
rect 628 5012 630 5073
rect 716 5052 718 5138
rect 736 5096 738 5138
rect 734 5095 740 5096
rect 734 5091 735 5095
rect 739 5091 740 5095
rect 734 5090 740 5091
rect 780 5079 782 5148
rect 972 5079 974 5148
rect 1142 5143 1148 5144
rect 1142 5139 1143 5143
rect 1147 5139 1148 5143
rect 1142 5138 1148 5139
rect 1144 5112 1146 5138
rect 1142 5111 1148 5112
rect 1142 5107 1143 5111
rect 1147 5107 1148 5111
rect 1142 5106 1148 5107
rect 1172 5079 1174 5148
rect 1260 5112 1262 5246
rect 1356 5244 1358 5305
rect 1476 5288 1478 5362
rect 1508 5311 1510 5372
rect 1560 5336 1562 5470
rect 1580 5468 1582 5529
rect 1706 5511 1712 5512
rect 1706 5507 1707 5511
rect 1711 5507 1712 5511
rect 1706 5506 1712 5507
rect 1708 5476 1710 5506
rect 1706 5475 1712 5476
rect 1706 5471 1707 5475
rect 1711 5471 1712 5475
rect 1706 5470 1712 5471
rect 1724 5468 1726 5529
rect 1846 5527 1847 5531
rect 1851 5527 1852 5531
rect 2346 5533 2352 5534
rect 1935 5529 1939 5530
rect 1974 5532 1980 5533
rect 1846 5526 1852 5527
rect 1848 5476 1850 5526
rect 1846 5475 1852 5476
rect 1846 5471 1847 5475
rect 1851 5471 1852 5475
rect 1846 5470 1852 5471
rect 1936 5469 1938 5529
rect 1974 5528 1975 5532
rect 1979 5528 1980 5532
rect 2346 5529 2347 5533
rect 2351 5529 2352 5533
rect 2346 5528 2352 5529
rect 2578 5533 2584 5534
rect 2578 5529 2579 5533
rect 2583 5529 2584 5533
rect 2578 5528 2584 5529
rect 1974 5527 1980 5528
rect 1934 5468 1940 5469
rect 1578 5467 1584 5468
rect 1578 5463 1579 5467
rect 1583 5463 1584 5467
rect 1578 5462 1584 5463
rect 1722 5467 1728 5468
rect 1722 5463 1723 5467
rect 1727 5463 1728 5467
rect 1934 5464 1935 5468
rect 1939 5464 1940 5468
rect 1934 5463 1940 5464
rect 1976 5463 1978 5527
rect 2348 5463 2350 5528
rect 2434 5491 2440 5492
rect 2434 5487 2435 5491
rect 2439 5487 2440 5491
rect 2434 5486 2440 5487
rect 1722 5462 1728 5463
rect 1975 5462 1979 5463
rect 1975 5457 1979 5458
rect 2347 5462 2351 5463
rect 2347 5457 2351 5458
rect 1606 5452 1612 5453
rect 1606 5448 1607 5452
rect 1611 5448 1612 5452
rect 1606 5447 1612 5448
rect 1750 5452 1756 5453
rect 1750 5448 1751 5452
rect 1755 5448 1756 5452
rect 1750 5447 1756 5448
rect 1934 5451 1940 5452
rect 1934 5447 1935 5451
rect 1939 5447 1940 5451
rect 1608 5423 1610 5447
rect 1752 5423 1754 5447
rect 1934 5446 1940 5447
rect 1936 5423 1938 5446
rect 1607 5422 1611 5423
rect 1607 5417 1611 5418
rect 1671 5422 1675 5423
rect 1671 5417 1675 5418
rect 1751 5422 1755 5423
rect 1751 5417 1755 5418
rect 1807 5422 1811 5423
rect 1807 5417 1811 5418
rect 1935 5422 1939 5423
rect 1935 5417 1939 5418
rect 1672 5393 1674 5417
rect 1808 5393 1810 5417
rect 1936 5394 1938 5417
rect 1976 5397 1978 5457
rect 2418 5439 2424 5440
rect 2418 5435 2419 5439
rect 2423 5435 2424 5439
rect 2418 5434 2424 5435
rect 1974 5396 1980 5397
rect 1934 5393 1940 5394
rect 1670 5392 1676 5393
rect 1670 5388 1671 5392
rect 1675 5388 1676 5392
rect 1670 5387 1676 5388
rect 1806 5392 1812 5393
rect 1806 5388 1807 5392
rect 1811 5388 1812 5392
rect 1934 5389 1935 5393
rect 1939 5389 1940 5393
rect 1974 5392 1975 5396
rect 1979 5392 1980 5396
rect 1974 5391 1980 5392
rect 1934 5388 1940 5389
rect 1806 5387 1812 5388
rect 1974 5379 1980 5380
rect 1642 5377 1648 5378
rect 1642 5373 1643 5377
rect 1647 5373 1648 5377
rect 1642 5372 1648 5373
rect 1778 5377 1784 5378
rect 1778 5373 1779 5377
rect 1783 5373 1784 5377
rect 1778 5372 1784 5373
rect 1934 5376 1940 5377
rect 1934 5372 1935 5376
rect 1939 5372 1940 5376
rect 1974 5375 1975 5379
rect 1979 5375 1980 5379
rect 1974 5374 1980 5375
rect 1558 5335 1564 5336
rect 1558 5331 1559 5335
rect 1563 5331 1564 5335
rect 1558 5330 1564 5331
rect 1644 5311 1646 5372
rect 1658 5367 1664 5368
rect 1658 5363 1659 5367
rect 1663 5363 1664 5367
rect 1658 5362 1664 5363
rect 1660 5336 1662 5362
rect 1658 5335 1664 5336
rect 1658 5331 1659 5335
rect 1663 5331 1664 5335
rect 1658 5330 1664 5331
rect 1780 5311 1782 5372
rect 1934 5371 1940 5372
rect 1794 5367 1800 5368
rect 1794 5363 1795 5367
rect 1799 5363 1800 5367
rect 1794 5362 1800 5363
rect 1796 5336 1798 5362
rect 1794 5335 1800 5336
rect 1794 5331 1795 5335
rect 1799 5331 1800 5335
rect 1794 5330 1800 5331
rect 1936 5311 1938 5371
rect 1976 5351 1978 5374
rect 1975 5350 1979 5351
rect 1975 5345 1979 5346
rect 2319 5350 2323 5351
rect 2319 5345 2323 5346
rect 1976 5322 1978 5345
rect 1974 5321 1980 5322
rect 2320 5321 2322 5345
rect 1974 5317 1975 5321
rect 1979 5317 1980 5321
rect 1974 5316 1980 5317
rect 2318 5320 2324 5321
rect 2318 5316 2319 5320
rect 2323 5316 2324 5320
rect 2318 5315 2324 5316
rect 1507 5310 1511 5311
rect 1507 5305 1511 5306
rect 1523 5310 1527 5311
rect 1523 5305 1527 5306
rect 1643 5310 1647 5311
rect 1643 5305 1647 5306
rect 1779 5310 1783 5311
rect 1779 5305 1783 5306
rect 1935 5310 1939 5311
rect 1935 5305 1939 5306
rect 2290 5305 2296 5306
rect 1474 5287 1480 5288
rect 1474 5283 1475 5287
rect 1479 5283 1480 5287
rect 1474 5282 1480 5283
rect 1524 5244 1526 5305
rect 1646 5251 1652 5252
rect 1646 5247 1647 5251
rect 1651 5247 1652 5251
rect 1646 5246 1652 5247
rect 1354 5243 1360 5244
rect 1354 5239 1355 5243
rect 1359 5239 1360 5243
rect 1354 5238 1360 5239
rect 1522 5243 1528 5244
rect 1522 5239 1523 5243
rect 1527 5239 1528 5243
rect 1522 5238 1528 5239
rect 1382 5228 1388 5229
rect 1382 5224 1383 5228
rect 1387 5224 1388 5228
rect 1382 5223 1388 5224
rect 1550 5228 1556 5229
rect 1550 5224 1551 5228
rect 1555 5224 1556 5228
rect 1550 5223 1556 5224
rect 1384 5199 1386 5223
rect 1552 5199 1554 5223
rect 1383 5198 1387 5199
rect 1383 5193 1387 5194
rect 1399 5198 1403 5199
rect 1399 5193 1403 5194
rect 1551 5198 1555 5199
rect 1551 5193 1555 5194
rect 1607 5198 1611 5199
rect 1607 5193 1611 5194
rect 1400 5169 1402 5193
rect 1608 5169 1610 5193
rect 1398 5168 1404 5169
rect 1398 5164 1399 5168
rect 1403 5164 1404 5168
rect 1398 5163 1404 5164
rect 1606 5168 1612 5169
rect 1606 5164 1607 5168
rect 1611 5164 1612 5168
rect 1606 5163 1612 5164
rect 1370 5153 1376 5154
rect 1370 5149 1371 5153
rect 1375 5149 1376 5153
rect 1370 5148 1376 5149
rect 1578 5153 1584 5154
rect 1578 5149 1579 5153
rect 1583 5149 1584 5153
rect 1578 5148 1584 5149
rect 1258 5111 1264 5112
rect 1258 5107 1259 5111
rect 1263 5107 1264 5111
rect 1258 5106 1264 5107
rect 1318 5079 1324 5080
rect 1372 5079 1374 5148
rect 1490 5143 1496 5144
rect 1490 5139 1491 5143
rect 1495 5139 1496 5143
rect 1490 5138 1496 5139
rect 1458 5135 1464 5136
rect 1458 5131 1459 5135
rect 1463 5131 1464 5135
rect 1458 5130 1464 5131
rect 1460 5112 1462 5130
rect 1458 5111 1464 5112
rect 1458 5107 1459 5111
rect 1463 5107 1464 5111
rect 1458 5106 1464 5107
rect 779 5078 783 5079
rect 779 5073 783 5074
rect 899 5078 903 5079
rect 899 5073 903 5074
rect 971 5078 975 5079
rect 971 5073 975 5074
rect 1171 5078 1175 5079
rect 1171 5073 1175 5074
rect 1195 5078 1199 5079
rect 1318 5075 1319 5079
rect 1323 5075 1324 5079
rect 1318 5074 1324 5075
rect 1371 5078 1375 5079
rect 1195 5073 1199 5074
rect 754 5055 760 5056
rect 714 5051 720 5052
rect 714 5047 715 5051
rect 719 5047 720 5051
rect 754 5051 755 5055
rect 759 5051 760 5055
rect 754 5050 760 5051
rect 714 5046 720 5047
rect 756 5020 758 5050
rect 754 5019 760 5020
rect 754 5015 755 5019
rect 759 5015 760 5019
rect 754 5014 760 5015
rect 900 5012 902 5073
rect 1118 5055 1124 5056
rect 1118 5051 1119 5055
rect 1123 5051 1124 5055
rect 1118 5050 1124 5051
rect 1120 5020 1122 5050
rect 1118 5019 1124 5020
rect 1118 5015 1119 5019
rect 1123 5015 1124 5019
rect 1118 5014 1124 5015
rect 1196 5012 1198 5073
rect 1320 5020 1322 5074
rect 1371 5073 1375 5074
rect 1492 5056 1494 5138
rect 1580 5079 1582 5148
rect 1648 5112 1650 5246
rect 1936 5245 1938 5305
rect 1974 5304 1980 5305
rect 1974 5300 1975 5304
rect 1979 5300 1980 5304
rect 2290 5301 2291 5305
rect 2295 5301 2296 5305
rect 2290 5300 2296 5301
rect 1974 5299 1980 5300
rect 1934 5244 1940 5245
rect 1934 5240 1935 5244
rect 1939 5240 1940 5244
rect 1934 5239 1940 5240
rect 1976 5235 1978 5299
rect 2292 5235 2294 5300
rect 2420 5296 2422 5434
rect 2436 5404 2438 5486
rect 2580 5463 2582 5528
rect 2652 5524 2654 5658
rect 2748 5624 2750 5685
rect 2874 5667 2880 5668
rect 2874 5663 2875 5667
rect 2879 5663 2880 5667
rect 2874 5662 2880 5663
rect 2876 5632 2878 5662
rect 2874 5631 2880 5632
rect 2874 5627 2875 5631
rect 2879 5627 2880 5631
rect 2874 5626 2880 5627
rect 2932 5624 2934 5685
rect 3058 5667 3064 5668
rect 3058 5663 3059 5667
rect 3063 5663 3064 5667
rect 3058 5662 3064 5663
rect 3060 5632 3062 5662
rect 3066 5651 3072 5652
rect 3066 5647 3067 5651
rect 3071 5647 3072 5651
rect 3066 5646 3072 5647
rect 3058 5631 3064 5632
rect 3058 5627 3059 5631
rect 3063 5627 3064 5631
rect 3058 5626 3064 5627
rect 2746 5623 2752 5624
rect 2746 5619 2747 5623
rect 2751 5619 2752 5623
rect 2746 5618 2752 5619
rect 2930 5623 2936 5624
rect 2930 5619 2931 5623
rect 2935 5619 2936 5623
rect 2930 5618 2936 5619
rect 2774 5608 2780 5609
rect 2774 5604 2775 5608
rect 2779 5604 2780 5608
rect 2774 5603 2780 5604
rect 2958 5608 2964 5609
rect 2958 5604 2959 5608
rect 2963 5604 2964 5608
rect 2958 5603 2964 5604
rect 2776 5579 2778 5603
rect 2960 5579 2962 5603
rect 2775 5578 2779 5579
rect 2775 5573 2779 5574
rect 2831 5578 2835 5579
rect 2831 5573 2835 5574
rect 2959 5578 2963 5579
rect 2959 5573 2963 5574
rect 3047 5578 3051 5579
rect 3047 5573 3051 5574
rect 2832 5549 2834 5573
rect 3048 5549 3050 5573
rect 2830 5548 2836 5549
rect 2830 5544 2831 5548
rect 2835 5544 2836 5548
rect 2830 5543 2836 5544
rect 3046 5548 3052 5549
rect 3046 5544 3047 5548
rect 3051 5544 3052 5548
rect 3046 5543 3052 5544
rect 2802 5533 2808 5534
rect 2802 5529 2803 5533
rect 2807 5529 2808 5533
rect 2802 5528 2808 5529
rect 3018 5533 3024 5534
rect 3018 5529 3019 5533
rect 3023 5529 3024 5533
rect 3018 5528 3024 5529
rect 2594 5523 2600 5524
rect 2594 5519 2595 5523
rect 2599 5519 2600 5523
rect 2594 5518 2600 5519
rect 2650 5523 2656 5524
rect 2650 5519 2651 5523
rect 2655 5519 2656 5523
rect 2650 5518 2656 5519
rect 2596 5492 2598 5518
rect 2594 5491 2600 5492
rect 2594 5487 2595 5491
rect 2599 5487 2600 5491
rect 2594 5486 2600 5487
rect 2804 5463 2806 5528
rect 2822 5491 2828 5492
rect 2822 5487 2823 5491
rect 2827 5487 2828 5491
rect 2822 5486 2828 5487
rect 2451 5462 2455 5463
rect 2451 5457 2455 5458
rect 2579 5462 2583 5463
rect 2579 5457 2583 5458
rect 2699 5462 2703 5463
rect 2699 5457 2703 5458
rect 2803 5462 2807 5463
rect 2803 5457 2807 5458
rect 2434 5403 2440 5404
rect 2434 5399 2435 5403
rect 2439 5399 2440 5403
rect 2434 5398 2440 5399
rect 2452 5396 2454 5457
rect 2700 5396 2702 5457
rect 2824 5404 2826 5486
rect 3020 5463 3022 5528
rect 3068 5524 3070 5646
rect 3108 5624 3110 5685
rect 3234 5667 3240 5668
rect 3234 5663 3235 5667
rect 3239 5663 3240 5667
rect 3234 5662 3240 5663
rect 3236 5632 3238 5662
rect 3234 5631 3240 5632
rect 3234 5627 3235 5631
rect 3239 5627 3240 5631
rect 3234 5626 3240 5627
rect 3276 5624 3278 5685
rect 3402 5667 3408 5668
rect 3402 5663 3403 5667
rect 3407 5663 3408 5667
rect 3402 5662 3408 5663
rect 3404 5632 3406 5662
rect 3402 5631 3408 5632
rect 3402 5627 3403 5631
rect 3407 5627 3408 5631
rect 3402 5626 3408 5627
rect 3444 5624 3446 5685
rect 3570 5667 3576 5668
rect 3570 5663 3571 5667
rect 3575 5663 3576 5667
rect 3570 5662 3576 5663
rect 3572 5632 3574 5662
rect 3570 5631 3576 5632
rect 3570 5627 3571 5631
rect 3575 5627 3576 5631
rect 3570 5626 3576 5627
rect 3620 5624 3622 5685
rect 3738 5631 3744 5632
rect 3738 5627 3739 5631
rect 3743 5627 3744 5631
rect 3738 5626 3744 5627
rect 3106 5623 3112 5624
rect 3106 5619 3107 5623
rect 3111 5619 3112 5623
rect 3106 5618 3112 5619
rect 3274 5623 3280 5624
rect 3274 5619 3275 5623
rect 3279 5619 3280 5623
rect 3274 5618 3280 5619
rect 3442 5623 3448 5624
rect 3442 5619 3443 5623
rect 3447 5619 3448 5623
rect 3442 5618 3448 5619
rect 3618 5623 3624 5624
rect 3618 5619 3619 5623
rect 3623 5619 3624 5623
rect 3618 5618 3624 5619
rect 3134 5608 3140 5609
rect 3134 5604 3135 5608
rect 3139 5604 3140 5608
rect 3134 5603 3140 5604
rect 3302 5608 3308 5609
rect 3302 5604 3303 5608
rect 3307 5604 3308 5608
rect 3302 5603 3308 5604
rect 3470 5608 3476 5609
rect 3470 5604 3471 5608
rect 3475 5604 3476 5608
rect 3470 5603 3476 5604
rect 3646 5608 3652 5609
rect 3646 5604 3647 5608
rect 3651 5604 3652 5608
rect 3646 5603 3652 5604
rect 3136 5579 3138 5603
rect 3304 5579 3306 5603
rect 3472 5579 3474 5603
rect 3648 5579 3650 5603
rect 3135 5578 3139 5579
rect 3135 5573 3139 5574
rect 3263 5578 3267 5579
rect 3263 5573 3267 5574
rect 3303 5578 3307 5579
rect 3303 5573 3307 5574
rect 3471 5578 3475 5579
rect 3471 5573 3475 5574
rect 3479 5578 3483 5579
rect 3479 5573 3483 5574
rect 3647 5578 3651 5579
rect 3647 5573 3651 5574
rect 3679 5578 3683 5579
rect 3679 5573 3683 5574
rect 3264 5549 3266 5573
rect 3480 5549 3482 5573
rect 3680 5549 3682 5573
rect 3262 5548 3268 5549
rect 3262 5544 3263 5548
rect 3267 5544 3268 5548
rect 3262 5543 3268 5544
rect 3478 5548 3484 5549
rect 3478 5544 3479 5548
rect 3483 5544 3484 5548
rect 3478 5543 3484 5544
rect 3678 5548 3684 5549
rect 3678 5544 3679 5548
rect 3683 5544 3684 5548
rect 3678 5543 3684 5544
rect 3234 5533 3240 5534
rect 3234 5529 3235 5533
rect 3239 5529 3240 5533
rect 3234 5528 3240 5529
rect 3450 5533 3456 5534
rect 3450 5529 3451 5533
rect 3455 5529 3456 5533
rect 3450 5528 3456 5529
rect 3650 5533 3656 5534
rect 3650 5529 3651 5533
rect 3655 5529 3656 5533
rect 3650 5528 3656 5529
rect 3034 5523 3040 5524
rect 3034 5519 3035 5523
rect 3039 5519 3040 5523
rect 3034 5518 3040 5519
rect 3066 5523 3072 5524
rect 3066 5519 3067 5523
rect 3071 5519 3072 5523
rect 3066 5518 3072 5519
rect 3036 5492 3038 5518
rect 3034 5491 3040 5492
rect 3034 5487 3035 5491
rect 3039 5487 3040 5491
rect 3034 5486 3040 5487
rect 3236 5463 3238 5528
rect 3322 5515 3328 5516
rect 3322 5511 3323 5515
rect 3327 5511 3328 5515
rect 3322 5510 3328 5511
rect 3324 5492 3326 5510
rect 3322 5491 3328 5492
rect 3322 5487 3323 5491
rect 3327 5487 3328 5491
rect 3322 5486 3328 5487
rect 3452 5463 3454 5528
rect 3466 5523 3472 5524
rect 3466 5519 3467 5523
rect 3471 5519 3472 5523
rect 3466 5518 3472 5519
rect 3578 5523 3584 5524
rect 3578 5519 3579 5523
rect 3583 5519 3584 5523
rect 3578 5518 3584 5519
rect 3468 5492 3470 5518
rect 3466 5491 3472 5492
rect 3466 5487 3467 5491
rect 3471 5487 3472 5491
rect 3466 5486 3472 5487
rect 2947 5462 2951 5463
rect 2947 5457 2951 5458
rect 3019 5462 3023 5463
rect 3019 5457 3023 5458
rect 3187 5462 3191 5463
rect 3187 5457 3191 5458
rect 3235 5462 3239 5463
rect 3235 5457 3239 5458
rect 3427 5462 3431 5463
rect 3427 5457 3431 5458
rect 3451 5462 3455 5463
rect 3451 5457 3455 5458
rect 2894 5439 2900 5440
rect 2894 5435 2895 5439
rect 2899 5435 2900 5439
rect 2894 5434 2900 5435
rect 2896 5404 2898 5434
rect 2822 5403 2828 5404
rect 2822 5399 2823 5403
rect 2827 5399 2828 5403
rect 2822 5398 2828 5399
rect 2894 5403 2900 5404
rect 2894 5399 2895 5403
rect 2899 5399 2900 5403
rect 2894 5398 2900 5399
rect 2948 5396 2950 5457
rect 3034 5435 3040 5436
rect 3034 5431 3035 5435
rect 3039 5431 3040 5435
rect 3034 5430 3040 5431
rect 2450 5395 2456 5396
rect 2450 5391 2451 5395
rect 2455 5391 2456 5395
rect 2450 5390 2456 5391
rect 2698 5395 2704 5396
rect 2698 5391 2699 5395
rect 2703 5391 2704 5395
rect 2698 5390 2704 5391
rect 2946 5395 2952 5396
rect 2946 5391 2947 5395
rect 2951 5391 2952 5395
rect 2946 5390 2952 5391
rect 2478 5380 2484 5381
rect 2478 5376 2479 5380
rect 2483 5376 2484 5380
rect 2478 5375 2484 5376
rect 2726 5380 2732 5381
rect 2726 5376 2727 5380
rect 2731 5376 2732 5380
rect 2726 5375 2732 5376
rect 2974 5380 2980 5381
rect 2974 5376 2975 5380
rect 2979 5376 2980 5380
rect 2974 5375 2980 5376
rect 2480 5351 2482 5375
rect 2728 5351 2730 5375
rect 2976 5351 2978 5375
rect 2479 5350 2483 5351
rect 2479 5345 2483 5346
rect 2519 5350 2523 5351
rect 2519 5345 2523 5346
rect 2719 5350 2723 5351
rect 2719 5345 2723 5346
rect 2727 5350 2731 5351
rect 2727 5345 2731 5346
rect 2919 5350 2923 5351
rect 2919 5345 2923 5346
rect 2975 5350 2979 5351
rect 2975 5345 2979 5346
rect 2520 5321 2522 5345
rect 2720 5321 2722 5345
rect 2920 5321 2922 5345
rect 2518 5320 2524 5321
rect 2518 5316 2519 5320
rect 2523 5316 2524 5320
rect 2518 5315 2524 5316
rect 2718 5320 2724 5321
rect 2718 5316 2719 5320
rect 2723 5316 2724 5320
rect 2718 5315 2724 5316
rect 2918 5320 2924 5321
rect 2918 5316 2919 5320
rect 2923 5316 2924 5320
rect 2918 5315 2924 5316
rect 2490 5305 2496 5306
rect 2490 5301 2491 5305
rect 2495 5301 2496 5305
rect 2490 5300 2496 5301
rect 2690 5305 2696 5306
rect 2690 5301 2691 5305
rect 2695 5301 2696 5305
rect 2690 5300 2696 5301
rect 2890 5305 2896 5306
rect 2890 5301 2891 5305
rect 2895 5301 2896 5305
rect 2890 5300 2896 5301
rect 2418 5295 2424 5296
rect 2418 5291 2419 5295
rect 2423 5291 2424 5295
rect 2418 5290 2424 5291
rect 2378 5287 2384 5288
rect 2378 5283 2379 5287
rect 2383 5283 2384 5287
rect 2378 5282 2384 5283
rect 2380 5264 2382 5282
rect 2378 5263 2384 5264
rect 2378 5259 2379 5263
rect 2383 5259 2384 5263
rect 2378 5258 2384 5259
rect 2492 5235 2494 5300
rect 2578 5263 2584 5264
rect 2578 5259 2579 5263
rect 2583 5259 2584 5263
rect 2578 5258 2584 5259
rect 1975 5234 1979 5235
rect 1975 5229 1979 5230
rect 2275 5234 2279 5235
rect 2275 5229 2279 5230
rect 2291 5234 2295 5235
rect 2291 5229 2295 5230
rect 2475 5234 2479 5235
rect 2475 5229 2479 5230
rect 2491 5234 2495 5235
rect 2491 5229 2495 5230
rect 1934 5227 1940 5228
rect 1934 5223 1935 5227
rect 1939 5223 1940 5227
rect 1934 5222 1940 5223
rect 1936 5199 1938 5222
rect 1815 5198 1819 5199
rect 1815 5193 1819 5194
rect 1935 5198 1939 5199
rect 1935 5193 1939 5194
rect 1816 5169 1818 5193
rect 1936 5170 1938 5193
rect 1934 5169 1940 5170
rect 1976 5169 1978 5229
rect 1814 5168 1820 5169
rect 1814 5164 1815 5168
rect 1819 5164 1820 5168
rect 1934 5165 1935 5169
rect 1939 5165 1940 5169
rect 1934 5164 1940 5165
rect 1974 5168 1980 5169
rect 2276 5168 2278 5229
rect 2402 5211 2408 5212
rect 2362 5207 2368 5208
rect 2362 5203 2363 5207
rect 2367 5203 2368 5207
rect 2402 5207 2403 5211
rect 2407 5207 2408 5211
rect 2402 5206 2408 5207
rect 2362 5202 2368 5203
rect 1974 5164 1975 5168
rect 1979 5164 1980 5168
rect 1814 5163 1820 5164
rect 1974 5163 1980 5164
rect 2274 5167 2280 5168
rect 2274 5163 2275 5167
rect 2279 5163 2280 5167
rect 2274 5162 2280 5163
rect 1786 5153 1792 5154
rect 1786 5149 1787 5153
rect 1791 5149 1792 5153
rect 1786 5148 1792 5149
rect 1934 5152 1940 5153
rect 2302 5152 2308 5153
rect 1934 5148 1935 5152
rect 1939 5148 1940 5152
rect 1646 5111 1652 5112
rect 1646 5107 1647 5111
rect 1651 5107 1652 5111
rect 1646 5106 1652 5107
rect 1788 5079 1790 5148
rect 1934 5147 1940 5148
rect 1974 5151 1980 5152
rect 1974 5147 1975 5151
rect 1979 5147 1980 5151
rect 2302 5148 2303 5152
rect 2307 5148 2308 5152
rect 2302 5147 2308 5148
rect 1802 5143 1808 5144
rect 1802 5139 1803 5143
rect 1807 5139 1808 5143
rect 1802 5138 1808 5139
rect 1804 5112 1806 5138
rect 1802 5111 1808 5112
rect 1802 5107 1803 5111
rect 1807 5107 1808 5111
rect 1802 5106 1808 5107
rect 1936 5079 1938 5147
rect 1974 5146 1980 5147
rect 1976 5107 1978 5146
rect 2304 5107 2306 5147
rect 2364 5115 2366 5202
rect 2404 5176 2406 5206
rect 2402 5175 2408 5176
rect 2402 5171 2403 5175
rect 2407 5171 2408 5175
rect 2402 5170 2408 5171
rect 2476 5168 2478 5229
rect 2580 5176 2582 5258
rect 2692 5235 2694 5300
rect 2706 5295 2712 5296
rect 2706 5291 2707 5295
rect 2711 5291 2712 5295
rect 2706 5290 2712 5291
rect 2708 5264 2710 5290
rect 2706 5263 2712 5264
rect 2706 5259 2707 5263
rect 2711 5259 2712 5263
rect 2706 5258 2712 5259
rect 2892 5235 2894 5300
rect 3036 5296 3038 5430
rect 3188 5396 3190 5457
rect 3314 5439 3320 5440
rect 3274 5435 3280 5436
rect 3274 5431 3275 5435
rect 3279 5431 3280 5435
rect 3314 5435 3315 5439
rect 3319 5435 3320 5439
rect 3314 5434 3320 5435
rect 3274 5430 3280 5431
rect 3276 5416 3278 5430
rect 3274 5415 3280 5416
rect 3274 5411 3275 5415
rect 3279 5411 3280 5415
rect 3274 5410 3280 5411
rect 3316 5404 3318 5434
rect 3314 5403 3320 5404
rect 3314 5399 3315 5403
rect 3319 5399 3320 5403
rect 3314 5398 3320 5399
rect 3428 5396 3430 5457
rect 3580 5440 3582 5518
rect 3652 5463 3654 5528
rect 3740 5492 3742 5626
rect 3800 5625 3802 5685
rect 3840 5629 3842 5689
rect 3838 5628 3844 5629
rect 4468 5628 4470 5689
rect 4554 5667 4560 5668
rect 4554 5663 4555 5667
rect 4559 5663 4560 5667
rect 4554 5662 4560 5663
rect 3798 5624 3804 5625
rect 3798 5620 3799 5624
rect 3803 5620 3804 5624
rect 3838 5624 3839 5628
rect 3843 5624 3844 5628
rect 3838 5623 3844 5624
rect 4466 5627 4472 5628
rect 4466 5623 4467 5627
rect 4471 5623 4472 5627
rect 4466 5622 4472 5623
rect 3798 5619 3804 5620
rect 4494 5612 4500 5613
rect 3838 5611 3844 5612
rect 3798 5607 3804 5608
rect 3798 5603 3799 5607
rect 3803 5603 3804 5607
rect 3838 5607 3839 5611
rect 3843 5607 3844 5611
rect 4494 5608 4495 5612
rect 4499 5608 4500 5612
rect 4494 5607 4500 5608
rect 3838 5606 3844 5607
rect 3798 5602 3804 5603
rect 3800 5579 3802 5602
rect 3840 5583 3842 5606
rect 4496 5583 4498 5607
rect 3839 5582 3843 5583
rect 3799 5578 3803 5579
rect 3839 5577 3843 5578
rect 4431 5582 4435 5583
rect 4431 5577 4435 5578
rect 4495 5582 4499 5583
rect 4495 5577 4499 5578
rect 3799 5573 3803 5574
rect 3800 5550 3802 5573
rect 3840 5554 3842 5577
rect 3838 5553 3844 5554
rect 4432 5553 4434 5577
rect 3798 5549 3804 5550
rect 3798 5545 3799 5549
rect 3803 5545 3804 5549
rect 3838 5549 3839 5553
rect 3843 5549 3844 5553
rect 3838 5548 3844 5549
rect 4430 5552 4436 5553
rect 4430 5548 4431 5552
rect 4435 5548 4436 5552
rect 4430 5547 4436 5548
rect 3798 5544 3804 5545
rect 4402 5537 4408 5538
rect 3838 5536 3844 5537
rect 3798 5532 3804 5533
rect 3798 5528 3799 5532
rect 3803 5528 3804 5532
rect 3838 5532 3839 5536
rect 3843 5532 3844 5536
rect 4402 5533 4403 5537
rect 4407 5533 4408 5537
rect 4402 5532 4408 5533
rect 4538 5537 4544 5538
rect 4538 5533 4539 5537
rect 4543 5533 4544 5537
rect 4538 5532 4544 5533
rect 3838 5531 3844 5532
rect 3798 5527 3804 5528
rect 3738 5491 3744 5492
rect 3738 5487 3739 5491
rect 3743 5487 3744 5491
rect 3738 5486 3744 5487
rect 3800 5463 3802 5527
rect 3840 5471 3842 5531
rect 4404 5471 4406 5532
rect 4490 5519 4496 5520
rect 4490 5515 4491 5519
rect 4495 5515 4496 5519
rect 4490 5514 4496 5515
rect 4492 5496 4494 5514
rect 4490 5495 4496 5496
rect 4490 5491 4491 5495
rect 4495 5491 4496 5495
rect 4490 5490 4496 5491
rect 4540 5471 4542 5532
rect 4556 5528 4558 5662
rect 4604 5628 4606 5689
rect 4740 5628 4742 5689
rect 4876 5628 4878 5689
rect 4910 5635 4916 5636
rect 4910 5631 4911 5635
rect 4915 5631 4916 5635
rect 4910 5630 4916 5631
rect 4602 5627 4608 5628
rect 4602 5623 4603 5627
rect 4607 5623 4608 5627
rect 4602 5622 4608 5623
rect 4738 5627 4744 5628
rect 4738 5623 4739 5627
rect 4743 5623 4744 5627
rect 4738 5622 4744 5623
rect 4874 5627 4880 5628
rect 4874 5623 4875 5627
rect 4879 5623 4880 5627
rect 4874 5622 4880 5623
rect 4630 5612 4636 5613
rect 4630 5608 4631 5612
rect 4635 5608 4636 5612
rect 4630 5607 4636 5608
rect 4766 5612 4772 5613
rect 4766 5608 4767 5612
rect 4771 5608 4772 5612
rect 4766 5607 4772 5608
rect 4902 5612 4908 5613
rect 4902 5608 4903 5612
rect 4907 5608 4908 5612
rect 4902 5607 4908 5608
rect 4632 5583 4634 5607
rect 4768 5583 4770 5607
rect 4904 5583 4906 5607
rect 4567 5582 4571 5583
rect 4567 5577 4571 5578
rect 4631 5582 4635 5583
rect 4631 5577 4635 5578
rect 4703 5582 4707 5583
rect 4703 5577 4707 5578
rect 4767 5582 4771 5583
rect 4767 5577 4771 5578
rect 4839 5582 4843 5583
rect 4839 5577 4843 5578
rect 4903 5582 4907 5583
rect 4903 5577 4907 5578
rect 4568 5553 4570 5577
rect 4704 5553 4706 5577
rect 4840 5553 4842 5577
rect 4566 5552 4572 5553
rect 4566 5548 4567 5552
rect 4571 5548 4572 5552
rect 4566 5547 4572 5548
rect 4702 5552 4708 5553
rect 4702 5548 4703 5552
rect 4707 5548 4708 5552
rect 4702 5547 4708 5548
rect 4838 5552 4844 5553
rect 4838 5548 4839 5552
rect 4843 5548 4844 5552
rect 4838 5547 4844 5548
rect 4674 5537 4680 5538
rect 4674 5533 4675 5537
rect 4679 5533 4680 5537
rect 4674 5532 4680 5533
rect 4810 5537 4816 5538
rect 4810 5533 4811 5537
rect 4815 5533 4816 5537
rect 4810 5532 4816 5533
rect 4554 5527 4560 5528
rect 4554 5523 4555 5527
rect 4559 5523 4560 5527
rect 4554 5522 4560 5523
rect 4626 5495 4632 5496
rect 4626 5491 4627 5495
rect 4631 5491 4632 5495
rect 4626 5490 4632 5491
rect 3839 5470 3843 5471
rect 3839 5465 3843 5466
rect 4403 5470 4407 5471
rect 4403 5465 4407 5466
rect 4427 5470 4431 5471
rect 4427 5465 4431 5466
rect 4539 5470 4543 5471
rect 4539 5465 4543 5466
rect 4587 5470 4591 5471
rect 4587 5465 4591 5466
rect 3651 5462 3655 5463
rect 3651 5457 3655 5458
rect 3799 5462 3803 5463
rect 3799 5457 3803 5458
rect 3578 5439 3584 5440
rect 3578 5435 3579 5439
rect 3583 5435 3584 5439
rect 3578 5434 3584 5435
rect 3550 5403 3556 5404
rect 3550 5399 3551 5403
rect 3555 5399 3556 5403
rect 3550 5398 3556 5399
rect 3186 5395 3192 5396
rect 3186 5391 3187 5395
rect 3191 5391 3192 5395
rect 3186 5390 3192 5391
rect 3426 5395 3432 5396
rect 3426 5391 3427 5395
rect 3431 5391 3432 5395
rect 3426 5390 3432 5391
rect 3214 5380 3220 5381
rect 3214 5376 3215 5380
rect 3219 5376 3220 5380
rect 3214 5375 3220 5376
rect 3454 5380 3460 5381
rect 3454 5376 3455 5380
rect 3459 5376 3460 5380
rect 3454 5375 3460 5376
rect 3216 5351 3218 5375
rect 3456 5351 3458 5375
rect 3119 5350 3123 5351
rect 3119 5345 3123 5346
rect 3215 5350 3219 5351
rect 3215 5345 3219 5346
rect 3327 5350 3331 5351
rect 3327 5345 3331 5346
rect 3455 5350 3459 5351
rect 3455 5345 3459 5346
rect 3535 5350 3539 5351
rect 3535 5345 3539 5346
rect 3120 5321 3122 5345
rect 3328 5321 3330 5345
rect 3536 5321 3538 5345
rect 3118 5320 3124 5321
rect 3118 5316 3119 5320
rect 3123 5316 3124 5320
rect 3118 5315 3124 5316
rect 3326 5320 3332 5321
rect 3326 5316 3327 5320
rect 3331 5316 3332 5320
rect 3326 5315 3332 5316
rect 3534 5320 3540 5321
rect 3534 5316 3535 5320
rect 3539 5316 3540 5320
rect 3534 5315 3540 5316
rect 3090 5305 3096 5306
rect 3090 5301 3091 5305
rect 3095 5301 3096 5305
rect 3090 5300 3096 5301
rect 3298 5305 3304 5306
rect 3298 5301 3299 5305
rect 3303 5301 3304 5305
rect 3298 5300 3304 5301
rect 3506 5305 3512 5306
rect 3506 5301 3507 5305
rect 3511 5301 3512 5305
rect 3506 5300 3512 5301
rect 3034 5295 3040 5296
rect 3034 5291 3035 5295
rect 3039 5291 3040 5295
rect 3034 5290 3040 5291
rect 2978 5263 2984 5264
rect 2978 5259 2979 5263
rect 2983 5259 2984 5263
rect 2978 5258 2984 5259
rect 2683 5234 2687 5235
rect 2683 5229 2687 5230
rect 2691 5234 2695 5235
rect 2691 5229 2695 5230
rect 2891 5234 2895 5235
rect 2891 5229 2895 5230
rect 2578 5175 2584 5176
rect 2578 5171 2579 5175
rect 2583 5171 2584 5175
rect 2578 5170 2584 5171
rect 2684 5168 2686 5229
rect 2810 5211 2816 5212
rect 2770 5207 2776 5208
rect 2770 5203 2771 5207
rect 2775 5203 2776 5207
rect 2810 5207 2811 5211
rect 2815 5207 2816 5211
rect 2810 5206 2816 5207
rect 2770 5202 2776 5203
rect 2474 5167 2480 5168
rect 2474 5163 2475 5167
rect 2479 5163 2480 5167
rect 2474 5162 2480 5163
rect 2682 5167 2688 5168
rect 2682 5163 2683 5167
rect 2687 5163 2688 5167
rect 2682 5162 2688 5163
rect 2502 5152 2508 5153
rect 2502 5148 2503 5152
rect 2507 5148 2508 5152
rect 2502 5147 2508 5148
rect 2710 5152 2716 5153
rect 2710 5148 2711 5152
rect 2715 5148 2716 5152
rect 2710 5147 2716 5148
rect 2356 5113 2366 5115
rect 1975 5106 1979 5107
rect 1975 5101 1979 5102
rect 2119 5106 2123 5107
rect 2119 5101 2123 5102
rect 2303 5106 2307 5107
rect 2303 5101 2307 5102
rect 2327 5106 2331 5107
rect 2327 5101 2331 5102
rect 1499 5078 1503 5079
rect 1499 5073 1503 5074
rect 1579 5078 1583 5079
rect 1579 5073 1583 5074
rect 1787 5078 1791 5079
rect 1787 5073 1791 5074
rect 1935 5078 1939 5079
rect 1976 5078 1978 5101
rect 1935 5073 1939 5074
rect 1974 5077 1980 5078
rect 2120 5077 2122 5101
rect 2328 5077 2330 5101
rect 1974 5073 1975 5077
rect 1979 5073 1980 5077
rect 1490 5055 1496 5056
rect 1490 5051 1491 5055
rect 1495 5051 1496 5055
rect 1490 5050 1496 5051
rect 1318 5019 1324 5020
rect 1318 5015 1319 5019
rect 1323 5015 1324 5019
rect 1318 5014 1324 5015
rect 1500 5012 1502 5073
rect 1626 5055 1632 5056
rect 1626 5051 1627 5055
rect 1631 5051 1632 5055
rect 1626 5050 1632 5051
rect 1628 5020 1630 5050
rect 1626 5019 1632 5020
rect 1626 5015 1627 5019
rect 1631 5015 1632 5019
rect 1626 5014 1632 5015
rect 1788 5012 1790 5073
rect 1936 5013 1938 5073
rect 1974 5072 1980 5073
rect 2118 5076 2124 5077
rect 2118 5072 2119 5076
rect 2123 5072 2124 5076
rect 2118 5071 2124 5072
rect 2326 5076 2332 5077
rect 2326 5072 2327 5076
rect 2331 5072 2332 5076
rect 2326 5071 2332 5072
rect 2090 5061 2096 5062
rect 1974 5060 1980 5061
rect 1974 5056 1975 5060
rect 1979 5056 1980 5060
rect 2090 5057 2091 5061
rect 2095 5057 2096 5061
rect 2090 5056 2096 5057
rect 2298 5061 2304 5062
rect 2298 5057 2299 5061
rect 2303 5057 2304 5061
rect 2298 5056 2304 5057
rect 1974 5055 1980 5056
rect 1934 5012 1940 5013
rect 626 5011 632 5012
rect 626 5007 627 5011
rect 631 5007 632 5011
rect 626 5006 632 5007
rect 898 5011 904 5012
rect 898 5007 899 5011
rect 903 5007 904 5011
rect 898 5006 904 5007
rect 1194 5011 1200 5012
rect 1194 5007 1195 5011
rect 1199 5007 1200 5011
rect 1194 5006 1200 5007
rect 1498 5011 1504 5012
rect 1498 5007 1499 5011
rect 1503 5007 1504 5011
rect 1498 5006 1504 5007
rect 1786 5011 1792 5012
rect 1786 5007 1787 5011
rect 1791 5007 1792 5011
rect 1934 5008 1935 5012
rect 1939 5008 1940 5012
rect 1934 5007 1940 5008
rect 1786 5006 1792 5007
rect 654 4996 660 4997
rect 654 4992 655 4996
rect 659 4992 660 4996
rect 654 4991 660 4992
rect 926 4996 932 4997
rect 926 4992 927 4996
rect 931 4992 932 4996
rect 926 4991 932 4992
rect 1222 4996 1228 4997
rect 1222 4992 1223 4996
rect 1227 4992 1228 4996
rect 1222 4991 1228 4992
rect 1526 4996 1532 4997
rect 1526 4992 1527 4996
rect 1531 4992 1532 4996
rect 1526 4991 1532 4992
rect 1814 4996 1820 4997
rect 1814 4992 1815 4996
rect 1819 4992 1820 4996
rect 1814 4991 1820 4992
rect 1934 4995 1940 4996
rect 1934 4991 1935 4995
rect 1939 4991 1940 4995
rect 656 4939 658 4991
rect 928 4939 930 4991
rect 1224 4939 1226 4991
rect 1528 4939 1530 4991
rect 1816 4939 1818 4991
rect 1934 4990 1940 4991
rect 1936 4939 1938 4990
rect 1976 4987 1978 5055
rect 2092 4987 2094 5056
rect 2178 5043 2184 5044
rect 2178 5039 2179 5043
rect 2183 5039 2184 5043
rect 2178 5038 2184 5039
rect 2180 5020 2182 5038
rect 2178 5019 2184 5020
rect 2178 5015 2179 5019
rect 2183 5015 2184 5019
rect 2178 5014 2184 5015
rect 2300 4987 2302 5056
rect 2356 5052 2358 5113
rect 2504 5107 2506 5147
rect 2712 5107 2714 5147
rect 2503 5106 2507 5107
rect 2503 5101 2507 5102
rect 2535 5106 2539 5107
rect 2535 5101 2539 5102
rect 2711 5106 2715 5107
rect 2711 5101 2715 5102
rect 2751 5106 2755 5107
rect 2751 5101 2755 5102
rect 2536 5077 2538 5101
rect 2752 5077 2754 5101
rect 2534 5076 2540 5077
rect 2534 5072 2535 5076
rect 2539 5072 2540 5076
rect 2534 5071 2540 5072
rect 2750 5076 2756 5077
rect 2750 5072 2751 5076
rect 2755 5072 2756 5076
rect 2750 5071 2756 5072
rect 2506 5061 2512 5062
rect 2506 5057 2507 5061
rect 2511 5057 2512 5061
rect 2506 5056 2512 5057
rect 2722 5061 2728 5062
rect 2722 5057 2723 5061
rect 2727 5057 2728 5061
rect 2722 5056 2728 5057
rect 2354 5051 2360 5052
rect 2354 5047 2355 5051
rect 2359 5047 2360 5051
rect 2354 5046 2360 5047
rect 2508 4987 2510 5056
rect 2724 4987 2726 5056
rect 2772 5052 2774 5202
rect 2812 5176 2814 5206
rect 2810 5175 2816 5176
rect 2810 5171 2811 5175
rect 2815 5171 2816 5175
rect 2810 5170 2816 5171
rect 2892 5168 2894 5229
rect 2980 5176 2982 5258
rect 3092 5235 3094 5300
rect 3178 5287 3184 5288
rect 3178 5283 3179 5287
rect 3183 5283 3184 5287
rect 3178 5282 3184 5283
rect 3180 5264 3182 5282
rect 3178 5263 3184 5264
rect 3178 5259 3179 5263
rect 3183 5259 3184 5263
rect 3178 5258 3184 5259
rect 3300 5235 3302 5300
rect 3314 5295 3320 5296
rect 3314 5291 3315 5295
rect 3319 5291 3320 5295
rect 3314 5290 3320 5291
rect 3410 5295 3416 5296
rect 3410 5291 3411 5295
rect 3415 5291 3416 5295
rect 3410 5290 3416 5291
rect 3316 5264 3318 5290
rect 3314 5263 3320 5264
rect 3314 5259 3315 5263
rect 3319 5259 3320 5263
rect 3314 5258 3320 5259
rect 3091 5234 3095 5235
rect 3091 5229 3095 5230
rect 3099 5234 3103 5235
rect 3099 5229 3103 5230
rect 3299 5234 3303 5235
rect 3299 5229 3303 5230
rect 3307 5234 3311 5235
rect 3307 5229 3311 5230
rect 2978 5175 2984 5176
rect 2978 5171 2979 5175
rect 2983 5171 2984 5175
rect 2978 5170 2984 5171
rect 3078 5175 3084 5176
rect 3078 5171 3079 5175
rect 3083 5171 3084 5175
rect 3078 5170 3084 5171
rect 2890 5167 2896 5168
rect 2890 5163 2891 5167
rect 2895 5163 2896 5167
rect 2890 5162 2896 5163
rect 2918 5152 2924 5153
rect 2918 5148 2919 5152
rect 2923 5148 2924 5152
rect 2918 5147 2924 5148
rect 2920 5107 2922 5147
rect 2919 5106 2923 5107
rect 2919 5101 2923 5102
rect 2975 5106 2979 5107
rect 2975 5101 2979 5102
rect 2976 5077 2978 5101
rect 2974 5076 2980 5077
rect 2974 5072 2975 5076
rect 2979 5072 2980 5076
rect 2974 5071 2980 5072
rect 2946 5061 2952 5062
rect 2946 5057 2947 5061
rect 2951 5057 2952 5061
rect 2946 5056 2952 5057
rect 2770 5051 2776 5052
rect 2770 5047 2771 5051
rect 2775 5047 2776 5051
rect 2770 5046 2776 5047
rect 2838 5003 2844 5004
rect 2838 4999 2839 5003
rect 2843 4999 2844 5003
rect 2838 4998 2844 4999
rect 1975 4986 1979 4987
rect 1975 4981 1979 4982
rect 1995 4986 1999 4987
rect 1995 4981 1999 4982
rect 2091 4986 2095 4987
rect 2091 4981 2095 4982
rect 2131 4986 2135 4987
rect 2131 4981 2135 4982
rect 2267 4986 2271 4987
rect 2267 4981 2271 4982
rect 2299 4986 2303 4987
rect 2299 4981 2303 4982
rect 2419 4986 2423 4987
rect 2419 4981 2423 4982
rect 2507 4986 2511 4987
rect 2507 4981 2511 4982
rect 2619 4986 2623 4987
rect 2619 4981 2623 4982
rect 2723 4986 2727 4987
rect 2723 4981 2727 4982
rect 567 4938 571 4939
rect 567 4933 571 4934
rect 655 4938 659 4939
rect 655 4933 659 4934
rect 703 4938 707 4939
rect 703 4933 707 4934
rect 927 4938 931 4939
rect 927 4933 931 4934
rect 1223 4938 1227 4939
rect 1223 4933 1227 4934
rect 1527 4938 1531 4939
rect 1527 4933 1531 4934
rect 1815 4938 1819 4939
rect 1815 4933 1819 4934
rect 1935 4938 1939 4939
rect 1935 4933 1939 4934
rect 568 4909 570 4933
rect 704 4909 706 4933
rect 1936 4910 1938 4933
rect 1976 4921 1978 4981
rect 1974 4920 1980 4921
rect 1996 4920 1998 4981
rect 2132 4920 2134 4981
rect 2268 4920 2270 4981
rect 2394 4963 2400 4964
rect 2394 4959 2395 4963
rect 2399 4959 2400 4963
rect 2394 4958 2400 4959
rect 2396 4928 2398 4958
rect 2394 4927 2400 4928
rect 2394 4923 2395 4927
rect 2399 4923 2400 4927
rect 2394 4922 2400 4923
rect 2420 4920 2422 4981
rect 2546 4963 2552 4964
rect 2546 4959 2547 4963
rect 2551 4959 2552 4963
rect 2546 4958 2552 4959
rect 2548 4928 2550 4958
rect 2546 4927 2552 4928
rect 2546 4923 2547 4927
rect 2551 4923 2552 4927
rect 2546 4922 2552 4923
rect 2620 4920 2622 4981
rect 2746 4963 2752 4964
rect 2746 4959 2747 4963
rect 2751 4959 2752 4963
rect 2746 4958 2752 4959
rect 2748 4928 2750 4958
rect 2840 4928 2842 4998
rect 2948 4987 2950 5056
rect 3080 5020 3082 5170
rect 3100 5168 3102 5229
rect 3308 5168 3310 5229
rect 3412 5212 3414 5290
rect 3508 5235 3510 5300
rect 3552 5264 3554 5398
rect 3652 5396 3654 5457
rect 3800 5397 3802 5457
rect 3840 5405 3842 5465
rect 3838 5404 3844 5405
rect 4428 5404 4430 5465
rect 4514 5443 4520 5444
rect 4514 5439 4515 5443
rect 4519 5439 4520 5443
rect 4514 5438 4520 5439
rect 3838 5400 3839 5404
rect 3843 5400 3844 5404
rect 3838 5399 3844 5400
rect 4426 5403 4432 5404
rect 4426 5399 4427 5403
rect 4431 5399 4432 5403
rect 4426 5398 4432 5399
rect 3798 5396 3804 5397
rect 3650 5395 3656 5396
rect 3650 5391 3651 5395
rect 3655 5391 3656 5395
rect 3798 5392 3799 5396
rect 3803 5392 3804 5396
rect 3798 5391 3804 5392
rect 3650 5390 3656 5391
rect 4454 5388 4460 5389
rect 3838 5387 3844 5388
rect 3838 5383 3839 5387
rect 3843 5383 3844 5387
rect 4454 5384 4455 5388
rect 4459 5384 4460 5388
rect 4454 5383 4460 5384
rect 3838 5382 3844 5383
rect 3678 5380 3684 5381
rect 3678 5376 3679 5380
rect 3683 5376 3684 5380
rect 3678 5375 3684 5376
rect 3798 5379 3804 5380
rect 3798 5375 3799 5379
rect 3803 5375 3804 5379
rect 3680 5351 3682 5375
rect 3798 5374 3804 5375
rect 3800 5351 3802 5374
rect 3840 5351 3842 5382
rect 4456 5351 4458 5383
rect 3679 5350 3683 5351
rect 3679 5345 3683 5346
rect 3799 5350 3803 5351
rect 3799 5345 3803 5346
rect 3839 5350 3843 5351
rect 3839 5345 3843 5346
rect 4431 5350 4435 5351
rect 4431 5345 4435 5346
rect 4455 5350 4459 5351
rect 4455 5345 4459 5346
rect 3800 5322 3802 5345
rect 3840 5322 3842 5345
rect 3798 5321 3804 5322
rect 3798 5317 3799 5321
rect 3803 5317 3804 5321
rect 3798 5316 3804 5317
rect 3838 5321 3844 5322
rect 4432 5321 4434 5345
rect 3838 5317 3839 5321
rect 3843 5317 3844 5321
rect 3838 5316 3844 5317
rect 4430 5320 4436 5321
rect 4430 5316 4431 5320
rect 4435 5316 4436 5320
rect 4430 5315 4436 5316
rect 4402 5305 4408 5306
rect 3798 5304 3804 5305
rect 3798 5300 3799 5304
rect 3803 5300 3804 5304
rect 3798 5299 3804 5300
rect 3838 5304 3844 5305
rect 3838 5300 3839 5304
rect 3843 5300 3844 5304
rect 4402 5301 4403 5305
rect 4407 5301 4408 5305
rect 4402 5300 4408 5301
rect 3838 5299 3844 5300
rect 3550 5263 3556 5264
rect 3550 5259 3551 5263
rect 3555 5259 3556 5263
rect 3550 5258 3556 5259
rect 3800 5235 3802 5299
rect 3507 5234 3511 5235
rect 3507 5229 3511 5230
rect 3799 5234 3803 5235
rect 3799 5229 3803 5230
rect 3410 5211 3416 5212
rect 3410 5207 3411 5211
rect 3415 5207 3416 5211
rect 3410 5206 3416 5207
rect 3800 5169 3802 5229
rect 3840 5223 3842 5299
rect 4404 5223 4406 5300
rect 4516 5296 4518 5438
rect 4588 5404 4590 5465
rect 4628 5412 4630 5490
rect 4676 5471 4678 5532
rect 4812 5471 4814 5532
rect 4826 5527 4832 5528
rect 4826 5523 4827 5527
rect 4831 5523 4832 5527
rect 4826 5522 4832 5523
rect 4828 5496 4830 5522
rect 4886 5519 4892 5520
rect 4886 5515 4887 5519
rect 4891 5515 4892 5519
rect 4886 5514 4892 5515
rect 4826 5495 4832 5496
rect 4826 5491 4827 5495
rect 4831 5491 4832 5495
rect 4826 5490 4832 5491
rect 4675 5470 4679 5471
rect 4675 5465 4679 5466
rect 4747 5470 4751 5471
rect 4747 5465 4751 5466
rect 4811 5470 4815 5471
rect 4811 5465 4815 5466
rect 4626 5411 4632 5412
rect 4626 5407 4627 5411
rect 4631 5407 4632 5411
rect 4626 5406 4632 5407
rect 4748 5404 4750 5465
rect 4888 5448 4890 5514
rect 4912 5512 4914 5630
rect 5664 5629 5666 5689
rect 5662 5628 5668 5629
rect 5662 5624 5663 5628
rect 5667 5624 5668 5628
rect 5662 5623 5668 5624
rect 5662 5611 5668 5612
rect 5662 5607 5663 5611
rect 5667 5607 5668 5611
rect 5662 5606 5668 5607
rect 5664 5583 5666 5606
rect 4975 5582 4979 5583
rect 4975 5577 4979 5578
rect 5111 5582 5115 5583
rect 5111 5577 5115 5578
rect 5663 5582 5667 5583
rect 5663 5577 5667 5578
rect 4976 5553 4978 5577
rect 5112 5553 5114 5577
rect 5664 5554 5666 5577
rect 5662 5553 5668 5554
rect 4974 5552 4980 5553
rect 4974 5548 4975 5552
rect 4979 5548 4980 5552
rect 4974 5547 4980 5548
rect 5110 5552 5116 5553
rect 5110 5548 5111 5552
rect 5115 5548 5116 5552
rect 5662 5549 5663 5553
rect 5667 5549 5668 5553
rect 5662 5548 5668 5549
rect 5110 5547 5116 5548
rect 4946 5537 4952 5538
rect 4946 5533 4947 5537
rect 4951 5533 4952 5537
rect 4946 5532 4952 5533
rect 5082 5537 5088 5538
rect 5082 5533 5083 5537
rect 5087 5533 5088 5537
rect 5082 5532 5088 5533
rect 5662 5536 5668 5537
rect 5662 5532 5663 5536
rect 5667 5532 5668 5536
rect 4910 5511 4916 5512
rect 4910 5507 4911 5511
rect 4915 5507 4916 5511
rect 4910 5506 4916 5507
rect 4948 5471 4950 5532
rect 4962 5527 4968 5528
rect 4962 5523 4963 5527
rect 4967 5523 4968 5527
rect 4962 5522 4968 5523
rect 4964 5496 4966 5522
rect 4962 5495 4968 5496
rect 4962 5491 4963 5495
rect 4967 5491 4968 5495
rect 4962 5490 4968 5491
rect 5084 5471 5086 5532
rect 5662 5531 5668 5532
rect 5098 5527 5104 5528
rect 5098 5523 5099 5527
rect 5103 5523 5104 5527
rect 5098 5522 5104 5523
rect 5100 5496 5102 5522
rect 5098 5495 5104 5496
rect 5098 5491 5099 5495
rect 5103 5491 5104 5495
rect 5098 5490 5104 5491
rect 5664 5471 5666 5531
rect 4907 5470 4911 5471
rect 4907 5465 4911 5466
rect 4947 5470 4951 5471
rect 4947 5465 4951 5466
rect 5075 5470 5079 5471
rect 5075 5465 5079 5466
rect 5083 5470 5087 5471
rect 5083 5465 5087 5466
rect 5663 5470 5667 5471
rect 5663 5465 5667 5466
rect 4886 5447 4892 5448
rect 4886 5443 4887 5447
rect 4891 5443 4892 5447
rect 4886 5442 4892 5443
rect 4908 5404 4910 5465
rect 5076 5404 5078 5465
rect 5198 5411 5204 5412
rect 5198 5407 5199 5411
rect 5203 5407 5204 5411
rect 5198 5406 5204 5407
rect 4586 5403 4592 5404
rect 4586 5399 4587 5403
rect 4591 5399 4592 5403
rect 4586 5398 4592 5399
rect 4746 5403 4752 5404
rect 4746 5399 4747 5403
rect 4751 5399 4752 5403
rect 4746 5398 4752 5399
rect 4906 5403 4912 5404
rect 4906 5399 4907 5403
rect 4911 5399 4912 5403
rect 4906 5398 4912 5399
rect 5074 5403 5080 5404
rect 5074 5399 5075 5403
rect 5079 5399 5080 5403
rect 5074 5398 5080 5399
rect 4614 5388 4620 5389
rect 4614 5384 4615 5388
rect 4619 5384 4620 5388
rect 4614 5383 4620 5384
rect 4774 5388 4780 5389
rect 4774 5384 4775 5388
rect 4779 5384 4780 5388
rect 4774 5383 4780 5384
rect 4934 5388 4940 5389
rect 4934 5384 4935 5388
rect 4939 5384 4940 5388
rect 4934 5383 4940 5384
rect 5102 5388 5108 5389
rect 5102 5384 5103 5388
rect 5107 5384 5108 5388
rect 5102 5383 5108 5384
rect 4616 5351 4618 5383
rect 4776 5351 4778 5383
rect 4936 5351 4938 5383
rect 5104 5351 5106 5383
rect 4615 5350 4619 5351
rect 4615 5345 4619 5346
rect 4775 5350 4779 5351
rect 4775 5345 4779 5346
rect 4799 5350 4803 5351
rect 4799 5345 4803 5346
rect 4935 5350 4939 5351
rect 4935 5345 4939 5346
rect 4983 5350 4987 5351
rect 4983 5345 4987 5346
rect 5103 5350 5107 5351
rect 5103 5345 5107 5346
rect 5175 5350 5179 5351
rect 5175 5345 5179 5346
rect 4616 5321 4618 5345
rect 4800 5321 4802 5345
rect 4984 5321 4986 5345
rect 5176 5321 5178 5345
rect 4614 5320 4620 5321
rect 4614 5316 4615 5320
rect 4619 5316 4620 5320
rect 4614 5315 4620 5316
rect 4798 5320 4804 5321
rect 4798 5316 4799 5320
rect 4803 5316 4804 5320
rect 4798 5315 4804 5316
rect 4982 5320 4988 5321
rect 4982 5316 4983 5320
rect 4987 5316 4988 5320
rect 4982 5315 4988 5316
rect 5174 5320 5180 5321
rect 5174 5316 5175 5320
rect 5179 5316 5180 5320
rect 5174 5315 5180 5316
rect 4586 5305 4592 5306
rect 4586 5301 4587 5305
rect 4591 5301 4592 5305
rect 4586 5300 4592 5301
rect 4770 5305 4776 5306
rect 4770 5301 4771 5305
rect 4775 5301 4776 5305
rect 4770 5300 4776 5301
rect 4954 5305 4960 5306
rect 4954 5301 4955 5305
rect 4959 5301 4960 5305
rect 4954 5300 4960 5301
rect 5146 5305 5152 5306
rect 5146 5301 5147 5305
rect 5151 5301 5152 5305
rect 5146 5300 5152 5301
rect 4514 5295 4520 5296
rect 4514 5291 4515 5295
rect 4519 5291 4520 5295
rect 4514 5290 4520 5291
rect 4566 5295 4572 5296
rect 4566 5291 4567 5295
rect 4571 5291 4572 5295
rect 4566 5290 4572 5291
rect 4568 5264 4570 5290
rect 4566 5263 4572 5264
rect 4566 5259 4567 5263
rect 4571 5259 4572 5263
rect 4566 5258 4572 5259
rect 4588 5223 4590 5300
rect 4602 5263 4608 5264
rect 4602 5259 4603 5263
rect 4607 5259 4608 5263
rect 4602 5258 4608 5259
rect 3839 5222 3843 5223
rect 3839 5217 3843 5218
rect 4403 5222 4407 5223
rect 4403 5217 4407 5218
rect 4435 5222 4439 5223
rect 4435 5217 4439 5218
rect 4587 5222 4591 5223
rect 4587 5217 4591 5218
rect 4595 5222 4599 5223
rect 4595 5217 4599 5218
rect 3798 5168 3804 5169
rect 3098 5167 3104 5168
rect 3098 5163 3099 5167
rect 3103 5163 3104 5167
rect 3098 5162 3104 5163
rect 3306 5167 3312 5168
rect 3306 5163 3307 5167
rect 3311 5163 3312 5167
rect 3798 5164 3799 5168
rect 3803 5164 3804 5168
rect 3798 5163 3804 5164
rect 3306 5162 3312 5163
rect 3840 5157 3842 5217
rect 4426 5199 4432 5200
rect 4426 5195 4427 5199
rect 4431 5195 4432 5199
rect 4426 5194 4432 5195
rect 3838 5156 3844 5157
rect 3126 5152 3132 5153
rect 3126 5148 3127 5152
rect 3131 5148 3132 5152
rect 3126 5147 3132 5148
rect 3334 5152 3340 5153
rect 3838 5152 3839 5156
rect 3843 5152 3844 5156
rect 3334 5148 3335 5152
rect 3339 5148 3340 5152
rect 3334 5147 3340 5148
rect 3798 5151 3804 5152
rect 3838 5151 3844 5152
rect 3798 5147 3799 5151
rect 3803 5147 3804 5151
rect 3128 5107 3130 5147
rect 3336 5107 3338 5147
rect 3798 5146 3804 5147
rect 3800 5107 3802 5146
rect 3838 5139 3844 5140
rect 3838 5135 3839 5139
rect 3843 5135 3844 5139
rect 3838 5134 3844 5135
rect 3127 5106 3131 5107
rect 3127 5101 3131 5102
rect 3207 5106 3211 5107
rect 3207 5101 3211 5102
rect 3335 5106 3339 5107
rect 3335 5101 3339 5102
rect 3799 5106 3803 5107
rect 3840 5103 3842 5134
rect 3799 5101 3803 5102
rect 3839 5102 3843 5103
rect 3208 5077 3210 5101
rect 3800 5078 3802 5101
rect 3839 5097 3843 5098
rect 3887 5102 3891 5103
rect 3887 5097 3891 5098
rect 4087 5102 4091 5103
rect 4087 5097 4091 5098
rect 4327 5102 4331 5103
rect 4327 5097 4331 5098
rect 3798 5077 3804 5078
rect 3206 5076 3212 5077
rect 3206 5072 3207 5076
rect 3211 5072 3212 5076
rect 3798 5073 3799 5077
rect 3803 5073 3804 5077
rect 3840 5074 3842 5097
rect 3798 5072 3804 5073
rect 3838 5073 3844 5074
rect 3888 5073 3890 5097
rect 4088 5073 4090 5097
rect 4328 5073 4330 5097
rect 3206 5071 3212 5072
rect 3838 5069 3839 5073
rect 3843 5069 3844 5073
rect 3838 5068 3844 5069
rect 3886 5072 3892 5073
rect 3886 5068 3887 5072
rect 3891 5068 3892 5072
rect 3886 5067 3892 5068
rect 4086 5072 4092 5073
rect 4086 5068 4087 5072
rect 4091 5068 4092 5072
rect 4086 5067 4092 5068
rect 4326 5072 4332 5073
rect 4326 5068 4327 5072
rect 4331 5068 4332 5072
rect 4326 5067 4332 5068
rect 3178 5061 3184 5062
rect 3178 5057 3179 5061
rect 3183 5057 3184 5061
rect 3178 5056 3184 5057
rect 3798 5060 3804 5061
rect 3798 5056 3799 5060
rect 3803 5056 3804 5060
rect 3858 5057 3864 5058
rect 3078 5019 3084 5020
rect 3078 5015 3079 5019
rect 3083 5015 3084 5019
rect 3078 5014 3084 5015
rect 3180 4987 3182 5056
rect 3798 5055 3804 5056
rect 3838 5056 3844 5057
rect 3194 5051 3200 5052
rect 3194 5047 3195 5051
rect 3199 5047 3200 5051
rect 3194 5046 3200 5047
rect 3196 5020 3198 5046
rect 3194 5019 3200 5020
rect 3194 5015 3195 5019
rect 3199 5015 3200 5019
rect 3194 5014 3200 5015
rect 3246 5003 3252 5004
rect 3246 4999 3247 5003
rect 3251 4999 3252 5003
rect 3246 4998 3252 4999
rect 2859 4986 2863 4987
rect 2859 4981 2863 4982
rect 2947 4986 2951 4987
rect 2947 4981 2951 4982
rect 3123 4986 3127 4987
rect 3123 4981 3127 4982
rect 3179 4986 3183 4987
rect 3179 4981 3183 4982
rect 2746 4927 2752 4928
rect 2746 4923 2747 4927
rect 2751 4923 2752 4927
rect 2746 4922 2752 4923
rect 2838 4927 2844 4928
rect 2838 4923 2839 4927
rect 2843 4923 2844 4927
rect 2838 4922 2844 4923
rect 2860 4920 2862 4981
rect 2962 4963 2968 4964
rect 2962 4959 2963 4963
rect 2967 4959 2968 4963
rect 2962 4958 2968 4959
rect 1974 4916 1975 4920
rect 1979 4916 1980 4920
rect 1974 4915 1980 4916
rect 1994 4919 2000 4920
rect 1994 4915 1995 4919
rect 1999 4915 2000 4919
rect 1994 4914 2000 4915
rect 2130 4919 2136 4920
rect 2130 4915 2131 4919
rect 2135 4915 2136 4919
rect 2130 4914 2136 4915
rect 2266 4919 2272 4920
rect 2266 4915 2267 4919
rect 2271 4915 2272 4919
rect 2266 4914 2272 4915
rect 2418 4919 2424 4920
rect 2418 4915 2419 4919
rect 2423 4915 2424 4919
rect 2418 4914 2424 4915
rect 2618 4919 2624 4920
rect 2618 4915 2619 4919
rect 2623 4915 2624 4919
rect 2618 4914 2624 4915
rect 2858 4919 2864 4920
rect 2858 4915 2859 4919
rect 2863 4915 2864 4919
rect 2858 4914 2864 4915
rect 1934 4909 1940 4910
rect 566 4908 572 4909
rect 566 4904 567 4908
rect 571 4904 572 4908
rect 566 4903 572 4904
rect 702 4908 708 4909
rect 702 4904 703 4908
rect 707 4904 708 4908
rect 1934 4905 1935 4909
rect 1939 4905 1940 4909
rect 1934 4904 1940 4905
rect 2022 4904 2028 4905
rect 702 4903 708 4904
rect 1974 4903 1980 4904
rect 1974 4899 1975 4903
rect 1979 4899 1980 4903
rect 2022 4900 2023 4904
rect 2027 4900 2028 4904
rect 2022 4899 2028 4900
rect 2158 4904 2164 4905
rect 2158 4900 2159 4904
rect 2163 4900 2164 4904
rect 2158 4899 2164 4900
rect 2294 4904 2300 4905
rect 2294 4900 2295 4904
rect 2299 4900 2300 4904
rect 2294 4899 2300 4900
rect 2446 4904 2452 4905
rect 2446 4900 2447 4904
rect 2451 4900 2452 4904
rect 2446 4899 2452 4900
rect 2646 4904 2652 4905
rect 2646 4900 2647 4904
rect 2651 4900 2652 4904
rect 2646 4899 2652 4900
rect 2886 4904 2892 4905
rect 2886 4900 2887 4904
rect 2891 4900 2892 4904
rect 2886 4899 2892 4900
rect 1974 4898 1980 4899
rect 538 4893 544 4894
rect 538 4889 539 4893
rect 543 4889 544 4893
rect 538 4888 544 4889
rect 674 4893 680 4894
rect 674 4889 675 4893
rect 679 4889 680 4893
rect 674 4888 680 4889
rect 1934 4892 1940 4893
rect 1934 4888 1935 4892
rect 1939 4888 1940 4892
rect 490 4851 496 4852
rect 490 4847 491 4851
rect 495 4847 496 4851
rect 490 4846 496 4847
rect 540 4815 542 4888
rect 554 4883 560 4884
rect 554 4879 555 4883
rect 559 4879 560 4883
rect 554 4878 560 4879
rect 556 4852 558 4878
rect 554 4851 560 4852
rect 554 4847 555 4851
rect 559 4847 560 4851
rect 554 4846 560 4847
rect 676 4815 678 4888
rect 1934 4887 1940 4888
rect 690 4883 696 4884
rect 690 4879 691 4883
rect 695 4879 696 4883
rect 690 4878 696 4879
rect 692 4852 694 4878
rect 690 4851 696 4852
rect 690 4847 691 4851
rect 695 4847 696 4851
rect 690 4846 696 4847
rect 1936 4815 1938 4887
rect 1976 4867 1978 4898
rect 2024 4867 2026 4899
rect 2160 4867 2162 4899
rect 2296 4867 2298 4899
rect 2448 4867 2450 4899
rect 2648 4867 2650 4899
rect 2888 4867 2890 4899
rect 1975 4866 1979 4867
rect 1975 4861 1979 4862
rect 2023 4866 2027 4867
rect 2023 4861 2027 4862
rect 2159 4866 2163 4867
rect 2159 4861 2163 4862
rect 2295 4866 2299 4867
rect 2295 4861 2299 4862
rect 2327 4866 2331 4867
rect 2327 4861 2331 4862
rect 2447 4866 2451 4867
rect 2447 4861 2451 4862
rect 2559 4866 2563 4867
rect 2559 4861 2563 4862
rect 2647 4866 2651 4867
rect 2647 4861 2651 4862
rect 2823 4866 2827 4867
rect 2823 4861 2827 4862
rect 2887 4866 2891 4867
rect 2887 4861 2891 4862
rect 1976 4838 1978 4861
rect 1974 4837 1980 4838
rect 2328 4837 2330 4861
rect 2560 4837 2562 4861
rect 2824 4837 2826 4861
rect 1974 4833 1975 4837
rect 1979 4833 1980 4837
rect 1974 4832 1980 4833
rect 2326 4836 2332 4837
rect 2326 4832 2327 4836
rect 2331 4832 2332 4836
rect 2326 4831 2332 4832
rect 2558 4836 2564 4837
rect 2558 4832 2559 4836
rect 2563 4832 2564 4836
rect 2558 4831 2564 4832
rect 2822 4836 2828 4837
rect 2822 4832 2823 4836
rect 2827 4832 2828 4836
rect 2822 4831 2828 4832
rect 2298 4821 2304 4822
rect 1974 4820 1980 4821
rect 1974 4816 1975 4820
rect 1979 4816 1980 4820
rect 2298 4817 2299 4821
rect 2303 4817 2304 4821
rect 2298 4816 2304 4817
rect 2530 4821 2536 4822
rect 2530 4817 2531 4821
rect 2535 4817 2536 4821
rect 2530 4816 2536 4817
rect 2794 4821 2800 4822
rect 2794 4817 2795 4821
rect 2799 4817 2800 4821
rect 2794 4816 2800 4817
rect 1974 4815 1980 4816
rect 267 4814 271 4815
rect 267 4809 271 4810
rect 403 4814 407 4815
rect 403 4809 407 4810
rect 539 4814 543 4815
rect 539 4809 543 4810
rect 675 4814 679 4815
rect 675 4809 679 4810
rect 1935 4814 1939 4815
rect 1935 4809 1939 4810
rect 234 4791 240 4792
rect 234 4787 235 4791
rect 239 4787 240 4791
rect 234 4786 240 4787
rect 258 4791 264 4792
rect 258 4787 259 4791
rect 263 4787 264 4791
rect 258 4786 264 4787
rect 218 4763 224 4764
rect 218 4759 219 4763
rect 223 4759 224 4763
rect 218 4758 224 4759
rect 110 4744 111 4748
rect 115 4744 116 4748
rect 110 4743 116 4744
rect 130 4747 136 4748
rect 130 4743 131 4747
rect 135 4743 136 4747
rect 130 4742 136 4743
rect 158 4732 164 4733
rect 110 4731 116 4732
rect 110 4727 111 4731
rect 115 4727 116 4731
rect 158 4728 159 4732
rect 163 4728 164 4732
rect 158 4727 164 4728
rect 110 4726 116 4727
rect 112 4699 114 4726
rect 160 4699 162 4727
rect 111 4698 115 4699
rect 111 4693 115 4694
rect 159 4698 163 4699
rect 159 4693 163 4694
rect 112 4670 114 4693
rect 110 4669 116 4670
rect 160 4669 162 4693
rect 110 4665 111 4669
rect 115 4665 116 4669
rect 110 4664 116 4665
rect 158 4668 164 4669
rect 158 4664 159 4668
rect 163 4664 164 4668
rect 158 4663 164 4664
rect 130 4653 136 4654
rect 110 4652 116 4653
rect 110 4648 111 4652
rect 115 4648 116 4652
rect 130 4649 131 4653
rect 135 4649 136 4653
rect 130 4648 136 4649
rect 110 4647 116 4648
rect 112 4575 114 4647
rect 132 4575 134 4648
rect 220 4612 222 4758
rect 260 4756 262 4786
rect 258 4755 264 4756
rect 258 4751 259 4755
rect 263 4751 264 4755
rect 258 4750 264 4751
rect 268 4748 270 4809
rect 394 4791 400 4792
rect 394 4787 395 4791
rect 399 4787 400 4791
rect 394 4786 400 4787
rect 396 4756 398 4786
rect 394 4755 400 4756
rect 394 4751 395 4755
rect 399 4751 400 4755
rect 394 4750 400 4751
rect 404 4748 406 4809
rect 530 4791 536 4792
rect 530 4787 531 4791
rect 535 4787 536 4791
rect 530 4786 536 4787
rect 532 4756 534 4786
rect 530 4755 536 4756
rect 530 4751 531 4755
rect 535 4751 536 4755
rect 530 4750 536 4751
rect 540 4748 542 4809
rect 666 4791 672 4792
rect 666 4787 667 4791
rect 671 4787 672 4791
rect 666 4786 672 4787
rect 668 4756 670 4786
rect 666 4755 672 4756
rect 666 4751 667 4755
rect 671 4751 672 4755
rect 666 4750 672 4751
rect 676 4748 678 4809
rect 1936 4749 1938 4809
rect 1934 4748 1940 4749
rect 266 4747 272 4748
rect 266 4743 267 4747
rect 271 4743 272 4747
rect 266 4742 272 4743
rect 402 4747 408 4748
rect 402 4743 403 4747
rect 407 4743 408 4747
rect 402 4742 408 4743
rect 538 4747 544 4748
rect 538 4743 539 4747
rect 543 4743 544 4747
rect 538 4742 544 4743
rect 674 4747 680 4748
rect 674 4743 675 4747
rect 679 4743 680 4747
rect 1934 4744 1935 4748
rect 1939 4744 1940 4748
rect 1934 4743 1940 4744
rect 1976 4743 1978 4815
rect 2300 4743 2302 4816
rect 2386 4779 2392 4780
rect 2386 4775 2387 4779
rect 2391 4775 2392 4779
rect 2386 4774 2392 4775
rect 674 4742 680 4743
rect 1975 4742 1979 4743
rect 1975 4737 1979 4738
rect 2019 4742 2023 4743
rect 2019 4737 2023 4738
rect 2195 4742 2199 4743
rect 2195 4737 2199 4738
rect 2299 4742 2303 4743
rect 2299 4737 2303 4738
rect 2371 4742 2375 4743
rect 2371 4737 2375 4738
rect 294 4732 300 4733
rect 294 4728 295 4732
rect 299 4728 300 4732
rect 294 4727 300 4728
rect 430 4732 436 4733
rect 430 4728 431 4732
rect 435 4728 436 4732
rect 430 4727 436 4728
rect 566 4732 572 4733
rect 566 4728 567 4732
rect 571 4728 572 4732
rect 566 4727 572 4728
rect 702 4732 708 4733
rect 702 4728 703 4732
rect 707 4728 708 4732
rect 702 4727 708 4728
rect 1934 4731 1940 4732
rect 1934 4727 1935 4731
rect 1939 4727 1940 4731
rect 296 4699 298 4727
rect 432 4699 434 4727
rect 568 4699 570 4727
rect 704 4699 706 4727
rect 1934 4726 1940 4727
rect 1936 4699 1938 4726
rect 295 4698 299 4699
rect 295 4693 299 4694
rect 431 4698 435 4699
rect 431 4693 435 4694
rect 567 4698 571 4699
rect 567 4693 571 4694
rect 703 4698 707 4699
rect 703 4693 707 4694
rect 1935 4698 1939 4699
rect 1935 4693 1939 4694
rect 296 4669 298 4693
rect 432 4669 434 4693
rect 568 4669 570 4693
rect 704 4669 706 4693
rect 1936 4670 1938 4693
rect 1976 4677 1978 4737
rect 1974 4676 1980 4677
rect 2020 4676 2022 4737
rect 2146 4719 2152 4720
rect 2106 4715 2112 4716
rect 2106 4711 2107 4715
rect 2111 4711 2112 4715
rect 2146 4715 2147 4719
rect 2151 4715 2152 4719
rect 2146 4714 2152 4715
rect 2106 4710 2112 4711
rect 1974 4672 1975 4676
rect 1979 4672 1980 4676
rect 1974 4671 1980 4672
rect 2018 4675 2024 4676
rect 2018 4671 2019 4675
rect 2023 4671 2024 4675
rect 2018 4670 2024 4671
rect 1934 4669 1940 4670
rect 294 4668 300 4669
rect 294 4664 295 4668
rect 299 4664 300 4668
rect 294 4663 300 4664
rect 430 4668 436 4669
rect 430 4664 431 4668
rect 435 4664 436 4668
rect 430 4663 436 4664
rect 566 4668 572 4669
rect 566 4664 567 4668
rect 571 4664 572 4668
rect 566 4663 572 4664
rect 702 4668 708 4669
rect 702 4664 703 4668
rect 707 4664 708 4668
rect 1934 4665 1935 4669
rect 1939 4665 1940 4669
rect 1934 4664 1940 4665
rect 702 4663 708 4664
rect 2046 4660 2052 4661
rect 1974 4659 1980 4660
rect 1974 4655 1975 4659
rect 1979 4655 1980 4659
rect 2046 4656 2047 4660
rect 2051 4656 2052 4660
rect 2046 4655 2052 4656
rect 1974 4654 1980 4655
rect 266 4653 272 4654
rect 266 4649 267 4653
rect 271 4649 272 4653
rect 266 4648 272 4649
rect 402 4653 408 4654
rect 402 4649 403 4653
rect 407 4649 408 4653
rect 402 4648 408 4649
rect 538 4653 544 4654
rect 538 4649 539 4653
rect 543 4649 544 4653
rect 538 4648 544 4649
rect 674 4653 680 4654
rect 674 4649 675 4653
rect 679 4649 680 4653
rect 674 4648 680 4649
rect 1934 4652 1940 4653
rect 1934 4648 1935 4652
rect 1939 4648 1940 4652
rect 218 4611 224 4612
rect 218 4607 219 4611
rect 223 4607 224 4611
rect 218 4606 224 4607
rect 268 4575 270 4648
rect 282 4643 288 4644
rect 282 4639 283 4643
rect 287 4639 288 4643
rect 282 4638 288 4639
rect 284 4612 286 4638
rect 282 4611 288 4612
rect 282 4607 283 4611
rect 287 4607 288 4611
rect 282 4606 288 4607
rect 404 4575 406 4648
rect 418 4643 424 4644
rect 418 4639 419 4643
rect 423 4639 424 4643
rect 418 4638 424 4639
rect 420 4612 422 4638
rect 418 4611 424 4612
rect 418 4607 419 4611
rect 423 4607 424 4611
rect 418 4606 424 4607
rect 540 4575 542 4648
rect 554 4643 560 4644
rect 554 4639 555 4643
rect 559 4639 560 4643
rect 554 4638 560 4639
rect 556 4612 558 4638
rect 554 4611 560 4612
rect 554 4607 555 4611
rect 559 4607 560 4611
rect 554 4606 560 4607
rect 676 4575 678 4648
rect 1934 4647 1940 4648
rect 690 4643 696 4644
rect 690 4639 691 4643
rect 695 4639 696 4643
rect 690 4638 696 4639
rect 754 4643 760 4644
rect 754 4639 755 4643
rect 759 4639 760 4643
rect 754 4638 760 4639
rect 692 4612 694 4638
rect 690 4611 696 4612
rect 690 4607 691 4611
rect 695 4607 696 4611
rect 690 4606 696 4607
rect 111 4574 115 4575
rect 111 4569 115 4570
rect 131 4574 135 4575
rect 131 4569 135 4570
rect 251 4574 255 4575
rect 251 4569 255 4570
rect 267 4574 271 4575
rect 267 4569 271 4570
rect 403 4574 407 4575
rect 403 4569 407 4570
rect 443 4574 447 4575
rect 443 4569 447 4570
rect 539 4574 543 4575
rect 651 4574 655 4575
rect 539 4569 543 4570
rect 578 4571 584 4572
rect 112 4509 114 4569
rect 110 4508 116 4509
rect 252 4508 254 4569
rect 378 4551 384 4552
rect 378 4547 379 4551
rect 383 4547 384 4551
rect 378 4546 384 4547
rect 380 4516 382 4546
rect 378 4515 384 4516
rect 378 4511 379 4515
rect 383 4511 384 4515
rect 378 4510 384 4511
rect 444 4508 446 4569
rect 578 4567 579 4571
rect 583 4567 584 4571
rect 651 4569 655 4570
rect 675 4574 679 4575
rect 675 4569 679 4570
rect 578 4566 584 4567
rect 566 4551 572 4552
rect 566 4547 567 4551
rect 571 4547 572 4551
rect 566 4546 572 4547
rect 568 4516 570 4546
rect 566 4515 572 4516
rect 566 4511 567 4515
rect 571 4511 572 4515
rect 566 4510 572 4511
rect 110 4504 111 4508
rect 115 4504 116 4508
rect 110 4503 116 4504
rect 250 4507 256 4508
rect 250 4503 251 4507
rect 255 4503 256 4507
rect 250 4502 256 4503
rect 442 4507 448 4508
rect 442 4503 443 4507
rect 447 4503 448 4507
rect 442 4502 448 4503
rect 278 4492 284 4493
rect 110 4491 116 4492
rect 110 4487 111 4491
rect 115 4487 116 4491
rect 278 4488 279 4492
rect 283 4488 284 4492
rect 278 4487 284 4488
rect 470 4492 476 4493
rect 470 4488 471 4492
rect 475 4488 476 4492
rect 470 4487 476 4488
rect 110 4486 116 4487
rect 112 4463 114 4486
rect 280 4463 282 4487
rect 472 4463 474 4487
rect 111 4462 115 4463
rect 111 4457 115 4458
rect 279 4462 283 4463
rect 279 4457 283 4458
rect 471 4462 475 4463
rect 471 4457 475 4458
rect 511 4462 515 4463
rect 511 4457 515 4458
rect 112 4434 114 4457
rect 110 4433 116 4434
rect 512 4433 514 4457
rect 110 4429 111 4433
rect 115 4429 116 4433
rect 110 4428 116 4429
rect 510 4432 516 4433
rect 510 4428 511 4432
rect 515 4428 516 4432
rect 510 4427 516 4428
rect 482 4417 488 4418
rect 110 4416 116 4417
rect 110 4412 111 4416
rect 115 4412 116 4416
rect 482 4413 483 4417
rect 487 4413 488 4417
rect 482 4412 488 4413
rect 110 4411 116 4412
rect 112 4347 114 4411
rect 484 4347 486 4412
rect 580 4376 582 4566
rect 652 4508 654 4569
rect 756 4564 758 4638
rect 1936 4575 1938 4647
rect 1976 4627 1978 4654
rect 2048 4627 2050 4655
rect 1975 4626 1979 4627
rect 1975 4621 1979 4622
rect 2023 4626 2027 4627
rect 2023 4621 2027 4622
rect 2047 4626 2051 4627
rect 2047 4621 2051 4622
rect 1976 4598 1978 4621
rect 1974 4597 1980 4598
rect 2024 4597 2026 4621
rect 1974 4593 1975 4597
rect 1979 4593 1980 4597
rect 1974 4592 1980 4593
rect 2022 4596 2028 4597
rect 2022 4592 2023 4596
rect 2027 4592 2028 4596
rect 2022 4591 2028 4592
rect 1994 4581 2000 4582
rect 1974 4580 1980 4581
rect 1974 4576 1975 4580
rect 1979 4576 1980 4580
rect 1994 4577 1995 4581
rect 1999 4577 2000 4581
rect 1994 4576 2000 4577
rect 1974 4575 1980 4576
rect 875 4574 879 4575
rect 875 4569 879 4570
rect 1099 4574 1103 4575
rect 1331 4574 1335 4575
rect 1099 4569 1103 4570
rect 1222 4571 1228 4572
rect 754 4563 760 4564
rect 754 4559 755 4563
rect 759 4559 760 4563
rect 754 4558 760 4559
rect 778 4551 784 4552
rect 778 4547 779 4551
rect 783 4547 784 4551
rect 778 4546 784 4547
rect 780 4516 782 4546
rect 778 4515 784 4516
rect 778 4511 779 4515
rect 783 4511 784 4515
rect 778 4510 784 4511
rect 876 4508 878 4569
rect 1002 4551 1008 4552
rect 1002 4547 1003 4551
rect 1007 4547 1008 4551
rect 1002 4546 1008 4547
rect 1004 4516 1006 4546
rect 1002 4515 1008 4516
rect 1002 4511 1003 4515
rect 1007 4511 1008 4515
rect 1002 4510 1008 4511
rect 1100 4508 1102 4569
rect 1222 4567 1223 4571
rect 1227 4567 1228 4571
rect 1331 4569 1335 4570
rect 1571 4574 1575 4575
rect 1571 4569 1575 4570
rect 1787 4574 1791 4575
rect 1787 4569 1791 4570
rect 1935 4574 1939 4575
rect 1935 4569 1939 4570
rect 1222 4566 1228 4567
rect 1224 4516 1226 4566
rect 1222 4515 1228 4516
rect 1222 4511 1223 4515
rect 1227 4511 1228 4515
rect 1222 4510 1228 4511
rect 1332 4508 1334 4569
rect 1522 4551 1528 4552
rect 1522 4547 1523 4551
rect 1527 4547 1528 4551
rect 1522 4546 1528 4547
rect 1524 4516 1526 4546
rect 1562 4543 1568 4544
rect 1562 4539 1563 4543
rect 1567 4539 1568 4543
rect 1562 4538 1568 4539
rect 1522 4515 1528 4516
rect 1522 4511 1523 4515
rect 1527 4511 1528 4515
rect 1522 4510 1528 4511
rect 650 4507 656 4508
rect 650 4503 651 4507
rect 655 4503 656 4507
rect 650 4502 656 4503
rect 874 4507 880 4508
rect 874 4503 875 4507
rect 879 4503 880 4507
rect 874 4502 880 4503
rect 1098 4507 1104 4508
rect 1098 4503 1099 4507
rect 1103 4503 1104 4507
rect 1098 4502 1104 4503
rect 1330 4507 1336 4508
rect 1330 4503 1331 4507
rect 1335 4503 1336 4507
rect 1330 4502 1336 4503
rect 678 4492 684 4493
rect 678 4488 679 4492
rect 683 4488 684 4492
rect 678 4487 684 4488
rect 902 4492 908 4493
rect 902 4488 903 4492
rect 907 4488 908 4492
rect 902 4487 908 4488
rect 1126 4492 1132 4493
rect 1126 4488 1127 4492
rect 1131 4488 1132 4492
rect 1126 4487 1132 4488
rect 1358 4492 1364 4493
rect 1358 4488 1359 4492
rect 1363 4488 1364 4492
rect 1358 4487 1364 4488
rect 680 4463 682 4487
rect 904 4463 906 4487
rect 1128 4463 1130 4487
rect 1360 4463 1362 4487
rect 679 4462 683 4463
rect 679 4457 683 4458
rect 687 4462 691 4463
rect 687 4457 691 4458
rect 871 4462 875 4463
rect 871 4457 875 4458
rect 903 4462 907 4463
rect 903 4457 907 4458
rect 1071 4462 1075 4463
rect 1071 4457 1075 4458
rect 1127 4462 1131 4463
rect 1127 4457 1131 4458
rect 1279 4462 1283 4463
rect 1279 4457 1283 4458
rect 1359 4462 1363 4463
rect 1359 4457 1363 4458
rect 1495 4462 1499 4463
rect 1495 4457 1499 4458
rect 688 4433 690 4457
rect 872 4433 874 4457
rect 1072 4433 1074 4457
rect 1280 4433 1282 4457
rect 1496 4433 1498 4457
rect 686 4432 692 4433
rect 686 4428 687 4432
rect 691 4428 692 4432
rect 686 4427 692 4428
rect 870 4432 876 4433
rect 870 4428 871 4432
rect 875 4428 876 4432
rect 870 4427 876 4428
rect 1070 4432 1076 4433
rect 1070 4428 1071 4432
rect 1075 4428 1076 4432
rect 1070 4427 1076 4428
rect 1278 4432 1284 4433
rect 1278 4428 1279 4432
rect 1283 4428 1284 4432
rect 1278 4427 1284 4428
rect 1494 4432 1500 4433
rect 1494 4428 1495 4432
rect 1499 4428 1500 4432
rect 1494 4427 1500 4428
rect 658 4417 664 4418
rect 658 4413 659 4417
rect 663 4413 664 4417
rect 658 4412 664 4413
rect 842 4417 848 4418
rect 842 4413 843 4417
rect 847 4413 848 4417
rect 842 4412 848 4413
rect 1042 4417 1048 4418
rect 1042 4413 1043 4417
rect 1047 4413 1048 4417
rect 1042 4412 1048 4413
rect 1250 4417 1256 4418
rect 1250 4413 1251 4417
rect 1255 4413 1256 4417
rect 1250 4412 1256 4413
rect 1466 4417 1472 4418
rect 1466 4413 1467 4417
rect 1471 4413 1472 4417
rect 1466 4412 1472 4413
rect 578 4375 584 4376
rect 578 4371 579 4375
rect 583 4371 584 4375
rect 578 4370 584 4371
rect 660 4347 662 4412
rect 674 4407 680 4408
rect 674 4403 675 4407
rect 679 4403 680 4407
rect 674 4402 680 4403
rect 676 4376 678 4402
rect 674 4375 680 4376
rect 674 4371 675 4375
rect 679 4371 680 4375
rect 674 4370 680 4371
rect 844 4347 846 4412
rect 858 4407 864 4408
rect 858 4403 859 4407
rect 863 4403 864 4407
rect 858 4402 864 4403
rect 860 4376 862 4402
rect 858 4375 864 4376
rect 858 4371 859 4375
rect 863 4371 864 4375
rect 858 4370 864 4371
rect 1044 4347 1046 4412
rect 1058 4407 1064 4408
rect 1058 4403 1059 4407
rect 1063 4403 1064 4407
rect 1058 4402 1064 4403
rect 1060 4376 1062 4402
rect 1058 4375 1064 4376
rect 1058 4371 1059 4375
rect 1063 4371 1064 4375
rect 1058 4370 1064 4371
rect 1252 4347 1254 4412
rect 1266 4407 1272 4408
rect 1266 4403 1267 4407
rect 1271 4403 1272 4407
rect 1266 4402 1272 4403
rect 1362 4407 1368 4408
rect 1362 4403 1363 4407
rect 1367 4403 1368 4407
rect 1362 4402 1368 4403
rect 1268 4376 1270 4402
rect 1266 4375 1272 4376
rect 1266 4371 1267 4375
rect 1271 4371 1272 4375
rect 1266 4370 1272 4371
rect 111 4346 115 4347
rect 111 4341 115 4342
rect 483 4346 487 4347
rect 483 4341 487 4342
rect 659 4346 663 4347
rect 659 4341 663 4342
rect 715 4346 719 4347
rect 715 4341 719 4342
rect 843 4346 847 4347
rect 843 4341 847 4342
rect 851 4346 855 4347
rect 851 4341 855 4342
rect 987 4346 991 4347
rect 987 4341 991 4342
rect 1043 4346 1047 4347
rect 1043 4341 1047 4342
rect 1123 4346 1127 4347
rect 1123 4341 1127 4342
rect 1251 4346 1255 4347
rect 1251 4341 1255 4342
rect 1259 4346 1263 4347
rect 1259 4341 1263 4342
rect 112 4281 114 4341
rect 110 4280 116 4281
rect 716 4280 718 4341
rect 852 4280 854 4341
rect 988 4280 990 4341
rect 1124 4280 1126 4341
rect 1260 4280 1262 4341
rect 1364 4336 1366 4402
rect 1468 4347 1470 4412
rect 1564 4408 1566 4538
rect 1572 4508 1574 4569
rect 1788 4508 1790 4569
rect 1936 4509 1938 4569
rect 1934 4508 1940 4509
rect 1570 4507 1576 4508
rect 1570 4503 1571 4507
rect 1575 4503 1576 4507
rect 1570 4502 1576 4503
rect 1786 4507 1792 4508
rect 1786 4503 1787 4507
rect 1791 4503 1792 4507
rect 1934 4504 1935 4508
rect 1939 4504 1940 4508
rect 1934 4503 1940 4504
rect 1976 4503 1978 4575
rect 1996 4503 1998 4576
rect 2108 4572 2110 4710
rect 2148 4684 2150 4714
rect 2146 4683 2152 4684
rect 2146 4679 2147 4683
rect 2151 4679 2152 4683
rect 2146 4678 2152 4679
rect 2196 4676 2198 4737
rect 2322 4719 2328 4720
rect 2322 4715 2323 4719
rect 2327 4715 2328 4719
rect 2322 4714 2328 4715
rect 2324 4684 2326 4714
rect 2322 4683 2328 4684
rect 2322 4679 2323 4683
rect 2327 4679 2328 4683
rect 2322 4678 2328 4679
rect 2372 4676 2374 4737
rect 2388 4684 2390 4774
rect 2532 4743 2534 4816
rect 2546 4811 2552 4812
rect 2546 4807 2547 4811
rect 2551 4807 2552 4811
rect 2546 4806 2552 4807
rect 2548 4780 2550 4806
rect 2666 4803 2672 4804
rect 2666 4799 2667 4803
rect 2671 4799 2672 4803
rect 2666 4798 2672 4799
rect 2546 4779 2552 4780
rect 2546 4775 2547 4779
rect 2551 4775 2552 4779
rect 2546 4774 2552 4775
rect 2531 4742 2535 4743
rect 2531 4737 2535 4738
rect 2547 4742 2551 4743
rect 2547 4737 2551 4738
rect 2386 4683 2392 4684
rect 2386 4679 2387 4683
rect 2391 4679 2392 4683
rect 2386 4678 2392 4679
rect 2548 4676 2550 4737
rect 2668 4720 2670 4798
rect 2796 4743 2798 4816
rect 2964 4812 2966 4958
rect 3124 4920 3126 4981
rect 3248 4928 3250 4998
rect 3800 4987 3802 5055
rect 3838 5052 3839 5056
rect 3843 5052 3844 5056
rect 3858 5053 3859 5057
rect 3863 5053 3864 5057
rect 3858 5052 3864 5053
rect 4058 5057 4064 5058
rect 4058 5053 4059 5057
rect 4063 5053 4064 5057
rect 4058 5052 4064 5053
rect 4298 5057 4304 5058
rect 4298 5053 4299 5057
rect 4303 5053 4304 5057
rect 4298 5052 4304 5053
rect 3838 5051 3844 5052
rect 3840 4991 3842 5051
rect 3860 4991 3862 5052
rect 4060 4991 4062 5052
rect 4074 5047 4080 5048
rect 4074 5043 4075 5047
rect 4079 5043 4080 5047
rect 4074 5042 4080 5043
rect 4218 5047 4224 5048
rect 4218 5043 4219 5047
rect 4223 5043 4224 5047
rect 4218 5042 4224 5043
rect 4076 5016 4078 5042
rect 4066 5015 4072 5016
rect 4066 5011 4067 5015
rect 4071 5011 4072 5015
rect 4066 5010 4072 5011
rect 4074 5015 4080 5016
rect 4074 5011 4075 5015
rect 4079 5011 4080 5015
rect 4074 5010 4080 5011
rect 3839 4990 3843 4991
rect 3395 4986 3399 4987
rect 3395 4981 3399 4982
rect 3651 4986 3655 4987
rect 3651 4981 3655 4982
rect 3799 4986 3803 4987
rect 3839 4985 3843 4986
rect 3859 4990 3863 4991
rect 3859 4985 3863 4986
rect 3995 4990 3999 4991
rect 3995 4985 3999 4986
rect 4059 4990 4063 4991
rect 4059 4985 4063 4986
rect 3799 4981 3803 4982
rect 3246 4927 3252 4928
rect 3246 4923 3247 4927
rect 3251 4923 3252 4927
rect 3246 4922 3252 4923
rect 3396 4920 3398 4981
rect 3458 4927 3464 4928
rect 3458 4923 3459 4927
rect 3463 4923 3464 4927
rect 3458 4922 3464 4923
rect 3122 4919 3128 4920
rect 3122 4915 3123 4919
rect 3127 4915 3128 4919
rect 3122 4914 3128 4915
rect 3394 4919 3400 4920
rect 3394 4915 3395 4919
rect 3399 4915 3400 4919
rect 3394 4914 3400 4915
rect 3150 4904 3156 4905
rect 3150 4900 3151 4904
rect 3155 4900 3156 4904
rect 3150 4899 3156 4900
rect 3422 4904 3428 4905
rect 3422 4900 3423 4904
rect 3427 4900 3428 4904
rect 3422 4899 3428 4900
rect 3152 4867 3154 4899
rect 3424 4867 3426 4899
rect 3103 4866 3107 4867
rect 3103 4861 3107 4862
rect 3151 4866 3155 4867
rect 3151 4861 3155 4862
rect 3399 4866 3403 4867
rect 3399 4861 3403 4862
rect 3423 4866 3427 4867
rect 3423 4861 3427 4862
rect 3104 4837 3106 4861
rect 3400 4837 3402 4861
rect 3102 4836 3108 4837
rect 3102 4832 3103 4836
rect 3107 4832 3108 4836
rect 3102 4831 3108 4832
rect 3398 4836 3404 4837
rect 3398 4832 3399 4836
rect 3403 4832 3404 4836
rect 3398 4831 3404 4832
rect 3074 4821 3080 4822
rect 3074 4817 3075 4821
rect 3079 4817 3080 4821
rect 3074 4816 3080 4817
rect 3370 4821 3376 4822
rect 3370 4817 3371 4821
rect 3375 4817 3376 4821
rect 3370 4816 3376 4817
rect 2810 4811 2816 4812
rect 2810 4807 2811 4811
rect 2815 4807 2816 4811
rect 2810 4806 2816 4807
rect 2962 4811 2968 4812
rect 2962 4807 2963 4811
rect 2967 4807 2968 4811
rect 2962 4806 2968 4807
rect 2812 4780 2814 4806
rect 2810 4779 2816 4780
rect 2810 4775 2811 4779
rect 2815 4775 2816 4779
rect 2810 4774 2816 4775
rect 3076 4743 3078 4816
rect 3372 4743 3374 4816
rect 3460 4780 3462 4922
rect 3652 4920 3654 4981
rect 3790 4967 3796 4968
rect 3790 4963 3791 4967
rect 3795 4963 3796 4967
rect 3790 4962 3796 4963
rect 3738 4959 3744 4960
rect 3738 4955 3739 4959
rect 3743 4955 3744 4959
rect 3738 4954 3744 4955
rect 3650 4919 3656 4920
rect 3650 4915 3651 4919
rect 3655 4915 3656 4919
rect 3650 4914 3656 4915
rect 3678 4904 3684 4905
rect 3678 4900 3679 4904
rect 3683 4900 3684 4904
rect 3678 4899 3684 4900
rect 3680 4867 3682 4899
rect 3679 4866 3683 4867
rect 3679 4861 3683 4862
rect 3680 4837 3682 4861
rect 3678 4836 3684 4837
rect 3678 4832 3679 4836
rect 3683 4832 3684 4836
rect 3678 4831 3684 4832
rect 3650 4821 3656 4822
rect 3650 4817 3651 4821
rect 3655 4817 3656 4821
rect 3650 4816 3656 4817
rect 3458 4779 3464 4780
rect 3458 4775 3459 4779
rect 3463 4775 3464 4779
rect 3458 4774 3464 4775
rect 3652 4743 3654 4816
rect 3740 4812 3742 4954
rect 3792 4928 3794 4962
rect 3790 4927 3796 4928
rect 3790 4923 3791 4927
rect 3795 4923 3796 4927
rect 3790 4922 3796 4923
rect 3800 4921 3802 4981
rect 3840 4925 3842 4985
rect 3838 4924 3844 4925
rect 3860 4924 3862 4985
rect 3986 4967 3992 4968
rect 3986 4963 3987 4967
rect 3991 4963 3992 4967
rect 3986 4962 3992 4963
rect 3988 4932 3990 4962
rect 3986 4931 3992 4932
rect 3986 4927 3987 4931
rect 3991 4927 3992 4931
rect 3986 4926 3992 4927
rect 3996 4924 3998 4985
rect 4068 4932 4070 5010
rect 4131 4990 4135 4991
rect 4131 4985 4135 4986
rect 4066 4931 4072 4932
rect 4066 4927 4067 4931
rect 4071 4927 4072 4931
rect 4066 4926 4072 4927
rect 4132 4924 4134 4985
rect 4220 4964 4222 5042
rect 4300 4991 4302 5052
rect 4428 5048 4430 5194
rect 4436 5156 4438 5217
rect 4596 5156 4598 5217
rect 4604 5164 4606 5258
rect 4772 5223 4774 5300
rect 4946 5295 4952 5296
rect 4946 5291 4947 5295
rect 4951 5291 4952 5295
rect 4946 5290 4952 5291
rect 4948 5264 4950 5290
rect 4946 5263 4952 5264
rect 4946 5259 4947 5263
rect 4951 5259 4952 5263
rect 4946 5258 4952 5259
rect 4956 5223 4958 5300
rect 5148 5223 5150 5300
rect 5200 5264 5202 5406
rect 5664 5405 5666 5465
rect 5662 5404 5668 5405
rect 5662 5400 5663 5404
rect 5667 5400 5668 5404
rect 5662 5399 5668 5400
rect 5662 5387 5668 5388
rect 5662 5383 5663 5387
rect 5667 5383 5668 5387
rect 5662 5382 5668 5383
rect 5664 5351 5666 5382
rect 5663 5350 5667 5351
rect 5663 5345 5667 5346
rect 5664 5322 5666 5345
rect 5662 5321 5668 5322
rect 5662 5317 5663 5321
rect 5667 5317 5668 5321
rect 5662 5316 5668 5317
rect 5662 5304 5668 5305
rect 5662 5300 5663 5304
rect 5667 5300 5668 5304
rect 5662 5299 5668 5300
rect 5198 5263 5204 5264
rect 5198 5259 5199 5263
rect 5203 5259 5204 5263
rect 5198 5258 5204 5259
rect 5664 5223 5666 5299
rect 4755 5222 4759 5223
rect 4755 5217 4759 5218
rect 4771 5222 4775 5223
rect 4771 5217 4775 5218
rect 4915 5222 4919 5223
rect 4915 5217 4919 5218
rect 4955 5222 4959 5223
rect 4955 5217 4959 5218
rect 5067 5222 5071 5223
rect 5067 5217 5071 5218
rect 5147 5222 5151 5223
rect 5147 5217 5151 5218
rect 5219 5222 5223 5223
rect 5219 5217 5223 5218
rect 5379 5222 5383 5223
rect 5379 5217 5383 5218
rect 5515 5222 5519 5223
rect 5515 5217 5519 5218
rect 5663 5222 5667 5223
rect 5663 5217 5667 5218
rect 4602 5163 4608 5164
rect 4602 5159 4603 5163
rect 4607 5159 4608 5163
rect 4602 5158 4608 5159
rect 4756 5156 4758 5217
rect 4916 5156 4918 5217
rect 5068 5156 5070 5217
rect 5220 5156 5222 5217
rect 5380 5156 5382 5217
rect 5516 5156 5518 5217
rect 5602 5163 5608 5164
rect 5602 5159 5603 5163
rect 5607 5159 5608 5163
rect 5602 5158 5608 5159
rect 4434 5155 4440 5156
rect 4434 5151 4435 5155
rect 4439 5151 4440 5155
rect 4434 5150 4440 5151
rect 4594 5155 4600 5156
rect 4594 5151 4595 5155
rect 4599 5151 4600 5155
rect 4594 5150 4600 5151
rect 4754 5155 4760 5156
rect 4754 5151 4755 5155
rect 4759 5151 4760 5155
rect 4754 5150 4760 5151
rect 4914 5155 4920 5156
rect 4914 5151 4915 5155
rect 4919 5151 4920 5155
rect 4914 5150 4920 5151
rect 5066 5155 5072 5156
rect 5066 5151 5067 5155
rect 5071 5151 5072 5155
rect 5066 5150 5072 5151
rect 5218 5155 5224 5156
rect 5218 5151 5219 5155
rect 5223 5151 5224 5155
rect 5218 5150 5224 5151
rect 5378 5155 5384 5156
rect 5378 5151 5379 5155
rect 5383 5151 5384 5155
rect 5378 5150 5384 5151
rect 5514 5155 5520 5156
rect 5514 5151 5515 5155
rect 5519 5151 5520 5155
rect 5514 5150 5520 5151
rect 4462 5140 4468 5141
rect 4462 5136 4463 5140
rect 4467 5136 4468 5140
rect 4462 5135 4468 5136
rect 4622 5140 4628 5141
rect 4622 5136 4623 5140
rect 4627 5136 4628 5140
rect 4622 5135 4628 5136
rect 4782 5140 4788 5141
rect 4782 5136 4783 5140
rect 4787 5136 4788 5140
rect 4782 5135 4788 5136
rect 4942 5140 4948 5141
rect 4942 5136 4943 5140
rect 4947 5136 4948 5140
rect 4942 5135 4948 5136
rect 5094 5140 5100 5141
rect 5094 5136 5095 5140
rect 5099 5136 5100 5140
rect 5094 5135 5100 5136
rect 5246 5140 5252 5141
rect 5246 5136 5247 5140
rect 5251 5136 5252 5140
rect 5246 5135 5252 5136
rect 5406 5140 5412 5141
rect 5406 5136 5407 5140
rect 5411 5136 5412 5140
rect 5406 5135 5412 5136
rect 5542 5140 5548 5141
rect 5542 5136 5543 5140
rect 5547 5136 5548 5140
rect 5542 5135 5548 5136
rect 4464 5103 4466 5135
rect 4624 5103 4626 5135
rect 4784 5103 4786 5135
rect 4944 5103 4946 5135
rect 5096 5103 5098 5135
rect 5248 5103 5250 5135
rect 5408 5103 5410 5135
rect 5544 5103 5546 5135
rect 4463 5102 4467 5103
rect 4463 5097 4467 5098
rect 4567 5102 4571 5103
rect 4567 5097 4571 5098
rect 4623 5102 4627 5103
rect 4623 5097 4627 5098
rect 4783 5102 4787 5103
rect 4783 5097 4787 5098
rect 4815 5102 4819 5103
rect 4815 5097 4819 5098
rect 4943 5102 4947 5103
rect 4943 5097 4947 5098
rect 5063 5102 5067 5103
rect 5063 5097 5067 5098
rect 5095 5102 5099 5103
rect 5095 5097 5099 5098
rect 5247 5102 5251 5103
rect 5247 5097 5251 5098
rect 5311 5102 5315 5103
rect 5311 5097 5315 5098
rect 5407 5102 5411 5103
rect 5407 5097 5411 5098
rect 5543 5102 5547 5103
rect 5543 5097 5547 5098
rect 4568 5073 4570 5097
rect 4816 5073 4818 5097
rect 5064 5073 5066 5097
rect 5312 5073 5314 5097
rect 5544 5073 5546 5097
rect 4566 5072 4572 5073
rect 4566 5068 4567 5072
rect 4571 5068 4572 5072
rect 4566 5067 4572 5068
rect 4814 5072 4820 5073
rect 4814 5068 4815 5072
rect 4819 5068 4820 5072
rect 4814 5067 4820 5068
rect 5062 5072 5068 5073
rect 5062 5068 5063 5072
rect 5067 5068 5068 5072
rect 5062 5067 5068 5068
rect 5310 5072 5316 5073
rect 5310 5068 5311 5072
rect 5315 5068 5316 5072
rect 5310 5067 5316 5068
rect 5542 5072 5548 5073
rect 5542 5068 5543 5072
rect 5547 5068 5548 5072
rect 5542 5067 5548 5068
rect 4538 5057 4544 5058
rect 4538 5053 4539 5057
rect 4543 5053 4544 5057
rect 4538 5052 4544 5053
rect 4786 5057 4792 5058
rect 4786 5053 4787 5057
rect 4791 5053 4792 5057
rect 4786 5052 4792 5053
rect 5034 5057 5040 5058
rect 5034 5053 5035 5057
rect 5039 5053 5040 5057
rect 5034 5052 5040 5053
rect 5282 5057 5288 5058
rect 5282 5053 5283 5057
rect 5287 5053 5288 5057
rect 5282 5052 5288 5053
rect 5514 5057 5520 5058
rect 5514 5053 5515 5057
rect 5519 5053 5520 5057
rect 5514 5052 5520 5053
rect 4426 5047 4432 5048
rect 4426 5043 4427 5047
rect 4431 5043 4432 5047
rect 4426 5042 4432 5043
rect 4458 5047 4464 5048
rect 4458 5043 4459 5047
rect 4463 5043 4464 5047
rect 4458 5042 4464 5043
rect 4460 5016 4462 5042
rect 4458 5015 4464 5016
rect 4458 5011 4459 5015
rect 4463 5011 4464 5015
rect 4458 5010 4464 5011
rect 4540 4991 4542 5052
rect 4682 5047 4688 5048
rect 4682 5043 4683 5047
rect 4687 5043 4688 5047
rect 4682 5042 4688 5043
rect 4684 5016 4686 5042
rect 4682 5015 4688 5016
rect 4682 5011 4683 5015
rect 4687 5011 4688 5015
rect 4682 5010 4688 5011
rect 4788 4991 4790 5052
rect 4874 5015 4880 5016
rect 4874 5011 4875 5015
rect 4879 5011 4880 5015
rect 4874 5010 4880 5011
rect 4267 4990 4271 4991
rect 4267 4985 4271 4986
rect 4299 4990 4303 4991
rect 4299 4985 4303 4986
rect 4403 4990 4407 4991
rect 4403 4985 4407 4986
rect 4539 4990 4543 4991
rect 4539 4985 4543 4986
rect 4675 4990 4679 4991
rect 4675 4985 4679 4986
rect 4787 4990 4791 4991
rect 4787 4985 4791 4986
rect 4811 4990 4815 4991
rect 4811 4985 4815 4986
rect 4218 4963 4224 4964
rect 4218 4959 4219 4963
rect 4223 4959 4224 4963
rect 4218 4958 4224 4959
rect 4268 4924 4270 4985
rect 4404 4924 4406 4985
rect 4540 4924 4542 4985
rect 4676 4924 4678 4985
rect 4802 4967 4808 4968
rect 4802 4963 4803 4967
rect 4807 4963 4808 4967
rect 4802 4962 4808 4963
rect 4804 4932 4806 4962
rect 4802 4931 4808 4932
rect 4802 4927 4803 4931
rect 4807 4927 4808 4931
rect 4802 4926 4808 4927
rect 4812 4924 4814 4985
rect 4876 4973 4878 5010
rect 5036 4991 5038 5052
rect 5122 5039 5128 5040
rect 5122 5035 5123 5039
rect 5127 5035 5128 5039
rect 5122 5034 5128 5035
rect 5124 5016 5126 5034
rect 5122 5015 5128 5016
rect 5122 5011 5123 5015
rect 5127 5011 5128 5015
rect 5122 5010 5128 5011
rect 5284 4991 5286 5052
rect 5298 5047 5304 5048
rect 5298 5043 5299 5047
rect 5303 5043 5304 5047
rect 5298 5042 5304 5043
rect 5370 5047 5376 5048
rect 5370 5043 5371 5047
rect 5375 5043 5376 5047
rect 5370 5042 5376 5043
rect 5300 5016 5302 5042
rect 5298 5015 5304 5016
rect 5298 5011 5299 5015
rect 5303 5011 5304 5015
rect 5298 5010 5304 5011
rect 4947 4990 4951 4991
rect 4947 4985 4951 4986
rect 5035 4990 5039 4991
rect 5035 4985 5039 4986
rect 5083 4990 5087 4991
rect 5083 4985 5087 4986
rect 5227 4990 5231 4991
rect 5227 4985 5231 4986
rect 5283 4990 5287 4991
rect 5283 4985 5287 4986
rect 4875 4972 4879 4973
rect 4875 4967 4879 4968
rect 4948 4924 4950 4985
rect 5084 4924 5086 4985
rect 5210 4967 5216 4968
rect 5210 4963 5211 4967
rect 5215 4963 5216 4967
rect 5210 4962 5216 4963
rect 5212 4932 5214 4962
rect 5210 4931 5216 4932
rect 5210 4927 5211 4931
rect 5215 4927 5216 4931
rect 5210 4926 5216 4927
rect 5228 4924 5230 4985
rect 5239 4972 5243 4973
rect 5372 4968 5374 5042
rect 5516 4991 5518 5052
rect 5604 5016 5606 5158
rect 5664 5157 5666 5217
rect 5662 5156 5668 5157
rect 5662 5152 5663 5156
rect 5667 5152 5668 5156
rect 5662 5151 5668 5152
rect 5662 5139 5668 5140
rect 5662 5135 5663 5139
rect 5667 5135 5668 5139
rect 5662 5134 5668 5135
rect 5664 5103 5666 5134
rect 5663 5102 5667 5103
rect 5663 5097 5667 5098
rect 5664 5074 5666 5097
rect 5662 5073 5668 5074
rect 5662 5069 5663 5073
rect 5667 5069 5668 5073
rect 5662 5068 5668 5069
rect 5662 5056 5668 5057
rect 5662 5052 5663 5056
rect 5667 5052 5668 5056
rect 5662 5051 5668 5052
rect 5602 5015 5608 5016
rect 5602 5011 5603 5015
rect 5607 5011 5608 5015
rect 5602 5010 5608 5011
rect 5664 4991 5666 5051
rect 5379 4990 5383 4991
rect 5379 4985 5383 4986
rect 5515 4990 5519 4991
rect 5515 4985 5519 4986
rect 5663 4990 5667 4991
rect 5663 4985 5667 4986
rect 5239 4967 5243 4968
rect 5370 4967 5376 4968
rect 5240 4932 5242 4967
rect 5370 4963 5371 4967
rect 5375 4963 5376 4967
rect 5370 4962 5376 4963
rect 5238 4931 5244 4932
rect 5238 4927 5239 4931
rect 5243 4927 5244 4931
rect 5238 4926 5244 4927
rect 5380 4924 5382 4985
rect 5516 4924 5518 4985
rect 5602 4931 5608 4932
rect 5602 4927 5603 4931
rect 5607 4927 5608 4931
rect 5602 4926 5608 4927
rect 3798 4920 3804 4921
rect 3798 4916 3799 4920
rect 3803 4916 3804 4920
rect 3838 4920 3839 4924
rect 3843 4920 3844 4924
rect 3838 4919 3844 4920
rect 3858 4923 3864 4924
rect 3858 4919 3859 4923
rect 3863 4919 3864 4923
rect 3858 4918 3864 4919
rect 3994 4923 4000 4924
rect 3994 4919 3995 4923
rect 3999 4919 4000 4923
rect 3994 4918 4000 4919
rect 4130 4923 4136 4924
rect 4130 4919 4131 4923
rect 4135 4919 4136 4923
rect 4130 4918 4136 4919
rect 4266 4923 4272 4924
rect 4266 4919 4267 4923
rect 4271 4919 4272 4923
rect 4266 4918 4272 4919
rect 4402 4923 4408 4924
rect 4402 4919 4403 4923
rect 4407 4919 4408 4923
rect 4402 4918 4408 4919
rect 4538 4923 4544 4924
rect 4538 4919 4539 4923
rect 4543 4919 4544 4923
rect 4538 4918 4544 4919
rect 4674 4923 4680 4924
rect 4674 4919 4675 4923
rect 4679 4919 4680 4923
rect 4674 4918 4680 4919
rect 4810 4923 4816 4924
rect 4810 4919 4811 4923
rect 4815 4919 4816 4923
rect 4810 4918 4816 4919
rect 4946 4923 4952 4924
rect 4946 4919 4947 4923
rect 4951 4919 4952 4923
rect 4946 4918 4952 4919
rect 5082 4923 5088 4924
rect 5082 4919 5083 4923
rect 5087 4919 5088 4923
rect 5082 4918 5088 4919
rect 5226 4923 5232 4924
rect 5226 4919 5227 4923
rect 5231 4919 5232 4923
rect 5226 4918 5232 4919
rect 5378 4923 5384 4924
rect 5378 4919 5379 4923
rect 5383 4919 5384 4923
rect 5378 4918 5384 4919
rect 5514 4923 5520 4924
rect 5514 4919 5515 4923
rect 5519 4919 5520 4923
rect 5514 4918 5520 4919
rect 3798 4915 3804 4916
rect 3886 4908 3892 4909
rect 3838 4907 3844 4908
rect 3798 4903 3804 4904
rect 3798 4899 3799 4903
rect 3803 4899 3804 4903
rect 3838 4903 3839 4907
rect 3843 4903 3844 4907
rect 3886 4904 3887 4908
rect 3891 4904 3892 4908
rect 3886 4903 3892 4904
rect 4022 4908 4028 4909
rect 4022 4904 4023 4908
rect 4027 4904 4028 4908
rect 4022 4903 4028 4904
rect 4158 4908 4164 4909
rect 4158 4904 4159 4908
rect 4163 4904 4164 4908
rect 4158 4903 4164 4904
rect 4294 4908 4300 4909
rect 4294 4904 4295 4908
rect 4299 4904 4300 4908
rect 4294 4903 4300 4904
rect 4430 4908 4436 4909
rect 4430 4904 4431 4908
rect 4435 4904 4436 4908
rect 4430 4903 4436 4904
rect 4566 4908 4572 4909
rect 4566 4904 4567 4908
rect 4571 4904 4572 4908
rect 4566 4903 4572 4904
rect 4702 4908 4708 4909
rect 4702 4904 4703 4908
rect 4707 4904 4708 4908
rect 4702 4903 4708 4904
rect 4838 4908 4844 4909
rect 4838 4904 4839 4908
rect 4843 4904 4844 4908
rect 4838 4903 4844 4904
rect 4974 4908 4980 4909
rect 4974 4904 4975 4908
rect 4979 4904 4980 4908
rect 4974 4903 4980 4904
rect 5110 4908 5116 4909
rect 5110 4904 5111 4908
rect 5115 4904 5116 4908
rect 5110 4903 5116 4904
rect 5254 4908 5260 4909
rect 5254 4904 5255 4908
rect 5259 4904 5260 4908
rect 5254 4903 5260 4904
rect 5406 4908 5412 4909
rect 5406 4904 5407 4908
rect 5411 4904 5412 4908
rect 5406 4903 5412 4904
rect 5542 4908 5548 4909
rect 5542 4904 5543 4908
rect 5547 4904 5548 4908
rect 5542 4903 5548 4904
rect 3838 4902 3844 4903
rect 3798 4898 3804 4899
rect 3800 4867 3802 4898
rect 3799 4866 3803 4867
rect 3799 4861 3803 4862
rect 3800 4838 3802 4861
rect 3798 4837 3804 4838
rect 3798 4833 3799 4837
rect 3803 4833 3804 4837
rect 3798 4832 3804 4833
rect 3798 4820 3804 4821
rect 3798 4816 3799 4820
rect 3803 4816 3804 4820
rect 3798 4815 3804 4816
rect 3738 4811 3744 4812
rect 3738 4807 3739 4811
rect 3743 4807 3744 4811
rect 3738 4806 3744 4807
rect 3738 4779 3744 4780
rect 3738 4775 3739 4779
rect 3743 4775 3744 4779
rect 3738 4774 3744 4775
rect 3740 4748 3742 4774
rect 3738 4747 3744 4748
rect 3738 4743 3739 4747
rect 3743 4743 3744 4747
rect 3800 4743 3802 4815
rect 3840 4803 3842 4902
rect 3888 4803 3890 4903
rect 4024 4803 4026 4903
rect 4160 4803 4162 4903
rect 4296 4803 4298 4903
rect 4432 4803 4434 4903
rect 4568 4803 4570 4903
rect 4704 4803 4706 4903
rect 4840 4803 4842 4903
rect 4976 4803 4978 4903
rect 5112 4803 5114 4903
rect 5256 4803 5258 4903
rect 5408 4803 5410 4903
rect 5544 4803 5546 4903
rect 3839 4802 3843 4803
rect 3839 4797 3843 4798
rect 3887 4802 3891 4803
rect 3887 4797 3891 4798
rect 4023 4802 4027 4803
rect 4023 4797 4027 4798
rect 4071 4802 4075 4803
rect 4071 4797 4075 4798
rect 4159 4802 4163 4803
rect 4159 4797 4163 4798
rect 4295 4802 4299 4803
rect 4295 4797 4299 4798
rect 4431 4802 4435 4803
rect 4431 4797 4435 4798
rect 4535 4802 4539 4803
rect 4535 4797 4539 4798
rect 4567 4802 4571 4803
rect 4567 4797 4571 4798
rect 4703 4802 4707 4803
rect 4703 4797 4707 4798
rect 4783 4802 4787 4803
rect 4783 4797 4787 4798
rect 4839 4802 4843 4803
rect 4839 4797 4843 4798
rect 4975 4802 4979 4803
rect 4975 4797 4979 4798
rect 5039 4802 5043 4803
rect 5039 4797 5043 4798
rect 5111 4802 5115 4803
rect 5111 4797 5115 4798
rect 5255 4802 5259 4803
rect 5255 4797 5259 4798
rect 5303 4802 5307 4803
rect 5303 4797 5307 4798
rect 5407 4802 5411 4803
rect 5407 4797 5411 4798
rect 5543 4802 5547 4803
rect 5543 4797 5547 4798
rect 3840 4774 3842 4797
rect 3838 4773 3844 4774
rect 3888 4773 3890 4797
rect 4072 4773 4074 4797
rect 4296 4773 4298 4797
rect 4536 4773 4538 4797
rect 4784 4773 4786 4797
rect 5040 4773 5042 4797
rect 5304 4773 5306 4797
rect 5544 4773 5546 4797
rect 3838 4769 3839 4773
rect 3843 4769 3844 4773
rect 3838 4768 3844 4769
rect 3886 4772 3892 4773
rect 3886 4768 3887 4772
rect 3891 4768 3892 4772
rect 3886 4767 3892 4768
rect 4070 4772 4076 4773
rect 4070 4768 4071 4772
rect 4075 4768 4076 4772
rect 4070 4767 4076 4768
rect 4294 4772 4300 4773
rect 4294 4768 4295 4772
rect 4299 4768 4300 4772
rect 4294 4767 4300 4768
rect 4534 4772 4540 4773
rect 4534 4768 4535 4772
rect 4539 4768 4540 4772
rect 4534 4767 4540 4768
rect 4782 4772 4788 4773
rect 4782 4768 4783 4772
rect 4787 4768 4788 4772
rect 4782 4767 4788 4768
rect 5038 4772 5044 4773
rect 5038 4768 5039 4772
rect 5043 4768 5044 4772
rect 5038 4767 5044 4768
rect 5302 4772 5308 4773
rect 5302 4768 5303 4772
rect 5307 4768 5308 4772
rect 5302 4767 5308 4768
rect 5542 4772 5548 4773
rect 5542 4768 5543 4772
rect 5547 4768 5548 4772
rect 5542 4767 5548 4768
rect 3858 4757 3864 4758
rect 3838 4756 3844 4757
rect 3838 4752 3839 4756
rect 3843 4752 3844 4756
rect 3858 4753 3859 4757
rect 3863 4753 3864 4757
rect 3858 4752 3864 4753
rect 4042 4757 4048 4758
rect 4042 4753 4043 4757
rect 4047 4753 4048 4757
rect 4042 4752 4048 4753
rect 4266 4757 4272 4758
rect 4266 4753 4267 4757
rect 4271 4753 4272 4757
rect 4266 4752 4272 4753
rect 4506 4757 4512 4758
rect 4506 4753 4507 4757
rect 4511 4753 4512 4757
rect 4506 4752 4512 4753
rect 4754 4757 4760 4758
rect 4754 4753 4755 4757
rect 4759 4753 4760 4757
rect 4754 4752 4760 4753
rect 5010 4757 5016 4758
rect 5010 4753 5011 4757
rect 5015 4753 5016 4757
rect 5010 4752 5016 4753
rect 5274 4757 5280 4758
rect 5274 4753 5275 4757
rect 5279 4753 5280 4757
rect 5274 4752 5280 4753
rect 5514 4757 5520 4758
rect 5514 4753 5515 4757
rect 5519 4753 5520 4757
rect 5514 4752 5520 4753
rect 3838 4751 3844 4752
rect 2723 4742 2727 4743
rect 2723 4737 2727 4738
rect 2795 4742 2799 4743
rect 2795 4737 2799 4738
rect 3075 4742 3079 4743
rect 3075 4737 3079 4738
rect 3371 4742 3375 4743
rect 3371 4737 3375 4738
rect 3651 4742 3655 4743
rect 3738 4742 3744 4743
rect 3799 4742 3803 4743
rect 3651 4737 3655 4738
rect 3799 4737 3803 4738
rect 2666 4719 2672 4720
rect 2666 4715 2667 4719
rect 2671 4715 2672 4719
rect 2666 4714 2672 4715
rect 2674 4719 2680 4720
rect 2674 4715 2675 4719
rect 2679 4715 2680 4719
rect 2674 4714 2680 4715
rect 2676 4684 2678 4714
rect 2674 4683 2680 4684
rect 2674 4679 2675 4683
rect 2679 4679 2680 4683
rect 2674 4678 2680 4679
rect 2724 4676 2726 4737
rect 2834 4683 2840 4684
rect 2834 4679 2835 4683
rect 2839 4679 2840 4683
rect 2834 4678 2840 4679
rect 2194 4675 2200 4676
rect 2194 4671 2195 4675
rect 2199 4671 2200 4675
rect 2194 4670 2200 4671
rect 2370 4675 2376 4676
rect 2370 4671 2371 4675
rect 2375 4671 2376 4675
rect 2370 4670 2376 4671
rect 2546 4675 2552 4676
rect 2546 4671 2547 4675
rect 2551 4671 2552 4675
rect 2546 4670 2552 4671
rect 2722 4675 2728 4676
rect 2722 4671 2723 4675
rect 2727 4671 2728 4675
rect 2722 4670 2728 4671
rect 2222 4660 2228 4661
rect 2222 4656 2223 4660
rect 2227 4656 2228 4660
rect 2222 4655 2228 4656
rect 2398 4660 2404 4661
rect 2398 4656 2399 4660
rect 2403 4656 2404 4660
rect 2398 4655 2404 4656
rect 2574 4660 2580 4661
rect 2574 4656 2575 4660
rect 2579 4656 2580 4660
rect 2574 4655 2580 4656
rect 2750 4660 2756 4661
rect 2750 4656 2751 4660
rect 2755 4656 2756 4660
rect 2750 4655 2756 4656
rect 2224 4627 2226 4655
rect 2400 4627 2402 4655
rect 2576 4627 2578 4655
rect 2752 4627 2754 4655
rect 2223 4626 2227 4627
rect 2223 4621 2227 4622
rect 2263 4626 2267 4627
rect 2263 4621 2267 4622
rect 2399 4626 2403 4627
rect 2399 4621 2403 4622
rect 2527 4626 2531 4627
rect 2527 4621 2531 4622
rect 2575 4626 2579 4627
rect 2575 4621 2579 4622
rect 2751 4626 2755 4627
rect 2751 4621 2755 4622
rect 2775 4626 2779 4627
rect 2775 4621 2779 4622
rect 2264 4597 2266 4621
rect 2528 4597 2530 4621
rect 2776 4597 2778 4621
rect 2262 4596 2268 4597
rect 2262 4592 2263 4596
rect 2267 4592 2268 4596
rect 2262 4591 2268 4592
rect 2526 4596 2532 4597
rect 2526 4592 2527 4596
rect 2531 4592 2532 4596
rect 2526 4591 2532 4592
rect 2774 4596 2780 4597
rect 2774 4592 2775 4596
rect 2779 4592 2780 4596
rect 2774 4591 2780 4592
rect 2234 4581 2240 4582
rect 2234 4577 2235 4581
rect 2239 4577 2240 4581
rect 2234 4576 2240 4577
rect 2498 4581 2504 4582
rect 2498 4577 2499 4581
rect 2503 4577 2504 4581
rect 2498 4576 2504 4577
rect 2746 4581 2752 4582
rect 2746 4577 2747 4581
rect 2751 4577 2752 4581
rect 2746 4576 2752 4577
rect 2106 4571 2112 4572
rect 2106 4567 2107 4571
rect 2111 4567 2112 4571
rect 2106 4566 2112 4567
rect 2010 4539 2016 4540
rect 2010 4535 2011 4539
rect 2015 4535 2016 4539
rect 2010 4534 2016 4535
rect 2012 4516 2014 4534
rect 2010 4515 2016 4516
rect 2010 4511 2011 4515
rect 2015 4511 2016 4515
rect 2010 4510 2016 4511
rect 2236 4503 2238 4576
rect 2322 4563 2328 4564
rect 2322 4559 2323 4563
rect 2327 4559 2328 4563
rect 2322 4558 2328 4559
rect 2324 4540 2326 4558
rect 2322 4539 2328 4540
rect 2322 4535 2323 4539
rect 2327 4535 2328 4539
rect 2322 4534 2328 4535
rect 2500 4503 2502 4576
rect 2514 4571 2520 4572
rect 2514 4567 2515 4571
rect 2519 4567 2520 4571
rect 2514 4566 2520 4567
rect 2618 4571 2624 4572
rect 2618 4567 2619 4571
rect 2623 4567 2624 4571
rect 2618 4566 2624 4567
rect 2516 4540 2518 4566
rect 2514 4539 2520 4540
rect 2514 4535 2515 4539
rect 2519 4535 2520 4539
rect 2514 4534 2520 4535
rect 1786 4502 1792 4503
rect 1975 4502 1979 4503
rect 1975 4497 1979 4498
rect 1995 4502 1999 4503
rect 1995 4497 1999 4498
rect 2235 4502 2239 4503
rect 2235 4497 2239 4498
rect 2267 4502 2271 4503
rect 2267 4497 2271 4498
rect 2499 4502 2503 4503
rect 2499 4497 2503 4498
rect 2515 4502 2519 4503
rect 2515 4497 2519 4498
rect 1598 4492 1604 4493
rect 1598 4488 1599 4492
rect 1603 4488 1604 4492
rect 1598 4487 1604 4488
rect 1814 4492 1820 4493
rect 1814 4488 1815 4492
rect 1819 4488 1820 4492
rect 1814 4487 1820 4488
rect 1934 4491 1940 4492
rect 1934 4487 1935 4491
rect 1939 4487 1940 4491
rect 1600 4463 1602 4487
rect 1816 4463 1818 4487
rect 1934 4486 1940 4487
rect 1936 4463 1938 4486
rect 1599 4462 1603 4463
rect 1599 4457 1603 4458
rect 1719 4462 1723 4463
rect 1719 4457 1723 4458
rect 1815 4462 1819 4463
rect 1815 4457 1819 4458
rect 1935 4462 1939 4463
rect 1935 4457 1939 4458
rect 1720 4433 1722 4457
rect 1936 4434 1938 4457
rect 1976 4437 1978 4497
rect 1974 4436 1980 4437
rect 2268 4436 2270 4497
rect 2494 4479 2500 4480
rect 2494 4475 2495 4479
rect 2499 4475 2500 4479
rect 2494 4474 2500 4475
rect 2496 4444 2498 4474
rect 2390 4443 2396 4444
rect 2390 4439 2391 4443
rect 2395 4439 2396 4443
rect 2390 4438 2396 4439
rect 2494 4443 2500 4444
rect 2494 4439 2495 4443
rect 2499 4439 2500 4443
rect 2494 4438 2500 4439
rect 1934 4433 1940 4434
rect 1718 4432 1724 4433
rect 1718 4428 1719 4432
rect 1723 4428 1724 4432
rect 1934 4429 1935 4433
rect 1939 4429 1940 4433
rect 1974 4432 1975 4436
rect 1979 4432 1980 4436
rect 1974 4431 1980 4432
rect 2266 4435 2272 4436
rect 2266 4431 2267 4435
rect 2271 4431 2272 4435
rect 2266 4430 2272 4431
rect 1934 4428 1940 4429
rect 1718 4427 1724 4428
rect 2294 4420 2300 4421
rect 1974 4419 1980 4420
rect 1690 4417 1696 4418
rect 1690 4413 1691 4417
rect 1695 4413 1696 4417
rect 1690 4412 1696 4413
rect 1934 4416 1940 4417
rect 1934 4412 1935 4416
rect 1939 4412 1940 4416
rect 1974 4415 1975 4419
rect 1979 4415 1980 4419
rect 2294 4416 2295 4420
rect 2299 4416 2300 4420
rect 2294 4415 2300 4416
rect 1974 4414 1980 4415
rect 1562 4407 1568 4408
rect 1562 4403 1563 4407
rect 1567 4403 1568 4407
rect 1562 4402 1568 4403
rect 1610 4407 1616 4408
rect 1610 4403 1611 4407
rect 1615 4403 1616 4407
rect 1610 4402 1616 4403
rect 1612 4376 1614 4402
rect 1610 4375 1616 4376
rect 1610 4371 1611 4375
rect 1615 4371 1616 4375
rect 1610 4370 1616 4371
rect 1692 4347 1694 4412
rect 1934 4411 1940 4412
rect 1778 4375 1784 4376
rect 1778 4371 1779 4375
rect 1783 4371 1784 4375
rect 1778 4370 1784 4371
rect 1395 4346 1399 4347
rect 1395 4341 1399 4342
rect 1467 4346 1471 4347
rect 1467 4341 1471 4342
rect 1531 4346 1535 4347
rect 1531 4341 1535 4342
rect 1667 4346 1671 4347
rect 1667 4341 1671 4342
rect 1691 4346 1695 4347
rect 1691 4341 1695 4342
rect 1362 4335 1368 4336
rect 1362 4331 1363 4335
rect 1367 4331 1368 4335
rect 1362 4330 1368 4331
rect 1330 4287 1336 4288
rect 1330 4283 1331 4287
rect 1335 4283 1336 4287
rect 1330 4282 1336 4283
rect 110 4276 111 4280
rect 115 4276 116 4280
rect 110 4275 116 4276
rect 714 4279 720 4280
rect 714 4275 715 4279
rect 719 4275 720 4279
rect 714 4274 720 4275
rect 850 4279 856 4280
rect 850 4275 851 4279
rect 855 4275 856 4279
rect 850 4274 856 4275
rect 986 4279 992 4280
rect 986 4275 987 4279
rect 991 4275 992 4279
rect 986 4274 992 4275
rect 1122 4279 1128 4280
rect 1122 4275 1123 4279
rect 1127 4275 1128 4279
rect 1122 4274 1128 4275
rect 1258 4279 1264 4280
rect 1258 4275 1259 4279
rect 1263 4275 1264 4279
rect 1258 4274 1264 4275
rect 742 4264 748 4265
rect 110 4263 116 4264
rect 110 4259 111 4263
rect 115 4259 116 4263
rect 742 4260 743 4264
rect 747 4260 748 4264
rect 742 4259 748 4260
rect 878 4264 884 4265
rect 878 4260 879 4264
rect 883 4260 884 4264
rect 878 4259 884 4260
rect 1014 4264 1020 4265
rect 1014 4260 1015 4264
rect 1019 4260 1020 4264
rect 1014 4259 1020 4260
rect 1150 4264 1156 4265
rect 1150 4260 1151 4264
rect 1155 4260 1156 4264
rect 1150 4259 1156 4260
rect 1286 4264 1292 4265
rect 1286 4260 1287 4264
rect 1291 4260 1292 4264
rect 1286 4259 1292 4260
rect 110 4258 116 4259
rect 112 4227 114 4258
rect 744 4227 746 4259
rect 880 4227 882 4259
rect 1016 4227 1018 4259
rect 1152 4227 1154 4259
rect 1288 4227 1290 4259
rect 111 4226 115 4227
rect 111 4221 115 4222
rect 727 4226 731 4227
rect 727 4221 731 4222
rect 743 4226 747 4227
rect 743 4221 747 4222
rect 863 4226 867 4227
rect 863 4221 867 4222
rect 879 4226 883 4227
rect 879 4221 883 4222
rect 999 4226 1003 4227
rect 999 4221 1003 4222
rect 1015 4226 1019 4227
rect 1015 4221 1019 4222
rect 1135 4226 1139 4227
rect 1135 4221 1139 4222
rect 1151 4226 1155 4227
rect 1151 4221 1155 4222
rect 1271 4226 1275 4227
rect 1271 4221 1275 4222
rect 1287 4226 1291 4227
rect 1287 4221 1291 4222
rect 112 4198 114 4221
rect 110 4197 116 4198
rect 728 4197 730 4221
rect 864 4197 866 4221
rect 1000 4197 1002 4221
rect 1136 4197 1138 4221
rect 1272 4197 1274 4221
rect 110 4193 111 4197
rect 115 4193 116 4197
rect 110 4192 116 4193
rect 726 4196 732 4197
rect 726 4192 727 4196
rect 731 4192 732 4196
rect 726 4191 732 4192
rect 862 4196 868 4197
rect 862 4192 863 4196
rect 867 4192 868 4196
rect 862 4191 868 4192
rect 998 4196 1004 4197
rect 998 4192 999 4196
rect 1003 4192 1004 4196
rect 998 4191 1004 4192
rect 1134 4196 1140 4197
rect 1134 4192 1135 4196
rect 1139 4192 1140 4196
rect 1134 4191 1140 4192
rect 1270 4196 1276 4197
rect 1270 4192 1271 4196
rect 1275 4192 1276 4196
rect 1270 4191 1276 4192
rect 698 4181 704 4182
rect 110 4180 116 4181
rect 110 4176 111 4180
rect 115 4176 116 4180
rect 698 4177 699 4181
rect 703 4177 704 4181
rect 698 4176 704 4177
rect 834 4181 840 4182
rect 834 4177 835 4181
rect 839 4177 840 4181
rect 834 4176 840 4177
rect 970 4181 976 4182
rect 970 4177 971 4181
rect 975 4177 976 4181
rect 970 4176 976 4177
rect 1106 4181 1112 4182
rect 1106 4177 1107 4181
rect 1111 4177 1112 4181
rect 1106 4176 1112 4177
rect 1242 4181 1248 4182
rect 1242 4177 1243 4181
rect 1247 4177 1248 4181
rect 1242 4176 1248 4177
rect 110 4175 116 4176
rect 112 4115 114 4175
rect 700 4115 702 4176
rect 786 4163 792 4164
rect 786 4159 787 4163
rect 791 4159 792 4163
rect 786 4158 792 4159
rect 788 4140 790 4158
rect 786 4139 792 4140
rect 786 4135 787 4139
rect 791 4135 792 4139
rect 786 4134 792 4135
rect 836 4115 838 4176
rect 850 4171 856 4172
rect 850 4167 851 4171
rect 855 4167 856 4171
rect 850 4166 856 4167
rect 962 4171 968 4172
rect 962 4167 963 4171
rect 967 4167 968 4171
rect 962 4166 968 4167
rect 852 4140 854 4166
rect 850 4139 856 4140
rect 850 4135 851 4139
rect 855 4135 856 4139
rect 850 4134 856 4135
rect 111 4114 115 4115
rect 111 4109 115 4110
rect 563 4114 567 4115
rect 563 4109 567 4110
rect 699 4114 703 4115
rect 699 4109 703 4110
rect 835 4114 839 4115
rect 835 4109 839 4110
rect 112 4049 114 4109
rect 110 4048 116 4049
rect 564 4048 566 4109
rect 650 4087 656 4088
rect 650 4083 651 4087
rect 655 4083 656 4087
rect 650 4082 656 4083
rect 652 4064 654 4082
rect 650 4063 656 4064
rect 650 4059 651 4063
rect 655 4059 656 4063
rect 650 4058 656 4059
rect 700 4048 702 4109
rect 836 4048 838 4109
rect 964 4092 966 4166
rect 972 4115 974 4176
rect 1108 4115 1110 4176
rect 1244 4115 1246 4176
rect 1332 4140 1334 4282
rect 1396 4280 1398 4341
rect 1522 4323 1528 4324
rect 1522 4319 1523 4323
rect 1527 4319 1528 4323
rect 1522 4318 1528 4319
rect 1524 4288 1526 4318
rect 1522 4287 1528 4288
rect 1522 4283 1523 4287
rect 1527 4283 1528 4287
rect 1522 4282 1528 4283
rect 1532 4280 1534 4341
rect 1658 4323 1664 4324
rect 1658 4319 1659 4323
rect 1663 4319 1664 4323
rect 1658 4318 1664 4319
rect 1618 4307 1624 4308
rect 1618 4303 1619 4307
rect 1623 4303 1624 4307
rect 1618 4302 1624 4303
rect 1394 4279 1400 4280
rect 1394 4275 1395 4279
rect 1399 4275 1400 4279
rect 1394 4274 1400 4275
rect 1530 4279 1536 4280
rect 1530 4275 1531 4279
rect 1535 4275 1536 4279
rect 1530 4274 1536 4275
rect 1422 4264 1428 4265
rect 1422 4260 1423 4264
rect 1427 4260 1428 4264
rect 1422 4259 1428 4260
rect 1558 4264 1564 4265
rect 1558 4260 1559 4264
rect 1563 4260 1564 4264
rect 1558 4259 1564 4260
rect 1424 4227 1426 4259
rect 1560 4227 1562 4259
rect 1407 4226 1411 4227
rect 1407 4221 1411 4222
rect 1423 4226 1427 4227
rect 1423 4221 1427 4222
rect 1543 4226 1547 4227
rect 1543 4221 1547 4222
rect 1559 4226 1563 4227
rect 1559 4221 1563 4222
rect 1408 4197 1410 4221
rect 1544 4197 1546 4221
rect 1406 4196 1412 4197
rect 1406 4192 1407 4196
rect 1411 4192 1412 4196
rect 1406 4191 1412 4192
rect 1542 4196 1548 4197
rect 1542 4192 1543 4196
rect 1547 4192 1548 4196
rect 1542 4191 1548 4192
rect 1378 4181 1384 4182
rect 1378 4177 1379 4181
rect 1383 4177 1384 4181
rect 1378 4176 1384 4177
rect 1514 4181 1520 4182
rect 1514 4177 1515 4181
rect 1519 4177 1520 4181
rect 1514 4176 1520 4177
rect 1330 4139 1336 4140
rect 1330 4135 1331 4139
rect 1335 4135 1336 4139
rect 1330 4134 1336 4135
rect 1380 4115 1382 4176
rect 1466 4139 1472 4140
rect 1466 4135 1467 4139
rect 1471 4135 1472 4139
rect 1466 4134 1472 4135
rect 971 4114 975 4115
rect 971 4109 975 4110
rect 1107 4114 1111 4115
rect 1107 4109 1111 4110
rect 1243 4114 1247 4115
rect 1243 4109 1247 4110
rect 1379 4114 1383 4115
rect 1379 4109 1383 4110
rect 962 4091 968 4092
rect 962 4087 963 4091
rect 967 4087 968 4091
rect 962 4086 968 4087
rect 958 4055 964 4056
rect 958 4051 959 4055
rect 963 4051 964 4055
rect 958 4050 964 4051
rect 110 4044 111 4048
rect 115 4044 116 4048
rect 110 4043 116 4044
rect 562 4047 568 4048
rect 562 4043 563 4047
rect 567 4043 568 4047
rect 562 4042 568 4043
rect 698 4047 704 4048
rect 698 4043 699 4047
rect 703 4043 704 4047
rect 698 4042 704 4043
rect 834 4047 840 4048
rect 834 4043 835 4047
rect 839 4043 840 4047
rect 834 4042 840 4043
rect 590 4032 596 4033
rect 110 4031 116 4032
rect 110 4027 111 4031
rect 115 4027 116 4031
rect 590 4028 591 4032
rect 595 4028 596 4032
rect 590 4027 596 4028
rect 726 4032 732 4033
rect 726 4028 727 4032
rect 731 4028 732 4032
rect 726 4027 732 4028
rect 862 4032 868 4033
rect 862 4028 863 4032
rect 867 4028 868 4032
rect 862 4027 868 4028
rect 110 4026 116 4027
rect 112 4003 114 4026
rect 592 4003 594 4027
rect 728 4003 730 4027
rect 864 4003 866 4027
rect 111 4002 115 4003
rect 111 3997 115 3998
rect 159 4002 163 4003
rect 159 3997 163 3998
rect 327 4002 331 4003
rect 327 3997 331 3998
rect 535 4002 539 4003
rect 535 3997 539 3998
rect 591 4002 595 4003
rect 591 3997 595 3998
rect 727 4002 731 4003
rect 727 3997 731 3998
rect 751 4002 755 4003
rect 751 3997 755 3998
rect 863 4002 867 4003
rect 863 3997 867 3998
rect 112 3974 114 3997
rect 110 3973 116 3974
rect 160 3973 162 3997
rect 328 3973 330 3997
rect 536 3973 538 3997
rect 752 3973 754 3997
rect 110 3969 111 3973
rect 115 3969 116 3973
rect 110 3968 116 3969
rect 158 3972 164 3973
rect 158 3968 159 3972
rect 163 3968 164 3972
rect 158 3967 164 3968
rect 326 3972 332 3973
rect 326 3968 327 3972
rect 331 3968 332 3972
rect 326 3967 332 3968
rect 534 3972 540 3973
rect 534 3968 535 3972
rect 539 3968 540 3972
rect 534 3967 540 3968
rect 750 3972 756 3973
rect 750 3968 751 3972
rect 755 3968 756 3972
rect 750 3967 756 3968
rect 130 3957 136 3958
rect 110 3956 116 3957
rect 110 3952 111 3956
rect 115 3952 116 3956
rect 130 3953 131 3957
rect 135 3953 136 3957
rect 130 3952 136 3953
rect 298 3957 304 3958
rect 298 3953 299 3957
rect 303 3953 304 3957
rect 298 3952 304 3953
rect 506 3957 512 3958
rect 506 3953 507 3957
rect 511 3953 512 3957
rect 506 3952 512 3953
rect 722 3957 728 3958
rect 722 3953 723 3957
rect 727 3953 728 3957
rect 722 3952 728 3953
rect 938 3957 944 3958
rect 938 3953 939 3957
rect 943 3953 944 3957
rect 938 3952 944 3953
rect 110 3951 116 3952
rect 112 3891 114 3951
rect 132 3891 134 3952
rect 234 3947 240 3948
rect 234 3943 235 3947
rect 239 3943 240 3947
rect 234 3942 240 3943
rect 286 3947 292 3948
rect 286 3943 287 3947
rect 291 3943 292 3947
rect 286 3942 292 3943
rect 111 3890 115 3891
rect 111 3885 115 3886
rect 131 3890 135 3891
rect 131 3885 135 3886
rect 112 3825 114 3885
rect 110 3824 116 3825
rect 132 3824 134 3885
rect 236 3868 238 3942
rect 288 3916 290 3942
rect 286 3915 292 3916
rect 286 3911 287 3915
rect 291 3911 292 3915
rect 286 3910 292 3911
rect 300 3891 302 3952
rect 450 3947 456 3948
rect 450 3943 451 3947
rect 455 3943 456 3947
rect 450 3942 456 3943
rect 452 3916 454 3942
rect 450 3915 456 3916
rect 450 3911 451 3915
rect 455 3911 456 3915
rect 450 3910 456 3911
rect 508 3891 510 3952
rect 702 3947 708 3948
rect 702 3943 703 3947
rect 707 3943 708 3947
rect 702 3942 708 3943
rect 704 3916 706 3942
rect 702 3915 708 3916
rect 702 3911 703 3915
rect 707 3911 708 3915
rect 702 3910 708 3911
rect 724 3891 726 3952
rect 878 3947 884 3948
rect 878 3943 879 3947
rect 883 3943 884 3947
rect 878 3942 884 3943
rect 880 3916 882 3942
rect 878 3915 884 3916
rect 878 3911 879 3915
rect 883 3911 884 3915
rect 878 3910 884 3911
rect 940 3891 942 3952
rect 960 3916 962 4050
rect 972 4048 974 4109
rect 1108 4048 1110 4109
rect 1244 4048 1246 4109
rect 1380 4048 1382 4109
rect 1468 4056 1470 4134
rect 1516 4115 1518 4176
rect 1620 4172 1622 4302
rect 1660 4288 1662 4318
rect 1658 4287 1664 4288
rect 1658 4283 1659 4287
rect 1663 4283 1664 4287
rect 1658 4282 1664 4283
rect 1668 4280 1670 4341
rect 1780 4288 1782 4370
rect 1936 4347 1938 4411
rect 1976 4379 1978 4414
rect 2296 4379 2298 4415
rect 1975 4378 1979 4379
rect 1975 4373 1979 4374
rect 2023 4378 2027 4379
rect 2023 4373 2027 4374
rect 2199 4378 2203 4379
rect 2199 4373 2203 4374
rect 2295 4378 2299 4379
rect 2295 4373 2299 4374
rect 1976 4350 1978 4373
rect 1974 4349 1980 4350
rect 2024 4349 2026 4373
rect 2200 4349 2202 4373
rect 1935 4346 1939 4347
rect 1974 4345 1975 4349
rect 1979 4345 1980 4349
rect 1974 4344 1980 4345
rect 2022 4348 2028 4349
rect 2022 4344 2023 4348
rect 2027 4344 2028 4348
rect 2022 4343 2028 4344
rect 2198 4348 2204 4349
rect 2198 4344 2199 4348
rect 2203 4344 2204 4348
rect 2198 4343 2204 4344
rect 1935 4341 1939 4342
rect 1778 4287 1784 4288
rect 1778 4283 1779 4287
rect 1783 4283 1784 4287
rect 1778 4282 1784 4283
rect 1936 4281 1938 4341
rect 1994 4333 2000 4334
rect 1974 4332 1980 4333
rect 1974 4328 1975 4332
rect 1979 4328 1980 4332
rect 1994 4329 1995 4333
rect 1999 4329 2000 4333
rect 1994 4328 2000 4329
rect 2170 4333 2176 4334
rect 2170 4329 2171 4333
rect 2175 4329 2176 4333
rect 2170 4328 2176 4329
rect 2370 4333 2376 4334
rect 2370 4329 2371 4333
rect 2375 4329 2376 4333
rect 2370 4328 2376 4329
rect 1974 4327 1980 4328
rect 1934 4280 1940 4281
rect 1666 4279 1672 4280
rect 1666 4275 1667 4279
rect 1671 4275 1672 4279
rect 1934 4276 1935 4280
rect 1939 4276 1940 4280
rect 1934 4275 1940 4276
rect 1666 4274 1672 4275
rect 1694 4264 1700 4265
rect 1694 4260 1695 4264
rect 1699 4260 1700 4264
rect 1694 4259 1700 4260
rect 1934 4263 1940 4264
rect 1976 4263 1978 4327
rect 1996 4263 1998 4328
rect 2098 4323 2104 4324
rect 2098 4319 2099 4323
rect 2103 4319 2104 4323
rect 2098 4318 2104 4319
rect 1934 4259 1935 4263
rect 1939 4259 1940 4263
rect 1696 4227 1698 4259
rect 1934 4258 1940 4259
rect 1975 4262 1979 4263
rect 1936 4227 1938 4258
rect 1975 4257 1979 4258
rect 1995 4262 1999 4263
rect 1995 4257 1999 4258
rect 1679 4226 1683 4227
rect 1679 4221 1683 4222
rect 1695 4226 1699 4227
rect 1695 4221 1699 4222
rect 1815 4226 1819 4227
rect 1815 4221 1819 4222
rect 1935 4226 1939 4227
rect 1935 4221 1939 4222
rect 1680 4197 1682 4221
rect 1816 4197 1818 4221
rect 1936 4198 1938 4221
rect 1946 4203 1952 4204
rect 1946 4199 1947 4203
rect 1951 4199 1952 4203
rect 1946 4198 1952 4199
rect 1934 4197 1940 4198
rect 1678 4196 1684 4197
rect 1678 4192 1679 4196
rect 1683 4192 1684 4196
rect 1678 4191 1684 4192
rect 1814 4196 1820 4197
rect 1814 4192 1815 4196
rect 1819 4192 1820 4196
rect 1934 4193 1935 4197
rect 1939 4193 1940 4197
rect 1934 4192 1940 4193
rect 1814 4191 1820 4192
rect 1650 4181 1656 4182
rect 1650 4177 1651 4181
rect 1655 4177 1656 4181
rect 1650 4176 1656 4177
rect 1786 4181 1792 4182
rect 1786 4177 1787 4181
rect 1791 4177 1792 4181
rect 1786 4176 1792 4177
rect 1934 4180 1940 4181
rect 1934 4176 1935 4180
rect 1939 4176 1940 4180
rect 1530 4171 1536 4172
rect 1530 4167 1531 4171
rect 1535 4167 1536 4171
rect 1530 4166 1536 4167
rect 1618 4171 1624 4172
rect 1618 4167 1619 4171
rect 1623 4167 1624 4171
rect 1618 4166 1624 4167
rect 1532 4140 1534 4166
rect 1530 4139 1536 4140
rect 1530 4135 1531 4139
rect 1535 4135 1536 4139
rect 1530 4134 1536 4135
rect 1652 4115 1654 4176
rect 1778 4171 1784 4172
rect 1778 4167 1779 4171
rect 1783 4167 1784 4171
rect 1778 4166 1784 4167
rect 1515 4114 1519 4115
rect 1515 4109 1519 4110
rect 1651 4114 1655 4115
rect 1651 4109 1655 4110
rect 1474 4075 1480 4076
rect 1474 4071 1475 4075
rect 1479 4071 1480 4075
rect 1474 4070 1480 4071
rect 1466 4055 1472 4056
rect 1466 4051 1467 4055
rect 1471 4051 1472 4055
rect 1466 4050 1472 4051
rect 970 4047 976 4048
rect 970 4043 971 4047
rect 975 4043 976 4047
rect 970 4042 976 4043
rect 1106 4047 1112 4048
rect 1106 4043 1107 4047
rect 1111 4043 1112 4047
rect 1106 4042 1112 4043
rect 1242 4047 1248 4048
rect 1242 4043 1243 4047
rect 1247 4043 1248 4047
rect 1242 4042 1248 4043
rect 1378 4047 1384 4048
rect 1378 4043 1379 4047
rect 1383 4043 1384 4047
rect 1378 4042 1384 4043
rect 998 4032 1004 4033
rect 998 4028 999 4032
rect 1003 4028 1004 4032
rect 998 4027 1004 4028
rect 1134 4032 1140 4033
rect 1134 4028 1135 4032
rect 1139 4028 1140 4032
rect 1134 4027 1140 4028
rect 1270 4032 1276 4033
rect 1270 4028 1271 4032
rect 1275 4028 1276 4032
rect 1270 4027 1276 4028
rect 1406 4032 1412 4033
rect 1406 4028 1407 4032
rect 1411 4028 1412 4032
rect 1406 4027 1412 4028
rect 1000 4003 1002 4027
rect 1136 4003 1138 4027
rect 1272 4003 1274 4027
rect 1408 4003 1410 4027
rect 967 4002 971 4003
rect 967 3997 971 3998
rect 999 4002 1003 4003
rect 999 3997 1003 3998
rect 1135 4002 1139 4003
rect 1135 3997 1139 3998
rect 1183 4002 1187 4003
rect 1183 3997 1187 3998
rect 1271 4002 1275 4003
rect 1271 3997 1275 3998
rect 1399 4002 1403 4003
rect 1399 3997 1403 3998
rect 1407 4002 1411 4003
rect 1407 3997 1411 3998
rect 968 3973 970 3997
rect 1184 3973 1186 3997
rect 1400 3973 1402 3997
rect 966 3972 972 3973
rect 966 3968 967 3972
rect 971 3968 972 3972
rect 966 3967 972 3968
rect 1182 3972 1188 3973
rect 1182 3968 1183 3972
rect 1187 3968 1188 3972
rect 1182 3967 1188 3968
rect 1398 3972 1404 3973
rect 1398 3968 1399 3972
rect 1403 3968 1404 3972
rect 1398 3967 1404 3968
rect 1154 3957 1160 3958
rect 1154 3953 1155 3957
rect 1159 3953 1160 3957
rect 1154 3952 1160 3953
rect 1370 3957 1376 3958
rect 1370 3953 1371 3957
rect 1375 3953 1376 3957
rect 1370 3952 1376 3953
rect 958 3915 964 3916
rect 958 3911 959 3915
rect 963 3911 964 3915
rect 958 3910 964 3911
rect 1156 3891 1158 3952
rect 1242 3915 1248 3916
rect 1242 3911 1243 3915
rect 1247 3911 1248 3915
rect 1242 3910 1248 3911
rect 299 3890 303 3891
rect 299 3885 303 3886
rect 355 3890 359 3891
rect 355 3885 359 3886
rect 507 3890 511 3891
rect 507 3885 511 3886
rect 619 3890 623 3891
rect 619 3885 623 3886
rect 723 3890 727 3891
rect 723 3885 727 3886
rect 899 3890 903 3891
rect 899 3885 903 3886
rect 939 3890 943 3891
rect 939 3885 943 3886
rect 1155 3890 1159 3891
rect 1155 3885 1159 3886
rect 1195 3890 1199 3891
rect 1195 3885 1199 3886
rect 234 3867 240 3868
rect 234 3863 235 3867
rect 239 3863 240 3867
rect 234 3862 240 3863
rect 258 3867 264 3868
rect 258 3863 259 3867
rect 263 3863 264 3867
rect 258 3862 264 3863
rect 260 3832 262 3862
rect 258 3831 264 3832
rect 258 3827 259 3831
rect 263 3827 264 3831
rect 258 3826 264 3827
rect 356 3824 358 3885
rect 482 3867 488 3868
rect 482 3863 483 3867
rect 487 3863 488 3867
rect 482 3862 488 3863
rect 484 3832 486 3862
rect 482 3831 488 3832
rect 482 3827 483 3831
rect 487 3827 488 3831
rect 482 3826 488 3827
rect 620 3824 622 3885
rect 746 3867 752 3868
rect 746 3863 747 3867
rect 751 3863 752 3867
rect 746 3862 752 3863
rect 748 3832 750 3862
rect 746 3831 752 3832
rect 746 3827 747 3831
rect 751 3827 752 3831
rect 746 3826 752 3827
rect 850 3831 856 3832
rect 850 3827 851 3831
rect 855 3827 856 3831
rect 850 3826 856 3827
rect 110 3820 111 3824
rect 115 3820 116 3824
rect 110 3819 116 3820
rect 130 3823 136 3824
rect 130 3819 131 3823
rect 135 3819 136 3823
rect 130 3818 136 3819
rect 354 3823 360 3824
rect 354 3819 355 3823
rect 359 3819 360 3823
rect 354 3818 360 3819
rect 618 3823 624 3824
rect 618 3819 619 3823
rect 623 3819 624 3823
rect 618 3818 624 3819
rect 158 3808 164 3809
rect 110 3807 116 3808
rect 110 3803 111 3807
rect 115 3803 116 3807
rect 158 3804 159 3808
rect 163 3804 164 3808
rect 158 3803 164 3804
rect 382 3808 388 3809
rect 382 3804 383 3808
rect 387 3804 388 3808
rect 382 3803 388 3804
rect 646 3808 652 3809
rect 646 3804 647 3808
rect 651 3804 652 3808
rect 646 3803 652 3804
rect 110 3802 116 3803
rect 112 3767 114 3802
rect 160 3767 162 3803
rect 384 3767 386 3803
rect 648 3767 650 3803
rect 111 3766 115 3767
rect 111 3761 115 3762
rect 159 3766 163 3767
rect 159 3761 163 3762
rect 247 3766 251 3767
rect 247 3761 251 3762
rect 383 3766 387 3767
rect 383 3761 387 3762
rect 519 3766 523 3767
rect 519 3761 523 3762
rect 647 3766 651 3767
rect 647 3761 651 3762
rect 791 3766 795 3767
rect 791 3761 795 3762
rect 112 3738 114 3761
rect 110 3737 116 3738
rect 248 3737 250 3761
rect 520 3737 522 3761
rect 792 3737 794 3761
rect 110 3733 111 3737
rect 115 3733 116 3737
rect 110 3732 116 3733
rect 246 3736 252 3737
rect 246 3732 247 3736
rect 251 3732 252 3736
rect 246 3731 252 3732
rect 518 3736 524 3737
rect 518 3732 519 3736
rect 523 3732 524 3736
rect 518 3731 524 3732
rect 790 3736 796 3737
rect 790 3732 791 3736
rect 795 3732 796 3736
rect 790 3731 796 3732
rect 218 3721 224 3722
rect 110 3720 116 3721
rect 110 3716 111 3720
rect 115 3716 116 3720
rect 218 3717 219 3721
rect 223 3717 224 3721
rect 218 3716 224 3717
rect 490 3721 496 3722
rect 490 3717 491 3721
rect 495 3717 496 3721
rect 490 3716 496 3717
rect 762 3721 768 3722
rect 762 3717 763 3721
rect 767 3717 768 3721
rect 762 3716 768 3717
rect 110 3715 116 3716
rect 112 3639 114 3715
rect 220 3639 222 3716
rect 306 3703 312 3704
rect 306 3699 307 3703
rect 311 3699 312 3703
rect 306 3698 312 3699
rect 308 3680 310 3698
rect 306 3679 312 3680
rect 306 3675 307 3679
rect 311 3675 312 3679
rect 306 3674 312 3675
rect 492 3639 494 3716
rect 506 3711 512 3712
rect 506 3707 507 3711
rect 511 3707 512 3711
rect 506 3706 512 3707
rect 594 3711 600 3712
rect 594 3707 595 3711
rect 599 3707 600 3711
rect 594 3706 600 3707
rect 508 3680 510 3706
rect 506 3679 512 3680
rect 506 3675 507 3679
rect 511 3675 512 3679
rect 506 3674 512 3675
rect 111 3638 115 3639
rect 111 3633 115 3634
rect 219 3638 223 3639
rect 219 3633 223 3634
rect 491 3638 495 3639
rect 491 3633 495 3634
rect 112 3573 114 3633
rect 110 3572 116 3573
rect 492 3572 494 3633
rect 596 3616 598 3706
rect 764 3639 766 3716
rect 852 3680 854 3826
rect 900 3824 902 3885
rect 1196 3824 1198 3885
rect 1244 3832 1246 3910
rect 1372 3891 1374 3952
rect 1476 3948 1478 4070
rect 1516 4048 1518 4109
rect 1638 4055 1644 4056
rect 1638 4051 1639 4055
rect 1643 4051 1644 4055
rect 1638 4050 1644 4051
rect 1514 4047 1520 4048
rect 1514 4043 1515 4047
rect 1519 4043 1520 4047
rect 1514 4042 1520 4043
rect 1542 4032 1548 4033
rect 1542 4028 1543 4032
rect 1547 4028 1548 4032
rect 1542 4027 1548 4028
rect 1544 4003 1546 4027
rect 1543 4002 1547 4003
rect 1543 3997 1547 3998
rect 1615 4002 1619 4003
rect 1615 3997 1619 3998
rect 1616 3973 1618 3997
rect 1614 3972 1620 3973
rect 1614 3968 1615 3972
rect 1619 3968 1620 3972
rect 1614 3967 1620 3968
rect 1586 3957 1592 3958
rect 1586 3953 1587 3957
rect 1591 3953 1592 3957
rect 1586 3952 1592 3953
rect 1386 3947 1392 3948
rect 1386 3943 1387 3947
rect 1391 3943 1392 3947
rect 1386 3942 1392 3943
rect 1474 3947 1480 3948
rect 1474 3943 1475 3947
rect 1479 3943 1480 3947
rect 1474 3942 1480 3943
rect 1388 3916 1390 3942
rect 1386 3915 1392 3916
rect 1386 3911 1387 3915
rect 1391 3911 1392 3915
rect 1386 3910 1392 3911
rect 1588 3891 1590 3952
rect 1640 3916 1642 4050
rect 1652 4048 1654 4109
rect 1780 4092 1782 4166
rect 1788 4115 1790 4176
rect 1934 4175 1940 4176
rect 1794 4171 1800 4172
rect 1794 4167 1795 4171
rect 1799 4167 1800 4171
rect 1794 4166 1800 4167
rect 1796 4140 1798 4166
rect 1794 4139 1800 4140
rect 1794 4135 1795 4139
rect 1799 4135 1800 4139
rect 1794 4134 1800 4135
rect 1936 4115 1938 4175
rect 1948 4140 1950 4198
rect 1976 4197 1978 4257
rect 1974 4196 1980 4197
rect 1996 4196 1998 4257
rect 2100 4240 2102 4318
rect 2172 4263 2174 4328
rect 2310 4323 2316 4324
rect 2310 4319 2311 4323
rect 2315 4319 2316 4323
rect 2310 4318 2316 4319
rect 2312 4292 2314 4318
rect 2310 4291 2316 4292
rect 2310 4287 2311 4291
rect 2315 4287 2316 4291
rect 2310 4286 2316 4287
rect 2372 4263 2374 4328
rect 2392 4292 2394 4438
rect 2516 4436 2518 4497
rect 2620 4480 2622 4566
rect 2748 4503 2750 4576
rect 2836 4540 2838 4678
rect 3800 4677 3802 4737
rect 3840 4691 3842 4751
rect 3860 4691 3862 4752
rect 4002 4747 4008 4748
rect 4002 4743 4003 4747
rect 4007 4743 4008 4747
rect 4002 4742 4008 4743
rect 4004 4716 4006 4742
rect 4002 4715 4008 4716
rect 4002 4711 4003 4715
rect 4007 4711 4008 4715
rect 4002 4710 4008 4711
rect 4044 4691 4046 4752
rect 4130 4739 4136 4740
rect 4130 4735 4131 4739
rect 4135 4735 4136 4739
rect 4130 4734 4136 4735
rect 4132 4716 4134 4734
rect 4130 4715 4136 4716
rect 4130 4711 4131 4715
rect 4135 4711 4136 4715
rect 4130 4710 4136 4711
rect 4138 4715 4144 4716
rect 4138 4711 4139 4715
rect 4143 4711 4144 4715
rect 4138 4710 4144 4711
rect 3839 4690 3843 4691
rect 3839 4685 3843 4686
rect 3859 4690 3863 4691
rect 3859 4685 3863 4686
rect 3995 4690 3999 4691
rect 3995 4685 3999 4686
rect 4043 4690 4047 4691
rect 4043 4685 4047 4686
rect 4131 4690 4135 4691
rect 4131 4685 4135 4686
rect 3798 4676 3804 4677
rect 3798 4672 3799 4676
rect 3803 4672 3804 4676
rect 3798 4671 3804 4672
rect 3778 4667 3784 4668
rect 3778 4663 3779 4667
rect 3783 4663 3784 4667
rect 3778 4662 3784 4663
rect 3015 4626 3019 4627
rect 3015 4621 3019 4622
rect 3247 4626 3251 4627
rect 3247 4621 3251 4622
rect 3471 4626 3475 4627
rect 3471 4621 3475 4622
rect 3679 4626 3683 4627
rect 3679 4621 3683 4622
rect 3016 4597 3018 4621
rect 3248 4597 3250 4621
rect 3472 4597 3474 4621
rect 3680 4597 3682 4621
rect 3014 4596 3020 4597
rect 3014 4592 3015 4596
rect 3019 4592 3020 4596
rect 3014 4591 3020 4592
rect 3246 4596 3252 4597
rect 3246 4592 3247 4596
rect 3251 4592 3252 4596
rect 3246 4591 3252 4592
rect 3470 4596 3476 4597
rect 3470 4592 3471 4596
rect 3475 4592 3476 4596
rect 3470 4591 3476 4592
rect 3678 4596 3684 4597
rect 3678 4592 3679 4596
rect 3683 4592 3684 4596
rect 3678 4591 3684 4592
rect 2986 4581 2992 4582
rect 2986 4577 2987 4581
rect 2991 4577 2992 4581
rect 2986 4576 2992 4577
rect 3218 4581 3224 4582
rect 3218 4577 3219 4581
rect 3223 4577 3224 4581
rect 3218 4576 3224 4577
rect 3442 4581 3448 4582
rect 3442 4577 3443 4581
rect 3447 4577 3448 4581
rect 3442 4576 3448 4577
rect 3650 4581 3656 4582
rect 3650 4577 3651 4581
rect 3655 4577 3656 4581
rect 3650 4576 3656 4577
rect 2834 4539 2840 4540
rect 2834 4535 2835 4539
rect 2839 4535 2840 4539
rect 2834 4534 2840 4535
rect 2988 4503 2990 4576
rect 3074 4539 3080 4540
rect 3074 4535 3075 4539
rect 3079 4535 3080 4539
rect 3074 4534 3080 4535
rect 2747 4502 2751 4503
rect 2747 4497 2751 4498
rect 2971 4502 2975 4503
rect 2971 4497 2975 4498
rect 2987 4502 2991 4503
rect 2987 4497 2991 4498
rect 2618 4479 2624 4480
rect 2618 4475 2619 4479
rect 2623 4475 2624 4479
rect 2618 4474 2624 4475
rect 2748 4436 2750 4497
rect 2874 4479 2880 4480
rect 2834 4475 2840 4476
rect 2834 4471 2835 4475
rect 2839 4471 2840 4475
rect 2874 4475 2875 4479
rect 2879 4475 2880 4479
rect 2874 4474 2880 4475
rect 2834 4470 2840 4471
rect 2514 4435 2520 4436
rect 2514 4431 2515 4435
rect 2519 4431 2520 4435
rect 2514 4430 2520 4431
rect 2746 4435 2752 4436
rect 2746 4431 2747 4435
rect 2751 4431 2752 4435
rect 2746 4430 2752 4431
rect 2542 4420 2548 4421
rect 2542 4416 2543 4420
rect 2547 4416 2548 4420
rect 2542 4415 2548 4416
rect 2774 4420 2780 4421
rect 2774 4416 2775 4420
rect 2779 4416 2780 4420
rect 2774 4415 2780 4416
rect 2544 4379 2546 4415
rect 2776 4379 2778 4415
rect 2399 4378 2403 4379
rect 2399 4373 2403 4374
rect 2543 4378 2547 4379
rect 2543 4373 2547 4374
rect 2591 4378 2595 4379
rect 2591 4373 2595 4374
rect 2775 4378 2779 4379
rect 2775 4373 2779 4374
rect 2400 4349 2402 4373
rect 2592 4349 2594 4373
rect 2776 4349 2778 4373
rect 2398 4348 2404 4349
rect 2398 4344 2399 4348
rect 2403 4344 2404 4348
rect 2398 4343 2404 4344
rect 2590 4348 2596 4349
rect 2590 4344 2591 4348
rect 2595 4344 2596 4348
rect 2590 4343 2596 4344
rect 2774 4348 2780 4349
rect 2774 4344 2775 4348
rect 2779 4344 2780 4348
rect 2774 4343 2780 4344
rect 2562 4333 2568 4334
rect 2562 4329 2563 4333
rect 2567 4329 2568 4333
rect 2562 4328 2568 4329
rect 2746 4333 2752 4334
rect 2746 4329 2747 4333
rect 2751 4329 2752 4333
rect 2746 4328 2752 4329
rect 2390 4291 2396 4292
rect 2390 4287 2391 4291
rect 2395 4287 2396 4291
rect 2390 4286 2396 4287
rect 2564 4263 2566 4328
rect 2630 4291 2636 4292
rect 2630 4287 2631 4291
rect 2635 4287 2636 4291
rect 2630 4286 2636 4287
rect 2171 4262 2175 4263
rect 2171 4257 2175 4258
rect 2243 4262 2247 4263
rect 2243 4257 2247 4258
rect 2371 4262 2375 4263
rect 2371 4257 2375 4258
rect 2507 4262 2511 4263
rect 2507 4257 2511 4258
rect 2563 4262 2567 4263
rect 2563 4257 2567 4258
rect 2098 4239 2104 4240
rect 2098 4235 2099 4239
rect 2103 4235 2104 4239
rect 2098 4234 2104 4235
rect 2244 4196 2246 4257
rect 2330 4235 2336 4236
rect 2330 4231 2331 4235
rect 2335 4231 2336 4235
rect 2330 4230 2336 4231
rect 2332 4212 2334 4230
rect 2330 4211 2336 4212
rect 2330 4207 2331 4211
rect 2335 4207 2336 4211
rect 2330 4206 2336 4207
rect 2508 4196 2510 4257
rect 2632 4204 2634 4286
rect 2748 4263 2750 4328
rect 2762 4323 2768 4324
rect 2762 4319 2763 4323
rect 2767 4319 2768 4323
rect 2762 4318 2768 4319
rect 2764 4292 2766 4318
rect 2836 4316 2838 4470
rect 2876 4444 2878 4474
rect 2874 4443 2880 4444
rect 2874 4439 2875 4443
rect 2879 4439 2880 4443
rect 2874 4438 2880 4439
rect 2972 4436 2974 4497
rect 3076 4493 3078 4534
rect 3220 4503 3222 4576
rect 3234 4571 3240 4572
rect 3234 4567 3235 4571
rect 3239 4567 3240 4571
rect 3234 4566 3240 4567
rect 3236 4540 3238 4566
rect 3234 4539 3240 4540
rect 3234 4535 3235 4539
rect 3239 4535 3240 4539
rect 3234 4534 3240 4535
rect 3444 4503 3446 4576
rect 3458 4571 3464 4572
rect 3458 4567 3459 4571
rect 3463 4567 3464 4571
rect 3458 4566 3464 4567
rect 3460 4540 3462 4566
rect 3458 4539 3464 4540
rect 3458 4535 3459 4539
rect 3463 4535 3464 4539
rect 3458 4534 3464 4535
rect 3652 4503 3654 4576
rect 3780 4572 3782 4662
rect 3798 4659 3804 4660
rect 3798 4655 3799 4659
rect 3803 4655 3804 4659
rect 3798 4654 3804 4655
rect 3800 4627 3802 4654
rect 3799 4626 3803 4627
rect 3840 4625 3842 4685
rect 3799 4621 3803 4622
rect 3838 4624 3844 4625
rect 3860 4624 3862 4685
rect 3986 4667 3992 4668
rect 3986 4663 3987 4667
rect 3991 4663 3992 4667
rect 3986 4662 3992 4663
rect 3988 4632 3990 4662
rect 3986 4631 3992 4632
rect 3986 4627 3987 4631
rect 3991 4627 3992 4631
rect 3986 4626 3992 4627
rect 3996 4624 3998 4685
rect 4132 4624 4134 4685
rect 4140 4632 4142 4710
rect 4268 4691 4270 4752
rect 4508 4691 4510 4752
rect 4522 4747 4528 4748
rect 4522 4743 4523 4747
rect 4527 4743 4528 4747
rect 4522 4742 4528 4743
rect 4524 4716 4526 4742
rect 4522 4715 4528 4716
rect 4522 4711 4523 4715
rect 4527 4711 4528 4715
rect 4522 4710 4528 4711
rect 4756 4691 4758 4752
rect 4770 4747 4776 4748
rect 4770 4743 4771 4747
rect 4775 4743 4776 4747
rect 4770 4742 4776 4743
rect 4772 4716 4774 4742
rect 4770 4715 4776 4716
rect 4770 4711 4771 4715
rect 4775 4711 4776 4715
rect 4770 4710 4776 4711
rect 5012 4691 5014 4752
rect 5098 4739 5104 4740
rect 5098 4735 5099 4739
rect 5103 4735 5104 4739
rect 5098 4734 5104 4735
rect 5100 4716 5102 4734
rect 5098 4715 5104 4716
rect 5098 4711 5099 4715
rect 5103 4711 5104 4715
rect 5098 4710 5104 4711
rect 5276 4691 5278 4752
rect 5290 4747 5296 4748
rect 5290 4743 5291 4747
rect 5295 4743 5296 4747
rect 5290 4742 5296 4743
rect 5370 4747 5376 4748
rect 5370 4743 5371 4747
rect 5375 4743 5376 4747
rect 5370 4742 5376 4743
rect 5292 4716 5294 4742
rect 5290 4715 5296 4716
rect 5290 4711 5291 4715
rect 5295 4711 5296 4715
rect 5290 4710 5296 4711
rect 4267 4690 4271 4691
rect 4267 4685 4271 4686
rect 4403 4690 4407 4691
rect 4403 4685 4407 4686
rect 4507 4690 4511 4691
rect 4507 4685 4511 4686
rect 4539 4690 4543 4691
rect 4539 4685 4543 4686
rect 4675 4690 4679 4691
rect 4675 4685 4679 4686
rect 4755 4690 4759 4691
rect 4755 4685 4759 4686
rect 4819 4690 4823 4691
rect 4819 4685 4823 4686
rect 4963 4690 4967 4691
rect 4963 4685 4967 4686
rect 5011 4690 5015 4691
rect 5011 4685 5015 4686
rect 5107 4690 5111 4691
rect 5107 4685 5111 4686
rect 5243 4690 5247 4691
rect 5243 4685 5247 4686
rect 5275 4690 5279 4691
rect 5275 4685 5279 4686
rect 4258 4667 4264 4668
rect 4218 4663 4224 4664
rect 4218 4659 4219 4663
rect 4223 4659 4224 4663
rect 4258 4663 4259 4667
rect 4263 4663 4264 4667
rect 4258 4662 4264 4663
rect 4218 4658 4224 4659
rect 4220 4640 4222 4658
rect 4218 4639 4224 4640
rect 4218 4635 4219 4639
rect 4223 4635 4224 4639
rect 4218 4634 4224 4635
rect 4260 4632 4262 4662
rect 4138 4631 4144 4632
rect 4138 4627 4139 4631
rect 4143 4627 4144 4631
rect 4138 4626 4144 4627
rect 4258 4631 4264 4632
rect 4258 4627 4259 4631
rect 4263 4627 4264 4631
rect 4258 4626 4264 4627
rect 4268 4624 4270 4685
rect 4394 4667 4400 4668
rect 4394 4663 4395 4667
rect 4399 4663 4400 4667
rect 4394 4662 4400 4663
rect 4396 4632 4398 4662
rect 4394 4631 4400 4632
rect 4394 4627 4395 4631
rect 4399 4627 4400 4631
rect 4394 4626 4400 4627
rect 4404 4624 4406 4685
rect 4540 4624 4542 4685
rect 4594 4631 4600 4632
rect 4594 4627 4595 4631
rect 4599 4627 4600 4631
rect 4594 4626 4600 4627
rect 3800 4598 3802 4621
rect 3838 4620 3839 4624
rect 3843 4620 3844 4624
rect 3838 4619 3844 4620
rect 3858 4623 3864 4624
rect 3858 4619 3859 4623
rect 3863 4619 3864 4623
rect 3858 4618 3864 4619
rect 3994 4623 4000 4624
rect 3994 4619 3995 4623
rect 3999 4619 4000 4623
rect 3994 4618 4000 4619
rect 4130 4623 4136 4624
rect 4130 4619 4131 4623
rect 4135 4619 4136 4623
rect 4130 4618 4136 4619
rect 4266 4623 4272 4624
rect 4266 4619 4267 4623
rect 4271 4619 4272 4623
rect 4266 4618 4272 4619
rect 4402 4623 4408 4624
rect 4402 4619 4403 4623
rect 4407 4619 4408 4623
rect 4402 4618 4408 4619
rect 4538 4623 4544 4624
rect 4538 4619 4539 4623
rect 4543 4619 4544 4623
rect 4538 4618 4544 4619
rect 3886 4608 3892 4609
rect 3838 4607 3844 4608
rect 3838 4603 3839 4607
rect 3843 4603 3844 4607
rect 3886 4604 3887 4608
rect 3891 4604 3892 4608
rect 3886 4603 3892 4604
rect 4022 4608 4028 4609
rect 4022 4604 4023 4608
rect 4027 4604 4028 4608
rect 4022 4603 4028 4604
rect 4158 4608 4164 4609
rect 4158 4604 4159 4608
rect 4163 4604 4164 4608
rect 4158 4603 4164 4604
rect 4294 4608 4300 4609
rect 4294 4604 4295 4608
rect 4299 4604 4300 4608
rect 4294 4603 4300 4604
rect 4430 4608 4436 4609
rect 4430 4604 4431 4608
rect 4435 4604 4436 4608
rect 4430 4603 4436 4604
rect 4566 4608 4572 4609
rect 4566 4604 4567 4608
rect 4571 4604 4572 4608
rect 4566 4603 4572 4604
rect 3838 4602 3844 4603
rect 3798 4597 3804 4598
rect 3798 4593 3799 4597
rect 3803 4593 3804 4597
rect 3798 4592 3804 4593
rect 3798 4580 3804 4581
rect 3798 4576 3799 4580
rect 3803 4576 3804 4580
rect 3840 4579 3842 4602
rect 3888 4579 3890 4603
rect 4024 4579 4026 4603
rect 4160 4579 4162 4603
rect 4296 4579 4298 4603
rect 4432 4579 4434 4603
rect 4568 4579 4570 4603
rect 3798 4575 3804 4576
rect 3839 4578 3843 4579
rect 3666 4571 3672 4572
rect 3666 4567 3667 4571
rect 3671 4567 3672 4571
rect 3666 4566 3672 4567
rect 3778 4571 3784 4572
rect 3778 4567 3779 4571
rect 3783 4567 3784 4571
rect 3778 4566 3784 4567
rect 3668 4540 3670 4566
rect 3666 4539 3672 4540
rect 3666 4535 3667 4539
rect 3671 4535 3672 4539
rect 3666 4534 3672 4535
rect 3800 4503 3802 4575
rect 3839 4573 3843 4574
rect 3887 4578 3891 4579
rect 3887 4573 3891 4574
rect 4023 4578 4027 4579
rect 4023 4573 4027 4574
rect 4159 4578 4163 4579
rect 4159 4573 4163 4574
rect 4295 4578 4299 4579
rect 4295 4573 4299 4574
rect 4431 4578 4435 4579
rect 4431 4573 4435 4574
rect 4567 4578 4571 4579
rect 4567 4573 4571 4574
rect 3840 4550 3842 4573
rect 3838 4549 3844 4550
rect 3838 4545 3839 4549
rect 3843 4545 3844 4549
rect 3838 4544 3844 4545
rect 3838 4532 3844 4533
rect 3838 4528 3839 4532
rect 3843 4528 3844 4532
rect 3838 4527 3844 4528
rect 3187 4502 3191 4503
rect 3187 4497 3191 4498
rect 3219 4502 3223 4503
rect 3219 4497 3223 4498
rect 3395 4502 3399 4503
rect 3395 4497 3399 4498
rect 3443 4502 3447 4503
rect 3443 4497 3447 4498
rect 3611 4502 3615 4503
rect 3611 4497 3615 4498
rect 3651 4502 3655 4503
rect 3651 4497 3655 4498
rect 3799 4502 3803 4503
rect 3799 4497 3803 4498
rect 3075 4492 3079 4493
rect 3075 4487 3079 4488
rect 3098 4479 3104 4480
rect 3098 4475 3099 4479
rect 3103 4475 3104 4479
rect 3098 4474 3104 4475
rect 3100 4444 3102 4474
rect 3098 4443 3104 4444
rect 3098 4439 3099 4443
rect 3103 4439 3104 4443
rect 3098 4438 3104 4439
rect 3188 4436 3190 4497
rect 3314 4479 3320 4480
rect 3314 4475 3315 4479
rect 3319 4475 3320 4479
rect 3314 4474 3320 4475
rect 3316 4444 3318 4474
rect 3314 4443 3320 4444
rect 3314 4439 3315 4443
rect 3319 4439 3320 4443
rect 3314 4438 3320 4439
rect 3396 4436 3398 4497
rect 3522 4479 3528 4480
rect 3522 4475 3523 4479
rect 3527 4475 3528 4479
rect 3522 4474 3528 4475
rect 3524 4444 3526 4474
rect 3522 4443 3528 4444
rect 3522 4439 3523 4443
rect 3527 4439 3528 4443
rect 3522 4438 3528 4439
rect 3612 4436 3614 4497
rect 3735 4492 3739 4493
rect 3735 4487 3739 4488
rect 3736 4444 3738 4487
rect 3734 4443 3740 4444
rect 3734 4439 3735 4443
rect 3739 4439 3740 4443
rect 3734 4438 3740 4439
rect 3800 4437 3802 4497
rect 3840 4463 3842 4527
rect 4596 4492 4598 4626
rect 4676 4624 4678 4685
rect 4820 4624 4822 4685
rect 4964 4624 4966 4685
rect 5108 4624 5110 4685
rect 5244 4624 5246 4685
rect 5372 4668 5374 4742
rect 5516 4691 5518 4752
rect 5604 4716 5606 4926
rect 5664 4925 5666 4985
rect 5662 4924 5668 4925
rect 5662 4920 5663 4924
rect 5667 4920 5668 4924
rect 5662 4919 5668 4920
rect 5662 4907 5668 4908
rect 5662 4903 5663 4907
rect 5667 4903 5668 4907
rect 5662 4902 5668 4903
rect 5664 4803 5666 4902
rect 5663 4802 5667 4803
rect 5663 4797 5667 4798
rect 5664 4774 5666 4797
rect 5662 4773 5668 4774
rect 5662 4769 5663 4773
rect 5667 4769 5668 4773
rect 5662 4768 5668 4769
rect 5662 4756 5668 4757
rect 5662 4752 5663 4756
rect 5667 4752 5668 4756
rect 5662 4751 5668 4752
rect 5602 4715 5608 4716
rect 5602 4711 5603 4715
rect 5607 4711 5608 4715
rect 5602 4710 5608 4711
rect 5664 4691 5666 4751
rect 5379 4690 5383 4691
rect 5379 4685 5383 4686
rect 5515 4690 5519 4691
rect 5515 4685 5519 4686
rect 5663 4690 5667 4691
rect 5663 4685 5667 4686
rect 5370 4667 5376 4668
rect 5330 4663 5336 4664
rect 5330 4659 5331 4663
rect 5335 4659 5336 4663
rect 5370 4663 5371 4667
rect 5375 4663 5376 4667
rect 5370 4662 5376 4663
rect 5330 4658 5336 4659
rect 5332 4640 5334 4658
rect 5330 4639 5336 4640
rect 5330 4635 5331 4639
rect 5335 4635 5336 4639
rect 5330 4634 5336 4635
rect 5380 4624 5382 4685
rect 5516 4624 5518 4685
rect 5664 4625 5666 4685
rect 5662 4624 5668 4625
rect 4674 4623 4680 4624
rect 4674 4619 4675 4623
rect 4679 4619 4680 4623
rect 4674 4618 4680 4619
rect 4818 4623 4824 4624
rect 4818 4619 4819 4623
rect 4823 4619 4824 4623
rect 4818 4618 4824 4619
rect 4962 4623 4968 4624
rect 4962 4619 4963 4623
rect 4967 4619 4968 4623
rect 4962 4618 4968 4619
rect 5106 4623 5112 4624
rect 5106 4619 5107 4623
rect 5111 4619 5112 4623
rect 5106 4618 5112 4619
rect 5242 4623 5248 4624
rect 5242 4619 5243 4623
rect 5247 4619 5248 4623
rect 5242 4618 5248 4619
rect 5378 4623 5384 4624
rect 5378 4619 5379 4623
rect 5383 4619 5384 4623
rect 5378 4618 5384 4619
rect 5514 4623 5520 4624
rect 5514 4619 5515 4623
rect 5519 4619 5520 4623
rect 5662 4620 5663 4624
rect 5667 4620 5668 4624
rect 5662 4619 5668 4620
rect 5514 4618 5520 4619
rect 4702 4608 4708 4609
rect 4702 4604 4703 4608
rect 4707 4604 4708 4608
rect 4702 4603 4708 4604
rect 4846 4608 4852 4609
rect 4846 4604 4847 4608
rect 4851 4604 4852 4608
rect 4846 4603 4852 4604
rect 4990 4608 4996 4609
rect 4990 4604 4991 4608
rect 4995 4604 4996 4608
rect 4990 4603 4996 4604
rect 5134 4608 5140 4609
rect 5134 4604 5135 4608
rect 5139 4604 5140 4608
rect 5134 4603 5140 4604
rect 5270 4608 5276 4609
rect 5270 4604 5271 4608
rect 5275 4604 5276 4608
rect 5270 4603 5276 4604
rect 5406 4608 5412 4609
rect 5406 4604 5407 4608
rect 5411 4604 5412 4608
rect 5406 4603 5412 4604
rect 5542 4608 5548 4609
rect 5542 4604 5543 4608
rect 5547 4604 5548 4608
rect 5542 4603 5548 4604
rect 5662 4607 5668 4608
rect 5662 4603 5663 4607
rect 5667 4603 5668 4607
rect 4704 4579 4706 4603
rect 4848 4579 4850 4603
rect 4992 4579 4994 4603
rect 5136 4579 5138 4603
rect 5272 4579 5274 4603
rect 5408 4579 5410 4603
rect 5544 4579 5546 4603
rect 5662 4602 5668 4603
rect 5664 4579 5666 4602
rect 4671 4578 4675 4579
rect 4671 4573 4675 4574
rect 4703 4578 4707 4579
rect 4703 4573 4707 4574
rect 4807 4578 4811 4579
rect 4807 4573 4811 4574
rect 4847 4578 4851 4579
rect 4847 4573 4851 4574
rect 4943 4578 4947 4579
rect 4943 4573 4947 4574
rect 4991 4578 4995 4579
rect 4991 4573 4995 4574
rect 5079 4578 5083 4579
rect 5079 4573 5083 4574
rect 5135 4578 5139 4579
rect 5135 4573 5139 4574
rect 5271 4578 5275 4579
rect 5271 4573 5275 4574
rect 5407 4578 5411 4579
rect 5407 4573 5411 4574
rect 5543 4578 5547 4579
rect 5543 4573 5547 4574
rect 5663 4578 5667 4579
rect 5663 4573 5667 4574
rect 4672 4549 4674 4573
rect 4808 4549 4810 4573
rect 4944 4549 4946 4573
rect 5080 4549 5082 4573
rect 5664 4550 5666 4573
rect 5662 4549 5668 4550
rect 4670 4548 4676 4549
rect 4670 4544 4671 4548
rect 4675 4544 4676 4548
rect 4670 4543 4676 4544
rect 4806 4548 4812 4549
rect 4806 4544 4807 4548
rect 4811 4544 4812 4548
rect 4806 4543 4812 4544
rect 4942 4548 4948 4549
rect 4942 4544 4943 4548
rect 4947 4544 4948 4548
rect 4942 4543 4948 4544
rect 5078 4548 5084 4549
rect 5078 4544 5079 4548
rect 5083 4544 5084 4548
rect 5662 4545 5663 4549
rect 5667 4545 5668 4549
rect 5662 4544 5668 4545
rect 5078 4543 5084 4544
rect 4642 4533 4648 4534
rect 4642 4529 4643 4533
rect 4647 4529 4648 4533
rect 4642 4528 4648 4529
rect 4778 4533 4784 4534
rect 4778 4529 4779 4533
rect 4783 4529 4784 4533
rect 4778 4528 4784 4529
rect 4914 4533 4920 4534
rect 4914 4529 4915 4533
rect 4919 4529 4920 4533
rect 4914 4528 4920 4529
rect 5050 4533 5056 4534
rect 5050 4529 5051 4533
rect 5055 4529 5056 4533
rect 5050 4528 5056 4529
rect 5662 4532 5668 4533
rect 5662 4528 5663 4532
rect 5667 4528 5668 4532
rect 4594 4491 4600 4492
rect 4594 4487 4595 4491
rect 4599 4487 4600 4491
rect 4594 4486 4600 4487
rect 4644 4463 4646 4528
rect 4780 4463 4782 4528
rect 4794 4523 4800 4524
rect 4794 4519 4795 4523
rect 4799 4519 4800 4523
rect 4794 4518 4800 4519
rect 4796 4492 4798 4518
rect 4794 4491 4800 4492
rect 4794 4487 4795 4491
rect 4799 4487 4800 4491
rect 4794 4486 4800 4487
rect 4916 4463 4918 4528
rect 4930 4523 4936 4524
rect 4930 4519 4931 4523
rect 4935 4519 4936 4523
rect 4930 4518 4936 4519
rect 4932 4492 4934 4518
rect 4930 4491 4936 4492
rect 4930 4487 4931 4491
rect 4935 4487 4936 4491
rect 4930 4486 4936 4487
rect 5052 4463 5054 4528
rect 5662 4527 5668 4528
rect 5066 4523 5072 4524
rect 5066 4519 5067 4523
rect 5071 4519 5072 4523
rect 5066 4518 5072 4519
rect 5074 4523 5080 4524
rect 5074 4519 5075 4523
rect 5079 4519 5080 4523
rect 5074 4518 5080 4519
rect 5068 4492 5070 4518
rect 5066 4491 5072 4492
rect 5066 4487 5067 4491
rect 5071 4487 5072 4491
rect 5066 4486 5072 4487
rect 3839 4462 3843 4463
rect 3839 4457 3843 4458
rect 4347 4462 4351 4463
rect 4347 4457 4351 4458
rect 4483 4462 4487 4463
rect 4483 4457 4487 4458
rect 4619 4462 4623 4463
rect 4619 4457 4623 4458
rect 4643 4462 4647 4463
rect 4643 4457 4647 4458
rect 4755 4462 4759 4463
rect 4755 4457 4759 4458
rect 4779 4462 4783 4463
rect 4779 4457 4783 4458
rect 4891 4462 4895 4463
rect 4891 4457 4895 4458
rect 4915 4462 4919 4463
rect 4915 4457 4919 4458
rect 5051 4462 5055 4463
rect 5051 4457 5055 4458
rect 3798 4436 3804 4437
rect 2970 4435 2976 4436
rect 2970 4431 2971 4435
rect 2975 4431 2976 4435
rect 2970 4430 2976 4431
rect 3186 4435 3192 4436
rect 3186 4431 3187 4435
rect 3191 4431 3192 4435
rect 3186 4430 3192 4431
rect 3394 4435 3400 4436
rect 3394 4431 3395 4435
rect 3399 4431 3400 4435
rect 3394 4430 3400 4431
rect 3610 4435 3616 4436
rect 3610 4431 3611 4435
rect 3615 4431 3616 4435
rect 3798 4432 3799 4436
rect 3803 4432 3804 4436
rect 3798 4431 3804 4432
rect 3610 4430 3616 4431
rect 2998 4420 3004 4421
rect 2998 4416 2999 4420
rect 3003 4416 3004 4420
rect 2998 4415 3004 4416
rect 3214 4420 3220 4421
rect 3214 4416 3215 4420
rect 3219 4416 3220 4420
rect 3214 4415 3220 4416
rect 3422 4420 3428 4421
rect 3422 4416 3423 4420
rect 3427 4416 3428 4420
rect 3422 4415 3428 4416
rect 3638 4420 3644 4421
rect 3638 4416 3639 4420
rect 3643 4416 3644 4420
rect 3638 4415 3644 4416
rect 3798 4419 3804 4420
rect 3798 4415 3799 4419
rect 3803 4415 3804 4419
rect 3000 4379 3002 4415
rect 3216 4379 3218 4415
rect 3424 4379 3426 4415
rect 3640 4379 3642 4415
rect 3798 4414 3804 4415
rect 3800 4379 3802 4414
rect 3840 4397 3842 4457
rect 3838 4396 3844 4397
rect 4348 4396 4350 4457
rect 4466 4403 4472 4404
rect 4466 4399 4467 4403
rect 4471 4399 4472 4403
rect 4466 4398 4472 4399
rect 3838 4392 3839 4396
rect 3843 4392 3844 4396
rect 3838 4391 3844 4392
rect 4346 4395 4352 4396
rect 4346 4391 4347 4395
rect 4351 4391 4352 4395
rect 4346 4390 4352 4391
rect 4374 4380 4380 4381
rect 3838 4379 3844 4380
rect 2951 4378 2955 4379
rect 2951 4373 2955 4374
rect 2999 4378 3003 4379
rect 2999 4373 3003 4374
rect 3135 4378 3139 4379
rect 3135 4373 3139 4374
rect 3215 4378 3219 4379
rect 3215 4373 3219 4374
rect 3319 4378 3323 4379
rect 3319 4373 3323 4374
rect 3423 4378 3427 4379
rect 3423 4373 3427 4374
rect 3639 4378 3643 4379
rect 3639 4373 3643 4374
rect 3799 4378 3803 4379
rect 3838 4375 3839 4379
rect 3843 4375 3844 4379
rect 4374 4376 4375 4380
rect 4379 4376 4380 4380
rect 4374 4375 4380 4376
rect 3838 4374 3844 4375
rect 3799 4373 3803 4374
rect 2952 4349 2954 4373
rect 3136 4349 3138 4373
rect 3320 4349 3322 4373
rect 3800 4350 3802 4373
rect 3798 4349 3804 4350
rect 2950 4348 2956 4349
rect 2950 4344 2951 4348
rect 2955 4344 2956 4348
rect 2950 4343 2956 4344
rect 3134 4348 3140 4349
rect 3134 4344 3135 4348
rect 3139 4344 3140 4348
rect 3134 4343 3140 4344
rect 3318 4348 3324 4349
rect 3318 4344 3319 4348
rect 3323 4344 3324 4348
rect 3798 4345 3799 4349
rect 3803 4345 3804 4349
rect 3798 4344 3804 4345
rect 3318 4343 3324 4344
rect 3840 4335 3842 4374
rect 4376 4335 4378 4375
rect 3839 4334 3843 4335
rect 2922 4333 2928 4334
rect 2922 4329 2923 4333
rect 2927 4329 2928 4333
rect 2922 4328 2928 4329
rect 3106 4333 3112 4334
rect 3106 4329 3107 4333
rect 3111 4329 3112 4333
rect 3106 4328 3112 4329
rect 3290 4333 3296 4334
rect 3290 4329 3291 4333
rect 3295 4329 3296 4333
rect 3290 4328 3296 4329
rect 3798 4332 3804 4333
rect 3798 4328 3799 4332
rect 3803 4328 3804 4332
rect 3839 4329 3843 4330
rect 4135 4334 4139 4335
rect 4135 4329 4139 4330
rect 4271 4334 4275 4335
rect 4271 4329 4275 4330
rect 4375 4334 4379 4335
rect 4375 4329 4379 4330
rect 4407 4334 4411 4335
rect 4407 4329 4411 4330
rect 2834 4315 2840 4316
rect 2834 4311 2835 4315
rect 2839 4311 2840 4315
rect 2834 4310 2840 4311
rect 2762 4291 2768 4292
rect 2762 4287 2763 4291
rect 2767 4287 2768 4291
rect 2762 4286 2768 4287
rect 2924 4263 2926 4328
rect 2938 4323 2944 4324
rect 2938 4319 2939 4323
rect 2943 4319 2944 4323
rect 2938 4318 2944 4319
rect 2940 4292 2942 4318
rect 2938 4291 2944 4292
rect 2938 4287 2939 4291
rect 2943 4287 2944 4291
rect 2938 4286 2944 4287
rect 3108 4263 3110 4328
rect 3122 4323 3128 4324
rect 3122 4319 3123 4323
rect 3127 4319 3128 4323
rect 3122 4318 3128 4319
rect 3124 4292 3126 4318
rect 3122 4291 3128 4292
rect 3122 4287 3123 4291
rect 3127 4287 3128 4291
rect 3122 4286 3128 4287
rect 3292 4263 3294 4328
rect 3798 4327 3804 4328
rect 3306 4323 3312 4324
rect 3306 4319 3307 4323
rect 3311 4319 3312 4323
rect 3306 4318 3312 4319
rect 3308 4292 3310 4318
rect 3306 4291 3312 4292
rect 3306 4287 3307 4291
rect 3311 4287 3312 4291
rect 3306 4286 3312 4287
rect 3800 4263 3802 4327
rect 3840 4306 3842 4329
rect 3838 4305 3844 4306
rect 4136 4305 4138 4329
rect 4272 4305 4274 4329
rect 4408 4305 4410 4329
rect 3838 4301 3839 4305
rect 3843 4301 3844 4305
rect 3838 4300 3844 4301
rect 4134 4304 4140 4305
rect 4134 4300 4135 4304
rect 4139 4300 4140 4304
rect 4134 4299 4140 4300
rect 4270 4304 4276 4305
rect 4270 4300 4271 4304
rect 4275 4300 4276 4304
rect 4270 4299 4276 4300
rect 4406 4304 4412 4305
rect 4406 4300 4407 4304
rect 4411 4300 4412 4304
rect 4406 4299 4412 4300
rect 4106 4289 4112 4290
rect 3838 4288 3844 4289
rect 3838 4284 3839 4288
rect 3843 4284 3844 4288
rect 4106 4285 4107 4289
rect 4111 4285 4112 4289
rect 4106 4284 4112 4285
rect 4242 4289 4248 4290
rect 4242 4285 4243 4289
rect 4247 4285 4248 4289
rect 4242 4284 4248 4285
rect 4378 4289 4384 4290
rect 4378 4285 4379 4289
rect 4383 4285 4384 4289
rect 4378 4284 4384 4285
rect 3838 4283 3844 4284
rect 2747 4262 2751 4263
rect 2747 4257 2751 4258
rect 2763 4262 2767 4263
rect 2763 4257 2767 4258
rect 2923 4262 2927 4263
rect 2923 4257 2927 4258
rect 3019 4262 3023 4263
rect 3019 4257 3023 4258
rect 3107 4262 3111 4263
rect 3107 4257 3111 4258
rect 3283 4262 3287 4263
rect 3283 4257 3287 4258
rect 3291 4262 3295 4263
rect 3291 4257 3295 4258
rect 3799 4262 3803 4263
rect 3799 4257 3803 4258
rect 2630 4203 2636 4204
rect 2630 4199 2631 4203
rect 2635 4199 2636 4203
rect 2630 4198 2636 4199
rect 2764 4196 2766 4257
rect 2958 4239 2964 4240
rect 2958 4235 2959 4239
rect 2963 4235 2964 4239
rect 2958 4234 2964 4235
rect 2960 4204 2962 4234
rect 2958 4203 2964 4204
rect 2958 4199 2959 4203
rect 2963 4199 2964 4203
rect 2958 4198 2964 4199
rect 3020 4196 3022 4257
rect 3284 4196 3286 4257
rect 3370 4235 3376 4236
rect 3370 4231 3371 4235
rect 3375 4231 3376 4235
rect 3370 4230 3376 4231
rect 1974 4192 1975 4196
rect 1979 4192 1980 4196
rect 1974 4191 1980 4192
rect 1994 4195 2000 4196
rect 1994 4191 1995 4195
rect 1999 4191 2000 4195
rect 1994 4190 2000 4191
rect 2242 4195 2248 4196
rect 2242 4191 2243 4195
rect 2247 4191 2248 4195
rect 2242 4190 2248 4191
rect 2506 4195 2512 4196
rect 2506 4191 2507 4195
rect 2511 4191 2512 4195
rect 2506 4190 2512 4191
rect 2762 4195 2768 4196
rect 2762 4191 2763 4195
rect 2767 4191 2768 4195
rect 2762 4190 2768 4191
rect 3018 4195 3024 4196
rect 3018 4191 3019 4195
rect 3023 4191 3024 4195
rect 3018 4190 3024 4191
rect 3282 4195 3288 4196
rect 3282 4191 3283 4195
rect 3287 4191 3288 4195
rect 3282 4190 3288 4191
rect 2022 4180 2028 4181
rect 1974 4179 1980 4180
rect 1974 4175 1975 4179
rect 1979 4175 1980 4179
rect 2022 4176 2023 4180
rect 2027 4176 2028 4180
rect 2022 4175 2028 4176
rect 2270 4180 2276 4181
rect 2270 4176 2271 4180
rect 2275 4176 2276 4180
rect 2270 4175 2276 4176
rect 2534 4180 2540 4181
rect 2534 4176 2535 4180
rect 2539 4176 2540 4180
rect 2534 4175 2540 4176
rect 2790 4180 2796 4181
rect 2790 4176 2791 4180
rect 2795 4176 2796 4180
rect 2790 4175 2796 4176
rect 3046 4180 3052 4181
rect 3046 4176 3047 4180
rect 3051 4176 3052 4180
rect 3046 4175 3052 4176
rect 3310 4180 3316 4181
rect 3310 4176 3311 4180
rect 3315 4176 3316 4180
rect 3310 4175 3316 4176
rect 1974 4174 1980 4175
rect 1946 4139 1952 4140
rect 1976 4139 1978 4174
rect 2024 4139 2026 4175
rect 2272 4139 2274 4175
rect 2536 4139 2538 4175
rect 2792 4139 2794 4175
rect 3048 4139 3050 4175
rect 3312 4139 3314 4175
rect 1946 4135 1947 4139
rect 1951 4135 1952 4139
rect 1946 4134 1952 4135
rect 1975 4138 1979 4139
rect 1975 4133 1979 4134
rect 2023 4138 2027 4139
rect 2023 4133 2027 4134
rect 2271 4138 2275 4139
rect 2271 4133 2275 4134
rect 2535 4138 2539 4139
rect 2535 4133 2539 4134
rect 2791 4138 2795 4139
rect 2791 4133 2795 4134
rect 3047 4138 3051 4139
rect 3047 4133 3051 4134
rect 3135 4138 3139 4139
rect 3135 4133 3139 4134
rect 3271 4138 3275 4139
rect 3271 4133 3275 4134
rect 3311 4138 3315 4139
rect 3311 4133 3315 4134
rect 1787 4114 1791 4115
rect 1787 4109 1791 4110
rect 1935 4114 1939 4115
rect 1976 4110 1978 4133
rect 1935 4109 1939 4110
rect 1974 4109 1980 4110
rect 3136 4109 3138 4133
rect 3272 4109 3274 4133
rect 1778 4091 1784 4092
rect 1778 4087 1779 4091
rect 1783 4087 1784 4091
rect 1778 4086 1784 4087
rect 1788 4048 1790 4109
rect 1936 4049 1938 4109
rect 1974 4105 1975 4109
rect 1979 4105 1980 4109
rect 1974 4104 1980 4105
rect 3134 4108 3140 4109
rect 3134 4104 3135 4108
rect 3139 4104 3140 4108
rect 3134 4103 3140 4104
rect 3270 4108 3276 4109
rect 3270 4104 3271 4108
rect 3275 4104 3276 4108
rect 3270 4103 3276 4104
rect 3106 4093 3112 4094
rect 1974 4092 1980 4093
rect 1974 4088 1975 4092
rect 1979 4088 1980 4092
rect 3106 4089 3107 4093
rect 3111 4089 3112 4093
rect 3106 4088 3112 4089
rect 3242 4093 3248 4094
rect 3242 4089 3243 4093
rect 3247 4089 3248 4093
rect 3242 4088 3248 4089
rect 1974 4087 1980 4088
rect 1934 4048 1940 4049
rect 1650 4047 1656 4048
rect 1650 4043 1651 4047
rect 1655 4043 1656 4047
rect 1650 4042 1656 4043
rect 1786 4047 1792 4048
rect 1786 4043 1787 4047
rect 1791 4043 1792 4047
rect 1934 4044 1935 4048
rect 1939 4044 1940 4048
rect 1934 4043 1940 4044
rect 1786 4042 1792 4043
rect 1678 4032 1684 4033
rect 1678 4028 1679 4032
rect 1683 4028 1684 4032
rect 1678 4027 1684 4028
rect 1814 4032 1820 4033
rect 1814 4028 1815 4032
rect 1819 4028 1820 4032
rect 1814 4027 1820 4028
rect 1934 4031 1940 4032
rect 1934 4027 1935 4031
rect 1939 4027 1940 4031
rect 1680 4003 1682 4027
rect 1816 4003 1818 4027
rect 1934 4026 1940 4027
rect 1936 4003 1938 4026
rect 1679 4002 1683 4003
rect 1679 3997 1683 3998
rect 1815 4002 1819 4003
rect 1815 3997 1819 3998
rect 1935 4002 1939 4003
rect 1935 3997 1939 3998
rect 1816 3973 1818 3997
rect 1936 3974 1938 3997
rect 1934 3973 1940 3974
rect 1814 3972 1820 3973
rect 1814 3968 1815 3972
rect 1819 3968 1820 3972
rect 1934 3969 1935 3973
rect 1939 3969 1940 3973
rect 1934 3968 1940 3969
rect 1814 3967 1820 3968
rect 1786 3957 1792 3958
rect 1786 3953 1787 3957
rect 1791 3953 1792 3957
rect 1786 3952 1792 3953
rect 1934 3956 1940 3957
rect 1934 3952 1935 3956
rect 1939 3952 1940 3956
rect 1638 3915 1644 3916
rect 1638 3911 1639 3915
rect 1643 3911 1644 3915
rect 1638 3910 1644 3911
rect 1788 3891 1790 3952
rect 1934 3951 1940 3952
rect 1802 3947 1808 3948
rect 1802 3943 1803 3947
rect 1807 3943 1808 3947
rect 1802 3942 1808 3943
rect 1890 3947 1896 3948
rect 1890 3943 1891 3947
rect 1895 3943 1896 3947
rect 1890 3942 1896 3943
rect 1804 3916 1806 3942
rect 1802 3915 1808 3916
rect 1802 3911 1803 3915
rect 1807 3911 1808 3915
rect 1802 3910 1808 3911
rect 1371 3890 1375 3891
rect 1371 3885 1375 3886
rect 1499 3890 1503 3891
rect 1499 3885 1503 3886
rect 1587 3890 1591 3891
rect 1587 3885 1591 3886
rect 1787 3890 1791 3891
rect 1787 3885 1791 3886
rect 1334 3867 1340 3868
rect 1334 3863 1335 3867
rect 1339 3863 1340 3867
rect 1334 3862 1340 3863
rect 1336 3832 1338 3862
rect 1242 3831 1248 3832
rect 1242 3827 1243 3831
rect 1247 3827 1248 3831
rect 1242 3826 1248 3827
rect 1334 3831 1340 3832
rect 1334 3827 1335 3831
rect 1339 3827 1340 3831
rect 1334 3826 1340 3827
rect 1500 3824 1502 3885
rect 1788 3824 1790 3885
rect 1892 3868 1894 3942
rect 1914 3911 1920 3912
rect 1914 3907 1915 3911
rect 1919 3907 1920 3911
rect 1914 3906 1920 3907
rect 1890 3867 1896 3868
rect 1890 3863 1891 3867
rect 1895 3863 1896 3867
rect 1890 3862 1896 3863
rect 1916 3832 1918 3906
rect 1936 3891 1938 3951
rect 1976 3935 1978 4087
rect 3108 3935 3110 4088
rect 3194 4075 3200 4076
rect 3194 4071 3195 4075
rect 3199 4071 3200 4075
rect 3194 4070 3200 4071
rect 3196 4052 3198 4070
rect 3194 4051 3200 4052
rect 3194 4047 3195 4051
rect 3199 4047 3200 4051
rect 3194 4046 3200 4047
rect 3244 3935 3246 4088
rect 3372 4084 3374 4230
rect 3800 4197 3802 4257
rect 3840 4211 3842 4283
rect 4108 4211 4110 4284
rect 4234 4279 4240 4280
rect 4234 4275 4235 4279
rect 4239 4275 4240 4279
rect 4234 4274 4240 4275
rect 3839 4210 3843 4211
rect 3839 4205 3843 4206
rect 3971 4210 3975 4211
rect 3971 4205 3975 4206
rect 4107 4210 4111 4211
rect 4107 4205 4111 4206
rect 3798 4196 3804 4197
rect 3798 4192 3799 4196
rect 3803 4192 3804 4196
rect 3798 4191 3804 4192
rect 3798 4179 3804 4180
rect 3798 4175 3799 4179
rect 3803 4175 3804 4179
rect 3798 4174 3804 4175
rect 3800 4139 3802 4174
rect 3840 4145 3842 4205
rect 3838 4144 3844 4145
rect 3972 4144 3974 4205
rect 4058 4183 4064 4184
rect 4058 4178 4059 4183
rect 4063 4178 4064 4183
rect 4059 4175 4063 4176
rect 4108 4144 4110 4205
rect 4236 4188 4238 4274
rect 4244 4211 4246 4284
rect 4250 4279 4256 4280
rect 4250 4275 4251 4279
rect 4255 4275 4256 4279
rect 4250 4274 4256 4275
rect 4252 4248 4254 4274
rect 4330 4271 4336 4272
rect 4330 4267 4331 4271
rect 4335 4267 4336 4271
rect 4330 4266 4336 4267
rect 4332 4248 4334 4266
rect 4250 4247 4256 4248
rect 4250 4243 4251 4247
rect 4255 4243 4256 4247
rect 4250 4242 4256 4243
rect 4330 4247 4336 4248
rect 4330 4243 4331 4247
rect 4335 4243 4336 4247
rect 4330 4242 4336 4243
rect 4380 4211 4382 4284
rect 4468 4248 4470 4398
rect 4484 4396 4486 4457
rect 4620 4396 4622 4457
rect 4756 4396 4758 4457
rect 4892 4396 4894 4457
rect 5076 4440 5078 4518
rect 5664 4463 5666 4527
rect 5663 4462 5667 4463
rect 5663 4457 5667 4458
rect 5074 4439 5080 4440
rect 5074 4435 5075 4439
rect 5079 4435 5080 4439
rect 5074 4434 5080 4435
rect 5664 4397 5666 4457
rect 5662 4396 5668 4397
rect 4482 4395 4488 4396
rect 4482 4391 4483 4395
rect 4487 4391 4488 4395
rect 4482 4390 4488 4391
rect 4618 4395 4624 4396
rect 4618 4391 4619 4395
rect 4623 4391 4624 4395
rect 4618 4390 4624 4391
rect 4754 4395 4760 4396
rect 4754 4391 4755 4395
rect 4759 4391 4760 4395
rect 4754 4390 4760 4391
rect 4890 4395 4896 4396
rect 4890 4391 4891 4395
rect 4895 4391 4896 4395
rect 5662 4392 5663 4396
rect 5667 4392 5668 4396
rect 5662 4391 5668 4392
rect 4890 4390 4896 4391
rect 4510 4380 4516 4381
rect 4510 4376 4511 4380
rect 4515 4376 4516 4380
rect 4510 4375 4516 4376
rect 4646 4380 4652 4381
rect 4646 4376 4647 4380
rect 4651 4376 4652 4380
rect 4646 4375 4652 4376
rect 4782 4380 4788 4381
rect 4782 4376 4783 4380
rect 4787 4376 4788 4380
rect 4782 4375 4788 4376
rect 4918 4380 4924 4381
rect 4918 4376 4919 4380
rect 4923 4376 4924 4380
rect 4918 4375 4924 4376
rect 5662 4379 5668 4380
rect 5662 4375 5663 4379
rect 5667 4375 5668 4379
rect 4512 4335 4514 4375
rect 4648 4335 4650 4375
rect 4784 4335 4786 4375
rect 4920 4335 4922 4375
rect 5662 4374 5668 4375
rect 5664 4335 5666 4374
rect 4511 4334 4515 4335
rect 4511 4329 4515 4330
rect 4543 4334 4547 4335
rect 4543 4329 4547 4330
rect 4647 4334 4651 4335
rect 4647 4329 4651 4330
rect 4679 4334 4683 4335
rect 4679 4329 4683 4330
rect 4783 4334 4787 4335
rect 4783 4329 4787 4330
rect 4919 4334 4923 4335
rect 4919 4329 4923 4330
rect 5663 4334 5667 4335
rect 5663 4329 5667 4330
rect 4544 4305 4546 4329
rect 4680 4305 4682 4329
rect 5664 4306 5666 4329
rect 5662 4305 5668 4306
rect 4542 4304 4548 4305
rect 4542 4300 4543 4304
rect 4547 4300 4548 4304
rect 4542 4299 4548 4300
rect 4678 4304 4684 4305
rect 4678 4300 4679 4304
rect 4683 4300 4684 4304
rect 5662 4301 5663 4305
rect 5667 4301 5668 4305
rect 5662 4300 5668 4301
rect 4678 4299 4684 4300
rect 4514 4289 4520 4290
rect 4514 4285 4515 4289
rect 4519 4285 4520 4289
rect 4514 4284 4520 4285
rect 4650 4289 4656 4290
rect 4650 4285 4651 4289
rect 4655 4285 4656 4289
rect 4650 4284 4656 4285
rect 5662 4288 5668 4289
rect 5662 4284 5663 4288
rect 5667 4284 5668 4288
rect 4466 4247 4472 4248
rect 4466 4243 4467 4247
rect 4471 4243 4472 4247
rect 4466 4242 4472 4243
rect 4516 4211 4518 4284
rect 4530 4279 4536 4280
rect 4530 4275 4531 4279
rect 4535 4275 4536 4279
rect 4530 4274 4536 4275
rect 4532 4248 4534 4274
rect 4530 4247 4536 4248
rect 4530 4243 4531 4247
rect 4535 4243 4536 4247
rect 4530 4242 4536 4243
rect 4652 4211 4654 4284
rect 5662 4283 5668 4284
rect 4666 4279 4672 4280
rect 4666 4275 4667 4279
rect 4671 4275 4672 4279
rect 4666 4274 4672 4275
rect 4668 4248 4670 4274
rect 4666 4247 4672 4248
rect 4666 4243 4667 4247
rect 4671 4243 4672 4247
rect 4666 4242 4672 4243
rect 5664 4211 5666 4283
rect 4243 4210 4247 4211
rect 4243 4205 4247 4206
rect 4379 4210 4383 4211
rect 4379 4205 4383 4206
rect 4515 4210 4519 4211
rect 4515 4205 4519 4206
rect 4651 4210 4655 4211
rect 4651 4205 4655 4206
rect 5663 4210 5667 4211
rect 5663 4205 5667 4206
rect 4234 4187 4240 4188
rect 4234 4183 4235 4187
rect 4239 4183 4240 4187
rect 4234 4182 4240 4183
rect 4244 4144 4246 4205
rect 4282 4151 4288 4152
rect 4282 4147 4283 4151
rect 4287 4147 4288 4151
rect 4282 4146 4288 4147
rect 3838 4140 3839 4144
rect 3843 4140 3844 4144
rect 3838 4139 3844 4140
rect 3970 4143 3976 4144
rect 3970 4139 3971 4143
rect 3975 4139 3976 4143
rect 3407 4138 3411 4139
rect 3407 4133 3411 4134
rect 3543 4138 3547 4139
rect 3543 4133 3547 4134
rect 3679 4138 3683 4139
rect 3679 4133 3683 4134
rect 3799 4138 3803 4139
rect 3970 4138 3976 4139
rect 4106 4143 4112 4144
rect 4106 4139 4107 4143
rect 4111 4139 4112 4143
rect 4106 4138 4112 4139
rect 4242 4143 4248 4144
rect 4242 4139 4243 4143
rect 4247 4139 4248 4143
rect 4242 4138 4248 4139
rect 3799 4133 3803 4134
rect 3408 4109 3410 4133
rect 3544 4109 3546 4133
rect 3680 4109 3682 4133
rect 3800 4110 3802 4133
rect 3998 4128 4004 4129
rect 3838 4127 3844 4128
rect 3838 4123 3839 4127
rect 3843 4123 3844 4127
rect 3998 4124 3999 4128
rect 4003 4124 4004 4128
rect 3998 4123 4004 4124
rect 4134 4128 4140 4129
rect 4134 4124 4135 4128
rect 4139 4124 4140 4128
rect 4134 4123 4140 4124
rect 4270 4128 4276 4129
rect 4270 4124 4271 4128
rect 4275 4124 4276 4128
rect 4270 4123 4276 4124
rect 3838 4122 3844 4123
rect 3798 4109 3804 4110
rect 3406 4108 3412 4109
rect 3406 4104 3407 4108
rect 3411 4104 3412 4108
rect 3406 4103 3412 4104
rect 3542 4108 3548 4109
rect 3542 4104 3543 4108
rect 3547 4104 3548 4108
rect 3542 4103 3548 4104
rect 3678 4108 3684 4109
rect 3678 4104 3679 4108
rect 3683 4104 3684 4108
rect 3798 4105 3799 4109
rect 3803 4105 3804 4109
rect 3798 4104 3804 4105
rect 3678 4103 3684 4104
rect 3378 4093 3384 4094
rect 3378 4089 3379 4093
rect 3383 4089 3384 4093
rect 3378 4088 3384 4089
rect 3514 4093 3520 4094
rect 3514 4089 3515 4093
rect 3519 4089 3520 4093
rect 3514 4088 3520 4089
rect 3650 4093 3656 4094
rect 3650 4089 3651 4093
rect 3655 4089 3656 4093
rect 3650 4088 3656 4089
rect 3798 4092 3804 4093
rect 3798 4088 3799 4092
rect 3803 4088 3804 4092
rect 3258 4083 3264 4084
rect 3258 4079 3259 4083
rect 3263 4079 3264 4083
rect 3258 4078 3264 4079
rect 3370 4083 3376 4084
rect 3370 4079 3371 4083
rect 3375 4079 3376 4083
rect 3370 4078 3376 4079
rect 3260 4052 3262 4078
rect 3258 4051 3264 4052
rect 3258 4047 3259 4051
rect 3263 4047 3264 4051
rect 3258 4046 3264 4047
rect 3380 3935 3382 4088
rect 3516 3935 3518 4088
rect 3652 3935 3654 4088
rect 3798 4087 3804 4088
rect 3738 4051 3744 4052
rect 3738 4047 3739 4051
rect 3743 4047 3744 4051
rect 3738 4046 3744 4047
rect 3740 4020 3742 4046
rect 3738 4019 3744 4020
rect 3738 4015 3739 4019
rect 3743 4015 3744 4019
rect 3738 4014 3744 4015
rect 3778 3939 3784 3940
rect 3778 3935 3779 3939
rect 3783 3935 3784 3939
rect 3800 3935 3802 4087
rect 3840 4075 3842 4122
rect 4000 4075 4002 4123
rect 4136 4075 4138 4123
rect 4272 4075 4274 4123
rect 3839 4074 3843 4075
rect 3839 4069 3843 4070
rect 3887 4074 3891 4075
rect 3887 4069 3891 4070
rect 3999 4074 4003 4075
rect 3999 4069 4003 4070
rect 4023 4074 4027 4075
rect 4023 4069 4027 4070
rect 4135 4074 4139 4075
rect 4135 4069 4139 4070
rect 4159 4074 4163 4075
rect 4159 4069 4163 4070
rect 4271 4074 4275 4075
rect 4271 4069 4275 4070
rect 3840 4046 3842 4069
rect 3838 4045 3844 4046
rect 3888 4045 3890 4069
rect 4024 4045 4026 4069
rect 4160 4045 4162 4069
rect 3838 4041 3839 4045
rect 3843 4041 3844 4045
rect 3838 4040 3844 4041
rect 3886 4044 3892 4045
rect 3886 4040 3887 4044
rect 3891 4040 3892 4044
rect 3886 4039 3892 4040
rect 4022 4044 4028 4045
rect 4022 4040 4023 4044
rect 4027 4040 4028 4044
rect 4022 4039 4028 4040
rect 4158 4044 4164 4045
rect 4158 4040 4159 4044
rect 4163 4040 4164 4044
rect 4158 4039 4164 4040
rect 3858 4029 3864 4030
rect 3838 4028 3844 4029
rect 3838 4024 3839 4028
rect 3843 4024 3844 4028
rect 3858 4025 3859 4029
rect 3863 4025 3864 4029
rect 3858 4024 3864 4025
rect 3994 4029 4000 4030
rect 3994 4025 3995 4029
rect 3999 4025 4000 4029
rect 3994 4024 4000 4025
rect 4130 4029 4136 4030
rect 4130 4025 4131 4029
rect 4135 4025 4136 4029
rect 4130 4024 4136 4025
rect 4266 4029 4272 4030
rect 4266 4025 4267 4029
rect 4271 4025 4272 4029
rect 4266 4024 4272 4025
rect 3838 4023 3844 4024
rect 3840 3963 3842 4023
rect 3860 3963 3862 4024
rect 3996 3963 3998 4024
rect 4002 4019 4008 4020
rect 4002 4015 4003 4019
rect 4007 4015 4008 4019
rect 4002 4014 4008 4015
rect 4004 3988 4006 4014
rect 4082 4011 4088 4012
rect 4082 4007 4083 4011
rect 4087 4007 4088 4011
rect 4082 4006 4088 4007
rect 4084 3988 4086 4006
rect 4002 3987 4008 3988
rect 4002 3983 4003 3987
rect 4007 3983 4008 3987
rect 4002 3982 4008 3983
rect 4082 3987 4088 3988
rect 4082 3983 4083 3987
rect 4087 3983 4088 3987
rect 4082 3982 4088 3983
rect 4122 3987 4128 3988
rect 4122 3983 4123 3987
rect 4127 3983 4128 3987
rect 4122 3982 4128 3983
rect 3839 3962 3843 3963
rect 3839 3957 3843 3958
rect 3859 3962 3863 3963
rect 3859 3957 3863 3958
rect 3995 3962 3999 3963
rect 3995 3957 3999 3958
rect 1975 3934 1979 3935
rect 1975 3929 1979 3930
rect 1995 3934 1999 3935
rect 1995 3929 1999 3930
rect 2403 3934 2407 3935
rect 2403 3929 2407 3930
rect 2827 3934 2831 3935
rect 2827 3929 2831 3930
rect 3107 3934 3111 3935
rect 3107 3929 3111 3930
rect 3243 3934 3247 3935
rect 3243 3929 3247 3930
rect 3251 3934 3255 3935
rect 3251 3929 3255 3930
rect 3379 3934 3383 3935
rect 3379 3929 3383 3930
rect 3515 3934 3519 3935
rect 3515 3929 3519 3930
rect 3651 3934 3655 3935
rect 3778 3934 3784 3935
rect 3799 3934 3803 3935
rect 3651 3929 3655 3930
rect 1935 3890 1939 3891
rect 1935 3885 1939 3886
rect 1914 3831 1920 3832
rect 1914 3827 1915 3831
rect 1919 3827 1920 3831
rect 1914 3826 1920 3827
rect 1936 3825 1938 3885
rect 1976 3869 1978 3929
rect 1974 3868 1980 3869
rect 1996 3868 1998 3929
rect 2082 3875 2088 3876
rect 2082 3871 2083 3875
rect 2087 3871 2088 3875
rect 2082 3870 2088 3871
rect 1974 3864 1975 3868
rect 1979 3864 1980 3868
rect 1974 3863 1980 3864
rect 1994 3867 2000 3868
rect 1994 3863 1995 3867
rect 1999 3863 2000 3867
rect 1994 3862 2000 3863
rect 2022 3852 2028 3853
rect 1974 3851 1980 3852
rect 1974 3847 1975 3851
rect 1979 3847 1980 3851
rect 2022 3848 2023 3852
rect 2027 3848 2028 3852
rect 2022 3847 2028 3848
rect 1974 3846 1980 3847
rect 1934 3824 1940 3825
rect 898 3823 904 3824
rect 898 3819 899 3823
rect 903 3819 904 3823
rect 898 3818 904 3819
rect 1194 3823 1200 3824
rect 1194 3819 1195 3823
rect 1199 3819 1200 3823
rect 1194 3818 1200 3819
rect 1498 3823 1504 3824
rect 1498 3819 1499 3823
rect 1503 3819 1504 3823
rect 1498 3818 1504 3819
rect 1786 3823 1792 3824
rect 1786 3819 1787 3823
rect 1791 3819 1792 3823
rect 1934 3820 1935 3824
rect 1939 3820 1940 3824
rect 1976 3823 1978 3846
rect 2024 3823 2026 3847
rect 1934 3819 1940 3820
rect 1975 3822 1979 3823
rect 1786 3818 1792 3819
rect 1975 3817 1979 3818
rect 2023 3822 2027 3823
rect 2023 3817 2027 3818
rect 926 3808 932 3809
rect 926 3804 927 3808
rect 931 3804 932 3808
rect 926 3803 932 3804
rect 1222 3808 1228 3809
rect 1222 3804 1223 3808
rect 1227 3804 1228 3808
rect 1222 3803 1228 3804
rect 1526 3808 1532 3809
rect 1526 3804 1527 3808
rect 1531 3804 1532 3808
rect 1526 3803 1532 3804
rect 1814 3808 1820 3809
rect 1814 3804 1815 3808
rect 1819 3804 1820 3808
rect 1814 3803 1820 3804
rect 1934 3807 1940 3808
rect 1934 3803 1935 3807
rect 1939 3803 1940 3807
rect 928 3767 930 3803
rect 1224 3767 1226 3803
rect 1528 3767 1530 3803
rect 1816 3767 1818 3803
rect 1934 3802 1940 3803
rect 1936 3767 1938 3802
rect 1976 3794 1978 3817
rect 1974 3793 1980 3794
rect 2024 3793 2026 3817
rect 1974 3789 1975 3793
rect 1979 3789 1980 3793
rect 1974 3788 1980 3789
rect 2022 3792 2028 3793
rect 2022 3788 2023 3792
rect 2027 3788 2028 3792
rect 2022 3787 2028 3788
rect 1994 3777 2000 3778
rect 1974 3776 1980 3777
rect 1974 3772 1975 3776
rect 1979 3772 1980 3776
rect 1994 3773 1995 3777
rect 1999 3773 2000 3777
rect 1994 3772 2000 3773
rect 1974 3771 1980 3772
rect 927 3766 931 3767
rect 927 3761 931 3762
rect 1063 3766 1067 3767
rect 1063 3761 1067 3762
rect 1223 3766 1227 3767
rect 1223 3761 1227 3762
rect 1343 3766 1347 3767
rect 1343 3761 1347 3762
rect 1527 3766 1531 3767
rect 1527 3761 1531 3762
rect 1815 3766 1819 3767
rect 1815 3761 1819 3762
rect 1935 3766 1939 3767
rect 1935 3761 1939 3762
rect 1064 3737 1066 3761
rect 1344 3737 1346 3761
rect 1936 3738 1938 3761
rect 1934 3737 1940 3738
rect 1062 3736 1068 3737
rect 1062 3732 1063 3736
rect 1067 3732 1068 3736
rect 1062 3731 1068 3732
rect 1342 3736 1348 3737
rect 1342 3732 1343 3736
rect 1347 3732 1348 3736
rect 1934 3733 1935 3737
rect 1939 3733 1940 3737
rect 1934 3732 1940 3733
rect 1342 3731 1348 3732
rect 1034 3721 1040 3722
rect 1034 3717 1035 3721
rect 1039 3717 1040 3721
rect 1034 3716 1040 3717
rect 1314 3721 1320 3722
rect 1314 3717 1315 3721
rect 1319 3717 1320 3721
rect 1314 3716 1320 3717
rect 1934 3720 1940 3721
rect 1934 3716 1935 3720
rect 1939 3716 1940 3720
rect 850 3679 856 3680
rect 850 3675 851 3679
rect 855 3675 856 3679
rect 850 3674 856 3675
rect 1036 3639 1038 3716
rect 1202 3679 1208 3680
rect 1202 3675 1203 3679
rect 1207 3675 1208 3679
rect 1202 3674 1208 3675
rect 635 3638 639 3639
rect 635 3633 639 3634
rect 763 3638 767 3639
rect 763 3633 767 3634
rect 779 3638 783 3639
rect 779 3633 783 3634
rect 923 3638 927 3639
rect 923 3633 927 3634
rect 1035 3638 1039 3639
rect 1035 3633 1039 3634
rect 1067 3638 1071 3639
rect 1067 3633 1071 3634
rect 594 3615 600 3616
rect 594 3611 595 3615
rect 599 3611 600 3615
rect 594 3610 600 3611
rect 636 3572 638 3633
rect 762 3615 768 3616
rect 762 3611 763 3615
rect 767 3611 768 3615
rect 762 3610 768 3611
rect 764 3580 766 3610
rect 762 3579 768 3580
rect 762 3575 763 3579
rect 767 3575 768 3579
rect 762 3574 768 3575
rect 780 3572 782 3633
rect 898 3579 904 3580
rect 898 3575 899 3579
rect 903 3575 904 3579
rect 898 3574 904 3575
rect 110 3568 111 3572
rect 115 3568 116 3572
rect 110 3567 116 3568
rect 490 3571 496 3572
rect 490 3567 491 3571
rect 495 3567 496 3571
rect 490 3566 496 3567
rect 634 3571 640 3572
rect 634 3567 635 3571
rect 639 3567 640 3571
rect 634 3566 640 3567
rect 778 3571 784 3572
rect 778 3567 779 3571
rect 783 3567 784 3571
rect 778 3566 784 3567
rect 518 3556 524 3557
rect 110 3555 116 3556
rect 110 3551 111 3555
rect 115 3551 116 3555
rect 518 3552 519 3556
rect 523 3552 524 3556
rect 518 3551 524 3552
rect 662 3556 668 3557
rect 662 3552 663 3556
rect 667 3552 668 3556
rect 662 3551 668 3552
rect 806 3556 812 3557
rect 806 3552 807 3556
rect 811 3552 812 3556
rect 806 3551 812 3552
rect 110 3550 116 3551
rect 112 3507 114 3550
rect 520 3507 522 3551
rect 664 3507 666 3551
rect 808 3507 810 3551
rect 111 3506 115 3507
rect 111 3501 115 3502
rect 431 3506 435 3507
rect 431 3501 435 3502
rect 519 3506 523 3507
rect 519 3501 523 3502
rect 567 3506 571 3507
rect 567 3501 571 3502
rect 663 3506 667 3507
rect 663 3501 667 3502
rect 703 3506 707 3507
rect 703 3501 707 3502
rect 807 3506 811 3507
rect 807 3501 811 3502
rect 839 3506 843 3507
rect 839 3501 843 3502
rect 112 3478 114 3501
rect 110 3477 116 3478
rect 432 3477 434 3501
rect 568 3477 570 3501
rect 704 3477 706 3501
rect 840 3477 842 3501
rect 110 3473 111 3477
rect 115 3473 116 3477
rect 110 3472 116 3473
rect 430 3476 436 3477
rect 430 3472 431 3476
rect 435 3472 436 3476
rect 430 3471 436 3472
rect 566 3476 572 3477
rect 566 3472 567 3476
rect 571 3472 572 3476
rect 566 3471 572 3472
rect 702 3476 708 3477
rect 702 3472 703 3476
rect 707 3472 708 3476
rect 702 3471 708 3472
rect 838 3476 844 3477
rect 838 3472 839 3476
rect 843 3472 844 3476
rect 838 3471 844 3472
rect 402 3461 408 3462
rect 110 3460 116 3461
rect 110 3456 111 3460
rect 115 3456 116 3460
rect 402 3457 403 3461
rect 407 3457 408 3461
rect 402 3456 408 3457
rect 538 3461 544 3462
rect 538 3457 539 3461
rect 543 3457 544 3461
rect 538 3456 544 3457
rect 674 3461 680 3462
rect 674 3457 675 3461
rect 679 3457 680 3461
rect 674 3456 680 3457
rect 810 3461 816 3462
rect 810 3457 811 3461
rect 815 3457 816 3461
rect 810 3456 816 3457
rect 110 3455 116 3456
rect 112 3387 114 3455
rect 404 3387 406 3456
rect 446 3419 452 3420
rect 446 3415 447 3419
rect 451 3415 452 3419
rect 446 3414 452 3415
rect 111 3386 115 3387
rect 111 3381 115 3382
rect 323 3386 327 3387
rect 323 3381 327 3382
rect 403 3386 407 3387
rect 403 3381 407 3382
rect 112 3321 114 3381
rect 110 3320 116 3321
rect 324 3320 326 3381
rect 448 3328 450 3414
rect 540 3387 542 3456
rect 618 3451 624 3452
rect 618 3447 619 3451
rect 623 3447 624 3451
rect 618 3446 624 3447
rect 620 3420 622 3446
rect 618 3419 624 3420
rect 618 3415 619 3419
rect 623 3415 624 3419
rect 618 3414 624 3415
rect 676 3387 678 3456
rect 690 3451 696 3452
rect 690 3447 691 3451
rect 695 3447 696 3451
rect 690 3446 696 3447
rect 692 3420 694 3446
rect 690 3419 696 3420
rect 690 3415 691 3419
rect 695 3415 696 3419
rect 690 3414 696 3415
rect 812 3387 814 3456
rect 818 3451 824 3452
rect 818 3447 819 3451
rect 823 3447 824 3451
rect 818 3446 824 3447
rect 459 3386 463 3387
rect 459 3381 463 3382
rect 539 3386 543 3387
rect 539 3381 543 3382
rect 595 3386 599 3387
rect 595 3381 599 3382
rect 675 3386 679 3387
rect 675 3381 679 3382
rect 731 3386 735 3387
rect 731 3381 735 3382
rect 811 3386 815 3387
rect 811 3381 815 3382
rect 446 3327 452 3328
rect 446 3323 447 3327
rect 451 3323 452 3327
rect 446 3322 452 3323
rect 460 3320 462 3381
rect 562 3363 568 3364
rect 562 3359 563 3363
rect 567 3359 568 3363
rect 562 3358 568 3359
rect 110 3316 111 3320
rect 115 3316 116 3320
rect 110 3315 116 3316
rect 322 3319 328 3320
rect 322 3315 323 3319
rect 327 3315 328 3319
rect 322 3314 328 3315
rect 458 3319 464 3320
rect 458 3315 459 3319
rect 463 3315 464 3319
rect 458 3314 464 3315
rect 350 3304 356 3305
rect 110 3303 116 3304
rect 110 3299 111 3303
rect 115 3299 116 3303
rect 350 3300 351 3304
rect 355 3300 356 3304
rect 350 3299 356 3300
rect 486 3304 492 3305
rect 486 3300 487 3304
rect 491 3300 492 3304
rect 486 3299 492 3300
rect 110 3298 116 3299
rect 112 3267 114 3298
rect 352 3267 354 3299
rect 488 3267 490 3299
rect 111 3266 115 3267
rect 111 3261 115 3262
rect 159 3266 163 3267
rect 159 3261 163 3262
rect 335 3266 339 3267
rect 335 3261 339 3262
rect 351 3266 355 3267
rect 351 3261 355 3262
rect 487 3266 491 3267
rect 487 3261 491 3262
rect 543 3266 547 3267
rect 543 3261 547 3262
rect 112 3238 114 3261
rect 110 3237 116 3238
rect 160 3237 162 3261
rect 336 3237 338 3261
rect 544 3237 546 3261
rect 110 3233 111 3237
rect 115 3233 116 3237
rect 110 3232 116 3233
rect 158 3236 164 3237
rect 158 3232 159 3236
rect 163 3232 164 3236
rect 158 3231 164 3232
rect 334 3236 340 3237
rect 334 3232 335 3236
rect 339 3232 340 3236
rect 334 3231 340 3232
rect 542 3236 548 3237
rect 542 3232 543 3236
rect 547 3232 548 3236
rect 542 3231 548 3232
rect 130 3221 136 3222
rect 110 3220 116 3221
rect 110 3216 111 3220
rect 115 3216 116 3220
rect 130 3217 131 3221
rect 135 3217 136 3221
rect 130 3216 136 3217
rect 306 3221 312 3222
rect 306 3217 307 3221
rect 311 3217 312 3221
rect 306 3216 312 3217
rect 514 3221 520 3222
rect 514 3217 515 3221
rect 519 3217 520 3221
rect 514 3216 520 3217
rect 110 3215 116 3216
rect 112 3139 114 3215
rect 132 3139 134 3216
rect 226 3179 232 3180
rect 226 3175 227 3179
rect 231 3175 232 3179
rect 226 3174 232 3175
rect 111 3138 115 3139
rect 111 3133 115 3134
rect 131 3138 135 3139
rect 131 3133 135 3134
rect 112 3073 114 3133
rect 110 3072 116 3073
rect 132 3072 134 3133
rect 228 3080 230 3174
rect 308 3139 310 3216
rect 322 3211 328 3212
rect 322 3207 323 3211
rect 327 3207 328 3211
rect 322 3206 328 3207
rect 324 3180 326 3206
rect 322 3179 328 3180
rect 322 3175 323 3179
rect 327 3175 328 3179
rect 322 3174 328 3175
rect 516 3139 518 3216
rect 564 3212 566 3358
rect 596 3320 598 3381
rect 682 3359 688 3360
rect 682 3355 683 3359
rect 687 3355 688 3359
rect 682 3354 688 3355
rect 684 3336 686 3354
rect 682 3335 688 3336
rect 682 3331 683 3335
rect 687 3331 688 3335
rect 682 3330 688 3331
rect 732 3320 734 3381
rect 820 3360 822 3446
rect 900 3420 902 3574
rect 924 3572 926 3633
rect 1050 3615 1056 3616
rect 1010 3611 1016 3612
rect 1010 3607 1011 3611
rect 1015 3607 1016 3611
rect 1050 3611 1051 3615
rect 1055 3611 1056 3615
rect 1050 3610 1056 3611
rect 1010 3606 1016 3607
rect 922 3571 928 3572
rect 922 3567 923 3571
rect 927 3567 928 3571
rect 922 3566 928 3567
rect 950 3556 956 3557
rect 950 3552 951 3556
rect 955 3552 956 3556
rect 950 3551 956 3552
rect 952 3507 954 3551
rect 951 3506 955 3507
rect 951 3501 955 3502
rect 975 3506 979 3507
rect 975 3501 979 3502
rect 976 3477 978 3501
rect 974 3476 980 3477
rect 974 3472 975 3476
rect 979 3472 980 3476
rect 974 3471 980 3472
rect 946 3461 952 3462
rect 946 3457 947 3461
rect 951 3457 952 3461
rect 946 3456 952 3457
rect 898 3419 904 3420
rect 898 3415 899 3419
rect 903 3415 904 3419
rect 898 3414 904 3415
rect 948 3387 950 3456
rect 1012 3452 1014 3606
rect 1052 3580 1054 3610
rect 1050 3579 1056 3580
rect 1050 3575 1051 3579
rect 1055 3575 1056 3579
rect 1050 3574 1056 3575
rect 1068 3572 1070 3633
rect 1194 3615 1200 3616
rect 1194 3611 1195 3615
rect 1199 3611 1200 3615
rect 1194 3610 1200 3611
rect 1196 3580 1198 3610
rect 1204 3580 1206 3674
rect 1316 3639 1318 3716
rect 1934 3715 1940 3716
rect 1330 3711 1336 3712
rect 1330 3707 1331 3711
rect 1335 3707 1336 3711
rect 1330 3706 1336 3707
rect 1332 3680 1334 3706
rect 1330 3679 1336 3680
rect 1330 3675 1331 3679
rect 1335 3675 1336 3679
rect 1330 3674 1336 3675
rect 1936 3639 1938 3715
rect 1976 3703 1978 3771
rect 1996 3703 1998 3772
rect 2084 3736 2086 3870
rect 2404 3868 2406 3929
rect 2522 3911 2528 3912
rect 2522 3907 2523 3911
rect 2527 3907 2528 3911
rect 2522 3906 2528 3907
rect 2530 3911 2536 3912
rect 2530 3907 2531 3911
rect 2535 3907 2536 3911
rect 2530 3906 2536 3907
rect 2402 3867 2408 3868
rect 2402 3863 2403 3867
rect 2407 3863 2408 3867
rect 2402 3862 2408 3863
rect 2430 3852 2436 3853
rect 2430 3848 2431 3852
rect 2435 3848 2436 3852
rect 2430 3847 2436 3848
rect 2432 3823 2434 3847
rect 2524 3836 2526 3906
rect 2532 3876 2534 3906
rect 2530 3875 2536 3876
rect 2530 3871 2531 3875
rect 2535 3871 2536 3875
rect 2530 3870 2536 3871
rect 2828 3868 2830 3929
rect 2954 3911 2960 3912
rect 2954 3907 2955 3911
rect 2959 3907 2960 3911
rect 2954 3906 2960 3907
rect 2956 3876 2958 3906
rect 2954 3875 2960 3876
rect 2954 3871 2955 3875
rect 2959 3871 2960 3875
rect 2954 3870 2960 3871
rect 3252 3868 3254 3929
rect 3378 3911 3384 3912
rect 3378 3907 3379 3911
rect 3383 3907 3384 3911
rect 3378 3906 3384 3907
rect 3380 3876 3382 3906
rect 3378 3875 3384 3876
rect 3378 3871 3379 3875
rect 3383 3871 3384 3875
rect 3378 3870 3384 3871
rect 3652 3868 3654 3929
rect 3780 3876 3782 3934
rect 3799 3929 3803 3930
rect 3778 3875 3784 3876
rect 3778 3871 3779 3875
rect 3783 3871 3784 3875
rect 3778 3870 3784 3871
rect 3800 3869 3802 3929
rect 3840 3897 3842 3957
rect 3838 3896 3844 3897
rect 3860 3896 3862 3957
rect 3986 3939 3992 3940
rect 3986 3935 3987 3939
rect 3991 3935 3992 3939
rect 3986 3934 3992 3935
rect 3988 3904 3990 3934
rect 3986 3903 3992 3904
rect 3986 3899 3987 3903
rect 3991 3899 3992 3903
rect 3986 3898 3992 3899
rect 3996 3896 3998 3957
rect 4124 3904 4126 3982
rect 4132 3963 4134 4024
rect 4268 3963 4270 4024
rect 4284 3988 4286 4146
rect 4380 4144 4382 4205
rect 4516 4144 4518 4205
rect 4523 4180 4527 4181
rect 4523 4175 4527 4176
rect 4524 4152 4526 4175
rect 4522 4151 4528 4152
rect 4522 4147 4523 4151
rect 4527 4147 4528 4151
rect 4522 4146 4528 4147
rect 5664 4145 5666 4205
rect 5662 4144 5668 4145
rect 4378 4143 4384 4144
rect 4378 4139 4379 4143
rect 4383 4139 4384 4143
rect 4378 4138 4384 4139
rect 4514 4143 4520 4144
rect 4514 4139 4515 4143
rect 4519 4139 4520 4143
rect 5662 4140 5663 4144
rect 5667 4140 5668 4144
rect 5662 4139 5668 4140
rect 4514 4138 4520 4139
rect 4406 4128 4412 4129
rect 4406 4124 4407 4128
rect 4411 4124 4412 4128
rect 4406 4123 4412 4124
rect 4542 4128 4548 4129
rect 4542 4124 4543 4128
rect 4547 4124 4548 4128
rect 4542 4123 4548 4124
rect 5662 4127 5668 4128
rect 5662 4123 5663 4127
rect 5667 4123 5668 4127
rect 4408 4075 4410 4123
rect 4544 4075 4546 4123
rect 5662 4122 5668 4123
rect 5664 4075 5666 4122
rect 4295 4074 4299 4075
rect 4295 4069 4299 4070
rect 4407 4074 4411 4075
rect 4407 4069 4411 4070
rect 4431 4074 4435 4075
rect 4431 4069 4435 4070
rect 4543 4074 4547 4075
rect 4543 4069 4547 4070
rect 4567 4074 4571 4075
rect 4567 4069 4571 4070
rect 4703 4074 4707 4075
rect 4703 4069 4707 4070
rect 4839 4074 4843 4075
rect 4839 4069 4843 4070
rect 5663 4074 5667 4075
rect 5663 4069 5667 4070
rect 4296 4045 4298 4069
rect 4432 4045 4434 4069
rect 4568 4045 4570 4069
rect 4704 4045 4706 4069
rect 4840 4045 4842 4069
rect 5664 4046 5666 4069
rect 5662 4045 5668 4046
rect 4294 4044 4300 4045
rect 4294 4040 4295 4044
rect 4299 4040 4300 4044
rect 4294 4039 4300 4040
rect 4430 4044 4436 4045
rect 4430 4040 4431 4044
rect 4435 4040 4436 4044
rect 4430 4039 4436 4040
rect 4566 4044 4572 4045
rect 4566 4040 4567 4044
rect 4571 4040 4572 4044
rect 4566 4039 4572 4040
rect 4702 4044 4708 4045
rect 4702 4040 4703 4044
rect 4707 4040 4708 4044
rect 4702 4039 4708 4040
rect 4838 4044 4844 4045
rect 4838 4040 4839 4044
rect 4843 4040 4844 4044
rect 5662 4041 5663 4045
rect 5667 4041 5668 4045
rect 5662 4040 5668 4041
rect 4838 4039 4844 4040
rect 4402 4029 4408 4030
rect 4402 4025 4403 4029
rect 4407 4025 4408 4029
rect 4402 4024 4408 4025
rect 4538 4029 4544 4030
rect 4538 4025 4539 4029
rect 4543 4025 4544 4029
rect 4538 4024 4544 4025
rect 4674 4029 4680 4030
rect 4674 4025 4675 4029
rect 4679 4025 4680 4029
rect 4674 4024 4680 4025
rect 4810 4029 4816 4030
rect 4810 4025 4811 4029
rect 4815 4025 4816 4029
rect 4810 4024 4816 4025
rect 5662 4028 5668 4029
rect 5662 4024 5663 4028
rect 5667 4024 5668 4028
rect 4282 3987 4288 3988
rect 4282 3983 4283 3987
rect 4287 3983 4288 3987
rect 4282 3982 4288 3983
rect 4404 3963 4406 4024
rect 4418 4019 4424 4020
rect 4418 4015 4419 4019
rect 4423 4015 4424 4019
rect 4418 4014 4424 4015
rect 4420 3988 4422 4014
rect 4418 3987 4424 3988
rect 4418 3983 4419 3987
rect 4423 3983 4424 3987
rect 4418 3982 4424 3983
rect 4540 3963 4542 4024
rect 4554 4019 4560 4020
rect 4554 4015 4555 4019
rect 4559 4015 4560 4019
rect 4554 4014 4560 4015
rect 4556 3988 4558 4014
rect 4554 3987 4560 3988
rect 4554 3983 4555 3987
rect 4559 3983 4560 3987
rect 4554 3982 4560 3983
rect 4676 3963 4678 4024
rect 4690 4019 4696 4020
rect 4690 4015 4691 4019
rect 4695 4015 4696 4019
rect 4690 4014 4696 4015
rect 4692 3988 4694 4014
rect 4690 3987 4696 3988
rect 4690 3983 4691 3987
rect 4695 3983 4696 3987
rect 4690 3982 4696 3983
rect 4812 3963 4814 4024
rect 5662 4023 5668 4024
rect 4826 4019 4832 4020
rect 4826 4015 4827 4019
rect 4831 4015 4832 4019
rect 4826 4014 4832 4015
rect 4828 3988 4830 4014
rect 4826 3987 4832 3988
rect 4826 3983 4827 3987
rect 4831 3983 4832 3987
rect 4826 3982 4832 3983
rect 5664 3963 5666 4023
rect 4131 3962 4135 3963
rect 4131 3957 4135 3958
rect 4147 3962 4151 3963
rect 4147 3957 4151 3958
rect 4267 3962 4271 3963
rect 4267 3957 4271 3958
rect 4299 3962 4303 3963
rect 4299 3957 4303 3958
rect 4403 3962 4407 3963
rect 4403 3957 4407 3958
rect 4459 3962 4463 3963
rect 4459 3957 4463 3958
rect 4539 3962 4543 3963
rect 4539 3957 4543 3958
rect 4619 3962 4623 3963
rect 4619 3957 4623 3958
rect 4675 3962 4679 3963
rect 4675 3957 4679 3958
rect 4779 3962 4783 3963
rect 4779 3957 4783 3958
rect 4811 3962 4815 3963
rect 4811 3957 4815 3958
rect 5663 3962 5667 3963
rect 5663 3957 5667 3958
rect 4122 3903 4128 3904
rect 4122 3899 4123 3903
rect 4127 3899 4128 3903
rect 4122 3898 4128 3899
rect 4148 3896 4150 3957
rect 4274 3939 4280 3940
rect 4274 3935 4275 3939
rect 4279 3935 4280 3939
rect 4274 3934 4280 3935
rect 4276 3904 4278 3934
rect 4274 3903 4280 3904
rect 4274 3899 4275 3903
rect 4279 3899 4280 3903
rect 4274 3898 4280 3899
rect 4300 3896 4302 3957
rect 4450 3939 4456 3940
rect 4450 3935 4451 3939
rect 4455 3935 4456 3939
rect 4450 3934 4456 3935
rect 4452 3904 4454 3934
rect 4450 3903 4456 3904
rect 4450 3899 4451 3903
rect 4455 3899 4456 3903
rect 4450 3898 4456 3899
rect 4460 3896 4462 3957
rect 4610 3939 4616 3940
rect 4610 3935 4611 3939
rect 4615 3935 4616 3939
rect 4610 3934 4616 3935
rect 4612 3904 4614 3934
rect 4610 3903 4616 3904
rect 4610 3899 4611 3903
rect 4615 3899 4616 3903
rect 4610 3898 4616 3899
rect 4620 3896 4622 3957
rect 4770 3939 4776 3940
rect 4770 3935 4771 3939
rect 4775 3935 4776 3939
rect 4770 3934 4776 3935
rect 4772 3904 4774 3934
rect 4770 3903 4776 3904
rect 4770 3899 4771 3903
rect 4775 3899 4776 3903
rect 4770 3898 4776 3899
rect 4780 3896 4782 3957
rect 4786 3903 4792 3904
rect 4786 3899 4787 3903
rect 4791 3899 4792 3903
rect 4786 3898 4792 3899
rect 3838 3892 3839 3896
rect 3843 3892 3844 3896
rect 3838 3891 3844 3892
rect 3858 3895 3864 3896
rect 3858 3891 3859 3895
rect 3863 3891 3864 3895
rect 3858 3890 3864 3891
rect 3994 3895 4000 3896
rect 3994 3891 3995 3895
rect 3999 3891 4000 3895
rect 3994 3890 4000 3891
rect 4146 3895 4152 3896
rect 4146 3891 4147 3895
rect 4151 3891 4152 3895
rect 4146 3890 4152 3891
rect 4298 3895 4304 3896
rect 4298 3891 4299 3895
rect 4303 3891 4304 3895
rect 4298 3890 4304 3891
rect 4458 3895 4464 3896
rect 4458 3891 4459 3895
rect 4463 3891 4464 3895
rect 4458 3890 4464 3891
rect 4618 3895 4624 3896
rect 4618 3891 4619 3895
rect 4623 3891 4624 3895
rect 4618 3890 4624 3891
rect 4778 3895 4784 3896
rect 4778 3891 4779 3895
rect 4783 3891 4784 3895
rect 4778 3890 4784 3891
rect 3886 3880 3892 3881
rect 3838 3879 3844 3880
rect 3838 3875 3839 3879
rect 3843 3875 3844 3879
rect 3886 3876 3887 3880
rect 3891 3876 3892 3880
rect 3886 3875 3892 3876
rect 4022 3880 4028 3881
rect 4022 3876 4023 3880
rect 4027 3876 4028 3880
rect 4022 3875 4028 3876
rect 4174 3880 4180 3881
rect 4174 3876 4175 3880
rect 4179 3876 4180 3880
rect 4174 3875 4180 3876
rect 4326 3880 4332 3881
rect 4326 3876 4327 3880
rect 4331 3876 4332 3880
rect 4326 3875 4332 3876
rect 4486 3880 4492 3881
rect 4486 3876 4487 3880
rect 4491 3876 4492 3880
rect 4486 3875 4492 3876
rect 4646 3880 4652 3881
rect 4646 3876 4647 3880
rect 4651 3876 4652 3880
rect 4646 3875 4652 3876
rect 3838 3874 3844 3875
rect 3798 3868 3804 3869
rect 2826 3867 2832 3868
rect 2826 3863 2827 3867
rect 2831 3863 2832 3867
rect 2826 3862 2832 3863
rect 3250 3867 3256 3868
rect 3250 3863 3251 3867
rect 3255 3863 3256 3867
rect 3250 3862 3256 3863
rect 3650 3867 3656 3868
rect 3650 3863 3651 3867
rect 3655 3863 3656 3867
rect 3798 3864 3799 3868
rect 3803 3864 3804 3868
rect 3798 3863 3804 3864
rect 3650 3862 3656 3863
rect 2854 3852 2860 3853
rect 2854 3848 2855 3852
rect 2859 3848 2860 3852
rect 2854 3847 2860 3848
rect 3278 3852 3284 3853
rect 3278 3848 3279 3852
rect 3283 3848 3284 3852
rect 3278 3847 3284 3848
rect 3678 3852 3684 3853
rect 3678 3848 3679 3852
rect 3683 3848 3684 3852
rect 3678 3847 3684 3848
rect 3798 3851 3804 3852
rect 3798 3847 3799 3851
rect 3803 3847 3804 3851
rect 2522 3835 2528 3836
rect 2522 3831 2523 3835
rect 2527 3831 2528 3835
rect 2522 3830 2528 3831
rect 2856 3823 2858 3847
rect 3280 3823 3282 3847
rect 3654 3835 3660 3836
rect 3654 3831 3655 3835
rect 3659 3831 3660 3835
rect 3654 3830 3660 3831
rect 2175 3822 2179 3823
rect 2175 3817 2179 3818
rect 2351 3822 2355 3823
rect 2351 3817 2355 3818
rect 2431 3822 2435 3823
rect 2431 3817 2435 3818
rect 2535 3822 2539 3823
rect 2535 3817 2539 3818
rect 2719 3822 2723 3823
rect 2719 3817 2723 3818
rect 2855 3822 2859 3823
rect 2855 3817 2859 3818
rect 2895 3822 2899 3823
rect 2895 3817 2899 3818
rect 3071 3822 3075 3823
rect 3071 3817 3075 3818
rect 3247 3822 3251 3823
rect 3247 3817 3251 3818
rect 3279 3822 3283 3823
rect 3279 3817 3283 3818
rect 3423 3822 3427 3823
rect 3423 3817 3427 3818
rect 3607 3822 3611 3823
rect 3607 3817 3611 3818
rect 2176 3793 2178 3817
rect 2352 3793 2354 3817
rect 2536 3793 2538 3817
rect 2720 3793 2722 3817
rect 2896 3793 2898 3817
rect 3072 3793 3074 3817
rect 3248 3793 3250 3817
rect 3424 3793 3426 3817
rect 3608 3793 3610 3817
rect 2174 3792 2180 3793
rect 2174 3788 2175 3792
rect 2179 3788 2180 3792
rect 2174 3787 2180 3788
rect 2350 3792 2356 3793
rect 2350 3788 2351 3792
rect 2355 3788 2356 3792
rect 2350 3787 2356 3788
rect 2534 3792 2540 3793
rect 2534 3788 2535 3792
rect 2539 3788 2540 3792
rect 2534 3787 2540 3788
rect 2718 3792 2724 3793
rect 2718 3788 2719 3792
rect 2723 3788 2724 3792
rect 2718 3787 2724 3788
rect 2894 3792 2900 3793
rect 2894 3788 2895 3792
rect 2899 3788 2900 3792
rect 2894 3787 2900 3788
rect 3070 3792 3076 3793
rect 3070 3788 3071 3792
rect 3075 3788 3076 3792
rect 3070 3787 3076 3788
rect 3246 3792 3252 3793
rect 3246 3788 3247 3792
rect 3251 3788 3252 3792
rect 3246 3787 3252 3788
rect 3422 3792 3428 3793
rect 3422 3788 3423 3792
rect 3427 3788 3428 3792
rect 3422 3787 3428 3788
rect 3606 3792 3612 3793
rect 3606 3788 3607 3792
rect 3611 3788 3612 3792
rect 3606 3787 3612 3788
rect 2146 3777 2152 3778
rect 2146 3773 2147 3777
rect 2151 3773 2152 3777
rect 2146 3772 2152 3773
rect 2322 3777 2328 3778
rect 2322 3773 2323 3777
rect 2327 3773 2328 3777
rect 2322 3772 2328 3773
rect 2506 3777 2512 3778
rect 2506 3773 2507 3777
rect 2511 3773 2512 3777
rect 2506 3772 2512 3773
rect 2690 3777 2696 3778
rect 2690 3773 2691 3777
rect 2695 3773 2696 3777
rect 2690 3772 2696 3773
rect 2866 3777 2872 3778
rect 2866 3773 2867 3777
rect 2871 3773 2872 3777
rect 2866 3772 2872 3773
rect 3042 3777 3048 3778
rect 3042 3773 3043 3777
rect 3047 3773 3048 3777
rect 3042 3772 3048 3773
rect 3218 3777 3224 3778
rect 3218 3773 3219 3777
rect 3223 3773 3224 3777
rect 3218 3772 3224 3773
rect 3394 3777 3400 3778
rect 3394 3773 3395 3777
rect 3399 3773 3400 3777
rect 3394 3772 3400 3773
rect 3578 3777 3584 3778
rect 3578 3773 3579 3777
rect 3583 3773 3584 3777
rect 3578 3772 3584 3773
rect 2082 3735 2088 3736
rect 2082 3731 2083 3735
rect 2087 3731 2088 3735
rect 2082 3730 2088 3731
rect 2148 3703 2150 3772
rect 2162 3767 2168 3768
rect 2162 3763 2163 3767
rect 2167 3763 2168 3767
rect 2162 3762 2168 3763
rect 2164 3736 2166 3762
rect 2162 3735 2168 3736
rect 2162 3731 2163 3735
rect 2167 3731 2168 3735
rect 2162 3730 2168 3731
rect 2324 3703 2326 3772
rect 2338 3767 2344 3768
rect 2338 3763 2339 3767
rect 2343 3763 2344 3767
rect 2338 3762 2344 3763
rect 2340 3736 2342 3762
rect 2338 3735 2344 3736
rect 2338 3731 2339 3735
rect 2343 3731 2344 3735
rect 2338 3730 2344 3731
rect 2508 3703 2510 3772
rect 2522 3767 2528 3768
rect 2522 3763 2523 3767
rect 2527 3763 2528 3767
rect 2522 3762 2528 3763
rect 2524 3736 2526 3762
rect 2522 3735 2528 3736
rect 2522 3731 2523 3735
rect 2527 3731 2528 3735
rect 2522 3730 2528 3731
rect 2692 3703 2694 3772
rect 2706 3767 2712 3768
rect 2706 3763 2707 3767
rect 2711 3763 2712 3767
rect 2706 3762 2712 3763
rect 2708 3736 2710 3762
rect 2706 3735 2712 3736
rect 2706 3731 2707 3735
rect 2711 3731 2712 3735
rect 2706 3730 2712 3731
rect 2868 3703 2870 3772
rect 3044 3703 3046 3772
rect 3058 3767 3064 3768
rect 3058 3763 3059 3767
rect 3063 3763 3064 3767
rect 3058 3762 3064 3763
rect 3060 3736 3062 3762
rect 3058 3735 3064 3736
rect 3058 3731 3059 3735
rect 3063 3731 3064 3735
rect 3058 3730 3064 3731
rect 3220 3703 3222 3772
rect 3234 3767 3240 3768
rect 3234 3763 3235 3767
rect 3239 3763 3240 3767
rect 3234 3762 3240 3763
rect 3236 3736 3238 3762
rect 3234 3735 3240 3736
rect 3234 3731 3235 3735
rect 3239 3731 3240 3735
rect 3234 3730 3240 3731
rect 3396 3703 3398 3772
rect 3410 3767 3416 3768
rect 3410 3763 3411 3767
rect 3415 3763 3416 3767
rect 3410 3762 3416 3763
rect 3412 3736 3414 3762
rect 3410 3735 3416 3736
rect 3410 3731 3411 3735
rect 3415 3731 3416 3735
rect 3410 3730 3416 3731
rect 3422 3719 3428 3720
rect 3422 3715 3423 3719
rect 3427 3715 3428 3719
rect 3422 3714 3428 3715
rect 1975 3702 1979 3703
rect 1975 3697 1979 3698
rect 1995 3702 1999 3703
rect 1995 3697 1999 3698
rect 2011 3702 2015 3703
rect 2011 3697 2015 3698
rect 2147 3702 2151 3703
rect 2147 3697 2151 3698
rect 2291 3702 2295 3703
rect 2291 3697 2295 3698
rect 2323 3702 2327 3703
rect 2323 3697 2327 3698
rect 2435 3702 2439 3703
rect 2435 3697 2439 3698
rect 2507 3702 2511 3703
rect 2507 3697 2511 3698
rect 2579 3702 2583 3703
rect 2579 3697 2583 3698
rect 2691 3702 2695 3703
rect 2691 3697 2695 3698
rect 2723 3702 2727 3703
rect 2723 3697 2727 3698
rect 2867 3702 2871 3703
rect 2867 3697 2871 3698
rect 3011 3702 3015 3703
rect 3011 3697 3015 3698
rect 3043 3702 3047 3703
rect 3043 3697 3047 3698
rect 3155 3702 3159 3703
rect 3155 3697 3159 3698
rect 3219 3702 3223 3703
rect 3219 3697 3223 3698
rect 3299 3702 3303 3703
rect 3299 3697 3303 3698
rect 3395 3702 3399 3703
rect 3395 3697 3399 3698
rect 1211 3638 1215 3639
rect 1211 3633 1215 3634
rect 1315 3638 1319 3639
rect 1315 3633 1319 3634
rect 1935 3638 1939 3639
rect 1976 3637 1978 3697
rect 1935 3633 1939 3634
rect 1974 3636 1980 3637
rect 2012 3636 2014 3697
rect 2148 3636 2150 3697
rect 2274 3679 2280 3680
rect 2274 3675 2275 3679
rect 2279 3675 2280 3679
rect 2274 3674 2280 3675
rect 2276 3644 2278 3674
rect 2274 3643 2280 3644
rect 2274 3639 2275 3643
rect 2279 3639 2280 3643
rect 2274 3638 2280 3639
rect 2292 3636 2294 3697
rect 2418 3679 2424 3680
rect 2418 3675 2419 3679
rect 2423 3675 2424 3679
rect 2418 3674 2424 3675
rect 2420 3644 2422 3674
rect 2418 3643 2424 3644
rect 2418 3639 2419 3643
rect 2423 3639 2424 3643
rect 2418 3638 2424 3639
rect 2436 3636 2438 3697
rect 2562 3679 2568 3680
rect 2562 3675 2563 3679
rect 2567 3675 2568 3679
rect 2562 3674 2568 3675
rect 2564 3644 2566 3674
rect 2562 3643 2568 3644
rect 2562 3639 2563 3643
rect 2567 3639 2568 3643
rect 2562 3638 2568 3639
rect 2580 3636 2582 3697
rect 2598 3643 2604 3644
rect 2598 3639 2599 3643
rect 2603 3639 2604 3643
rect 2598 3638 2604 3639
rect 1194 3579 1200 3580
rect 1194 3575 1195 3579
rect 1199 3575 1200 3579
rect 1194 3574 1200 3575
rect 1202 3579 1208 3580
rect 1202 3575 1203 3579
rect 1207 3575 1208 3579
rect 1202 3574 1208 3575
rect 1212 3572 1214 3633
rect 1936 3573 1938 3633
rect 1974 3632 1975 3636
rect 1979 3632 1980 3636
rect 1974 3631 1980 3632
rect 2010 3635 2016 3636
rect 2010 3631 2011 3635
rect 2015 3631 2016 3635
rect 2010 3630 2016 3631
rect 2146 3635 2152 3636
rect 2146 3631 2147 3635
rect 2151 3631 2152 3635
rect 2146 3630 2152 3631
rect 2290 3635 2296 3636
rect 2290 3631 2291 3635
rect 2295 3631 2296 3635
rect 2290 3630 2296 3631
rect 2434 3635 2440 3636
rect 2434 3631 2435 3635
rect 2439 3631 2440 3635
rect 2434 3630 2440 3631
rect 2578 3635 2584 3636
rect 2578 3631 2579 3635
rect 2583 3631 2584 3635
rect 2578 3630 2584 3631
rect 2038 3620 2044 3621
rect 1974 3619 1980 3620
rect 1974 3615 1975 3619
rect 1979 3615 1980 3619
rect 2038 3616 2039 3620
rect 2043 3616 2044 3620
rect 2038 3615 2044 3616
rect 2174 3620 2180 3621
rect 2174 3616 2175 3620
rect 2179 3616 2180 3620
rect 2174 3615 2180 3616
rect 2318 3620 2324 3621
rect 2318 3616 2319 3620
rect 2323 3616 2324 3620
rect 2318 3615 2324 3616
rect 2462 3620 2468 3621
rect 2462 3616 2463 3620
rect 2467 3616 2468 3620
rect 2462 3615 2468 3616
rect 1974 3614 1980 3615
rect 1976 3583 1978 3614
rect 2040 3583 2042 3615
rect 2176 3583 2178 3615
rect 2320 3583 2322 3615
rect 2464 3583 2466 3615
rect 1975 3582 1979 3583
rect 1975 3577 1979 3578
rect 2039 3582 2043 3583
rect 2039 3577 2043 3578
rect 2175 3582 2179 3583
rect 2175 3577 2179 3578
rect 2239 3582 2243 3583
rect 2239 3577 2243 3578
rect 2319 3582 2323 3583
rect 2319 3577 2323 3578
rect 2375 3582 2379 3583
rect 2375 3577 2379 3578
rect 2463 3582 2467 3583
rect 2463 3577 2467 3578
rect 2511 3582 2515 3583
rect 2511 3577 2515 3578
rect 1934 3572 1940 3573
rect 1066 3571 1072 3572
rect 1066 3567 1067 3571
rect 1071 3567 1072 3571
rect 1066 3566 1072 3567
rect 1210 3571 1216 3572
rect 1210 3567 1211 3571
rect 1215 3567 1216 3571
rect 1934 3568 1935 3572
rect 1939 3568 1940 3572
rect 1934 3567 1940 3568
rect 1210 3566 1216 3567
rect 1094 3556 1100 3557
rect 1094 3552 1095 3556
rect 1099 3552 1100 3556
rect 1094 3551 1100 3552
rect 1238 3556 1244 3557
rect 1238 3552 1239 3556
rect 1243 3552 1244 3556
rect 1238 3551 1244 3552
rect 1934 3555 1940 3556
rect 1934 3551 1935 3555
rect 1939 3551 1940 3555
rect 1976 3554 1978 3577
rect 1096 3507 1098 3551
rect 1240 3507 1242 3551
rect 1934 3550 1940 3551
rect 1974 3553 1980 3554
rect 2240 3553 2242 3577
rect 2376 3553 2378 3577
rect 2512 3553 2514 3577
rect 1936 3507 1938 3550
rect 1974 3549 1975 3553
rect 1979 3549 1980 3553
rect 1974 3548 1980 3549
rect 2238 3552 2244 3553
rect 2238 3548 2239 3552
rect 2243 3548 2244 3552
rect 2238 3547 2244 3548
rect 2374 3552 2380 3553
rect 2374 3548 2375 3552
rect 2379 3548 2380 3552
rect 2374 3547 2380 3548
rect 2510 3552 2516 3553
rect 2510 3548 2511 3552
rect 2515 3548 2516 3552
rect 2510 3547 2516 3548
rect 2210 3537 2216 3538
rect 1974 3536 1980 3537
rect 1974 3532 1975 3536
rect 1979 3532 1980 3536
rect 2210 3533 2211 3537
rect 2215 3533 2216 3537
rect 2210 3532 2216 3533
rect 2346 3537 2352 3538
rect 2346 3533 2347 3537
rect 2351 3533 2352 3537
rect 2346 3532 2352 3533
rect 2482 3537 2488 3538
rect 2482 3533 2483 3537
rect 2487 3533 2488 3537
rect 2482 3532 2488 3533
rect 1974 3531 1980 3532
rect 1095 3506 1099 3507
rect 1095 3501 1099 3502
rect 1239 3506 1243 3507
rect 1239 3501 1243 3502
rect 1935 3506 1939 3507
rect 1935 3501 1939 3502
rect 1936 3478 1938 3501
rect 1934 3477 1940 3478
rect 1934 3473 1935 3477
rect 1939 3473 1940 3477
rect 1934 3472 1940 3473
rect 1976 3467 1978 3531
rect 2212 3467 2214 3532
rect 2348 3467 2350 3532
rect 2362 3527 2368 3528
rect 2362 3523 2363 3527
rect 2367 3523 2368 3527
rect 2362 3522 2368 3523
rect 2364 3496 2366 3522
rect 2362 3495 2368 3496
rect 2362 3491 2363 3495
rect 2367 3491 2368 3495
rect 2362 3490 2368 3491
rect 2484 3467 2486 3532
rect 2498 3527 2504 3528
rect 2498 3523 2499 3527
rect 2503 3523 2504 3527
rect 2498 3522 2504 3523
rect 2500 3496 2502 3522
rect 2600 3512 2602 3638
rect 2724 3636 2726 3697
rect 2850 3679 2856 3680
rect 2850 3675 2851 3679
rect 2855 3675 2856 3679
rect 2850 3674 2856 3675
rect 2852 3644 2854 3674
rect 2850 3643 2856 3644
rect 2850 3639 2851 3643
rect 2855 3639 2856 3643
rect 2850 3638 2856 3639
rect 2868 3636 2870 3697
rect 2994 3679 3000 3680
rect 2994 3675 2995 3679
rect 2999 3675 3000 3679
rect 2994 3674 3000 3675
rect 2954 3663 2960 3664
rect 2954 3659 2955 3663
rect 2959 3659 2960 3663
rect 2954 3658 2960 3659
rect 2722 3635 2728 3636
rect 2722 3631 2723 3635
rect 2727 3631 2728 3635
rect 2722 3630 2728 3631
rect 2866 3635 2872 3636
rect 2866 3631 2867 3635
rect 2871 3631 2872 3635
rect 2866 3630 2872 3631
rect 2606 3620 2612 3621
rect 2606 3616 2607 3620
rect 2611 3616 2612 3620
rect 2606 3615 2612 3616
rect 2750 3620 2756 3621
rect 2750 3616 2751 3620
rect 2755 3616 2756 3620
rect 2750 3615 2756 3616
rect 2894 3620 2900 3621
rect 2894 3616 2895 3620
rect 2899 3616 2900 3620
rect 2894 3615 2900 3616
rect 2608 3583 2610 3615
rect 2752 3583 2754 3615
rect 2896 3583 2898 3615
rect 2607 3582 2611 3583
rect 2607 3577 2611 3578
rect 2647 3582 2651 3583
rect 2647 3577 2651 3578
rect 2751 3582 2755 3583
rect 2751 3577 2755 3578
rect 2783 3582 2787 3583
rect 2783 3577 2787 3578
rect 2895 3582 2899 3583
rect 2895 3577 2899 3578
rect 2919 3582 2923 3583
rect 2919 3577 2923 3578
rect 2648 3553 2650 3577
rect 2784 3553 2786 3577
rect 2920 3553 2922 3577
rect 2646 3552 2652 3553
rect 2646 3548 2647 3552
rect 2651 3548 2652 3552
rect 2646 3547 2652 3548
rect 2782 3552 2788 3553
rect 2782 3548 2783 3552
rect 2787 3548 2788 3552
rect 2782 3547 2788 3548
rect 2918 3552 2924 3553
rect 2918 3548 2919 3552
rect 2923 3548 2924 3552
rect 2918 3547 2924 3548
rect 2618 3537 2624 3538
rect 2618 3533 2619 3537
rect 2623 3533 2624 3537
rect 2618 3532 2624 3533
rect 2754 3537 2760 3538
rect 2754 3533 2755 3537
rect 2759 3533 2760 3537
rect 2754 3532 2760 3533
rect 2890 3537 2896 3538
rect 2890 3533 2891 3537
rect 2895 3533 2896 3537
rect 2890 3532 2896 3533
rect 2598 3511 2604 3512
rect 2598 3507 2599 3511
rect 2603 3507 2604 3511
rect 2598 3506 2604 3507
rect 2498 3495 2504 3496
rect 2498 3491 2499 3495
rect 2503 3491 2504 3495
rect 2498 3490 2504 3491
rect 2620 3467 2622 3532
rect 2634 3527 2640 3528
rect 2634 3523 2635 3527
rect 2639 3523 2640 3527
rect 2634 3522 2640 3523
rect 2636 3496 2638 3522
rect 2634 3495 2640 3496
rect 2634 3491 2635 3495
rect 2639 3491 2640 3495
rect 2634 3490 2640 3491
rect 2756 3467 2758 3532
rect 2770 3527 2776 3528
rect 2770 3523 2771 3527
rect 2775 3523 2776 3527
rect 2770 3522 2776 3523
rect 2802 3527 2808 3528
rect 2802 3523 2803 3527
rect 2807 3523 2808 3527
rect 2802 3522 2808 3523
rect 2772 3496 2774 3522
rect 2770 3495 2776 3496
rect 2770 3491 2771 3495
rect 2775 3491 2776 3495
rect 2770 3490 2776 3491
rect 1975 3466 1979 3467
rect 1975 3461 1979 3462
rect 2171 3466 2175 3467
rect 2171 3461 2175 3462
rect 2211 3466 2215 3467
rect 2211 3461 2215 3462
rect 2347 3466 2351 3467
rect 2347 3461 2351 3462
rect 2483 3466 2487 3467
rect 2483 3461 2487 3462
rect 2531 3466 2535 3467
rect 2531 3461 2535 3462
rect 2619 3466 2623 3467
rect 2619 3461 2623 3462
rect 2715 3466 2719 3467
rect 2715 3461 2719 3462
rect 2755 3466 2759 3467
rect 2755 3461 2759 3462
rect 1934 3460 1940 3461
rect 1934 3456 1935 3460
rect 1939 3456 1940 3460
rect 1934 3455 1940 3456
rect 962 3451 968 3452
rect 962 3447 963 3451
rect 967 3447 968 3451
rect 962 3446 968 3447
rect 1010 3451 1016 3452
rect 1010 3447 1011 3451
rect 1015 3447 1016 3451
rect 1010 3446 1016 3447
rect 964 3420 966 3446
rect 962 3419 968 3420
rect 962 3415 963 3419
rect 967 3415 968 3419
rect 962 3414 968 3415
rect 1936 3387 1938 3455
rect 1976 3401 1978 3461
rect 1974 3400 1980 3401
rect 2172 3400 2174 3461
rect 2318 3443 2324 3444
rect 2318 3439 2319 3443
rect 2323 3439 2324 3443
rect 2318 3438 2324 3439
rect 2326 3443 2332 3444
rect 2326 3439 2327 3443
rect 2331 3439 2332 3443
rect 2326 3438 2332 3439
rect 2320 3416 2322 3438
rect 2318 3415 2324 3416
rect 2318 3411 2319 3415
rect 2323 3411 2324 3415
rect 2318 3410 2324 3411
rect 2328 3408 2330 3438
rect 2326 3407 2332 3408
rect 2326 3403 2327 3407
rect 2331 3403 2332 3407
rect 2326 3402 2332 3403
rect 2348 3400 2350 3461
rect 2474 3443 2480 3444
rect 2474 3439 2475 3443
rect 2479 3439 2480 3443
rect 2474 3438 2480 3439
rect 2476 3408 2478 3438
rect 2474 3407 2480 3408
rect 2474 3403 2475 3407
rect 2479 3403 2480 3407
rect 2474 3402 2480 3403
rect 2532 3400 2534 3461
rect 2716 3400 2718 3461
rect 2804 3440 2806 3522
rect 2892 3467 2894 3532
rect 2956 3528 2958 3658
rect 2996 3644 2998 3674
rect 2994 3643 3000 3644
rect 2994 3639 2995 3643
rect 2999 3639 3000 3643
rect 2994 3638 3000 3639
rect 3012 3636 3014 3697
rect 3156 3636 3158 3697
rect 3282 3679 3288 3680
rect 3282 3675 3283 3679
rect 3287 3675 3288 3679
rect 3282 3674 3288 3675
rect 3284 3644 3286 3674
rect 3282 3643 3288 3644
rect 3282 3639 3283 3643
rect 3287 3639 3288 3643
rect 3282 3638 3288 3639
rect 3300 3636 3302 3697
rect 3424 3644 3426 3714
rect 3580 3703 3582 3772
rect 3656 3768 3658 3830
rect 3680 3823 3682 3847
rect 3798 3846 3804 3847
rect 3800 3823 3802 3846
rect 3840 3823 3842 3874
rect 3888 3823 3890 3875
rect 4024 3823 4026 3875
rect 4176 3823 4178 3875
rect 4328 3823 4330 3875
rect 4488 3823 4490 3875
rect 4648 3823 4650 3875
rect 3679 3822 3683 3823
rect 3679 3817 3683 3818
rect 3799 3822 3803 3823
rect 3799 3817 3803 3818
rect 3839 3822 3843 3823
rect 3839 3817 3843 3818
rect 3887 3822 3891 3823
rect 3887 3817 3891 3818
rect 4023 3822 4027 3823
rect 4023 3817 4027 3818
rect 4175 3822 4179 3823
rect 4175 3817 4179 3818
rect 4327 3822 4331 3823
rect 4327 3817 4331 3818
rect 4487 3822 4491 3823
rect 4487 3817 4491 3818
rect 4503 3822 4507 3823
rect 4503 3817 4507 3818
rect 4639 3822 4643 3823
rect 4639 3817 4643 3818
rect 4647 3822 4651 3823
rect 4647 3817 4651 3818
rect 4775 3822 4779 3823
rect 4775 3817 4779 3818
rect 3800 3794 3802 3817
rect 3840 3794 3842 3817
rect 3798 3793 3804 3794
rect 3798 3789 3799 3793
rect 3803 3789 3804 3793
rect 3798 3788 3804 3789
rect 3838 3793 3844 3794
rect 4504 3793 4506 3817
rect 4640 3793 4642 3817
rect 4776 3793 4778 3817
rect 3838 3789 3839 3793
rect 3843 3789 3844 3793
rect 3838 3788 3844 3789
rect 4502 3792 4508 3793
rect 4502 3788 4503 3792
rect 4507 3788 4508 3792
rect 4502 3787 4508 3788
rect 4638 3792 4644 3793
rect 4638 3788 4639 3792
rect 4643 3788 4644 3792
rect 4638 3787 4644 3788
rect 4774 3792 4780 3793
rect 4774 3788 4775 3792
rect 4779 3788 4780 3792
rect 4774 3787 4780 3788
rect 4474 3777 4480 3778
rect 3798 3776 3804 3777
rect 3798 3772 3799 3776
rect 3803 3772 3804 3776
rect 3798 3771 3804 3772
rect 3838 3776 3844 3777
rect 3838 3772 3839 3776
rect 3843 3772 3844 3776
rect 4474 3773 4475 3777
rect 4479 3773 4480 3777
rect 4474 3772 4480 3773
rect 4610 3777 4616 3778
rect 4610 3773 4611 3777
rect 4615 3773 4616 3777
rect 4610 3772 4616 3773
rect 4746 3777 4752 3778
rect 4746 3773 4747 3777
rect 4751 3773 4752 3777
rect 4746 3772 4752 3773
rect 3838 3771 3844 3772
rect 3594 3767 3600 3768
rect 3594 3763 3595 3767
rect 3599 3763 3600 3767
rect 3594 3762 3600 3763
rect 3654 3767 3660 3768
rect 3654 3763 3655 3767
rect 3659 3763 3660 3767
rect 3654 3762 3660 3763
rect 3596 3736 3598 3762
rect 3594 3735 3600 3736
rect 3594 3731 3595 3735
rect 3599 3731 3600 3735
rect 3594 3730 3600 3731
rect 3800 3703 3802 3771
rect 3579 3702 3583 3703
rect 3579 3697 3583 3698
rect 3799 3702 3803 3703
rect 3799 3697 3803 3698
rect 3422 3643 3428 3644
rect 3422 3639 3423 3643
rect 3427 3639 3428 3643
rect 3422 3638 3428 3639
rect 3800 3637 3802 3697
rect 3840 3691 3842 3771
rect 4122 3759 4128 3760
rect 4122 3755 4123 3759
rect 4127 3755 4128 3759
rect 4122 3754 4128 3755
rect 3839 3690 3843 3691
rect 3839 3685 3843 3686
rect 4019 3690 4023 3691
rect 4019 3685 4023 3686
rect 3798 3636 3804 3637
rect 3010 3635 3016 3636
rect 3010 3631 3011 3635
rect 3015 3631 3016 3635
rect 3010 3630 3016 3631
rect 3154 3635 3160 3636
rect 3154 3631 3155 3635
rect 3159 3631 3160 3635
rect 3154 3630 3160 3631
rect 3298 3635 3304 3636
rect 3298 3631 3299 3635
rect 3303 3631 3304 3635
rect 3798 3632 3799 3636
rect 3803 3632 3804 3636
rect 3798 3631 3804 3632
rect 3298 3630 3304 3631
rect 3840 3625 3842 3685
rect 3838 3624 3844 3625
rect 4020 3624 4022 3685
rect 4124 3668 4126 3754
rect 4476 3691 4478 3772
rect 4612 3691 4614 3772
rect 4626 3767 4632 3768
rect 4626 3763 4627 3767
rect 4631 3763 4632 3767
rect 4626 3762 4632 3763
rect 4628 3736 4630 3762
rect 4626 3735 4632 3736
rect 4626 3731 4627 3735
rect 4631 3731 4632 3735
rect 4626 3730 4632 3731
rect 4748 3691 4750 3772
rect 4762 3767 4768 3768
rect 4762 3763 4763 3767
rect 4767 3763 4768 3767
rect 4762 3762 4768 3763
rect 4764 3736 4766 3762
rect 4788 3752 4790 3898
rect 5664 3897 5666 3957
rect 5662 3896 5668 3897
rect 5662 3892 5663 3896
rect 5667 3892 5668 3896
rect 5662 3891 5668 3892
rect 4806 3880 4812 3881
rect 4806 3876 4807 3880
rect 4811 3876 4812 3880
rect 4806 3875 4812 3876
rect 5662 3879 5668 3880
rect 5662 3875 5663 3879
rect 5667 3875 5668 3879
rect 4808 3823 4810 3875
rect 5662 3874 5668 3875
rect 5664 3823 5666 3874
rect 4807 3822 4811 3823
rect 4807 3817 4811 3818
rect 4911 3822 4915 3823
rect 4911 3817 4915 3818
rect 5047 3822 5051 3823
rect 5047 3817 5051 3818
rect 5663 3822 5667 3823
rect 5663 3817 5667 3818
rect 4912 3793 4914 3817
rect 5048 3793 5050 3817
rect 5664 3794 5666 3817
rect 5662 3793 5668 3794
rect 4910 3792 4916 3793
rect 4910 3788 4911 3792
rect 4915 3788 4916 3792
rect 4910 3787 4916 3788
rect 5046 3792 5052 3793
rect 5046 3788 5047 3792
rect 5051 3788 5052 3792
rect 5662 3789 5663 3793
rect 5667 3789 5668 3793
rect 5662 3788 5668 3789
rect 5046 3787 5052 3788
rect 4882 3777 4888 3778
rect 4882 3773 4883 3777
rect 4887 3773 4888 3777
rect 4882 3772 4888 3773
rect 5018 3777 5024 3778
rect 5018 3773 5019 3777
rect 5023 3773 5024 3777
rect 5018 3772 5024 3773
rect 5662 3776 5668 3777
rect 5662 3772 5663 3776
rect 5667 3772 5668 3776
rect 4786 3751 4792 3752
rect 4786 3747 4787 3751
rect 4791 3747 4792 3751
rect 4786 3746 4792 3747
rect 4762 3735 4768 3736
rect 4762 3731 4763 3735
rect 4767 3731 4768 3735
rect 4762 3730 4768 3731
rect 4884 3691 4886 3772
rect 4898 3767 4904 3768
rect 4898 3763 4899 3767
rect 4903 3763 4904 3767
rect 4898 3762 4904 3763
rect 4900 3736 4902 3762
rect 4898 3735 4904 3736
rect 4898 3731 4899 3735
rect 4903 3731 4904 3735
rect 4898 3730 4904 3731
rect 5020 3691 5022 3772
rect 5662 3771 5668 3772
rect 5034 3767 5040 3768
rect 5034 3763 5035 3767
rect 5039 3763 5040 3767
rect 5034 3762 5040 3763
rect 5036 3736 5038 3762
rect 5034 3735 5040 3736
rect 5034 3731 5035 3735
rect 5039 3731 5040 3735
rect 5034 3730 5040 3731
rect 5664 3691 5666 3771
rect 4155 3690 4159 3691
rect 4155 3685 4159 3686
rect 4291 3690 4295 3691
rect 4291 3685 4295 3686
rect 4427 3690 4431 3691
rect 4427 3685 4431 3686
rect 4475 3690 4479 3691
rect 4475 3685 4479 3686
rect 4563 3690 4567 3691
rect 4563 3685 4567 3686
rect 4611 3690 4615 3691
rect 4611 3685 4615 3686
rect 4699 3690 4703 3691
rect 4699 3685 4703 3686
rect 4747 3690 4751 3691
rect 4747 3685 4751 3686
rect 4835 3690 4839 3691
rect 4835 3685 4839 3686
rect 4883 3690 4887 3691
rect 4883 3685 4887 3686
rect 4971 3690 4975 3691
rect 4971 3685 4975 3686
rect 5019 3690 5023 3691
rect 5019 3685 5023 3686
rect 5107 3690 5111 3691
rect 5107 3685 5111 3686
rect 5243 3690 5247 3691
rect 5243 3685 5247 3686
rect 5379 3690 5383 3691
rect 5379 3685 5383 3686
rect 5515 3690 5519 3691
rect 5515 3685 5519 3686
rect 5663 3690 5667 3691
rect 5663 3685 5667 3686
rect 4122 3667 4128 3668
rect 4122 3663 4123 3667
rect 4127 3663 4128 3667
rect 4122 3662 4128 3663
rect 4146 3667 4152 3668
rect 4146 3663 4147 3667
rect 4151 3663 4152 3667
rect 4146 3662 4152 3663
rect 4148 3632 4150 3662
rect 4146 3631 4152 3632
rect 4146 3627 4147 3631
rect 4151 3627 4152 3631
rect 4146 3626 4152 3627
rect 4156 3624 4158 3685
rect 4282 3667 4288 3668
rect 4282 3663 4283 3667
rect 4287 3663 4288 3667
rect 4282 3662 4288 3663
rect 4284 3632 4286 3662
rect 4282 3631 4288 3632
rect 4282 3627 4283 3631
rect 4287 3627 4288 3631
rect 4282 3626 4288 3627
rect 4292 3624 4294 3685
rect 4418 3667 4424 3668
rect 4418 3663 4419 3667
rect 4423 3663 4424 3667
rect 4418 3662 4424 3663
rect 4420 3632 4422 3662
rect 4418 3631 4424 3632
rect 4418 3627 4419 3631
rect 4423 3627 4424 3631
rect 4418 3626 4424 3627
rect 4428 3624 4430 3685
rect 4554 3667 4560 3668
rect 4554 3663 4555 3667
rect 4559 3663 4560 3667
rect 4554 3662 4560 3663
rect 4556 3632 4558 3662
rect 4554 3631 4560 3632
rect 4554 3627 4555 3631
rect 4559 3627 4560 3631
rect 4554 3626 4560 3627
rect 4564 3624 4566 3685
rect 4690 3667 4696 3668
rect 4690 3663 4691 3667
rect 4695 3663 4696 3667
rect 4690 3662 4696 3663
rect 4692 3632 4694 3662
rect 4690 3631 4696 3632
rect 4690 3627 4691 3631
rect 4695 3627 4696 3631
rect 4690 3626 4696 3627
rect 4700 3624 4702 3685
rect 4826 3667 4832 3668
rect 4826 3663 4827 3667
rect 4831 3663 4832 3667
rect 4826 3662 4832 3663
rect 4828 3632 4830 3662
rect 4826 3631 4832 3632
rect 4826 3627 4827 3631
rect 4831 3627 4832 3631
rect 4826 3626 4832 3627
rect 4836 3624 4838 3685
rect 4972 3624 4974 3685
rect 5108 3624 5110 3685
rect 5244 3624 5246 3685
rect 5380 3624 5382 3685
rect 5516 3624 5518 3685
rect 5550 3631 5556 3632
rect 5550 3627 5551 3631
rect 5555 3627 5556 3631
rect 5550 3626 5556 3627
rect 3038 3620 3044 3621
rect 3038 3616 3039 3620
rect 3043 3616 3044 3620
rect 3038 3615 3044 3616
rect 3182 3620 3188 3621
rect 3182 3616 3183 3620
rect 3187 3616 3188 3620
rect 3182 3615 3188 3616
rect 3326 3620 3332 3621
rect 3838 3620 3839 3624
rect 3843 3620 3844 3624
rect 3326 3616 3327 3620
rect 3331 3616 3332 3620
rect 3326 3615 3332 3616
rect 3798 3619 3804 3620
rect 3838 3619 3844 3620
rect 4018 3623 4024 3624
rect 4018 3619 4019 3623
rect 4023 3619 4024 3623
rect 3798 3615 3799 3619
rect 3803 3615 3804 3619
rect 4018 3618 4024 3619
rect 4154 3623 4160 3624
rect 4154 3619 4155 3623
rect 4159 3619 4160 3623
rect 4154 3618 4160 3619
rect 4290 3623 4296 3624
rect 4290 3619 4291 3623
rect 4295 3619 4296 3623
rect 4290 3618 4296 3619
rect 4426 3623 4432 3624
rect 4426 3619 4427 3623
rect 4431 3619 4432 3623
rect 4426 3618 4432 3619
rect 4562 3623 4568 3624
rect 4562 3619 4563 3623
rect 4567 3619 4568 3623
rect 4562 3618 4568 3619
rect 4698 3623 4704 3624
rect 4698 3619 4699 3623
rect 4703 3619 4704 3623
rect 4698 3618 4704 3619
rect 4834 3623 4840 3624
rect 4834 3619 4835 3623
rect 4839 3619 4840 3623
rect 4834 3618 4840 3619
rect 4970 3623 4976 3624
rect 4970 3619 4971 3623
rect 4975 3619 4976 3623
rect 4970 3618 4976 3619
rect 5106 3623 5112 3624
rect 5106 3619 5107 3623
rect 5111 3619 5112 3623
rect 5106 3618 5112 3619
rect 5242 3623 5248 3624
rect 5242 3619 5243 3623
rect 5247 3619 5248 3623
rect 5242 3618 5248 3619
rect 5378 3623 5384 3624
rect 5378 3619 5379 3623
rect 5383 3619 5384 3623
rect 5378 3618 5384 3619
rect 5514 3623 5520 3624
rect 5514 3619 5515 3623
rect 5519 3619 5520 3623
rect 5514 3618 5520 3619
rect 3040 3583 3042 3615
rect 3184 3583 3186 3615
rect 3328 3583 3330 3615
rect 3798 3614 3804 3615
rect 3800 3583 3802 3614
rect 4046 3608 4052 3609
rect 3838 3607 3844 3608
rect 3838 3603 3839 3607
rect 3843 3603 3844 3607
rect 4046 3604 4047 3608
rect 4051 3604 4052 3608
rect 4046 3603 4052 3604
rect 4182 3608 4188 3609
rect 4182 3604 4183 3608
rect 4187 3604 4188 3608
rect 4182 3603 4188 3604
rect 4318 3608 4324 3609
rect 4318 3604 4319 3608
rect 4323 3604 4324 3608
rect 4318 3603 4324 3604
rect 4454 3608 4460 3609
rect 4454 3604 4455 3608
rect 4459 3604 4460 3608
rect 4454 3603 4460 3604
rect 4590 3608 4596 3609
rect 4590 3604 4591 3608
rect 4595 3604 4596 3608
rect 4590 3603 4596 3604
rect 4726 3608 4732 3609
rect 4726 3604 4727 3608
rect 4731 3604 4732 3608
rect 4726 3603 4732 3604
rect 4862 3608 4868 3609
rect 4862 3604 4863 3608
rect 4867 3604 4868 3608
rect 4862 3603 4868 3604
rect 4998 3608 5004 3609
rect 4998 3604 4999 3608
rect 5003 3604 5004 3608
rect 4998 3603 5004 3604
rect 5134 3608 5140 3609
rect 5134 3604 5135 3608
rect 5139 3604 5140 3608
rect 5134 3603 5140 3604
rect 5270 3608 5276 3609
rect 5270 3604 5271 3608
rect 5275 3604 5276 3608
rect 5270 3603 5276 3604
rect 5406 3608 5412 3609
rect 5406 3604 5407 3608
rect 5411 3604 5412 3608
rect 5406 3603 5412 3604
rect 5542 3608 5548 3609
rect 5542 3604 5543 3608
rect 5547 3604 5548 3608
rect 5542 3603 5548 3604
rect 3838 3602 3844 3603
rect 3039 3582 3043 3583
rect 3039 3577 3043 3578
rect 3055 3582 3059 3583
rect 3055 3577 3059 3578
rect 3183 3582 3187 3583
rect 3183 3577 3187 3578
rect 3191 3582 3195 3583
rect 3191 3577 3195 3578
rect 3327 3582 3331 3583
rect 3327 3577 3331 3578
rect 3463 3582 3467 3583
rect 3463 3577 3467 3578
rect 3799 3582 3803 3583
rect 3799 3577 3803 3578
rect 3056 3553 3058 3577
rect 3192 3553 3194 3577
rect 3328 3553 3330 3577
rect 3464 3553 3466 3577
rect 3800 3554 3802 3577
rect 3798 3553 3804 3554
rect 3054 3552 3060 3553
rect 3054 3548 3055 3552
rect 3059 3548 3060 3552
rect 3054 3547 3060 3548
rect 3190 3552 3196 3553
rect 3190 3548 3191 3552
rect 3195 3548 3196 3552
rect 3190 3547 3196 3548
rect 3326 3552 3332 3553
rect 3326 3548 3327 3552
rect 3331 3548 3332 3552
rect 3326 3547 3332 3548
rect 3462 3552 3468 3553
rect 3462 3548 3463 3552
rect 3467 3548 3468 3552
rect 3798 3549 3799 3553
rect 3803 3549 3804 3553
rect 3798 3548 3804 3549
rect 3462 3547 3468 3548
rect 3026 3537 3032 3538
rect 3026 3533 3027 3537
rect 3031 3533 3032 3537
rect 3026 3532 3032 3533
rect 3162 3537 3168 3538
rect 3162 3533 3163 3537
rect 3167 3533 3168 3537
rect 3162 3532 3168 3533
rect 3298 3537 3304 3538
rect 3298 3533 3299 3537
rect 3303 3533 3304 3537
rect 3298 3532 3304 3533
rect 3434 3537 3440 3538
rect 3434 3533 3435 3537
rect 3439 3533 3440 3537
rect 3434 3532 3440 3533
rect 3798 3536 3804 3537
rect 3798 3532 3799 3536
rect 3803 3532 3804 3536
rect 2954 3527 2960 3528
rect 2954 3523 2955 3527
rect 2959 3523 2960 3527
rect 2954 3522 2960 3523
rect 3028 3467 3030 3532
rect 3164 3467 3166 3532
rect 3170 3527 3176 3528
rect 3170 3523 3171 3527
rect 3175 3523 3176 3527
rect 3170 3522 3176 3523
rect 3172 3496 3174 3522
rect 3250 3519 3256 3520
rect 3250 3515 3251 3519
rect 3255 3515 3256 3519
rect 3250 3514 3256 3515
rect 3252 3496 3254 3514
rect 3170 3495 3176 3496
rect 3170 3491 3171 3495
rect 3175 3491 3176 3495
rect 3170 3490 3176 3491
rect 3250 3495 3256 3496
rect 3250 3491 3251 3495
rect 3255 3491 3256 3495
rect 3250 3490 3256 3491
rect 3300 3467 3302 3532
rect 3386 3495 3392 3496
rect 3386 3491 3387 3495
rect 3391 3491 3392 3495
rect 3386 3490 3392 3491
rect 2891 3466 2895 3467
rect 2891 3461 2895 3462
rect 2907 3466 2911 3467
rect 2907 3461 2911 3462
rect 3027 3466 3031 3467
rect 3027 3461 3031 3462
rect 3099 3466 3103 3467
rect 3099 3461 3103 3462
rect 3163 3466 3167 3467
rect 3163 3461 3167 3462
rect 3291 3466 3295 3467
rect 3291 3461 3295 3462
rect 3299 3466 3303 3467
rect 3299 3461 3303 3462
rect 2818 3443 2824 3444
rect 2802 3439 2808 3440
rect 2802 3435 2803 3439
rect 2807 3435 2808 3439
rect 2818 3439 2819 3443
rect 2823 3439 2824 3443
rect 2818 3438 2824 3439
rect 2802 3434 2808 3435
rect 2820 3408 2822 3438
rect 2818 3407 2824 3408
rect 2818 3403 2819 3407
rect 2823 3403 2824 3407
rect 2818 3402 2824 3403
rect 2908 3400 2910 3461
rect 3030 3407 3036 3408
rect 3030 3403 3031 3407
rect 3035 3403 3036 3407
rect 3030 3402 3036 3403
rect 1974 3396 1975 3400
rect 1979 3396 1980 3400
rect 1974 3395 1980 3396
rect 2170 3399 2176 3400
rect 2170 3395 2171 3399
rect 2175 3395 2176 3399
rect 2170 3394 2176 3395
rect 2346 3399 2352 3400
rect 2346 3395 2347 3399
rect 2351 3395 2352 3399
rect 2346 3394 2352 3395
rect 2530 3399 2536 3400
rect 2530 3395 2531 3399
rect 2535 3395 2536 3399
rect 2530 3394 2536 3395
rect 2714 3399 2720 3400
rect 2714 3395 2715 3399
rect 2719 3395 2720 3399
rect 2714 3394 2720 3395
rect 2906 3399 2912 3400
rect 2906 3395 2907 3399
rect 2911 3395 2912 3399
rect 2906 3394 2912 3395
rect 867 3386 871 3387
rect 867 3381 871 3382
rect 947 3386 951 3387
rect 947 3381 951 3382
rect 1935 3386 1939 3387
rect 2198 3384 2204 3385
rect 1935 3381 1939 3382
rect 1974 3383 1980 3384
rect 818 3359 824 3360
rect 818 3355 819 3359
rect 823 3355 824 3359
rect 818 3354 824 3355
rect 738 3327 744 3328
rect 738 3323 739 3327
rect 743 3323 744 3327
rect 738 3322 744 3323
rect 594 3319 600 3320
rect 594 3315 595 3319
rect 599 3315 600 3319
rect 594 3314 600 3315
rect 730 3319 736 3320
rect 730 3315 731 3319
rect 735 3315 736 3319
rect 730 3314 736 3315
rect 622 3304 628 3305
rect 622 3300 623 3304
rect 627 3300 628 3304
rect 622 3299 628 3300
rect 624 3267 626 3299
rect 623 3266 627 3267
rect 623 3261 627 3262
rect 722 3221 728 3222
rect 722 3217 723 3221
rect 727 3217 728 3221
rect 722 3216 728 3217
rect 530 3211 536 3212
rect 530 3207 531 3211
rect 535 3207 536 3211
rect 530 3206 536 3207
rect 562 3211 568 3212
rect 562 3207 563 3211
rect 567 3207 568 3211
rect 562 3206 568 3207
rect 532 3180 534 3206
rect 530 3179 536 3180
rect 530 3175 531 3179
rect 535 3175 536 3179
rect 530 3174 536 3175
rect 724 3139 726 3216
rect 740 3180 742 3322
rect 868 3320 870 3381
rect 1936 3321 1938 3381
rect 1974 3379 1975 3383
rect 1979 3379 1980 3383
rect 2198 3380 2199 3384
rect 2203 3380 2204 3384
rect 2198 3379 2204 3380
rect 2374 3384 2380 3385
rect 2374 3380 2375 3384
rect 2379 3380 2380 3384
rect 2374 3379 2380 3380
rect 2558 3384 2564 3385
rect 2558 3380 2559 3384
rect 2563 3380 2564 3384
rect 2558 3379 2564 3380
rect 2742 3384 2748 3385
rect 2742 3380 2743 3384
rect 2747 3380 2748 3384
rect 2742 3379 2748 3380
rect 2934 3384 2940 3385
rect 2934 3380 2935 3384
rect 2939 3380 2940 3384
rect 2934 3379 2940 3380
rect 1974 3378 1980 3379
rect 1976 3331 1978 3378
rect 2200 3331 2202 3379
rect 2376 3331 2378 3379
rect 2560 3331 2562 3379
rect 2744 3331 2746 3379
rect 2936 3331 2938 3379
rect 1975 3330 1979 3331
rect 1975 3325 1979 3326
rect 2151 3330 2155 3331
rect 2151 3325 2155 3326
rect 2199 3330 2203 3331
rect 2199 3325 2203 3326
rect 2375 3330 2379 3331
rect 2375 3325 2379 3326
rect 2399 3330 2403 3331
rect 2399 3325 2403 3326
rect 2559 3330 2563 3331
rect 2559 3325 2563 3326
rect 2687 3330 2691 3331
rect 2687 3325 2691 3326
rect 2743 3330 2747 3331
rect 2743 3325 2747 3326
rect 2935 3330 2939 3331
rect 2935 3325 2939 3326
rect 3015 3330 3019 3331
rect 3015 3325 3019 3326
rect 1934 3320 1940 3321
rect 866 3319 872 3320
rect 866 3315 867 3319
rect 871 3315 872 3319
rect 1934 3316 1935 3320
rect 1939 3316 1940 3320
rect 1934 3315 1940 3316
rect 866 3314 872 3315
rect 758 3304 764 3305
rect 758 3300 759 3304
rect 763 3300 764 3304
rect 758 3299 764 3300
rect 894 3304 900 3305
rect 894 3300 895 3304
rect 899 3300 900 3304
rect 894 3299 900 3300
rect 1934 3303 1940 3304
rect 1934 3299 1935 3303
rect 1939 3299 1940 3303
rect 1976 3302 1978 3325
rect 760 3267 762 3299
rect 896 3267 898 3299
rect 1934 3298 1940 3299
rect 1974 3301 1980 3302
rect 2152 3301 2154 3325
rect 2400 3301 2402 3325
rect 2688 3301 2690 3325
rect 3016 3301 3018 3325
rect 1936 3267 1938 3298
rect 1974 3297 1975 3301
rect 1979 3297 1980 3301
rect 1974 3296 1980 3297
rect 2150 3300 2156 3301
rect 2150 3296 2151 3300
rect 2155 3296 2156 3300
rect 2150 3295 2156 3296
rect 2398 3300 2404 3301
rect 2398 3296 2399 3300
rect 2403 3296 2404 3300
rect 2398 3295 2404 3296
rect 2686 3300 2692 3301
rect 2686 3296 2687 3300
rect 2691 3296 2692 3300
rect 2686 3295 2692 3296
rect 3014 3300 3020 3301
rect 3014 3296 3015 3300
rect 3019 3296 3020 3300
rect 3014 3295 3020 3296
rect 2122 3285 2128 3286
rect 1974 3284 1980 3285
rect 1974 3280 1975 3284
rect 1979 3280 1980 3284
rect 2122 3281 2123 3285
rect 2127 3281 2128 3285
rect 2122 3280 2128 3281
rect 2370 3285 2376 3286
rect 2370 3281 2371 3285
rect 2375 3281 2376 3285
rect 2370 3280 2376 3281
rect 2658 3285 2664 3286
rect 2658 3281 2659 3285
rect 2663 3281 2664 3285
rect 2658 3280 2664 3281
rect 2986 3285 2992 3286
rect 2986 3281 2987 3285
rect 2991 3281 2992 3285
rect 2986 3280 2992 3281
rect 1974 3279 1980 3280
rect 751 3266 755 3267
rect 751 3261 755 3262
rect 759 3266 763 3267
rect 759 3261 763 3262
rect 895 3266 899 3267
rect 895 3261 899 3262
rect 959 3266 963 3267
rect 959 3261 963 3262
rect 1935 3266 1939 3267
rect 1935 3261 1939 3262
rect 752 3237 754 3261
rect 960 3237 962 3261
rect 1936 3238 1938 3261
rect 1934 3237 1940 3238
rect 750 3236 756 3237
rect 750 3232 751 3236
rect 755 3232 756 3236
rect 750 3231 756 3232
rect 958 3236 964 3237
rect 958 3232 959 3236
rect 963 3232 964 3236
rect 1934 3233 1935 3237
rect 1939 3233 1940 3237
rect 1934 3232 1940 3233
rect 958 3231 964 3232
rect 930 3221 936 3222
rect 930 3217 931 3221
rect 935 3217 936 3221
rect 930 3216 936 3217
rect 1934 3220 1940 3221
rect 1934 3216 1935 3220
rect 1939 3216 1940 3220
rect 1976 3219 1978 3279
rect 2124 3219 2126 3280
rect 2290 3243 2296 3244
rect 2290 3239 2291 3243
rect 2295 3239 2296 3243
rect 2290 3238 2296 3239
rect 738 3179 744 3180
rect 738 3175 739 3179
rect 743 3175 744 3179
rect 738 3174 744 3175
rect 932 3139 934 3216
rect 1934 3215 1940 3216
rect 1975 3218 1979 3219
rect 946 3211 952 3212
rect 946 3207 947 3211
rect 951 3207 952 3211
rect 946 3206 952 3207
rect 1058 3211 1064 3212
rect 1058 3207 1059 3211
rect 1063 3207 1064 3211
rect 1058 3206 1064 3207
rect 948 3180 950 3206
rect 946 3179 952 3180
rect 946 3175 947 3179
rect 951 3175 952 3179
rect 946 3174 952 3175
rect 307 3138 311 3139
rect 307 3133 311 3134
rect 371 3138 375 3139
rect 371 3133 375 3134
rect 515 3138 519 3139
rect 515 3133 519 3134
rect 627 3138 631 3139
rect 627 3133 631 3134
rect 723 3138 727 3139
rect 723 3133 727 3134
rect 875 3138 879 3139
rect 875 3133 879 3134
rect 931 3138 935 3139
rect 931 3133 935 3134
rect 330 3115 336 3116
rect 330 3111 331 3115
rect 335 3111 336 3115
rect 330 3110 336 3111
rect 226 3079 232 3080
rect 226 3075 227 3079
rect 231 3075 232 3079
rect 226 3074 232 3075
rect 110 3068 111 3072
rect 115 3068 116 3072
rect 110 3067 116 3068
rect 130 3071 136 3072
rect 130 3067 131 3071
rect 135 3067 136 3071
rect 130 3066 136 3067
rect 158 3056 164 3057
rect 110 3055 116 3056
rect 110 3051 111 3055
rect 115 3051 116 3055
rect 158 3052 159 3056
rect 163 3052 164 3056
rect 158 3051 164 3052
rect 110 3050 116 3051
rect 112 3027 114 3050
rect 160 3027 162 3051
rect 111 3026 115 3027
rect 111 3021 115 3022
rect 159 3026 163 3027
rect 159 3021 163 3022
rect 175 3026 179 3027
rect 175 3021 179 3022
rect 112 2998 114 3021
rect 110 2997 116 2998
rect 176 2997 178 3021
rect 110 2993 111 2997
rect 115 2993 116 2997
rect 110 2992 116 2993
rect 174 2996 180 2997
rect 174 2992 175 2996
rect 179 2992 180 2996
rect 174 2991 180 2992
rect 146 2981 152 2982
rect 110 2980 116 2981
rect 110 2976 111 2980
rect 115 2976 116 2980
rect 146 2977 147 2981
rect 151 2977 152 2981
rect 146 2976 152 2977
rect 110 2975 116 2976
rect 112 2911 114 2975
rect 148 2911 150 2976
rect 332 2972 334 3110
rect 372 3072 374 3133
rect 628 3072 630 3133
rect 822 3115 828 3116
rect 822 3111 823 3115
rect 827 3111 828 3115
rect 822 3110 828 3111
rect 824 3080 826 3110
rect 682 3079 688 3080
rect 682 3075 683 3079
rect 687 3075 688 3079
rect 682 3074 688 3075
rect 822 3079 828 3080
rect 822 3075 823 3079
rect 827 3075 828 3079
rect 822 3074 828 3075
rect 370 3071 376 3072
rect 370 3067 371 3071
rect 375 3067 376 3071
rect 370 3066 376 3067
rect 626 3071 632 3072
rect 626 3067 627 3071
rect 631 3067 632 3071
rect 626 3066 632 3067
rect 398 3056 404 3057
rect 398 3052 399 3056
rect 403 3052 404 3056
rect 398 3051 404 3052
rect 654 3056 660 3057
rect 654 3052 655 3056
rect 659 3052 660 3056
rect 654 3051 660 3052
rect 400 3027 402 3051
rect 656 3027 658 3051
rect 399 3026 403 3027
rect 399 3021 403 3022
rect 407 3026 411 3027
rect 407 3021 411 3022
rect 623 3026 627 3027
rect 623 3021 627 3022
rect 655 3026 659 3027
rect 655 3021 659 3022
rect 408 2997 410 3021
rect 624 2997 626 3021
rect 406 2996 412 2997
rect 406 2992 407 2996
rect 411 2992 412 2996
rect 406 2991 412 2992
rect 622 2996 628 2997
rect 622 2992 623 2996
rect 627 2992 628 2996
rect 622 2991 628 2992
rect 378 2981 384 2982
rect 378 2977 379 2981
rect 383 2977 384 2981
rect 378 2976 384 2977
rect 594 2981 600 2982
rect 594 2977 595 2981
rect 599 2977 600 2981
rect 594 2976 600 2977
rect 330 2971 336 2972
rect 330 2967 331 2971
rect 335 2967 336 2971
rect 330 2966 336 2967
rect 338 2971 344 2972
rect 338 2967 339 2971
rect 343 2967 344 2971
rect 338 2966 344 2967
rect 340 2940 342 2966
rect 338 2939 344 2940
rect 338 2935 339 2939
rect 343 2935 344 2939
rect 338 2934 344 2935
rect 380 2911 382 2976
rect 466 2939 472 2940
rect 466 2935 467 2939
rect 471 2935 472 2939
rect 466 2934 472 2935
rect 111 2910 115 2911
rect 111 2905 115 2906
rect 147 2910 151 2911
rect 147 2905 151 2906
rect 379 2910 383 2911
rect 379 2905 383 2906
rect 395 2910 399 2911
rect 395 2905 399 2906
rect 112 2845 114 2905
rect 110 2844 116 2845
rect 396 2844 398 2905
rect 468 2852 470 2934
rect 596 2911 598 2976
rect 684 2940 686 3074
rect 876 3072 878 3133
rect 1060 3116 1062 3206
rect 1914 3195 1920 3196
rect 1914 3191 1915 3195
rect 1919 3191 1920 3195
rect 1914 3190 1920 3191
rect 1115 3138 1119 3139
rect 1115 3133 1119 3134
rect 1347 3138 1351 3139
rect 1347 3133 1351 3134
rect 1579 3138 1583 3139
rect 1579 3133 1583 3134
rect 1787 3138 1791 3139
rect 1787 3133 1791 3134
rect 1050 3115 1056 3116
rect 1050 3111 1051 3115
rect 1055 3111 1056 3115
rect 1050 3110 1056 3111
rect 1058 3115 1064 3116
rect 1058 3111 1059 3115
rect 1063 3111 1064 3115
rect 1058 3110 1064 3111
rect 1052 3080 1054 3110
rect 1050 3079 1056 3080
rect 1050 3075 1051 3079
rect 1055 3075 1056 3079
rect 1050 3074 1056 3075
rect 1116 3072 1118 3133
rect 1348 3072 1350 3133
rect 1450 3115 1456 3116
rect 1450 3111 1451 3115
rect 1455 3111 1456 3115
rect 1450 3110 1456 3111
rect 1474 3115 1480 3116
rect 1474 3111 1475 3115
rect 1479 3111 1480 3115
rect 1474 3110 1480 3111
rect 874 3071 880 3072
rect 874 3067 875 3071
rect 879 3067 880 3071
rect 874 3066 880 3067
rect 1114 3071 1120 3072
rect 1114 3067 1115 3071
rect 1119 3067 1120 3071
rect 1114 3066 1120 3067
rect 1346 3071 1352 3072
rect 1346 3067 1347 3071
rect 1351 3067 1352 3071
rect 1346 3066 1352 3067
rect 902 3056 908 3057
rect 902 3052 903 3056
rect 907 3052 908 3056
rect 902 3051 908 3052
rect 1142 3056 1148 3057
rect 1142 3052 1143 3056
rect 1147 3052 1148 3056
rect 1142 3051 1148 3052
rect 1374 3056 1380 3057
rect 1374 3052 1375 3056
rect 1379 3052 1380 3056
rect 1374 3051 1380 3052
rect 904 3027 906 3051
rect 1144 3027 1146 3051
rect 1376 3027 1378 3051
rect 823 3026 827 3027
rect 823 3021 827 3022
rect 903 3026 907 3027
rect 903 3021 907 3022
rect 1007 3026 1011 3027
rect 1007 3021 1011 3022
rect 1143 3026 1147 3027
rect 1143 3021 1147 3022
rect 1183 3026 1187 3027
rect 1183 3021 1187 3022
rect 1351 3026 1355 3027
rect 1351 3021 1355 3022
rect 1375 3026 1379 3027
rect 1375 3021 1379 3022
rect 824 2997 826 3021
rect 1008 2997 1010 3021
rect 1184 2997 1186 3021
rect 1352 2997 1354 3021
rect 1452 3012 1454 3110
rect 1476 3080 1478 3110
rect 1474 3079 1480 3080
rect 1474 3075 1475 3079
rect 1479 3075 1480 3079
rect 1474 3074 1480 3075
rect 1580 3072 1582 3133
rect 1706 3115 1712 3116
rect 1706 3111 1707 3115
rect 1711 3111 1712 3115
rect 1706 3110 1712 3111
rect 1708 3080 1710 3110
rect 1706 3079 1712 3080
rect 1706 3075 1707 3079
rect 1711 3075 1712 3079
rect 1706 3074 1712 3075
rect 1788 3072 1790 3133
rect 1916 3080 1918 3190
rect 1936 3139 1938 3215
rect 1975 3213 1979 3214
rect 1995 3218 1999 3219
rect 1995 3213 1999 3214
rect 2123 3218 2127 3219
rect 2123 3213 2127 3214
rect 2147 3218 2151 3219
rect 2147 3213 2151 3214
rect 1976 3153 1978 3213
rect 1974 3152 1980 3153
rect 1996 3152 1998 3213
rect 2122 3195 2128 3196
rect 2122 3191 2123 3195
rect 2127 3191 2128 3195
rect 2122 3190 2128 3191
rect 2124 3160 2126 3190
rect 2122 3159 2128 3160
rect 2122 3155 2123 3159
rect 2127 3155 2128 3159
rect 2122 3154 2128 3155
rect 2148 3152 2150 3213
rect 2274 3195 2280 3196
rect 2274 3191 2275 3195
rect 2279 3191 2280 3195
rect 2274 3190 2280 3191
rect 2276 3160 2278 3190
rect 2292 3160 2294 3238
rect 2372 3219 2374 3280
rect 2386 3275 2392 3276
rect 2386 3271 2387 3275
rect 2391 3271 2392 3275
rect 2386 3270 2392 3271
rect 2388 3244 2390 3270
rect 2386 3243 2392 3244
rect 2386 3239 2387 3243
rect 2391 3239 2392 3243
rect 2386 3238 2392 3239
rect 2660 3219 2662 3280
rect 2674 3275 2680 3276
rect 2674 3271 2675 3275
rect 2679 3271 2680 3275
rect 2674 3270 2680 3271
rect 2682 3275 2688 3276
rect 2682 3271 2683 3275
rect 2687 3271 2688 3275
rect 2682 3270 2688 3271
rect 2676 3244 2678 3270
rect 2674 3243 2680 3244
rect 2674 3239 2675 3243
rect 2679 3239 2680 3243
rect 2674 3238 2680 3239
rect 2347 3218 2351 3219
rect 2347 3213 2351 3214
rect 2371 3218 2375 3219
rect 2371 3213 2375 3214
rect 2555 3218 2559 3219
rect 2555 3213 2559 3214
rect 2659 3218 2663 3219
rect 2659 3213 2663 3214
rect 2274 3159 2280 3160
rect 2274 3155 2275 3159
rect 2279 3155 2280 3159
rect 2274 3154 2280 3155
rect 2290 3159 2296 3160
rect 2290 3155 2291 3159
rect 2295 3155 2296 3159
rect 2290 3154 2296 3155
rect 2348 3152 2350 3213
rect 2556 3152 2558 3213
rect 2684 3204 2686 3270
rect 2988 3219 2990 3280
rect 3032 3244 3034 3402
rect 3100 3400 3102 3461
rect 3226 3443 3232 3444
rect 3186 3439 3192 3440
rect 3186 3435 3187 3439
rect 3191 3435 3192 3439
rect 3226 3439 3227 3443
rect 3231 3439 3232 3443
rect 3226 3438 3232 3439
rect 3186 3434 3192 3435
rect 3188 3416 3190 3434
rect 3186 3415 3192 3416
rect 3186 3411 3187 3415
rect 3191 3411 3192 3415
rect 3186 3410 3192 3411
rect 3228 3408 3230 3438
rect 3226 3407 3232 3408
rect 3226 3403 3227 3407
rect 3231 3403 3232 3407
rect 3226 3402 3232 3403
rect 3292 3400 3294 3461
rect 3388 3408 3390 3490
rect 3436 3467 3438 3532
rect 3798 3531 3804 3532
rect 3840 3531 3842 3602
rect 4048 3531 4050 3603
rect 4184 3531 4186 3603
rect 4320 3531 4322 3603
rect 4456 3531 4458 3603
rect 4592 3531 4594 3603
rect 4728 3531 4730 3603
rect 4864 3531 4866 3603
rect 5000 3531 5002 3603
rect 5136 3531 5138 3603
rect 5272 3531 5274 3603
rect 5408 3531 5410 3603
rect 5544 3531 5546 3603
rect 3450 3527 3456 3528
rect 3450 3523 3451 3527
rect 3455 3523 3456 3527
rect 3450 3522 3456 3523
rect 3452 3496 3454 3522
rect 3450 3495 3456 3496
rect 3450 3491 3451 3495
rect 3455 3491 3456 3495
rect 3450 3490 3456 3491
rect 3800 3467 3802 3531
rect 3839 3530 3843 3531
rect 3839 3525 3843 3526
rect 4047 3530 4051 3531
rect 4047 3525 4051 3526
rect 4183 3530 4187 3531
rect 4183 3525 4187 3526
rect 4319 3530 4323 3531
rect 4319 3525 4323 3526
rect 4455 3530 4459 3531
rect 4455 3525 4459 3526
rect 4591 3530 4595 3531
rect 4591 3525 4595 3526
rect 4727 3530 4731 3531
rect 4727 3525 4731 3526
rect 4863 3530 4867 3531
rect 4863 3525 4867 3526
rect 4999 3530 5003 3531
rect 4999 3525 5003 3526
rect 5135 3530 5139 3531
rect 5135 3525 5139 3526
rect 5271 3530 5275 3531
rect 5271 3525 5275 3526
rect 5407 3530 5411 3531
rect 5407 3525 5411 3526
rect 5543 3530 5547 3531
rect 5543 3525 5547 3526
rect 3840 3502 3842 3525
rect 3838 3501 3844 3502
rect 5408 3501 5410 3525
rect 5544 3501 5546 3525
rect 3838 3497 3839 3501
rect 3843 3497 3844 3501
rect 3838 3496 3844 3497
rect 5406 3500 5412 3501
rect 5406 3496 5407 3500
rect 5411 3496 5412 3500
rect 5406 3495 5412 3496
rect 5542 3500 5548 3501
rect 5542 3496 5543 3500
rect 5547 3496 5548 3500
rect 5542 3495 5548 3496
rect 5378 3485 5384 3486
rect 3838 3484 3844 3485
rect 3838 3480 3839 3484
rect 3843 3480 3844 3484
rect 5378 3481 5379 3485
rect 5383 3481 5384 3485
rect 5378 3480 5384 3481
rect 5514 3485 5520 3486
rect 5514 3481 5515 3485
rect 5519 3481 5520 3485
rect 5514 3480 5520 3481
rect 3838 3479 3844 3480
rect 3435 3466 3439 3467
rect 3435 3461 3439 3462
rect 3483 3466 3487 3467
rect 3483 3461 3487 3462
rect 3651 3466 3655 3467
rect 3651 3461 3655 3462
rect 3799 3466 3803 3467
rect 3799 3461 3803 3462
rect 3386 3407 3392 3408
rect 3386 3403 3387 3407
rect 3391 3403 3392 3407
rect 3386 3402 3392 3403
rect 3484 3400 3486 3461
rect 3638 3443 3644 3444
rect 3638 3439 3639 3443
rect 3643 3439 3644 3443
rect 3638 3438 3644 3439
rect 3640 3408 3642 3438
rect 3638 3407 3644 3408
rect 3638 3403 3639 3407
rect 3643 3403 3644 3407
rect 3638 3402 3644 3403
rect 3652 3400 3654 3461
rect 3738 3439 3744 3440
rect 3738 3435 3739 3439
rect 3743 3435 3744 3439
rect 3738 3434 3744 3435
rect 3098 3399 3104 3400
rect 3098 3395 3099 3399
rect 3103 3395 3104 3399
rect 3098 3394 3104 3395
rect 3290 3399 3296 3400
rect 3290 3395 3291 3399
rect 3295 3395 3296 3399
rect 3290 3394 3296 3395
rect 3482 3399 3488 3400
rect 3482 3395 3483 3399
rect 3487 3395 3488 3399
rect 3482 3394 3488 3395
rect 3650 3399 3656 3400
rect 3650 3395 3651 3399
rect 3655 3395 3656 3399
rect 3650 3394 3656 3395
rect 3126 3384 3132 3385
rect 3126 3380 3127 3384
rect 3131 3380 3132 3384
rect 3126 3379 3132 3380
rect 3318 3384 3324 3385
rect 3318 3380 3319 3384
rect 3323 3380 3324 3384
rect 3318 3379 3324 3380
rect 3510 3384 3516 3385
rect 3510 3380 3511 3384
rect 3515 3380 3516 3384
rect 3510 3379 3516 3380
rect 3678 3384 3684 3385
rect 3678 3380 3679 3384
rect 3683 3380 3684 3384
rect 3678 3379 3684 3380
rect 3128 3331 3130 3379
rect 3320 3331 3322 3379
rect 3512 3331 3514 3379
rect 3680 3331 3682 3379
rect 3740 3352 3742 3434
rect 3800 3401 3802 3461
rect 3840 3411 3842 3479
rect 5380 3411 5382 3480
rect 5516 3411 5518 3480
rect 5530 3475 5536 3476
rect 5530 3471 5531 3475
rect 5535 3471 5536 3475
rect 5530 3470 5536 3471
rect 5532 3444 5534 3470
rect 5552 3460 5554 3626
rect 5664 3625 5666 3685
rect 5662 3624 5668 3625
rect 5662 3620 5663 3624
rect 5667 3620 5668 3624
rect 5662 3619 5668 3620
rect 5662 3607 5668 3608
rect 5662 3603 5663 3607
rect 5667 3603 5668 3607
rect 5662 3602 5668 3603
rect 5664 3531 5666 3602
rect 5663 3530 5667 3531
rect 5663 3525 5667 3526
rect 5664 3502 5666 3525
rect 5662 3501 5668 3502
rect 5662 3497 5663 3501
rect 5667 3497 5668 3501
rect 5662 3496 5668 3497
rect 5662 3484 5668 3485
rect 5662 3480 5663 3484
rect 5667 3480 5668 3484
rect 5662 3479 5668 3480
rect 5602 3475 5608 3476
rect 5602 3471 5603 3475
rect 5607 3471 5608 3475
rect 5602 3470 5608 3471
rect 5550 3459 5556 3460
rect 5550 3455 5551 3459
rect 5555 3455 5556 3459
rect 5550 3454 5556 3455
rect 5530 3443 5536 3444
rect 5530 3439 5531 3443
rect 5535 3439 5536 3443
rect 5530 3438 5536 3439
rect 3839 3410 3843 3411
rect 3839 3405 3843 3406
rect 3859 3410 3863 3411
rect 3859 3405 3863 3406
rect 4099 3410 4103 3411
rect 4099 3405 4103 3406
rect 4347 3410 4351 3411
rect 4347 3405 4351 3406
rect 4587 3410 4591 3411
rect 4587 3405 4591 3406
rect 4811 3410 4815 3411
rect 4811 3405 4815 3406
rect 5027 3410 5031 3411
rect 5027 3405 5031 3406
rect 5235 3410 5239 3411
rect 5235 3405 5239 3406
rect 5379 3410 5383 3411
rect 5379 3405 5383 3406
rect 5451 3410 5455 3411
rect 5451 3405 5455 3406
rect 5515 3410 5519 3411
rect 5515 3405 5519 3406
rect 3798 3400 3804 3401
rect 3798 3396 3799 3400
rect 3803 3396 3804 3400
rect 3798 3395 3804 3396
rect 3798 3383 3804 3384
rect 3798 3379 3799 3383
rect 3803 3379 3804 3383
rect 3798 3378 3804 3379
rect 3738 3351 3744 3352
rect 3738 3347 3739 3351
rect 3743 3347 3744 3351
rect 3738 3346 3744 3347
rect 3800 3331 3802 3378
rect 3840 3345 3842 3405
rect 3838 3344 3844 3345
rect 3860 3344 3862 3405
rect 4100 3344 4102 3405
rect 4226 3387 4232 3388
rect 4226 3383 4227 3387
rect 4231 3383 4232 3387
rect 4226 3382 4232 3383
rect 3838 3340 3839 3344
rect 3843 3340 3844 3344
rect 3838 3339 3844 3340
rect 3858 3343 3864 3344
rect 3858 3339 3859 3343
rect 3863 3339 3864 3343
rect 3858 3338 3864 3339
rect 4098 3343 4104 3344
rect 4098 3339 4099 3343
rect 4103 3339 4104 3343
rect 4098 3338 4104 3339
rect 3127 3330 3131 3331
rect 3127 3325 3131 3326
rect 3319 3330 3323 3331
rect 3319 3325 3323 3326
rect 3359 3330 3363 3331
rect 3359 3325 3363 3326
rect 3511 3330 3515 3331
rect 3511 3325 3515 3326
rect 3679 3330 3683 3331
rect 3679 3325 3683 3326
rect 3799 3330 3803 3331
rect 3886 3328 3892 3329
rect 3799 3325 3803 3326
rect 3838 3327 3844 3328
rect 3360 3301 3362 3325
rect 3680 3301 3682 3325
rect 3800 3302 3802 3325
rect 3838 3323 3839 3327
rect 3843 3323 3844 3327
rect 3886 3324 3887 3328
rect 3891 3324 3892 3328
rect 3886 3323 3892 3324
rect 4126 3328 4132 3329
rect 4126 3324 4127 3328
rect 4131 3324 4132 3328
rect 4126 3323 4132 3324
rect 3838 3322 3844 3323
rect 3798 3301 3804 3302
rect 3358 3300 3364 3301
rect 3358 3296 3359 3300
rect 3363 3296 3364 3300
rect 3358 3295 3364 3296
rect 3678 3300 3684 3301
rect 3678 3296 3679 3300
rect 3683 3296 3684 3300
rect 3798 3297 3799 3301
rect 3803 3297 3804 3301
rect 3840 3299 3842 3322
rect 3888 3299 3890 3323
rect 4128 3299 4130 3323
rect 3798 3296 3804 3297
rect 3839 3298 3843 3299
rect 3678 3295 3684 3296
rect 3839 3293 3843 3294
rect 3887 3298 3891 3299
rect 3887 3293 3891 3294
rect 4127 3298 4131 3299
rect 4127 3293 4131 3294
rect 3330 3285 3336 3286
rect 3330 3281 3331 3285
rect 3335 3281 3336 3285
rect 3330 3280 3336 3281
rect 3650 3285 3656 3286
rect 3650 3281 3651 3285
rect 3655 3281 3656 3285
rect 3650 3280 3656 3281
rect 3798 3284 3804 3285
rect 3798 3280 3799 3284
rect 3803 3280 3804 3284
rect 3182 3275 3188 3276
rect 3182 3271 3183 3275
rect 3187 3271 3188 3275
rect 3182 3270 3188 3271
rect 3184 3244 3186 3270
rect 3030 3243 3036 3244
rect 3030 3239 3031 3243
rect 3035 3239 3036 3243
rect 3030 3238 3036 3239
rect 3182 3243 3188 3244
rect 3182 3239 3183 3243
rect 3187 3239 3188 3243
rect 3182 3238 3188 3239
rect 3332 3219 3334 3280
rect 3652 3219 3654 3280
rect 3798 3279 3804 3280
rect 3778 3275 3784 3276
rect 3778 3271 3779 3275
rect 3783 3271 3784 3275
rect 3778 3270 3784 3271
rect 3738 3243 3744 3244
rect 3738 3239 3739 3243
rect 3743 3239 3744 3243
rect 3738 3238 3744 3239
rect 2771 3218 2775 3219
rect 2771 3213 2775 3214
rect 2987 3218 2991 3219
rect 2987 3213 2991 3214
rect 3211 3218 3215 3219
rect 3211 3213 3215 3214
rect 3331 3218 3335 3219
rect 3331 3213 3335 3214
rect 3443 3218 3447 3219
rect 3443 3213 3447 3214
rect 3651 3218 3655 3219
rect 3651 3213 3655 3214
rect 2682 3203 2688 3204
rect 2682 3199 2683 3203
rect 2687 3199 2688 3203
rect 2682 3198 2688 3199
rect 2682 3195 2688 3196
rect 2682 3191 2683 3195
rect 2687 3191 2688 3195
rect 2682 3190 2688 3191
rect 2684 3160 2686 3190
rect 2682 3159 2688 3160
rect 2682 3155 2683 3159
rect 2687 3155 2688 3159
rect 2682 3154 2688 3155
rect 2772 3152 2774 3213
rect 2914 3159 2920 3160
rect 2914 3155 2915 3159
rect 2919 3155 2920 3159
rect 2914 3154 2920 3155
rect 1974 3148 1975 3152
rect 1979 3148 1980 3152
rect 1974 3147 1980 3148
rect 1994 3151 2000 3152
rect 1994 3147 1995 3151
rect 1999 3147 2000 3151
rect 1994 3146 2000 3147
rect 2146 3151 2152 3152
rect 2146 3147 2147 3151
rect 2151 3147 2152 3151
rect 2146 3146 2152 3147
rect 2346 3151 2352 3152
rect 2346 3147 2347 3151
rect 2351 3147 2352 3151
rect 2346 3146 2352 3147
rect 2554 3151 2560 3152
rect 2554 3147 2555 3151
rect 2559 3147 2560 3151
rect 2554 3146 2560 3147
rect 2770 3151 2776 3152
rect 2770 3147 2771 3151
rect 2775 3147 2776 3151
rect 2770 3146 2776 3147
rect 1935 3138 1939 3139
rect 2022 3136 2028 3137
rect 1935 3133 1939 3134
rect 1974 3135 1980 3136
rect 1914 3079 1920 3080
rect 1914 3075 1915 3079
rect 1919 3075 1920 3079
rect 1914 3074 1920 3075
rect 1936 3073 1938 3133
rect 1974 3131 1975 3135
rect 1979 3131 1980 3135
rect 2022 3132 2023 3136
rect 2027 3132 2028 3136
rect 2022 3131 2028 3132
rect 2174 3136 2180 3137
rect 2174 3132 2175 3136
rect 2179 3132 2180 3136
rect 2174 3131 2180 3132
rect 2374 3136 2380 3137
rect 2374 3132 2375 3136
rect 2379 3132 2380 3136
rect 2374 3131 2380 3132
rect 2582 3136 2588 3137
rect 2582 3132 2583 3136
rect 2587 3132 2588 3136
rect 2582 3131 2588 3132
rect 2798 3136 2804 3137
rect 2798 3132 2799 3136
rect 2803 3132 2804 3136
rect 2798 3131 2804 3132
rect 1974 3130 1980 3131
rect 1976 3107 1978 3130
rect 2024 3107 2026 3131
rect 2176 3107 2178 3131
rect 2376 3107 2378 3131
rect 2584 3107 2586 3131
rect 2800 3107 2802 3131
rect 1975 3106 1979 3107
rect 1975 3101 1979 3102
rect 2023 3106 2027 3107
rect 2023 3101 2027 3102
rect 2175 3106 2179 3107
rect 2175 3101 2179 3102
rect 2375 3106 2379 3107
rect 2375 3101 2379 3102
rect 2583 3106 2587 3107
rect 2583 3101 2587 3102
rect 2647 3106 2651 3107
rect 2647 3101 2651 3102
rect 2783 3106 2787 3107
rect 2783 3101 2787 3102
rect 2799 3106 2803 3107
rect 2799 3101 2803 3102
rect 1976 3078 1978 3101
rect 1974 3077 1980 3078
rect 2648 3077 2650 3101
rect 2784 3077 2786 3101
rect 1974 3073 1975 3077
rect 1979 3073 1980 3077
rect 1934 3072 1940 3073
rect 1974 3072 1980 3073
rect 2646 3076 2652 3077
rect 2646 3072 2647 3076
rect 2651 3072 2652 3076
rect 1578 3071 1584 3072
rect 1578 3067 1579 3071
rect 1583 3067 1584 3071
rect 1578 3066 1584 3067
rect 1786 3071 1792 3072
rect 1786 3067 1787 3071
rect 1791 3067 1792 3071
rect 1934 3068 1935 3072
rect 1939 3068 1940 3072
rect 2646 3071 2652 3072
rect 2782 3076 2788 3077
rect 2782 3072 2783 3076
rect 2787 3072 2788 3076
rect 2782 3071 2788 3072
rect 1934 3067 1940 3068
rect 1786 3066 1792 3067
rect 2618 3061 2624 3062
rect 1974 3060 1980 3061
rect 1606 3056 1612 3057
rect 1606 3052 1607 3056
rect 1611 3052 1612 3056
rect 1606 3051 1612 3052
rect 1814 3056 1820 3057
rect 1974 3056 1975 3060
rect 1979 3056 1980 3060
rect 2618 3057 2619 3061
rect 2623 3057 2624 3061
rect 2618 3056 2624 3057
rect 2754 3061 2760 3062
rect 2754 3057 2755 3061
rect 2759 3057 2760 3061
rect 2754 3056 2760 3057
rect 2898 3061 2904 3062
rect 2898 3057 2899 3061
rect 2903 3057 2904 3061
rect 2898 3056 2904 3057
rect 1814 3052 1815 3056
rect 1819 3052 1820 3056
rect 1814 3051 1820 3052
rect 1934 3055 1940 3056
rect 1974 3055 1980 3056
rect 1934 3051 1935 3055
rect 1939 3051 1940 3055
rect 1608 3027 1610 3051
rect 1816 3027 1818 3051
rect 1934 3050 1940 3051
rect 1936 3027 1938 3050
rect 1511 3026 1515 3027
rect 1511 3021 1515 3022
rect 1607 3026 1611 3027
rect 1607 3021 1611 3022
rect 1671 3026 1675 3027
rect 1671 3021 1675 3022
rect 1815 3026 1819 3027
rect 1815 3021 1819 3022
rect 1935 3026 1939 3027
rect 1935 3021 1939 3022
rect 1450 3011 1456 3012
rect 1450 3007 1451 3011
rect 1455 3007 1456 3011
rect 1450 3006 1456 3007
rect 1512 2997 1514 3021
rect 1672 2997 1674 3021
rect 1816 2997 1818 3021
rect 1910 3011 1916 3012
rect 1910 3007 1911 3011
rect 1915 3007 1916 3011
rect 1910 3006 1916 3007
rect 822 2996 828 2997
rect 822 2992 823 2996
rect 827 2992 828 2996
rect 822 2991 828 2992
rect 1006 2996 1012 2997
rect 1006 2992 1007 2996
rect 1011 2992 1012 2996
rect 1006 2991 1012 2992
rect 1182 2996 1188 2997
rect 1182 2992 1183 2996
rect 1187 2992 1188 2996
rect 1182 2991 1188 2992
rect 1350 2996 1356 2997
rect 1350 2992 1351 2996
rect 1355 2992 1356 2996
rect 1350 2991 1356 2992
rect 1510 2996 1516 2997
rect 1510 2992 1511 2996
rect 1515 2992 1516 2996
rect 1510 2991 1516 2992
rect 1670 2996 1676 2997
rect 1670 2992 1671 2996
rect 1675 2992 1676 2996
rect 1670 2991 1676 2992
rect 1814 2996 1820 2997
rect 1814 2992 1815 2996
rect 1819 2992 1820 2996
rect 1814 2991 1820 2992
rect 794 2981 800 2982
rect 794 2977 795 2981
rect 799 2977 800 2981
rect 794 2976 800 2977
rect 978 2981 984 2982
rect 978 2977 979 2981
rect 983 2977 984 2981
rect 978 2976 984 2977
rect 1154 2981 1160 2982
rect 1154 2977 1155 2981
rect 1159 2977 1160 2981
rect 1154 2976 1160 2977
rect 1322 2981 1328 2982
rect 1322 2977 1323 2981
rect 1327 2977 1328 2981
rect 1322 2976 1328 2977
rect 1482 2981 1488 2982
rect 1482 2977 1483 2981
rect 1487 2977 1488 2981
rect 1482 2976 1488 2977
rect 1642 2981 1648 2982
rect 1642 2977 1643 2981
rect 1647 2977 1648 2981
rect 1642 2976 1648 2977
rect 1786 2981 1792 2982
rect 1786 2977 1787 2981
rect 1791 2977 1792 2981
rect 1786 2976 1792 2977
rect 682 2939 688 2940
rect 682 2935 683 2939
rect 687 2935 688 2939
rect 682 2934 688 2935
rect 796 2911 798 2976
rect 810 2971 816 2972
rect 810 2967 811 2971
rect 815 2967 816 2971
rect 810 2966 816 2967
rect 812 2940 814 2966
rect 906 2963 912 2964
rect 906 2959 907 2963
rect 911 2959 912 2963
rect 906 2958 912 2959
rect 810 2939 816 2940
rect 810 2935 811 2939
rect 815 2935 816 2939
rect 810 2934 816 2935
rect 595 2910 599 2911
rect 595 2905 599 2906
rect 787 2910 791 2911
rect 787 2905 791 2906
rect 795 2910 799 2911
rect 795 2905 799 2906
rect 466 2851 472 2852
rect 466 2847 467 2851
rect 471 2847 472 2851
rect 466 2846 472 2847
rect 596 2844 598 2905
rect 682 2883 688 2884
rect 682 2879 683 2883
rect 687 2879 688 2883
rect 682 2878 688 2879
rect 110 2840 111 2844
rect 115 2840 116 2844
rect 110 2839 116 2840
rect 394 2843 400 2844
rect 394 2839 395 2843
rect 399 2839 400 2843
rect 394 2838 400 2839
rect 594 2843 600 2844
rect 594 2839 595 2843
rect 599 2839 600 2843
rect 594 2838 600 2839
rect 422 2828 428 2829
rect 110 2827 116 2828
rect 110 2823 111 2827
rect 115 2823 116 2827
rect 422 2824 423 2828
rect 427 2824 428 2828
rect 422 2823 428 2824
rect 622 2828 628 2829
rect 622 2824 623 2828
rect 627 2824 628 2828
rect 622 2823 628 2824
rect 110 2822 116 2823
rect 112 2787 114 2822
rect 424 2787 426 2823
rect 624 2787 626 2823
rect 111 2786 115 2787
rect 111 2781 115 2782
rect 423 2786 427 2787
rect 423 2781 427 2782
rect 623 2786 627 2787
rect 623 2781 627 2782
rect 655 2786 659 2787
rect 655 2781 659 2782
rect 112 2758 114 2781
rect 110 2757 116 2758
rect 656 2757 658 2781
rect 110 2753 111 2757
rect 115 2753 116 2757
rect 110 2752 116 2753
rect 654 2756 660 2757
rect 654 2752 655 2756
rect 659 2752 660 2756
rect 654 2751 660 2752
rect 626 2741 632 2742
rect 110 2740 116 2741
rect 110 2736 111 2740
rect 115 2736 116 2740
rect 626 2737 627 2741
rect 631 2737 632 2741
rect 626 2736 632 2737
rect 110 2735 116 2736
rect 112 2675 114 2735
rect 628 2675 630 2736
rect 684 2732 686 2878
rect 788 2844 790 2905
rect 908 2888 910 2958
rect 980 2911 982 2976
rect 994 2971 1000 2972
rect 994 2967 995 2971
rect 999 2967 1000 2971
rect 994 2966 1000 2967
rect 996 2940 998 2966
rect 994 2939 1000 2940
rect 994 2935 995 2939
rect 999 2935 1000 2939
rect 994 2934 1000 2935
rect 1156 2911 1158 2976
rect 1324 2911 1326 2976
rect 1338 2971 1344 2972
rect 1338 2967 1339 2971
rect 1343 2967 1344 2971
rect 1338 2966 1344 2967
rect 1340 2940 1342 2966
rect 1338 2939 1344 2940
rect 1338 2935 1339 2939
rect 1343 2935 1344 2939
rect 1338 2934 1344 2935
rect 1484 2911 1486 2976
rect 1498 2971 1504 2972
rect 1498 2967 1499 2971
rect 1503 2967 1504 2971
rect 1498 2966 1504 2967
rect 1500 2940 1502 2966
rect 1498 2939 1504 2940
rect 1498 2935 1499 2939
rect 1503 2935 1504 2939
rect 1498 2934 1504 2935
rect 1644 2911 1646 2976
rect 1658 2971 1664 2972
rect 1658 2967 1659 2971
rect 1663 2967 1664 2971
rect 1658 2966 1664 2967
rect 1660 2940 1662 2966
rect 1658 2939 1664 2940
rect 1658 2935 1659 2939
rect 1663 2935 1664 2939
rect 1658 2934 1664 2935
rect 1788 2911 1790 2976
rect 1912 2972 1914 3006
rect 1936 2998 1938 3021
rect 1934 2997 1940 2998
rect 1934 2993 1935 2997
rect 1939 2993 1940 2997
rect 1976 2995 1978 3055
rect 2620 2995 2622 3056
rect 2756 2995 2758 3056
rect 2770 3051 2776 3052
rect 2770 3047 2771 3051
rect 2775 3047 2776 3051
rect 2770 3046 2776 3047
rect 2890 3051 2896 3052
rect 2890 3047 2891 3051
rect 2895 3047 2896 3051
rect 2890 3046 2896 3047
rect 2772 3020 2774 3046
rect 2770 3019 2776 3020
rect 2770 3015 2771 3019
rect 2775 3015 2776 3019
rect 2770 3014 2776 3015
rect 1934 2992 1940 2993
rect 1975 2994 1979 2995
rect 1975 2989 1979 2990
rect 2619 2994 2623 2995
rect 2619 2989 2623 2990
rect 2755 2994 2759 2995
rect 2755 2989 2759 2990
rect 2803 2994 2807 2995
rect 2803 2989 2807 2990
rect 1934 2980 1940 2981
rect 1934 2976 1935 2980
rect 1939 2976 1940 2980
rect 1934 2975 1940 2976
rect 1802 2971 1808 2972
rect 1802 2967 1803 2971
rect 1807 2967 1808 2971
rect 1802 2966 1808 2967
rect 1910 2971 1916 2972
rect 1910 2967 1911 2971
rect 1915 2967 1916 2971
rect 1910 2966 1916 2967
rect 1804 2940 1806 2966
rect 1802 2939 1808 2940
rect 1802 2935 1803 2939
rect 1807 2935 1808 2939
rect 1802 2934 1808 2935
rect 1936 2911 1938 2975
rect 1976 2929 1978 2989
rect 1974 2928 1980 2929
rect 2804 2928 2806 2989
rect 2892 2968 2894 3046
rect 2900 2995 2902 3056
rect 2916 3020 2918 3154
rect 2988 3152 2990 3213
rect 3022 3159 3028 3160
rect 3022 3155 3023 3159
rect 3027 3155 3028 3159
rect 3022 3154 3028 3155
rect 2986 3151 2992 3152
rect 2986 3147 2987 3151
rect 2991 3147 2992 3151
rect 2986 3146 2992 3147
rect 3014 3136 3020 3137
rect 3014 3132 3015 3136
rect 3019 3132 3020 3136
rect 3014 3131 3020 3132
rect 3016 3107 3018 3131
rect 2927 3106 2931 3107
rect 2927 3101 2931 3102
rect 3015 3106 3019 3107
rect 3015 3101 3019 3102
rect 2928 3077 2930 3101
rect 2926 3076 2932 3077
rect 2926 3072 2927 3076
rect 2931 3072 2932 3076
rect 2926 3071 2932 3072
rect 3024 3036 3026 3154
rect 3212 3152 3214 3213
rect 3414 3195 3420 3196
rect 3414 3191 3415 3195
rect 3419 3191 3420 3195
rect 3414 3190 3420 3191
rect 3382 3187 3388 3188
rect 3382 3183 3383 3187
rect 3387 3183 3388 3187
rect 3382 3182 3388 3183
rect 3210 3151 3216 3152
rect 3210 3147 3211 3151
rect 3215 3147 3216 3151
rect 3210 3146 3216 3147
rect 3238 3136 3244 3137
rect 3238 3132 3239 3136
rect 3243 3132 3244 3136
rect 3238 3131 3244 3132
rect 3240 3107 3242 3131
rect 3079 3106 3083 3107
rect 3079 3101 3083 3102
rect 3239 3106 3243 3107
rect 3239 3101 3243 3102
rect 3080 3077 3082 3101
rect 3240 3077 3242 3101
rect 3078 3076 3084 3077
rect 3078 3072 3079 3076
rect 3083 3072 3084 3076
rect 3078 3071 3084 3072
rect 3238 3076 3244 3077
rect 3238 3072 3239 3076
rect 3243 3072 3244 3076
rect 3238 3071 3244 3072
rect 3050 3061 3056 3062
rect 3050 3057 3051 3061
rect 3055 3057 3056 3061
rect 3050 3056 3056 3057
rect 3210 3061 3216 3062
rect 3210 3057 3211 3061
rect 3215 3057 3216 3061
rect 3210 3056 3216 3057
rect 3370 3061 3376 3062
rect 3370 3057 3371 3061
rect 3375 3057 3376 3061
rect 3370 3056 3376 3057
rect 3022 3035 3028 3036
rect 3022 3031 3023 3035
rect 3027 3031 3028 3035
rect 3022 3030 3028 3031
rect 2914 3019 2920 3020
rect 2914 3015 2915 3019
rect 2919 3015 2920 3019
rect 2914 3014 2920 3015
rect 3052 2995 3054 3056
rect 3066 3051 3072 3052
rect 3066 3047 3067 3051
rect 3071 3047 3072 3051
rect 3066 3046 3072 3047
rect 3068 3020 3070 3046
rect 3066 3019 3072 3020
rect 3066 3015 3067 3019
rect 3071 3015 3072 3019
rect 3066 3014 3072 3015
rect 3212 2995 3214 3056
rect 3226 3051 3232 3052
rect 3226 3047 3227 3051
rect 3231 3047 3232 3051
rect 3226 3046 3232 3047
rect 3228 3020 3230 3046
rect 3226 3019 3232 3020
rect 3226 3015 3227 3019
rect 3231 3015 3232 3019
rect 3226 3014 3232 3015
rect 3372 2995 3374 3056
rect 3384 3052 3386 3182
rect 3416 3160 3418 3190
rect 3414 3159 3420 3160
rect 3414 3155 3415 3159
rect 3419 3155 3420 3159
rect 3414 3154 3420 3155
rect 3444 3152 3446 3213
rect 3570 3195 3576 3196
rect 3570 3191 3571 3195
rect 3575 3191 3576 3195
rect 3570 3190 3576 3191
rect 3572 3160 3574 3190
rect 3570 3159 3576 3160
rect 3570 3155 3571 3159
rect 3575 3155 3576 3159
rect 3570 3154 3576 3155
rect 3652 3152 3654 3213
rect 3740 3160 3742 3238
rect 3780 3212 3782 3270
rect 3800 3219 3802 3279
rect 3840 3270 3842 3293
rect 3838 3269 3844 3270
rect 3888 3269 3890 3293
rect 4128 3269 4130 3293
rect 3838 3265 3839 3269
rect 3843 3265 3844 3269
rect 3838 3264 3844 3265
rect 3886 3268 3892 3269
rect 3886 3264 3887 3268
rect 3891 3264 3892 3268
rect 3886 3263 3892 3264
rect 4126 3268 4132 3269
rect 4126 3264 4127 3268
rect 4131 3264 4132 3268
rect 4126 3263 4132 3264
rect 3858 3253 3864 3254
rect 3838 3252 3844 3253
rect 3838 3248 3839 3252
rect 3843 3248 3844 3252
rect 3858 3249 3859 3253
rect 3863 3249 3864 3253
rect 3858 3248 3864 3249
rect 4098 3253 4104 3254
rect 4098 3249 4099 3253
rect 4103 3249 4104 3253
rect 4098 3248 4104 3249
rect 3838 3247 3844 3248
rect 3799 3218 3803 3219
rect 3799 3213 3803 3214
rect 3778 3211 3784 3212
rect 3778 3207 3779 3211
rect 3783 3207 3784 3211
rect 3778 3206 3784 3207
rect 3738 3159 3744 3160
rect 3738 3155 3739 3159
rect 3743 3155 3744 3159
rect 3738 3154 3744 3155
rect 3800 3153 3802 3213
rect 3840 3171 3842 3247
rect 3860 3171 3862 3248
rect 4100 3171 4102 3248
rect 4228 3244 4230 3382
rect 4294 3379 4300 3380
rect 4294 3375 4295 3379
rect 4299 3375 4300 3379
rect 4294 3374 4300 3375
rect 4296 3352 4298 3374
rect 4294 3351 4300 3352
rect 4294 3347 4295 3351
rect 4299 3347 4300 3351
rect 4294 3346 4300 3347
rect 4348 3344 4350 3405
rect 4588 3344 4590 3405
rect 4674 3383 4680 3384
rect 4674 3379 4675 3383
rect 4679 3379 4680 3383
rect 4674 3378 4680 3379
rect 4676 3360 4678 3378
rect 4674 3359 4680 3360
rect 4674 3355 4675 3359
rect 4679 3355 4680 3359
rect 4674 3354 4680 3355
rect 4802 3351 4808 3352
rect 4802 3347 4803 3351
rect 4807 3347 4808 3351
rect 4802 3346 4808 3347
rect 4346 3343 4352 3344
rect 4346 3339 4347 3343
rect 4351 3339 4352 3343
rect 4346 3338 4352 3339
rect 4586 3343 4592 3344
rect 4586 3339 4587 3343
rect 4591 3339 4592 3343
rect 4586 3338 4592 3339
rect 4374 3328 4380 3329
rect 4374 3324 4375 3328
rect 4379 3324 4380 3328
rect 4374 3323 4380 3324
rect 4614 3328 4620 3329
rect 4614 3324 4615 3328
rect 4619 3324 4620 3328
rect 4614 3323 4620 3324
rect 4376 3299 4378 3323
rect 4616 3299 4618 3323
rect 4375 3298 4379 3299
rect 4375 3293 4379 3294
rect 4607 3298 4611 3299
rect 4607 3293 4611 3294
rect 4615 3298 4619 3299
rect 4615 3293 4619 3294
rect 4376 3269 4378 3293
rect 4608 3269 4610 3293
rect 4374 3268 4380 3269
rect 4374 3264 4375 3268
rect 4379 3264 4380 3268
rect 4374 3263 4380 3264
rect 4606 3268 4612 3269
rect 4606 3264 4607 3268
rect 4611 3264 4612 3268
rect 4606 3263 4612 3264
rect 4346 3253 4352 3254
rect 4346 3249 4347 3253
rect 4351 3249 4352 3253
rect 4346 3248 4352 3249
rect 4578 3253 4584 3254
rect 4578 3249 4579 3253
rect 4583 3249 4584 3253
rect 4578 3248 4584 3249
rect 4786 3253 4792 3254
rect 4786 3249 4787 3253
rect 4791 3249 4792 3253
rect 4786 3248 4792 3249
rect 4114 3243 4120 3244
rect 4114 3239 4115 3243
rect 4119 3239 4120 3243
rect 4114 3238 4120 3239
rect 4226 3243 4232 3244
rect 4226 3239 4227 3243
rect 4231 3239 4232 3243
rect 4226 3238 4232 3239
rect 4116 3212 4118 3238
rect 4114 3211 4120 3212
rect 4114 3207 4115 3211
rect 4119 3207 4120 3211
rect 4114 3206 4120 3207
rect 4348 3171 4350 3248
rect 4434 3235 4440 3236
rect 4434 3231 4435 3235
rect 4439 3231 4440 3235
rect 4434 3230 4440 3231
rect 4436 3212 4438 3230
rect 4434 3211 4440 3212
rect 4434 3207 4435 3211
rect 4439 3207 4440 3211
rect 4434 3206 4440 3207
rect 4580 3171 4582 3248
rect 4594 3243 4600 3244
rect 4594 3239 4595 3243
rect 4599 3239 4600 3243
rect 4594 3238 4600 3239
rect 4758 3243 4764 3244
rect 4758 3239 4759 3243
rect 4763 3239 4764 3243
rect 4758 3238 4764 3239
rect 4596 3212 4598 3238
rect 4594 3211 4600 3212
rect 4594 3207 4595 3211
rect 4599 3207 4600 3211
rect 4594 3206 4600 3207
rect 3839 3170 3843 3171
rect 3839 3165 3843 3166
rect 3859 3170 3863 3171
rect 3859 3165 3863 3166
rect 4099 3170 4103 3171
rect 4099 3165 4103 3166
rect 4347 3170 4351 3171
rect 4347 3165 4351 3166
rect 4467 3170 4471 3171
rect 4467 3165 4471 3166
rect 4579 3170 4583 3171
rect 4579 3165 4583 3166
rect 4651 3170 4655 3171
rect 4651 3165 4655 3166
rect 3798 3152 3804 3153
rect 3442 3151 3448 3152
rect 3442 3147 3443 3151
rect 3447 3147 3448 3151
rect 3442 3146 3448 3147
rect 3650 3151 3656 3152
rect 3650 3147 3651 3151
rect 3655 3147 3656 3151
rect 3798 3148 3799 3152
rect 3803 3148 3804 3152
rect 3798 3147 3804 3148
rect 3650 3146 3656 3147
rect 3470 3136 3476 3137
rect 3470 3132 3471 3136
rect 3475 3132 3476 3136
rect 3470 3131 3476 3132
rect 3678 3136 3684 3137
rect 3678 3132 3679 3136
rect 3683 3132 3684 3136
rect 3678 3131 3684 3132
rect 3798 3135 3804 3136
rect 3798 3131 3799 3135
rect 3803 3131 3804 3135
rect 3472 3107 3474 3131
rect 3680 3107 3682 3131
rect 3798 3130 3804 3131
rect 3800 3107 3802 3130
rect 3399 3106 3403 3107
rect 3399 3101 3403 3102
rect 3471 3106 3475 3107
rect 3471 3101 3475 3102
rect 3567 3106 3571 3107
rect 3567 3101 3571 3102
rect 3679 3106 3683 3107
rect 3679 3101 3683 3102
rect 3799 3106 3803 3107
rect 3840 3105 3842 3165
rect 3799 3101 3803 3102
rect 3838 3104 3844 3105
rect 4468 3104 4470 3165
rect 4554 3143 4560 3144
rect 4554 3139 4555 3143
rect 4559 3139 4560 3143
rect 4554 3138 4560 3139
rect 4556 3120 4558 3138
rect 4554 3119 4560 3120
rect 4554 3115 4555 3119
rect 4559 3115 4560 3119
rect 4554 3114 4560 3115
rect 4652 3104 4654 3165
rect 4760 3148 4762 3238
rect 4788 3171 4790 3248
rect 4804 3212 4806 3346
rect 4812 3344 4814 3405
rect 4990 3387 4996 3388
rect 4990 3383 4991 3387
rect 4995 3383 4996 3387
rect 4990 3382 4996 3383
rect 4992 3352 4994 3382
rect 4990 3351 4996 3352
rect 4990 3347 4991 3351
rect 4995 3347 4996 3351
rect 4990 3346 4996 3347
rect 5028 3344 5030 3405
rect 5236 3344 5238 3405
rect 5414 3387 5420 3388
rect 5414 3383 5415 3387
rect 5419 3383 5420 3387
rect 5414 3382 5420 3383
rect 5442 3387 5448 3388
rect 5442 3383 5443 3387
rect 5447 3383 5448 3387
rect 5442 3382 5448 3383
rect 5416 3352 5418 3382
rect 5414 3351 5420 3352
rect 5414 3347 5415 3351
rect 5419 3347 5420 3351
rect 5414 3346 5420 3347
rect 4810 3343 4816 3344
rect 4810 3339 4811 3343
rect 4815 3339 4816 3343
rect 4810 3338 4816 3339
rect 5026 3343 5032 3344
rect 5026 3339 5027 3343
rect 5031 3339 5032 3343
rect 5026 3338 5032 3339
rect 5234 3343 5240 3344
rect 5234 3339 5235 3343
rect 5239 3339 5240 3343
rect 5234 3338 5240 3339
rect 4838 3328 4844 3329
rect 4838 3324 4839 3328
rect 4843 3324 4844 3328
rect 4838 3323 4844 3324
rect 5054 3328 5060 3329
rect 5054 3324 5055 3328
rect 5059 3324 5060 3328
rect 5054 3323 5060 3324
rect 5262 3328 5268 3329
rect 5262 3324 5263 3328
rect 5267 3324 5268 3328
rect 5262 3323 5268 3324
rect 4840 3299 4842 3323
rect 5056 3299 5058 3323
rect 5264 3299 5266 3323
rect 4815 3298 4819 3299
rect 4815 3293 4819 3294
rect 4839 3298 4843 3299
rect 4839 3293 4843 3294
rect 5015 3298 5019 3299
rect 5015 3293 5019 3294
rect 5055 3298 5059 3299
rect 5055 3293 5059 3294
rect 5199 3298 5203 3299
rect 5199 3293 5203 3294
rect 5263 3298 5267 3299
rect 5263 3293 5267 3294
rect 5383 3298 5387 3299
rect 5383 3293 5387 3294
rect 4816 3269 4818 3293
rect 5016 3269 5018 3293
rect 5200 3269 5202 3293
rect 5384 3269 5386 3293
rect 4814 3268 4820 3269
rect 4814 3264 4815 3268
rect 4819 3264 4820 3268
rect 4814 3263 4820 3264
rect 5014 3268 5020 3269
rect 5014 3264 5015 3268
rect 5019 3264 5020 3268
rect 5014 3263 5020 3264
rect 5198 3268 5204 3269
rect 5198 3264 5199 3268
rect 5203 3264 5204 3268
rect 5198 3263 5204 3264
rect 5382 3268 5388 3269
rect 5382 3264 5383 3268
rect 5387 3264 5388 3268
rect 5382 3263 5388 3264
rect 4986 3253 4992 3254
rect 4986 3249 4987 3253
rect 4991 3249 4992 3253
rect 4986 3248 4992 3249
rect 5170 3253 5176 3254
rect 5170 3249 5171 3253
rect 5175 3249 5176 3253
rect 5170 3248 5176 3249
rect 5354 3253 5360 3254
rect 5354 3249 5355 3253
rect 5359 3249 5360 3253
rect 5354 3248 5360 3249
rect 4802 3211 4808 3212
rect 4802 3207 4803 3211
rect 4807 3207 4808 3211
rect 4802 3206 4808 3207
rect 4988 3171 4990 3248
rect 5002 3243 5008 3244
rect 5002 3239 5003 3243
rect 5007 3239 5008 3243
rect 5002 3238 5008 3239
rect 5004 3212 5006 3238
rect 5002 3211 5008 3212
rect 5002 3207 5003 3211
rect 5007 3207 5008 3211
rect 5002 3206 5008 3207
rect 5172 3171 5174 3248
rect 5356 3171 5358 3248
rect 5444 3244 5446 3382
rect 5452 3344 5454 3405
rect 5450 3343 5456 3344
rect 5450 3339 5451 3343
rect 5455 3339 5456 3343
rect 5450 3338 5456 3339
rect 5478 3328 5484 3329
rect 5478 3324 5479 3328
rect 5483 3324 5484 3328
rect 5478 3323 5484 3324
rect 5480 3299 5482 3323
rect 5479 3298 5483 3299
rect 5479 3293 5483 3294
rect 5543 3298 5547 3299
rect 5543 3293 5547 3294
rect 5544 3269 5546 3293
rect 5542 3268 5548 3269
rect 5542 3264 5543 3268
rect 5547 3264 5548 3268
rect 5542 3263 5548 3264
rect 5514 3253 5520 3254
rect 5514 3249 5515 3253
rect 5519 3249 5520 3253
rect 5514 3248 5520 3249
rect 5370 3243 5376 3244
rect 5370 3239 5371 3243
rect 5375 3239 5376 3243
rect 5370 3238 5376 3239
rect 5442 3243 5448 3244
rect 5442 3239 5443 3243
rect 5447 3239 5448 3243
rect 5442 3238 5448 3239
rect 5372 3212 5374 3238
rect 5362 3211 5368 3212
rect 5362 3207 5363 3211
rect 5367 3207 5368 3211
rect 5362 3206 5368 3207
rect 5370 3211 5376 3212
rect 5370 3207 5371 3211
rect 5375 3207 5376 3211
rect 5370 3206 5376 3207
rect 4787 3170 4791 3171
rect 4787 3165 4791 3166
rect 4859 3170 4863 3171
rect 4859 3165 4863 3166
rect 4987 3170 4991 3171
rect 4987 3165 4991 3166
rect 5075 3170 5079 3171
rect 5075 3165 5079 3166
rect 5171 3170 5175 3171
rect 5171 3165 5175 3166
rect 5307 3170 5311 3171
rect 5307 3165 5311 3166
rect 5355 3170 5359 3171
rect 5355 3165 5359 3166
rect 4758 3147 4764 3148
rect 4758 3143 4759 3147
rect 4763 3143 4764 3147
rect 4758 3142 4764 3143
rect 4658 3111 4664 3112
rect 4658 3107 4659 3111
rect 4663 3107 4664 3111
rect 4658 3106 4664 3107
rect 3400 3077 3402 3101
rect 3568 3077 3570 3101
rect 3800 3078 3802 3101
rect 3838 3100 3839 3104
rect 3843 3100 3844 3104
rect 3838 3099 3844 3100
rect 4466 3103 4472 3104
rect 4466 3099 4467 3103
rect 4471 3099 4472 3103
rect 4466 3098 4472 3099
rect 4650 3103 4656 3104
rect 4650 3099 4651 3103
rect 4655 3099 4656 3103
rect 4650 3098 4656 3099
rect 4494 3088 4500 3089
rect 3838 3087 3844 3088
rect 3838 3083 3839 3087
rect 3843 3083 3844 3087
rect 4494 3084 4495 3088
rect 4499 3084 4500 3088
rect 4494 3083 4500 3084
rect 3838 3082 3844 3083
rect 3798 3077 3804 3078
rect 3398 3076 3404 3077
rect 3398 3072 3399 3076
rect 3403 3072 3404 3076
rect 3398 3071 3404 3072
rect 3566 3076 3572 3077
rect 3566 3072 3567 3076
rect 3571 3072 3572 3076
rect 3798 3073 3799 3077
rect 3803 3073 3804 3077
rect 3798 3072 3804 3073
rect 3566 3071 3572 3072
rect 3538 3061 3544 3062
rect 3538 3057 3539 3061
rect 3543 3057 3544 3061
rect 3538 3056 3544 3057
rect 3798 3060 3804 3061
rect 3798 3056 3799 3060
rect 3803 3056 3804 3060
rect 3840 3059 3842 3082
rect 4496 3059 4498 3083
rect 3382 3051 3388 3052
rect 3382 3047 3383 3051
rect 3387 3047 3388 3051
rect 3382 3046 3388 3047
rect 3526 3051 3532 3052
rect 3526 3047 3527 3051
rect 3531 3047 3532 3051
rect 3526 3046 3532 3047
rect 3528 3020 3530 3046
rect 3526 3019 3532 3020
rect 3526 3015 3527 3019
rect 3531 3015 3532 3019
rect 3526 3014 3532 3015
rect 3540 2995 3542 3056
rect 3798 3055 3804 3056
rect 3839 3058 3843 3059
rect 3606 3019 3612 3020
rect 3606 3015 3607 3019
rect 3611 3015 3612 3019
rect 3606 3014 3612 3015
rect 2899 2994 2903 2995
rect 2899 2989 2903 2990
rect 2939 2994 2943 2995
rect 2939 2989 2943 2990
rect 3051 2994 3055 2995
rect 3051 2989 3055 2990
rect 3075 2994 3079 2995
rect 3075 2989 3079 2990
rect 3211 2994 3215 2995
rect 3211 2989 3215 2990
rect 3347 2994 3351 2995
rect 3347 2989 3351 2990
rect 3371 2994 3375 2995
rect 3371 2989 3375 2990
rect 3483 2994 3487 2995
rect 3483 2989 3487 2990
rect 3539 2994 3543 2995
rect 3539 2989 3543 2990
rect 2890 2967 2896 2968
rect 2890 2963 2891 2967
rect 2895 2963 2896 2967
rect 2890 2962 2896 2963
rect 2940 2928 2942 2989
rect 3058 2935 3064 2936
rect 3058 2931 3059 2935
rect 3063 2931 3064 2935
rect 3058 2930 3064 2931
rect 1974 2924 1975 2928
rect 1979 2924 1980 2928
rect 1974 2923 1980 2924
rect 2802 2927 2808 2928
rect 2802 2923 2803 2927
rect 2807 2923 2808 2927
rect 2802 2922 2808 2923
rect 2938 2927 2944 2928
rect 2938 2923 2939 2927
rect 2943 2923 2944 2927
rect 2938 2922 2944 2923
rect 2830 2912 2836 2913
rect 1974 2911 1980 2912
rect 971 2910 975 2911
rect 971 2905 975 2906
rect 979 2910 983 2911
rect 979 2905 983 2906
rect 1147 2910 1151 2911
rect 1147 2905 1151 2906
rect 1155 2910 1159 2911
rect 1155 2905 1159 2906
rect 1315 2910 1319 2911
rect 1315 2905 1319 2906
rect 1323 2910 1327 2911
rect 1323 2905 1327 2906
rect 1483 2910 1487 2911
rect 1483 2905 1487 2906
rect 1643 2910 1647 2911
rect 1643 2905 1647 2906
rect 1787 2910 1791 2911
rect 1787 2905 1791 2906
rect 1935 2910 1939 2911
rect 1974 2907 1975 2911
rect 1979 2907 1980 2911
rect 2830 2908 2831 2912
rect 2835 2908 2836 2912
rect 2830 2907 2836 2908
rect 2966 2912 2972 2913
rect 2966 2908 2967 2912
rect 2971 2908 2972 2912
rect 2966 2907 2972 2908
rect 1974 2906 1980 2907
rect 1935 2905 1939 2906
rect 906 2887 912 2888
rect 906 2883 907 2887
rect 911 2883 912 2887
rect 906 2882 912 2883
rect 914 2887 920 2888
rect 914 2883 915 2887
rect 919 2883 920 2887
rect 914 2882 920 2883
rect 916 2852 918 2882
rect 914 2851 920 2852
rect 914 2847 915 2851
rect 919 2847 920 2851
rect 914 2846 920 2847
rect 972 2844 974 2905
rect 1098 2887 1104 2888
rect 1098 2883 1099 2887
rect 1103 2883 1104 2887
rect 1098 2882 1104 2883
rect 1100 2852 1102 2882
rect 1098 2851 1104 2852
rect 1098 2847 1099 2851
rect 1103 2847 1104 2851
rect 1098 2846 1104 2847
rect 1148 2844 1150 2905
rect 1202 2851 1208 2852
rect 1202 2847 1203 2851
rect 1207 2847 1208 2851
rect 1202 2846 1208 2847
rect 786 2843 792 2844
rect 786 2839 787 2843
rect 791 2839 792 2843
rect 786 2838 792 2839
rect 970 2843 976 2844
rect 970 2839 971 2843
rect 975 2839 976 2843
rect 970 2838 976 2839
rect 1146 2843 1152 2844
rect 1146 2839 1147 2843
rect 1151 2839 1152 2843
rect 1146 2838 1152 2839
rect 814 2828 820 2829
rect 814 2824 815 2828
rect 819 2824 820 2828
rect 814 2823 820 2824
rect 998 2828 1004 2829
rect 998 2824 999 2828
rect 1003 2824 1004 2828
rect 998 2823 1004 2824
rect 1174 2828 1180 2829
rect 1174 2824 1175 2828
rect 1179 2824 1180 2828
rect 1174 2823 1180 2824
rect 816 2787 818 2823
rect 1000 2787 1002 2823
rect 1176 2787 1178 2823
rect 815 2786 819 2787
rect 815 2781 819 2782
rect 975 2786 979 2787
rect 975 2781 979 2782
rect 999 2786 1003 2787
rect 999 2781 1003 2782
rect 1143 2786 1147 2787
rect 1143 2781 1147 2782
rect 1175 2786 1179 2787
rect 1175 2781 1179 2782
rect 816 2757 818 2781
rect 976 2757 978 2781
rect 1144 2757 1146 2781
rect 814 2756 820 2757
rect 814 2752 815 2756
rect 819 2752 820 2756
rect 814 2751 820 2752
rect 974 2756 980 2757
rect 974 2752 975 2756
rect 979 2752 980 2756
rect 974 2751 980 2752
rect 1142 2756 1148 2757
rect 1142 2752 1143 2756
rect 1147 2752 1148 2756
rect 1142 2751 1148 2752
rect 786 2741 792 2742
rect 786 2737 787 2741
rect 791 2737 792 2741
rect 786 2736 792 2737
rect 946 2741 952 2742
rect 946 2737 947 2741
rect 951 2737 952 2741
rect 946 2736 952 2737
rect 1114 2741 1120 2742
rect 1114 2737 1115 2741
rect 1119 2737 1120 2741
rect 1114 2736 1120 2737
rect 682 2731 688 2732
rect 682 2727 683 2731
rect 687 2727 688 2731
rect 682 2726 688 2727
rect 788 2675 790 2736
rect 948 2675 950 2736
rect 1030 2699 1036 2700
rect 1030 2695 1031 2699
rect 1035 2695 1036 2699
rect 1030 2694 1036 2695
rect 111 2674 115 2675
rect 111 2669 115 2670
rect 627 2674 631 2675
rect 627 2669 631 2670
rect 771 2674 775 2675
rect 771 2669 775 2670
rect 787 2674 791 2675
rect 787 2669 791 2670
rect 907 2674 911 2675
rect 907 2669 911 2670
rect 947 2674 951 2675
rect 947 2669 951 2670
rect 112 2609 114 2669
rect 110 2608 116 2609
rect 772 2608 774 2669
rect 858 2647 864 2648
rect 858 2643 859 2647
rect 863 2643 864 2647
rect 858 2642 864 2643
rect 860 2624 862 2642
rect 858 2623 864 2624
rect 858 2619 859 2623
rect 863 2619 864 2623
rect 858 2618 864 2619
rect 908 2608 910 2669
rect 1032 2616 1034 2694
rect 1116 2675 1118 2736
rect 1204 2700 1206 2846
rect 1316 2844 1318 2905
rect 1484 2844 1486 2905
rect 1644 2844 1646 2905
rect 1788 2844 1790 2905
rect 1874 2883 1880 2884
rect 1874 2879 1875 2883
rect 1879 2879 1880 2883
rect 1874 2878 1880 2879
rect 1314 2843 1320 2844
rect 1314 2839 1315 2843
rect 1319 2839 1320 2843
rect 1314 2838 1320 2839
rect 1482 2843 1488 2844
rect 1482 2839 1483 2843
rect 1487 2839 1488 2843
rect 1482 2838 1488 2839
rect 1642 2843 1648 2844
rect 1642 2839 1643 2843
rect 1647 2839 1648 2843
rect 1642 2838 1648 2839
rect 1786 2843 1792 2844
rect 1786 2839 1787 2843
rect 1791 2839 1792 2843
rect 1786 2838 1792 2839
rect 1342 2828 1348 2829
rect 1342 2824 1343 2828
rect 1347 2824 1348 2828
rect 1342 2823 1348 2824
rect 1510 2828 1516 2829
rect 1510 2824 1511 2828
rect 1515 2824 1516 2828
rect 1510 2823 1516 2824
rect 1670 2828 1676 2829
rect 1670 2824 1671 2828
rect 1675 2824 1676 2828
rect 1670 2823 1676 2824
rect 1814 2828 1820 2829
rect 1814 2824 1815 2828
rect 1819 2824 1820 2828
rect 1814 2823 1820 2824
rect 1344 2787 1346 2823
rect 1512 2787 1514 2823
rect 1672 2787 1674 2823
rect 1816 2787 1818 2823
rect 1311 2786 1315 2787
rect 1311 2781 1315 2782
rect 1343 2786 1347 2787
rect 1343 2781 1347 2782
rect 1479 2786 1483 2787
rect 1479 2781 1483 2782
rect 1511 2786 1515 2787
rect 1511 2781 1515 2782
rect 1671 2786 1675 2787
rect 1671 2781 1675 2782
rect 1815 2786 1819 2787
rect 1815 2781 1819 2782
rect 1312 2757 1314 2781
rect 1480 2757 1482 2781
rect 1876 2776 1878 2878
rect 1936 2845 1938 2905
rect 1934 2844 1940 2845
rect 1934 2840 1935 2844
rect 1939 2840 1940 2844
rect 1934 2839 1940 2840
rect 1976 2831 1978 2906
rect 2832 2831 2834 2907
rect 2968 2831 2970 2907
rect 1975 2830 1979 2831
rect 1934 2827 1940 2828
rect 1934 2823 1935 2827
rect 1939 2823 1940 2827
rect 1975 2825 1979 2826
rect 2023 2830 2027 2831
rect 2023 2825 2027 2826
rect 2167 2830 2171 2831
rect 2167 2825 2171 2826
rect 2335 2830 2339 2831
rect 2335 2825 2339 2826
rect 2495 2830 2499 2831
rect 2495 2825 2499 2826
rect 2663 2830 2667 2831
rect 2663 2825 2667 2826
rect 2831 2830 2835 2831
rect 2831 2825 2835 2826
rect 2967 2830 2971 2831
rect 2967 2825 2971 2826
rect 2999 2830 3003 2831
rect 2999 2825 3003 2826
rect 1934 2822 1940 2823
rect 1936 2787 1938 2822
rect 1976 2802 1978 2825
rect 1974 2801 1980 2802
rect 2024 2801 2026 2825
rect 2168 2801 2170 2825
rect 2336 2801 2338 2825
rect 2496 2801 2498 2825
rect 2664 2801 2666 2825
rect 2832 2801 2834 2825
rect 3000 2801 3002 2825
rect 1974 2797 1975 2801
rect 1979 2797 1980 2801
rect 1974 2796 1980 2797
rect 2022 2800 2028 2801
rect 2022 2796 2023 2800
rect 2027 2796 2028 2800
rect 2022 2795 2028 2796
rect 2166 2800 2172 2801
rect 2166 2796 2167 2800
rect 2171 2796 2172 2800
rect 2166 2795 2172 2796
rect 2334 2800 2340 2801
rect 2334 2796 2335 2800
rect 2339 2796 2340 2800
rect 2334 2795 2340 2796
rect 2494 2800 2500 2801
rect 2494 2796 2495 2800
rect 2499 2796 2500 2800
rect 2494 2795 2500 2796
rect 2662 2800 2668 2801
rect 2662 2796 2663 2800
rect 2667 2796 2668 2800
rect 2662 2795 2668 2796
rect 2830 2800 2836 2801
rect 2830 2796 2831 2800
rect 2835 2796 2836 2800
rect 2830 2795 2836 2796
rect 2998 2800 3004 2801
rect 2998 2796 2999 2800
rect 3003 2796 3004 2800
rect 2998 2795 3004 2796
rect 1935 2786 1939 2787
rect 1994 2785 2000 2786
rect 1935 2781 1939 2782
rect 1974 2784 1980 2785
rect 1874 2775 1880 2776
rect 1874 2771 1875 2775
rect 1879 2771 1880 2775
rect 1874 2770 1880 2771
rect 1936 2758 1938 2781
rect 1974 2780 1975 2784
rect 1979 2780 1980 2784
rect 1994 2781 1995 2785
rect 1999 2781 2000 2785
rect 1994 2780 2000 2781
rect 2138 2785 2144 2786
rect 2138 2781 2139 2785
rect 2143 2781 2144 2785
rect 2138 2780 2144 2781
rect 2306 2785 2312 2786
rect 2306 2781 2307 2785
rect 2311 2781 2312 2785
rect 2306 2780 2312 2781
rect 2466 2785 2472 2786
rect 2466 2781 2467 2785
rect 2471 2781 2472 2785
rect 2466 2780 2472 2781
rect 2634 2785 2640 2786
rect 2634 2781 2635 2785
rect 2639 2781 2640 2785
rect 2634 2780 2640 2781
rect 2802 2785 2808 2786
rect 2802 2781 2803 2785
rect 2807 2781 2808 2785
rect 2802 2780 2808 2781
rect 2970 2785 2976 2786
rect 2970 2781 2971 2785
rect 2975 2781 2976 2785
rect 2970 2780 2976 2781
rect 1974 2779 1980 2780
rect 1934 2757 1940 2758
rect 1310 2756 1316 2757
rect 1310 2752 1311 2756
rect 1315 2752 1316 2756
rect 1310 2751 1316 2752
rect 1478 2756 1484 2757
rect 1478 2752 1479 2756
rect 1483 2752 1484 2756
rect 1934 2753 1935 2757
rect 1939 2753 1940 2757
rect 1934 2752 1940 2753
rect 1478 2751 1484 2752
rect 1282 2741 1288 2742
rect 1282 2737 1283 2741
rect 1287 2737 1288 2741
rect 1282 2736 1288 2737
rect 1450 2741 1456 2742
rect 1450 2737 1451 2741
rect 1455 2737 1456 2741
rect 1450 2736 1456 2737
rect 1934 2740 1940 2741
rect 1934 2736 1935 2740
rect 1939 2736 1940 2740
rect 1202 2699 1208 2700
rect 1202 2695 1203 2699
rect 1207 2695 1208 2699
rect 1202 2694 1208 2695
rect 1284 2675 1286 2736
rect 1298 2731 1304 2732
rect 1298 2727 1299 2731
rect 1303 2727 1304 2731
rect 1298 2726 1304 2727
rect 1300 2700 1302 2726
rect 1298 2699 1304 2700
rect 1298 2695 1299 2699
rect 1303 2695 1304 2699
rect 1298 2694 1304 2695
rect 1452 2675 1454 2736
rect 1934 2735 1940 2736
rect 1466 2731 1472 2732
rect 1466 2727 1467 2731
rect 1471 2727 1472 2731
rect 1466 2726 1472 2727
rect 1554 2731 1560 2732
rect 1554 2727 1555 2731
rect 1559 2727 1560 2731
rect 1554 2726 1560 2727
rect 1468 2700 1470 2726
rect 1466 2699 1472 2700
rect 1466 2695 1467 2699
rect 1471 2695 1472 2699
rect 1466 2694 1472 2695
rect 1043 2674 1047 2675
rect 1043 2669 1047 2670
rect 1115 2674 1119 2675
rect 1115 2669 1119 2670
rect 1179 2674 1183 2675
rect 1179 2669 1183 2670
rect 1283 2674 1287 2675
rect 1283 2669 1287 2670
rect 1315 2674 1319 2675
rect 1315 2669 1319 2670
rect 1451 2674 1455 2675
rect 1451 2669 1455 2670
rect 1030 2615 1036 2616
rect 1030 2611 1031 2615
rect 1035 2611 1036 2615
rect 1030 2610 1036 2611
rect 1044 2608 1046 2669
rect 1180 2608 1182 2669
rect 1316 2608 1318 2669
rect 1402 2647 1408 2648
rect 1402 2643 1403 2647
rect 1407 2643 1408 2647
rect 1402 2642 1408 2643
rect 110 2604 111 2608
rect 115 2604 116 2608
rect 110 2603 116 2604
rect 770 2607 776 2608
rect 770 2603 771 2607
rect 775 2603 776 2607
rect 770 2602 776 2603
rect 906 2607 912 2608
rect 906 2603 907 2607
rect 911 2603 912 2607
rect 906 2602 912 2603
rect 1042 2607 1048 2608
rect 1042 2603 1043 2607
rect 1047 2603 1048 2607
rect 1042 2602 1048 2603
rect 1178 2607 1184 2608
rect 1178 2603 1179 2607
rect 1183 2603 1184 2607
rect 1178 2602 1184 2603
rect 1314 2607 1320 2608
rect 1314 2603 1315 2607
rect 1319 2603 1320 2607
rect 1314 2602 1320 2603
rect 798 2592 804 2593
rect 110 2591 116 2592
rect 110 2587 111 2591
rect 115 2587 116 2591
rect 798 2588 799 2592
rect 803 2588 804 2592
rect 798 2587 804 2588
rect 934 2592 940 2593
rect 934 2588 935 2592
rect 939 2588 940 2592
rect 934 2587 940 2588
rect 1070 2592 1076 2593
rect 1070 2588 1071 2592
rect 1075 2588 1076 2592
rect 1070 2587 1076 2588
rect 1206 2592 1212 2593
rect 1206 2588 1207 2592
rect 1211 2588 1212 2592
rect 1206 2587 1212 2588
rect 1342 2592 1348 2593
rect 1342 2588 1343 2592
rect 1347 2588 1348 2592
rect 1342 2587 1348 2588
rect 110 2586 116 2587
rect 112 2547 114 2586
rect 800 2547 802 2587
rect 936 2547 938 2587
rect 1072 2547 1074 2587
rect 1208 2547 1210 2587
rect 1344 2547 1346 2587
rect 111 2546 115 2547
rect 111 2541 115 2542
rect 551 2546 555 2547
rect 551 2541 555 2542
rect 687 2546 691 2547
rect 687 2541 691 2542
rect 799 2546 803 2547
rect 799 2541 803 2542
rect 831 2546 835 2547
rect 831 2541 835 2542
rect 935 2546 939 2547
rect 935 2541 939 2542
rect 983 2546 987 2547
rect 983 2541 987 2542
rect 1071 2546 1075 2547
rect 1071 2541 1075 2542
rect 1135 2546 1139 2547
rect 1135 2541 1139 2542
rect 1207 2546 1211 2547
rect 1207 2541 1211 2542
rect 1295 2546 1299 2547
rect 1295 2541 1299 2542
rect 1343 2546 1347 2547
rect 1343 2541 1347 2542
rect 112 2518 114 2541
rect 110 2517 116 2518
rect 552 2517 554 2541
rect 688 2517 690 2541
rect 832 2517 834 2541
rect 984 2517 986 2541
rect 1136 2517 1138 2541
rect 1296 2517 1298 2541
rect 110 2513 111 2517
rect 115 2513 116 2517
rect 110 2512 116 2513
rect 550 2516 556 2517
rect 550 2512 551 2516
rect 555 2512 556 2516
rect 550 2511 556 2512
rect 686 2516 692 2517
rect 686 2512 687 2516
rect 691 2512 692 2516
rect 686 2511 692 2512
rect 830 2516 836 2517
rect 830 2512 831 2516
rect 835 2512 836 2516
rect 830 2511 836 2512
rect 982 2516 988 2517
rect 982 2512 983 2516
rect 987 2512 988 2516
rect 982 2511 988 2512
rect 1134 2516 1140 2517
rect 1134 2512 1135 2516
rect 1139 2512 1140 2516
rect 1134 2511 1140 2512
rect 1294 2516 1300 2517
rect 1294 2512 1295 2516
rect 1299 2512 1300 2516
rect 1294 2511 1300 2512
rect 522 2501 528 2502
rect 110 2500 116 2501
rect 110 2496 111 2500
rect 115 2496 116 2500
rect 522 2497 523 2501
rect 527 2497 528 2501
rect 522 2496 528 2497
rect 658 2501 664 2502
rect 658 2497 659 2501
rect 663 2497 664 2501
rect 658 2496 664 2497
rect 802 2501 808 2502
rect 802 2497 803 2501
rect 807 2497 808 2501
rect 802 2496 808 2497
rect 954 2501 960 2502
rect 954 2497 955 2501
rect 959 2497 960 2501
rect 954 2496 960 2497
rect 1106 2501 1112 2502
rect 1106 2497 1107 2501
rect 1111 2497 1112 2501
rect 1106 2496 1112 2497
rect 1266 2501 1272 2502
rect 1266 2497 1267 2501
rect 1271 2497 1272 2501
rect 1266 2496 1272 2497
rect 110 2495 116 2496
rect 112 2423 114 2495
rect 524 2423 526 2496
rect 660 2423 662 2496
rect 674 2491 680 2492
rect 674 2487 675 2491
rect 679 2487 680 2491
rect 674 2486 680 2487
rect 676 2460 678 2486
rect 666 2459 672 2460
rect 666 2455 667 2459
rect 671 2455 672 2459
rect 666 2454 672 2455
rect 674 2459 680 2460
rect 674 2455 675 2459
rect 679 2455 680 2459
rect 674 2454 680 2455
rect 111 2422 115 2423
rect 111 2417 115 2418
rect 131 2422 135 2423
rect 131 2417 135 2418
rect 339 2422 343 2423
rect 339 2417 343 2418
rect 523 2422 527 2423
rect 523 2417 527 2418
rect 563 2422 567 2423
rect 563 2417 567 2418
rect 659 2422 663 2423
rect 659 2417 663 2418
rect 112 2357 114 2417
rect 110 2356 116 2357
rect 132 2356 134 2417
rect 306 2399 312 2400
rect 218 2395 224 2396
rect 218 2391 219 2395
rect 223 2391 224 2395
rect 306 2395 307 2399
rect 311 2395 312 2399
rect 306 2394 312 2395
rect 218 2390 224 2391
rect 110 2352 111 2356
rect 115 2352 116 2356
rect 110 2351 116 2352
rect 130 2355 136 2356
rect 130 2351 131 2355
rect 135 2351 136 2355
rect 130 2350 136 2351
rect 158 2340 164 2341
rect 110 2339 116 2340
rect 110 2335 111 2339
rect 115 2335 116 2339
rect 158 2336 159 2340
rect 163 2336 164 2340
rect 158 2335 164 2336
rect 110 2334 116 2335
rect 112 2307 114 2334
rect 160 2307 162 2335
rect 111 2306 115 2307
rect 111 2301 115 2302
rect 159 2306 163 2307
rect 159 2301 163 2302
rect 112 2278 114 2301
rect 110 2277 116 2278
rect 160 2277 162 2301
rect 110 2273 111 2277
rect 115 2273 116 2277
rect 110 2272 116 2273
rect 158 2276 164 2277
rect 158 2272 159 2276
rect 163 2272 164 2276
rect 158 2271 164 2272
rect 130 2261 136 2262
rect 110 2260 116 2261
rect 110 2256 111 2260
rect 115 2256 116 2260
rect 130 2257 131 2261
rect 135 2257 136 2261
rect 130 2256 136 2257
rect 110 2255 116 2256
rect 112 2171 114 2255
rect 132 2171 134 2256
rect 220 2244 222 2390
rect 308 2364 310 2394
rect 306 2363 312 2364
rect 306 2359 307 2363
rect 311 2359 312 2363
rect 306 2358 312 2359
rect 340 2356 342 2417
rect 466 2399 472 2400
rect 466 2395 467 2399
rect 471 2395 472 2399
rect 466 2394 472 2395
rect 468 2364 470 2394
rect 466 2363 472 2364
rect 466 2359 467 2363
rect 471 2359 472 2363
rect 466 2358 472 2359
rect 564 2356 566 2417
rect 668 2372 670 2454
rect 804 2423 806 2496
rect 818 2491 824 2492
rect 818 2487 819 2491
rect 823 2487 824 2491
rect 818 2486 824 2487
rect 820 2460 822 2486
rect 818 2459 824 2460
rect 818 2455 819 2459
rect 823 2455 824 2459
rect 818 2454 824 2455
rect 956 2423 958 2496
rect 970 2491 976 2492
rect 970 2487 971 2491
rect 975 2487 976 2491
rect 970 2486 976 2487
rect 972 2460 974 2486
rect 970 2459 976 2460
rect 970 2455 971 2459
rect 975 2455 976 2459
rect 970 2454 976 2455
rect 1108 2423 1110 2496
rect 1122 2491 1128 2492
rect 1122 2487 1123 2491
rect 1127 2487 1128 2491
rect 1122 2486 1128 2487
rect 1124 2460 1126 2486
rect 1122 2459 1128 2460
rect 1122 2455 1123 2459
rect 1127 2455 1128 2459
rect 1122 2454 1128 2455
rect 1268 2423 1270 2496
rect 1404 2492 1406 2642
rect 1452 2608 1454 2669
rect 1556 2652 1558 2726
rect 1936 2675 1938 2735
rect 1976 2719 1978 2779
rect 1996 2719 1998 2780
rect 2140 2719 2142 2780
rect 2308 2719 2310 2780
rect 2468 2719 2470 2780
rect 2502 2743 2508 2744
rect 2502 2739 2503 2743
rect 2507 2739 2508 2743
rect 2502 2738 2508 2739
rect 1975 2718 1979 2719
rect 1975 2713 1979 2714
rect 1995 2718 1999 2719
rect 1995 2713 1999 2714
rect 2139 2718 2143 2719
rect 2139 2713 2143 2714
rect 2307 2718 2311 2719
rect 2307 2713 2311 2714
rect 2379 2718 2383 2719
rect 2379 2713 2383 2714
rect 2467 2718 2471 2719
rect 2467 2713 2471 2714
rect 1587 2674 1591 2675
rect 1587 2669 1591 2670
rect 1723 2674 1727 2675
rect 1723 2669 1727 2670
rect 1935 2674 1939 2675
rect 1935 2669 1939 2670
rect 1554 2651 1560 2652
rect 1554 2647 1555 2651
rect 1559 2647 1560 2651
rect 1554 2646 1560 2647
rect 1588 2608 1590 2669
rect 1724 2608 1726 2669
rect 1842 2615 1848 2616
rect 1842 2611 1843 2615
rect 1847 2611 1848 2615
rect 1842 2610 1848 2611
rect 1450 2607 1456 2608
rect 1450 2603 1451 2607
rect 1455 2603 1456 2607
rect 1450 2602 1456 2603
rect 1586 2607 1592 2608
rect 1586 2603 1587 2607
rect 1591 2603 1592 2607
rect 1586 2602 1592 2603
rect 1722 2607 1728 2608
rect 1722 2603 1723 2607
rect 1727 2603 1728 2607
rect 1722 2602 1728 2603
rect 1478 2592 1484 2593
rect 1478 2588 1479 2592
rect 1483 2588 1484 2592
rect 1478 2587 1484 2588
rect 1614 2592 1620 2593
rect 1614 2588 1615 2592
rect 1619 2588 1620 2592
rect 1614 2587 1620 2588
rect 1750 2592 1756 2593
rect 1750 2588 1751 2592
rect 1755 2588 1756 2592
rect 1750 2587 1756 2588
rect 1480 2547 1482 2587
rect 1616 2547 1618 2587
rect 1752 2547 1754 2587
rect 1455 2546 1459 2547
rect 1455 2541 1459 2542
rect 1479 2546 1483 2547
rect 1479 2541 1483 2542
rect 1615 2546 1619 2547
rect 1615 2541 1619 2542
rect 1751 2546 1755 2547
rect 1751 2541 1755 2542
rect 1783 2546 1787 2547
rect 1783 2541 1787 2542
rect 1456 2517 1458 2541
rect 1616 2517 1618 2541
rect 1784 2517 1786 2541
rect 1454 2516 1460 2517
rect 1454 2512 1455 2516
rect 1459 2512 1460 2516
rect 1454 2511 1460 2512
rect 1614 2516 1620 2517
rect 1614 2512 1615 2516
rect 1619 2512 1620 2516
rect 1614 2511 1620 2512
rect 1782 2516 1788 2517
rect 1782 2512 1783 2516
rect 1787 2512 1788 2516
rect 1782 2511 1788 2512
rect 1426 2501 1432 2502
rect 1426 2497 1427 2501
rect 1431 2497 1432 2501
rect 1426 2496 1432 2497
rect 1586 2501 1592 2502
rect 1586 2497 1587 2501
rect 1591 2497 1592 2501
rect 1586 2496 1592 2497
rect 1754 2501 1760 2502
rect 1754 2497 1755 2501
rect 1759 2497 1760 2501
rect 1754 2496 1760 2497
rect 1282 2491 1288 2492
rect 1282 2487 1283 2491
rect 1287 2487 1288 2491
rect 1282 2486 1288 2487
rect 1402 2491 1408 2492
rect 1402 2487 1403 2491
rect 1407 2487 1408 2491
rect 1402 2486 1408 2487
rect 1410 2491 1416 2492
rect 1410 2487 1411 2491
rect 1415 2487 1416 2491
rect 1410 2486 1416 2487
rect 1284 2460 1286 2486
rect 1282 2459 1288 2460
rect 1282 2455 1283 2459
rect 1287 2455 1288 2459
rect 1282 2454 1288 2455
rect 803 2422 807 2423
rect 803 2417 807 2418
rect 955 2422 959 2423
rect 955 2417 959 2418
rect 1043 2422 1047 2423
rect 1043 2417 1047 2418
rect 1107 2422 1111 2423
rect 1107 2417 1111 2418
rect 1267 2422 1271 2423
rect 1267 2417 1271 2418
rect 1291 2422 1295 2423
rect 1291 2417 1295 2418
rect 690 2399 696 2400
rect 690 2395 691 2399
rect 695 2395 696 2399
rect 690 2394 696 2395
rect 666 2371 672 2372
rect 666 2367 667 2371
rect 671 2367 672 2371
rect 666 2366 672 2367
rect 692 2364 694 2394
rect 690 2363 696 2364
rect 690 2359 691 2363
rect 695 2359 696 2363
rect 690 2358 696 2359
rect 804 2356 806 2417
rect 930 2399 936 2400
rect 930 2395 931 2399
rect 935 2395 936 2399
rect 930 2394 936 2395
rect 932 2364 934 2394
rect 930 2363 936 2364
rect 930 2359 931 2363
rect 935 2359 936 2363
rect 930 2358 936 2359
rect 1044 2356 1046 2417
rect 1292 2356 1294 2417
rect 1412 2400 1414 2486
rect 1428 2423 1430 2496
rect 1588 2423 1590 2496
rect 1742 2491 1748 2492
rect 1742 2487 1743 2491
rect 1747 2487 1748 2491
rect 1742 2486 1748 2487
rect 1744 2460 1746 2486
rect 1742 2459 1748 2460
rect 1742 2455 1743 2459
rect 1747 2455 1748 2459
rect 1742 2454 1748 2455
rect 1756 2423 1758 2496
rect 1844 2460 1846 2610
rect 1936 2609 1938 2669
rect 1976 2653 1978 2713
rect 1974 2652 1980 2653
rect 2380 2652 2382 2713
rect 2504 2660 2506 2738
rect 2636 2719 2638 2780
rect 2746 2775 2752 2776
rect 2746 2771 2747 2775
rect 2751 2771 2752 2775
rect 2746 2770 2752 2771
rect 2790 2775 2796 2776
rect 2790 2771 2791 2775
rect 2795 2771 2796 2775
rect 2790 2770 2796 2771
rect 2515 2718 2519 2719
rect 2515 2713 2519 2714
rect 2635 2718 2639 2719
rect 2635 2713 2639 2714
rect 2659 2718 2663 2719
rect 2659 2713 2663 2714
rect 2502 2659 2508 2660
rect 2502 2655 2503 2659
rect 2507 2655 2508 2659
rect 2502 2654 2508 2655
rect 2516 2652 2518 2713
rect 2602 2691 2608 2692
rect 2602 2687 2603 2691
rect 2607 2687 2608 2691
rect 2602 2686 2608 2687
rect 1974 2648 1975 2652
rect 1979 2648 1980 2652
rect 1974 2647 1980 2648
rect 2378 2651 2384 2652
rect 2378 2647 2379 2651
rect 2383 2647 2384 2651
rect 2378 2646 2384 2647
rect 2514 2651 2520 2652
rect 2514 2647 2515 2651
rect 2519 2647 2520 2651
rect 2514 2646 2520 2647
rect 2406 2636 2412 2637
rect 1974 2635 1980 2636
rect 1974 2631 1975 2635
rect 1979 2631 1980 2635
rect 2406 2632 2407 2636
rect 2411 2632 2412 2636
rect 2406 2631 2412 2632
rect 2542 2636 2548 2637
rect 2542 2632 2543 2636
rect 2547 2632 2548 2636
rect 2542 2631 2548 2632
rect 1974 2630 1980 2631
rect 1934 2608 1940 2609
rect 1934 2604 1935 2608
rect 1939 2604 1940 2608
rect 1934 2603 1940 2604
rect 1976 2603 1978 2630
rect 2408 2603 2410 2631
rect 2544 2603 2546 2631
rect 1975 2602 1979 2603
rect 1975 2597 1979 2598
rect 2407 2602 2411 2603
rect 2407 2597 2411 2598
rect 2511 2602 2515 2603
rect 2511 2597 2515 2598
rect 2543 2602 2547 2603
rect 2543 2597 2547 2598
rect 1934 2591 1940 2592
rect 1934 2587 1935 2591
rect 1939 2587 1940 2591
rect 1934 2586 1940 2587
rect 1936 2547 1938 2586
rect 1976 2574 1978 2597
rect 1974 2573 1980 2574
rect 2512 2573 2514 2597
rect 1974 2569 1975 2573
rect 1979 2569 1980 2573
rect 1974 2568 1980 2569
rect 2510 2572 2516 2573
rect 2510 2568 2511 2572
rect 2515 2568 2516 2572
rect 2510 2567 2516 2568
rect 2482 2557 2488 2558
rect 1974 2556 1980 2557
rect 1974 2552 1975 2556
rect 1979 2552 1980 2556
rect 2482 2553 2483 2557
rect 2487 2553 2488 2557
rect 2482 2552 2488 2553
rect 1974 2551 1980 2552
rect 1935 2546 1939 2547
rect 1935 2541 1939 2542
rect 1936 2518 1938 2541
rect 1934 2517 1940 2518
rect 1934 2513 1935 2517
rect 1939 2513 1940 2517
rect 1934 2512 1940 2513
rect 1934 2500 1940 2501
rect 1934 2496 1935 2500
rect 1939 2496 1940 2500
rect 1934 2495 1940 2496
rect 1842 2459 1848 2460
rect 1842 2455 1843 2459
rect 1847 2455 1848 2459
rect 1842 2454 1848 2455
rect 1936 2423 1938 2495
rect 1976 2475 1978 2551
rect 2484 2475 2486 2552
rect 2604 2548 2606 2686
rect 2660 2652 2662 2713
rect 2748 2692 2750 2770
rect 2792 2744 2794 2770
rect 2790 2743 2796 2744
rect 2790 2739 2791 2743
rect 2795 2739 2796 2743
rect 2790 2738 2796 2739
rect 2804 2719 2806 2780
rect 2890 2767 2896 2768
rect 2890 2763 2891 2767
rect 2895 2763 2896 2767
rect 2890 2762 2896 2763
rect 2892 2744 2894 2762
rect 2890 2743 2896 2744
rect 2890 2739 2891 2743
rect 2895 2739 2896 2743
rect 2890 2738 2896 2739
rect 2972 2719 2974 2780
rect 3060 2744 3062 2930
rect 3076 2928 3078 2989
rect 3212 2928 3214 2989
rect 3348 2928 3350 2989
rect 3484 2928 3486 2989
rect 3608 2936 3610 3014
rect 3800 2995 3802 3055
rect 3839 3053 3843 3054
rect 4255 3058 4259 3059
rect 4255 3053 4259 3054
rect 4455 3058 4459 3059
rect 4455 3053 4459 3054
rect 4495 3058 4499 3059
rect 4495 3053 4499 3054
rect 3840 3030 3842 3053
rect 3838 3029 3844 3030
rect 4256 3029 4258 3053
rect 4358 3043 4364 3044
rect 4358 3039 4359 3043
rect 4363 3039 4364 3043
rect 4358 3038 4364 3039
rect 3838 3025 3839 3029
rect 3843 3025 3844 3029
rect 3838 3024 3844 3025
rect 4254 3028 4260 3029
rect 4254 3024 4255 3028
rect 4259 3024 4260 3028
rect 4254 3023 4260 3024
rect 4226 3013 4232 3014
rect 3838 3012 3844 3013
rect 3838 3008 3839 3012
rect 3843 3008 3844 3012
rect 4226 3009 4227 3013
rect 4231 3009 4232 3013
rect 4226 3008 4232 3009
rect 3838 3007 3844 3008
rect 3799 2994 3803 2995
rect 3799 2989 3803 2990
rect 3606 2935 3612 2936
rect 3606 2931 3607 2935
rect 3611 2931 3612 2935
rect 3606 2930 3612 2931
rect 3800 2929 3802 2989
rect 3798 2928 3804 2929
rect 3074 2927 3080 2928
rect 3074 2923 3075 2927
rect 3079 2923 3080 2927
rect 3074 2922 3080 2923
rect 3210 2927 3216 2928
rect 3210 2923 3211 2927
rect 3215 2923 3216 2927
rect 3210 2922 3216 2923
rect 3346 2927 3352 2928
rect 3346 2923 3347 2927
rect 3351 2923 3352 2927
rect 3346 2922 3352 2923
rect 3482 2927 3488 2928
rect 3482 2923 3483 2927
rect 3487 2923 3488 2927
rect 3798 2924 3799 2928
rect 3803 2924 3804 2928
rect 3798 2923 3804 2924
rect 3840 2923 3842 3007
rect 4228 2923 4230 3008
rect 4360 2972 4362 3038
rect 4456 3029 4458 3053
rect 4454 3028 4460 3029
rect 4454 3024 4455 3028
rect 4459 3024 4460 3028
rect 4454 3023 4460 3024
rect 4426 3013 4432 3014
rect 4426 3009 4427 3013
rect 4431 3009 4432 3013
rect 4426 3008 4432 3009
rect 4642 3013 4648 3014
rect 4642 3009 4643 3013
rect 4647 3009 4648 3013
rect 4642 3008 4648 3009
rect 4358 2971 4364 2972
rect 4358 2967 4359 2971
rect 4363 2967 4364 2971
rect 4358 2966 4364 2967
rect 4428 2923 4430 3008
rect 4442 3003 4448 3004
rect 4442 2999 4443 3003
rect 4447 2999 4448 3003
rect 4442 2998 4448 2999
rect 4546 3003 4552 3004
rect 4546 2999 4547 3003
rect 4551 2999 4552 3003
rect 4546 2998 4552 2999
rect 4444 2972 4446 2998
rect 4442 2971 4448 2972
rect 4442 2967 4443 2971
rect 4447 2967 4448 2971
rect 4442 2966 4448 2967
rect 3482 2922 3488 2923
rect 3839 2922 3843 2923
rect 3839 2917 3843 2918
rect 3995 2922 3999 2923
rect 3995 2917 3999 2918
rect 4211 2922 4215 2923
rect 4211 2917 4215 2918
rect 4227 2922 4231 2923
rect 4227 2917 4231 2918
rect 4427 2922 4431 2923
rect 4427 2917 4431 2918
rect 4443 2922 4447 2923
rect 4443 2917 4447 2918
rect 3102 2912 3108 2913
rect 3102 2908 3103 2912
rect 3107 2908 3108 2912
rect 3102 2907 3108 2908
rect 3238 2912 3244 2913
rect 3238 2908 3239 2912
rect 3243 2908 3244 2912
rect 3238 2907 3244 2908
rect 3374 2912 3380 2913
rect 3374 2908 3375 2912
rect 3379 2908 3380 2912
rect 3374 2907 3380 2908
rect 3510 2912 3516 2913
rect 3510 2908 3511 2912
rect 3515 2908 3516 2912
rect 3510 2907 3516 2908
rect 3798 2911 3804 2912
rect 3798 2907 3799 2911
rect 3803 2907 3804 2911
rect 3104 2831 3106 2907
rect 3240 2831 3242 2907
rect 3376 2831 3378 2907
rect 3512 2831 3514 2907
rect 3798 2906 3804 2907
rect 3800 2831 3802 2906
rect 3840 2857 3842 2917
rect 3978 2863 3984 2864
rect 3978 2859 3979 2863
rect 3983 2859 3984 2863
rect 3978 2858 3984 2859
rect 3838 2856 3844 2857
rect 3838 2852 3839 2856
rect 3843 2852 3844 2856
rect 3838 2851 3844 2852
rect 3838 2839 3844 2840
rect 3838 2835 3839 2839
rect 3843 2835 3844 2839
rect 3838 2834 3844 2835
rect 3103 2830 3107 2831
rect 3103 2825 3107 2826
rect 3167 2830 3171 2831
rect 3167 2825 3171 2826
rect 3239 2830 3243 2831
rect 3239 2825 3243 2826
rect 3375 2830 3379 2831
rect 3375 2825 3379 2826
rect 3511 2830 3515 2831
rect 3511 2825 3515 2826
rect 3799 2830 3803 2831
rect 3799 2825 3803 2826
rect 3168 2801 3170 2825
rect 3800 2802 3802 2825
rect 3840 2807 3842 2834
rect 3839 2806 3843 2807
rect 3798 2801 3804 2802
rect 3839 2801 3843 2802
rect 3919 2806 3923 2807
rect 3919 2801 3923 2802
rect 3166 2800 3172 2801
rect 3166 2796 3167 2800
rect 3171 2796 3172 2800
rect 3798 2797 3799 2801
rect 3803 2797 3804 2801
rect 3798 2796 3804 2797
rect 3166 2795 3172 2796
rect 3138 2785 3144 2786
rect 3138 2781 3139 2785
rect 3143 2781 3144 2785
rect 3138 2780 3144 2781
rect 3798 2784 3804 2785
rect 3798 2780 3799 2784
rect 3803 2780 3804 2784
rect 3058 2743 3064 2744
rect 3058 2739 3059 2743
rect 3063 2739 3064 2743
rect 3058 2738 3064 2739
rect 3140 2719 3142 2780
rect 3798 2779 3804 2780
rect 3154 2775 3160 2776
rect 3154 2771 3155 2775
rect 3159 2771 3160 2775
rect 3154 2770 3160 2771
rect 3156 2744 3158 2770
rect 3154 2743 3160 2744
rect 3154 2739 3155 2743
rect 3159 2739 3160 2743
rect 3154 2738 3160 2739
rect 3800 2719 3802 2779
rect 3840 2778 3842 2801
rect 3838 2777 3844 2778
rect 3920 2777 3922 2801
rect 3838 2773 3839 2777
rect 3843 2773 3844 2777
rect 3838 2772 3844 2773
rect 3918 2776 3924 2777
rect 3918 2772 3919 2776
rect 3923 2772 3924 2776
rect 3918 2771 3924 2772
rect 3890 2761 3896 2762
rect 3838 2760 3844 2761
rect 3838 2756 3839 2760
rect 3843 2756 3844 2760
rect 3890 2757 3891 2761
rect 3895 2757 3896 2761
rect 3890 2756 3896 2757
rect 3838 2755 3844 2756
rect 2803 2718 2807 2719
rect 2803 2713 2807 2714
rect 2947 2718 2951 2719
rect 2947 2713 2951 2714
rect 2971 2718 2975 2719
rect 2971 2713 2975 2714
rect 3091 2718 3095 2719
rect 3091 2713 3095 2714
rect 3139 2718 3143 2719
rect 3139 2713 3143 2714
rect 3235 2718 3239 2719
rect 3235 2713 3239 2714
rect 3799 2718 3803 2719
rect 3799 2713 3803 2714
rect 2786 2695 2792 2696
rect 2746 2691 2752 2692
rect 2746 2687 2747 2691
rect 2751 2687 2752 2691
rect 2786 2691 2787 2695
rect 2791 2691 2792 2695
rect 2786 2690 2792 2691
rect 2746 2686 2752 2687
rect 2788 2660 2790 2690
rect 2786 2659 2792 2660
rect 2786 2655 2787 2659
rect 2791 2655 2792 2659
rect 2786 2654 2792 2655
rect 2804 2652 2806 2713
rect 2930 2695 2936 2696
rect 2930 2691 2931 2695
rect 2935 2691 2936 2695
rect 2930 2690 2936 2691
rect 2932 2660 2934 2690
rect 2930 2659 2936 2660
rect 2930 2655 2931 2659
rect 2935 2655 2936 2659
rect 2930 2654 2936 2655
rect 2948 2652 2950 2713
rect 3074 2695 3080 2696
rect 3074 2691 3075 2695
rect 3079 2691 3080 2695
rect 3074 2690 3080 2691
rect 3076 2660 3078 2690
rect 3074 2659 3080 2660
rect 3074 2655 3075 2659
rect 3079 2655 3080 2659
rect 3074 2654 3080 2655
rect 3092 2652 3094 2713
rect 3218 2695 3224 2696
rect 3218 2691 3219 2695
rect 3223 2691 3224 2695
rect 3218 2690 3224 2691
rect 3220 2660 3222 2690
rect 3218 2659 3224 2660
rect 3218 2655 3219 2659
rect 3223 2655 3224 2659
rect 3218 2654 3224 2655
rect 3236 2652 3238 2713
rect 3270 2659 3276 2660
rect 3270 2655 3271 2659
rect 3275 2655 3276 2659
rect 3270 2654 3276 2655
rect 2658 2651 2664 2652
rect 2658 2647 2659 2651
rect 2663 2647 2664 2651
rect 2658 2646 2664 2647
rect 2802 2651 2808 2652
rect 2802 2647 2803 2651
rect 2807 2647 2808 2651
rect 2802 2646 2808 2647
rect 2946 2651 2952 2652
rect 2946 2647 2947 2651
rect 2951 2647 2952 2651
rect 2946 2646 2952 2647
rect 3090 2651 3096 2652
rect 3090 2647 3091 2651
rect 3095 2647 3096 2651
rect 3090 2646 3096 2647
rect 3234 2651 3240 2652
rect 3234 2647 3235 2651
rect 3239 2647 3240 2651
rect 3234 2646 3240 2647
rect 2686 2636 2692 2637
rect 2686 2632 2687 2636
rect 2691 2632 2692 2636
rect 2686 2631 2692 2632
rect 2830 2636 2836 2637
rect 2830 2632 2831 2636
rect 2835 2632 2836 2636
rect 2830 2631 2836 2632
rect 2974 2636 2980 2637
rect 2974 2632 2975 2636
rect 2979 2632 2980 2636
rect 2974 2631 2980 2632
rect 3118 2636 3124 2637
rect 3118 2632 3119 2636
rect 3123 2632 3124 2636
rect 3118 2631 3124 2632
rect 3262 2636 3268 2637
rect 3262 2632 3263 2636
rect 3267 2632 3268 2636
rect 3262 2631 3268 2632
rect 2688 2603 2690 2631
rect 2832 2603 2834 2631
rect 2976 2603 2978 2631
rect 3120 2603 3122 2631
rect 3264 2603 3266 2631
rect 2647 2602 2651 2603
rect 2647 2597 2651 2598
rect 2687 2602 2691 2603
rect 2687 2597 2691 2598
rect 2783 2602 2787 2603
rect 2783 2597 2787 2598
rect 2831 2602 2835 2603
rect 2831 2597 2835 2598
rect 2919 2602 2923 2603
rect 2919 2597 2923 2598
rect 2975 2602 2979 2603
rect 2975 2597 2979 2598
rect 3055 2602 3059 2603
rect 3055 2597 3059 2598
rect 3119 2602 3123 2603
rect 3119 2597 3123 2598
rect 3191 2602 3195 2603
rect 3191 2597 3195 2598
rect 3263 2602 3267 2603
rect 3263 2597 3267 2598
rect 2648 2573 2650 2597
rect 2784 2573 2786 2597
rect 2920 2573 2922 2597
rect 3056 2573 3058 2597
rect 3192 2573 3194 2597
rect 2646 2572 2652 2573
rect 2646 2568 2647 2572
rect 2651 2568 2652 2572
rect 2646 2567 2652 2568
rect 2782 2572 2788 2573
rect 2782 2568 2783 2572
rect 2787 2568 2788 2572
rect 2782 2567 2788 2568
rect 2918 2572 2924 2573
rect 2918 2568 2919 2572
rect 2923 2568 2924 2572
rect 2918 2567 2924 2568
rect 3054 2572 3060 2573
rect 3054 2568 3055 2572
rect 3059 2568 3060 2572
rect 3054 2567 3060 2568
rect 3190 2572 3196 2573
rect 3190 2568 3191 2572
rect 3195 2568 3196 2572
rect 3190 2567 3196 2568
rect 2618 2557 2624 2558
rect 2618 2553 2619 2557
rect 2623 2553 2624 2557
rect 2618 2552 2624 2553
rect 2754 2557 2760 2558
rect 2754 2553 2755 2557
rect 2759 2553 2760 2557
rect 2754 2552 2760 2553
rect 2890 2557 2896 2558
rect 2890 2553 2891 2557
rect 2895 2553 2896 2557
rect 2890 2552 2896 2553
rect 3026 2557 3032 2558
rect 3026 2553 3027 2557
rect 3031 2553 3032 2557
rect 3026 2552 3032 2553
rect 3162 2557 3168 2558
rect 3162 2553 3163 2557
rect 3167 2553 3168 2557
rect 3162 2552 3168 2553
rect 2602 2547 2608 2548
rect 2602 2543 2603 2547
rect 2607 2543 2608 2547
rect 2602 2542 2608 2543
rect 2620 2475 2622 2552
rect 2756 2475 2758 2552
rect 2838 2515 2844 2516
rect 2838 2511 2839 2515
rect 2843 2511 2844 2515
rect 2838 2510 2844 2511
rect 1975 2474 1979 2475
rect 1975 2469 1979 2470
rect 2307 2474 2311 2475
rect 2307 2469 2311 2470
rect 2483 2474 2487 2475
rect 2483 2469 2487 2470
rect 2515 2474 2519 2475
rect 2515 2469 2519 2470
rect 2619 2474 2623 2475
rect 2619 2469 2623 2470
rect 2715 2474 2719 2475
rect 2715 2469 2719 2470
rect 2755 2474 2759 2475
rect 2755 2469 2759 2470
rect 1427 2422 1431 2423
rect 1427 2417 1431 2418
rect 1547 2422 1551 2423
rect 1547 2417 1551 2418
rect 1587 2422 1591 2423
rect 1587 2417 1591 2418
rect 1755 2422 1759 2423
rect 1755 2417 1759 2418
rect 1787 2422 1791 2423
rect 1787 2417 1791 2418
rect 1935 2422 1939 2423
rect 1935 2417 1939 2418
rect 1410 2399 1416 2400
rect 1410 2395 1411 2399
rect 1415 2395 1416 2399
rect 1410 2394 1416 2395
rect 1438 2399 1444 2400
rect 1438 2395 1439 2399
rect 1443 2395 1444 2399
rect 1438 2394 1444 2395
rect 1440 2364 1442 2394
rect 1438 2363 1444 2364
rect 1438 2359 1439 2363
rect 1443 2359 1444 2363
rect 1438 2358 1444 2359
rect 1548 2356 1550 2417
rect 1674 2399 1680 2400
rect 1674 2395 1675 2399
rect 1679 2395 1680 2399
rect 1674 2394 1680 2395
rect 1676 2364 1678 2394
rect 1674 2363 1680 2364
rect 1674 2359 1675 2363
rect 1679 2359 1680 2363
rect 1674 2358 1680 2359
rect 1788 2356 1790 2417
rect 1874 2363 1880 2364
rect 1874 2359 1875 2363
rect 1879 2359 1880 2363
rect 1874 2358 1880 2359
rect 338 2355 344 2356
rect 338 2351 339 2355
rect 343 2351 344 2355
rect 338 2350 344 2351
rect 562 2355 568 2356
rect 562 2351 563 2355
rect 567 2351 568 2355
rect 562 2350 568 2351
rect 802 2355 808 2356
rect 802 2351 803 2355
rect 807 2351 808 2355
rect 802 2350 808 2351
rect 1042 2355 1048 2356
rect 1042 2351 1043 2355
rect 1047 2351 1048 2355
rect 1042 2350 1048 2351
rect 1290 2355 1296 2356
rect 1290 2351 1291 2355
rect 1295 2351 1296 2355
rect 1290 2350 1296 2351
rect 1546 2355 1552 2356
rect 1546 2351 1547 2355
rect 1551 2351 1552 2355
rect 1546 2350 1552 2351
rect 1786 2355 1792 2356
rect 1786 2351 1787 2355
rect 1791 2351 1792 2355
rect 1786 2350 1792 2351
rect 366 2340 372 2341
rect 366 2336 367 2340
rect 371 2336 372 2340
rect 366 2335 372 2336
rect 590 2340 596 2341
rect 590 2336 591 2340
rect 595 2336 596 2340
rect 590 2335 596 2336
rect 830 2340 836 2341
rect 830 2336 831 2340
rect 835 2336 836 2340
rect 830 2335 836 2336
rect 1070 2340 1076 2341
rect 1070 2336 1071 2340
rect 1075 2336 1076 2340
rect 1070 2335 1076 2336
rect 1318 2340 1324 2341
rect 1318 2336 1319 2340
rect 1323 2336 1324 2340
rect 1318 2335 1324 2336
rect 1574 2340 1580 2341
rect 1574 2336 1575 2340
rect 1579 2336 1580 2340
rect 1574 2335 1580 2336
rect 1814 2340 1820 2341
rect 1814 2336 1815 2340
rect 1819 2336 1820 2340
rect 1814 2335 1820 2336
rect 368 2307 370 2335
rect 592 2307 594 2335
rect 832 2307 834 2335
rect 1072 2307 1074 2335
rect 1320 2307 1322 2335
rect 1576 2307 1578 2335
rect 1816 2307 1818 2335
rect 319 2306 323 2307
rect 319 2301 323 2302
rect 367 2306 371 2307
rect 367 2301 371 2302
rect 551 2306 555 2307
rect 551 2301 555 2302
rect 591 2306 595 2307
rect 591 2301 595 2302
rect 831 2306 835 2307
rect 831 2301 835 2302
rect 1071 2306 1075 2307
rect 1071 2301 1075 2302
rect 1151 2306 1155 2307
rect 1151 2301 1155 2302
rect 1319 2306 1323 2307
rect 1319 2301 1323 2302
rect 1495 2306 1499 2307
rect 1495 2301 1499 2302
rect 1575 2306 1579 2307
rect 1575 2301 1579 2302
rect 1815 2306 1819 2307
rect 1815 2301 1819 2302
rect 320 2277 322 2301
rect 552 2277 554 2301
rect 832 2277 834 2301
rect 1152 2277 1154 2301
rect 1246 2291 1252 2292
rect 1246 2287 1247 2291
rect 1251 2287 1252 2291
rect 1246 2286 1252 2287
rect 318 2276 324 2277
rect 318 2272 319 2276
rect 323 2272 324 2276
rect 318 2271 324 2272
rect 550 2276 556 2277
rect 550 2272 551 2276
rect 555 2272 556 2276
rect 550 2271 556 2272
rect 830 2276 836 2277
rect 830 2272 831 2276
rect 835 2272 836 2276
rect 830 2271 836 2272
rect 1150 2276 1156 2277
rect 1150 2272 1151 2276
rect 1155 2272 1156 2276
rect 1150 2271 1156 2272
rect 290 2261 296 2262
rect 290 2257 291 2261
rect 295 2257 296 2261
rect 290 2256 296 2257
rect 522 2261 528 2262
rect 522 2257 523 2261
rect 527 2257 528 2261
rect 522 2256 528 2257
rect 802 2261 808 2262
rect 802 2257 803 2261
rect 807 2257 808 2261
rect 802 2256 808 2257
rect 1122 2261 1128 2262
rect 1122 2257 1123 2261
rect 1127 2257 1128 2261
rect 1122 2256 1128 2257
rect 218 2243 224 2244
rect 218 2239 219 2243
rect 223 2239 224 2243
rect 218 2238 224 2239
rect 292 2171 294 2256
rect 306 2251 312 2252
rect 306 2247 307 2251
rect 311 2247 312 2251
rect 306 2246 312 2247
rect 308 2220 310 2246
rect 306 2219 312 2220
rect 306 2215 307 2219
rect 311 2215 312 2219
rect 306 2214 312 2215
rect 524 2171 526 2256
rect 538 2251 544 2252
rect 538 2247 539 2251
rect 543 2247 544 2251
rect 538 2246 544 2247
rect 540 2220 542 2246
rect 538 2219 544 2220
rect 538 2215 539 2219
rect 543 2215 544 2219
rect 538 2214 544 2215
rect 804 2171 806 2256
rect 818 2251 824 2252
rect 818 2247 819 2251
rect 823 2247 824 2251
rect 818 2246 824 2247
rect 820 2220 822 2246
rect 818 2219 824 2220
rect 818 2215 819 2219
rect 823 2215 824 2219
rect 818 2214 824 2215
rect 1124 2171 1126 2256
rect 1248 2252 1250 2286
rect 1496 2277 1498 2301
rect 1816 2277 1818 2301
rect 1494 2276 1500 2277
rect 1494 2272 1495 2276
rect 1499 2272 1500 2276
rect 1494 2271 1500 2272
rect 1814 2276 1820 2277
rect 1814 2272 1815 2276
rect 1819 2272 1820 2276
rect 1814 2271 1820 2272
rect 1466 2261 1472 2262
rect 1466 2257 1467 2261
rect 1471 2257 1472 2261
rect 1466 2256 1472 2257
rect 1786 2261 1792 2262
rect 1786 2257 1787 2261
rect 1791 2257 1792 2261
rect 1786 2256 1792 2257
rect 1246 2251 1252 2252
rect 1246 2247 1247 2251
rect 1251 2247 1252 2251
rect 1246 2246 1252 2247
rect 1266 2251 1272 2252
rect 1266 2247 1267 2251
rect 1271 2247 1272 2251
rect 1266 2246 1272 2247
rect 1268 2220 1270 2246
rect 1266 2219 1272 2220
rect 1266 2215 1267 2219
rect 1271 2215 1272 2219
rect 1266 2214 1272 2215
rect 1274 2219 1280 2220
rect 1274 2215 1275 2219
rect 1279 2215 1280 2219
rect 1274 2214 1280 2215
rect 111 2170 115 2171
rect 111 2165 115 2166
rect 131 2170 135 2171
rect 131 2165 135 2166
rect 291 2170 295 2171
rect 291 2165 295 2166
rect 483 2170 487 2171
rect 483 2165 487 2166
rect 523 2170 527 2171
rect 523 2165 527 2166
rect 691 2170 695 2171
rect 691 2165 695 2166
rect 803 2170 807 2171
rect 803 2165 807 2166
rect 915 2170 919 2171
rect 915 2165 919 2166
rect 1123 2170 1127 2171
rect 1123 2165 1127 2166
rect 1147 2170 1151 2171
rect 1147 2165 1151 2166
rect 112 2105 114 2165
rect 110 2104 116 2105
rect 292 2104 294 2165
rect 418 2147 424 2148
rect 418 2143 419 2147
rect 423 2143 424 2147
rect 418 2142 424 2143
rect 420 2112 422 2142
rect 418 2111 424 2112
rect 418 2107 419 2111
rect 423 2107 424 2111
rect 418 2106 424 2107
rect 484 2104 486 2165
rect 692 2104 694 2165
rect 814 2131 820 2132
rect 814 2127 815 2131
rect 819 2127 820 2131
rect 814 2126 820 2127
rect 816 2112 818 2126
rect 814 2111 820 2112
rect 814 2107 815 2111
rect 819 2107 820 2111
rect 814 2106 820 2107
rect 916 2104 918 2165
rect 1018 2147 1024 2148
rect 1002 2143 1008 2144
rect 1002 2139 1003 2143
rect 1007 2139 1008 2143
rect 1018 2143 1019 2147
rect 1023 2143 1024 2147
rect 1018 2142 1024 2143
rect 1002 2138 1008 2139
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 290 2103 296 2104
rect 290 2099 291 2103
rect 295 2099 296 2103
rect 290 2098 296 2099
rect 482 2103 488 2104
rect 482 2099 483 2103
rect 487 2099 488 2103
rect 482 2098 488 2099
rect 690 2103 696 2104
rect 690 2099 691 2103
rect 695 2099 696 2103
rect 690 2098 696 2099
rect 914 2103 920 2104
rect 914 2099 915 2103
rect 919 2099 920 2103
rect 914 2098 920 2099
rect 318 2088 324 2089
rect 110 2087 116 2088
rect 110 2083 111 2087
rect 115 2083 116 2087
rect 318 2084 319 2088
rect 323 2084 324 2088
rect 318 2083 324 2084
rect 510 2088 516 2089
rect 510 2084 511 2088
rect 515 2084 516 2088
rect 510 2083 516 2084
rect 718 2088 724 2089
rect 718 2084 719 2088
rect 723 2084 724 2088
rect 718 2083 724 2084
rect 942 2088 948 2089
rect 942 2084 943 2088
rect 947 2084 948 2088
rect 942 2083 948 2084
rect 110 2082 116 2083
rect 112 2055 114 2082
rect 320 2055 322 2083
rect 512 2055 514 2083
rect 720 2055 722 2083
rect 944 2055 946 2083
rect 111 2054 115 2055
rect 111 2049 115 2050
rect 263 2054 267 2055
rect 263 2049 267 2050
rect 319 2054 323 2055
rect 319 2049 323 2050
rect 399 2054 403 2055
rect 399 2049 403 2050
rect 511 2054 515 2055
rect 511 2049 515 2050
rect 535 2054 539 2055
rect 535 2049 539 2050
rect 679 2054 683 2055
rect 679 2049 683 2050
rect 719 2054 723 2055
rect 719 2049 723 2050
rect 823 2054 827 2055
rect 823 2049 827 2050
rect 943 2054 947 2055
rect 943 2049 947 2050
rect 967 2054 971 2055
rect 967 2049 971 2050
rect 112 2026 114 2049
rect 110 2025 116 2026
rect 264 2025 266 2049
rect 400 2025 402 2049
rect 536 2025 538 2049
rect 680 2025 682 2049
rect 824 2025 826 2049
rect 968 2025 970 2049
rect 110 2021 111 2025
rect 115 2021 116 2025
rect 110 2020 116 2021
rect 262 2024 268 2025
rect 262 2020 263 2024
rect 267 2020 268 2024
rect 262 2019 268 2020
rect 398 2024 404 2025
rect 398 2020 399 2024
rect 403 2020 404 2024
rect 398 2019 404 2020
rect 534 2024 540 2025
rect 534 2020 535 2024
rect 539 2020 540 2024
rect 534 2019 540 2020
rect 678 2024 684 2025
rect 678 2020 679 2024
rect 683 2020 684 2024
rect 678 2019 684 2020
rect 822 2024 828 2025
rect 822 2020 823 2024
rect 827 2020 828 2024
rect 822 2019 828 2020
rect 966 2024 972 2025
rect 966 2020 967 2024
rect 971 2020 972 2024
rect 966 2019 972 2020
rect 234 2009 240 2010
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 234 2005 235 2009
rect 239 2005 240 2009
rect 234 2004 240 2005
rect 370 2009 376 2010
rect 370 2005 371 2009
rect 375 2005 376 2009
rect 370 2004 376 2005
rect 506 2009 512 2010
rect 506 2005 507 2009
rect 511 2005 512 2009
rect 506 2004 512 2005
rect 650 2009 656 2010
rect 650 2005 651 2009
rect 655 2005 656 2009
rect 650 2004 656 2005
rect 794 2009 800 2010
rect 794 2005 795 2009
rect 799 2005 800 2009
rect 794 2004 800 2005
rect 938 2009 944 2010
rect 938 2005 939 2009
rect 943 2005 944 2009
rect 938 2004 944 2005
rect 110 2003 116 2004
rect 112 1931 114 2003
rect 236 1931 238 2004
rect 372 1931 374 2004
rect 386 1999 392 2000
rect 386 1995 387 1999
rect 391 1995 392 1999
rect 386 1994 392 1995
rect 388 1968 390 1994
rect 386 1967 392 1968
rect 386 1963 387 1967
rect 391 1963 392 1967
rect 386 1962 392 1963
rect 508 1931 510 2004
rect 522 1999 528 2000
rect 522 1995 523 1999
rect 527 1995 528 1999
rect 522 1994 528 1995
rect 524 1968 526 1994
rect 522 1967 528 1968
rect 522 1963 523 1967
rect 527 1963 528 1967
rect 522 1962 528 1963
rect 652 1931 654 2004
rect 666 1999 672 2000
rect 666 1995 667 1999
rect 671 1995 672 1999
rect 666 1994 672 1995
rect 668 1968 670 1994
rect 666 1967 672 1968
rect 666 1963 667 1967
rect 671 1963 672 1967
rect 666 1962 672 1963
rect 750 1951 756 1952
rect 750 1947 751 1951
rect 755 1947 756 1951
rect 750 1946 756 1947
rect 111 1930 115 1931
rect 111 1925 115 1926
rect 235 1930 239 1931
rect 235 1925 239 1926
rect 371 1930 375 1931
rect 371 1925 375 1926
rect 435 1930 439 1931
rect 435 1925 439 1926
rect 507 1930 511 1931
rect 507 1925 511 1926
rect 627 1930 631 1931
rect 627 1925 631 1926
rect 651 1930 655 1931
rect 651 1925 655 1926
rect 112 1865 114 1925
rect 110 1864 116 1865
rect 236 1864 238 1925
rect 362 1907 368 1908
rect 322 1903 328 1904
rect 322 1899 323 1903
rect 327 1899 328 1903
rect 362 1903 363 1907
rect 367 1903 368 1907
rect 362 1902 368 1903
rect 322 1898 328 1899
rect 110 1860 111 1864
rect 115 1860 116 1864
rect 110 1859 116 1860
rect 234 1863 240 1864
rect 234 1859 235 1863
rect 239 1859 240 1863
rect 234 1858 240 1859
rect 262 1848 268 1849
rect 110 1847 116 1848
rect 110 1843 111 1847
rect 115 1843 116 1847
rect 262 1844 263 1848
rect 267 1844 268 1848
rect 262 1843 268 1844
rect 110 1842 116 1843
rect 112 1807 114 1842
rect 264 1807 266 1843
rect 111 1806 115 1807
rect 111 1801 115 1802
rect 223 1806 227 1807
rect 223 1801 227 1802
rect 263 1806 267 1807
rect 263 1801 267 1802
rect 112 1778 114 1801
rect 110 1777 116 1778
rect 224 1777 226 1801
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 110 1772 116 1773
rect 222 1776 228 1777
rect 222 1772 223 1776
rect 227 1772 228 1776
rect 222 1771 228 1772
rect 194 1761 200 1762
rect 110 1760 116 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 194 1757 195 1761
rect 199 1757 200 1761
rect 194 1756 200 1757
rect 110 1755 116 1756
rect 112 1683 114 1755
rect 196 1683 198 1756
rect 324 1752 326 1898
rect 364 1872 366 1902
rect 362 1871 368 1872
rect 362 1867 363 1871
rect 367 1867 368 1871
rect 362 1866 368 1867
rect 436 1864 438 1925
rect 562 1907 568 1908
rect 562 1903 563 1907
rect 567 1903 568 1907
rect 562 1902 568 1903
rect 564 1872 566 1902
rect 562 1871 568 1872
rect 562 1867 563 1871
rect 567 1867 568 1871
rect 562 1866 568 1867
rect 628 1864 630 1925
rect 752 1872 754 1946
rect 796 1931 798 2004
rect 810 1999 816 2000
rect 810 1995 811 1999
rect 815 1995 816 1999
rect 810 1994 816 1995
rect 812 1968 814 1994
rect 930 1991 936 1992
rect 930 1987 931 1991
rect 935 1987 936 1991
rect 930 1986 936 1987
rect 810 1967 816 1968
rect 810 1963 811 1967
rect 815 1963 816 1967
rect 810 1962 816 1963
rect 795 1930 799 1931
rect 795 1925 799 1926
rect 811 1930 815 1931
rect 811 1925 815 1926
rect 750 1871 756 1872
rect 750 1867 751 1871
rect 755 1867 756 1871
rect 750 1866 756 1867
rect 812 1864 814 1925
rect 932 1908 934 1986
rect 940 1931 942 2004
rect 1004 2000 1006 2138
rect 1020 2120 1022 2142
rect 1018 2119 1024 2120
rect 1018 2115 1019 2119
rect 1023 2115 1024 2119
rect 1018 2114 1024 2115
rect 1148 2104 1150 2165
rect 1276 2112 1278 2214
rect 1468 2171 1470 2256
rect 1788 2171 1790 2256
rect 1876 2220 1878 2358
rect 1936 2357 1938 2417
rect 1976 2409 1978 2469
rect 2298 2451 2304 2452
rect 2298 2447 2299 2451
rect 2303 2447 2304 2451
rect 2298 2446 2304 2447
rect 1974 2408 1980 2409
rect 1974 2404 1975 2408
rect 1979 2404 1980 2408
rect 1974 2403 1980 2404
rect 1974 2391 1980 2392
rect 1974 2387 1975 2391
rect 1979 2387 1980 2391
rect 1974 2386 1980 2387
rect 1934 2356 1940 2357
rect 1934 2352 1935 2356
rect 1939 2352 1940 2356
rect 1976 2355 1978 2386
rect 1934 2351 1940 2352
rect 1975 2354 1979 2355
rect 1975 2349 1979 2350
rect 2223 2354 2227 2355
rect 2223 2349 2227 2350
rect 1934 2339 1940 2340
rect 1934 2335 1935 2339
rect 1939 2335 1940 2339
rect 1934 2334 1940 2335
rect 1936 2307 1938 2334
rect 1976 2326 1978 2349
rect 1974 2325 1980 2326
rect 2224 2325 2226 2349
rect 1974 2321 1975 2325
rect 1979 2321 1980 2325
rect 1974 2320 1980 2321
rect 2222 2324 2228 2325
rect 2222 2320 2223 2324
rect 2227 2320 2228 2324
rect 2222 2319 2228 2320
rect 2194 2309 2200 2310
rect 1974 2308 1980 2309
rect 1935 2306 1939 2307
rect 1974 2304 1975 2308
rect 1979 2304 1980 2308
rect 2194 2305 2195 2309
rect 2199 2305 2200 2309
rect 2194 2304 2200 2305
rect 1974 2303 1980 2304
rect 1935 2301 1939 2302
rect 1936 2278 1938 2301
rect 1934 2277 1940 2278
rect 1934 2273 1935 2277
rect 1939 2273 1940 2277
rect 1934 2272 1940 2273
rect 1934 2260 1940 2261
rect 1934 2256 1935 2260
rect 1939 2256 1940 2260
rect 1934 2255 1940 2256
rect 1914 2251 1920 2252
rect 1914 2247 1915 2251
rect 1919 2247 1920 2251
rect 1914 2246 1920 2247
rect 1916 2220 1918 2246
rect 1874 2219 1880 2220
rect 1874 2215 1875 2219
rect 1879 2215 1880 2219
rect 1874 2214 1880 2215
rect 1914 2219 1920 2220
rect 1914 2215 1915 2219
rect 1919 2215 1920 2219
rect 1914 2214 1920 2215
rect 1936 2171 1938 2255
rect 1976 2243 1978 2303
rect 2196 2243 2198 2304
rect 2300 2300 2302 2446
rect 2308 2408 2310 2469
rect 2434 2451 2440 2452
rect 2434 2447 2435 2451
rect 2439 2447 2440 2451
rect 2434 2446 2440 2447
rect 2436 2416 2438 2446
rect 2434 2415 2440 2416
rect 2434 2411 2435 2415
rect 2439 2411 2440 2415
rect 2434 2410 2440 2411
rect 2516 2408 2518 2469
rect 2642 2451 2648 2452
rect 2642 2447 2643 2451
rect 2647 2447 2648 2451
rect 2642 2446 2648 2447
rect 2644 2416 2646 2446
rect 2642 2415 2648 2416
rect 2642 2411 2643 2415
rect 2647 2411 2648 2415
rect 2642 2410 2648 2411
rect 2716 2408 2718 2469
rect 2840 2416 2842 2510
rect 2892 2475 2894 2552
rect 2978 2539 2984 2540
rect 2978 2535 2979 2539
rect 2983 2535 2984 2539
rect 2978 2534 2984 2535
rect 2980 2516 2982 2534
rect 3014 2531 3020 2532
rect 3014 2527 3015 2531
rect 3019 2527 3020 2531
rect 3014 2526 3020 2527
rect 2978 2515 2984 2516
rect 2978 2511 2979 2515
rect 2983 2511 2984 2515
rect 2978 2510 2984 2511
rect 2891 2474 2895 2475
rect 2891 2469 2895 2470
rect 2907 2474 2911 2475
rect 2907 2469 2911 2470
rect 2838 2415 2844 2416
rect 2838 2411 2839 2415
rect 2843 2411 2844 2415
rect 2838 2410 2844 2411
rect 2908 2408 2910 2469
rect 3016 2452 3018 2526
rect 3028 2475 3030 2552
rect 3042 2547 3048 2548
rect 3042 2543 3043 2547
rect 3047 2543 3048 2547
rect 3042 2542 3048 2543
rect 3044 2516 3046 2542
rect 3042 2515 3048 2516
rect 3042 2511 3043 2515
rect 3047 2511 3048 2515
rect 3042 2510 3048 2511
rect 3164 2475 3166 2552
rect 3178 2547 3184 2548
rect 3178 2543 3179 2547
rect 3183 2543 3184 2547
rect 3178 2542 3184 2543
rect 3180 2516 3182 2542
rect 3272 2540 3274 2654
rect 3800 2653 3802 2713
rect 3840 2683 3842 2755
rect 3892 2683 3894 2756
rect 3980 2720 3982 2858
rect 3996 2856 3998 2917
rect 4174 2899 4180 2900
rect 4174 2895 4175 2899
rect 4179 2895 4180 2899
rect 4174 2894 4180 2895
rect 4176 2864 4178 2894
rect 4174 2863 4180 2864
rect 4174 2859 4175 2863
rect 4179 2859 4180 2863
rect 4174 2858 4180 2859
rect 4212 2856 4214 2917
rect 4298 2895 4304 2896
rect 4298 2891 4299 2895
rect 4303 2891 4304 2895
rect 4298 2890 4304 2891
rect 4300 2872 4302 2890
rect 4298 2871 4304 2872
rect 4298 2867 4299 2871
rect 4303 2867 4304 2871
rect 4298 2866 4304 2867
rect 4444 2856 4446 2917
rect 4548 2900 4550 2998
rect 4644 2923 4646 3008
rect 4660 2972 4662 3106
rect 4860 3104 4862 3165
rect 4986 3147 4992 3148
rect 4986 3143 4987 3147
rect 4991 3143 4992 3147
rect 4986 3142 4992 3143
rect 4988 3112 4990 3142
rect 4986 3111 4992 3112
rect 4986 3107 4987 3111
rect 4991 3107 4992 3111
rect 4986 3106 4992 3107
rect 5076 3104 5078 3165
rect 5202 3147 5208 3148
rect 5202 3143 5203 3147
rect 5207 3143 5208 3147
rect 5202 3142 5208 3143
rect 5204 3112 5206 3142
rect 5202 3111 5208 3112
rect 5202 3107 5203 3111
rect 5207 3107 5208 3111
rect 5202 3106 5208 3107
rect 5308 3104 5310 3165
rect 4858 3103 4864 3104
rect 4858 3099 4859 3103
rect 4863 3099 4864 3103
rect 4858 3098 4864 3099
rect 5074 3103 5080 3104
rect 5074 3099 5075 3103
rect 5079 3099 5080 3103
rect 5074 3098 5080 3099
rect 5306 3103 5312 3104
rect 5306 3099 5307 3103
rect 5311 3099 5312 3103
rect 5306 3098 5312 3099
rect 4678 3088 4684 3089
rect 4678 3084 4679 3088
rect 4683 3084 4684 3088
rect 4678 3083 4684 3084
rect 4886 3088 4892 3089
rect 4886 3084 4887 3088
rect 4891 3084 4892 3088
rect 4886 3083 4892 3084
rect 5102 3088 5108 3089
rect 5102 3084 5103 3088
rect 5107 3084 5108 3088
rect 5102 3083 5108 3084
rect 5334 3088 5340 3089
rect 5334 3084 5335 3088
rect 5339 3084 5340 3088
rect 5334 3083 5340 3084
rect 4680 3059 4682 3083
rect 4888 3059 4890 3083
rect 5104 3059 5106 3083
rect 5336 3059 5338 3083
rect 4671 3058 4675 3059
rect 4671 3053 4675 3054
rect 4679 3058 4683 3059
rect 4679 3053 4683 3054
rect 4887 3058 4891 3059
rect 4887 3053 4891 3054
rect 4911 3058 4915 3059
rect 4911 3053 4915 3054
rect 5103 3058 5107 3059
rect 5103 3053 5107 3054
rect 5167 3058 5171 3059
rect 5167 3053 5171 3054
rect 5335 3058 5339 3059
rect 5335 3053 5339 3054
rect 4672 3029 4674 3053
rect 4912 3029 4914 3053
rect 5168 3029 5170 3053
rect 5262 3043 5268 3044
rect 5262 3039 5263 3043
rect 5267 3039 5268 3043
rect 5262 3038 5268 3039
rect 4670 3028 4676 3029
rect 4670 3024 4671 3028
rect 4675 3024 4676 3028
rect 4670 3023 4676 3024
rect 4910 3028 4916 3029
rect 4910 3024 4911 3028
rect 4915 3024 4916 3028
rect 4910 3023 4916 3024
rect 5166 3028 5172 3029
rect 5166 3024 5167 3028
rect 5171 3024 5172 3028
rect 5166 3023 5172 3024
rect 4882 3013 4888 3014
rect 4882 3009 4883 3013
rect 4887 3009 4888 3013
rect 4882 3008 4888 3009
rect 5138 3013 5144 3014
rect 5138 3009 5139 3013
rect 5143 3009 5144 3013
rect 5138 3008 5144 3009
rect 4658 2971 4664 2972
rect 4658 2967 4659 2971
rect 4663 2967 4664 2971
rect 4658 2966 4664 2967
rect 4884 2923 4886 3008
rect 4898 3003 4904 3004
rect 4898 2999 4899 3003
rect 4903 2999 4904 3003
rect 4898 2998 4904 2999
rect 4900 2972 4902 2998
rect 4898 2971 4904 2972
rect 4898 2967 4899 2971
rect 4903 2967 4904 2971
rect 4898 2966 4904 2967
rect 5140 2923 5142 3008
rect 5264 3004 5266 3038
rect 5364 3004 5366 3206
rect 5516 3171 5518 3248
rect 5604 3212 5606 3470
rect 5664 3411 5666 3479
rect 5663 3410 5667 3411
rect 5663 3405 5667 3406
rect 5664 3345 5666 3405
rect 5662 3344 5668 3345
rect 5662 3340 5663 3344
rect 5667 3340 5668 3344
rect 5662 3339 5668 3340
rect 5662 3327 5668 3328
rect 5662 3323 5663 3327
rect 5667 3323 5668 3327
rect 5662 3322 5668 3323
rect 5664 3299 5666 3322
rect 5663 3298 5667 3299
rect 5663 3293 5667 3294
rect 5664 3270 5666 3293
rect 5662 3269 5668 3270
rect 5662 3265 5663 3269
rect 5667 3265 5668 3269
rect 5662 3264 5668 3265
rect 5662 3252 5668 3253
rect 5662 3248 5663 3252
rect 5667 3248 5668 3252
rect 5662 3247 5668 3248
rect 5618 3243 5624 3244
rect 5618 3239 5619 3243
rect 5623 3239 5624 3243
rect 5618 3238 5624 3239
rect 5602 3211 5608 3212
rect 5602 3207 5603 3211
rect 5607 3207 5608 3211
rect 5602 3206 5608 3207
rect 5515 3170 5519 3171
rect 5515 3165 5519 3166
rect 5430 3131 5436 3132
rect 5430 3127 5431 3131
rect 5435 3127 5436 3131
rect 5430 3126 5436 3127
rect 5432 3112 5434 3126
rect 5430 3111 5436 3112
rect 5430 3107 5431 3111
rect 5435 3107 5436 3111
rect 5430 3106 5436 3107
rect 5516 3104 5518 3165
rect 5620 3148 5622 3238
rect 5664 3171 5666 3247
rect 5663 3170 5667 3171
rect 5663 3165 5667 3166
rect 5618 3147 5624 3148
rect 5618 3143 5619 3147
rect 5623 3143 5624 3147
rect 5618 3142 5624 3143
rect 5618 3111 5624 3112
rect 5618 3107 5619 3111
rect 5623 3107 5624 3111
rect 5618 3106 5624 3107
rect 5514 3103 5520 3104
rect 5514 3099 5515 3103
rect 5519 3099 5520 3103
rect 5514 3098 5520 3099
rect 5542 3088 5548 3089
rect 5542 3084 5543 3088
rect 5547 3084 5548 3088
rect 5542 3083 5548 3084
rect 5544 3059 5546 3083
rect 5423 3058 5427 3059
rect 5423 3053 5427 3054
rect 5543 3058 5547 3059
rect 5543 3053 5547 3054
rect 5424 3029 5426 3053
rect 5422 3028 5428 3029
rect 5422 3024 5423 3028
rect 5427 3024 5428 3028
rect 5422 3023 5428 3024
rect 5394 3013 5400 3014
rect 5394 3009 5395 3013
rect 5399 3009 5400 3013
rect 5394 3008 5400 3009
rect 5154 3003 5160 3004
rect 5154 2999 5155 3003
rect 5159 2999 5160 3003
rect 5154 2998 5160 2999
rect 5262 3003 5268 3004
rect 5262 2999 5263 3003
rect 5267 2999 5268 3003
rect 5262 2998 5268 2999
rect 5362 3003 5368 3004
rect 5362 2999 5363 3003
rect 5367 2999 5368 3003
rect 5362 2998 5368 2999
rect 5156 2972 5158 2998
rect 5154 2971 5160 2972
rect 5154 2967 5155 2971
rect 5159 2967 5160 2971
rect 5154 2966 5160 2967
rect 5396 2923 5398 3008
rect 5410 2971 5416 2972
rect 5410 2967 5411 2971
rect 5415 2967 5416 2971
rect 5410 2966 5416 2967
rect 4643 2922 4647 2923
rect 4643 2917 4647 2918
rect 4699 2922 4703 2923
rect 4699 2917 4703 2918
rect 4883 2922 4887 2923
rect 4883 2917 4887 2918
rect 4971 2922 4975 2923
rect 4971 2917 4975 2918
rect 5139 2922 5143 2923
rect 5139 2917 5143 2918
rect 5251 2922 5255 2923
rect 5251 2917 5255 2918
rect 5395 2922 5399 2923
rect 5395 2917 5399 2918
rect 4546 2899 4552 2900
rect 4546 2895 4547 2899
rect 4551 2895 4552 2899
rect 4546 2894 4552 2895
rect 4570 2899 4576 2900
rect 4570 2895 4571 2899
rect 4575 2895 4576 2899
rect 4570 2894 4576 2895
rect 4572 2864 4574 2894
rect 4570 2863 4576 2864
rect 4570 2859 4571 2863
rect 4575 2859 4576 2863
rect 4570 2858 4576 2859
rect 4700 2856 4702 2917
rect 4826 2899 4832 2900
rect 4826 2895 4827 2899
rect 4831 2895 4832 2899
rect 4826 2894 4832 2895
rect 4828 2864 4830 2894
rect 4826 2863 4832 2864
rect 4826 2859 4827 2863
rect 4831 2859 4832 2863
rect 4826 2858 4832 2859
rect 4972 2856 4974 2917
rect 5252 2856 5254 2917
rect 5338 2895 5344 2896
rect 5338 2891 5339 2895
rect 5343 2891 5344 2895
rect 5338 2890 5344 2891
rect 3994 2855 4000 2856
rect 3994 2851 3995 2855
rect 3999 2851 4000 2855
rect 3994 2850 4000 2851
rect 4210 2855 4216 2856
rect 4210 2851 4211 2855
rect 4215 2851 4216 2855
rect 4210 2850 4216 2851
rect 4442 2855 4448 2856
rect 4442 2851 4443 2855
rect 4447 2851 4448 2855
rect 4442 2850 4448 2851
rect 4698 2855 4704 2856
rect 4698 2851 4699 2855
rect 4703 2851 4704 2855
rect 4698 2850 4704 2851
rect 4970 2855 4976 2856
rect 4970 2851 4971 2855
rect 4975 2851 4976 2855
rect 4970 2850 4976 2851
rect 5250 2855 5256 2856
rect 5250 2851 5251 2855
rect 5255 2851 5256 2855
rect 5250 2850 5256 2851
rect 4022 2840 4028 2841
rect 4022 2836 4023 2840
rect 4027 2836 4028 2840
rect 4022 2835 4028 2836
rect 4238 2840 4244 2841
rect 4238 2836 4239 2840
rect 4243 2836 4244 2840
rect 4238 2835 4244 2836
rect 4470 2840 4476 2841
rect 4470 2836 4471 2840
rect 4475 2836 4476 2840
rect 4470 2835 4476 2836
rect 4726 2840 4732 2841
rect 4726 2836 4727 2840
rect 4731 2836 4732 2840
rect 4726 2835 4732 2836
rect 4998 2840 5004 2841
rect 4998 2836 4999 2840
rect 5003 2836 5004 2840
rect 4998 2835 5004 2836
rect 5278 2840 5284 2841
rect 5278 2836 5279 2840
rect 5283 2836 5284 2840
rect 5278 2835 5284 2836
rect 4024 2807 4026 2835
rect 4240 2807 4242 2835
rect 4472 2807 4474 2835
rect 4728 2807 4730 2835
rect 5000 2807 5002 2835
rect 5280 2807 5282 2835
rect 4023 2806 4027 2807
rect 4023 2801 4027 2802
rect 4055 2806 4059 2807
rect 4055 2801 4059 2802
rect 4191 2806 4195 2807
rect 4191 2801 4195 2802
rect 4239 2806 4243 2807
rect 4239 2801 4243 2802
rect 4327 2806 4331 2807
rect 4327 2801 4331 2802
rect 4463 2806 4467 2807
rect 4463 2801 4467 2802
rect 4471 2806 4475 2807
rect 4471 2801 4475 2802
rect 4727 2806 4731 2807
rect 4727 2801 4731 2802
rect 4999 2806 5003 2807
rect 4999 2801 5003 2802
rect 5279 2806 5283 2807
rect 5279 2801 5283 2802
rect 4056 2777 4058 2801
rect 4192 2777 4194 2801
rect 4328 2777 4330 2801
rect 4464 2777 4466 2801
rect 4054 2776 4060 2777
rect 4054 2772 4055 2776
rect 4059 2772 4060 2776
rect 4054 2771 4060 2772
rect 4190 2776 4196 2777
rect 4190 2772 4191 2776
rect 4195 2772 4196 2776
rect 4190 2771 4196 2772
rect 4326 2776 4332 2777
rect 4326 2772 4327 2776
rect 4331 2772 4332 2776
rect 4326 2771 4332 2772
rect 4462 2776 4468 2777
rect 4462 2772 4463 2776
rect 4467 2772 4468 2776
rect 4462 2771 4468 2772
rect 4026 2761 4032 2762
rect 4026 2757 4027 2761
rect 4031 2757 4032 2761
rect 4026 2756 4032 2757
rect 4162 2761 4168 2762
rect 4162 2757 4163 2761
rect 4167 2757 4168 2761
rect 4162 2756 4168 2757
rect 4298 2761 4304 2762
rect 4298 2757 4299 2761
rect 4303 2757 4304 2761
rect 4298 2756 4304 2757
rect 4434 2761 4440 2762
rect 4434 2757 4435 2761
rect 4439 2757 4440 2761
rect 4434 2756 4440 2757
rect 3978 2719 3984 2720
rect 3978 2715 3979 2719
rect 3983 2715 3984 2719
rect 3978 2714 3984 2715
rect 4028 2683 4030 2756
rect 4042 2751 4048 2752
rect 4042 2747 4043 2751
rect 4047 2747 4048 2751
rect 4042 2746 4048 2747
rect 4044 2720 4046 2746
rect 4042 2719 4048 2720
rect 4042 2715 4043 2719
rect 4047 2715 4048 2719
rect 4042 2714 4048 2715
rect 4164 2683 4166 2756
rect 4178 2751 4184 2752
rect 4178 2747 4179 2751
rect 4183 2747 4184 2751
rect 4178 2746 4184 2747
rect 4180 2720 4182 2746
rect 4218 2743 4224 2744
rect 4218 2739 4219 2743
rect 4223 2739 4224 2743
rect 4218 2738 4224 2739
rect 4178 2719 4184 2720
rect 4178 2715 4179 2719
rect 4183 2715 4184 2719
rect 4178 2714 4184 2715
rect 3839 2682 3843 2683
rect 3839 2677 3843 2678
rect 3891 2682 3895 2683
rect 3891 2677 3895 2678
rect 4027 2682 4031 2683
rect 4027 2677 4031 2678
rect 4099 2682 4103 2683
rect 4099 2677 4103 2678
rect 4163 2682 4167 2683
rect 4163 2677 4167 2678
rect 3798 2652 3804 2653
rect 3798 2648 3799 2652
rect 3803 2648 3804 2652
rect 3798 2647 3804 2648
rect 3798 2635 3804 2636
rect 3798 2631 3799 2635
rect 3803 2631 3804 2635
rect 3798 2630 3804 2631
rect 3800 2603 3802 2630
rect 3840 2617 3842 2677
rect 3838 2616 3844 2617
rect 4100 2616 4102 2677
rect 4220 2660 4222 2738
rect 4300 2683 4302 2756
rect 4314 2751 4320 2752
rect 4314 2747 4315 2751
rect 4319 2747 4320 2751
rect 4314 2746 4320 2747
rect 4316 2720 4318 2746
rect 4314 2719 4320 2720
rect 4314 2715 4315 2719
rect 4319 2715 4320 2719
rect 4314 2714 4320 2715
rect 4436 2683 4438 2756
rect 4450 2751 4456 2752
rect 4450 2747 4451 2751
rect 4455 2747 4456 2751
rect 4450 2746 4456 2747
rect 4452 2720 4454 2746
rect 4450 2719 4456 2720
rect 4450 2715 4451 2719
rect 4455 2715 4456 2719
rect 4450 2714 4456 2715
rect 4299 2682 4303 2683
rect 4299 2677 4303 2678
rect 4435 2682 4439 2683
rect 4435 2677 4439 2678
rect 4515 2682 4519 2683
rect 4515 2677 4519 2678
rect 4755 2682 4759 2683
rect 4755 2677 4759 2678
rect 5011 2682 5015 2683
rect 5011 2677 5015 2678
rect 5275 2682 5279 2683
rect 5275 2677 5279 2678
rect 4218 2659 4224 2660
rect 4218 2655 4219 2659
rect 4223 2655 4224 2659
rect 4218 2654 4224 2655
rect 4226 2659 4232 2660
rect 4226 2655 4227 2659
rect 4231 2655 4232 2659
rect 4226 2654 4232 2655
rect 4228 2624 4230 2654
rect 4226 2623 4232 2624
rect 4226 2619 4227 2623
rect 4231 2619 4232 2623
rect 4226 2618 4232 2619
rect 4300 2616 4302 2677
rect 4426 2659 4432 2660
rect 4426 2655 4427 2659
rect 4431 2655 4432 2659
rect 4426 2654 4432 2655
rect 4428 2624 4430 2654
rect 4426 2623 4432 2624
rect 4426 2619 4427 2623
rect 4431 2619 4432 2623
rect 4426 2618 4432 2619
rect 4516 2616 4518 2677
rect 4642 2659 4648 2660
rect 4642 2655 4643 2659
rect 4647 2655 4648 2659
rect 4642 2654 4648 2655
rect 4644 2624 4646 2654
rect 4642 2623 4648 2624
rect 4642 2619 4643 2623
rect 4647 2619 4648 2623
rect 4642 2618 4648 2619
rect 4756 2616 4758 2677
rect 4882 2659 4888 2660
rect 4882 2655 4883 2659
rect 4887 2655 4888 2659
rect 4882 2654 4888 2655
rect 4884 2624 4886 2654
rect 4882 2623 4888 2624
rect 4882 2619 4883 2623
rect 4887 2619 4888 2623
rect 4882 2618 4888 2619
rect 4998 2623 5004 2624
rect 4998 2619 4999 2623
rect 5003 2619 5004 2623
rect 4998 2618 5004 2619
rect 3838 2612 3839 2616
rect 3843 2612 3844 2616
rect 3838 2611 3844 2612
rect 4098 2615 4104 2616
rect 4098 2611 4099 2615
rect 4103 2611 4104 2615
rect 4098 2610 4104 2611
rect 4298 2615 4304 2616
rect 4298 2611 4299 2615
rect 4303 2611 4304 2615
rect 4298 2610 4304 2611
rect 4514 2615 4520 2616
rect 4514 2611 4515 2615
rect 4519 2611 4520 2615
rect 4514 2610 4520 2611
rect 4754 2615 4760 2616
rect 4754 2611 4755 2615
rect 4759 2611 4760 2615
rect 4754 2610 4760 2611
rect 3327 2602 3331 2603
rect 3327 2597 3331 2598
rect 3463 2602 3467 2603
rect 3463 2597 3467 2598
rect 3799 2602 3803 2603
rect 4126 2600 4132 2601
rect 3799 2597 3803 2598
rect 3838 2599 3844 2600
rect 3328 2573 3330 2597
rect 3464 2573 3466 2597
rect 3800 2574 3802 2597
rect 3838 2595 3839 2599
rect 3843 2595 3844 2599
rect 4126 2596 4127 2600
rect 4131 2596 4132 2600
rect 4126 2595 4132 2596
rect 4326 2600 4332 2601
rect 4326 2596 4327 2600
rect 4331 2596 4332 2600
rect 4326 2595 4332 2596
rect 4542 2600 4548 2601
rect 4542 2596 4543 2600
rect 4547 2596 4548 2600
rect 4542 2595 4548 2596
rect 4782 2600 4788 2601
rect 4782 2596 4783 2600
rect 4787 2596 4788 2600
rect 4782 2595 4788 2596
rect 3838 2594 3844 2595
rect 3798 2573 3804 2574
rect 3326 2572 3332 2573
rect 3326 2568 3327 2572
rect 3331 2568 3332 2572
rect 3326 2567 3332 2568
rect 3462 2572 3468 2573
rect 3462 2568 3463 2572
rect 3467 2568 3468 2572
rect 3798 2569 3799 2573
rect 3803 2569 3804 2573
rect 3798 2568 3804 2569
rect 3462 2567 3468 2568
rect 3840 2567 3842 2594
rect 4128 2567 4130 2595
rect 4328 2567 4330 2595
rect 4544 2567 4546 2595
rect 4784 2567 4786 2595
rect 3839 2566 3843 2567
rect 3839 2561 3843 2562
rect 4127 2566 4131 2567
rect 4127 2561 4131 2562
rect 4327 2566 4331 2567
rect 4327 2561 4331 2562
rect 4495 2566 4499 2567
rect 4495 2561 4499 2562
rect 4543 2566 4547 2567
rect 4543 2561 4547 2562
rect 4631 2566 4635 2567
rect 4631 2561 4635 2562
rect 4767 2566 4771 2567
rect 4767 2561 4771 2562
rect 4783 2566 4787 2567
rect 4783 2561 4787 2562
rect 4903 2566 4907 2567
rect 4903 2561 4907 2562
rect 3298 2557 3304 2558
rect 3298 2553 3299 2557
rect 3303 2553 3304 2557
rect 3298 2552 3304 2553
rect 3434 2557 3440 2558
rect 3434 2553 3435 2557
rect 3439 2553 3440 2557
rect 3434 2552 3440 2553
rect 3798 2556 3804 2557
rect 3798 2552 3799 2556
rect 3803 2552 3804 2556
rect 3270 2539 3276 2540
rect 3270 2535 3271 2539
rect 3275 2535 3276 2539
rect 3270 2534 3276 2535
rect 3178 2515 3184 2516
rect 3178 2511 3179 2515
rect 3183 2511 3184 2515
rect 3178 2510 3184 2511
rect 3300 2475 3302 2552
rect 3314 2547 3320 2548
rect 3314 2543 3315 2547
rect 3319 2543 3320 2547
rect 3314 2542 3320 2543
rect 3316 2516 3318 2542
rect 3314 2515 3320 2516
rect 3314 2511 3315 2515
rect 3319 2511 3320 2515
rect 3314 2510 3320 2511
rect 3436 2475 3438 2552
rect 3798 2551 3804 2552
rect 3450 2547 3456 2548
rect 3450 2543 3451 2547
rect 3455 2543 3456 2547
rect 3450 2542 3456 2543
rect 3452 2516 3454 2542
rect 3450 2515 3456 2516
rect 3450 2511 3451 2515
rect 3455 2511 3456 2515
rect 3450 2510 3456 2511
rect 3800 2475 3802 2551
rect 3840 2538 3842 2561
rect 3838 2537 3844 2538
rect 4496 2537 4498 2561
rect 4632 2537 4634 2561
rect 4768 2537 4770 2561
rect 4904 2537 4906 2561
rect 3838 2533 3839 2537
rect 3843 2533 3844 2537
rect 3838 2532 3844 2533
rect 4494 2536 4500 2537
rect 4494 2532 4495 2536
rect 4499 2532 4500 2536
rect 4494 2531 4500 2532
rect 4630 2536 4636 2537
rect 4630 2532 4631 2536
rect 4635 2532 4636 2536
rect 4630 2531 4636 2532
rect 4766 2536 4772 2537
rect 4766 2532 4767 2536
rect 4771 2532 4772 2536
rect 4766 2531 4772 2532
rect 4902 2536 4908 2537
rect 4902 2532 4903 2536
rect 4907 2532 4908 2536
rect 4902 2531 4908 2532
rect 4466 2521 4472 2522
rect 3838 2520 3844 2521
rect 3838 2516 3839 2520
rect 3843 2516 3844 2520
rect 4466 2517 4467 2521
rect 4471 2517 4472 2521
rect 4466 2516 4472 2517
rect 4602 2521 4608 2522
rect 4602 2517 4603 2521
rect 4607 2517 4608 2521
rect 4602 2516 4608 2517
rect 4738 2521 4744 2522
rect 4738 2517 4739 2521
rect 4743 2517 4744 2521
rect 4738 2516 4744 2517
rect 4874 2521 4880 2522
rect 4874 2517 4875 2521
rect 4879 2517 4880 2521
rect 4874 2516 4880 2517
rect 3838 2515 3844 2516
rect 3027 2474 3031 2475
rect 3027 2469 3031 2470
rect 3099 2474 3103 2475
rect 3099 2469 3103 2470
rect 3163 2474 3167 2475
rect 3163 2469 3167 2470
rect 3283 2474 3287 2475
rect 3283 2469 3287 2470
rect 3299 2474 3303 2475
rect 3299 2469 3303 2470
rect 3435 2474 3439 2475
rect 3435 2469 3439 2470
rect 3467 2474 3471 2475
rect 3467 2469 3471 2470
rect 3651 2474 3655 2475
rect 3651 2469 3655 2470
rect 3799 2474 3803 2475
rect 3799 2469 3803 2470
rect 3014 2451 3020 2452
rect 3014 2447 3015 2451
rect 3019 2447 3020 2451
rect 3014 2446 3020 2447
rect 3034 2451 3040 2452
rect 3034 2447 3035 2451
rect 3039 2447 3040 2451
rect 3034 2446 3040 2447
rect 3036 2416 3038 2446
rect 3034 2415 3040 2416
rect 3034 2411 3035 2415
rect 3039 2411 3040 2415
rect 3034 2410 3040 2411
rect 3100 2408 3102 2469
rect 3226 2451 3232 2452
rect 3226 2447 3227 2451
rect 3231 2447 3232 2451
rect 3226 2446 3232 2447
rect 3228 2416 3230 2446
rect 3226 2415 3232 2416
rect 3226 2411 3227 2415
rect 3231 2411 3232 2415
rect 3226 2410 3232 2411
rect 3284 2408 3286 2469
rect 3410 2451 3416 2452
rect 3410 2447 3411 2451
rect 3415 2447 3416 2451
rect 3410 2446 3416 2447
rect 3412 2416 3414 2446
rect 3410 2415 3416 2416
rect 3410 2411 3411 2415
rect 3415 2411 3416 2415
rect 3410 2410 3416 2411
rect 3468 2408 3470 2469
rect 3594 2451 3600 2452
rect 3594 2447 3595 2451
rect 3599 2447 3600 2451
rect 3594 2446 3600 2447
rect 3596 2416 3598 2446
rect 3594 2415 3600 2416
rect 3594 2411 3595 2415
rect 3599 2411 3600 2415
rect 3594 2410 3600 2411
rect 3652 2408 3654 2469
rect 3738 2415 3744 2416
rect 3738 2411 3739 2415
rect 3743 2411 3744 2415
rect 3738 2410 3744 2411
rect 2306 2407 2312 2408
rect 2306 2403 2307 2407
rect 2311 2403 2312 2407
rect 2306 2402 2312 2403
rect 2514 2407 2520 2408
rect 2514 2403 2515 2407
rect 2519 2403 2520 2407
rect 2514 2402 2520 2403
rect 2714 2407 2720 2408
rect 2714 2403 2715 2407
rect 2719 2403 2720 2407
rect 2714 2402 2720 2403
rect 2906 2407 2912 2408
rect 2906 2403 2907 2407
rect 2911 2403 2912 2407
rect 2906 2402 2912 2403
rect 3098 2407 3104 2408
rect 3098 2403 3099 2407
rect 3103 2403 3104 2407
rect 3098 2402 3104 2403
rect 3282 2407 3288 2408
rect 3282 2403 3283 2407
rect 3287 2403 3288 2407
rect 3282 2402 3288 2403
rect 3466 2407 3472 2408
rect 3466 2403 3467 2407
rect 3471 2403 3472 2407
rect 3466 2402 3472 2403
rect 3650 2407 3656 2408
rect 3650 2403 3651 2407
rect 3655 2403 3656 2407
rect 3650 2402 3656 2403
rect 2334 2392 2340 2393
rect 2334 2388 2335 2392
rect 2339 2388 2340 2392
rect 2334 2387 2340 2388
rect 2542 2392 2548 2393
rect 2542 2388 2543 2392
rect 2547 2388 2548 2392
rect 2542 2387 2548 2388
rect 2742 2392 2748 2393
rect 2742 2388 2743 2392
rect 2747 2388 2748 2392
rect 2742 2387 2748 2388
rect 2934 2392 2940 2393
rect 2934 2388 2935 2392
rect 2939 2388 2940 2392
rect 2934 2387 2940 2388
rect 3126 2392 3132 2393
rect 3126 2388 3127 2392
rect 3131 2388 3132 2392
rect 3126 2387 3132 2388
rect 3310 2392 3316 2393
rect 3310 2388 3311 2392
rect 3315 2388 3316 2392
rect 3310 2387 3316 2388
rect 3494 2392 3500 2393
rect 3494 2388 3495 2392
rect 3499 2388 3500 2392
rect 3494 2387 3500 2388
rect 3678 2392 3684 2393
rect 3678 2388 3679 2392
rect 3683 2388 3684 2392
rect 3678 2387 3684 2388
rect 2336 2355 2338 2387
rect 2544 2355 2546 2387
rect 2744 2355 2746 2387
rect 2936 2355 2938 2387
rect 3128 2355 3130 2387
rect 3312 2355 3314 2387
rect 3496 2355 3498 2387
rect 3680 2355 3682 2387
rect 2335 2354 2339 2355
rect 2335 2349 2339 2350
rect 2503 2354 2507 2355
rect 2503 2349 2507 2350
rect 2543 2354 2547 2355
rect 2543 2349 2547 2350
rect 2743 2354 2747 2355
rect 2743 2349 2747 2350
rect 2767 2354 2771 2355
rect 2767 2349 2771 2350
rect 2935 2354 2939 2355
rect 2935 2349 2939 2350
rect 3007 2354 3011 2355
rect 3007 2349 3011 2350
rect 3127 2354 3131 2355
rect 3127 2349 3131 2350
rect 3239 2354 3243 2355
rect 3239 2349 3243 2350
rect 3311 2354 3315 2355
rect 3311 2349 3315 2350
rect 3471 2354 3475 2355
rect 3471 2349 3475 2350
rect 3495 2354 3499 2355
rect 3495 2349 3499 2350
rect 3679 2354 3683 2355
rect 3679 2349 3683 2350
rect 2504 2325 2506 2349
rect 2768 2325 2770 2349
rect 3008 2325 3010 2349
rect 3240 2325 3242 2349
rect 3472 2325 3474 2349
rect 3680 2325 3682 2349
rect 2502 2324 2508 2325
rect 2502 2320 2503 2324
rect 2507 2320 2508 2324
rect 2502 2319 2508 2320
rect 2766 2324 2772 2325
rect 2766 2320 2767 2324
rect 2771 2320 2772 2324
rect 2766 2319 2772 2320
rect 3006 2324 3012 2325
rect 3006 2320 3007 2324
rect 3011 2320 3012 2324
rect 3006 2319 3012 2320
rect 3238 2324 3244 2325
rect 3238 2320 3239 2324
rect 3243 2320 3244 2324
rect 3238 2319 3244 2320
rect 3470 2324 3476 2325
rect 3470 2320 3471 2324
rect 3475 2320 3476 2324
rect 3470 2319 3476 2320
rect 3678 2324 3684 2325
rect 3678 2320 3679 2324
rect 3683 2320 3684 2324
rect 3678 2319 3684 2320
rect 2474 2309 2480 2310
rect 2474 2305 2475 2309
rect 2479 2305 2480 2309
rect 2474 2304 2480 2305
rect 2738 2309 2744 2310
rect 2738 2305 2739 2309
rect 2743 2305 2744 2309
rect 2738 2304 2744 2305
rect 2978 2309 2984 2310
rect 2978 2305 2979 2309
rect 2983 2305 2984 2309
rect 2978 2304 2984 2305
rect 3210 2309 3216 2310
rect 3210 2305 3211 2309
rect 3215 2305 3216 2309
rect 3210 2304 3216 2305
rect 3442 2309 3448 2310
rect 3442 2305 3443 2309
rect 3447 2305 3448 2309
rect 3442 2304 3448 2305
rect 3650 2309 3656 2310
rect 3650 2305 3651 2309
rect 3655 2305 3656 2309
rect 3650 2304 3656 2305
rect 2298 2299 2304 2300
rect 2298 2295 2299 2299
rect 2303 2295 2304 2299
rect 2298 2294 2304 2295
rect 2334 2299 2340 2300
rect 2334 2295 2335 2299
rect 2339 2295 2340 2299
rect 2334 2294 2340 2295
rect 2336 2268 2338 2294
rect 2334 2267 2340 2268
rect 2334 2263 2335 2267
rect 2339 2263 2340 2267
rect 2334 2262 2340 2263
rect 2476 2243 2478 2304
rect 2562 2267 2568 2268
rect 2562 2263 2563 2267
rect 2567 2263 2568 2267
rect 2562 2262 2568 2263
rect 1975 2242 1979 2243
rect 1975 2237 1979 2238
rect 1995 2242 1999 2243
rect 1995 2237 1999 2238
rect 2155 2242 2159 2243
rect 2155 2237 2159 2238
rect 2195 2242 2199 2243
rect 2195 2237 2199 2238
rect 2387 2242 2391 2243
rect 2387 2237 2391 2238
rect 2475 2242 2479 2243
rect 2475 2237 2479 2238
rect 1976 2177 1978 2237
rect 1974 2176 1980 2177
rect 1996 2176 1998 2237
rect 2122 2219 2128 2220
rect 2122 2215 2123 2219
rect 2127 2215 2128 2219
rect 2122 2214 2128 2215
rect 2124 2184 2126 2214
rect 2122 2183 2128 2184
rect 2122 2179 2123 2183
rect 2127 2179 2128 2183
rect 2122 2178 2128 2179
rect 2156 2176 2158 2237
rect 2388 2176 2390 2237
rect 2514 2219 2520 2220
rect 2514 2215 2515 2219
rect 2519 2215 2520 2219
rect 2514 2214 2520 2215
rect 2516 2184 2518 2214
rect 2564 2192 2566 2262
rect 2740 2243 2742 2304
rect 2826 2291 2832 2292
rect 2826 2287 2827 2291
rect 2831 2287 2832 2291
rect 2826 2286 2832 2287
rect 2828 2268 2830 2286
rect 2826 2267 2832 2268
rect 2826 2263 2827 2267
rect 2831 2263 2832 2267
rect 2826 2262 2832 2263
rect 2980 2243 2982 2304
rect 2994 2299 3000 2300
rect 2994 2295 2995 2299
rect 2999 2295 3000 2299
rect 2994 2294 3000 2295
rect 2996 2268 2998 2294
rect 2994 2267 3000 2268
rect 2994 2263 2995 2267
rect 2999 2263 3000 2267
rect 2994 2262 3000 2263
rect 3212 2243 3214 2304
rect 3226 2299 3232 2300
rect 3226 2295 3227 2299
rect 3231 2295 3232 2299
rect 3226 2294 3232 2295
rect 3228 2268 3230 2294
rect 3226 2267 3232 2268
rect 3226 2263 3227 2267
rect 3231 2263 3232 2267
rect 3226 2262 3232 2263
rect 3444 2243 3446 2304
rect 3458 2299 3464 2300
rect 3458 2295 3459 2299
rect 3463 2295 3464 2299
rect 3458 2294 3464 2295
rect 3460 2268 3462 2294
rect 3458 2267 3464 2268
rect 3458 2263 3459 2267
rect 3463 2263 3464 2267
rect 3458 2262 3464 2263
rect 3652 2243 3654 2304
rect 3666 2299 3672 2300
rect 3666 2295 3667 2299
rect 3671 2295 3672 2299
rect 3666 2294 3672 2295
rect 3668 2268 3670 2294
rect 3740 2292 3742 2410
rect 3800 2409 3802 2469
rect 3840 2439 3842 2515
rect 4468 2439 4470 2516
rect 4604 2439 4606 2516
rect 4618 2511 4624 2512
rect 4618 2507 4619 2511
rect 4623 2507 4624 2511
rect 4618 2506 4624 2507
rect 4620 2480 4622 2506
rect 4618 2479 4624 2480
rect 4618 2475 4619 2479
rect 4623 2475 4624 2479
rect 4618 2474 4624 2475
rect 4740 2439 4742 2516
rect 4754 2511 4760 2512
rect 4754 2507 4755 2511
rect 4759 2507 4760 2511
rect 4754 2506 4760 2507
rect 4756 2480 4758 2506
rect 4818 2503 4824 2504
rect 4818 2499 4819 2503
rect 4823 2499 4824 2503
rect 4818 2498 4824 2499
rect 4754 2479 4760 2480
rect 4754 2475 4755 2479
rect 4759 2475 4760 2479
rect 4754 2474 4760 2475
rect 3839 2438 3843 2439
rect 3839 2433 3843 2434
rect 4467 2438 4471 2439
rect 4467 2433 4471 2434
rect 4603 2438 4607 2439
rect 4603 2433 4607 2434
rect 4699 2438 4703 2439
rect 4699 2433 4703 2434
rect 4739 2438 4743 2439
rect 4739 2433 4743 2434
rect 3798 2408 3804 2409
rect 3798 2404 3799 2408
rect 3803 2404 3804 2408
rect 3798 2403 3804 2404
rect 3798 2391 3804 2392
rect 3798 2387 3799 2391
rect 3803 2387 3804 2391
rect 3798 2386 3804 2387
rect 3800 2355 3802 2386
rect 3840 2373 3842 2433
rect 3838 2372 3844 2373
rect 4700 2372 4702 2433
rect 4820 2416 4822 2498
rect 4876 2439 4878 2516
rect 4890 2511 4896 2512
rect 4890 2507 4891 2511
rect 4895 2507 4896 2511
rect 4890 2506 4896 2507
rect 4892 2480 4894 2506
rect 5000 2496 5002 2618
rect 5012 2616 5014 2677
rect 5276 2616 5278 2677
rect 5340 2624 5342 2890
rect 5412 2864 5414 2966
rect 5515 2922 5519 2923
rect 5515 2917 5519 2918
rect 5410 2863 5416 2864
rect 5410 2859 5411 2863
rect 5415 2859 5416 2863
rect 5410 2858 5416 2859
rect 5516 2856 5518 2917
rect 5620 2900 5622 3106
rect 5664 3105 5666 3165
rect 5662 3104 5668 3105
rect 5662 3100 5663 3104
rect 5667 3100 5668 3104
rect 5662 3099 5668 3100
rect 5662 3087 5668 3088
rect 5662 3083 5663 3087
rect 5667 3083 5668 3087
rect 5662 3082 5668 3083
rect 5664 3059 5666 3082
rect 5663 3058 5667 3059
rect 5663 3053 5667 3054
rect 5664 3030 5666 3053
rect 5662 3029 5668 3030
rect 5662 3025 5663 3029
rect 5667 3025 5668 3029
rect 5662 3024 5668 3025
rect 5662 3012 5668 3013
rect 5662 3008 5663 3012
rect 5667 3008 5668 3012
rect 5662 3007 5668 3008
rect 5664 2923 5666 3007
rect 5663 2922 5667 2923
rect 5663 2917 5667 2918
rect 5618 2899 5624 2900
rect 5618 2895 5619 2899
rect 5623 2895 5624 2899
rect 5618 2894 5624 2895
rect 5618 2863 5624 2864
rect 5618 2859 5619 2863
rect 5623 2859 5624 2863
rect 5618 2858 5624 2859
rect 5514 2855 5520 2856
rect 5514 2851 5515 2855
rect 5519 2851 5520 2855
rect 5514 2850 5520 2851
rect 5542 2840 5548 2841
rect 5542 2836 5543 2840
rect 5547 2836 5548 2840
rect 5542 2835 5548 2836
rect 5544 2807 5546 2835
rect 5543 2806 5547 2807
rect 5543 2801 5547 2802
rect 5515 2682 5519 2683
rect 5515 2677 5519 2678
rect 5398 2659 5404 2660
rect 5398 2655 5399 2659
rect 5403 2655 5404 2659
rect 5398 2654 5404 2655
rect 5338 2623 5344 2624
rect 5338 2619 5339 2623
rect 5343 2619 5344 2623
rect 5338 2618 5344 2619
rect 5010 2615 5016 2616
rect 5010 2611 5011 2615
rect 5015 2611 5016 2615
rect 5010 2610 5016 2611
rect 5274 2615 5280 2616
rect 5274 2611 5275 2615
rect 5279 2611 5280 2615
rect 5274 2610 5280 2611
rect 5038 2600 5044 2601
rect 5038 2596 5039 2600
rect 5043 2596 5044 2600
rect 5038 2595 5044 2596
rect 5302 2600 5308 2601
rect 5302 2596 5303 2600
rect 5307 2596 5308 2600
rect 5302 2595 5308 2596
rect 5040 2567 5042 2595
rect 5304 2567 5306 2595
rect 5039 2566 5043 2567
rect 5039 2561 5043 2562
rect 5303 2566 5307 2567
rect 5303 2561 5307 2562
rect 5040 2537 5042 2561
rect 5038 2536 5044 2537
rect 5038 2532 5039 2536
rect 5043 2532 5044 2536
rect 5038 2531 5044 2532
rect 5010 2521 5016 2522
rect 5010 2517 5011 2521
rect 5015 2517 5016 2521
rect 5010 2516 5016 2517
rect 4998 2495 5004 2496
rect 4998 2491 4999 2495
rect 5003 2491 5004 2495
rect 4998 2490 5004 2491
rect 4890 2479 4896 2480
rect 4890 2475 4891 2479
rect 4895 2475 4896 2479
rect 4890 2474 4896 2475
rect 5012 2439 5014 2516
rect 5026 2511 5032 2512
rect 5026 2507 5027 2511
rect 5031 2507 5032 2511
rect 5026 2506 5032 2507
rect 5028 2480 5030 2506
rect 5026 2479 5032 2480
rect 5026 2475 5027 2479
rect 5031 2475 5032 2479
rect 5026 2474 5032 2475
rect 4835 2438 4839 2439
rect 4835 2433 4839 2434
rect 4875 2438 4879 2439
rect 4875 2433 4879 2434
rect 4971 2438 4975 2439
rect 4971 2433 4975 2434
rect 5011 2438 5015 2439
rect 5011 2433 5015 2434
rect 5107 2438 5111 2439
rect 5107 2433 5111 2434
rect 5243 2438 5247 2439
rect 5243 2433 5247 2434
rect 5379 2438 5383 2439
rect 5379 2433 5383 2434
rect 4818 2415 4824 2416
rect 4818 2411 4819 2415
rect 4823 2411 4824 2415
rect 4818 2410 4824 2411
rect 4826 2415 4832 2416
rect 4826 2411 4827 2415
rect 4831 2411 4832 2415
rect 4826 2410 4832 2411
rect 4828 2380 4830 2410
rect 4826 2379 4832 2380
rect 4826 2375 4827 2379
rect 4831 2375 4832 2379
rect 4826 2374 4832 2375
rect 4836 2372 4838 2433
rect 4972 2372 4974 2433
rect 5108 2372 5110 2433
rect 5244 2372 5246 2433
rect 5370 2379 5376 2380
rect 5370 2375 5371 2379
rect 5375 2375 5376 2379
rect 5370 2374 5376 2375
rect 3838 2368 3839 2372
rect 3843 2368 3844 2372
rect 3838 2367 3844 2368
rect 4698 2371 4704 2372
rect 4698 2367 4699 2371
rect 4703 2367 4704 2371
rect 4698 2366 4704 2367
rect 4834 2371 4840 2372
rect 4834 2367 4835 2371
rect 4839 2367 4840 2371
rect 4834 2366 4840 2367
rect 4970 2371 4976 2372
rect 4970 2367 4971 2371
rect 4975 2367 4976 2371
rect 4970 2366 4976 2367
rect 5106 2371 5112 2372
rect 5106 2367 5107 2371
rect 5111 2367 5112 2371
rect 5106 2366 5112 2367
rect 5242 2371 5248 2372
rect 5242 2367 5243 2371
rect 5247 2367 5248 2371
rect 5242 2366 5248 2367
rect 4726 2356 4732 2357
rect 3838 2355 3844 2356
rect 3799 2354 3803 2355
rect 3838 2351 3839 2355
rect 3843 2351 3844 2355
rect 4726 2352 4727 2356
rect 4731 2352 4732 2356
rect 4726 2351 4732 2352
rect 4862 2356 4868 2357
rect 4862 2352 4863 2356
rect 4867 2352 4868 2356
rect 4862 2351 4868 2352
rect 4998 2356 5004 2357
rect 4998 2352 4999 2356
rect 5003 2352 5004 2356
rect 4998 2351 5004 2352
rect 5134 2356 5140 2357
rect 5134 2352 5135 2356
rect 5139 2352 5140 2356
rect 5134 2351 5140 2352
rect 5270 2356 5276 2357
rect 5270 2352 5271 2356
rect 5275 2352 5276 2356
rect 5270 2351 5276 2352
rect 3838 2350 3844 2351
rect 3799 2349 3803 2350
rect 3800 2326 3802 2349
rect 3798 2325 3804 2326
rect 3798 2321 3799 2325
rect 3803 2321 3804 2325
rect 3798 2320 3804 2321
rect 3840 2315 3842 2350
rect 4728 2315 4730 2351
rect 4864 2315 4866 2351
rect 5000 2315 5002 2351
rect 5136 2315 5138 2351
rect 5272 2315 5274 2351
rect 3839 2314 3843 2315
rect 3839 2309 3843 2310
rect 3887 2314 3891 2315
rect 3887 2309 3891 2310
rect 4183 2314 4187 2315
rect 4183 2309 4187 2310
rect 4495 2314 4499 2315
rect 4495 2309 4499 2310
rect 4727 2314 4731 2315
rect 4727 2309 4731 2310
rect 4791 2314 4795 2315
rect 4791 2309 4795 2310
rect 4863 2314 4867 2315
rect 4863 2309 4867 2310
rect 4999 2314 5003 2315
rect 4999 2309 5003 2310
rect 5087 2314 5091 2315
rect 5087 2309 5091 2310
rect 5135 2314 5139 2315
rect 5135 2309 5139 2310
rect 5271 2314 5275 2315
rect 5271 2309 5275 2310
rect 3798 2308 3804 2309
rect 3798 2304 3799 2308
rect 3803 2304 3804 2308
rect 3798 2303 3804 2304
rect 3754 2299 3760 2300
rect 3754 2295 3755 2299
rect 3759 2295 3760 2299
rect 3754 2294 3760 2295
rect 3738 2291 3744 2292
rect 3738 2287 3739 2291
rect 3743 2287 3744 2291
rect 3738 2286 3744 2287
rect 3666 2267 3672 2268
rect 3666 2263 3667 2267
rect 3671 2263 3672 2267
rect 3666 2262 3672 2263
rect 2667 2242 2671 2243
rect 2667 2237 2671 2238
rect 2739 2242 2743 2243
rect 2739 2237 2743 2238
rect 2979 2242 2983 2243
rect 2979 2237 2983 2238
rect 2987 2242 2991 2243
rect 2987 2237 2991 2238
rect 3211 2242 3215 2243
rect 3211 2237 3215 2238
rect 3331 2242 3335 2243
rect 3331 2237 3335 2238
rect 3443 2242 3447 2243
rect 3443 2237 3447 2238
rect 3651 2242 3655 2243
rect 3651 2237 3655 2238
rect 2562 2191 2568 2192
rect 2562 2187 2563 2191
rect 2567 2187 2568 2191
rect 2562 2186 2568 2187
rect 2514 2183 2520 2184
rect 2514 2179 2515 2183
rect 2519 2179 2520 2183
rect 2514 2178 2520 2179
rect 2668 2176 2670 2237
rect 2794 2219 2800 2220
rect 2794 2215 2795 2219
rect 2799 2215 2800 2219
rect 2794 2214 2800 2215
rect 2796 2184 2798 2214
rect 2794 2183 2800 2184
rect 2794 2179 2795 2183
rect 2799 2179 2800 2183
rect 2794 2178 2800 2179
rect 2988 2176 2990 2237
rect 3114 2219 3120 2220
rect 3114 2215 3115 2219
rect 3119 2215 3120 2219
rect 3114 2214 3120 2215
rect 3116 2184 3118 2214
rect 3114 2183 3120 2184
rect 3114 2179 3115 2183
rect 3119 2179 3120 2183
rect 3114 2178 3120 2179
rect 3332 2176 3334 2237
rect 3652 2176 3654 2237
rect 3756 2220 3758 2294
rect 3800 2243 3802 2303
rect 3840 2286 3842 2309
rect 3838 2285 3844 2286
rect 3888 2285 3890 2309
rect 4184 2285 4186 2309
rect 4496 2285 4498 2309
rect 4792 2285 4794 2309
rect 5088 2285 5090 2309
rect 3838 2281 3839 2285
rect 3843 2281 3844 2285
rect 3838 2280 3844 2281
rect 3886 2284 3892 2285
rect 3886 2280 3887 2284
rect 3891 2280 3892 2284
rect 3886 2279 3892 2280
rect 4182 2284 4188 2285
rect 4182 2280 4183 2284
rect 4187 2280 4188 2284
rect 4182 2279 4188 2280
rect 4494 2284 4500 2285
rect 4494 2280 4495 2284
rect 4499 2280 4500 2284
rect 4494 2279 4500 2280
rect 4790 2284 4796 2285
rect 4790 2280 4791 2284
rect 4795 2280 4796 2284
rect 4790 2279 4796 2280
rect 5086 2284 5092 2285
rect 5086 2280 5087 2284
rect 5091 2280 5092 2284
rect 5086 2279 5092 2280
rect 3858 2269 3864 2270
rect 3838 2268 3844 2269
rect 3838 2264 3839 2268
rect 3843 2264 3844 2268
rect 3858 2265 3859 2269
rect 3863 2265 3864 2269
rect 3858 2264 3864 2265
rect 4154 2269 4160 2270
rect 4154 2265 4155 2269
rect 4159 2265 4160 2269
rect 4154 2264 4160 2265
rect 4466 2269 4472 2270
rect 4466 2265 4467 2269
rect 4471 2265 4472 2269
rect 4466 2264 4472 2265
rect 4762 2269 4768 2270
rect 4762 2265 4763 2269
rect 4767 2265 4768 2269
rect 4762 2264 4768 2265
rect 5058 2269 5064 2270
rect 5058 2265 5059 2269
rect 5063 2265 5064 2269
rect 5058 2264 5064 2265
rect 5354 2269 5360 2270
rect 5354 2265 5355 2269
rect 5359 2265 5360 2269
rect 5354 2264 5360 2265
rect 3838 2263 3844 2264
rect 3799 2242 3803 2243
rect 3799 2237 3803 2238
rect 3778 2227 3784 2228
rect 3778 2223 3779 2227
rect 3783 2223 3784 2227
rect 3778 2222 3784 2223
rect 3754 2219 3760 2220
rect 3754 2215 3755 2219
rect 3759 2215 3760 2219
rect 3754 2214 3760 2215
rect 3780 2184 3782 2222
rect 3778 2183 3784 2184
rect 3778 2179 3779 2183
rect 3783 2179 3784 2183
rect 3778 2178 3784 2179
rect 3800 2177 3802 2237
rect 3840 2199 3842 2263
rect 3860 2199 3862 2264
rect 3962 2259 3968 2260
rect 3962 2255 3963 2259
rect 3967 2255 3968 2259
rect 3962 2254 3968 2255
rect 3839 2198 3843 2199
rect 3839 2193 3843 2194
rect 3859 2198 3863 2199
rect 3859 2193 3863 2194
rect 3798 2176 3804 2177
rect 1974 2172 1975 2176
rect 1979 2172 1980 2176
rect 1974 2171 1980 2172
rect 1994 2175 2000 2176
rect 1994 2171 1995 2175
rect 1999 2171 2000 2175
rect 1387 2170 1391 2171
rect 1387 2165 1391 2166
rect 1467 2170 1471 2171
rect 1467 2165 1471 2166
rect 1635 2170 1639 2171
rect 1635 2165 1639 2166
rect 1787 2170 1791 2171
rect 1787 2165 1791 2166
rect 1935 2170 1939 2171
rect 1994 2170 2000 2171
rect 2154 2175 2160 2176
rect 2154 2171 2155 2175
rect 2159 2171 2160 2175
rect 2154 2170 2160 2171
rect 2386 2175 2392 2176
rect 2386 2171 2387 2175
rect 2391 2171 2392 2175
rect 2386 2170 2392 2171
rect 2666 2175 2672 2176
rect 2666 2171 2667 2175
rect 2671 2171 2672 2175
rect 2666 2170 2672 2171
rect 2986 2175 2992 2176
rect 2986 2171 2987 2175
rect 2991 2171 2992 2175
rect 2986 2170 2992 2171
rect 3330 2175 3336 2176
rect 3330 2171 3331 2175
rect 3335 2171 3336 2175
rect 3330 2170 3336 2171
rect 3650 2175 3656 2176
rect 3650 2171 3651 2175
rect 3655 2171 3656 2175
rect 3798 2172 3799 2176
rect 3803 2172 3804 2176
rect 3798 2171 3804 2172
rect 3650 2170 3656 2171
rect 1935 2165 1939 2166
rect 1274 2111 1280 2112
rect 1274 2107 1275 2111
rect 1279 2107 1280 2111
rect 1274 2106 1280 2107
rect 1388 2104 1390 2165
rect 1614 2147 1620 2148
rect 1614 2143 1615 2147
rect 1619 2143 1620 2147
rect 1614 2142 1620 2143
rect 1626 2147 1632 2148
rect 1626 2143 1627 2147
rect 1631 2143 1632 2147
rect 1626 2142 1632 2143
rect 1616 2112 1618 2142
rect 1458 2111 1464 2112
rect 1458 2107 1459 2111
rect 1463 2107 1464 2111
rect 1458 2106 1464 2107
rect 1614 2111 1620 2112
rect 1614 2107 1615 2111
rect 1619 2107 1620 2111
rect 1614 2106 1620 2107
rect 1146 2103 1152 2104
rect 1146 2099 1147 2103
rect 1151 2099 1152 2103
rect 1146 2098 1152 2099
rect 1386 2103 1392 2104
rect 1386 2099 1387 2103
rect 1391 2099 1392 2103
rect 1386 2098 1392 2099
rect 1174 2088 1180 2089
rect 1174 2084 1175 2088
rect 1179 2084 1180 2088
rect 1174 2083 1180 2084
rect 1414 2088 1420 2089
rect 1414 2084 1415 2088
rect 1419 2084 1420 2088
rect 1414 2083 1420 2084
rect 1176 2055 1178 2083
rect 1416 2055 1418 2083
rect 1111 2054 1115 2055
rect 1111 2049 1115 2050
rect 1175 2054 1179 2055
rect 1175 2049 1179 2050
rect 1255 2054 1259 2055
rect 1255 2049 1259 2050
rect 1399 2054 1403 2055
rect 1399 2049 1403 2050
rect 1415 2054 1419 2055
rect 1415 2049 1419 2050
rect 1112 2025 1114 2049
rect 1256 2025 1258 2049
rect 1400 2025 1402 2049
rect 1110 2024 1116 2025
rect 1110 2020 1111 2024
rect 1115 2020 1116 2024
rect 1110 2019 1116 2020
rect 1254 2024 1260 2025
rect 1254 2020 1255 2024
rect 1259 2020 1260 2024
rect 1254 2019 1260 2020
rect 1398 2024 1404 2025
rect 1398 2020 1399 2024
rect 1403 2020 1404 2024
rect 1398 2019 1404 2020
rect 1082 2009 1088 2010
rect 1082 2005 1083 2009
rect 1087 2005 1088 2009
rect 1082 2004 1088 2005
rect 1226 2009 1232 2010
rect 1226 2005 1227 2009
rect 1231 2005 1232 2009
rect 1226 2004 1232 2005
rect 1370 2009 1376 2010
rect 1370 2005 1371 2009
rect 1375 2005 1376 2009
rect 1370 2004 1376 2005
rect 954 1999 960 2000
rect 954 1995 955 1999
rect 959 1995 960 1999
rect 954 1994 960 1995
rect 1002 1999 1008 2000
rect 1002 1995 1003 1999
rect 1007 1995 1008 1999
rect 1002 1994 1008 1995
rect 956 1968 958 1994
rect 954 1967 960 1968
rect 954 1963 955 1967
rect 959 1963 960 1967
rect 954 1962 960 1963
rect 1084 1931 1086 2004
rect 1228 1931 1230 2004
rect 1372 1931 1374 2004
rect 1460 1968 1462 2106
rect 1543 2054 1547 2055
rect 1543 2049 1547 2050
rect 1544 2025 1546 2049
rect 1542 2024 1548 2025
rect 1542 2020 1543 2024
rect 1547 2020 1548 2024
rect 1542 2019 1548 2020
rect 1514 2009 1520 2010
rect 1514 2005 1515 2009
rect 1519 2005 1520 2009
rect 1514 2004 1520 2005
rect 1458 1967 1464 1968
rect 1458 1963 1459 1967
rect 1463 1963 1464 1967
rect 1458 1962 1464 1963
rect 1516 1931 1518 2004
rect 1628 2000 1630 2142
rect 1636 2104 1638 2165
rect 1936 2105 1938 2165
rect 2022 2160 2028 2161
rect 1974 2159 1980 2160
rect 1974 2155 1975 2159
rect 1979 2155 1980 2159
rect 2022 2156 2023 2160
rect 2027 2156 2028 2160
rect 2022 2155 2028 2156
rect 2182 2160 2188 2161
rect 2182 2156 2183 2160
rect 2187 2156 2188 2160
rect 2182 2155 2188 2156
rect 2414 2160 2420 2161
rect 2414 2156 2415 2160
rect 2419 2156 2420 2160
rect 2414 2155 2420 2156
rect 2694 2160 2700 2161
rect 2694 2156 2695 2160
rect 2699 2156 2700 2160
rect 2694 2155 2700 2156
rect 3014 2160 3020 2161
rect 3014 2156 3015 2160
rect 3019 2156 3020 2160
rect 3014 2155 3020 2156
rect 3358 2160 3364 2161
rect 3358 2156 3359 2160
rect 3363 2156 3364 2160
rect 3358 2155 3364 2156
rect 3678 2160 3684 2161
rect 3678 2156 3679 2160
rect 3683 2156 3684 2160
rect 3678 2155 3684 2156
rect 3798 2159 3804 2160
rect 3798 2155 3799 2159
rect 3803 2155 3804 2159
rect 1974 2154 1980 2155
rect 1934 2104 1940 2105
rect 1634 2103 1640 2104
rect 1634 2099 1635 2103
rect 1639 2099 1640 2103
rect 1934 2100 1935 2104
rect 1939 2100 1940 2104
rect 1934 2099 1940 2100
rect 1634 2098 1640 2099
rect 1662 2088 1668 2089
rect 1662 2084 1663 2088
rect 1667 2084 1668 2088
rect 1662 2083 1668 2084
rect 1934 2087 1940 2088
rect 1934 2083 1935 2087
rect 1939 2083 1940 2087
rect 1664 2055 1666 2083
rect 1934 2082 1940 2083
rect 1936 2055 1938 2082
rect 1663 2054 1667 2055
rect 1663 2049 1667 2050
rect 1679 2054 1683 2055
rect 1679 2049 1683 2050
rect 1815 2054 1819 2055
rect 1815 2049 1819 2050
rect 1935 2054 1939 2055
rect 1935 2049 1939 2050
rect 1680 2025 1682 2049
rect 1816 2025 1818 2049
rect 1936 2026 1938 2049
rect 1934 2025 1940 2026
rect 1678 2024 1684 2025
rect 1678 2020 1679 2024
rect 1683 2020 1684 2024
rect 1678 2019 1684 2020
rect 1814 2024 1820 2025
rect 1814 2020 1815 2024
rect 1819 2020 1820 2024
rect 1934 2021 1935 2025
rect 1939 2021 1940 2025
rect 1934 2020 1940 2021
rect 1814 2019 1820 2020
rect 1650 2009 1656 2010
rect 1650 2005 1651 2009
rect 1655 2005 1656 2009
rect 1650 2004 1656 2005
rect 1786 2009 1792 2010
rect 1786 2005 1787 2009
rect 1791 2005 1792 2009
rect 1786 2004 1792 2005
rect 1934 2008 1940 2009
rect 1934 2004 1935 2008
rect 1939 2004 1940 2008
rect 1626 1999 1632 2000
rect 1626 1995 1627 1999
rect 1631 1995 1632 1999
rect 1626 1994 1632 1995
rect 1602 1991 1608 1992
rect 1602 1987 1603 1991
rect 1607 1987 1608 1991
rect 1602 1986 1608 1987
rect 1604 1968 1606 1986
rect 1602 1967 1608 1968
rect 1602 1963 1603 1967
rect 1607 1963 1608 1967
rect 1602 1962 1608 1963
rect 1652 1931 1654 2004
rect 1738 1967 1744 1968
rect 1738 1963 1739 1967
rect 1743 1963 1744 1967
rect 1738 1962 1744 1963
rect 939 1930 943 1931
rect 939 1925 943 1926
rect 987 1930 991 1931
rect 987 1925 991 1926
rect 1083 1930 1087 1931
rect 1083 1925 1087 1926
rect 1155 1930 1159 1931
rect 1155 1925 1159 1926
rect 1227 1930 1231 1931
rect 1227 1925 1231 1926
rect 1323 1930 1327 1931
rect 1323 1925 1327 1926
rect 1371 1930 1375 1931
rect 1371 1925 1375 1926
rect 1483 1930 1487 1931
rect 1483 1925 1487 1926
rect 1515 1930 1519 1931
rect 1515 1925 1519 1926
rect 1643 1930 1647 1931
rect 1643 1925 1647 1926
rect 1651 1930 1655 1931
rect 1651 1925 1655 1926
rect 930 1907 936 1908
rect 930 1903 931 1907
rect 935 1903 936 1907
rect 930 1902 936 1903
rect 938 1907 944 1908
rect 938 1903 939 1907
rect 943 1903 944 1907
rect 938 1902 944 1903
rect 940 1872 942 1902
rect 938 1871 944 1872
rect 938 1867 939 1871
rect 943 1867 944 1871
rect 938 1866 944 1867
rect 988 1864 990 1925
rect 1114 1907 1120 1908
rect 1114 1903 1115 1907
rect 1119 1903 1120 1907
rect 1114 1902 1120 1903
rect 1116 1872 1118 1902
rect 1114 1871 1120 1872
rect 1114 1867 1115 1871
rect 1119 1867 1120 1871
rect 1114 1866 1120 1867
rect 1156 1864 1158 1925
rect 1324 1864 1326 1925
rect 1450 1907 1456 1908
rect 1410 1903 1416 1904
rect 1410 1899 1411 1903
rect 1415 1899 1416 1903
rect 1450 1903 1451 1907
rect 1455 1903 1456 1907
rect 1450 1902 1456 1903
rect 1410 1898 1416 1899
rect 1412 1880 1414 1898
rect 1410 1879 1416 1880
rect 1410 1875 1411 1879
rect 1415 1875 1416 1879
rect 1410 1874 1416 1875
rect 1452 1872 1454 1902
rect 1378 1871 1384 1872
rect 1378 1867 1379 1871
rect 1383 1867 1384 1871
rect 1378 1866 1384 1867
rect 1450 1871 1456 1872
rect 1450 1867 1451 1871
rect 1455 1867 1456 1871
rect 1450 1866 1456 1867
rect 434 1863 440 1864
rect 434 1859 435 1863
rect 439 1859 440 1863
rect 434 1858 440 1859
rect 626 1863 632 1864
rect 626 1859 627 1863
rect 631 1859 632 1863
rect 626 1858 632 1859
rect 810 1863 816 1864
rect 810 1859 811 1863
rect 815 1859 816 1863
rect 810 1858 816 1859
rect 986 1863 992 1864
rect 986 1859 987 1863
rect 991 1859 992 1863
rect 986 1858 992 1859
rect 1154 1863 1160 1864
rect 1154 1859 1155 1863
rect 1159 1859 1160 1863
rect 1154 1858 1160 1859
rect 1322 1863 1328 1864
rect 1322 1859 1323 1863
rect 1327 1859 1328 1863
rect 1322 1858 1328 1859
rect 462 1848 468 1849
rect 462 1844 463 1848
rect 467 1844 468 1848
rect 462 1843 468 1844
rect 654 1848 660 1849
rect 654 1844 655 1848
rect 659 1844 660 1848
rect 654 1843 660 1844
rect 838 1848 844 1849
rect 838 1844 839 1848
rect 843 1844 844 1848
rect 838 1843 844 1844
rect 1014 1848 1020 1849
rect 1014 1844 1015 1848
rect 1019 1844 1020 1848
rect 1014 1843 1020 1844
rect 1182 1848 1188 1849
rect 1182 1844 1183 1848
rect 1187 1844 1188 1848
rect 1182 1843 1188 1844
rect 1350 1848 1356 1849
rect 1350 1844 1351 1848
rect 1355 1844 1356 1848
rect 1350 1843 1356 1844
rect 464 1807 466 1843
rect 656 1807 658 1843
rect 840 1807 842 1843
rect 1016 1807 1018 1843
rect 1184 1807 1186 1843
rect 1352 1807 1354 1843
rect 463 1806 467 1807
rect 463 1801 467 1802
rect 655 1806 659 1807
rect 655 1801 659 1802
rect 695 1806 699 1807
rect 695 1801 699 1802
rect 839 1806 843 1807
rect 839 1801 843 1802
rect 927 1806 931 1807
rect 927 1801 931 1802
rect 1015 1806 1019 1807
rect 1015 1801 1019 1802
rect 1159 1806 1163 1807
rect 1159 1801 1163 1802
rect 1183 1806 1187 1807
rect 1183 1801 1187 1802
rect 1351 1806 1355 1807
rect 1351 1801 1355 1802
rect 464 1777 466 1801
rect 696 1777 698 1801
rect 928 1777 930 1801
rect 1160 1777 1162 1801
rect 462 1776 468 1777
rect 462 1772 463 1776
rect 467 1772 468 1776
rect 462 1771 468 1772
rect 694 1776 700 1777
rect 694 1772 695 1776
rect 699 1772 700 1776
rect 694 1771 700 1772
rect 926 1776 932 1777
rect 926 1772 927 1776
rect 931 1772 932 1776
rect 926 1771 932 1772
rect 1158 1776 1164 1777
rect 1158 1772 1159 1776
rect 1163 1772 1164 1776
rect 1158 1771 1164 1772
rect 434 1761 440 1762
rect 434 1757 435 1761
rect 439 1757 440 1761
rect 434 1756 440 1757
rect 666 1761 672 1762
rect 666 1757 667 1761
rect 671 1757 672 1761
rect 666 1756 672 1757
rect 898 1761 904 1762
rect 898 1757 899 1761
rect 903 1757 904 1761
rect 898 1756 904 1757
rect 1130 1761 1136 1762
rect 1130 1757 1131 1761
rect 1135 1757 1136 1761
rect 1130 1756 1136 1757
rect 1362 1761 1368 1762
rect 1362 1757 1363 1761
rect 1367 1757 1368 1761
rect 1362 1756 1368 1757
rect 322 1751 328 1752
rect 322 1747 323 1751
rect 327 1747 328 1751
rect 322 1746 328 1747
rect 436 1683 438 1756
rect 486 1719 492 1720
rect 486 1715 487 1719
rect 491 1715 492 1719
rect 486 1714 492 1715
rect 111 1682 115 1683
rect 111 1677 115 1678
rect 131 1682 135 1683
rect 131 1677 135 1678
rect 195 1682 199 1683
rect 195 1677 199 1678
rect 363 1682 367 1683
rect 363 1677 367 1678
rect 435 1682 439 1683
rect 435 1677 439 1678
rect 112 1617 114 1677
rect 110 1616 116 1617
rect 132 1616 134 1677
rect 258 1659 264 1660
rect 218 1655 224 1656
rect 218 1651 219 1655
rect 223 1651 224 1655
rect 258 1655 259 1659
rect 263 1655 264 1659
rect 258 1654 264 1655
rect 218 1650 224 1651
rect 110 1612 111 1616
rect 115 1612 116 1616
rect 110 1611 116 1612
rect 130 1615 136 1616
rect 130 1611 131 1615
rect 135 1611 136 1615
rect 130 1610 136 1611
rect 158 1600 164 1601
rect 110 1599 116 1600
rect 110 1595 111 1599
rect 115 1595 116 1599
rect 158 1596 159 1600
rect 163 1596 164 1600
rect 158 1595 164 1596
rect 110 1594 116 1595
rect 112 1559 114 1594
rect 160 1559 162 1595
rect 111 1558 115 1559
rect 111 1553 115 1554
rect 159 1558 163 1559
rect 159 1553 163 1554
rect 112 1530 114 1553
rect 110 1529 116 1530
rect 160 1529 162 1553
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 158 1528 164 1529
rect 158 1524 159 1528
rect 163 1524 164 1528
rect 158 1523 164 1524
rect 130 1513 136 1514
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 130 1509 131 1513
rect 135 1509 136 1513
rect 130 1508 136 1509
rect 110 1507 116 1508
rect 112 1435 114 1507
rect 132 1435 134 1508
rect 220 1504 222 1650
rect 260 1624 262 1654
rect 258 1623 264 1624
rect 258 1619 259 1623
rect 263 1619 264 1623
rect 258 1618 264 1619
rect 364 1616 366 1677
rect 488 1624 490 1714
rect 668 1683 670 1756
rect 754 1743 760 1744
rect 754 1739 755 1743
rect 759 1739 760 1743
rect 754 1738 760 1739
rect 756 1720 758 1738
rect 754 1719 760 1720
rect 754 1715 755 1719
rect 759 1715 760 1719
rect 754 1714 760 1715
rect 900 1683 902 1756
rect 914 1751 920 1752
rect 914 1747 915 1751
rect 919 1747 920 1751
rect 914 1746 920 1747
rect 916 1720 918 1746
rect 914 1719 920 1720
rect 914 1715 915 1719
rect 919 1715 920 1719
rect 914 1714 920 1715
rect 1132 1683 1134 1756
rect 1146 1751 1152 1752
rect 1146 1747 1147 1751
rect 1151 1747 1152 1751
rect 1146 1746 1152 1747
rect 1242 1751 1248 1752
rect 1242 1747 1243 1751
rect 1247 1747 1248 1751
rect 1242 1746 1248 1747
rect 1148 1720 1150 1746
rect 1146 1719 1152 1720
rect 1146 1715 1147 1719
rect 1151 1715 1152 1719
rect 1146 1714 1152 1715
rect 619 1682 623 1683
rect 619 1677 623 1678
rect 667 1682 671 1683
rect 667 1677 671 1678
rect 875 1682 879 1683
rect 875 1677 879 1678
rect 899 1682 903 1683
rect 899 1677 903 1678
rect 1131 1682 1135 1683
rect 1131 1677 1135 1678
rect 1139 1682 1143 1683
rect 1139 1677 1143 1678
rect 486 1623 492 1624
rect 486 1619 487 1623
rect 491 1619 492 1623
rect 486 1618 492 1619
rect 570 1623 576 1624
rect 570 1619 571 1623
rect 575 1619 576 1623
rect 570 1618 576 1619
rect 362 1615 368 1616
rect 362 1611 363 1615
rect 367 1611 368 1615
rect 362 1610 368 1611
rect 390 1600 396 1601
rect 390 1596 391 1600
rect 395 1596 396 1600
rect 390 1595 396 1596
rect 392 1559 394 1595
rect 327 1558 331 1559
rect 327 1553 331 1554
rect 391 1558 395 1559
rect 391 1553 395 1554
rect 511 1558 515 1559
rect 511 1553 515 1554
rect 328 1529 330 1553
rect 512 1529 514 1553
rect 326 1528 332 1529
rect 326 1524 327 1528
rect 331 1524 332 1528
rect 326 1523 332 1524
rect 510 1528 516 1529
rect 510 1524 511 1528
rect 515 1524 516 1528
rect 510 1523 516 1524
rect 298 1513 304 1514
rect 298 1509 299 1513
rect 303 1509 304 1513
rect 298 1508 304 1509
rect 482 1513 488 1514
rect 482 1509 483 1513
rect 487 1509 488 1513
rect 482 1508 488 1509
rect 218 1503 224 1504
rect 218 1499 219 1503
rect 223 1499 224 1503
rect 218 1498 224 1499
rect 286 1503 292 1504
rect 286 1499 287 1503
rect 291 1499 292 1503
rect 286 1498 292 1499
rect 288 1472 290 1498
rect 286 1471 292 1472
rect 286 1467 287 1471
rect 291 1467 292 1471
rect 286 1466 292 1467
rect 300 1435 302 1508
rect 386 1471 392 1472
rect 386 1467 387 1471
rect 391 1467 392 1471
rect 386 1466 392 1467
rect 111 1434 115 1435
rect 111 1429 115 1430
rect 131 1434 135 1435
rect 131 1429 135 1430
rect 299 1434 303 1435
rect 299 1429 303 1430
rect 112 1369 114 1429
rect 110 1368 116 1369
rect 132 1368 134 1429
rect 258 1411 264 1412
rect 218 1407 224 1408
rect 218 1403 219 1407
rect 223 1403 224 1407
rect 258 1407 259 1411
rect 263 1407 264 1411
rect 258 1406 264 1407
rect 218 1402 224 1403
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 130 1367 136 1368
rect 130 1363 131 1367
rect 135 1363 136 1367
rect 130 1362 136 1363
rect 158 1352 164 1353
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 158 1348 159 1352
rect 163 1348 164 1352
rect 158 1347 164 1348
rect 110 1346 116 1347
rect 112 1323 114 1346
rect 160 1323 162 1347
rect 111 1322 115 1323
rect 111 1317 115 1318
rect 159 1322 163 1323
rect 159 1317 163 1318
rect 112 1294 114 1317
rect 110 1293 116 1294
rect 160 1293 162 1317
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 158 1292 164 1293
rect 158 1288 159 1292
rect 163 1288 164 1292
rect 158 1287 164 1288
rect 130 1277 136 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 130 1273 131 1277
rect 135 1273 136 1277
rect 130 1272 136 1273
rect 110 1271 116 1272
rect 112 1187 114 1271
rect 132 1187 134 1272
rect 220 1268 222 1402
rect 260 1376 262 1406
rect 388 1376 390 1466
rect 484 1435 486 1508
rect 572 1472 574 1618
rect 620 1616 622 1677
rect 876 1616 878 1677
rect 962 1655 968 1656
rect 962 1651 963 1655
rect 967 1651 968 1655
rect 962 1650 968 1651
rect 964 1636 966 1650
rect 962 1635 968 1636
rect 962 1631 963 1635
rect 967 1631 968 1635
rect 962 1630 968 1631
rect 1140 1616 1142 1677
rect 1244 1660 1246 1746
rect 1364 1683 1366 1756
rect 1380 1720 1382 1866
rect 1484 1864 1486 1925
rect 1610 1907 1616 1908
rect 1610 1903 1611 1907
rect 1615 1903 1616 1907
rect 1610 1902 1616 1903
rect 1612 1872 1614 1902
rect 1610 1871 1616 1872
rect 1610 1867 1611 1871
rect 1615 1867 1616 1871
rect 1610 1866 1616 1867
rect 1644 1864 1646 1925
rect 1740 1872 1742 1962
rect 1788 1931 1790 2004
rect 1934 2003 1940 2004
rect 1802 1999 1808 2000
rect 1802 1995 1803 1999
rect 1807 1995 1808 1999
rect 1802 1994 1808 1995
rect 1804 1968 1806 1994
rect 1802 1967 1808 1968
rect 1802 1963 1803 1967
rect 1807 1963 1808 1967
rect 1802 1962 1808 1963
rect 1936 1931 1938 2003
rect 1976 1931 1978 2154
rect 2024 1931 2026 2155
rect 2184 1931 2186 2155
rect 2416 1931 2418 2155
rect 2696 1931 2698 2155
rect 3016 1931 3018 2155
rect 3360 1931 3362 2155
rect 3680 1931 3682 2155
rect 3798 2154 3804 2155
rect 3800 1931 3802 2154
rect 3840 2133 3842 2193
rect 3838 2132 3844 2133
rect 3860 2132 3862 2193
rect 3964 2176 3966 2254
rect 4156 2199 4158 2264
rect 4242 2251 4248 2252
rect 4242 2247 4243 2251
rect 4247 2247 4248 2251
rect 4242 2246 4248 2247
rect 4244 2228 4246 2246
rect 4242 2227 4248 2228
rect 4242 2223 4243 2227
rect 4247 2223 4248 2227
rect 4242 2222 4248 2223
rect 4468 2199 4470 2264
rect 4482 2259 4488 2260
rect 4482 2255 4483 2259
rect 4487 2255 4488 2259
rect 4482 2254 4488 2255
rect 4626 2259 4632 2260
rect 4626 2255 4627 2259
rect 4631 2255 4632 2259
rect 4626 2254 4632 2255
rect 4484 2228 4486 2254
rect 4482 2227 4488 2228
rect 4482 2223 4483 2227
rect 4487 2223 4488 2227
rect 4482 2222 4488 2223
rect 3995 2198 3999 2199
rect 3995 2193 3999 2194
rect 4131 2198 4135 2199
rect 4131 2193 4135 2194
rect 4155 2198 4159 2199
rect 4155 2193 4159 2194
rect 4267 2198 4271 2199
rect 4267 2193 4271 2194
rect 4403 2198 4407 2199
rect 4403 2193 4407 2194
rect 4467 2198 4471 2199
rect 4467 2193 4471 2194
rect 4539 2198 4543 2199
rect 4539 2193 4543 2194
rect 3962 2175 3968 2176
rect 3962 2171 3963 2175
rect 3967 2171 3968 2175
rect 3962 2170 3968 2171
rect 3986 2175 3992 2176
rect 3986 2171 3987 2175
rect 3991 2171 3992 2175
rect 3986 2170 3992 2171
rect 3988 2140 3990 2170
rect 3986 2139 3992 2140
rect 3986 2135 3987 2139
rect 3991 2135 3992 2139
rect 3986 2134 3992 2135
rect 3996 2132 3998 2193
rect 4132 2132 4134 2193
rect 4268 2132 4270 2193
rect 4404 2132 4406 2193
rect 4490 2139 4496 2140
rect 4490 2135 4491 2139
rect 4495 2135 4496 2139
rect 4490 2134 4496 2135
rect 3838 2128 3839 2132
rect 3843 2128 3844 2132
rect 3838 2127 3844 2128
rect 3858 2131 3864 2132
rect 3858 2127 3859 2131
rect 3863 2127 3864 2131
rect 3858 2126 3864 2127
rect 3994 2131 4000 2132
rect 3994 2127 3995 2131
rect 3999 2127 4000 2131
rect 3994 2126 4000 2127
rect 4130 2131 4136 2132
rect 4130 2127 4131 2131
rect 4135 2127 4136 2131
rect 4130 2126 4136 2127
rect 4266 2131 4272 2132
rect 4266 2127 4267 2131
rect 4271 2127 4272 2131
rect 4266 2126 4272 2127
rect 4402 2131 4408 2132
rect 4402 2127 4403 2131
rect 4407 2127 4408 2131
rect 4402 2126 4408 2127
rect 3886 2116 3892 2117
rect 3838 2115 3844 2116
rect 3838 2111 3839 2115
rect 3843 2111 3844 2115
rect 3886 2112 3887 2116
rect 3891 2112 3892 2116
rect 3886 2111 3892 2112
rect 4022 2116 4028 2117
rect 4022 2112 4023 2116
rect 4027 2112 4028 2116
rect 4022 2111 4028 2112
rect 4158 2116 4164 2117
rect 4158 2112 4159 2116
rect 4163 2112 4164 2116
rect 4158 2111 4164 2112
rect 4294 2116 4300 2117
rect 4294 2112 4295 2116
rect 4299 2112 4300 2116
rect 4294 2111 4300 2112
rect 4430 2116 4436 2117
rect 4430 2112 4431 2116
rect 4435 2112 4436 2116
rect 4430 2111 4436 2112
rect 3838 2110 3844 2111
rect 3840 2067 3842 2110
rect 3888 2067 3890 2111
rect 4024 2067 4026 2111
rect 4160 2067 4162 2111
rect 4296 2067 4298 2111
rect 4432 2067 4434 2111
rect 3839 2066 3843 2067
rect 3839 2061 3843 2062
rect 3887 2066 3891 2067
rect 3887 2061 3891 2062
rect 4023 2066 4027 2067
rect 4023 2061 4027 2062
rect 4159 2066 4163 2067
rect 4159 2061 4163 2062
rect 4295 2066 4299 2067
rect 4295 2061 4299 2062
rect 4431 2066 4435 2067
rect 4431 2061 4435 2062
rect 3840 2038 3842 2061
rect 3838 2037 3844 2038
rect 3888 2037 3890 2061
rect 4024 2037 4026 2061
rect 4160 2037 4162 2061
rect 4296 2037 4298 2061
rect 4432 2037 4434 2061
rect 3838 2033 3839 2037
rect 3843 2033 3844 2037
rect 3838 2032 3844 2033
rect 3886 2036 3892 2037
rect 3886 2032 3887 2036
rect 3891 2032 3892 2036
rect 3886 2031 3892 2032
rect 4022 2036 4028 2037
rect 4022 2032 4023 2036
rect 4027 2032 4028 2036
rect 4022 2031 4028 2032
rect 4158 2036 4164 2037
rect 4158 2032 4159 2036
rect 4163 2032 4164 2036
rect 4158 2031 4164 2032
rect 4294 2036 4300 2037
rect 4294 2032 4295 2036
rect 4299 2032 4300 2036
rect 4294 2031 4300 2032
rect 4430 2036 4436 2037
rect 4430 2032 4431 2036
rect 4435 2032 4436 2036
rect 4430 2031 4436 2032
rect 3858 2021 3864 2022
rect 3838 2020 3844 2021
rect 3838 2016 3839 2020
rect 3843 2016 3844 2020
rect 3858 2017 3859 2021
rect 3863 2017 3864 2021
rect 3858 2016 3864 2017
rect 3994 2021 4000 2022
rect 3994 2017 3995 2021
rect 3999 2017 4000 2021
rect 3994 2016 4000 2017
rect 4130 2021 4136 2022
rect 4130 2017 4131 2021
rect 4135 2017 4136 2021
rect 4130 2016 4136 2017
rect 4266 2021 4272 2022
rect 4266 2017 4267 2021
rect 4271 2017 4272 2021
rect 4266 2016 4272 2017
rect 4402 2021 4408 2022
rect 4402 2017 4403 2021
rect 4407 2017 4408 2021
rect 4402 2016 4408 2017
rect 3838 2015 3844 2016
rect 3840 1955 3842 2015
rect 3860 1955 3862 2016
rect 3962 2011 3968 2012
rect 3962 2007 3963 2011
rect 3967 2007 3968 2011
rect 3962 2006 3968 2007
rect 3839 1954 3843 1955
rect 3839 1949 3843 1950
rect 3859 1954 3863 1955
rect 3859 1949 3863 1950
rect 1787 1930 1791 1931
rect 1787 1925 1791 1926
rect 1935 1930 1939 1931
rect 1935 1925 1939 1926
rect 1975 1930 1979 1931
rect 1975 1925 1979 1926
rect 2023 1930 2027 1931
rect 2023 1925 2027 1926
rect 2183 1930 2187 1931
rect 2183 1925 2187 1926
rect 2415 1930 2419 1931
rect 2415 1925 2419 1926
rect 2695 1930 2699 1931
rect 2695 1925 2699 1926
rect 3015 1930 3019 1931
rect 3015 1925 3019 1926
rect 3135 1930 3139 1931
rect 3135 1925 3139 1926
rect 3271 1930 3275 1931
rect 3271 1925 3275 1926
rect 3359 1930 3363 1931
rect 3359 1925 3363 1926
rect 3407 1930 3411 1931
rect 3407 1925 3411 1926
rect 3543 1930 3547 1931
rect 3543 1925 3547 1926
rect 3679 1930 3683 1931
rect 3679 1925 3683 1926
rect 3799 1930 3803 1931
rect 3799 1925 3803 1926
rect 1738 1871 1744 1872
rect 1738 1867 1739 1871
rect 1743 1867 1744 1871
rect 1738 1866 1744 1867
rect 1788 1864 1790 1925
rect 1936 1865 1938 1925
rect 1976 1902 1978 1925
rect 2002 1907 2008 1908
rect 2002 1903 2003 1907
rect 2007 1903 2008 1907
rect 2002 1902 2008 1903
rect 1974 1901 1980 1902
rect 1974 1897 1975 1901
rect 1979 1897 1980 1901
rect 1974 1896 1980 1897
rect 1974 1884 1980 1885
rect 1974 1880 1975 1884
rect 1979 1880 1980 1884
rect 1974 1879 1980 1880
rect 1934 1864 1940 1865
rect 1482 1863 1488 1864
rect 1482 1859 1483 1863
rect 1487 1859 1488 1863
rect 1482 1858 1488 1859
rect 1642 1863 1648 1864
rect 1642 1859 1643 1863
rect 1647 1859 1648 1863
rect 1642 1858 1648 1859
rect 1786 1863 1792 1864
rect 1786 1859 1787 1863
rect 1791 1859 1792 1863
rect 1934 1860 1935 1864
rect 1939 1860 1940 1864
rect 1934 1859 1940 1860
rect 1786 1858 1792 1859
rect 1510 1848 1516 1849
rect 1510 1844 1511 1848
rect 1515 1844 1516 1848
rect 1510 1843 1516 1844
rect 1670 1848 1676 1849
rect 1670 1844 1671 1848
rect 1675 1844 1676 1848
rect 1670 1843 1676 1844
rect 1814 1848 1820 1849
rect 1814 1844 1815 1848
rect 1819 1844 1820 1848
rect 1814 1843 1820 1844
rect 1934 1847 1940 1848
rect 1934 1843 1935 1847
rect 1939 1843 1940 1847
rect 1512 1807 1514 1843
rect 1672 1807 1674 1843
rect 1816 1807 1818 1843
rect 1934 1842 1940 1843
rect 1936 1807 1938 1842
rect 1976 1807 1978 1879
rect 1391 1806 1395 1807
rect 1391 1801 1395 1802
rect 1511 1806 1515 1807
rect 1511 1801 1515 1802
rect 1671 1806 1675 1807
rect 1671 1801 1675 1802
rect 1815 1806 1819 1807
rect 1815 1801 1819 1802
rect 1935 1806 1939 1807
rect 1935 1801 1939 1802
rect 1975 1806 1979 1807
rect 1975 1801 1979 1802
rect 1995 1806 1999 1807
rect 1995 1801 1999 1802
rect 1392 1777 1394 1801
rect 1936 1778 1938 1801
rect 1934 1777 1940 1778
rect 1390 1776 1396 1777
rect 1390 1772 1391 1776
rect 1395 1772 1396 1776
rect 1934 1773 1935 1777
rect 1939 1773 1940 1777
rect 1934 1772 1940 1773
rect 1390 1771 1396 1772
rect 1934 1760 1940 1761
rect 1934 1756 1935 1760
rect 1939 1756 1940 1760
rect 1934 1755 1940 1756
rect 1378 1719 1384 1720
rect 1378 1715 1379 1719
rect 1383 1715 1384 1719
rect 1378 1714 1384 1715
rect 1936 1683 1938 1755
rect 1976 1741 1978 1801
rect 1974 1740 1980 1741
rect 1996 1740 1998 1801
rect 2004 1748 2006 1902
rect 3136 1901 3138 1925
rect 3272 1901 3274 1925
rect 3408 1901 3410 1925
rect 3544 1901 3546 1925
rect 3680 1901 3682 1925
rect 3800 1902 3802 1925
rect 3798 1901 3804 1902
rect 3134 1900 3140 1901
rect 3134 1896 3135 1900
rect 3139 1896 3140 1900
rect 3134 1895 3140 1896
rect 3270 1900 3276 1901
rect 3270 1896 3271 1900
rect 3275 1896 3276 1900
rect 3270 1895 3276 1896
rect 3406 1900 3412 1901
rect 3406 1896 3407 1900
rect 3411 1896 3412 1900
rect 3406 1895 3412 1896
rect 3542 1900 3548 1901
rect 3542 1896 3543 1900
rect 3547 1896 3548 1900
rect 3542 1895 3548 1896
rect 3678 1900 3684 1901
rect 3678 1896 3679 1900
rect 3683 1896 3684 1900
rect 3798 1897 3799 1901
rect 3803 1897 3804 1901
rect 3798 1896 3804 1897
rect 3678 1895 3684 1896
rect 3822 1895 3828 1896
rect 3822 1891 3823 1895
rect 3827 1891 3828 1895
rect 3822 1890 3828 1891
rect 3106 1885 3112 1886
rect 3106 1881 3107 1885
rect 3111 1881 3112 1885
rect 3106 1880 3112 1881
rect 3242 1885 3248 1886
rect 3242 1881 3243 1885
rect 3247 1881 3248 1885
rect 3242 1880 3248 1881
rect 3378 1885 3384 1886
rect 3378 1881 3379 1885
rect 3383 1881 3384 1885
rect 3378 1880 3384 1881
rect 3514 1885 3520 1886
rect 3514 1881 3515 1885
rect 3519 1881 3520 1885
rect 3514 1880 3520 1881
rect 3650 1885 3656 1886
rect 3650 1881 3651 1885
rect 3655 1881 3656 1885
rect 3650 1880 3656 1881
rect 3798 1884 3804 1885
rect 3798 1880 3799 1884
rect 3803 1880 3804 1884
rect 3108 1807 3110 1880
rect 3194 1867 3200 1868
rect 3194 1863 3195 1867
rect 3199 1863 3200 1867
rect 3194 1862 3200 1863
rect 3196 1844 3198 1862
rect 3194 1843 3200 1844
rect 3194 1839 3195 1843
rect 3199 1839 3200 1843
rect 3194 1838 3200 1839
rect 3244 1807 3246 1880
rect 3258 1875 3264 1876
rect 3258 1871 3259 1875
rect 3263 1871 3264 1875
rect 3258 1870 3264 1871
rect 3346 1875 3352 1876
rect 3346 1871 3347 1875
rect 3351 1871 3352 1875
rect 3346 1870 3352 1871
rect 3260 1844 3262 1870
rect 3258 1843 3264 1844
rect 3258 1839 3259 1843
rect 3263 1839 3264 1843
rect 3258 1838 3264 1839
rect 2131 1806 2135 1807
rect 2131 1801 2135 1802
rect 2267 1806 2271 1807
rect 2267 1801 2271 1802
rect 2419 1806 2423 1807
rect 2419 1801 2423 1802
rect 2579 1806 2583 1807
rect 2579 1801 2583 1802
rect 2739 1806 2743 1807
rect 2739 1801 2743 1802
rect 2899 1806 2903 1807
rect 2899 1801 2903 1802
rect 3051 1806 3055 1807
rect 3051 1801 3055 1802
rect 3107 1806 3111 1807
rect 3107 1801 3111 1802
rect 3203 1806 3207 1807
rect 3203 1801 3207 1802
rect 3243 1806 3247 1807
rect 3243 1801 3247 1802
rect 2002 1747 2008 1748
rect 2002 1743 2003 1747
rect 2007 1743 2008 1747
rect 2002 1742 2008 1743
rect 2132 1740 2134 1801
rect 2268 1740 2270 1801
rect 2420 1740 2422 1801
rect 2580 1740 2582 1801
rect 2722 1783 2728 1784
rect 2722 1779 2723 1783
rect 2727 1779 2728 1783
rect 2722 1778 2728 1779
rect 2730 1783 2736 1784
rect 2730 1779 2731 1783
rect 2735 1779 2736 1783
rect 2730 1778 2736 1779
rect 2724 1748 2726 1778
rect 2722 1747 2728 1748
rect 2722 1743 2723 1747
rect 2727 1743 2728 1747
rect 2722 1742 2728 1743
rect 1974 1736 1975 1740
rect 1979 1736 1980 1740
rect 1974 1735 1980 1736
rect 1994 1739 2000 1740
rect 1994 1735 1995 1739
rect 1999 1735 2000 1739
rect 1994 1734 2000 1735
rect 2130 1739 2136 1740
rect 2130 1735 2131 1739
rect 2135 1735 2136 1739
rect 2130 1734 2136 1735
rect 2266 1739 2272 1740
rect 2266 1735 2267 1739
rect 2271 1735 2272 1739
rect 2266 1734 2272 1735
rect 2418 1739 2424 1740
rect 2418 1735 2419 1739
rect 2423 1735 2424 1739
rect 2418 1734 2424 1735
rect 2578 1739 2584 1740
rect 2578 1735 2579 1739
rect 2583 1735 2584 1739
rect 2578 1734 2584 1735
rect 2022 1724 2028 1725
rect 1974 1723 1980 1724
rect 1974 1719 1975 1723
rect 1979 1719 1980 1723
rect 2022 1720 2023 1724
rect 2027 1720 2028 1724
rect 2022 1719 2028 1720
rect 2158 1724 2164 1725
rect 2158 1720 2159 1724
rect 2163 1720 2164 1724
rect 2158 1719 2164 1720
rect 2294 1724 2300 1725
rect 2294 1720 2295 1724
rect 2299 1720 2300 1724
rect 2294 1719 2300 1720
rect 2446 1724 2452 1725
rect 2446 1720 2447 1724
rect 2451 1720 2452 1724
rect 2446 1719 2452 1720
rect 2606 1724 2612 1725
rect 2606 1720 2607 1724
rect 2611 1720 2612 1724
rect 2606 1719 2612 1720
rect 1974 1718 1980 1719
rect 1976 1683 1978 1718
rect 2024 1683 2026 1719
rect 2160 1683 2162 1719
rect 2296 1683 2298 1719
rect 2448 1683 2450 1719
rect 2608 1683 2610 1719
rect 1363 1682 1367 1683
rect 1363 1677 1367 1678
rect 1935 1682 1939 1683
rect 1935 1677 1939 1678
rect 1975 1682 1979 1683
rect 1975 1677 1979 1678
rect 2023 1682 2027 1683
rect 2023 1677 2027 1678
rect 2159 1682 2163 1683
rect 2159 1677 2163 1678
rect 2167 1682 2171 1683
rect 2167 1677 2171 1678
rect 2295 1682 2299 1683
rect 2295 1677 2299 1678
rect 2319 1682 2323 1683
rect 2319 1677 2323 1678
rect 2447 1682 2451 1683
rect 2447 1677 2451 1678
rect 2479 1682 2483 1683
rect 2479 1677 2483 1678
rect 2607 1682 2611 1683
rect 2607 1677 2611 1678
rect 2639 1682 2643 1683
rect 2639 1677 2643 1678
rect 1242 1659 1248 1660
rect 1242 1655 1243 1659
rect 1247 1655 1248 1659
rect 1242 1654 1248 1655
rect 1936 1617 1938 1677
rect 1976 1654 1978 1677
rect 1974 1653 1980 1654
rect 2024 1653 2026 1677
rect 2168 1653 2170 1677
rect 2320 1653 2322 1677
rect 2480 1653 2482 1677
rect 2640 1653 2642 1677
rect 1974 1649 1975 1653
rect 1979 1649 1980 1653
rect 1974 1648 1980 1649
rect 2022 1652 2028 1653
rect 2022 1648 2023 1652
rect 2027 1648 2028 1652
rect 2022 1647 2028 1648
rect 2166 1652 2172 1653
rect 2166 1648 2167 1652
rect 2171 1648 2172 1652
rect 2166 1647 2172 1648
rect 2318 1652 2324 1653
rect 2318 1648 2319 1652
rect 2323 1648 2324 1652
rect 2318 1647 2324 1648
rect 2478 1652 2484 1653
rect 2478 1648 2479 1652
rect 2483 1648 2484 1652
rect 2478 1647 2484 1648
rect 2638 1652 2644 1653
rect 2638 1648 2639 1652
rect 2643 1648 2644 1652
rect 2638 1647 2644 1648
rect 1994 1637 2000 1638
rect 1974 1636 1980 1637
rect 1974 1632 1975 1636
rect 1979 1632 1980 1636
rect 1994 1633 1995 1637
rect 1999 1633 2000 1637
rect 1994 1632 2000 1633
rect 2138 1637 2144 1638
rect 2138 1633 2139 1637
rect 2143 1633 2144 1637
rect 2138 1632 2144 1633
rect 2290 1637 2296 1638
rect 2290 1633 2291 1637
rect 2295 1633 2296 1637
rect 2290 1632 2296 1633
rect 2450 1637 2456 1638
rect 2450 1633 2451 1637
rect 2455 1633 2456 1637
rect 2450 1632 2456 1633
rect 2610 1637 2616 1638
rect 2610 1633 2611 1637
rect 2615 1633 2616 1637
rect 2610 1632 2616 1633
rect 1974 1631 1980 1632
rect 1934 1616 1940 1617
rect 618 1615 624 1616
rect 618 1611 619 1615
rect 623 1611 624 1615
rect 618 1610 624 1611
rect 874 1615 880 1616
rect 874 1611 875 1615
rect 879 1611 880 1615
rect 874 1610 880 1611
rect 1138 1615 1144 1616
rect 1138 1611 1139 1615
rect 1143 1611 1144 1615
rect 1934 1612 1935 1616
rect 1939 1612 1940 1616
rect 1934 1611 1940 1612
rect 1138 1610 1144 1611
rect 646 1600 652 1601
rect 646 1596 647 1600
rect 651 1596 652 1600
rect 646 1595 652 1596
rect 902 1600 908 1601
rect 902 1596 903 1600
rect 907 1596 908 1600
rect 902 1595 908 1596
rect 1166 1600 1172 1601
rect 1166 1596 1167 1600
rect 1171 1596 1172 1600
rect 1166 1595 1172 1596
rect 1934 1599 1940 1600
rect 1934 1595 1935 1599
rect 1939 1595 1940 1599
rect 648 1559 650 1595
rect 904 1559 906 1595
rect 1168 1559 1170 1595
rect 1934 1594 1940 1595
rect 1936 1559 1938 1594
rect 1976 1559 1978 1631
rect 1996 1559 1998 1632
rect 2090 1595 2096 1596
rect 2090 1591 2091 1595
rect 2095 1591 2096 1595
rect 2090 1590 2096 1591
rect 647 1558 651 1559
rect 647 1553 651 1554
rect 695 1558 699 1559
rect 695 1553 699 1554
rect 887 1558 891 1559
rect 887 1553 891 1554
rect 903 1558 907 1559
rect 903 1553 907 1554
rect 1079 1558 1083 1559
rect 1079 1553 1083 1554
rect 1167 1558 1171 1559
rect 1167 1553 1171 1554
rect 1935 1558 1939 1559
rect 1935 1553 1939 1554
rect 1975 1558 1979 1559
rect 1975 1553 1979 1554
rect 1995 1558 1999 1559
rect 1995 1553 1999 1554
rect 696 1529 698 1553
rect 888 1529 890 1553
rect 1080 1529 1082 1553
rect 1936 1530 1938 1553
rect 1934 1529 1940 1530
rect 694 1528 700 1529
rect 694 1524 695 1528
rect 699 1524 700 1528
rect 694 1523 700 1524
rect 886 1528 892 1529
rect 886 1524 887 1528
rect 891 1524 892 1528
rect 886 1523 892 1524
rect 1078 1528 1084 1529
rect 1078 1524 1079 1528
rect 1083 1524 1084 1528
rect 1934 1525 1935 1529
rect 1939 1525 1940 1529
rect 1934 1524 1940 1525
rect 1078 1523 1084 1524
rect 666 1513 672 1514
rect 666 1509 667 1513
rect 671 1509 672 1513
rect 666 1508 672 1509
rect 858 1513 864 1514
rect 858 1509 859 1513
rect 863 1509 864 1513
rect 858 1508 864 1509
rect 1050 1513 1056 1514
rect 1050 1509 1051 1513
rect 1055 1509 1056 1513
rect 1050 1508 1056 1509
rect 1934 1512 1940 1513
rect 1934 1508 1935 1512
rect 1939 1508 1940 1512
rect 570 1471 576 1472
rect 570 1467 571 1471
rect 575 1467 576 1471
rect 570 1466 576 1467
rect 668 1435 670 1508
rect 682 1503 688 1504
rect 682 1499 683 1503
rect 687 1499 688 1503
rect 682 1498 688 1499
rect 684 1472 686 1498
rect 802 1495 808 1496
rect 802 1491 803 1495
rect 807 1491 808 1495
rect 802 1490 808 1491
rect 682 1471 688 1472
rect 682 1467 683 1471
rect 687 1467 688 1471
rect 682 1466 688 1467
rect 395 1434 399 1435
rect 395 1429 399 1430
rect 483 1434 487 1435
rect 483 1429 487 1430
rect 667 1434 671 1435
rect 667 1429 671 1430
rect 683 1434 687 1435
rect 683 1429 687 1430
rect 258 1375 264 1376
rect 258 1371 259 1375
rect 263 1371 264 1375
rect 258 1370 264 1371
rect 386 1375 392 1376
rect 386 1371 387 1375
rect 391 1371 392 1375
rect 386 1370 392 1371
rect 396 1368 398 1429
rect 684 1368 686 1429
rect 804 1412 806 1490
rect 860 1435 862 1508
rect 874 1503 880 1504
rect 874 1499 875 1503
rect 879 1499 880 1503
rect 874 1498 880 1499
rect 876 1472 878 1498
rect 874 1471 880 1472
rect 874 1467 875 1471
rect 879 1467 880 1471
rect 874 1466 880 1467
rect 1052 1435 1054 1508
rect 1934 1507 1940 1508
rect 1066 1503 1072 1504
rect 1066 1499 1067 1503
rect 1071 1499 1072 1503
rect 1066 1498 1072 1499
rect 1068 1472 1070 1498
rect 1066 1471 1072 1472
rect 1066 1467 1067 1471
rect 1071 1467 1072 1471
rect 1066 1466 1072 1467
rect 1936 1435 1938 1507
rect 1976 1493 1978 1553
rect 1974 1492 1980 1493
rect 1996 1492 1998 1553
rect 2092 1500 2094 1590
rect 2140 1559 2142 1632
rect 2154 1627 2160 1628
rect 2154 1623 2155 1627
rect 2159 1623 2160 1627
rect 2154 1622 2160 1623
rect 2156 1596 2158 1622
rect 2154 1595 2160 1596
rect 2154 1591 2155 1595
rect 2159 1591 2160 1595
rect 2154 1590 2160 1591
rect 2292 1559 2294 1632
rect 2306 1627 2312 1628
rect 2306 1623 2307 1627
rect 2311 1623 2312 1627
rect 2306 1622 2312 1623
rect 2308 1596 2310 1622
rect 2306 1595 2312 1596
rect 2306 1591 2307 1595
rect 2311 1591 2312 1595
rect 2306 1590 2312 1591
rect 2452 1559 2454 1632
rect 2466 1627 2472 1628
rect 2466 1623 2467 1627
rect 2471 1623 2472 1627
rect 2466 1622 2472 1623
rect 2468 1596 2470 1622
rect 2466 1595 2472 1596
rect 2466 1591 2467 1595
rect 2471 1591 2472 1595
rect 2466 1590 2472 1591
rect 2612 1559 2614 1632
rect 2732 1628 2734 1778
rect 2740 1740 2742 1801
rect 2900 1740 2902 1801
rect 3023 1788 3027 1789
rect 3022 1783 3028 1784
rect 3022 1779 3023 1783
rect 3027 1779 3028 1783
rect 3022 1778 3028 1779
rect 3052 1740 3054 1801
rect 3178 1783 3184 1784
rect 3178 1779 3179 1783
rect 3183 1779 3184 1783
rect 3178 1778 3184 1779
rect 3180 1748 3182 1778
rect 3178 1747 3184 1748
rect 3178 1743 3179 1747
rect 3183 1743 3184 1747
rect 3178 1742 3184 1743
rect 3204 1740 3206 1801
rect 3348 1784 3350 1870
rect 3380 1807 3382 1880
rect 3516 1807 3518 1880
rect 3652 1807 3654 1880
rect 3798 1879 3804 1880
rect 3800 1807 3802 1879
rect 3824 1844 3826 1890
rect 3840 1889 3842 1949
rect 3838 1888 3844 1889
rect 3860 1888 3862 1949
rect 3964 1932 3966 2006
rect 3996 1955 3998 2016
rect 4132 1955 4134 2016
rect 4268 1955 4270 2016
rect 4404 1955 4406 2016
rect 4492 1980 4494 2134
rect 4540 2132 4542 2193
rect 4628 2172 4630 2254
rect 4764 2199 4766 2264
rect 5002 2259 5008 2260
rect 5002 2255 5003 2259
rect 5007 2255 5008 2259
rect 5002 2254 5008 2255
rect 5004 2228 5006 2254
rect 5002 2227 5008 2228
rect 5002 2223 5003 2227
rect 5007 2223 5008 2227
rect 5002 2222 5008 2223
rect 5060 2199 5062 2264
rect 5278 2259 5284 2260
rect 5278 2255 5279 2259
rect 5283 2255 5284 2259
rect 5278 2254 5284 2255
rect 5280 2228 5282 2254
rect 5278 2227 5284 2228
rect 5278 2223 5279 2227
rect 5283 2223 5284 2227
rect 5278 2222 5284 2223
rect 5356 2199 5358 2264
rect 5372 2228 5374 2374
rect 5380 2372 5382 2433
rect 5400 2380 5402 2654
rect 5516 2616 5518 2677
rect 5620 2660 5622 2858
rect 5664 2857 5666 2917
rect 5662 2856 5668 2857
rect 5662 2852 5663 2856
rect 5667 2852 5668 2856
rect 5662 2851 5668 2852
rect 5662 2839 5668 2840
rect 5662 2835 5663 2839
rect 5667 2835 5668 2839
rect 5662 2834 5668 2835
rect 5664 2807 5666 2834
rect 5663 2806 5667 2807
rect 5663 2801 5667 2802
rect 5664 2778 5666 2801
rect 5662 2777 5668 2778
rect 5662 2773 5663 2777
rect 5667 2773 5668 2777
rect 5662 2772 5668 2773
rect 5662 2760 5668 2761
rect 5662 2756 5663 2760
rect 5667 2756 5668 2760
rect 5662 2755 5668 2756
rect 5664 2683 5666 2755
rect 5663 2682 5667 2683
rect 5663 2677 5667 2678
rect 5618 2659 5624 2660
rect 5618 2655 5619 2659
rect 5623 2655 5624 2659
rect 5618 2654 5624 2655
rect 5618 2623 5624 2624
rect 5618 2619 5619 2623
rect 5623 2619 5624 2623
rect 5618 2618 5624 2619
rect 5514 2615 5520 2616
rect 5514 2611 5515 2615
rect 5519 2611 5520 2615
rect 5514 2610 5520 2611
rect 5542 2600 5548 2601
rect 5542 2596 5543 2600
rect 5547 2596 5548 2600
rect 5542 2595 5548 2596
rect 5544 2567 5546 2595
rect 5543 2566 5547 2567
rect 5543 2561 5547 2562
rect 5515 2438 5519 2439
rect 5515 2433 5519 2434
rect 5466 2411 5472 2412
rect 5466 2407 5467 2411
rect 5471 2407 5472 2411
rect 5466 2406 5472 2407
rect 5468 2388 5470 2406
rect 5466 2387 5472 2388
rect 5466 2383 5467 2387
rect 5471 2383 5472 2387
rect 5466 2382 5472 2383
rect 5398 2379 5404 2380
rect 5398 2375 5399 2379
rect 5403 2375 5404 2379
rect 5398 2374 5404 2375
rect 5516 2372 5518 2433
rect 5620 2416 5622 2618
rect 5664 2617 5666 2677
rect 5662 2616 5668 2617
rect 5662 2612 5663 2616
rect 5667 2612 5668 2616
rect 5662 2611 5668 2612
rect 5662 2599 5668 2600
rect 5662 2595 5663 2599
rect 5667 2595 5668 2599
rect 5662 2594 5668 2595
rect 5664 2567 5666 2594
rect 5663 2566 5667 2567
rect 5663 2561 5667 2562
rect 5664 2538 5666 2561
rect 5662 2537 5668 2538
rect 5662 2533 5663 2537
rect 5667 2533 5668 2537
rect 5662 2532 5668 2533
rect 5662 2520 5668 2521
rect 5662 2516 5663 2520
rect 5667 2516 5668 2520
rect 5662 2515 5668 2516
rect 5664 2439 5666 2515
rect 5663 2438 5667 2439
rect 5663 2433 5667 2434
rect 5618 2415 5624 2416
rect 5618 2411 5619 2415
rect 5623 2411 5624 2415
rect 5618 2410 5624 2411
rect 5550 2387 5556 2388
rect 5550 2383 5551 2387
rect 5555 2383 5556 2387
rect 5550 2382 5556 2383
rect 5378 2371 5384 2372
rect 5378 2367 5379 2371
rect 5383 2367 5384 2371
rect 5378 2366 5384 2367
rect 5514 2371 5520 2372
rect 5514 2367 5515 2371
rect 5519 2367 5520 2371
rect 5514 2366 5520 2367
rect 5406 2356 5412 2357
rect 5406 2352 5407 2356
rect 5411 2352 5412 2356
rect 5406 2351 5412 2352
rect 5542 2356 5548 2357
rect 5542 2352 5543 2356
rect 5547 2352 5548 2356
rect 5542 2351 5548 2352
rect 5408 2315 5410 2351
rect 5544 2315 5546 2351
rect 5383 2314 5387 2315
rect 5383 2309 5387 2310
rect 5407 2314 5411 2315
rect 5407 2309 5411 2310
rect 5543 2314 5547 2315
rect 5543 2309 5547 2310
rect 5384 2285 5386 2309
rect 5382 2284 5388 2285
rect 5382 2280 5383 2284
rect 5387 2280 5388 2284
rect 5382 2279 5388 2280
rect 5370 2227 5376 2228
rect 5370 2223 5371 2227
rect 5375 2223 5376 2227
rect 5370 2222 5376 2223
rect 4699 2198 4703 2199
rect 4699 2193 4703 2194
rect 4763 2198 4767 2199
rect 4763 2193 4767 2194
rect 4891 2198 4895 2199
rect 4891 2193 4895 2194
rect 5059 2198 5063 2199
rect 5059 2193 5063 2194
rect 5099 2198 5103 2199
rect 5099 2193 5103 2194
rect 5315 2198 5319 2199
rect 5315 2193 5319 2194
rect 5355 2198 5359 2199
rect 5355 2193 5359 2194
rect 5515 2198 5519 2199
rect 5515 2193 5519 2194
rect 4666 2175 4672 2176
rect 4626 2171 4632 2172
rect 4626 2167 4627 2171
rect 4631 2167 4632 2171
rect 4666 2171 4667 2175
rect 4671 2171 4672 2175
rect 4666 2170 4672 2171
rect 4626 2166 4632 2167
rect 4668 2140 4670 2170
rect 4666 2139 4672 2140
rect 4666 2135 4667 2139
rect 4671 2135 4672 2139
rect 4666 2134 4672 2135
rect 4700 2132 4702 2193
rect 4826 2175 4832 2176
rect 4826 2171 4827 2175
rect 4831 2171 4832 2175
rect 4826 2170 4832 2171
rect 4828 2140 4830 2170
rect 4826 2139 4832 2140
rect 4826 2135 4827 2139
rect 4831 2135 4832 2139
rect 4826 2134 4832 2135
rect 4892 2132 4894 2193
rect 5018 2175 5024 2176
rect 5018 2171 5019 2175
rect 5023 2171 5024 2175
rect 5018 2170 5024 2171
rect 5020 2140 5022 2170
rect 5018 2139 5024 2140
rect 5018 2135 5019 2139
rect 5023 2135 5024 2139
rect 5018 2134 5024 2135
rect 5100 2132 5102 2193
rect 5316 2132 5318 2193
rect 5354 2139 5360 2140
rect 5354 2135 5355 2139
rect 5359 2135 5360 2139
rect 5354 2134 5360 2135
rect 4538 2131 4544 2132
rect 4538 2127 4539 2131
rect 4543 2127 4544 2131
rect 4538 2126 4544 2127
rect 4698 2131 4704 2132
rect 4698 2127 4699 2131
rect 4703 2127 4704 2131
rect 4698 2126 4704 2127
rect 4890 2131 4896 2132
rect 4890 2127 4891 2131
rect 4895 2127 4896 2131
rect 4890 2126 4896 2127
rect 5098 2131 5104 2132
rect 5098 2127 5099 2131
rect 5103 2127 5104 2131
rect 5098 2126 5104 2127
rect 5314 2131 5320 2132
rect 5314 2127 5315 2131
rect 5319 2127 5320 2131
rect 5314 2126 5320 2127
rect 4566 2116 4572 2117
rect 4566 2112 4567 2116
rect 4571 2112 4572 2116
rect 4566 2111 4572 2112
rect 4726 2116 4732 2117
rect 4726 2112 4727 2116
rect 4731 2112 4732 2116
rect 4726 2111 4732 2112
rect 4918 2116 4924 2117
rect 4918 2112 4919 2116
rect 4923 2112 4924 2116
rect 4918 2111 4924 2112
rect 5126 2116 5132 2117
rect 5126 2112 5127 2116
rect 5131 2112 5132 2116
rect 5126 2111 5132 2112
rect 5342 2116 5348 2117
rect 5342 2112 5343 2116
rect 5347 2112 5348 2116
rect 5342 2111 5348 2112
rect 4568 2067 4570 2111
rect 4728 2067 4730 2111
rect 4920 2067 4922 2111
rect 5128 2067 5130 2111
rect 5344 2067 5346 2111
rect 4567 2066 4571 2067
rect 4567 2061 4571 2062
rect 4719 2066 4723 2067
rect 4719 2061 4723 2062
rect 4727 2066 4731 2067
rect 4727 2061 4731 2062
rect 4895 2066 4899 2067
rect 4895 2061 4899 2062
rect 4919 2066 4923 2067
rect 4919 2061 4923 2062
rect 5087 2066 5091 2067
rect 5087 2061 5091 2062
rect 5127 2066 5131 2067
rect 5127 2061 5131 2062
rect 5279 2066 5283 2067
rect 5279 2061 5283 2062
rect 5343 2066 5347 2067
rect 5343 2061 5347 2062
rect 4568 2037 4570 2061
rect 4720 2037 4722 2061
rect 4896 2037 4898 2061
rect 5088 2037 5090 2061
rect 5280 2037 5282 2061
rect 4566 2036 4572 2037
rect 4566 2032 4567 2036
rect 4571 2032 4572 2036
rect 4566 2031 4572 2032
rect 4718 2036 4724 2037
rect 4718 2032 4719 2036
rect 4723 2032 4724 2036
rect 4718 2031 4724 2032
rect 4894 2036 4900 2037
rect 4894 2032 4895 2036
rect 4899 2032 4900 2036
rect 4894 2031 4900 2032
rect 5086 2036 5092 2037
rect 5086 2032 5087 2036
rect 5091 2032 5092 2036
rect 5086 2031 5092 2032
rect 5278 2036 5284 2037
rect 5278 2032 5279 2036
rect 5283 2032 5284 2036
rect 5278 2031 5284 2032
rect 4538 2021 4544 2022
rect 4538 2017 4539 2021
rect 4543 2017 4544 2021
rect 4538 2016 4544 2017
rect 4690 2021 4696 2022
rect 4690 2017 4691 2021
rect 4695 2017 4696 2021
rect 4690 2016 4696 2017
rect 4866 2021 4872 2022
rect 4866 2017 4867 2021
rect 4871 2017 4872 2021
rect 4866 2016 4872 2017
rect 5058 2021 5064 2022
rect 5058 2017 5059 2021
rect 5063 2017 5064 2021
rect 5058 2016 5064 2017
rect 5250 2021 5256 2022
rect 5250 2017 5251 2021
rect 5255 2017 5256 2021
rect 5250 2016 5256 2017
rect 4490 1979 4496 1980
rect 4490 1975 4491 1979
rect 4495 1975 4496 1979
rect 4490 1974 4496 1975
rect 4540 1955 4542 2016
rect 4682 2011 4688 2012
rect 4682 2007 4683 2011
rect 4687 2007 4688 2011
rect 4682 2006 4688 2007
rect 4684 1980 4686 2006
rect 4682 1979 4688 1980
rect 4682 1975 4683 1979
rect 4687 1975 4688 1979
rect 4682 1974 4688 1975
rect 4692 1955 4694 2016
rect 4834 2011 4840 2012
rect 4834 2007 4835 2011
rect 4839 2007 4840 2011
rect 4834 2006 4840 2007
rect 4836 1980 4838 2006
rect 4834 1979 4840 1980
rect 4834 1975 4835 1979
rect 4839 1975 4840 1979
rect 4834 1974 4840 1975
rect 4868 1955 4870 2016
rect 5060 1955 5062 2016
rect 5252 1955 5254 2016
rect 5356 1980 5358 2134
rect 5516 2132 5518 2193
rect 5514 2131 5520 2132
rect 5514 2127 5515 2131
rect 5519 2127 5520 2131
rect 5514 2126 5520 2127
rect 5542 2116 5548 2117
rect 5542 2112 5543 2116
rect 5547 2112 5548 2116
rect 5542 2111 5548 2112
rect 5544 2067 5546 2111
rect 5479 2066 5483 2067
rect 5479 2061 5483 2062
rect 5543 2066 5547 2067
rect 5543 2061 5547 2062
rect 5480 2037 5482 2061
rect 5478 2036 5484 2037
rect 5478 2032 5479 2036
rect 5483 2032 5484 2036
rect 5478 2031 5484 2032
rect 5450 2021 5456 2022
rect 5450 2017 5451 2021
rect 5455 2017 5456 2021
rect 5450 2016 5456 2017
rect 5354 1979 5360 1980
rect 5354 1975 5355 1979
rect 5359 1975 5360 1979
rect 5354 1974 5360 1975
rect 5452 1955 5454 2016
rect 5552 2012 5554 2382
rect 5618 2379 5624 2380
rect 5618 2375 5619 2379
rect 5623 2375 5624 2379
rect 5618 2374 5624 2375
rect 5620 2176 5622 2374
rect 5664 2373 5666 2433
rect 5662 2372 5668 2373
rect 5662 2368 5663 2372
rect 5667 2368 5668 2372
rect 5662 2367 5668 2368
rect 5662 2355 5668 2356
rect 5662 2351 5663 2355
rect 5667 2351 5668 2355
rect 5662 2350 5668 2351
rect 5664 2315 5666 2350
rect 5663 2314 5667 2315
rect 5663 2309 5667 2310
rect 5664 2286 5666 2309
rect 5662 2285 5668 2286
rect 5662 2281 5663 2285
rect 5667 2281 5668 2285
rect 5662 2280 5668 2281
rect 5662 2268 5668 2269
rect 5662 2264 5663 2268
rect 5667 2264 5668 2268
rect 5662 2263 5668 2264
rect 5664 2199 5666 2263
rect 5663 2198 5667 2199
rect 5663 2193 5667 2194
rect 5618 2175 5624 2176
rect 5618 2171 5619 2175
rect 5623 2171 5624 2175
rect 5618 2170 5624 2171
rect 5618 2139 5624 2140
rect 5618 2135 5619 2139
rect 5623 2135 5624 2139
rect 5618 2134 5624 2135
rect 5550 2011 5556 2012
rect 5550 2007 5551 2011
rect 5555 2007 5556 2011
rect 5550 2006 5556 2007
rect 5502 1979 5508 1980
rect 5502 1975 5503 1979
rect 5507 1975 5508 1979
rect 5502 1974 5508 1975
rect 3995 1954 3999 1955
rect 3995 1949 3999 1950
rect 4043 1954 4047 1955
rect 4043 1949 4047 1950
rect 4131 1954 4135 1955
rect 4131 1949 4135 1950
rect 4267 1954 4271 1955
rect 4267 1949 4271 1950
rect 4283 1954 4287 1955
rect 4283 1949 4287 1950
rect 4403 1954 4407 1955
rect 4403 1949 4407 1950
rect 4539 1954 4543 1955
rect 4539 1949 4543 1950
rect 4563 1954 4567 1955
rect 4563 1949 4567 1950
rect 4691 1954 4695 1955
rect 4691 1949 4695 1950
rect 4867 1954 4871 1955
rect 4867 1949 4871 1950
rect 4875 1954 4879 1955
rect 4875 1949 4879 1950
rect 5059 1954 5063 1955
rect 5059 1949 5063 1950
rect 5203 1954 5207 1955
rect 5203 1949 5207 1950
rect 5251 1954 5255 1955
rect 5251 1949 5255 1950
rect 5451 1954 5455 1955
rect 5451 1949 5455 1950
rect 3962 1931 3968 1932
rect 3962 1927 3963 1931
rect 3967 1927 3968 1931
rect 3962 1926 3968 1927
rect 4044 1888 4046 1949
rect 4170 1931 4176 1932
rect 4170 1927 4171 1931
rect 4175 1927 4176 1931
rect 4170 1926 4176 1927
rect 4172 1896 4174 1926
rect 4170 1895 4176 1896
rect 4170 1891 4171 1895
rect 4175 1891 4176 1895
rect 4170 1890 4176 1891
rect 4284 1888 4286 1949
rect 4410 1931 4416 1932
rect 4410 1927 4411 1931
rect 4415 1927 4416 1931
rect 4410 1926 4416 1927
rect 4412 1896 4414 1926
rect 4410 1895 4416 1896
rect 4410 1891 4411 1895
rect 4415 1891 4416 1895
rect 4410 1890 4416 1891
rect 4466 1895 4472 1896
rect 4466 1891 4467 1895
rect 4471 1891 4472 1895
rect 4466 1890 4472 1891
rect 3838 1884 3839 1888
rect 3843 1884 3844 1888
rect 3838 1883 3844 1884
rect 3858 1887 3864 1888
rect 3858 1883 3859 1887
rect 3863 1883 3864 1887
rect 3858 1882 3864 1883
rect 4042 1887 4048 1888
rect 4042 1883 4043 1887
rect 4047 1883 4048 1887
rect 4042 1882 4048 1883
rect 4282 1887 4288 1888
rect 4282 1883 4283 1887
rect 4287 1883 4288 1887
rect 4282 1882 4288 1883
rect 3886 1872 3892 1873
rect 3838 1871 3844 1872
rect 3838 1867 3839 1871
rect 3843 1867 3844 1871
rect 3886 1868 3887 1872
rect 3891 1868 3892 1872
rect 3886 1867 3892 1868
rect 4070 1872 4076 1873
rect 4070 1868 4071 1872
rect 4075 1868 4076 1872
rect 4070 1867 4076 1868
rect 4310 1872 4316 1873
rect 4310 1868 4311 1872
rect 4315 1868 4316 1872
rect 4310 1867 4316 1868
rect 3838 1866 3844 1867
rect 3822 1843 3828 1844
rect 3840 1843 3842 1866
rect 3888 1843 3890 1867
rect 4072 1843 4074 1867
rect 4312 1843 4314 1867
rect 3822 1839 3823 1843
rect 3827 1839 3828 1843
rect 3822 1838 3828 1839
rect 3839 1842 3843 1843
rect 3839 1837 3843 1838
rect 3887 1842 3891 1843
rect 3887 1837 3891 1838
rect 4071 1842 4075 1843
rect 4071 1837 4075 1838
rect 4311 1842 4315 1843
rect 4311 1837 4315 1838
rect 4407 1842 4411 1843
rect 4407 1837 4411 1838
rect 3840 1814 3842 1837
rect 3838 1813 3844 1814
rect 4408 1813 4410 1837
rect 3838 1809 3839 1813
rect 3843 1809 3844 1813
rect 3838 1808 3844 1809
rect 4406 1812 4412 1813
rect 4406 1808 4407 1812
rect 4411 1808 4412 1812
rect 4406 1807 4412 1808
rect 3355 1806 3359 1807
rect 3355 1801 3359 1802
rect 3379 1806 3383 1807
rect 3379 1801 3383 1802
rect 3515 1806 3519 1807
rect 3515 1801 3519 1802
rect 3651 1806 3655 1807
rect 3651 1801 3655 1802
rect 3799 1806 3803 1807
rect 3799 1801 3803 1802
rect 3346 1783 3352 1784
rect 3346 1779 3347 1783
rect 3351 1779 3352 1783
rect 3346 1778 3352 1779
rect 3322 1747 3328 1748
rect 3322 1743 3323 1747
rect 3327 1743 3328 1747
rect 3322 1742 3328 1743
rect 2738 1739 2744 1740
rect 2738 1735 2739 1739
rect 2743 1735 2744 1739
rect 2738 1734 2744 1735
rect 2898 1739 2904 1740
rect 2898 1735 2899 1739
rect 2903 1735 2904 1739
rect 2898 1734 2904 1735
rect 3050 1739 3056 1740
rect 3050 1735 3051 1739
rect 3055 1735 3056 1739
rect 3050 1734 3056 1735
rect 3202 1739 3208 1740
rect 3202 1735 3203 1739
rect 3207 1735 3208 1739
rect 3202 1734 3208 1735
rect 2766 1724 2772 1725
rect 2766 1720 2767 1724
rect 2771 1720 2772 1724
rect 2766 1719 2772 1720
rect 2926 1724 2932 1725
rect 2926 1720 2927 1724
rect 2931 1720 2932 1724
rect 2926 1719 2932 1720
rect 3078 1724 3084 1725
rect 3078 1720 3079 1724
rect 3083 1720 3084 1724
rect 3078 1719 3084 1720
rect 3230 1724 3236 1725
rect 3230 1720 3231 1724
rect 3235 1720 3236 1724
rect 3230 1719 3236 1720
rect 2768 1683 2770 1719
rect 2928 1683 2930 1719
rect 3080 1683 3082 1719
rect 3232 1683 3234 1719
rect 2767 1682 2771 1683
rect 2767 1677 2771 1678
rect 2791 1682 2795 1683
rect 2791 1677 2795 1678
rect 2927 1682 2931 1683
rect 2927 1677 2931 1678
rect 2943 1682 2947 1683
rect 2943 1677 2947 1678
rect 3079 1682 3083 1683
rect 3079 1677 3083 1678
rect 3103 1682 3107 1683
rect 3103 1677 3107 1678
rect 3231 1682 3235 1683
rect 3231 1677 3235 1678
rect 3263 1682 3267 1683
rect 3263 1677 3267 1678
rect 2792 1653 2794 1677
rect 2944 1653 2946 1677
rect 3104 1653 3106 1677
rect 3264 1653 3266 1677
rect 2790 1652 2796 1653
rect 2790 1648 2791 1652
rect 2795 1648 2796 1652
rect 2790 1647 2796 1648
rect 2942 1652 2948 1653
rect 2942 1648 2943 1652
rect 2947 1648 2948 1652
rect 2942 1647 2948 1648
rect 3102 1652 3108 1653
rect 3102 1648 3103 1652
rect 3107 1648 3108 1652
rect 3102 1647 3108 1648
rect 3262 1652 3268 1653
rect 3262 1648 3263 1652
rect 3267 1648 3268 1652
rect 3262 1647 3268 1648
rect 2762 1637 2768 1638
rect 2762 1633 2763 1637
rect 2767 1633 2768 1637
rect 2762 1632 2768 1633
rect 2914 1637 2920 1638
rect 2914 1633 2915 1637
rect 2919 1633 2920 1637
rect 2914 1632 2920 1633
rect 3074 1637 3080 1638
rect 3074 1633 3075 1637
rect 3079 1633 3080 1637
rect 3074 1632 3080 1633
rect 3234 1637 3240 1638
rect 3234 1633 3235 1637
rect 3239 1633 3240 1637
rect 3234 1632 3240 1633
rect 2626 1627 2632 1628
rect 2626 1623 2627 1627
rect 2631 1623 2632 1627
rect 2626 1622 2632 1623
rect 2730 1627 2736 1628
rect 2730 1623 2731 1627
rect 2735 1623 2736 1627
rect 2730 1622 2736 1623
rect 2628 1596 2630 1622
rect 2626 1595 2632 1596
rect 2626 1591 2627 1595
rect 2631 1591 2632 1595
rect 2626 1590 2632 1591
rect 2764 1559 2766 1632
rect 2850 1619 2856 1620
rect 2850 1615 2851 1619
rect 2855 1615 2856 1619
rect 2850 1614 2856 1615
rect 2852 1596 2854 1614
rect 2850 1595 2856 1596
rect 2850 1591 2851 1595
rect 2855 1591 2856 1595
rect 2850 1590 2856 1591
rect 2916 1559 2918 1632
rect 2930 1627 2936 1628
rect 2930 1623 2931 1627
rect 2935 1623 2936 1627
rect 2930 1622 2936 1623
rect 2932 1596 2934 1622
rect 2930 1595 2936 1596
rect 2930 1591 2931 1595
rect 2935 1591 2936 1595
rect 2930 1590 2936 1591
rect 3076 1559 3078 1632
rect 3090 1627 3096 1628
rect 3090 1623 3091 1627
rect 3095 1623 3096 1627
rect 3090 1622 3096 1623
rect 3092 1596 3094 1622
rect 3090 1595 3096 1596
rect 3090 1591 3091 1595
rect 3095 1591 3096 1595
rect 3090 1590 3096 1591
rect 3236 1559 3238 1632
rect 3324 1596 3326 1742
rect 3356 1740 3358 1801
rect 3482 1783 3488 1784
rect 3482 1779 3483 1783
rect 3487 1779 3488 1783
rect 3482 1778 3488 1779
rect 3484 1748 3486 1778
rect 3482 1747 3488 1748
rect 3482 1743 3483 1747
rect 3487 1743 3488 1747
rect 3482 1742 3488 1743
rect 3516 1740 3518 1801
rect 3652 1740 3654 1801
rect 3771 1788 3775 1789
rect 3771 1783 3775 1784
rect 3772 1748 3774 1783
rect 3770 1747 3776 1748
rect 3770 1743 3771 1747
rect 3775 1743 3776 1747
rect 3770 1742 3776 1743
rect 3800 1741 3802 1801
rect 4378 1797 4384 1798
rect 3838 1796 3844 1797
rect 3838 1792 3839 1796
rect 3843 1792 3844 1796
rect 4378 1793 4379 1797
rect 4383 1793 4384 1797
rect 4378 1792 4384 1793
rect 3838 1791 3844 1792
rect 3798 1740 3804 1741
rect 3354 1739 3360 1740
rect 3354 1735 3355 1739
rect 3359 1735 3360 1739
rect 3354 1734 3360 1735
rect 3514 1739 3520 1740
rect 3514 1735 3515 1739
rect 3519 1735 3520 1739
rect 3514 1734 3520 1735
rect 3650 1739 3656 1740
rect 3650 1735 3651 1739
rect 3655 1735 3656 1739
rect 3798 1736 3799 1740
rect 3803 1736 3804 1740
rect 3798 1735 3804 1736
rect 3650 1734 3656 1735
rect 3382 1724 3388 1725
rect 3382 1720 3383 1724
rect 3387 1720 3388 1724
rect 3382 1719 3388 1720
rect 3542 1724 3548 1725
rect 3542 1720 3543 1724
rect 3547 1720 3548 1724
rect 3542 1719 3548 1720
rect 3678 1724 3684 1725
rect 3678 1720 3679 1724
rect 3683 1720 3684 1724
rect 3678 1719 3684 1720
rect 3798 1723 3804 1724
rect 3798 1719 3799 1723
rect 3803 1719 3804 1723
rect 3384 1683 3386 1719
rect 3544 1683 3546 1719
rect 3680 1683 3682 1719
rect 3798 1718 3804 1719
rect 3800 1683 3802 1718
rect 3840 1715 3842 1791
rect 4380 1715 4382 1792
rect 4468 1756 4470 1890
rect 4564 1888 4566 1949
rect 4666 1943 4672 1944
rect 4666 1939 4667 1943
rect 4671 1939 4672 1943
rect 4666 1938 4672 1939
rect 4668 1896 4670 1938
rect 4690 1931 4696 1932
rect 4690 1927 4691 1931
rect 4695 1927 4696 1931
rect 4690 1926 4696 1927
rect 4692 1896 4694 1926
rect 4666 1895 4672 1896
rect 4666 1891 4667 1895
rect 4671 1891 4672 1895
rect 4666 1890 4672 1891
rect 4690 1895 4696 1896
rect 4690 1891 4691 1895
rect 4695 1891 4696 1895
rect 4690 1890 4696 1891
rect 4876 1888 4878 1949
rect 5002 1931 5008 1932
rect 5002 1927 5003 1931
rect 5007 1927 5008 1931
rect 5002 1926 5008 1927
rect 5004 1896 5006 1926
rect 5002 1895 5008 1896
rect 5002 1891 5003 1895
rect 5007 1891 5008 1895
rect 5002 1890 5008 1891
rect 5204 1888 5206 1949
rect 5326 1943 5332 1944
rect 5326 1939 5327 1943
rect 5331 1939 5332 1943
rect 5326 1938 5332 1939
rect 5328 1896 5330 1938
rect 5326 1895 5332 1896
rect 5326 1891 5327 1895
rect 5331 1891 5332 1895
rect 5326 1890 5332 1891
rect 4562 1887 4568 1888
rect 4562 1883 4563 1887
rect 4567 1883 4568 1887
rect 4562 1882 4568 1883
rect 4874 1887 4880 1888
rect 4874 1883 4875 1887
rect 4879 1883 4880 1887
rect 4874 1882 4880 1883
rect 5202 1887 5208 1888
rect 5202 1883 5203 1887
rect 5207 1883 5208 1887
rect 5202 1882 5208 1883
rect 4590 1872 4596 1873
rect 4590 1868 4591 1872
rect 4595 1868 4596 1872
rect 4590 1867 4596 1868
rect 4902 1872 4908 1873
rect 4902 1868 4903 1872
rect 4907 1868 4908 1872
rect 4902 1867 4908 1868
rect 5230 1872 5236 1873
rect 5230 1868 5231 1872
rect 5235 1868 5236 1872
rect 5230 1867 5236 1868
rect 4592 1843 4594 1867
rect 4904 1843 4906 1867
rect 5232 1843 5234 1867
rect 4543 1842 4547 1843
rect 4543 1837 4547 1838
rect 4591 1842 4595 1843
rect 4591 1837 4595 1838
rect 4679 1842 4683 1843
rect 4679 1837 4683 1838
rect 4815 1842 4819 1843
rect 4815 1837 4819 1838
rect 4903 1842 4907 1843
rect 4903 1837 4907 1838
rect 4951 1842 4955 1843
rect 4951 1837 4955 1838
rect 5231 1842 5235 1843
rect 5231 1837 5235 1838
rect 4544 1813 4546 1837
rect 4680 1813 4682 1837
rect 4816 1813 4818 1837
rect 4952 1813 4954 1837
rect 4542 1812 4548 1813
rect 4542 1808 4543 1812
rect 4547 1808 4548 1812
rect 4542 1807 4548 1808
rect 4678 1812 4684 1813
rect 4678 1808 4679 1812
rect 4683 1808 4684 1812
rect 4678 1807 4684 1808
rect 4814 1812 4820 1813
rect 4814 1808 4815 1812
rect 4819 1808 4820 1812
rect 4814 1807 4820 1808
rect 4950 1812 4956 1813
rect 4950 1808 4951 1812
rect 4955 1808 4956 1812
rect 4950 1807 4956 1808
rect 4514 1797 4520 1798
rect 4514 1793 4515 1797
rect 4519 1793 4520 1797
rect 4514 1792 4520 1793
rect 4650 1797 4656 1798
rect 4650 1793 4651 1797
rect 4655 1793 4656 1797
rect 4650 1792 4656 1793
rect 4786 1797 4792 1798
rect 4786 1793 4787 1797
rect 4791 1793 4792 1797
rect 4786 1792 4792 1793
rect 4922 1797 4928 1798
rect 4922 1793 4923 1797
rect 4927 1793 4928 1797
rect 4922 1792 4928 1793
rect 4466 1755 4472 1756
rect 4466 1751 4467 1755
rect 4471 1751 4472 1755
rect 4466 1750 4472 1751
rect 4516 1715 4518 1792
rect 4530 1787 4536 1788
rect 4530 1783 4531 1787
rect 4535 1783 4536 1787
rect 4530 1782 4536 1783
rect 4532 1756 4534 1782
rect 4530 1755 4536 1756
rect 4530 1751 4531 1755
rect 4535 1751 4536 1755
rect 4530 1750 4536 1751
rect 4652 1715 4654 1792
rect 4666 1787 4672 1788
rect 4666 1783 4667 1787
rect 4671 1783 4672 1787
rect 4666 1782 4672 1783
rect 4668 1756 4670 1782
rect 4666 1755 4672 1756
rect 4666 1751 4667 1755
rect 4671 1751 4672 1755
rect 4666 1750 4672 1751
rect 4788 1715 4790 1792
rect 4802 1787 4808 1788
rect 4802 1783 4803 1787
rect 4807 1783 4808 1787
rect 4802 1782 4808 1783
rect 4804 1756 4806 1782
rect 4802 1755 4808 1756
rect 4802 1751 4803 1755
rect 4807 1751 4808 1755
rect 4802 1750 4808 1751
rect 4924 1715 4926 1792
rect 4938 1787 4944 1788
rect 4938 1783 4939 1787
rect 4943 1783 4944 1787
rect 4938 1782 4944 1783
rect 4950 1787 4956 1788
rect 4950 1783 4951 1787
rect 4955 1783 4956 1787
rect 4950 1782 4956 1783
rect 4940 1756 4942 1782
rect 4938 1755 4944 1756
rect 4938 1751 4939 1755
rect 4943 1751 4944 1755
rect 4938 1750 4944 1751
rect 3839 1714 3843 1715
rect 3839 1709 3843 1710
rect 4379 1714 4383 1715
rect 4379 1709 4383 1710
rect 4515 1714 4519 1715
rect 4515 1709 4519 1710
rect 4563 1714 4567 1715
rect 4563 1709 4567 1710
rect 4651 1714 4655 1715
rect 4651 1709 4655 1710
rect 4699 1714 4703 1715
rect 4699 1709 4703 1710
rect 4787 1714 4791 1715
rect 4787 1709 4791 1710
rect 4835 1714 4839 1715
rect 4835 1709 4839 1710
rect 4923 1714 4927 1715
rect 4923 1709 4927 1710
rect 3383 1682 3387 1683
rect 3383 1677 3387 1678
rect 3423 1682 3427 1683
rect 3423 1677 3427 1678
rect 3543 1682 3547 1683
rect 3543 1677 3547 1678
rect 3679 1682 3683 1683
rect 3679 1677 3683 1678
rect 3799 1682 3803 1683
rect 3799 1677 3803 1678
rect 3424 1653 3426 1677
rect 3800 1654 3802 1677
rect 3798 1653 3804 1654
rect 3422 1652 3428 1653
rect 3422 1648 3423 1652
rect 3427 1648 3428 1652
rect 3798 1649 3799 1653
rect 3803 1649 3804 1653
rect 3840 1649 3842 1709
rect 3798 1648 3804 1649
rect 3838 1648 3844 1649
rect 4564 1648 4566 1709
rect 4650 1655 4656 1656
rect 4650 1651 4651 1655
rect 4655 1651 4656 1655
rect 4650 1650 4656 1651
rect 3422 1647 3428 1648
rect 3838 1644 3839 1648
rect 3843 1644 3844 1648
rect 3838 1643 3844 1644
rect 4562 1647 4568 1648
rect 4562 1643 4563 1647
rect 4567 1643 4568 1647
rect 4562 1642 4568 1643
rect 3394 1637 3400 1638
rect 3394 1633 3395 1637
rect 3399 1633 3400 1637
rect 3394 1632 3400 1633
rect 3798 1636 3804 1637
rect 3798 1632 3799 1636
rect 3803 1632 3804 1636
rect 4590 1632 4596 1633
rect 3322 1595 3328 1596
rect 3322 1591 3323 1595
rect 3327 1591 3328 1595
rect 3322 1590 3328 1591
rect 3396 1559 3398 1632
rect 3798 1631 3804 1632
rect 3838 1631 3844 1632
rect 3410 1627 3416 1628
rect 3410 1623 3411 1627
rect 3415 1623 3416 1627
rect 3410 1622 3416 1623
rect 3412 1596 3414 1622
rect 3410 1595 3416 1596
rect 3410 1591 3411 1595
rect 3415 1591 3416 1595
rect 3410 1590 3416 1591
rect 3800 1559 3802 1631
rect 3838 1627 3839 1631
rect 3843 1627 3844 1631
rect 4590 1628 4591 1632
rect 4595 1628 4596 1632
rect 4590 1627 4596 1628
rect 3838 1626 3844 1627
rect 3840 1587 3842 1626
rect 4592 1587 4594 1627
rect 3839 1586 3843 1587
rect 3839 1581 3843 1582
rect 4591 1586 4595 1587
rect 4591 1581 4595 1582
rect 2131 1558 2135 1559
rect 2131 1553 2135 1554
rect 2139 1558 2143 1559
rect 2139 1553 2143 1554
rect 2267 1558 2271 1559
rect 2267 1553 2271 1554
rect 2291 1558 2295 1559
rect 2291 1553 2295 1554
rect 2403 1558 2407 1559
rect 2403 1553 2407 1554
rect 2451 1558 2455 1559
rect 2451 1553 2455 1554
rect 2539 1558 2543 1559
rect 2539 1553 2543 1554
rect 2611 1558 2615 1559
rect 2611 1553 2615 1554
rect 2675 1558 2679 1559
rect 2675 1553 2679 1554
rect 2763 1558 2767 1559
rect 2763 1553 2767 1554
rect 2811 1558 2815 1559
rect 2811 1553 2815 1554
rect 2915 1558 2919 1559
rect 2915 1553 2919 1554
rect 2947 1558 2951 1559
rect 2947 1553 2951 1554
rect 3075 1558 3079 1559
rect 3075 1553 3079 1554
rect 3083 1558 3087 1559
rect 3083 1553 3087 1554
rect 3219 1558 3223 1559
rect 3219 1553 3223 1554
rect 3235 1558 3239 1559
rect 3235 1553 3239 1554
rect 3355 1558 3359 1559
rect 3355 1553 3359 1554
rect 3395 1558 3399 1559
rect 3395 1553 3399 1554
rect 3491 1558 3495 1559
rect 3491 1553 3495 1554
rect 3799 1558 3803 1559
rect 3840 1558 3842 1581
rect 3799 1553 3803 1554
rect 3838 1557 3844 1558
rect 4592 1557 4594 1581
rect 3838 1553 3839 1557
rect 3843 1553 3844 1557
rect 2090 1499 2096 1500
rect 2090 1495 2091 1499
rect 2095 1495 2096 1499
rect 2090 1494 2096 1495
rect 2132 1492 2134 1553
rect 2258 1535 2264 1536
rect 2258 1531 2259 1535
rect 2263 1531 2264 1535
rect 2258 1530 2264 1531
rect 1974 1488 1975 1492
rect 1979 1488 1980 1492
rect 1974 1487 1980 1488
rect 1994 1491 2000 1492
rect 1994 1487 1995 1491
rect 1999 1487 2000 1491
rect 1994 1486 2000 1487
rect 2130 1491 2136 1492
rect 2130 1487 2131 1491
rect 2135 1487 2136 1491
rect 2130 1486 2136 1487
rect 2022 1476 2028 1477
rect 1974 1475 1980 1476
rect 1974 1471 1975 1475
rect 1979 1471 1980 1475
rect 2022 1472 2023 1476
rect 2027 1472 2028 1476
rect 2022 1471 2028 1472
rect 2158 1476 2164 1477
rect 2158 1472 2159 1476
rect 2163 1472 2164 1476
rect 2158 1471 2164 1472
rect 1974 1470 1980 1471
rect 1976 1435 1978 1470
rect 2024 1435 2026 1471
rect 2160 1435 2162 1471
rect 859 1434 863 1435
rect 859 1429 863 1430
rect 971 1434 975 1435
rect 971 1429 975 1430
rect 1051 1434 1055 1435
rect 1051 1429 1055 1430
rect 1259 1434 1263 1435
rect 1259 1429 1263 1430
rect 1935 1434 1939 1435
rect 1935 1429 1939 1430
rect 1975 1434 1979 1435
rect 1975 1429 1979 1430
rect 2023 1434 2027 1435
rect 2023 1429 2027 1430
rect 2159 1434 2163 1435
rect 2159 1429 2163 1430
rect 2167 1434 2171 1435
rect 2167 1429 2171 1430
rect 802 1411 808 1412
rect 802 1407 803 1411
rect 807 1407 808 1411
rect 802 1406 808 1407
rect 810 1411 816 1412
rect 810 1407 811 1411
rect 815 1407 816 1411
rect 810 1406 816 1407
rect 812 1376 814 1406
rect 810 1375 816 1376
rect 810 1371 811 1375
rect 815 1371 816 1375
rect 810 1370 816 1371
rect 972 1368 974 1429
rect 1098 1411 1104 1412
rect 1098 1407 1099 1411
rect 1103 1407 1104 1411
rect 1098 1406 1104 1407
rect 1100 1376 1102 1406
rect 1098 1375 1104 1376
rect 1098 1371 1099 1375
rect 1103 1371 1104 1375
rect 1098 1370 1104 1371
rect 1260 1368 1262 1429
rect 1410 1375 1416 1376
rect 1410 1371 1411 1375
rect 1415 1371 1416 1375
rect 1410 1370 1416 1371
rect 394 1367 400 1368
rect 394 1363 395 1367
rect 399 1363 400 1367
rect 394 1362 400 1363
rect 682 1367 688 1368
rect 682 1363 683 1367
rect 687 1363 688 1367
rect 682 1362 688 1363
rect 970 1367 976 1368
rect 970 1363 971 1367
rect 975 1363 976 1367
rect 970 1362 976 1363
rect 1258 1367 1264 1368
rect 1258 1363 1259 1367
rect 1263 1363 1264 1367
rect 1258 1362 1264 1363
rect 422 1352 428 1353
rect 422 1348 423 1352
rect 427 1348 428 1352
rect 422 1347 428 1348
rect 710 1352 716 1353
rect 710 1348 711 1352
rect 715 1348 716 1352
rect 710 1347 716 1348
rect 998 1352 1004 1353
rect 998 1348 999 1352
rect 1003 1348 1004 1352
rect 998 1347 1004 1348
rect 1286 1352 1292 1353
rect 1286 1348 1287 1352
rect 1291 1348 1292 1352
rect 1286 1347 1292 1348
rect 424 1323 426 1347
rect 712 1323 714 1347
rect 1000 1323 1002 1347
rect 1288 1323 1290 1347
rect 423 1322 427 1323
rect 423 1317 427 1318
rect 455 1322 459 1323
rect 455 1317 459 1318
rect 711 1322 715 1323
rect 711 1317 715 1318
rect 775 1322 779 1323
rect 775 1317 779 1318
rect 999 1322 1003 1323
rect 999 1317 1003 1318
rect 1095 1322 1099 1323
rect 1095 1317 1099 1318
rect 1287 1322 1291 1323
rect 1287 1317 1291 1318
rect 456 1293 458 1317
rect 776 1293 778 1317
rect 1096 1293 1098 1317
rect 454 1292 460 1293
rect 454 1288 455 1292
rect 459 1288 460 1292
rect 454 1287 460 1288
rect 774 1292 780 1293
rect 774 1288 775 1292
rect 779 1288 780 1292
rect 774 1287 780 1288
rect 1094 1292 1100 1293
rect 1094 1288 1095 1292
rect 1099 1288 1100 1292
rect 1094 1287 1100 1288
rect 426 1277 432 1278
rect 426 1273 427 1277
rect 431 1273 432 1277
rect 426 1272 432 1273
rect 746 1277 752 1278
rect 746 1273 747 1277
rect 751 1273 752 1277
rect 746 1272 752 1273
rect 1066 1277 1072 1278
rect 1066 1273 1067 1277
rect 1071 1273 1072 1277
rect 1066 1272 1072 1273
rect 1394 1277 1400 1278
rect 1394 1273 1395 1277
rect 1399 1273 1400 1277
rect 1394 1272 1400 1273
rect 218 1267 224 1268
rect 218 1263 219 1267
rect 223 1263 224 1267
rect 218 1262 224 1263
rect 298 1267 304 1268
rect 298 1263 299 1267
rect 303 1263 304 1267
rect 298 1262 304 1263
rect 300 1236 302 1262
rect 298 1235 304 1236
rect 298 1231 299 1235
rect 303 1231 304 1235
rect 298 1230 304 1231
rect 428 1187 430 1272
rect 514 1235 520 1236
rect 514 1231 515 1235
rect 519 1231 520 1235
rect 514 1230 520 1231
rect 111 1186 115 1187
rect 111 1181 115 1182
rect 131 1186 135 1187
rect 131 1181 135 1182
rect 331 1186 335 1187
rect 331 1181 335 1182
rect 427 1186 431 1187
rect 427 1181 431 1182
rect 112 1121 114 1181
rect 110 1120 116 1121
rect 132 1120 134 1181
rect 258 1163 264 1164
rect 258 1159 259 1163
rect 263 1159 264 1163
rect 258 1158 264 1159
rect 260 1128 262 1158
rect 270 1155 276 1156
rect 270 1151 271 1155
rect 275 1151 276 1155
rect 270 1150 276 1151
rect 258 1127 264 1128
rect 258 1123 259 1127
rect 263 1123 264 1127
rect 258 1122 264 1123
rect 110 1116 111 1120
rect 115 1116 116 1120
rect 110 1115 116 1116
rect 130 1119 136 1120
rect 130 1115 131 1119
rect 135 1115 136 1119
rect 130 1114 136 1115
rect 158 1104 164 1105
rect 110 1103 116 1104
rect 110 1099 111 1103
rect 115 1099 116 1103
rect 158 1100 159 1104
rect 163 1100 164 1104
rect 158 1099 164 1100
rect 110 1098 116 1099
rect 112 1075 114 1098
rect 160 1075 162 1099
rect 111 1074 115 1075
rect 111 1069 115 1070
rect 159 1074 163 1075
rect 159 1069 163 1070
rect 263 1074 267 1075
rect 263 1069 267 1070
rect 112 1046 114 1069
rect 110 1045 116 1046
rect 264 1045 266 1069
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 262 1044 268 1045
rect 262 1040 263 1044
rect 267 1040 268 1044
rect 262 1039 268 1040
rect 234 1029 240 1030
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 234 1025 235 1029
rect 239 1025 240 1029
rect 234 1024 240 1025
rect 110 1023 116 1024
rect 112 959 114 1023
rect 236 959 238 1024
rect 272 1020 274 1150
rect 332 1120 334 1181
rect 458 1163 464 1164
rect 458 1159 459 1163
rect 463 1159 464 1163
rect 458 1158 464 1159
rect 460 1128 462 1158
rect 516 1128 518 1230
rect 748 1187 750 1272
rect 834 1259 840 1260
rect 834 1255 835 1259
rect 839 1255 840 1259
rect 834 1254 840 1255
rect 836 1236 838 1254
rect 834 1235 840 1236
rect 834 1231 835 1235
rect 839 1231 840 1235
rect 834 1230 840 1231
rect 1068 1187 1070 1272
rect 1082 1267 1088 1268
rect 1082 1263 1083 1267
rect 1087 1263 1088 1267
rect 1082 1262 1088 1263
rect 1084 1236 1086 1262
rect 1082 1235 1088 1236
rect 1082 1231 1083 1235
rect 1087 1231 1088 1235
rect 1082 1230 1088 1231
rect 1396 1187 1398 1272
rect 1412 1236 1414 1370
rect 1936 1369 1938 1429
rect 1976 1406 1978 1429
rect 1974 1405 1980 1406
rect 2168 1405 2170 1429
rect 1974 1401 1975 1405
rect 1979 1401 1980 1405
rect 1974 1400 1980 1401
rect 2166 1404 2172 1405
rect 2166 1400 2167 1404
rect 2171 1400 2172 1404
rect 2166 1399 2172 1400
rect 2138 1389 2144 1390
rect 1974 1388 1980 1389
rect 1974 1384 1975 1388
rect 1979 1384 1980 1388
rect 2138 1385 2139 1389
rect 2143 1385 2144 1389
rect 2138 1384 2144 1385
rect 1974 1383 1980 1384
rect 1934 1368 1940 1369
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 1934 1363 1940 1364
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 1934 1346 1940 1347
rect 1936 1323 1938 1346
rect 1976 1323 1978 1383
rect 2140 1323 2142 1384
rect 2260 1380 2262 1530
rect 2268 1492 2270 1553
rect 2404 1492 2406 1553
rect 2540 1492 2542 1553
rect 2626 1531 2632 1532
rect 2626 1527 2627 1531
rect 2631 1527 2632 1531
rect 2626 1526 2632 1527
rect 2628 1500 2630 1526
rect 2626 1499 2632 1500
rect 2626 1495 2627 1499
rect 2631 1495 2632 1499
rect 2626 1494 2632 1495
rect 2634 1499 2640 1500
rect 2634 1495 2635 1499
rect 2639 1495 2640 1499
rect 2634 1494 2640 1495
rect 2266 1491 2272 1492
rect 2266 1487 2267 1491
rect 2271 1487 2272 1491
rect 2266 1486 2272 1487
rect 2402 1491 2408 1492
rect 2402 1487 2403 1491
rect 2407 1487 2408 1491
rect 2402 1486 2408 1487
rect 2538 1491 2544 1492
rect 2538 1487 2539 1491
rect 2543 1487 2544 1491
rect 2538 1486 2544 1487
rect 2294 1476 2300 1477
rect 2294 1472 2295 1476
rect 2299 1472 2300 1476
rect 2294 1471 2300 1472
rect 2430 1476 2436 1477
rect 2430 1472 2431 1476
rect 2435 1472 2436 1476
rect 2430 1471 2436 1472
rect 2566 1476 2572 1477
rect 2566 1472 2567 1476
rect 2571 1472 2572 1476
rect 2566 1471 2572 1472
rect 2296 1435 2298 1471
rect 2432 1435 2434 1471
rect 2568 1435 2570 1471
rect 2295 1434 2299 1435
rect 2295 1429 2299 1430
rect 2303 1434 2307 1435
rect 2303 1429 2307 1430
rect 2431 1434 2435 1435
rect 2431 1429 2435 1430
rect 2439 1434 2443 1435
rect 2439 1429 2443 1430
rect 2567 1434 2571 1435
rect 2567 1429 2571 1430
rect 2575 1434 2579 1435
rect 2575 1429 2579 1430
rect 2304 1405 2306 1429
rect 2440 1405 2442 1429
rect 2576 1405 2578 1429
rect 2302 1404 2308 1405
rect 2302 1400 2303 1404
rect 2307 1400 2308 1404
rect 2302 1399 2308 1400
rect 2438 1404 2444 1405
rect 2438 1400 2439 1404
rect 2443 1400 2444 1404
rect 2438 1399 2444 1400
rect 2574 1404 2580 1405
rect 2574 1400 2575 1404
rect 2579 1400 2580 1404
rect 2574 1399 2580 1400
rect 2274 1389 2280 1390
rect 2274 1385 2275 1389
rect 2279 1385 2280 1389
rect 2274 1384 2280 1385
rect 2410 1389 2416 1390
rect 2410 1385 2411 1389
rect 2415 1385 2416 1389
rect 2410 1384 2416 1385
rect 2546 1389 2552 1390
rect 2546 1385 2547 1389
rect 2551 1385 2552 1389
rect 2546 1384 2552 1385
rect 2258 1379 2264 1380
rect 2258 1375 2259 1379
rect 2263 1375 2264 1379
rect 2258 1374 2264 1375
rect 2276 1323 2278 1384
rect 2412 1323 2414 1384
rect 2418 1379 2424 1380
rect 2418 1375 2419 1379
rect 2423 1375 2424 1379
rect 2418 1374 2424 1375
rect 2420 1348 2422 1374
rect 2418 1347 2424 1348
rect 2418 1343 2419 1347
rect 2423 1343 2424 1347
rect 2418 1342 2424 1343
rect 2498 1347 2504 1348
rect 2498 1343 2499 1347
rect 2503 1343 2504 1347
rect 2498 1342 2504 1343
rect 1423 1322 1427 1323
rect 1423 1317 1427 1318
rect 1935 1322 1939 1323
rect 1935 1317 1939 1318
rect 1975 1322 1979 1323
rect 1975 1317 1979 1318
rect 2131 1322 2135 1323
rect 2131 1317 2135 1318
rect 2139 1322 2143 1323
rect 2139 1317 2143 1318
rect 2267 1322 2271 1323
rect 2267 1317 2271 1318
rect 2275 1322 2279 1323
rect 2275 1317 2279 1318
rect 2403 1322 2407 1323
rect 2403 1317 2407 1318
rect 2411 1322 2415 1323
rect 2411 1317 2415 1318
rect 1424 1293 1426 1317
rect 1936 1294 1938 1317
rect 1934 1293 1940 1294
rect 1422 1292 1428 1293
rect 1422 1288 1423 1292
rect 1427 1288 1428 1292
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 1934 1288 1940 1289
rect 1422 1287 1428 1288
rect 1934 1276 1940 1277
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 1934 1271 1940 1272
rect 1410 1235 1416 1236
rect 1410 1231 1411 1235
rect 1415 1231 1416 1235
rect 1410 1230 1416 1231
rect 1936 1187 1938 1271
rect 1976 1257 1978 1317
rect 1974 1256 1980 1257
rect 2132 1256 2134 1317
rect 2246 1299 2252 1300
rect 2246 1295 2247 1299
rect 2251 1295 2252 1299
rect 2246 1294 2252 1295
rect 2258 1299 2264 1300
rect 2258 1295 2259 1299
rect 2263 1295 2264 1299
rect 2258 1294 2264 1295
rect 1974 1252 1975 1256
rect 1979 1252 1980 1256
rect 1974 1251 1980 1252
rect 2130 1255 2136 1256
rect 2130 1251 2131 1255
rect 2135 1251 2136 1255
rect 2130 1250 2136 1251
rect 2158 1240 2164 1241
rect 1974 1239 1980 1240
rect 1974 1235 1975 1239
rect 1979 1235 1980 1239
rect 2158 1236 2159 1240
rect 2163 1236 2164 1240
rect 2158 1235 2164 1236
rect 1974 1234 1980 1235
rect 1976 1211 1978 1234
rect 2160 1211 2162 1235
rect 2248 1216 2250 1294
rect 2260 1264 2262 1294
rect 2258 1263 2264 1264
rect 2258 1259 2259 1263
rect 2263 1259 2264 1263
rect 2258 1258 2264 1259
rect 2268 1256 2270 1317
rect 2404 1256 2406 1317
rect 2500 1301 2502 1342
rect 2548 1323 2550 1384
rect 2636 1348 2638 1494
rect 2676 1492 2678 1553
rect 2798 1519 2804 1520
rect 2798 1515 2799 1519
rect 2803 1515 2804 1519
rect 2798 1514 2804 1515
rect 2800 1500 2802 1514
rect 2798 1499 2804 1500
rect 2798 1495 2799 1499
rect 2803 1495 2804 1499
rect 2798 1494 2804 1495
rect 2812 1492 2814 1553
rect 2948 1492 2950 1553
rect 3084 1492 3086 1553
rect 3220 1492 3222 1553
rect 3356 1492 3358 1553
rect 3492 1492 3494 1553
rect 3614 1519 3620 1520
rect 3614 1515 3615 1519
rect 3619 1515 3620 1519
rect 3614 1514 3620 1515
rect 3616 1500 3618 1514
rect 3614 1499 3620 1500
rect 3614 1495 3615 1499
rect 3619 1495 3620 1499
rect 3614 1494 3620 1495
rect 3800 1493 3802 1553
rect 3838 1552 3844 1553
rect 4590 1556 4596 1557
rect 4590 1552 4591 1556
rect 4595 1552 4596 1556
rect 4590 1551 4596 1552
rect 4562 1541 4568 1542
rect 3838 1540 3844 1541
rect 3838 1536 3839 1540
rect 3843 1536 3844 1540
rect 4562 1537 4563 1541
rect 4567 1537 4568 1541
rect 4562 1536 4568 1537
rect 3838 1535 3844 1536
rect 3798 1492 3804 1493
rect 2674 1491 2680 1492
rect 2674 1487 2675 1491
rect 2679 1487 2680 1491
rect 2674 1486 2680 1487
rect 2810 1491 2816 1492
rect 2810 1487 2811 1491
rect 2815 1487 2816 1491
rect 2810 1486 2816 1487
rect 2946 1491 2952 1492
rect 2946 1487 2947 1491
rect 2951 1487 2952 1491
rect 2946 1486 2952 1487
rect 3082 1491 3088 1492
rect 3082 1487 3083 1491
rect 3087 1487 3088 1491
rect 3082 1486 3088 1487
rect 3218 1491 3224 1492
rect 3218 1487 3219 1491
rect 3223 1487 3224 1491
rect 3218 1486 3224 1487
rect 3354 1491 3360 1492
rect 3354 1487 3355 1491
rect 3359 1487 3360 1491
rect 3354 1486 3360 1487
rect 3490 1491 3496 1492
rect 3490 1487 3491 1491
rect 3495 1487 3496 1491
rect 3798 1488 3799 1492
rect 3803 1488 3804 1492
rect 3798 1487 3804 1488
rect 3490 1486 3496 1487
rect 2702 1476 2708 1477
rect 2702 1472 2703 1476
rect 2707 1472 2708 1476
rect 2702 1471 2708 1472
rect 2838 1476 2844 1477
rect 2838 1472 2839 1476
rect 2843 1472 2844 1476
rect 2838 1471 2844 1472
rect 2974 1476 2980 1477
rect 2974 1472 2975 1476
rect 2979 1472 2980 1476
rect 2974 1471 2980 1472
rect 3110 1476 3116 1477
rect 3110 1472 3111 1476
rect 3115 1472 3116 1476
rect 3110 1471 3116 1472
rect 3246 1476 3252 1477
rect 3246 1472 3247 1476
rect 3251 1472 3252 1476
rect 3246 1471 3252 1472
rect 3382 1476 3388 1477
rect 3382 1472 3383 1476
rect 3387 1472 3388 1476
rect 3382 1471 3388 1472
rect 3518 1476 3524 1477
rect 3518 1472 3519 1476
rect 3523 1472 3524 1476
rect 3518 1471 3524 1472
rect 3798 1475 3804 1476
rect 3798 1471 3799 1475
rect 3803 1471 3804 1475
rect 2704 1435 2706 1471
rect 2840 1435 2842 1471
rect 2976 1435 2978 1471
rect 3112 1435 3114 1471
rect 3248 1435 3250 1471
rect 3384 1435 3386 1471
rect 3520 1435 3522 1471
rect 3798 1470 3804 1471
rect 3800 1435 3802 1470
rect 2703 1434 2707 1435
rect 2703 1429 2707 1430
rect 2711 1434 2715 1435
rect 2711 1429 2715 1430
rect 2839 1434 2843 1435
rect 2839 1429 2843 1430
rect 2847 1434 2851 1435
rect 2847 1429 2851 1430
rect 2975 1434 2979 1435
rect 2975 1429 2979 1430
rect 2983 1434 2987 1435
rect 2983 1429 2987 1430
rect 3111 1434 3115 1435
rect 3111 1429 3115 1430
rect 3119 1434 3123 1435
rect 3119 1429 3123 1430
rect 3247 1434 3251 1435
rect 3247 1429 3251 1430
rect 3255 1434 3259 1435
rect 3255 1429 3259 1430
rect 3383 1434 3387 1435
rect 3383 1429 3387 1430
rect 3519 1434 3523 1435
rect 3519 1429 3523 1430
rect 3799 1434 3803 1435
rect 3799 1429 3803 1430
rect 2712 1405 2714 1429
rect 2848 1405 2850 1429
rect 2984 1405 2986 1429
rect 3120 1405 3122 1429
rect 3256 1405 3258 1429
rect 3800 1406 3802 1429
rect 3798 1405 3804 1406
rect 2710 1404 2716 1405
rect 2710 1400 2711 1404
rect 2715 1400 2716 1404
rect 2710 1399 2716 1400
rect 2846 1404 2852 1405
rect 2846 1400 2847 1404
rect 2851 1400 2852 1404
rect 2846 1399 2852 1400
rect 2982 1404 2988 1405
rect 2982 1400 2983 1404
rect 2987 1400 2988 1404
rect 2982 1399 2988 1400
rect 3118 1404 3124 1405
rect 3118 1400 3119 1404
rect 3123 1400 3124 1404
rect 3118 1399 3124 1400
rect 3254 1404 3260 1405
rect 3254 1400 3255 1404
rect 3259 1400 3260 1404
rect 3798 1401 3799 1405
rect 3803 1401 3804 1405
rect 3840 1403 3842 1535
rect 4564 1403 4566 1536
rect 4652 1500 4654 1650
rect 4700 1648 4702 1709
rect 4836 1648 4838 1709
rect 4952 1692 4954 1782
rect 4971 1714 4975 1715
rect 4971 1709 4975 1710
rect 5107 1714 5111 1715
rect 5107 1709 5111 1710
rect 5243 1714 5247 1715
rect 5243 1709 5247 1710
rect 5379 1714 5383 1715
rect 5379 1709 5383 1710
rect 4950 1691 4956 1692
rect 4950 1687 4951 1691
rect 4955 1687 4956 1691
rect 4950 1686 4956 1687
rect 4972 1648 4974 1709
rect 5098 1691 5104 1692
rect 5098 1687 5099 1691
rect 5103 1687 5104 1691
rect 5098 1686 5104 1687
rect 5100 1656 5102 1686
rect 5098 1655 5104 1656
rect 5098 1651 5099 1655
rect 5103 1651 5104 1655
rect 5098 1650 5104 1651
rect 5108 1648 5110 1709
rect 5244 1648 5246 1709
rect 5370 1691 5376 1692
rect 5330 1687 5336 1688
rect 5330 1683 5331 1687
rect 5335 1683 5336 1687
rect 5370 1687 5371 1691
rect 5375 1687 5376 1691
rect 5370 1686 5376 1687
rect 5330 1682 5336 1683
rect 5332 1664 5334 1682
rect 5330 1663 5336 1664
rect 5330 1659 5331 1663
rect 5335 1659 5336 1663
rect 5330 1658 5336 1659
rect 5372 1656 5374 1686
rect 5338 1655 5344 1656
rect 5338 1651 5339 1655
rect 5343 1651 5344 1655
rect 5338 1650 5344 1651
rect 5370 1655 5376 1656
rect 5370 1651 5371 1655
rect 5375 1651 5376 1655
rect 5370 1650 5376 1651
rect 4698 1647 4704 1648
rect 4698 1643 4699 1647
rect 4703 1643 4704 1647
rect 4698 1642 4704 1643
rect 4834 1647 4840 1648
rect 4834 1643 4835 1647
rect 4839 1643 4840 1647
rect 4834 1642 4840 1643
rect 4970 1647 4976 1648
rect 4970 1643 4971 1647
rect 4975 1643 4976 1647
rect 4970 1642 4976 1643
rect 5106 1647 5112 1648
rect 5106 1643 5107 1647
rect 5111 1643 5112 1647
rect 5106 1642 5112 1643
rect 5242 1647 5248 1648
rect 5242 1643 5243 1647
rect 5247 1643 5248 1647
rect 5242 1642 5248 1643
rect 4726 1632 4732 1633
rect 4726 1628 4727 1632
rect 4731 1628 4732 1632
rect 4726 1627 4732 1628
rect 4862 1632 4868 1633
rect 4862 1628 4863 1632
rect 4867 1628 4868 1632
rect 4862 1627 4868 1628
rect 4998 1632 5004 1633
rect 4998 1628 4999 1632
rect 5003 1628 5004 1632
rect 4998 1627 5004 1628
rect 5134 1632 5140 1633
rect 5134 1628 5135 1632
rect 5139 1628 5140 1632
rect 5134 1627 5140 1628
rect 5270 1632 5276 1633
rect 5270 1628 5271 1632
rect 5275 1628 5276 1632
rect 5270 1627 5276 1628
rect 4728 1587 4730 1627
rect 4864 1587 4866 1627
rect 5000 1587 5002 1627
rect 5136 1587 5138 1627
rect 5272 1587 5274 1627
rect 4727 1586 4731 1587
rect 4727 1581 4731 1582
rect 4863 1586 4867 1587
rect 4863 1581 4867 1582
rect 4999 1586 5003 1587
rect 4999 1581 5003 1582
rect 5135 1586 5139 1587
rect 5135 1581 5139 1582
rect 5271 1586 5275 1587
rect 5271 1581 5275 1582
rect 4728 1557 4730 1581
rect 4864 1557 4866 1581
rect 5000 1557 5002 1581
rect 5136 1557 5138 1581
rect 5272 1557 5274 1581
rect 4726 1556 4732 1557
rect 4726 1552 4727 1556
rect 4731 1552 4732 1556
rect 4726 1551 4732 1552
rect 4862 1556 4868 1557
rect 4862 1552 4863 1556
rect 4867 1552 4868 1556
rect 4862 1551 4868 1552
rect 4998 1556 5004 1557
rect 4998 1552 4999 1556
rect 5003 1552 5004 1556
rect 4998 1551 5004 1552
rect 5134 1556 5140 1557
rect 5134 1552 5135 1556
rect 5139 1552 5140 1556
rect 5134 1551 5140 1552
rect 5270 1556 5276 1557
rect 5270 1552 5271 1556
rect 5275 1552 5276 1556
rect 5270 1551 5276 1552
rect 4698 1541 4704 1542
rect 4698 1537 4699 1541
rect 4703 1537 4704 1541
rect 4698 1536 4704 1537
rect 4834 1541 4840 1542
rect 4834 1537 4835 1541
rect 4839 1537 4840 1541
rect 4834 1536 4840 1537
rect 4970 1541 4976 1542
rect 4970 1537 4971 1541
rect 4975 1537 4976 1541
rect 4970 1536 4976 1537
rect 5106 1541 5112 1542
rect 5106 1537 5107 1541
rect 5111 1537 5112 1541
rect 5106 1536 5112 1537
rect 5242 1541 5248 1542
rect 5242 1537 5243 1541
rect 5247 1537 5248 1541
rect 5242 1536 5248 1537
rect 4650 1499 4656 1500
rect 4650 1495 4651 1499
rect 4655 1495 4656 1499
rect 4650 1494 4656 1495
rect 4700 1403 4702 1536
rect 4714 1531 4720 1532
rect 4714 1527 4715 1531
rect 4719 1527 4720 1531
rect 4714 1526 4720 1527
rect 4716 1500 4718 1526
rect 4714 1499 4720 1500
rect 4714 1495 4715 1499
rect 4719 1495 4720 1499
rect 4714 1494 4720 1495
rect 4836 1403 4838 1536
rect 4850 1531 4856 1532
rect 4850 1527 4851 1531
rect 4855 1527 4856 1531
rect 4850 1526 4856 1527
rect 4852 1500 4854 1526
rect 4850 1499 4856 1500
rect 4850 1495 4851 1499
rect 4855 1495 4856 1499
rect 4850 1494 4856 1495
rect 4972 1403 4974 1536
rect 4986 1531 4992 1532
rect 4986 1527 4987 1531
rect 4991 1527 4992 1531
rect 4986 1526 4992 1527
rect 4988 1500 4990 1526
rect 4986 1499 4992 1500
rect 4986 1495 4987 1499
rect 4991 1495 4992 1499
rect 4986 1494 4992 1495
rect 5108 1403 5110 1536
rect 5122 1531 5128 1532
rect 5122 1527 5123 1531
rect 5127 1527 5128 1531
rect 5122 1526 5128 1527
rect 5124 1500 5126 1526
rect 5122 1499 5128 1500
rect 5122 1495 5123 1499
rect 5127 1495 5128 1499
rect 5122 1494 5128 1495
rect 5244 1403 5246 1536
rect 5258 1531 5264 1532
rect 5258 1527 5259 1531
rect 5263 1527 5264 1531
rect 5258 1526 5264 1527
rect 5260 1500 5262 1526
rect 5340 1500 5342 1650
rect 5380 1648 5382 1709
rect 5504 1656 5506 1974
rect 5515 1954 5519 1955
rect 5515 1949 5519 1950
rect 5516 1888 5518 1949
rect 5620 1932 5622 2134
rect 5664 2133 5666 2193
rect 5662 2132 5668 2133
rect 5662 2128 5663 2132
rect 5667 2128 5668 2132
rect 5662 2127 5668 2128
rect 5662 2115 5668 2116
rect 5662 2111 5663 2115
rect 5667 2111 5668 2115
rect 5662 2110 5668 2111
rect 5664 2067 5666 2110
rect 5663 2066 5667 2067
rect 5663 2061 5667 2062
rect 5664 2038 5666 2061
rect 5662 2037 5668 2038
rect 5662 2033 5663 2037
rect 5667 2033 5668 2037
rect 5662 2032 5668 2033
rect 5662 2020 5668 2021
rect 5662 2016 5663 2020
rect 5667 2016 5668 2020
rect 5662 2015 5668 2016
rect 5664 1955 5666 2015
rect 5663 1954 5667 1955
rect 5663 1949 5667 1950
rect 5618 1931 5624 1932
rect 5618 1927 5619 1931
rect 5623 1927 5624 1931
rect 5618 1926 5624 1927
rect 5618 1895 5624 1896
rect 5618 1891 5619 1895
rect 5623 1891 5624 1895
rect 5618 1890 5624 1891
rect 5514 1887 5520 1888
rect 5514 1883 5515 1887
rect 5519 1883 5520 1887
rect 5514 1882 5520 1883
rect 5542 1872 5548 1873
rect 5542 1868 5543 1872
rect 5547 1868 5548 1872
rect 5542 1867 5548 1868
rect 5544 1843 5546 1867
rect 5543 1842 5547 1843
rect 5543 1837 5547 1838
rect 5515 1714 5519 1715
rect 5515 1709 5519 1710
rect 5502 1655 5508 1656
rect 5502 1651 5503 1655
rect 5507 1651 5508 1655
rect 5502 1650 5508 1651
rect 5516 1648 5518 1709
rect 5620 1692 5622 1890
rect 5664 1889 5666 1949
rect 5662 1888 5668 1889
rect 5662 1884 5663 1888
rect 5667 1884 5668 1888
rect 5662 1883 5668 1884
rect 5662 1871 5668 1872
rect 5662 1867 5663 1871
rect 5667 1867 5668 1871
rect 5662 1866 5668 1867
rect 5664 1843 5666 1866
rect 5663 1842 5667 1843
rect 5663 1837 5667 1838
rect 5664 1814 5666 1837
rect 5662 1813 5668 1814
rect 5662 1809 5663 1813
rect 5667 1809 5668 1813
rect 5662 1808 5668 1809
rect 5662 1796 5668 1797
rect 5662 1792 5663 1796
rect 5667 1792 5668 1796
rect 5662 1791 5668 1792
rect 5664 1715 5666 1791
rect 5663 1714 5667 1715
rect 5663 1709 5667 1710
rect 5618 1691 5624 1692
rect 5618 1687 5619 1691
rect 5623 1687 5624 1691
rect 5618 1686 5624 1687
rect 5664 1649 5666 1709
rect 5662 1648 5668 1649
rect 5378 1647 5384 1648
rect 5378 1643 5379 1647
rect 5383 1643 5384 1647
rect 5378 1642 5384 1643
rect 5514 1647 5520 1648
rect 5514 1643 5515 1647
rect 5519 1643 5520 1647
rect 5662 1644 5663 1648
rect 5667 1644 5668 1648
rect 5662 1643 5668 1644
rect 5514 1642 5520 1643
rect 5406 1632 5412 1633
rect 5406 1628 5407 1632
rect 5411 1628 5412 1632
rect 5406 1627 5412 1628
rect 5542 1632 5548 1633
rect 5542 1628 5543 1632
rect 5547 1628 5548 1632
rect 5542 1627 5548 1628
rect 5662 1631 5668 1632
rect 5662 1627 5663 1631
rect 5667 1627 5668 1631
rect 5408 1587 5410 1627
rect 5544 1587 5546 1627
rect 5662 1626 5668 1627
rect 5664 1587 5666 1626
rect 5407 1586 5411 1587
rect 5407 1581 5411 1582
rect 5543 1586 5547 1587
rect 5543 1581 5547 1582
rect 5663 1586 5667 1587
rect 5663 1581 5667 1582
rect 5408 1557 5410 1581
rect 5544 1557 5546 1581
rect 5664 1558 5666 1581
rect 5662 1557 5668 1558
rect 5406 1556 5412 1557
rect 5406 1552 5407 1556
rect 5411 1552 5412 1556
rect 5406 1551 5412 1552
rect 5542 1556 5548 1557
rect 5542 1552 5543 1556
rect 5547 1552 5548 1556
rect 5662 1553 5663 1557
rect 5667 1553 5668 1557
rect 5662 1552 5668 1553
rect 5542 1551 5548 1552
rect 5378 1541 5384 1542
rect 5378 1537 5379 1541
rect 5383 1537 5384 1541
rect 5378 1536 5384 1537
rect 5514 1541 5520 1542
rect 5514 1537 5515 1541
rect 5519 1537 5520 1541
rect 5514 1536 5520 1537
rect 5662 1540 5668 1541
rect 5662 1536 5663 1540
rect 5667 1536 5668 1540
rect 5258 1499 5264 1500
rect 5258 1495 5259 1499
rect 5263 1495 5264 1499
rect 5258 1494 5264 1495
rect 5338 1499 5344 1500
rect 5338 1495 5339 1499
rect 5343 1495 5344 1499
rect 5338 1494 5344 1495
rect 5380 1403 5382 1536
rect 5516 1403 5518 1536
rect 5662 1535 5668 1536
rect 5530 1531 5536 1532
rect 5530 1527 5531 1531
rect 5535 1527 5536 1531
rect 5530 1526 5536 1527
rect 5532 1500 5534 1526
rect 5530 1499 5536 1500
rect 5530 1495 5531 1499
rect 5535 1495 5536 1499
rect 5530 1494 5536 1495
rect 5664 1403 5666 1535
rect 3798 1400 3804 1401
rect 3839 1402 3843 1403
rect 3254 1399 3260 1400
rect 3839 1397 3843 1398
rect 4563 1402 4567 1403
rect 4563 1397 4567 1398
rect 4699 1402 4703 1403
rect 4699 1397 4703 1398
rect 4811 1402 4815 1403
rect 4811 1397 4815 1398
rect 4835 1402 4839 1403
rect 4835 1397 4839 1398
rect 4947 1402 4951 1403
rect 4947 1397 4951 1398
rect 4971 1402 4975 1403
rect 4971 1397 4975 1398
rect 5083 1402 5087 1403
rect 5083 1397 5087 1398
rect 5107 1402 5111 1403
rect 5107 1397 5111 1398
rect 5219 1402 5223 1403
rect 5219 1397 5223 1398
rect 5243 1402 5247 1403
rect 5243 1397 5247 1398
rect 5355 1402 5359 1403
rect 5355 1397 5359 1398
rect 5379 1402 5383 1403
rect 5379 1397 5383 1398
rect 5491 1402 5495 1403
rect 5491 1397 5495 1398
rect 5515 1402 5519 1403
rect 5515 1397 5519 1398
rect 5663 1402 5667 1403
rect 5663 1397 5667 1398
rect 2682 1389 2688 1390
rect 2682 1385 2683 1389
rect 2687 1385 2688 1389
rect 2682 1384 2688 1385
rect 2818 1389 2824 1390
rect 2818 1385 2819 1389
rect 2823 1385 2824 1389
rect 2818 1384 2824 1385
rect 2954 1389 2960 1390
rect 2954 1385 2955 1389
rect 2959 1385 2960 1389
rect 2954 1384 2960 1385
rect 3090 1389 3096 1390
rect 3090 1385 3091 1389
rect 3095 1385 3096 1389
rect 3090 1384 3096 1385
rect 3226 1389 3232 1390
rect 3226 1385 3227 1389
rect 3231 1385 3232 1389
rect 3226 1384 3232 1385
rect 3798 1388 3804 1389
rect 3798 1384 3799 1388
rect 3803 1384 3804 1388
rect 2634 1347 2640 1348
rect 2634 1343 2635 1347
rect 2639 1343 2640 1347
rect 2634 1342 2640 1343
rect 2684 1323 2686 1384
rect 2698 1379 2704 1380
rect 2698 1375 2699 1379
rect 2703 1375 2704 1379
rect 2698 1374 2704 1375
rect 2700 1348 2702 1374
rect 2698 1347 2704 1348
rect 2698 1343 2699 1347
rect 2703 1343 2704 1347
rect 2698 1342 2704 1343
rect 2820 1323 2822 1384
rect 2834 1379 2840 1380
rect 2834 1375 2835 1379
rect 2839 1375 2840 1379
rect 2834 1374 2840 1375
rect 2836 1348 2838 1374
rect 2834 1347 2840 1348
rect 2834 1343 2835 1347
rect 2839 1343 2840 1347
rect 2834 1342 2840 1343
rect 2956 1323 2958 1384
rect 2970 1379 2976 1380
rect 2970 1375 2971 1379
rect 2975 1375 2976 1379
rect 2970 1374 2976 1375
rect 2972 1348 2974 1374
rect 2970 1347 2976 1348
rect 2970 1343 2971 1347
rect 2975 1343 2976 1347
rect 2970 1342 2976 1343
rect 3092 1323 3094 1384
rect 3106 1379 3112 1380
rect 3106 1375 3107 1379
rect 3111 1375 3112 1379
rect 3106 1374 3112 1375
rect 3108 1348 3110 1374
rect 3106 1347 3112 1348
rect 3106 1343 3107 1347
rect 3111 1343 3112 1347
rect 3106 1342 3112 1343
rect 3228 1323 3230 1384
rect 3798 1383 3804 1384
rect 3242 1379 3248 1380
rect 3242 1375 3243 1379
rect 3247 1375 3248 1379
rect 3242 1374 3248 1375
rect 3354 1379 3360 1380
rect 3354 1375 3355 1379
rect 3359 1375 3360 1379
rect 3354 1374 3360 1375
rect 3244 1348 3246 1374
rect 3242 1347 3248 1348
rect 3242 1343 3243 1347
rect 3247 1343 3248 1347
rect 3242 1342 3248 1343
rect 2547 1322 2551 1323
rect 2547 1317 2551 1318
rect 2555 1322 2559 1323
rect 2555 1317 2559 1318
rect 2683 1322 2687 1323
rect 2683 1317 2687 1318
rect 2715 1322 2719 1323
rect 2715 1317 2719 1318
rect 2819 1322 2823 1323
rect 2819 1317 2823 1318
rect 2891 1322 2895 1323
rect 2891 1317 2895 1318
rect 2955 1322 2959 1323
rect 2955 1317 2959 1318
rect 3075 1322 3079 1323
rect 3075 1317 3079 1318
rect 3091 1322 3095 1323
rect 3091 1317 3095 1318
rect 3227 1322 3231 1323
rect 3227 1317 3231 1318
rect 3267 1322 3271 1323
rect 3267 1317 3271 1318
rect 2499 1300 2503 1301
rect 2499 1295 2503 1296
rect 2530 1299 2536 1300
rect 2530 1295 2531 1299
rect 2535 1295 2536 1299
rect 2530 1294 2536 1295
rect 2532 1264 2534 1294
rect 2530 1263 2536 1264
rect 2530 1259 2531 1263
rect 2535 1259 2536 1263
rect 2530 1258 2536 1259
rect 2556 1256 2558 1317
rect 2706 1299 2712 1300
rect 2706 1295 2707 1299
rect 2711 1295 2712 1299
rect 2706 1294 2712 1295
rect 2708 1264 2710 1294
rect 2706 1263 2712 1264
rect 2706 1259 2707 1263
rect 2711 1259 2712 1263
rect 2706 1258 2712 1259
rect 2716 1256 2718 1317
rect 2723 1300 2727 1301
rect 2723 1295 2727 1296
rect 2724 1264 2726 1295
rect 2722 1263 2728 1264
rect 2722 1259 2723 1263
rect 2727 1259 2728 1263
rect 2722 1258 2728 1259
rect 2892 1256 2894 1317
rect 3014 1263 3020 1264
rect 3014 1259 3015 1263
rect 3019 1259 3020 1263
rect 3014 1258 3020 1259
rect 2266 1255 2272 1256
rect 2266 1251 2267 1255
rect 2271 1251 2272 1255
rect 2266 1250 2272 1251
rect 2402 1255 2408 1256
rect 2402 1251 2403 1255
rect 2407 1251 2408 1255
rect 2402 1250 2408 1251
rect 2554 1255 2560 1256
rect 2554 1251 2555 1255
rect 2559 1251 2560 1255
rect 2554 1250 2560 1251
rect 2714 1255 2720 1256
rect 2714 1251 2715 1255
rect 2719 1251 2720 1255
rect 2714 1250 2720 1251
rect 2890 1255 2896 1256
rect 2890 1251 2891 1255
rect 2895 1251 2896 1255
rect 2890 1250 2896 1251
rect 2294 1240 2300 1241
rect 2294 1236 2295 1240
rect 2299 1236 2300 1240
rect 2294 1235 2300 1236
rect 2430 1240 2436 1241
rect 2430 1236 2431 1240
rect 2435 1236 2436 1240
rect 2430 1235 2436 1236
rect 2582 1240 2588 1241
rect 2582 1236 2583 1240
rect 2587 1236 2588 1240
rect 2582 1235 2588 1236
rect 2742 1240 2748 1241
rect 2742 1236 2743 1240
rect 2747 1236 2748 1240
rect 2742 1235 2748 1236
rect 2918 1240 2924 1241
rect 2918 1236 2919 1240
rect 2923 1236 2924 1240
rect 2918 1235 2924 1236
rect 2246 1215 2252 1216
rect 2246 1211 2247 1215
rect 2251 1211 2252 1215
rect 2296 1211 2298 1235
rect 2432 1211 2434 1235
rect 2584 1211 2586 1235
rect 2744 1211 2746 1235
rect 2920 1211 2922 1235
rect 1975 1210 1979 1211
rect 1975 1205 1979 1206
rect 2023 1210 2027 1211
rect 2023 1205 2027 1206
rect 2159 1210 2163 1211
rect 2159 1205 2163 1206
rect 2239 1210 2243 1211
rect 2246 1210 2252 1211
rect 2295 1210 2299 1211
rect 2239 1205 2243 1206
rect 2295 1205 2299 1206
rect 2431 1210 2435 1211
rect 2431 1205 2435 1206
rect 2479 1210 2483 1211
rect 2479 1205 2483 1206
rect 2583 1210 2587 1211
rect 2583 1205 2587 1206
rect 2719 1210 2723 1211
rect 2719 1205 2723 1206
rect 2743 1210 2747 1211
rect 2919 1210 2923 1211
rect 2743 1205 2747 1206
rect 2810 1207 2816 1208
rect 563 1186 567 1187
rect 563 1181 567 1182
rect 747 1186 751 1187
rect 747 1181 751 1182
rect 803 1186 807 1187
rect 803 1181 807 1182
rect 1043 1186 1047 1187
rect 1043 1181 1047 1182
rect 1067 1186 1071 1187
rect 1067 1181 1071 1182
rect 1283 1186 1287 1187
rect 1283 1181 1287 1182
rect 1395 1186 1399 1187
rect 1395 1181 1399 1182
rect 1523 1186 1527 1187
rect 1523 1181 1527 1182
rect 1771 1186 1775 1187
rect 1771 1181 1775 1182
rect 1935 1186 1939 1187
rect 1976 1182 1978 1205
rect 1935 1181 1939 1182
rect 1974 1181 1980 1182
rect 2024 1181 2026 1205
rect 2240 1181 2242 1205
rect 2480 1181 2482 1205
rect 2720 1181 2722 1205
rect 2810 1203 2811 1207
rect 2815 1203 2816 1207
rect 2919 1205 2923 1206
rect 2959 1210 2963 1211
rect 2959 1205 2963 1206
rect 2810 1202 2816 1203
rect 458 1127 464 1128
rect 458 1123 459 1127
rect 463 1123 464 1127
rect 458 1122 464 1123
rect 514 1127 520 1128
rect 514 1123 515 1127
rect 519 1123 520 1127
rect 514 1122 520 1123
rect 564 1120 566 1181
rect 804 1120 806 1181
rect 938 1127 944 1128
rect 938 1123 939 1127
rect 943 1123 944 1127
rect 938 1122 944 1123
rect 330 1119 336 1120
rect 330 1115 331 1119
rect 335 1115 336 1119
rect 330 1114 336 1115
rect 562 1119 568 1120
rect 562 1115 563 1119
rect 567 1115 568 1119
rect 562 1114 568 1115
rect 802 1119 808 1120
rect 802 1115 803 1119
rect 807 1115 808 1119
rect 802 1114 808 1115
rect 358 1104 364 1105
rect 358 1100 359 1104
rect 363 1100 364 1104
rect 358 1099 364 1100
rect 590 1104 596 1105
rect 590 1100 591 1104
rect 595 1100 596 1104
rect 590 1099 596 1100
rect 830 1104 836 1105
rect 830 1100 831 1104
rect 835 1100 836 1104
rect 830 1099 836 1100
rect 360 1075 362 1099
rect 592 1075 594 1099
rect 832 1075 834 1099
rect 359 1074 363 1075
rect 359 1069 363 1070
rect 439 1074 443 1075
rect 439 1069 443 1070
rect 591 1074 595 1075
rect 591 1069 595 1070
rect 615 1074 619 1075
rect 615 1069 619 1070
rect 783 1074 787 1075
rect 783 1069 787 1070
rect 831 1074 835 1075
rect 831 1069 835 1070
rect 440 1045 442 1069
rect 616 1045 618 1069
rect 784 1045 786 1069
rect 438 1044 444 1045
rect 438 1040 439 1044
rect 443 1040 444 1044
rect 438 1039 444 1040
rect 614 1044 620 1045
rect 614 1040 615 1044
rect 619 1040 620 1044
rect 614 1039 620 1040
rect 782 1044 788 1045
rect 782 1040 783 1044
rect 787 1040 788 1044
rect 782 1039 788 1040
rect 410 1029 416 1030
rect 410 1025 411 1029
rect 415 1025 416 1029
rect 410 1024 416 1025
rect 586 1029 592 1030
rect 586 1025 587 1029
rect 591 1025 592 1029
rect 586 1024 592 1025
rect 754 1029 760 1030
rect 754 1025 755 1029
rect 759 1025 760 1029
rect 754 1024 760 1025
rect 922 1029 928 1030
rect 922 1025 923 1029
rect 927 1025 928 1029
rect 922 1024 928 1025
rect 270 1019 276 1020
rect 270 1015 271 1019
rect 275 1015 276 1019
rect 270 1014 276 1015
rect 412 959 414 1024
rect 498 987 504 988
rect 498 983 499 987
rect 503 983 504 987
rect 498 982 504 983
rect 111 958 115 959
rect 111 953 115 954
rect 227 958 231 959
rect 227 953 231 954
rect 235 958 239 959
rect 235 953 239 954
rect 379 958 383 959
rect 379 953 383 954
rect 411 958 415 959
rect 411 953 415 954
rect 112 893 114 953
rect 110 892 116 893
rect 228 892 230 953
rect 354 935 360 936
rect 314 931 320 932
rect 314 927 315 931
rect 319 927 320 931
rect 354 931 355 935
rect 359 931 360 935
rect 354 930 360 931
rect 314 926 320 927
rect 110 888 111 892
rect 115 888 116 892
rect 110 887 116 888
rect 226 891 232 892
rect 226 887 227 891
rect 231 887 232 891
rect 226 886 232 887
rect 254 876 260 877
rect 110 875 116 876
rect 110 871 111 875
rect 115 871 116 875
rect 254 872 255 876
rect 259 872 260 876
rect 254 871 260 872
rect 110 870 116 871
rect 112 831 114 870
rect 256 831 258 871
rect 111 830 115 831
rect 111 825 115 826
rect 255 830 259 831
rect 255 825 259 826
rect 112 802 114 825
rect 110 801 116 802
rect 110 797 111 801
rect 115 797 116 801
rect 110 796 116 797
rect 110 784 116 785
rect 110 780 111 784
rect 115 780 116 784
rect 110 779 116 780
rect 112 719 114 779
rect 316 768 318 926
rect 356 900 358 930
rect 354 899 360 900
rect 354 895 355 899
rect 359 895 360 899
rect 354 894 360 895
rect 380 892 382 953
rect 500 900 502 982
rect 588 959 590 1024
rect 658 1019 664 1020
rect 658 1015 659 1019
rect 663 1015 664 1019
rect 658 1014 664 1015
rect 746 1019 752 1020
rect 746 1015 747 1019
rect 751 1015 752 1019
rect 746 1014 752 1015
rect 539 958 543 959
rect 539 953 543 954
rect 587 958 591 959
rect 587 953 591 954
rect 498 899 504 900
rect 498 895 499 899
rect 503 895 504 899
rect 498 894 504 895
rect 540 892 542 953
rect 660 936 662 1014
rect 748 988 750 1014
rect 746 987 752 988
rect 746 983 747 987
rect 751 983 752 987
rect 746 982 752 983
rect 756 959 758 1024
rect 910 1019 916 1020
rect 910 1015 911 1019
rect 915 1015 916 1019
rect 910 1014 916 1015
rect 912 988 914 1014
rect 910 987 916 988
rect 910 983 911 987
rect 915 983 916 987
rect 910 982 916 983
rect 924 959 926 1024
rect 940 988 942 1122
rect 1044 1120 1046 1181
rect 1284 1120 1286 1181
rect 1524 1120 1526 1181
rect 1650 1163 1656 1164
rect 1650 1159 1651 1163
rect 1655 1159 1656 1163
rect 1650 1158 1656 1159
rect 1652 1128 1654 1158
rect 1758 1155 1764 1156
rect 1758 1151 1759 1155
rect 1763 1151 1764 1155
rect 1758 1150 1764 1151
rect 1650 1127 1656 1128
rect 1650 1123 1651 1127
rect 1655 1123 1656 1127
rect 1650 1122 1656 1123
rect 1042 1119 1048 1120
rect 1042 1115 1043 1119
rect 1047 1115 1048 1119
rect 1042 1114 1048 1115
rect 1282 1119 1288 1120
rect 1282 1115 1283 1119
rect 1287 1115 1288 1119
rect 1282 1114 1288 1115
rect 1522 1119 1528 1120
rect 1522 1115 1523 1119
rect 1527 1115 1528 1119
rect 1522 1114 1528 1115
rect 1070 1104 1076 1105
rect 1070 1100 1071 1104
rect 1075 1100 1076 1104
rect 1070 1099 1076 1100
rect 1310 1104 1316 1105
rect 1310 1100 1311 1104
rect 1315 1100 1316 1104
rect 1310 1099 1316 1100
rect 1550 1104 1556 1105
rect 1550 1100 1551 1104
rect 1555 1100 1556 1104
rect 1550 1099 1556 1100
rect 1072 1075 1074 1099
rect 1312 1075 1314 1099
rect 1552 1075 1554 1099
rect 951 1074 955 1075
rect 951 1069 955 1070
rect 1071 1074 1075 1075
rect 1071 1069 1075 1070
rect 1111 1074 1115 1075
rect 1111 1069 1115 1070
rect 1271 1074 1275 1075
rect 1271 1069 1275 1070
rect 1311 1074 1315 1075
rect 1311 1069 1315 1070
rect 1431 1074 1435 1075
rect 1431 1069 1435 1070
rect 1551 1074 1555 1075
rect 1551 1069 1555 1070
rect 1591 1074 1595 1075
rect 1591 1069 1595 1070
rect 1751 1074 1755 1075
rect 1751 1069 1755 1070
rect 952 1045 954 1069
rect 1112 1045 1114 1069
rect 1272 1045 1274 1069
rect 1432 1045 1434 1069
rect 1592 1045 1594 1069
rect 1752 1045 1754 1069
rect 950 1044 956 1045
rect 950 1040 951 1044
rect 955 1040 956 1044
rect 950 1039 956 1040
rect 1110 1044 1116 1045
rect 1110 1040 1111 1044
rect 1115 1040 1116 1044
rect 1110 1039 1116 1040
rect 1270 1044 1276 1045
rect 1270 1040 1271 1044
rect 1275 1040 1276 1044
rect 1270 1039 1276 1040
rect 1430 1044 1436 1045
rect 1430 1040 1431 1044
rect 1435 1040 1436 1044
rect 1430 1039 1436 1040
rect 1590 1044 1596 1045
rect 1590 1040 1591 1044
rect 1595 1040 1596 1044
rect 1590 1039 1596 1040
rect 1750 1044 1756 1045
rect 1750 1040 1751 1044
rect 1755 1040 1756 1044
rect 1750 1039 1756 1040
rect 1082 1029 1088 1030
rect 1082 1025 1083 1029
rect 1087 1025 1088 1029
rect 1082 1024 1088 1025
rect 1242 1029 1248 1030
rect 1242 1025 1243 1029
rect 1247 1025 1248 1029
rect 1242 1024 1248 1025
rect 1402 1029 1408 1030
rect 1402 1025 1403 1029
rect 1407 1025 1408 1029
rect 1402 1024 1408 1025
rect 1562 1029 1568 1030
rect 1562 1025 1563 1029
rect 1567 1025 1568 1029
rect 1562 1024 1568 1025
rect 1722 1029 1728 1030
rect 1722 1025 1723 1029
rect 1727 1025 1728 1029
rect 1722 1024 1728 1025
rect 938 987 944 988
rect 938 983 939 987
rect 943 983 944 987
rect 938 982 944 983
rect 1084 959 1086 1024
rect 1244 959 1246 1024
rect 1258 1019 1264 1020
rect 1258 1015 1259 1019
rect 1263 1015 1264 1019
rect 1258 1014 1264 1015
rect 1260 988 1262 1014
rect 1258 987 1264 988
rect 1258 983 1259 987
rect 1263 983 1264 987
rect 1258 982 1264 983
rect 1404 959 1406 1024
rect 1418 1019 1424 1020
rect 1418 1015 1419 1019
rect 1423 1015 1424 1019
rect 1418 1014 1424 1015
rect 1420 988 1422 1014
rect 1418 987 1424 988
rect 1418 983 1419 987
rect 1423 983 1424 987
rect 1418 982 1424 983
rect 1564 959 1566 1024
rect 1578 1019 1584 1020
rect 1578 1015 1579 1019
rect 1583 1015 1584 1019
rect 1578 1014 1584 1015
rect 1580 988 1582 1014
rect 1578 987 1584 988
rect 1578 983 1579 987
rect 1583 983 1584 987
rect 1578 982 1584 983
rect 1724 959 1726 1024
rect 1760 1020 1762 1150
rect 1772 1120 1774 1181
rect 1936 1121 1938 1181
rect 1974 1177 1975 1181
rect 1979 1177 1980 1181
rect 1974 1176 1980 1177
rect 2022 1180 2028 1181
rect 2022 1176 2023 1180
rect 2027 1176 2028 1180
rect 2022 1175 2028 1176
rect 2238 1180 2244 1181
rect 2238 1176 2239 1180
rect 2243 1176 2244 1180
rect 2238 1175 2244 1176
rect 2478 1180 2484 1181
rect 2478 1176 2479 1180
rect 2483 1176 2484 1180
rect 2478 1175 2484 1176
rect 2718 1180 2724 1181
rect 2718 1176 2719 1180
rect 2723 1176 2724 1180
rect 2718 1175 2724 1176
rect 1994 1165 2000 1166
rect 1974 1164 1980 1165
rect 1974 1160 1975 1164
rect 1979 1160 1980 1164
rect 1994 1161 1995 1165
rect 1999 1161 2000 1165
rect 1994 1160 2000 1161
rect 2210 1165 2216 1166
rect 2210 1161 2211 1165
rect 2215 1161 2216 1165
rect 2210 1160 2216 1161
rect 2450 1165 2456 1166
rect 2450 1161 2451 1165
rect 2455 1161 2456 1165
rect 2450 1160 2456 1161
rect 2690 1165 2696 1166
rect 2690 1161 2691 1165
rect 2695 1161 2696 1165
rect 2690 1160 2696 1161
rect 1974 1159 1980 1160
rect 1934 1120 1940 1121
rect 1770 1119 1776 1120
rect 1770 1115 1771 1119
rect 1775 1115 1776 1119
rect 1934 1116 1935 1120
rect 1939 1116 1940 1120
rect 1934 1115 1940 1116
rect 1770 1114 1776 1115
rect 1798 1104 1804 1105
rect 1798 1100 1799 1104
rect 1803 1100 1804 1104
rect 1798 1099 1804 1100
rect 1934 1103 1940 1104
rect 1934 1099 1935 1103
rect 1939 1099 1940 1103
rect 1800 1075 1802 1099
rect 1934 1098 1940 1099
rect 1936 1075 1938 1098
rect 1976 1075 1978 1159
rect 1996 1075 1998 1160
rect 2212 1075 2214 1160
rect 2226 1155 2232 1156
rect 2226 1151 2227 1155
rect 2231 1151 2232 1155
rect 2226 1150 2232 1151
rect 2228 1124 2230 1150
rect 2226 1123 2232 1124
rect 2226 1119 2227 1123
rect 2231 1119 2232 1123
rect 2226 1118 2232 1119
rect 2452 1075 2454 1160
rect 2466 1155 2472 1156
rect 2466 1151 2467 1155
rect 2471 1151 2472 1155
rect 2466 1150 2472 1151
rect 2468 1124 2470 1150
rect 2466 1123 2472 1124
rect 2466 1119 2467 1123
rect 2471 1119 2472 1123
rect 2466 1118 2472 1119
rect 2692 1075 2694 1160
rect 2812 1156 2814 1202
rect 2960 1181 2962 1205
rect 2958 1180 2964 1181
rect 2958 1176 2959 1180
rect 2963 1176 2964 1180
rect 2958 1175 2964 1176
rect 2930 1165 2936 1166
rect 2930 1161 2931 1165
rect 2935 1161 2936 1165
rect 2930 1160 2936 1161
rect 2706 1155 2712 1156
rect 2706 1151 2707 1155
rect 2711 1151 2712 1155
rect 2706 1150 2712 1151
rect 2810 1155 2816 1156
rect 2810 1151 2811 1155
rect 2815 1151 2816 1155
rect 2810 1150 2816 1151
rect 2708 1124 2710 1150
rect 2706 1123 2712 1124
rect 2706 1119 2707 1123
rect 2711 1119 2712 1123
rect 2706 1118 2712 1119
rect 2932 1075 2934 1160
rect 3016 1124 3018 1258
rect 3076 1256 3078 1317
rect 3268 1256 3270 1317
rect 3356 1296 3358 1374
rect 3800 1323 3802 1383
rect 3840 1337 3842 1397
rect 3838 1336 3844 1337
rect 4812 1336 4814 1397
rect 4934 1343 4940 1344
rect 4934 1339 4935 1343
rect 4939 1339 4940 1343
rect 4934 1338 4940 1339
rect 3838 1332 3839 1336
rect 3843 1332 3844 1336
rect 3838 1331 3844 1332
rect 4810 1335 4816 1336
rect 4810 1331 4811 1335
rect 4815 1331 4816 1335
rect 4810 1330 4816 1331
rect 3467 1322 3471 1323
rect 3467 1317 3471 1318
rect 3651 1322 3655 1323
rect 3651 1317 3655 1318
rect 3799 1322 3803 1323
rect 4838 1320 4844 1321
rect 3799 1317 3803 1318
rect 3838 1319 3844 1320
rect 3354 1295 3360 1296
rect 3354 1291 3355 1295
rect 3359 1291 3360 1295
rect 3354 1290 3360 1291
rect 3468 1256 3470 1317
rect 3594 1299 3600 1300
rect 3554 1295 3560 1296
rect 3554 1291 3555 1295
rect 3559 1291 3560 1295
rect 3594 1295 3595 1299
rect 3599 1295 3600 1299
rect 3594 1294 3600 1295
rect 3554 1290 3560 1291
rect 3074 1255 3080 1256
rect 3074 1251 3075 1255
rect 3079 1251 3080 1255
rect 3074 1250 3080 1251
rect 3266 1255 3272 1256
rect 3266 1251 3267 1255
rect 3271 1251 3272 1255
rect 3266 1250 3272 1251
rect 3466 1255 3472 1256
rect 3466 1251 3467 1255
rect 3471 1251 3472 1255
rect 3466 1250 3472 1251
rect 3102 1240 3108 1241
rect 3102 1236 3103 1240
rect 3107 1236 3108 1240
rect 3102 1235 3108 1236
rect 3294 1240 3300 1241
rect 3294 1236 3295 1240
rect 3299 1236 3300 1240
rect 3294 1235 3300 1236
rect 3494 1240 3500 1241
rect 3494 1236 3495 1240
rect 3499 1236 3500 1240
rect 3494 1235 3500 1236
rect 3104 1211 3106 1235
rect 3296 1211 3298 1235
rect 3496 1211 3498 1235
rect 3103 1210 3107 1211
rect 3103 1205 3107 1206
rect 3207 1210 3211 1211
rect 3207 1205 3211 1206
rect 3295 1210 3299 1211
rect 3295 1205 3299 1206
rect 3455 1210 3459 1211
rect 3455 1205 3459 1206
rect 3495 1210 3499 1211
rect 3495 1205 3499 1206
rect 3208 1181 3210 1205
rect 3456 1181 3458 1205
rect 3206 1180 3212 1181
rect 3206 1176 3207 1180
rect 3211 1176 3212 1180
rect 3206 1175 3212 1176
rect 3454 1180 3460 1181
rect 3454 1176 3455 1180
rect 3459 1176 3460 1180
rect 3454 1175 3460 1176
rect 3178 1165 3184 1166
rect 3178 1161 3179 1165
rect 3183 1161 3184 1165
rect 3178 1160 3184 1161
rect 3426 1165 3432 1166
rect 3426 1161 3427 1165
rect 3431 1161 3432 1165
rect 3426 1160 3432 1161
rect 3082 1155 3088 1156
rect 3082 1151 3083 1155
rect 3087 1151 3088 1155
rect 3082 1150 3088 1151
rect 3014 1123 3020 1124
rect 3014 1119 3015 1123
rect 3019 1119 3020 1123
rect 3014 1118 3020 1119
rect 1799 1074 1803 1075
rect 1799 1069 1803 1070
rect 1935 1074 1939 1075
rect 1935 1069 1939 1070
rect 1975 1074 1979 1075
rect 1975 1069 1979 1070
rect 1995 1074 1999 1075
rect 1995 1069 1999 1070
rect 2211 1074 2215 1075
rect 2211 1069 2215 1070
rect 2451 1074 2455 1075
rect 2451 1069 2455 1070
rect 2691 1074 2695 1075
rect 2691 1069 2695 1070
rect 2931 1074 2935 1075
rect 2931 1069 2935 1070
rect 1936 1046 1938 1069
rect 1934 1045 1940 1046
rect 1934 1041 1935 1045
rect 1939 1041 1940 1045
rect 1934 1040 1940 1041
rect 1934 1028 1940 1029
rect 1934 1024 1935 1028
rect 1939 1024 1940 1028
rect 1934 1023 1940 1024
rect 1738 1019 1744 1020
rect 1738 1015 1739 1019
rect 1743 1015 1744 1019
rect 1738 1014 1744 1015
rect 1758 1019 1764 1020
rect 1758 1015 1759 1019
rect 1763 1015 1764 1019
rect 1758 1014 1764 1015
rect 1740 988 1742 1014
rect 1738 987 1744 988
rect 1738 983 1739 987
rect 1743 983 1744 987
rect 1738 982 1744 983
rect 1936 959 1938 1023
rect 1976 1009 1978 1069
rect 3084 1052 3086 1150
rect 3180 1075 3182 1160
rect 3378 1123 3384 1124
rect 3378 1119 3379 1123
rect 3383 1119 3384 1123
rect 3378 1118 3384 1119
rect 3091 1074 3095 1075
rect 3091 1069 3095 1070
rect 3179 1074 3183 1075
rect 3179 1069 3183 1070
rect 3243 1074 3247 1075
rect 3243 1069 3247 1070
rect 3082 1051 3088 1052
rect 3082 1047 3083 1051
rect 3087 1047 3088 1051
rect 3082 1046 3088 1047
rect 2986 1015 2992 1016
rect 2986 1011 2987 1015
rect 2991 1011 2992 1015
rect 2986 1010 2992 1011
rect 1974 1008 1980 1009
rect 1974 1004 1975 1008
rect 1979 1004 1980 1008
rect 1974 1003 1980 1004
rect 1974 991 1980 992
rect 1974 987 1975 991
rect 1979 987 1980 991
rect 1974 986 1980 987
rect 715 958 719 959
rect 715 953 719 954
rect 755 958 759 959
rect 755 953 759 954
rect 891 958 895 959
rect 891 953 895 954
rect 923 958 927 959
rect 923 953 927 954
rect 1075 958 1079 959
rect 1075 953 1079 954
rect 1083 958 1087 959
rect 1083 953 1087 954
rect 1243 958 1247 959
rect 1243 953 1247 954
rect 1259 958 1263 959
rect 1259 953 1263 954
rect 1403 958 1407 959
rect 1403 953 1407 954
rect 1443 958 1447 959
rect 1443 953 1447 954
rect 1563 958 1567 959
rect 1563 953 1567 954
rect 1627 958 1631 959
rect 1627 953 1631 954
rect 1723 958 1727 959
rect 1723 953 1727 954
rect 1787 958 1791 959
rect 1787 953 1791 954
rect 1935 958 1939 959
rect 1935 953 1939 954
rect 658 935 664 936
rect 658 931 659 935
rect 663 931 664 935
rect 658 930 664 931
rect 666 935 672 936
rect 666 931 667 935
rect 671 931 672 935
rect 666 930 672 931
rect 668 900 670 930
rect 666 899 672 900
rect 666 895 667 899
rect 671 895 672 899
rect 666 894 672 895
rect 716 892 718 953
rect 842 935 848 936
rect 842 931 843 935
rect 847 931 848 935
rect 842 930 848 931
rect 844 900 846 930
rect 842 899 848 900
rect 842 895 843 899
rect 847 895 848 899
rect 842 894 848 895
rect 892 892 894 953
rect 1018 935 1024 936
rect 1018 931 1019 935
rect 1023 931 1024 935
rect 1018 930 1024 931
rect 1020 900 1022 930
rect 1018 899 1024 900
rect 1018 895 1019 899
rect 1023 895 1024 899
rect 1018 894 1024 895
rect 1076 892 1078 953
rect 1226 899 1232 900
rect 1226 895 1227 899
rect 1231 895 1232 899
rect 1226 894 1232 895
rect 378 891 384 892
rect 378 887 379 891
rect 383 887 384 891
rect 378 886 384 887
rect 538 891 544 892
rect 538 887 539 891
rect 543 887 544 891
rect 538 886 544 887
rect 714 891 720 892
rect 714 887 715 891
rect 719 887 720 891
rect 714 886 720 887
rect 890 891 896 892
rect 890 887 891 891
rect 895 887 896 891
rect 890 886 896 887
rect 1074 891 1080 892
rect 1074 887 1075 891
rect 1079 887 1080 891
rect 1074 886 1080 887
rect 406 876 412 877
rect 406 872 407 876
rect 411 872 412 876
rect 406 871 412 872
rect 566 876 572 877
rect 566 872 567 876
rect 571 872 572 876
rect 566 871 572 872
rect 742 876 748 877
rect 742 872 743 876
rect 747 872 748 876
rect 742 871 748 872
rect 918 876 924 877
rect 918 872 919 876
rect 923 872 924 876
rect 918 871 924 872
rect 1102 876 1108 877
rect 1102 872 1103 876
rect 1107 872 1108 876
rect 1102 871 1108 872
rect 408 831 410 871
rect 568 831 570 871
rect 744 831 746 871
rect 920 831 922 871
rect 1104 831 1106 871
rect 375 830 379 831
rect 375 825 379 826
rect 407 830 411 831
rect 407 825 411 826
rect 567 830 571 831
rect 567 825 571 826
rect 655 830 659 831
rect 655 825 659 826
rect 743 830 747 831
rect 743 825 747 826
rect 919 830 923 831
rect 919 825 923 826
rect 943 830 947 831
rect 943 825 947 826
rect 1103 830 1107 831
rect 1103 825 1107 826
rect 376 801 378 825
rect 656 801 658 825
rect 944 801 946 825
rect 374 800 380 801
rect 374 796 375 800
rect 379 796 380 800
rect 374 795 380 796
rect 654 800 660 801
rect 654 796 655 800
rect 659 796 660 800
rect 654 795 660 796
rect 942 800 948 801
rect 942 796 943 800
rect 947 796 948 800
rect 942 795 948 796
rect 346 785 352 786
rect 346 781 347 785
rect 351 781 352 785
rect 346 780 352 781
rect 626 785 632 786
rect 626 781 627 785
rect 631 781 632 785
rect 626 780 632 781
rect 914 785 920 786
rect 914 781 915 785
rect 919 781 920 785
rect 914 780 920 781
rect 1210 785 1216 786
rect 1210 781 1211 785
rect 1215 781 1216 785
rect 1210 780 1216 781
rect 314 767 320 768
rect 314 763 315 767
rect 319 763 320 767
rect 314 762 320 763
rect 348 719 350 780
rect 430 743 436 744
rect 430 739 431 743
rect 435 739 436 743
rect 430 738 436 739
rect 111 718 115 719
rect 111 713 115 714
rect 131 718 135 719
rect 131 713 135 714
rect 307 718 311 719
rect 307 713 311 714
rect 347 718 351 719
rect 347 713 351 714
rect 112 653 114 713
rect 110 652 116 653
rect 132 652 134 713
rect 258 695 264 696
rect 258 691 259 695
rect 263 691 264 695
rect 258 690 264 691
rect 260 660 262 690
rect 258 659 264 660
rect 258 655 259 659
rect 263 655 264 659
rect 258 654 264 655
rect 308 652 310 713
rect 432 660 434 738
rect 628 719 630 780
rect 642 775 648 776
rect 642 771 643 775
rect 647 771 648 775
rect 642 770 648 771
rect 644 744 646 770
rect 642 743 648 744
rect 642 739 643 743
rect 647 739 648 743
rect 642 738 648 739
rect 916 719 918 780
rect 1018 775 1024 776
rect 1018 771 1019 775
rect 1023 771 1024 775
rect 1018 770 1024 771
rect 1134 775 1140 776
rect 1134 771 1135 775
rect 1139 771 1140 775
rect 1134 770 1140 771
rect 499 718 503 719
rect 499 713 503 714
rect 627 718 631 719
rect 627 713 631 714
rect 683 718 687 719
rect 683 713 687 714
rect 859 718 863 719
rect 859 713 863 714
rect 915 718 919 719
rect 915 713 919 714
rect 474 695 480 696
rect 474 691 475 695
rect 479 691 480 695
rect 474 690 480 691
rect 430 659 436 660
rect 430 655 431 659
rect 435 655 436 659
rect 430 654 436 655
rect 110 648 111 652
rect 115 648 116 652
rect 110 647 116 648
rect 130 651 136 652
rect 130 647 131 651
rect 135 647 136 651
rect 130 646 136 647
rect 306 651 312 652
rect 306 647 307 651
rect 311 647 312 651
rect 306 646 312 647
rect 158 636 164 637
rect 110 635 116 636
rect 110 631 111 635
rect 115 631 116 635
rect 158 632 159 636
rect 163 632 164 636
rect 158 631 164 632
rect 334 636 340 637
rect 334 632 335 636
rect 339 632 340 636
rect 334 631 340 632
rect 110 630 116 631
rect 112 607 114 630
rect 160 607 162 631
rect 336 607 338 631
rect 111 606 115 607
rect 111 601 115 602
rect 159 606 163 607
rect 159 601 163 602
rect 335 606 339 607
rect 335 601 339 602
rect 375 606 379 607
rect 375 601 379 602
rect 112 578 114 601
rect 110 577 116 578
rect 160 577 162 601
rect 376 577 378 601
rect 110 573 111 577
rect 115 573 116 577
rect 110 572 116 573
rect 158 576 164 577
rect 158 572 159 576
rect 163 572 164 576
rect 158 571 164 572
rect 374 576 380 577
rect 374 572 375 576
rect 379 572 380 576
rect 374 571 380 572
rect 130 561 136 562
rect 110 560 116 561
rect 110 556 111 560
rect 115 556 116 560
rect 130 557 131 561
rect 135 557 136 561
rect 130 556 136 557
rect 346 561 352 562
rect 346 557 347 561
rect 351 557 352 561
rect 346 556 352 557
rect 110 555 116 556
rect 112 495 114 555
rect 132 495 134 556
rect 226 519 232 520
rect 226 515 227 519
rect 231 515 232 519
rect 226 514 232 515
rect 111 494 115 495
rect 111 489 115 490
rect 131 494 135 495
rect 131 489 135 490
rect 112 429 114 489
rect 110 428 116 429
rect 132 428 134 489
rect 228 436 230 514
rect 348 495 350 556
rect 476 552 478 690
rect 500 652 502 713
rect 684 652 686 713
rect 810 695 816 696
rect 810 691 811 695
rect 815 691 816 695
rect 810 690 816 691
rect 812 660 814 690
rect 810 659 816 660
rect 810 655 811 659
rect 815 655 816 659
rect 810 654 816 655
rect 860 652 862 713
rect 1020 696 1022 770
rect 1136 744 1138 770
rect 1134 743 1140 744
rect 1134 739 1135 743
rect 1139 739 1140 743
rect 1134 738 1140 739
rect 1212 719 1214 780
rect 1228 744 1230 894
rect 1260 892 1262 953
rect 1444 892 1446 953
rect 1606 935 1612 936
rect 1606 931 1607 935
rect 1611 931 1612 935
rect 1606 930 1612 931
rect 1608 900 1610 930
rect 1606 899 1612 900
rect 1606 895 1607 899
rect 1611 895 1612 899
rect 1606 894 1612 895
rect 1628 892 1630 953
rect 1788 892 1790 953
rect 1936 893 1938 953
rect 1976 935 1978 986
rect 1975 934 1979 935
rect 1975 929 1979 930
rect 2047 934 2051 935
rect 2047 929 2051 930
rect 2351 934 2355 935
rect 2351 929 2355 930
rect 2647 934 2651 935
rect 2647 929 2651 930
rect 2927 934 2931 935
rect 2927 929 2931 930
rect 1976 906 1978 929
rect 1974 905 1980 906
rect 2048 905 2050 929
rect 2352 905 2354 929
rect 2648 905 2650 929
rect 2928 905 2930 929
rect 1974 901 1975 905
rect 1979 901 1980 905
rect 1974 900 1980 901
rect 2046 904 2052 905
rect 2046 900 2047 904
rect 2051 900 2052 904
rect 2046 899 2052 900
rect 2350 904 2356 905
rect 2350 900 2351 904
rect 2355 900 2356 904
rect 2350 899 2356 900
rect 2646 904 2652 905
rect 2646 900 2647 904
rect 2651 900 2652 904
rect 2646 899 2652 900
rect 2926 904 2932 905
rect 2926 900 2927 904
rect 2931 900 2932 904
rect 2926 899 2932 900
rect 1934 892 1940 893
rect 1258 891 1264 892
rect 1258 887 1259 891
rect 1263 887 1264 891
rect 1258 886 1264 887
rect 1442 891 1448 892
rect 1442 887 1443 891
rect 1447 887 1448 891
rect 1442 886 1448 887
rect 1626 891 1632 892
rect 1626 887 1627 891
rect 1631 887 1632 891
rect 1626 886 1632 887
rect 1786 891 1792 892
rect 1786 887 1787 891
rect 1791 887 1792 891
rect 1934 888 1935 892
rect 1939 888 1940 892
rect 2018 889 2024 890
rect 1934 887 1940 888
rect 1974 888 1980 889
rect 1786 886 1792 887
rect 1974 884 1975 888
rect 1979 884 1980 888
rect 2018 885 2019 889
rect 2023 885 2024 889
rect 2018 884 2024 885
rect 2322 889 2328 890
rect 2322 885 2323 889
rect 2327 885 2328 889
rect 2322 884 2328 885
rect 2618 889 2624 890
rect 2618 885 2619 889
rect 2623 885 2624 889
rect 2618 884 2624 885
rect 2898 889 2904 890
rect 2898 885 2899 889
rect 2903 885 2904 889
rect 2898 884 2904 885
rect 1974 883 1980 884
rect 1286 876 1292 877
rect 1286 872 1287 876
rect 1291 872 1292 876
rect 1286 871 1292 872
rect 1470 876 1476 877
rect 1470 872 1471 876
rect 1475 872 1476 876
rect 1470 871 1476 872
rect 1654 876 1660 877
rect 1654 872 1655 876
rect 1659 872 1660 876
rect 1654 871 1660 872
rect 1814 876 1820 877
rect 1814 872 1815 876
rect 1819 872 1820 876
rect 1814 871 1820 872
rect 1934 875 1940 876
rect 1934 871 1935 875
rect 1939 871 1940 875
rect 1288 831 1290 871
rect 1472 831 1474 871
rect 1656 831 1658 871
rect 1816 831 1818 871
rect 1934 870 1940 871
rect 1936 831 1938 870
rect 1239 830 1243 831
rect 1239 825 1243 826
rect 1287 830 1291 831
rect 1287 825 1291 826
rect 1471 830 1475 831
rect 1471 825 1475 826
rect 1535 830 1539 831
rect 1535 825 1539 826
rect 1655 830 1659 831
rect 1655 825 1659 826
rect 1815 830 1819 831
rect 1815 825 1819 826
rect 1935 830 1939 831
rect 1935 825 1939 826
rect 1240 801 1242 825
rect 1536 801 1538 825
rect 1816 801 1818 825
rect 1936 802 1938 825
rect 1976 823 1978 883
rect 2020 823 2022 884
rect 2166 879 2172 880
rect 2166 875 2167 879
rect 2171 875 2172 879
rect 2166 874 2172 875
rect 2168 848 2170 874
rect 2166 847 2172 848
rect 2166 843 2167 847
rect 2171 843 2172 847
rect 2166 842 2172 843
rect 2324 823 2326 884
rect 2410 847 2416 848
rect 2410 843 2411 847
rect 2415 843 2416 847
rect 2410 842 2416 843
rect 1975 822 1979 823
rect 1975 817 1979 818
rect 1995 822 1999 823
rect 1995 817 1999 818
rect 2019 822 2023 823
rect 2019 817 2023 818
rect 2251 822 2255 823
rect 2251 817 2255 818
rect 2323 822 2327 823
rect 2323 817 2327 818
rect 1934 801 1940 802
rect 1238 800 1244 801
rect 1238 796 1239 800
rect 1243 796 1244 800
rect 1238 795 1244 796
rect 1534 800 1540 801
rect 1534 796 1535 800
rect 1539 796 1540 800
rect 1534 795 1540 796
rect 1814 800 1820 801
rect 1814 796 1815 800
rect 1819 796 1820 800
rect 1934 797 1935 801
rect 1939 797 1940 801
rect 1934 796 1940 797
rect 1942 799 1948 800
rect 1814 795 1820 796
rect 1942 795 1943 799
rect 1947 795 1948 799
rect 1942 794 1948 795
rect 1506 785 1512 786
rect 1506 781 1507 785
rect 1511 781 1512 785
rect 1506 780 1512 781
rect 1786 785 1792 786
rect 1786 781 1787 785
rect 1791 781 1792 785
rect 1786 780 1792 781
rect 1934 784 1940 785
rect 1934 780 1935 784
rect 1939 780 1940 784
rect 1226 743 1232 744
rect 1226 739 1227 743
rect 1231 739 1232 743
rect 1226 738 1232 739
rect 1508 719 1510 780
rect 1788 719 1790 780
rect 1934 779 1940 780
rect 1802 775 1808 776
rect 1802 771 1803 775
rect 1807 771 1808 775
rect 1802 770 1808 771
rect 1804 744 1806 770
rect 1910 759 1916 760
rect 1910 755 1911 759
rect 1915 755 1916 759
rect 1910 754 1916 755
rect 1802 743 1808 744
rect 1802 739 1803 743
rect 1807 739 1808 743
rect 1802 738 1808 739
rect 1027 718 1031 719
rect 1027 713 1031 714
rect 1187 718 1191 719
rect 1187 713 1191 714
rect 1211 718 1215 719
rect 1211 713 1215 714
rect 1339 718 1343 719
rect 1339 713 1343 714
rect 1491 718 1495 719
rect 1491 713 1495 714
rect 1507 718 1511 719
rect 1507 713 1511 714
rect 1651 718 1655 719
rect 1651 713 1655 714
rect 1787 718 1791 719
rect 1787 713 1791 714
rect 1018 695 1024 696
rect 1018 691 1019 695
rect 1023 691 1024 695
rect 1018 690 1024 691
rect 986 659 992 660
rect 986 655 987 659
rect 991 655 992 659
rect 986 654 992 655
rect 498 651 504 652
rect 498 647 499 651
rect 503 647 504 651
rect 498 646 504 647
rect 682 651 688 652
rect 682 647 683 651
rect 687 647 688 651
rect 682 646 688 647
rect 858 651 864 652
rect 858 647 859 651
rect 863 647 864 651
rect 858 646 864 647
rect 526 636 532 637
rect 526 632 527 636
rect 531 632 532 636
rect 526 631 532 632
rect 710 636 716 637
rect 710 632 711 636
rect 715 632 716 636
rect 710 631 716 632
rect 886 636 892 637
rect 886 632 887 636
rect 891 632 892 636
rect 886 631 892 632
rect 528 607 530 631
rect 712 607 714 631
rect 888 607 890 631
rect 527 606 531 607
rect 527 601 531 602
rect 599 606 603 607
rect 599 601 603 602
rect 711 606 715 607
rect 711 601 715 602
rect 807 606 811 607
rect 807 601 811 602
rect 887 606 891 607
rect 887 601 891 602
rect 600 577 602 601
rect 808 577 810 601
rect 598 576 604 577
rect 598 572 599 576
rect 603 572 604 576
rect 598 571 604 572
rect 806 576 812 577
rect 806 572 807 576
rect 811 572 812 576
rect 806 571 812 572
rect 570 561 576 562
rect 570 557 571 561
rect 575 557 576 561
rect 570 556 576 557
rect 778 561 784 562
rect 778 557 779 561
rect 783 557 784 561
rect 778 556 784 557
rect 970 561 976 562
rect 970 557 971 561
rect 975 557 976 561
rect 970 556 976 557
rect 362 551 368 552
rect 362 547 363 551
rect 367 547 368 551
rect 362 546 368 547
rect 474 551 480 552
rect 474 547 475 551
rect 479 547 480 551
rect 474 546 480 547
rect 364 520 366 546
rect 362 519 368 520
rect 362 515 363 519
rect 367 515 368 519
rect 362 514 368 515
rect 572 495 574 556
rect 698 551 704 552
rect 698 547 699 551
rect 703 547 704 551
rect 698 546 704 547
rect 347 494 351 495
rect 347 489 351 490
rect 427 494 431 495
rect 427 489 431 490
rect 571 494 575 495
rect 571 489 575 490
rect 350 471 356 472
rect 350 467 351 471
rect 355 467 356 471
rect 350 466 356 467
rect 352 436 354 466
rect 226 435 232 436
rect 226 431 227 435
rect 231 431 232 435
rect 226 430 232 431
rect 350 435 356 436
rect 350 431 351 435
rect 355 431 356 435
rect 350 430 356 431
rect 428 428 430 489
rect 700 472 702 546
rect 780 495 782 556
rect 972 495 974 556
rect 988 520 990 654
rect 1028 652 1030 713
rect 1150 679 1156 680
rect 1150 675 1151 679
rect 1155 675 1156 679
rect 1150 674 1156 675
rect 1152 660 1154 674
rect 1150 659 1156 660
rect 1150 655 1151 659
rect 1155 655 1156 659
rect 1150 654 1156 655
rect 1188 652 1190 713
rect 1274 691 1280 692
rect 1274 687 1275 691
rect 1279 687 1280 691
rect 1274 686 1280 687
rect 1026 651 1032 652
rect 1026 647 1027 651
rect 1031 647 1032 651
rect 1026 646 1032 647
rect 1186 651 1192 652
rect 1186 647 1187 651
rect 1191 647 1192 651
rect 1186 646 1192 647
rect 1054 636 1060 637
rect 1054 632 1055 636
rect 1059 632 1060 636
rect 1054 631 1060 632
rect 1214 636 1220 637
rect 1214 632 1215 636
rect 1219 632 1220 636
rect 1214 631 1220 632
rect 1056 607 1058 631
rect 1216 607 1218 631
rect 999 606 1003 607
rect 999 601 1003 602
rect 1055 606 1059 607
rect 1055 601 1059 602
rect 1175 606 1179 607
rect 1175 601 1179 602
rect 1215 606 1219 607
rect 1215 601 1219 602
rect 1000 577 1002 601
rect 1176 577 1178 601
rect 998 576 1004 577
rect 998 572 999 576
rect 1003 572 1004 576
rect 998 571 1004 572
rect 1174 576 1180 577
rect 1174 572 1175 576
rect 1179 572 1180 576
rect 1174 571 1180 572
rect 1146 561 1152 562
rect 1146 557 1147 561
rect 1151 557 1152 561
rect 1146 556 1152 557
rect 986 519 992 520
rect 986 515 987 519
rect 991 515 992 519
rect 986 514 992 515
rect 1148 495 1150 556
rect 1276 552 1278 686
rect 1340 652 1342 713
rect 1492 652 1494 713
rect 1652 652 1654 713
rect 1788 652 1790 713
rect 1912 660 1914 754
rect 1936 719 1938 779
rect 1944 776 1946 794
rect 1942 775 1948 776
rect 1942 771 1943 775
rect 1947 771 1948 775
rect 1942 770 1948 771
rect 1976 757 1978 817
rect 1974 756 1980 757
rect 1996 756 1998 817
rect 2122 799 2128 800
rect 2122 795 2123 799
rect 2127 795 2128 799
rect 2122 794 2128 795
rect 2124 764 2126 794
rect 2122 763 2128 764
rect 2122 759 2123 763
rect 2127 759 2128 763
rect 2122 758 2128 759
rect 2252 756 2254 817
rect 2378 799 2384 800
rect 2378 795 2379 799
rect 2383 795 2384 799
rect 2378 794 2384 795
rect 2380 764 2382 794
rect 2412 764 2414 842
rect 2620 823 2622 884
rect 2746 879 2752 880
rect 2746 875 2747 879
rect 2751 875 2752 879
rect 2746 874 2752 875
rect 2830 879 2836 880
rect 2830 875 2831 879
rect 2835 875 2836 879
rect 2830 874 2836 875
rect 2523 822 2527 823
rect 2523 817 2527 818
rect 2619 822 2623 823
rect 2619 817 2623 818
rect 2378 763 2384 764
rect 2378 759 2379 763
rect 2383 759 2384 763
rect 2378 758 2384 759
rect 2410 763 2416 764
rect 2410 759 2411 763
rect 2415 759 2416 763
rect 2410 758 2416 759
rect 2524 756 2526 817
rect 2748 800 2750 874
rect 2832 848 2834 874
rect 2830 847 2836 848
rect 2830 843 2831 847
rect 2835 843 2836 847
rect 2830 842 2836 843
rect 2900 823 2902 884
rect 2988 848 2990 1010
rect 3092 1008 3094 1069
rect 3244 1008 3246 1069
rect 3370 1051 3376 1052
rect 3330 1047 3336 1048
rect 3330 1043 3331 1047
rect 3335 1043 3336 1047
rect 3370 1047 3371 1051
rect 3375 1047 3376 1051
rect 3370 1046 3376 1047
rect 3330 1042 3336 1043
rect 3090 1007 3096 1008
rect 3090 1003 3091 1007
rect 3095 1003 3096 1007
rect 3090 1002 3096 1003
rect 3242 1007 3248 1008
rect 3242 1003 3243 1007
rect 3247 1003 3248 1007
rect 3242 1002 3248 1003
rect 3118 992 3124 993
rect 3118 988 3119 992
rect 3123 988 3124 992
rect 3118 987 3124 988
rect 3270 992 3276 993
rect 3270 988 3271 992
rect 3275 988 3276 992
rect 3270 987 3276 988
rect 3120 935 3122 987
rect 3272 935 3274 987
rect 3119 934 3123 935
rect 3119 929 3123 930
rect 3207 934 3211 935
rect 3207 929 3211 930
rect 3271 934 3275 935
rect 3271 929 3275 930
rect 3208 905 3210 929
rect 3206 904 3212 905
rect 3206 900 3207 904
rect 3211 900 3212 904
rect 3206 899 3212 900
rect 3178 889 3184 890
rect 3178 885 3179 889
rect 3183 885 3184 889
rect 3178 884 3184 885
rect 2986 847 2992 848
rect 2986 843 2987 847
rect 2991 843 2992 847
rect 2986 842 2992 843
rect 3180 823 3182 884
rect 3332 880 3334 1042
rect 3372 1016 3374 1046
rect 3380 1016 3382 1118
rect 3428 1075 3430 1160
rect 3556 1156 3558 1290
rect 3596 1264 3598 1294
rect 3594 1263 3600 1264
rect 3594 1259 3595 1263
rect 3599 1259 3600 1263
rect 3594 1258 3600 1259
rect 3652 1256 3654 1317
rect 3738 1263 3744 1264
rect 3738 1259 3739 1263
rect 3743 1259 3744 1263
rect 3738 1258 3744 1259
rect 3650 1255 3656 1256
rect 3650 1251 3651 1255
rect 3655 1251 3656 1255
rect 3650 1250 3656 1251
rect 3678 1240 3684 1241
rect 3678 1236 3679 1240
rect 3683 1236 3684 1240
rect 3678 1235 3684 1236
rect 3680 1211 3682 1235
rect 3679 1210 3683 1211
rect 3679 1205 3683 1206
rect 3680 1181 3682 1205
rect 3678 1180 3684 1181
rect 3678 1176 3679 1180
rect 3683 1176 3684 1180
rect 3678 1175 3684 1176
rect 3650 1165 3656 1166
rect 3650 1161 3651 1165
rect 3655 1161 3656 1165
rect 3650 1160 3656 1161
rect 3442 1155 3448 1156
rect 3442 1151 3443 1155
rect 3447 1151 3448 1155
rect 3442 1150 3448 1151
rect 3554 1155 3560 1156
rect 3554 1151 3555 1155
rect 3559 1151 3560 1155
rect 3554 1150 3560 1151
rect 3444 1124 3446 1150
rect 3442 1123 3448 1124
rect 3442 1119 3443 1123
rect 3447 1119 3448 1123
rect 3442 1118 3448 1119
rect 3652 1075 3654 1160
rect 3740 1124 3742 1258
rect 3800 1257 3802 1317
rect 3838 1315 3839 1319
rect 3843 1315 3844 1319
rect 4838 1316 4839 1320
rect 4843 1316 4844 1320
rect 4838 1315 4844 1316
rect 3838 1314 3844 1315
rect 3840 1287 3842 1314
rect 4840 1287 4842 1315
rect 3839 1286 3843 1287
rect 3839 1281 3843 1282
rect 4735 1286 4739 1287
rect 4735 1281 4739 1282
rect 4839 1286 4843 1287
rect 4839 1281 4843 1282
rect 4879 1286 4883 1287
rect 4879 1281 4883 1282
rect 3840 1258 3842 1281
rect 3838 1257 3844 1258
rect 4736 1257 4738 1281
rect 4880 1257 4882 1281
rect 3798 1256 3804 1257
rect 3798 1252 3799 1256
rect 3803 1252 3804 1256
rect 3838 1253 3839 1257
rect 3843 1253 3844 1257
rect 3838 1252 3844 1253
rect 4734 1256 4740 1257
rect 4734 1252 4735 1256
rect 4739 1252 4740 1256
rect 3798 1251 3804 1252
rect 4734 1251 4740 1252
rect 4878 1256 4884 1257
rect 4878 1252 4879 1256
rect 4883 1252 4884 1256
rect 4878 1251 4884 1252
rect 4706 1241 4712 1242
rect 3838 1240 3844 1241
rect 3798 1239 3804 1240
rect 3798 1235 3799 1239
rect 3803 1235 3804 1239
rect 3838 1236 3839 1240
rect 3843 1236 3844 1240
rect 4706 1237 4707 1241
rect 4711 1237 4712 1241
rect 4706 1236 4712 1237
rect 4850 1241 4856 1242
rect 4850 1237 4851 1241
rect 4855 1237 4856 1241
rect 4850 1236 4856 1237
rect 3838 1235 3844 1236
rect 3798 1234 3804 1235
rect 3800 1211 3802 1234
rect 3799 1210 3803 1211
rect 3799 1205 3803 1206
rect 3800 1182 3802 1205
rect 3798 1181 3804 1182
rect 3798 1177 3799 1181
rect 3803 1177 3804 1181
rect 3798 1176 3804 1177
rect 3840 1167 3842 1235
rect 4708 1167 4710 1236
rect 4794 1223 4800 1224
rect 4794 1219 4795 1223
rect 4799 1219 4800 1223
rect 4794 1218 4800 1219
rect 4796 1200 4798 1218
rect 4794 1199 4800 1200
rect 4794 1195 4795 1199
rect 4799 1195 4800 1199
rect 4794 1194 4800 1195
rect 4852 1167 4854 1236
rect 4858 1231 4864 1232
rect 4858 1227 4859 1231
rect 4863 1227 4864 1231
rect 4858 1226 4864 1227
rect 4860 1187 4862 1226
rect 4936 1200 4938 1338
rect 4948 1336 4950 1397
rect 5084 1336 5086 1397
rect 5220 1336 5222 1397
rect 5306 1375 5312 1376
rect 5306 1371 5307 1375
rect 5311 1371 5312 1375
rect 5306 1370 5312 1371
rect 4946 1335 4952 1336
rect 4946 1331 4947 1335
rect 4951 1331 4952 1335
rect 4946 1330 4952 1331
rect 5082 1335 5088 1336
rect 5082 1331 5083 1335
rect 5087 1331 5088 1335
rect 5082 1330 5088 1331
rect 5218 1335 5224 1336
rect 5218 1331 5219 1335
rect 5223 1331 5224 1335
rect 5218 1330 5224 1331
rect 4974 1320 4980 1321
rect 4974 1316 4975 1320
rect 4979 1316 4980 1320
rect 4974 1315 4980 1316
rect 5110 1320 5116 1321
rect 5110 1316 5111 1320
rect 5115 1316 5116 1320
rect 5110 1315 5116 1316
rect 5246 1320 5252 1321
rect 5246 1316 5247 1320
rect 5251 1316 5252 1320
rect 5246 1315 5252 1316
rect 4976 1287 4978 1315
rect 5112 1287 5114 1315
rect 5248 1287 5250 1315
rect 4975 1286 4979 1287
rect 4975 1281 4979 1282
rect 5031 1286 5035 1287
rect 5031 1281 5035 1282
rect 5111 1286 5115 1287
rect 5111 1281 5115 1282
rect 5191 1286 5195 1287
rect 5191 1281 5195 1282
rect 5247 1286 5251 1287
rect 5247 1281 5251 1282
rect 5032 1257 5034 1281
rect 5192 1257 5194 1281
rect 5030 1256 5036 1257
rect 5030 1252 5031 1256
rect 5035 1252 5036 1256
rect 5030 1251 5036 1252
rect 5190 1256 5196 1257
rect 5190 1252 5191 1256
rect 5195 1252 5196 1256
rect 5190 1251 5196 1252
rect 5002 1241 5008 1242
rect 5002 1237 5003 1241
rect 5007 1237 5008 1241
rect 5002 1236 5008 1237
rect 5162 1241 5168 1242
rect 5162 1237 5163 1241
rect 5167 1237 5168 1241
rect 5162 1236 5168 1237
rect 4934 1199 4940 1200
rect 4934 1195 4935 1199
rect 4939 1195 4940 1199
rect 4934 1194 4940 1195
rect 4860 1185 4870 1187
rect 3839 1166 3843 1167
rect 3798 1164 3804 1165
rect 3798 1160 3799 1164
rect 3803 1160 3804 1164
rect 3839 1161 3843 1162
rect 3859 1166 3863 1167
rect 3859 1161 3863 1162
rect 4067 1166 4071 1167
rect 4067 1161 4071 1162
rect 4299 1166 4303 1167
rect 4299 1161 4303 1162
rect 4539 1166 4543 1167
rect 4539 1161 4543 1162
rect 4707 1166 4711 1167
rect 4707 1161 4711 1162
rect 4779 1166 4783 1167
rect 4779 1161 4783 1162
rect 4851 1166 4855 1167
rect 4851 1161 4855 1162
rect 3798 1159 3804 1160
rect 3738 1123 3744 1124
rect 3738 1119 3739 1123
rect 3743 1119 3744 1123
rect 3738 1118 3744 1119
rect 3800 1075 3802 1159
rect 3840 1101 3842 1161
rect 3838 1100 3844 1101
rect 3860 1100 3862 1161
rect 4034 1143 4040 1144
rect 4034 1139 4035 1143
rect 4039 1139 4040 1143
rect 4034 1138 4040 1139
rect 4036 1108 4038 1138
rect 4034 1107 4040 1108
rect 4034 1103 4035 1107
rect 4039 1103 4040 1107
rect 4034 1102 4040 1103
rect 4068 1100 4070 1161
rect 4130 1107 4136 1108
rect 4130 1103 4131 1107
rect 4135 1103 4136 1107
rect 4130 1102 4136 1103
rect 3838 1096 3839 1100
rect 3843 1096 3844 1100
rect 3838 1095 3844 1096
rect 3858 1099 3864 1100
rect 3858 1095 3859 1099
rect 3863 1095 3864 1099
rect 3858 1094 3864 1095
rect 4066 1099 4072 1100
rect 4066 1095 4067 1099
rect 4071 1095 4072 1099
rect 4066 1094 4072 1095
rect 3886 1084 3892 1085
rect 3838 1083 3844 1084
rect 3838 1079 3839 1083
rect 3843 1079 3844 1083
rect 3886 1080 3887 1084
rect 3891 1080 3892 1084
rect 3886 1079 3892 1080
rect 4094 1084 4100 1085
rect 4094 1080 4095 1084
rect 4099 1080 4100 1084
rect 4094 1079 4100 1080
rect 3838 1078 3844 1079
rect 3395 1074 3399 1075
rect 3395 1069 3399 1070
rect 3427 1074 3431 1075
rect 3427 1069 3431 1070
rect 3651 1074 3655 1075
rect 3651 1069 3655 1070
rect 3799 1074 3803 1075
rect 3799 1069 3803 1070
rect 3370 1015 3376 1016
rect 3370 1011 3371 1015
rect 3375 1011 3376 1015
rect 3370 1010 3376 1011
rect 3378 1015 3384 1016
rect 3378 1011 3379 1015
rect 3383 1011 3384 1015
rect 3378 1010 3384 1011
rect 3396 1008 3398 1069
rect 3800 1009 3802 1069
rect 3840 1055 3842 1078
rect 3888 1055 3890 1079
rect 4096 1055 4098 1079
rect 3839 1054 3843 1055
rect 3839 1049 3843 1050
rect 3887 1054 3891 1055
rect 3887 1049 3891 1050
rect 4071 1054 4075 1055
rect 4071 1049 4075 1050
rect 4095 1054 4099 1055
rect 4095 1049 4099 1050
rect 3840 1026 3842 1049
rect 3838 1025 3844 1026
rect 3888 1025 3890 1049
rect 4072 1025 4074 1049
rect 3838 1021 3839 1025
rect 3843 1021 3844 1025
rect 3838 1020 3844 1021
rect 3886 1024 3892 1025
rect 3886 1020 3887 1024
rect 3891 1020 3892 1024
rect 3886 1019 3892 1020
rect 4070 1024 4076 1025
rect 4070 1020 4071 1024
rect 4075 1020 4076 1024
rect 4070 1019 4076 1020
rect 3858 1009 3864 1010
rect 3798 1008 3804 1009
rect 3394 1007 3400 1008
rect 3394 1003 3395 1007
rect 3399 1003 3400 1007
rect 3798 1004 3799 1008
rect 3803 1004 3804 1008
rect 3798 1003 3804 1004
rect 3838 1008 3844 1009
rect 3838 1004 3839 1008
rect 3843 1004 3844 1008
rect 3858 1005 3859 1009
rect 3863 1005 3864 1009
rect 3858 1004 3864 1005
rect 4042 1009 4048 1010
rect 4042 1005 4043 1009
rect 4047 1005 4048 1009
rect 4042 1004 4048 1005
rect 3838 1003 3844 1004
rect 3394 1002 3400 1003
rect 3422 992 3428 993
rect 3422 988 3423 992
rect 3427 988 3428 992
rect 3422 987 3428 988
rect 3798 991 3804 992
rect 3798 987 3799 991
rect 3803 987 3804 991
rect 3424 935 3426 987
rect 3798 986 3804 987
rect 3800 935 3802 986
rect 3840 943 3842 1003
rect 3860 943 3862 1004
rect 3962 999 3968 1000
rect 3962 995 3963 999
rect 3967 995 3968 999
rect 3962 994 3968 995
rect 4018 999 4024 1000
rect 4018 995 4019 999
rect 4023 995 4024 999
rect 4018 994 4024 995
rect 3839 942 3843 943
rect 3839 937 3843 938
rect 3859 942 3863 943
rect 3859 937 3863 938
rect 3423 934 3427 935
rect 3423 929 3427 930
rect 3495 934 3499 935
rect 3495 929 3499 930
rect 3799 934 3803 935
rect 3799 929 3803 930
rect 3496 905 3498 929
rect 3800 906 3802 929
rect 3798 905 3804 906
rect 3494 904 3500 905
rect 3494 900 3495 904
rect 3499 900 3500 904
rect 3798 901 3799 905
rect 3803 901 3804 905
rect 3798 900 3804 901
rect 3494 899 3500 900
rect 3466 889 3472 890
rect 3466 885 3467 889
rect 3471 885 3472 889
rect 3466 884 3472 885
rect 3798 888 3804 889
rect 3798 884 3799 888
rect 3803 884 3804 888
rect 3330 879 3336 880
rect 3330 875 3331 879
rect 3335 875 3336 879
rect 3330 874 3336 875
rect 3378 879 3384 880
rect 3378 875 3379 879
rect 3383 875 3384 879
rect 3378 874 3384 875
rect 3380 848 3382 874
rect 3378 847 3384 848
rect 3378 843 3379 847
rect 3383 843 3384 847
rect 3378 842 3384 843
rect 3468 823 3470 884
rect 3798 883 3804 884
rect 3554 847 3560 848
rect 3554 843 3555 847
rect 3559 843 3560 847
rect 3554 842 3560 843
rect 2771 822 2775 823
rect 2771 817 2775 818
rect 2899 822 2903 823
rect 2899 817 2903 818
rect 3003 822 3007 823
rect 3003 817 3007 818
rect 3179 822 3183 823
rect 3179 817 3183 818
rect 3227 822 3231 823
rect 3227 817 3231 818
rect 3451 822 3455 823
rect 3451 817 3455 818
rect 3467 822 3471 823
rect 3467 817 3471 818
rect 2746 799 2752 800
rect 2746 795 2747 799
rect 2751 795 2752 799
rect 2746 794 2752 795
rect 2772 756 2774 817
rect 2898 799 2904 800
rect 2898 795 2899 799
rect 2903 795 2904 799
rect 2898 794 2904 795
rect 2900 764 2902 794
rect 2898 763 2904 764
rect 2898 759 2899 763
rect 2903 759 2904 763
rect 2898 758 2904 759
rect 3004 756 3006 817
rect 3228 756 3230 817
rect 3354 799 3360 800
rect 3314 795 3320 796
rect 3314 791 3315 795
rect 3319 791 3320 795
rect 3354 795 3355 799
rect 3359 795 3360 799
rect 3354 794 3360 795
rect 3314 790 3320 791
rect 3316 772 3318 790
rect 3314 771 3320 772
rect 3314 767 3315 771
rect 3319 767 3320 771
rect 3314 766 3320 767
rect 3356 764 3358 794
rect 3298 763 3304 764
rect 3298 759 3299 763
rect 3303 759 3304 763
rect 3298 758 3304 759
rect 3354 763 3360 764
rect 3354 759 3355 763
rect 3359 759 3360 763
rect 3354 758 3360 759
rect 1974 752 1975 756
rect 1979 752 1980 756
rect 1974 751 1980 752
rect 1994 755 2000 756
rect 1994 751 1995 755
rect 1999 751 2000 755
rect 1994 750 2000 751
rect 2250 755 2256 756
rect 2250 751 2251 755
rect 2255 751 2256 755
rect 2250 750 2256 751
rect 2522 755 2528 756
rect 2522 751 2523 755
rect 2527 751 2528 755
rect 2522 750 2528 751
rect 2770 755 2776 756
rect 2770 751 2771 755
rect 2775 751 2776 755
rect 2770 750 2776 751
rect 3002 755 3008 756
rect 3002 751 3003 755
rect 3007 751 3008 755
rect 3002 750 3008 751
rect 3226 755 3232 756
rect 3226 751 3227 755
rect 3231 751 3232 755
rect 3226 750 3232 751
rect 2022 740 2028 741
rect 1974 739 1980 740
rect 1974 735 1975 739
rect 1979 735 1980 739
rect 2022 736 2023 740
rect 2027 736 2028 740
rect 2022 735 2028 736
rect 2278 740 2284 741
rect 2278 736 2279 740
rect 2283 736 2284 740
rect 2278 735 2284 736
rect 2550 740 2556 741
rect 2550 736 2551 740
rect 2555 736 2556 740
rect 2550 735 2556 736
rect 2798 740 2804 741
rect 2798 736 2799 740
rect 2803 736 2804 740
rect 2798 735 2804 736
rect 3030 740 3036 741
rect 3030 736 3031 740
rect 3035 736 3036 740
rect 3030 735 3036 736
rect 3254 740 3260 741
rect 3254 736 3255 740
rect 3259 736 3260 740
rect 3254 735 3260 736
rect 1974 734 1980 735
rect 1935 718 1939 719
rect 1935 713 1939 714
rect 1910 659 1916 660
rect 1910 655 1911 659
rect 1915 655 1916 659
rect 1910 654 1916 655
rect 1936 653 1938 713
rect 1934 652 1940 653
rect 1338 651 1344 652
rect 1338 647 1339 651
rect 1343 647 1344 651
rect 1338 646 1344 647
rect 1490 651 1496 652
rect 1490 647 1491 651
rect 1495 647 1496 651
rect 1490 646 1496 647
rect 1650 651 1656 652
rect 1650 647 1651 651
rect 1655 647 1656 651
rect 1650 646 1656 647
rect 1786 651 1792 652
rect 1786 647 1787 651
rect 1791 647 1792 651
rect 1934 648 1935 652
rect 1939 648 1940 652
rect 1934 647 1940 648
rect 1786 646 1792 647
rect 1366 636 1372 637
rect 1366 632 1367 636
rect 1371 632 1372 636
rect 1366 631 1372 632
rect 1518 636 1524 637
rect 1518 632 1519 636
rect 1523 632 1524 636
rect 1518 631 1524 632
rect 1678 636 1684 637
rect 1678 632 1679 636
rect 1683 632 1684 636
rect 1678 631 1684 632
rect 1814 636 1820 637
rect 1814 632 1815 636
rect 1819 632 1820 636
rect 1814 631 1820 632
rect 1934 635 1940 636
rect 1934 631 1935 635
rect 1939 631 1940 635
rect 1368 607 1370 631
rect 1520 607 1522 631
rect 1680 607 1682 631
rect 1816 607 1818 631
rect 1934 630 1940 631
rect 1936 607 1938 630
rect 1343 606 1347 607
rect 1343 601 1347 602
rect 1367 606 1371 607
rect 1367 601 1371 602
rect 1511 606 1515 607
rect 1511 601 1515 602
rect 1519 606 1523 607
rect 1519 601 1523 602
rect 1671 606 1675 607
rect 1671 601 1675 602
rect 1679 606 1683 607
rect 1679 601 1683 602
rect 1815 606 1819 607
rect 1815 601 1819 602
rect 1935 606 1939 607
rect 1935 601 1939 602
rect 1344 577 1346 601
rect 1512 577 1514 601
rect 1672 577 1674 601
rect 1816 577 1818 601
rect 1936 578 1938 601
rect 1976 579 1978 734
rect 2024 579 2026 735
rect 2280 579 2282 735
rect 2552 579 2554 735
rect 2800 579 2802 735
rect 3032 579 3034 735
rect 3256 579 3258 735
rect 1975 578 1979 579
rect 1934 577 1940 578
rect 1342 576 1348 577
rect 1342 572 1343 576
rect 1347 572 1348 576
rect 1342 571 1348 572
rect 1510 576 1516 577
rect 1510 572 1511 576
rect 1515 572 1516 576
rect 1510 571 1516 572
rect 1670 576 1676 577
rect 1670 572 1671 576
rect 1675 572 1676 576
rect 1670 571 1676 572
rect 1814 576 1820 577
rect 1814 572 1815 576
rect 1819 572 1820 576
rect 1934 573 1935 577
rect 1939 573 1940 577
rect 1975 573 1979 574
rect 2023 578 2027 579
rect 2023 573 2027 574
rect 2279 578 2283 579
rect 2279 573 2283 574
rect 2551 578 2555 579
rect 2551 573 2555 574
rect 2799 578 2803 579
rect 2799 573 2803 574
rect 3031 578 3035 579
rect 3031 573 3035 574
rect 3255 578 3259 579
rect 3255 573 3259 574
rect 1934 572 1940 573
rect 1814 571 1820 572
rect 1314 561 1320 562
rect 1314 557 1315 561
rect 1319 557 1320 561
rect 1314 556 1320 557
rect 1482 561 1488 562
rect 1482 557 1483 561
rect 1487 557 1488 561
rect 1482 556 1488 557
rect 1642 561 1648 562
rect 1642 557 1643 561
rect 1647 557 1648 561
rect 1642 556 1648 557
rect 1786 561 1792 562
rect 1786 557 1787 561
rect 1791 557 1792 561
rect 1786 556 1792 557
rect 1934 560 1940 561
rect 1934 556 1935 560
rect 1939 556 1940 560
rect 1274 551 1280 552
rect 1274 547 1275 551
rect 1279 547 1280 551
rect 1274 546 1280 547
rect 1302 551 1308 552
rect 1302 547 1303 551
rect 1307 547 1308 551
rect 1302 546 1308 547
rect 1304 520 1306 546
rect 1302 519 1308 520
rect 1302 515 1303 519
rect 1307 515 1308 519
rect 1302 514 1308 515
rect 1316 495 1318 556
rect 1484 495 1486 556
rect 1490 551 1496 552
rect 1490 547 1491 551
rect 1495 547 1496 551
rect 1490 546 1496 547
rect 1492 520 1494 546
rect 1490 519 1496 520
rect 1490 515 1491 519
rect 1495 515 1496 519
rect 1490 514 1496 515
rect 1644 495 1646 556
rect 1778 551 1784 552
rect 1778 547 1779 551
rect 1783 547 1784 551
rect 1778 546 1784 547
rect 1780 520 1782 546
rect 1778 519 1784 520
rect 1778 515 1779 519
rect 1783 515 1784 519
rect 1778 514 1784 515
rect 1788 495 1790 556
rect 1934 555 1940 556
rect 1882 519 1888 520
rect 1882 515 1883 519
rect 1887 515 1888 519
rect 1882 514 1888 515
rect 763 494 767 495
rect 763 489 767 490
rect 779 494 783 495
rect 779 489 783 490
rect 971 494 975 495
rect 971 489 975 490
rect 1107 494 1111 495
rect 1107 489 1111 490
rect 1147 494 1151 495
rect 1147 489 1151 490
rect 1315 494 1319 495
rect 1315 489 1319 490
rect 1459 494 1463 495
rect 1459 489 1463 490
rect 1483 494 1487 495
rect 1483 489 1487 490
rect 1643 494 1647 495
rect 1643 489 1647 490
rect 1787 494 1791 495
rect 1787 489 1791 490
rect 558 471 564 472
rect 558 467 559 471
rect 563 467 564 471
rect 558 466 564 467
rect 698 471 704 472
rect 698 467 699 471
rect 703 467 704 471
rect 698 466 704 467
rect 110 424 111 428
rect 115 424 116 428
rect 110 423 116 424
rect 130 427 136 428
rect 130 423 131 427
rect 135 423 136 427
rect 130 422 136 423
rect 426 427 432 428
rect 426 423 427 427
rect 431 423 432 427
rect 426 422 432 423
rect 158 412 164 413
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 158 408 159 412
rect 163 408 164 412
rect 158 407 164 408
rect 454 412 460 413
rect 454 408 455 412
rect 459 408 460 412
rect 454 407 460 408
rect 110 406 116 407
rect 112 367 114 406
rect 160 367 162 407
rect 456 367 458 407
rect 111 366 115 367
rect 111 361 115 362
rect 159 366 163 367
rect 159 361 163 362
rect 239 366 243 367
rect 239 361 243 362
rect 391 366 395 367
rect 391 361 395 362
rect 455 366 459 367
rect 455 361 459 362
rect 551 366 555 367
rect 551 361 555 362
rect 112 338 114 361
rect 110 337 116 338
rect 240 337 242 361
rect 392 337 394 361
rect 552 337 554 361
rect 110 333 111 337
rect 115 333 116 337
rect 110 332 116 333
rect 238 336 244 337
rect 238 332 239 336
rect 243 332 244 336
rect 238 331 244 332
rect 390 336 396 337
rect 390 332 391 336
rect 395 332 396 336
rect 390 331 396 332
rect 550 336 556 337
rect 550 332 551 336
rect 555 332 556 336
rect 550 331 556 332
rect 210 321 216 322
rect 110 320 116 321
rect 110 316 111 320
rect 115 316 116 320
rect 210 317 211 321
rect 215 317 216 321
rect 210 316 216 317
rect 362 321 368 322
rect 362 317 363 321
rect 367 317 368 321
rect 362 316 368 317
rect 522 321 528 322
rect 522 317 523 321
rect 527 317 528 321
rect 522 316 528 317
rect 110 315 116 316
rect 112 223 114 315
rect 212 223 214 316
rect 270 279 276 280
rect 270 275 271 279
rect 275 275 276 279
rect 270 274 276 275
rect 111 222 115 223
rect 111 217 115 218
rect 147 222 151 223
rect 147 217 151 218
rect 211 222 215 223
rect 211 217 215 218
rect 112 157 114 217
rect 110 156 116 157
rect 148 156 150 217
rect 272 164 274 274
rect 364 223 366 316
rect 378 311 384 312
rect 378 307 379 311
rect 383 307 384 311
rect 378 306 384 307
rect 380 280 382 306
rect 378 279 384 280
rect 378 275 379 279
rect 383 275 384 279
rect 378 274 384 275
rect 524 223 526 316
rect 560 312 562 466
rect 764 428 766 489
rect 890 471 896 472
rect 890 467 891 471
rect 895 467 896 471
rect 890 466 896 467
rect 892 436 894 466
rect 890 435 896 436
rect 890 431 891 435
rect 895 431 896 435
rect 890 430 896 431
rect 1108 428 1110 489
rect 1234 471 1240 472
rect 1234 467 1235 471
rect 1239 467 1240 471
rect 1234 466 1240 467
rect 1236 436 1238 466
rect 1234 435 1240 436
rect 1234 431 1235 435
rect 1239 431 1240 435
rect 1234 430 1240 431
rect 1460 428 1462 489
rect 1518 435 1524 436
rect 1518 431 1519 435
rect 1523 431 1524 435
rect 1518 430 1524 431
rect 762 427 768 428
rect 762 423 763 427
rect 767 423 768 427
rect 762 422 768 423
rect 1106 427 1112 428
rect 1106 423 1107 427
rect 1111 423 1112 427
rect 1106 422 1112 423
rect 1458 427 1464 428
rect 1458 423 1459 427
rect 1463 423 1464 427
rect 1458 422 1464 423
rect 790 412 796 413
rect 790 408 791 412
rect 795 408 796 412
rect 790 407 796 408
rect 1134 412 1140 413
rect 1134 408 1135 412
rect 1139 408 1140 412
rect 1134 407 1140 408
rect 1486 412 1492 413
rect 1486 408 1487 412
rect 1491 408 1492 412
rect 1486 407 1492 408
rect 792 367 794 407
rect 1136 367 1138 407
rect 1488 367 1490 407
rect 711 366 715 367
rect 711 361 715 362
rect 791 366 795 367
rect 791 361 795 362
rect 871 366 875 367
rect 871 361 875 362
rect 1031 366 1035 367
rect 1031 361 1035 362
rect 1135 366 1139 367
rect 1135 361 1139 362
rect 1487 366 1491 367
rect 1487 361 1491 362
rect 712 337 714 361
rect 872 337 874 361
rect 1032 337 1034 361
rect 710 336 716 337
rect 710 332 711 336
rect 715 332 716 336
rect 710 331 716 332
rect 870 336 876 337
rect 870 332 871 336
rect 875 332 876 336
rect 870 331 876 332
rect 1030 336 1036 337
rect 1030 332 1031 336
rect 1035 332 1036 336
rect 1030 331 1036 332
rect 682 321 688 322
rect 682 317 683 321
rect 687 317 688 321
rect 682 316 688 317
rect 842 321 848 322
rect 842 317 843 321
rect 847 317 848 321
rect 842 316 848 317
rect 1002 321 1008 322
rect 1002 317 1003 321
rect 1007 317 1008 321
rect 1002 316 1008 317
rect 538 311 544 312
rect 538 307 539 311
rect 543 307 544 311
rect 538 306 544 307
rect 558 311 564 312
rect 558 307 559 311
rect 563 307 564 311
rect 558 306 564 307
rect 540 280 542 306
rect 538 279 544 280
rect 538 275 539 279
rect 543 275 544 279
rect 538 274 544 275
rect 684 223 686 316
rect 810 311 816 312
rect 810 307 811 311
rect 815 307 816 311
rect 810 306 816 307
rect 283 222 287 223
rect 283 217 287 218
rect 363 222 367 223
rect 363 217 367 218
rect 419 222 423 223
rect 419 217 423 218
rect 523 222 527 223
rect 523 217 527 218
rect 555 222 559 223
rect 555 217 559 218
rect 683 222 687 223
rect 683 217 687 218
rect 691 222 695 223
rect 691 217 695 218
rect 270 163 276 164
rect 270 159 271 163
rect 275 159 276 163
rect 270 158 276 159
rect 284 156 286 217
rect 420 156 422 217
rect 556 156 558 217
rect 692 156 694 217
rect 812 200 814 306
rect 844 223 846 316
rect 1004 223 1006 316
rect 1520 280 1522 430
rect 1788 428 1790 489
rect 1884 436 1886 514
rect 1936 495 1938 555
rect 1976 550 1978 573
rect 1974 549 1980 550
rect 1974 545 1975 549
rect 1979 545 1980 549
rect 1974 544 1980 545
rect 3282 533 3288 534
rect 1974 532 1980 533
rect 1974 528 1975 532
rect 1979 528 1980 532
rect 3282 529 3283 533
rect 3287 529 3288 533
rect 3282 528 3288 529
rect 1974 527 1980 528
rect 1935 494 1939 495
rect 1935 489 1939 490
rect 1882 435 1888 436
rect 1882 431 1883 435
rect 1887 431 1888 435
rect 1882 430 1888 431
rect 1936 429 1938 489
rect 1976 467 1978 527
rect 3284 467 3286 528
rect 3300 492 3302 758
rect 3452 756 3454 817
rect 3556 764 3558 842
rect 3800 823 3802 883
rect 3840 877 3842 937
rect 3964 920 3966 994
rect 4020 968 4022 994
rect 4018 967 4024 968
rect 4018 963 4019 967
rect 4023 963 4024 967
rect 4018 962 4024 963
rect 4044 943 4046 1004
rect 4132 968 4134 1102
rect 4300 1100 4302 1161
rect 4426 1143 4432 1144
rect 4386 1139 4392 1140
rect 4386 1135 4387 1139
rect 4391 1135 4392 1139
rect 4426 1139 4427 1143
rect 4431 1139 4432 1143
rect 4426 1138 4432 1139
rect 4386 1134 4392 1135
rect 4388 1116 4390 1134
rect 4386 1115 4392 1116
rect 4386 1111 4387 1115
rect 4391 1111 4392 1115
rect 4386 1110 4392 1111
rect 4428 1108 4430 1138
rect 4426 1107 4432 1108
rect 4426 1103 4427 1107
rect 4431 1103 4432 1107
rect 4426 1102 4432 1103
rect 4540 1100 4542 1161
rect 4746 1107 4752 1108
rect 4746 1103 4747 1107
rect 4751 1103 4752 1107
rect 4746 1102 4752 1103
rect 4298 1099 4304 1100
rect 4298 1095 4299 1099
rect 4303 1095 4304 1099
rect 4298 1094 4304 1095
rect 4538 1099 4544 1100
rect 4538 1095 4539 1099
rect 4543 1095 4544 1099
rect 4538 1094 4544 1095
rect 4326 1084 4332 1085
rect 4326 1080 4327 1084
rect 4331 1080 4332 1084
rect 4326 1079 4332 1080
rect 4566 1084 4572 1085
rect 4566 1080 4567 1084
rect 4571 1080 4572 1084
rect 4566 1079 4572 1080
rect 4328 1055 4330 1079
rect 4568 1055 4570 1079
rect 4279 1054 4283 1055
rect 4279 1049 4283 1050
rect 4327 1054 4331 1055
rect 4327 1049 4331 1050
rect 4511 1054 4515 1055
rect 4511 1049 4515 1050
rect 4567 1054 4571 1055
rect 4567 1049 4571 1050
rect 4280 1025 4282 1049
rect 4512 1025 4514 1049
rect 4278 1024 4284 1025
rect 4278 1020 4279 1024
rect 4283 1020 4284 1024
rect 4278 1019 4284 1020
rect 4510 1024 4516 1025
rect 4510 1020 4511 1024
rect 4515 1020 4516 1024
rect 4510 1019 4516 1020
rect 4250 1009 4256 1010
rect 4250 1005 4251 1009
rect 4255 1005 4256 1009
rect 4250 1004 4256 1005
rect 4482 1009 4488 1010
rect 4482 1005 4483 1009
rect 4487 1005 4488 1009
rect 4482 1004 4488 1005
rect 4730 1009 4736 1010
rect 4730 1005 4731 1009
rect 4735 1005 4736 1009
rect 4730 1004 4736 1005
rect 4130 967 4136 968
rect 4130 963 4131 967
rect 4135 963 4136 967
rect 4130 962 4136 963
rect 4252 943 4254 1004
rect 4338 991 4344 992
rect 4338 987 4339 991
rect 4343 987 4344 991
rect 4338 986 4344 987
rect 4340 968 4342 986
rect 4338 967 4344 968
rect 4338 963 4339 967
rect 4343 963 4344 967
rect 4338 962 4344 963
rect 4484 943 4486 1004
rect 4498 999 4504 1000
rect 4498 995 4499 999
rect 4503 995 4504 999
rect 4498 994 4504 995
rect 4610 999 4616 1000
rect 4610 995 4611 999
rect 4615 995 4616 999
rect 4610 994 4616 995
rect 4500 968 4502 994
rect 4498 967 4504 968
rect 4498 963 4499 967
rect 4503 963 4504 967
rect 4498 962 4504 963
rect 3971 942 3975 943
rect 3971 937 3975 938
rect 4043 942 4047 943
rect 4043 937 4047 938
rect 4179 942 4183 943
rect 4179 937 4183 938
rect 4251 942 4255 943
rect 4251 937 4255 938
rect 4403 942 4407 943
rect 4403 937 4407 938
rect 4483 942 4487 943
rect 4483 937 4487 938
rect 3962 919 3968 920
rect 3962 915 3963 919
rect 3967 915 3968 919
rect 3962 914 3968 915
rect 3838 876 3844 877
rect 3972 876 3974 937
rect 4180 876 4182 937
rect 4306 919 4312 920
rect 4266 915 4272 916
rect 4266 911 4267 915
rect 4271 911 4272 915
rect 4306 915 4307 919
rect 4311 915 4312 919
rect 4306 914 4312 915
rect 4266 910 4272 911
rect 4268 892 4270 910
rect 4266 891 4272 892
rect 4266 887 4267 891
rect 4271 887 4272 891
rect 4266 886 4272 887
rect 4308 884 4310 914
rect 4266 883 4272 884
rect 4266 879 4267 883
rect 4271 879 4272 883
rect 4266 878 4272 879
rect 4306 883 4312 884
rect 4306 879 4307 883
rect 4311 879 4312 883
rect 4306 878 4312 879
rect 3838 872 3839 876
rect 3843 872 3844 876
rect 3838 871 3844 872
rect 3970 875 3976 876
rect 3970 871 3971 875
rect 3975 871 3976 875
rect 3970 870 3976 871
rect 4178 875 4184 876
rect 4178 871 4179 875
rect 4183 871 4184 875
rect 4178 870 4184 871
rect 3998 860 4004 861
rect 3838 859 3844 860
rect 3838 855 3839 859
rect 3843 855 3844 859
rect 3998 856 3999 860
rect 4003 856 4004 860
rect 3998 855 4004 856
rect 4206 860 4212 861
rect 4206 856 4207 860
rect 4211 856 4212 860
rect 4206 855 4212 856
rect 3838 854 3844 855
rect 3840 831 3842 854
rect 4000 831 4002 855
rect 4208 831 4210 855
rect 3839 830 3843 831
rect 3839 825 3843 826
rect 3887 830 3891 831
rect 3887 825 3891 826
rect 3999 830 4003 831
rect 3999 825 4003 826
rect 4047 830 4051 831
rect 4047 825 4051 826
rect 4207 830 4211 831
rect 4207 825 4211 826
rect 3651 822 3655 823
rect 3651 817 3655 818
rect 3799 822 3803 823
rect 3799 817 3803 818
rect 3554 763 3560 764
rect 3554 759 3555 763
rect 3559 759 3560 763
rect 3554 758 3560 759
rect 3652 756 3654 817
rect 3800 757 3802 817
rect 3840 802 3842 825
rect 3838 801 3844 802
rect 3888 801 3890 825
rect 4048 801 4050 825
rect 3838 797 3839 801
rect 3843 797 3844 801
rect 3838 796 3844 797
rect 3886 800 3892 801
rect 3886 796 3887 800
rect 3891 796 3892 800
rect 3866 795 3872 796
rect 3886 795 3892 796
rect 4046 800 4052 801
rect 4046 796 4047 800
rect 4051 796 4052 800
rect 4046 795 4052 796
rect 3866 791 3867 795
rect 3871 791 3872 795
rect 3866 790 3872 791
rect 3858 785 3864 786
rect 3838 784 3844 785
rect 3838 780 3839 784
rect 3843 780 3844 784
rect 3858 781 3859 785
rect 3863 781 3864 785
rect 3858 780 3864 781
rect 3838 779 3844 780
rect 3798 756 3804 757
rect 3450 755 3456 756
rect 3450 751 3451 755
rect 3455 751 3456 755
rect 3450 750 3456 751
rect 3650 755 3656 756
rect 3650 751 3651 755
rect 3655 751 3656 755
rect 3798 752 3799 756
rect 3803 752 3804 756
rect 3798 751 3804 752
rect 3650 750 3656 751
rect 3478 740 3484 741
rect 3478 736 3479 740
rect 3483 736 3484 740
rect 3478 735 3484 736
rect 3678 740 3684 741
rect 3678 736 3679 740
rect 3683 736 3684 740
rect 3678 735 3684 736
rect 3798 739 3804 740
rect 3798 735 3799 739
rect 3803 735 3804 739
rect 3480 579 3482 735
rect 3680 579 3682 735
rect 3798 734 3804 735
rect 3800 579 3802 734
rect 3840 711 3842 779
rect 3860 711 3862 780
rect 3839 710 3843 711
rect 3839 705 3843 706
rect 3859 710 3863 711
rect 3859 705 3863 706
rect 3840 645 3842 705
rect 3838 644 3844 645
rect 3860 644 3862 705
rect 3868 652 3870 790
rect 4018 785 4024 786
rect 4018 781 4019 785
rect 4023 781 4024 785
rect 4018 780 4024 781
rect 4250 785 4256 786
rect 4250 781 4251 785
rect 4255 781 4256 785
rect 4250 780 4256 781
rect 3986 775 3992 776
rect 3986 771 3987 775
rect 3991 771 3992 775
rect 3986 770 3992 771
rect 3988 688 3990 770
rect 4020 711 4022 780
rect 4026 775 4032 776
rect 4026 771 4027 775
rect 4031 771 4032 775
rect 4026 770 4032 771
rect 4028 744 4030 770
rect 4026 743 4032 744
rect 4026 739 4027 743
rect 4031 739 4032 743
rect 4026 738 4032 739
rect 4252 711 4254 780
rect 4268 744 4270 878
rect 4404 876 4406 937
rect 4612 920 4614 994
rect 4732 943 4734 1004
rect 4748 968 4750 1102
rect 4780 1100 4782 1161
rect 4868 1140 4870 1185
rect 5004 1167 5006 1236
rect 5018 1231 5024 1232
rect 5018 1227 5019 1231
rect 5023 1227 5024 1231
rect 5018 1226 5024 1227
rect 5020 1200 5022 1226
rect 5018 1199 5024 1200
rect 5018 1195 5019 1199
rect 5023 1195 5024 1199
rect 5018 1194 5024 1195
rect 5164 1167 5166 1236
rect 5308 1232 5310 1370
rect 5356 1336 5358 1397
rect 5482 1379 5488 1380
rect 5482 1375 5483 1379
rect 5487 1375 5488 1379
rect 5482 1374 5488 1375
rect 5484 1344 5486 1374
rect 5482 1343 5488 1344
rect 5482 1339 5483 1343
rect 5487 1339 5488 1343
rect 5482 1338 5488 1339
rect 5492 1336 5494 1397
rect 5586 1343 5592 1344
rect 5586 1339 5587 1343
rect 5591 1339 5592 1343
rect 5586 1338 5592 1339
rect 5354 1335 5360 1336
rect 5354 1331 5355 1335
rect 5359 1331 5360 1335
rect 5354 1330 5360 1331
rect 5490 1335 5496 1336
rect 5490 1331 5491 1335
rect 5495 1331 5496 1335
rect 5490 1330 5496 1331
rect 5382 1320 5388 1321
rect 5382 1316 5383 1320
rect 5387 1316 5388 1320
rect 5382 1315 5388 1316
rect 5518 1320 5524 1321
rect 5518 1316 5519 1320
rect 5523 1316 5524 1320
rect 5518 1315 5524 1316
rect 5384 1287 5386 1315
rect 5520 1287 5522 1315
rect 5359 1286 5363 1287
rect 5359 1281 5363 1282
rect 5383 1286 5387 1287
rect 5383 1281 5387 1282
rect 5519 1286 5523 1287
rect 5519 1281 5523 1282
rect 5527 1286 5531 1287
rect 5527 1281 5531 1282
rect 5360 1257 5362 1281
rect 5528 1257 5530 1281
rect 5358 1256 5364 1257
rect 5358 1252 5359 1256
rect 5363 1252 5364 1256
rect 5358 1251 5364 1252
rect 5526 1256 5532 1257
rect 5526 1252 5527 1256
rect 5531 1252 5532 1256
rect 5526 1251 5532 1252
rect 5330 1241 5336 1242
rect 5330 1237 5331 1241
rect 5335 1237 5336 1241
rect 5330 1236 5336 1237
rect 5498 1241 5504 1242
rect 5498 1237 5499 1241
rect 5503 1237 5504 1241
rect 5498 1236 5504 1237
rect 5306 1231 5312 1232
rect 5306 1227 5307 1231
rect 5311 1227 5312 1231
rect 5306 1226 5312 1227
rect 5318 1231 5324 1232
rect 5318 1227 5319 1231
rect 5323 1227 5324 1231
rect 5318 1226 5324 1227
rect 5320 1200 5322 1226
rect 5318 1199 5324 1200
rect 5318 1195 5319 1199
rect 5323 1195 5324 1199
rect 5318 1194 5324 1195
rect 5332 1167 5334 1236
rect 5406 1199 5412 1200
rect 5406 1195 5407 1199
rect 5411 1195 5412 1199
rect 5406 1194 5412 1195
rect 5003 1166 5007 1167
rect 5003 1161 5007 1162
rect 5027 1166 5031 1167
rect 5027 1161 5031 1162
rect 5163 1166 5167 1167
rect 5163 1161 5167 1162
rect 5283 1166 5287 1167
rect 5283 1161 5287 1162
rect 5331 1166 5335 1167
rect 5331 1161 5335 1162
rect 4906 1143 4912 1144
rect 4866 1139 4872 1140
rect 4866 1135 4867 1139
rect 4871 1135 4872 1139
rect 4906 1139 4907 1143
rect 4911 1139 4912 1143
rect 4906 1138 4912 1139
rect 4866 1134 4872 1135
rect 4908 1108 4910 1138
rect 4906 1107 4912 1108
rect 4906 1103 4907 1107
rect 4911 1103 4912 1107
rect 4906 1102 4912 1103
rect 5028 1100 5030 1161
rect 5284 1100 5286 1161
rect 5370 1139 5376 1140
rect 5370 1135 5371 1139
rect 5375 1135 5376 1139
rect 5370 1134 5376 1135
rect 4778 1099 4784 1100
rect 4778 1095 4779 1099
rect 4783 1095 4784 1099
rect 4778 1094 4784 1095
rect 5026 1099 5032 1100
rect 5026 1095 5027 1099
rect 5031 1095 5032 1099
rect 5026 1094 5032 1095
rect 5282 1099 5288 1100
rect 5282 1095 5283 1099
rect 5287 1095 5288 1099
rect 5282 1094 5288 1095
rect 4806 1084 4812 1085
rect 4806 1080 4807 1084
rect 4811 1080 4812 1084
rect 4806 1079 4812 1080
rect 5054 1084 5060 1085
rect 5054 1080 5055 1084
rect 5059 1080 5060 1084
rect 5054 1079 5060 1080
rect 5310 1084 5316 1085
rect 5310 1080 5311 1084
rect 5315 1080 5316 1084
rect 5310 1079 5316 1080
rect 4808 1055 4810 1079
rect 5056 1055 5058 1079
rect 5312 1055 5314 1079
rect 4759 1054 4763 1055
rect 4759 1049 4763 1050
rect 4807 1054 4811 1055
rect 4807 1049 4811 1050
rect 5023 1054 5027 1055
rect 5023 1049 5027 1050
rect 5055 1054 5059 1055
rect 5055 1049 5059 1050
rect 5295 1054 5299 1055
rect 5295 1049 5299 1050
rect 5311 1054 5315 1055
rect 5311 1049 5315 1050
rect 4760 1025 4762 1049
rect 5024 1025 5026 1049
rect 5296 1025 5298 1049
rect 4758 1024 4764 1025
rect 4758 1020 4759 1024
rect 4763 1020 4764 1024
rect 4758 1019 4764 1020
rect 5022 1024 5028 1025
rect 5022 1020 5023 1024
rect 5027 1020 5028 1024
rect 5022 1019 5028 1020
rect 5294 1024 5300 1025
rect 5294 1020 5295 1024
rect 5299 1020 5300 1024
rect 5294 1019 5300 1020
rect 4994 1009 5000 1010
rect 4994 1005 4995 1009
rect 4999 1005 5000 1009
rect 4994 1004 5000 1005
rect 5266 1009 5272 1010
rect 5266 1005 5267 1009
rect 5271 1005 5272 1009
rect 5266 1004 5272 1005
rect 4746 967 4752 968
rect 4746 963 4747 967
rect 4751 963 4752 967
rect 4746 962 4752 963
rect 4996 943 4998 1004
rect 5010 999 5016 1000
rect 5010 995 5011 999
rect 5015 995 5016 999
rect 5010 994 5016 995
rect 5012 968 5014 994
rect 5010 967 5016 968
rect 5010 963 5011 967
rect 5015 963 5016 967
rect 5010 962 5016 963
rect 5268 943 5270 1004
rect 5372 1000 5374 1134
rect 5408 1108 5410 1194
rect 5500 1167 5502 1236
rect 5588 1200 5590 1338
rect 5664 1337 5666 1397
rect 5662 1336 5668 1337
rect 5662 1332 5663 1336
rect 5667 1332 5668 1336
rect 5662 1331 5668 1332
rect 5662 1319 5668 1320
rect 5662 1315 5663 1319
rect 5667 1315 5668 1319
rect 5662 1314 5668 1315
rect 5664 1287 5666 1314
rect 5663 1286 5667 1287
rect 5663 1281 5667 1282
rect 5664 1258 5666 1281
rect 5662 1257 5668 1258
rect 5662 1253 5663 1257
rect 5667 1253 5668 1257
rect 5662 1252 5668 1253
rect 5662 1240 5668 1241
rect 5662 1236 5663 1240
rect 5667 1236 5668 1240
rect 5662 1235 5668 1236
rect 5618 1231 5624 1232
rect 5618 1227 5619 1231
rect 5623 1227 5624 1231
rect 5618 1226 5624 1227
rect 5586 1199 5592 1200
rect 5586 1195 5587 1199
rect 5591 1195 5592 1199
rect 5586 1194 5592 1195
rect 5499 1166 5503 1167
rect 5499 1161 5503 1162
rect 5515 1166 5519 1167
rect 5515 1161 5519 1162
rect 5406 1107 5412 1108
rect 5406 1103 5407 1107
rect 5411 1103 5412 1107
rect 5406 1102 5412 1103
rect 5516 1100 5518 1161
rect 5620 1144 5622 1226
rect 5664 1167 5666 1235
rect 5663 1166 5667 1167
rect 5663 1161 5667 1162
rect 5618 1143 5624 1144
rect 5618 1139 5619 1143
rect 5623 1139 5624 1143
rect 5618 1138 5624 1139
rect 5602 1107 5608 1108
rect 5602 1103 5603 1107
rect 5607 1103 5608 1107
rect 5602 1102 5608 1103
rect 5514 1099 5520 1100
rect 5514 1095 5515 1099
rect 5519 1095 5520 1099
rect 5514 1094 5520 1095
rect 5542 1084 5548 1085
rect 5542 1080 5543 1084
rect 5547 1080 5548 1084
rect 5542 1079 5548 1080
rect 5544 1055 5546 1079
rect 5543 1054 5547 1055
rect 5543 1049 5547 1050
rect 5544 1025 5546 1049
rect 5542 1024 5548 1025
rect 5542 1020 5543 1024
rect 5547 1020 5548 1024
rect 5542 1019 5548 1020
rect 5514 1009 5520 1010
rect 5514 1005 5515 1009
rect 5519 1005 5520 1009
rect 5514 1004 5520 1005
rect 5370 999 5376 1000
rect 5370 995 5371 999
rect 5375 995 5376 999
rect 5370 994 5376 995
rect 5294 967 5300 968
rect 5294 963 5295 967
rect 5299 963 5300 967
rect 5294 962 5300 963
rect 4643 942 4647 943
rect 4643 937 4647 938
rect 4731 942 4735 943
rect 4731 937 4735 938
rect 4899 942 4903 943
rect 4899 937 4903 938
rect 4995 942 4999 943
rect 4995 937 4999 938
rect 5171 942 5175 943
rect 5171 937 5175 938
rect 5267 942 5271 943
rect 5267 937 5271 938
rect 4610 919 4616 920
rect 4610 915 4611 919
rect 4615 915 4616 919
rect 4610 914 4616 915
rect 4546 883 4552 884
rect 4546 879 4547 883
rect 4551 879 4552 883
rect 4546 878 4552 879
rect 4402 875 4408 876
rect 4402 871 4403 875
rect 4407 871 4408 875
rect 4402 870 4408 871
rect 4430 860 4436 861
rect 4430 856 4431 860
rect 4435 856 4436 860
rect 4430 855 4436 856
rect 4432 831 4434 855
rect 4279 830 4283 831
rect 4279 825 4283 826
rect 4431 830 4435 831
rect 4431 825 4435 826
rect 4280 801 4282 825
rect 4278 800 4284 801
rect 4278 796 4279 800
rect 4283 796 4284 800
rect 4278 795 4284 796
rect 4530 785 4536 786
rect 4530 781 4531 785
rect 4535 781 4536 785
rect 4530 780 4536 781
rect 4266 743 4272 744
rect 4266 739 4267 743
rect 4271 739 4272 743
rect 4266 738 4272 739
rect 4532 711 4534 780
rect 4548 744 4550 878
rect 4644 876 4646 937
rect 4866 919 4872 920
rect 4866 915 4867 919
rect 4871 915 4872 919
rect 4866 914 4872 915
rect 4868 880 4870 914
rect 4866 879 4872 880
rect 4642 875 4648 876
rect 4642 871 4643 875
rect 4647 871 4648 875
rect 4866 875 4867 879
rect 4871 875 4872 879
rect 4900 876 4902 937
rect 5172 876 5174 937
rect 5296 884 5298 962
rect 5516 943 5518 1004
rect 5604 968 5606 1102
rect 5664 1101 5666 1161
rect 5662 1100 5668 1101
rect 5662 1096 5663 1100
rect 5667 1096 5668 1100
rect 5662 1095 5668 1096
rect 5662 1083 5668 1084
rect 5662 1079 5663 1083
rect 5667 1079 5668 1083
rect 5662 1078 5668 1079
rect 5664 1055 5666 1078
rect 5663 1054 5667 1055
rect 5663 1049 5667 1050
rect 5664 1026 5666 1049
rect 5662 1025 5668 1026
rect 5662 1021 5663 1025
rect 5667 1021 5668 1025
rect 5662 1020 5668 1021
rect 5662 1008 5668 1009
rect 5662 1004 5663 1008
rect 5667 1004 5668 1008
rect 5662 1003 5668 1004
rect 5610 999 5616 1000
rect 5610 995 5611 999
rect 5615 995 5616 999
rect 5610 994 5616 995
rect 5602 967 5608 968
rect 5602 963 5603 967
rect 5607 963 5608 967
rect 5602 962 5608 963
rect 5443 942 5447 943
rect 5443 937 5447 938
rect 5515 942 5519 943
rect 5515 937 5519 938
rect 5294 883 5300 884
rect 5294 879 5295 883
rect 5299 879 5300 883
rect 5294 878 5300 879
rect 5444 876 5446 937
rect 5530 915 5536 916
rect 5530 911 5531 915
rect 5535 911 5536 915
rect 5530 910 5536 911
rect 4866 874 4872 875
rect 4898 875 4904 876
rect 4642 870 4648 871
rect 4898 871 4899 875
rect 4903 871 4904 875
rect 4898 870 4904 871
rect 5170 875 5176 876
rect 5170 871 5171 875
rect 5175 871 5176 875
rect 5170 870 5176 871
rect 5442 875 5448 876
rect 5442 871 5443 875
rect 5447 871 5448 875
rect 5442 870 5448 871
rect 4670 860 4676 861
rect 4670 856 4671 860
rect 4675 856 4676 860
rect 4670 855 4676 856
rect 4926 860 4932 861
rect 4926 856 4927 860
rect 4931 856 4932 860
rect 4926 855 4932 856
rect 5198 860 5204 861
rect 5198 856 5199 860
rect 5203 856 5204 860
rect 5198 855 5204 856
rect 5470 860 5476 861
rect 5470 856 5471 860
rect 5475 856 5476 860
rect 5470 855 5476 856
rect 4672 831 4674 855
rect 4928 831 4930 855
rect 5200 831 5202 855
rect 5472 831 5474 855
rect 4559 830 4563 831
rect 4559 825 4563 826
rect 4671 830 4675 831
rect 4671 825 4675 826
rect 4879 830 4883 831
rect 4879 825 4883 826
rect 4927 830 4931 831
rect 4927 825 4931 826
rect 5199 830 5203 831
rect 5199 825 5203 826
rect 5223 830 5227 831
rect 5223 825 5227 826
rect 5471 830 5475 831
rect 5471 825 5475 826
rect 4560 801 4562 825
rect 4880 801 4882 825
rect 5224 801 5226 825
rect 4558 800 4564 801
rect 4558 796 4559 800
rect 4563 796 4564 800
rect 4558 795 4564 796
rect 4878 800 4884 801
rect 4878 796 4879 800
rect 4883 796 4884 800
rect 4878 795 4884 796
rect 5222 800 5228 801
rect 5222 796 5223 800
rect 5227 796 5228 800
rect 5222 795 5228 796
rect 4850 785 4856 786
rect 4850 781 4851 785
rect 4855 781 4856 785
rect 4850 780 4856 781
rect 5194 785 5200 786
rect 5194 781 5195 785
rect 5199 781 5200 785
rect 5194 780 5200 781
rect 5514 785 5520 786
rect 5514 781 5515 785
rect 5519 781 5520 785
rect 5514 780 5520 781
rect 4546 743 4552 744
rect 4546 739 4547 743
rect 4551 739 4552 743
rect 4546 738 4552 739
rect 4852 711 4854 780
rect 4866 775 4872 776
rect 4866 771 4867 775
rect 4871 771 4872 775
rect 4866 770 4872 771
rect 4868 744 4870 770
rect 4866 743 4872 744
rect 4866 739 4867 743
rect 4871 739 4872 743
rect 4866 738 4872 739
rect 5196 711 5198 780
rect 5210 775 5216 776
rect 5210 771 5211 775
rect 5215 771 5216 775
rect 5210 770 5216 771
rect 5212 744 5214 770
rect 5210 743 5216 744
rect 5210 739 5211 743
rect 5215 739 5216 743
rect 5210 738 5216 739
rect 5516 711 5518 780
rect 5532 776 5534 910
rect 5543 830 5547 831
rect 5543 825 5547 826
rect 5544 801 5546 825
rect 5542 800 5548 801
rect 5542 796 5543 800
rect 5547 796 5548 800
rect 5542 795 5548 796
rect 5530 775 5536 776
rect 5530 771 5531 775
rect 5535 771 5536 775
rect 5530 770 5536 771
rect 5612 744 5614 994
rect 5664 943 5666 1003
rect 5663 942 5667 943
rect 5663 937 5667 938
rect 5664 877 5666 937
rect 5662 876 5668 877
rect 5662 872 5663 876
rect 5667 872 5668 876
rect 5662 871 5668 872
rect 5662 859 5668 860
rect 5662 855 5663 859
rect 5667 855 5668 859
rect 5662 854 5668 855
rect 5664 831 5666 854
rect 5663 830 5667 831
rect 5663 825 5667 826
rect 5664 802 5666 825
rect 5662 801 5668 802
rect 5662 797 5663 801
rect 5667 797 5668 801
rect 5662 796 5668 797
rect 5662 784 5668 785
rect 5662 780 5663 784
rect 5667 780 5668 784
rect 5662 779 5668 780
rect 5610 743 5616 744
rect 5610 739 5611 743
rect 5615 739 5616 743
rect 5610 738 5616 739
rect 5664 711 5666 779
rect 3995 710 3999 711
rect 3995 705 3999 706
rect 4019 710 4023 711
rect 4019 705 4023 706
rect 4131 710 4135 711
rect 4131 705 4135 706
rect 4251 710 4255 711
rect 4251 705 4255 706
rect 4267 710 4271 711
rect 4267 705 4271 706
rect 4403 710 4407 711
rect 4403 705 4407 706
rect 4531 710 4535 711
rect 4531 705 4535 706
rect 4571 710 4575 711
rect 4571 705 4575 706
rect 4771 710 4775 711
rect 4771 705 4775 706
rect 4851 710 4855 711
rect 4851 705 4855 706
rect 4995 710 4999 711
rect 4995 705 4999 706
rect 5195 710 5199 711
rect 5195 705 5199 706
rect 5227 710 5231 711
rect 5227 705 5231 706
rect 5459 710 5463 711
rect 5459 705 5463 706
rect 5515 710 5519 711
rect 5515 705 5519 706
rect 5663 710 5667 711
rect 5663 705 5667 706
rect 3986 687 3992 688
rect 3946 683 3952 684
rect 3946 679 3947 683
rect 3951 679 3952 683
rect 3986 683 3987 687
rect 3991 683 3992 687
rect 3986 682 3992 683
rect 3946 678 3952 679
rect 3866 651 3872 652
rect 3866 647 3867 651
rect 3871 647 3872 651
rect 3866 646 3872 647
rect 3838 640 3839 644
rect 3843 640 3844 644
rect 3838 639 3844 640
rect 3858 643 3864 644
rect 3858 639 3859 643
rect 3863 639 3864 643
rect 3858 638 3864 639
rect 3886 628 3892 629
rect 3838 627 3844 628
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3886 624 3887 628
rect 3891 624 3892 628
rect 3886 623 3892 624
rect 3838 622 3844 623
rect 3840 599 3842 622
rect 3888 599 3890 623
rect 3839 598 3843 599
rect 3839 593 3843 594
rect 3887 598 3891 599
rect 3887 593 3891 594
rect 3311 578 3315 579
rect 3311 573 3315 574
rect 3447 578 3451 579
rect 3447 573 3451 574
rect 3479 578 3483 579
rect 3479 573 3483 574
rect 3583 578 3587 579
rect 3583 573 3587 574
rect 3679 578 3683 579
rect 3679 573 3683 574
rect 3799 578 3803 579
rect 3799 573 3803 574
rect 3312 549 3314 573
rect 3448 549 3450 573
rect 3584 549 3586 573
rect 3800 550 3802 573
rect 3840 570 3842 593
rect 3838 569 3844 570
rect 3888 569 3890 593
rect 3838 565 3839 569
rect 3843 565 3844 569
rect 3838 564 3844 565
rect 3886 568 3892 569
rect 3886 564 3887 568
rect 3891 564 3892 568
rect 3886 563 3892 564
rect 3858 553 3864 554
rect 3838 552 3844 553
rect 3798 549 3804 550
rect 3310 548 3316 549
rect 3310 544 3311 548
rect 3315 544 3316 548
rect 3310 543 3316 544
rect 3446 548 3452 549
rect 3446 544 3447 548
rect 3451 544 3452 548
rect 3446 543 3452 544
rect 3582 548 3588 549
rect 3582 544 3583 548
rect 3587 544 3588 548
rect 3798 545 3799 549
rect 3803 545 3804 549
rect 3838 548 3839 552
rect 3843 548 3844 552
rect 3858 549 3859 553
rect 3863 549 3864 553
rect 3858 548 3864 549
rect 3838 547 3844 548
rect 3798 544 3804 545
rect 3582 543 3588 544
rect 3418 533 3424 534
rect 3418 529 3419 533
rect 3423 529 3424 533
rect 3418 528 3424 529
rect 3554 533 3560 534
rect 3554 529 3555 533
rect 3559 529 3560 533
rect 3554 528 3560 529
rect 3798 532 3804 533
rect 3798 528 3799 532
rect 3803 528 3804 532
rect 3298 491 3304 492
rect 3298 487 3299 491
rect 3303 487 3304 491
rect 3298 486 3304 487
rect 3420 467 3422 528
rect 3434 523 3440 524
rect 3434 519 3435 523
rect 3439 519 3440 523
rect 3434 518 3440 519
rect 3436 492 3438 518
rect 3434 491 3440 492
rect 3434 487 3435 491
rect 3439 487 3440 491
rect 3434 486 3440 487
rect 3556 467 3558 528
rect 3798 527 3804 528
rect 3570 523 3576 524
rect 3570 519 3571 523
rect 3575 519 3576 523
rect 3570 518 3576 519
rect 3642 523 3648 524
rect 3642 519 3643 523
rect 3647 519 3648 523
rect 3642 518 3648 519
rect 3572 492 3574 518
rect 3570 491 3576 492
rect 3570 487 3571 491
rect 3575 487 3576 491
rect 3570 486 3576 487
rect 1975 466 1979 467
rect 1975 461 1979 462
rect 1995 466 1999 467
rect 1995 461 1999 462
rect 2155 466 2159 467
rect 2155 461 2159 462
rect 2347 466 2351 467
rect 2347 461 2351 462
rect 2539 466 2543 467
rect 2539 461 2543 462
rect 2731 466 2735 467
rect 2731 461 2735 462
rect 2923 466 2927 467
rect 2923 461 2927 462
rect 3115 466 3119 467
rect 3115 461 3119 462
rect 3283 466 3287 467
rect 3283 461 3287 462
rect 3299 466 3303 467
rect 3299 461 3303 462
rect 3419 466 3423 467
rect 3419 461 3423 462
rect 3483 466 3487 467
rect 3483 461 3487 462
rect 3555 466 3559 467
rect 3555 461 3559 462
rect 1934 428 1940 429
rect 1786 427 1792 428
rect 1786 423 1787 427
rect 1791 423 1792 427
rect 1934 424 1935 428
rect 1939 424 1940 428
rect 1934 423 1940 424
rect 1786 422 1792 423
rect 1814 412 1820 413
rect 1814 408 1815 412
rect 1819 408 1820 412
rect 1814 407 1820 408
rect 1934 411 1940 412
rect 1934 407 1935 411
rect 1939 407 1940 411
rect 1816 367 1818 407
rect 1934 406 1940 407
rect 1936 367 1938 406
rect 1976 401 1978 461
rect 1974 400 1980 401
rect 1996 400 1998 461
rect 2156 400 2158 461
rect 2258 443 2264 444
rect 2258 439 2259 443
rect 2263 439 2264 443
rect 2258 438 2264 439
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 1994 399 2000 400
rect 1994 395 1995 399
rect 1999 395 2000 399
rect 1994 394 2000 395
rect 2154 399 2160 400
rect 2154 395 2155 399
rect 2159 395 2160 399
rect 2154 394 2160 395
rect 2022 384 2028 385
rect 1974 383 1980 384
rect 1974 379 1975 383
rect 1979 379 1980 383
rect 2022 380 2023 384
rect 2027 380 2028 384
rect 2022 379 2028 380
rect 2182 384 2188 385
rect 2182 380 2183 384
rect 2187 380 2188 384
rect 2182 379 2188 380
rect 1974 378 1980 379
rect 1815 366 1819 367
rect 1815 361 1819 362
rect 1935 366 1939 367
rect 1935 361 1939 362
rect 1936 338 1938 361
rect 1934 337 1940 338
rect 1934 333 1935 337
rect 1939 333 1940 337
rect 1934 332 1940 333
rect 1976 331 1978 378
rect 2024 331 2026 379
rect 2184 331 2186 379
rect 1975 330 1979 331
rect 1975 325 1979 326
rect 2023 330 2027 331
rect 2023 325 2027 326
rect 2047 330 2051 331
rect 2047 325 2051 326
rect 2183 330 2187 331
rect 2183 325 2187 326
rect 1934 320 1940 321
rect 1934 316 1935 320
rect 1939 316 1940 320
rect 1934 315 1940 316
rect 1518 279 1524 280
rect 1518 275 1519 279
rect 1523 275 1524 279
rect 1518 274 1524 275
rect 1936 223 1938 315
rect 1976 302 1978 325
rect 1974 301 1980 302
rect 2048 301 2050 325
rect 2184 301 2186 325
rect 1974 297 1975 301
rect 1979 297 1980 301
rect 1974 296 1980 297
rect 2046 300 2052 301
rect 2046 296 2047 300
rect 2051 296 2052 300
rect 2046 295 2052 296
rect 2182 300 2188 301
rect 2182 296 2183 300
rect 2187 296 2188 300
rect 2182 295 2188 296
rect 2018 285 2024 286
rect 1974 284 1980 285
rect 1974 280 1975 284
rect 1979 280 1980 284
rect 2018 281 2019 285
rect 2023 281 2024 285
rect 2018 280 2024 281
rect 2154 285 2160 286
rect 2154 281 2155 285
rect 2159 281 2160 285
rect 2154 280 2160 281
rect 1974 279 1980 280
rect 827 222 831 223
rect 827 217 831 218
rect 843 222 847 223
rect 843 217 847 218
rect 963 222 967 223
rect 963 217 967 218
rect 1003 222 1007 223
rect 1003 217 1007 218
rect 1099 222 1103 223
rect 1099 217 1103 218
rect 1935 222 1939 223
rect 1935 217 1939 218
rect 810 199 816 200
rect 810 195 811 199
rect 815 195 816 199
rect 810 194 816 195
rect 828 156 830 217
rect 964 156 966 217
rect 1100 156 1102 217
rect 1202 211 1208 212
rect 1202 207 1203 211
rect 1207 207 1208 211
rect 1202 206 1208 207
rect 1204 164 1206 206
rect 1202 163 1208 164
rect 1202 159 1203 163
rect 1207 159 1208 163
rect 1202 158 1208 159
rect 1936 157 1938 217
rect 1976 203 1978 279
rect 2020 203 2022 280
rect 2106 243 2112 244
rect 2106 239 2107 243
rect 2111 239 2112 243
rect 2106 238 2112 239
rect 1975 202 1979 203
rect 1975 197 1979 198
rect 1995 202 1999 203
rect 1995 197 1999 198
rect 2019 202 2023 203
rect 2019 197 2023 198
rect 1934 156 1940 157
rect 110 152 111 156
rect 115 152 116 156
rect 110 151 116 152
rect 146 155 152 156
rect 146 151 147 155
rect 151 151 152 155
rect 146 150 152 151
rect 282 155 288 156
rect 282 151 283 155
rect 287 151 288 155
rect 282 150 288 151
rect 418 155 424 156
rect 418 151 419 155
rect 423 151 424 155
rect 418 150 424 151
rect 554 155 560 156
rect 554 151 555 155
rect 559 151 560 155
rect 554 150 560 151
rect 690 155 696 156
rect 690 151 691 155
rect 695 151 696 155
rect 690 150 696 151
rect 826 155 832 156
rect 826 151 827 155
rect 831 151 832 155
rect 826 150 832 151
rect 962 155 968 156
rect 962 151 963 155
rect 967 151 968 155
rect 962 150 968 151
rect 1098 155 1104 156
rect 1098 151 1099 155
rect 1103 151 1104 155
rect 1934 152 1935 156
rect 1939 152 1940 156
rect 1934 151 1940 152
rect 1098 150 1104 151
rect 174 140 180 141
rect 110 139 116 140
rect 110 135 111 139
rect 115 135 116 139
rect 174 136 175 140
rect 179 136 180 140
rect 174 135 180 136
rect 310 140 316 141
rect 310 136 311 140
rect 315 136 316 140
rect 310 135 316 136
rect 446 140 452 141
rect 446 136 447 140
rect 451 136 452 140
rect 446 135 452 136
rect 582 140 588 141
rect 582 136 583 140
rect 587 136 588 140
rect 582 135 588 136
rect 718 140 724 141
rect 718 136 719 140
rect 723 136 724 140
rect 718 135 724 136
rect 854 140 860 141
rect 854 136 855 140
rect 859 136 860 140
rect 854 135 860 136
rect 990 140 996 141
rect 990 136 991 140
rect 995 136 996 140
rect 990 135 996 136
rect 1126 140 1132 141
rect 1126 136 1127 140
rect 1131 136 1132 140
rect 1126 135 1132 136
rect 1934 139 1940 140
rect 1934 135 1935 139
rect 1939 135 1940 139
rect 1976 137 1978 197
rect 110 134 116 135
rect 112 111 114 134
rect 176 111 178 135
rect 312 111 314 135
rect 448 111 450 135
rect 584 111 586 135
rect 720 111 722 135
rect 856 111 858 135
rect 992 111 994 135
rect 1128 111 1130 135
rect 1934 134 1940 135
rect 1974 136 1980 137
rect 1996 136 1998 197
rect 2108 144 2110 238
rect 2156 203 2158 280
rect 2260 276 2262 438
rect 2348 400 2350 461
rect 2474 443 2480 444
rect 2474 439 2475 443
rect 2479 439 2480 443
rect 2474 438 2480 439
rect 2476 408 2478 438
rect 2474 407 2480 408
rect 2474 403 2475 407
rect 2479 403 2480 407
rect 2474 402 2480 403
rect 2540 400 2542 461
rect 2666 443 2672 444
rect 2666 439 2667 443
rect 2671 439 2672 443
rect 2666 438 2672 439
rect 2668 408 2670 438
rect 2666 407 2672 408
rect 2666 403 2667 407
rect 2671 403 2672 407
rect 2666 402 2672 403
rect 2732 400 2734 461
rect 2854 427 2860 428
rect 2854 423 2855 427
rect 2859 423 2860 427
rect 2854 422 2860 423
rect 2856 408 2858 422
rect 2854 407 2860 408
rect 2854 403 2855 407
rect 2859 403 2860 407
rect 2854 402 2860 403
rect 2924 400 2926 461
rect 3050 443 3056 444
rect 3010 439 3016 440
rect 3010 435 3011 439
rect 3015 435 3016 439
rect 3050 439 3051 443
rect 3055 439 3056 443
rect 3050 438 3056 439
rect 3010 434 3016 435
rect 3012 416 3014 434
rect 3010 415 3016 416
rect 3010 411 3011 415
rect 3015 411 3016 415
rect 3010 410 3016 411
rect 3052 408 3054 438
rect 3050 407 3056 408
rect 3050 403 3051 407
rect 3055 403 3056 407
rect 3050 402 3056 403
rect 3116 400 3118 461
rect 3242 443 3248 444
rect 3242 439 3243 443
rect 3247 439 3248 443
rect 3242 438 3248 439
rect 3244 408 3246 438
rect 3242 407 3248 408
rect 3242 403 3243 407
rect 3247 403 3248 407
rect 3242 402 3248 403
rect 3300 400 3302 461
rect 3422 407 3428 408
rect 3422 403 3423 407
rect 3427 403 3428 407
rect 3422 402 3428 403
rect 2346 399 2352 400
rect 2346 395 2347 399
rect 2351 395 2352 399
rect 2346 394 2352 395
rect 2538 399 2544 400
rect 2538 395 2539 399
rect 2543 395 2544 399
rect 2538 394 2544 395
rect 2730 399 2736 400
rect 2730 395 2731 399
rect 2735 395 2736 399
rect 2730 394 2736 395
rect 2922 399 2928 400
rect 2922 395 2923 399
rect 2927 395 2928 399
rect 2922 394 2928 395
rect 3114 399 3120 400
rect 3114 395 3115 399
rect 3119 395 3120 399
rect 3114 394 3120 395
rect 3298 399 3304 400
rect 3298 395 3299 399
rect 3303 395 3304 399
rect 3298 394 3304 395
rect 2374 384 2380 385
rect 2374 380 2375 384
rect 2379 380 2380 384
rect 2374 379 2380 380
rect 2566 384 2572 385
rect 2566 380 2567 384
rect 2571 380 2572 384
rect 2566 379 2572 380
rect 2758 384 2764 385
rect 2758 380 2759 384
rect 2763 380 2764 384
rect 2758 379 2764 380
rect 2950 384 2956 385
rect 2950 380 2951 384
rect 2955 380 2956 384
rect 2950 379 2956 380
rect 3142 384 3148 385
rect 3142 380 3143 384
rect 3147 380 3148 384
rect 3142 379 3148 380
rect 3326 384 3332 385
rect 3326 380 3327 384
rect 3331 380 3332 384
rect 3326 379 3332 380
rect 2376 331 2378 379
rect 2568 331 2570 379
rect 2760 331 2762 379
rect 2952 331 2954 379
rect 3144 331 3146 379
rect 3328 331 3330 379
rect 2319 330 2323 331
rect 2319 325 2323 326
rect 2375 330 2379 331
rect 2375 325 2379 326
rect 2455 330 2459 331
rect 2455 325 2459 326
rect 2567 330 2571 331
rect 2567 325 2571 326
rect 2591 330 2595 331
rect 2591 325 2595 326
rect 2727 330 2731 331
rect 2727 325 2731 326
rect 2759 330 2763 331
rect 2759 325 2763 326
rect 2863 330 2867 331
rect 2863 325 2867 326
rect 2951 330 2955 331
rect 2951 325 2955 326
rect 2999 330 3003 331
rect 2999 325 3003 326
rect 3135 330 3139 331
rect 3135 325 3139 326
rect 3143 330 3147 331
rect 3143 325 3147 326
rect 3271 330 3275 331
rect 3271 325 3275 326
rect 3327 330 3331 331
rect 3327 325 3331 326
rect 3407 330 3411 331
rect 3407 325 3411 326
rect 2320 301 2322 325
rect 2456 301 2458 325
rect 2592 301 2594 325
rect 2728 301 2730 325
rect 2864 301 2866 325
rect 3000 301 3002 325
rect 3136 301 3138 325
rect 3272 301 3274 325
rect 3408 301 3410 325
rect 2318 300 2324 301
rect 2318 296 2319 300
rect 2323 296 2324 300
rect 2318 295 2324 296
rect 2454 300 2460 301
rect 2454 296 2455 300
rect 2459 296 2460 300
rect 2454 295 2460 296
rect 2590 300 2596 301
rect 2590 296 2591 300
rect 2595 296 2596 300
rect 2590 295 2596 296
rect 2726 300 2732 301
rect 2726 296 2727 300
rect 2731 296 2732 300
rect 2726 295 2732 296
rect 2862 300 2868 301
rect 2862 296 2863 300
rect 2867 296 2868 300
rect 2862 295 2868 296
rect 2998 300 3004 301
rect 2998 296 2999 300
rect 3003 296 3004 300
rect 2998 295 3004 296
rect 3134 300 3140 301
rect 3134 296 3135 300
rect 3139 296 3140 300
rect 3134 295 3140 296
rect 3270 300 3276 301
rect 3270 296 3271 300
rect 3275 296 3276 300
rect 3270 295 3276 296
rect 3406 300 3412 301
rect 3406 296 3407 300
rect 3411 296 3412 300
rect 3406 295 3412 296
rect 2290 285 2296 286
rect 2290 281 2291 285
rect 2295 281 2296 285
rect 2290 280 2296 281
rect 2426 285 2432 286
rect 2426 281 2427 285
rect 2431 281 2432 285
rect 2426 280 2432 281
rect 2562 285 2568 286
rect 2562 281 2563 285
rect 2567 281 2568 285
rect 2562 280 2568 281
rect 2698 285 2704 286
rect 2698 281 2699 285
rect 2703 281 2704 285
rect 2698 280 2704 281
rect 2834 285 2840 286
rect 2834 281 2835 285
rect 2839 281 2840 285
rect 2834 280 2840 281
rect 2970 285 2976 286
rect 2970 281 2971 285
rect 2975 281 2976 285
rect 2970 280 2976 281
rect 3106 285 3112 286
rect 3106 281 3107 285
rect 3111 281 3112 285
rect 3106 280 3112 281
rect 3242 285 3248 286
rect 3242 281 3243 285
rect 3247 281 3248 285
rect 3242 280 3248 281
rect 3378 285 3384 286
rect 3378 281 3379 285
rect 3383 281 3384 285
rect 3378 280 3384 281
rect 2258 275 2264 276
rect 2258 271 2259 275
rect 2263 271 2264 275
rect 2258 270 2264 271
rect 2292 203 2294 280
rect 2306 275 2312 276
rect 2306 271 2307 275
rect 2311 271 2312 275
rect 2306 270 2312 271
rect 2308 244 2310 270
rect 2306 243 2312 244
rect 2306 239 2307 243
rect 2311 239 2312 243
rect 2306 238 2312 239
rect 2428 203 2430 280
rect 2442 275 2448 276
rect 2442 271 2443 275
rect 2447 271 2448 275
rect 2442 270 2448 271
rect 2530 275 2536 276
rect 2530 271 2531 275
rect 2535 271 2536 275
rect 2530 270 2536 271
rect 2444 244 2446 270
rect 2442 243 2448 244
rect 2442 239 2443 243
rect 2447 239 2448 243
rect 2442 238 2448 239
rect 2131 202 2135 203
rect 2131 197 2135 198
rect 2155 202 2159 203
rect 2155 197 2159 198
rect 2267 202 2271 203
rect 2267 197 2271 198
rect 2291 202 2295 203
rect 2291 197 2295 198
rect 2403 202 2407 203
rect 2403 197 2407 198
rect 2427 202 2431 203
rect 2427 197 2431 198
rect 2106 143 2112 144
rect 2106 139 2107 143
rect 2111 139 2112 143
rect 2106 138 2112 139
rect 2132 136 2134 197
rect 2268 136 2270 197
rect 2404 136 2406 197
rect 2532 180 2534 270
rect 2564 203 2566 280
rect 2700 203 2702 280
rect 2836 203 2838 280
rect 2922 267 2928 268
rect 2922 263 2923 267
rect 2927 263 2928 267
rect 2922 262 2928 263
rect 2924 244 2926 262
rect 2842 243 2848 244
rect 2842 239 2843 243
rect 2847 239 2848 243
rect 2842 238 2848 239
rect 2922 243 2928 244
rect 2922 239 2923 243
rect 2927 239 2928 243
rect 2922 238 2928 239
rect 2539 202 2543 203
rect 2539 197 2543 198
rect 2563 202 2567 203
rect 2563 197 2567 198
rect 2675 202 2679 203
rect 2675 197 2679 198
rect 2699 202 2703 203
rect 2699 197 2703 198
rect 2811 202 2815 203
rect 2811 197 2815 198
rect 2835 202 2839 203
rect 2835 197 2839 198
rect 2530 179 2536 180
rect 2490 175 2496 176
rect 2490 171 2491 175
rect 2495 171 2496 175
rect 2530 175 2531 179
rect 2535 175 2536 179
rect 2530 174 2536 175
rect 2490 170 2496 171
rect 2492 152 2494 170
rect 2490 151 2496 152
rect 2490 147 2491 151
rect 2495 147 2496 151
rect 2490 146 2496 147
rect 2540 136 2542 197
rect 2676 136 2678 197
rect 2812 136 2814 197
rect 2844 152 2846 238
rect 2972 203 2974 280
rect 2986 275 2992 276
rect 2986 271 2987 275
rect 2991 271 2992 275
rect 2986 270 2992 271
rect 2988 244 2990 270
rect 2986 243 2992 244
rect 2986 239 2987 243
rect 2991 239 2992 243
rect 2986 238 2992 239
rect 3108 203 3110 280
rect 3122 275 3128 276
rect 3122 271 3123 275
rect 3127 271 3128 275
rect 3122 270 3128 271
rect 3234 275 3240 276
rect 3234 271 3235 275
rect 3239 271 3240 275
rect 3234 270 3240 271
rect 3124 244 3126 270
rect 3122 243 3128 244
rect 3122 239 3123 243
rect 3127 239 3128 243
rect 3122 238 3128 239
rect 2947 202 2951 203
rect 2947 197 2951 198
rect 2971 202 2975 203
rect 2971 197 2975 198
rect 3083 202 3087 203
rect 3083 197 3087 198
rect 3107 202 3111 203
rect 3107 197 3111 198
rect 3219 202 3223 203
rect 3219 197 3223 198
rect 2842 151 2848 152
rect 2842 147 2843 151
rect 2847 147 2848 151
rect 2842 146 2848 147
rect 2948 136 2950 197
rect 3084 136 3086 197
rect 3220 136 3222 197
rect 3236 196 3238 270
rect 3244 203 3246 280
rect 3330 267 3336 268
rect 3330 263 3331 267
rect 3335 263 3336 267
rect 3330 262 3336 263
rect 3332 244 3334 262
rect 3330 243 3336 244
rect 3330 239 3331 243
rect 3335 239 3336 243
rect 3330 238 3336 239
rect 3380 203 3382 280
rect 3424 244 3426 402
rect 3484 400 3486 461
rect 3644 444 3646 518
rect 3800 467 3802 527
rect 3840 475 3842 547
rect 3860 475 3862 548
rect 3948 544 3950 678
rect 3996 644 3998 705
rect 4132 644 4134 705
rect 4218 659 4224 660
rect 4218 655 4219 659
rect 4223 655 4224 659
rect 4218 654 4224 655
rect 3994 643 4000 644
rect 3994 639 3995 643
rect 3999 639 4000 643
rect 3994 638 4000 639
rect 4130 643 4136 644
rect 4130 639 4131 643
rect 4135 639 4136 643
rect 4130 638 4136 639
rect 4022 628 4028 629
rect 4022 624 4023 628
rect 4027 624 4028 628
rect 4022 623 4028 624
rect 4158 628 4164 629
rect 4158 624 4159 628
rect 4163 624 4164 628
rect 4158 623 4164 624
rect 4024 599 4026 623
rect 4160 599 4162 623
rect 4023 598 4027 599
rect 4023 593 4027 594
rect 4159 598 4163 599
rect 4159 593 4163 594
rect 4024 569 4026 593
rect 4160 569 4162 593
rect 4022 568 4028 569
rect 4022 564 4023 568
rect 4027 564 4028 568
rect 4022 563 4028 564
rect 4158 568 4164 569
rect 4158 564 4159 568
rect 4163 564 4164 568
rect 4158 563 4164 564
rect 3994 553 4000 554
rect 3994 549 3995 553
rect 3999 549 4000 553
rect 3994 548 4000 549
rect 4130 553 4136 554
rect 4130 549 4131 553
rect 4135 549 4136 553
rect 4130 548 4136 549
rect 3946 543 3952 544
rect 3946 539 3947 543
rect 3951 539 3952 543
rect 3946 538 3952 539
rect 3996 475 3998 548
rect 4002 543 4008 544
rect 4002 539 4003 543
rect 4007 539 4008 543
rect 4002 538 4008 539
rect 4004 512 4006 538
rect 4002 511 4008 512
rect 4002 507 4003 511
rect 4007 507 4008 511
rect 4002 506 4008 507
rect 4132 475 4134 548
rect 4220 512 4222 654
rect 4268 644 4270 705
rect 4404 644 4406 705
rect 4572 644 4574 705
rect 4698 687 4704 688
rect 4698 683 4699 687
rect 4703 683 4704 687
rect 4698 682 4704 683
rect 4700 652 4702 682
rect 4698 651 4704 652
rect 4698 647 4699 651
rect 4703 647 4704 651
rect 4698 646 4704 647
rect 4772 644 4774 705
rect 4898 687 4904 688
rect 4898 683 4899 687
rect 4903 683 4904 687
rect 4898 682 4904 683
rect 4900 652 4902 682
rect 4898 651 4904 652
rect 4898 647 4899 651
rect 4903 647 4904 651
rect 4898 646 4904 647
rect 4996 644 4998 705
rect 5122 687 5128 688
rect 5122 683 5123 687
rect 5127 683 5128 687
rect 5122 682 5128 683
rect 5124 652 5126 682
rect 5122 651 5128 652
rect 5122 647 5123 651
rect 5127 647 5128 651
rect 5122 646 5128 647
rect 5228 644 5230 705
rect 5334 651 5340 652
rect 5334 647 5335 651
rect 5339 647 5340 651
rect 5334 646 5340 647
rect 4266 643 4272 644
rect 4266 639 4267 643
rect 4271 639 4272 643
rect 4266 638 4272 639
rect 4402 643 4408 644
rect 4402 639 4403 643
rect 4407 639 4408 643
rect 4402 638 4408 639
rect 4570 643 4576 644
rect 4570 639 4571 643
rect 4575 639 4576 643
rect 4570 638 4576 639
rect 4770 643 4776 644
rect 4770 639 4771 643
rect 4775 639 4776 643
rect 4770 638 4776 639
rect 4994 643 5000 644
rect 4994 639 4995 643
rect 4999 639 5000 643
rect 4994 638 5000 639
rect 5226 643 5232 644
rect 5226 639 5227 643
rect 5231 639 5232 643
rect 5226 638 5232 639
rect 4294 628 4300 629
rect 4294 624 4295 628
rect 4299 624 4300 628
rect 4294 623 4300 624
rect 4430 628 4436 629
rect 4430 624 4431 628
rect 4435 624 4436 628
rect 4430 623 4436 624
rect 4598 628 4604 629
rect 4598 624 4599 628
rect 4603 624 4604 628
rect 4598 623 4604 624
rect 4798 628 4804 629
rect 4798 624 4799 628
rect 4803 624 4804 628
rect 4798 623 4804 624
rect 5022 628 5028 629
rect 5022 624 5023 628
rect 5027 624 5028 628
rect 5022 623 5028 624
rect 5254 628 5260 629
rect 5254 624 5255 628
rect 5259 624 5260 628
rect 5254 623 5260 624
rect 4296 599 4298 623
rect 4432 599 4434 623
rect 4600 599 4602 623
rect 4800 599 4802 623
rect 5024 599 5026 623
rect 5256 599 5258 623
rect 5336 612 5338 646
rect 5460 644 5462 705
rect 5546 683 5552 684
rect 5546 679 5547 683
rect 5551 679 5552 683
rect 5546 678 5552 679
rect 5458 643 5464 644
rect 5458 639 5459 643
rect 5463 639 5464 643
rect 5458 638 5464 639
rect 5486 628 5492 629
rect 5486 624 5487 628
rect 5491 624 5492 628
rect 5486 623 5492 624
rect 5334 611 5340 612
rect 5334 607 5335 611
rect 5339 607 5340 611
rect 5334 606 5340 607
rect 5488 599 5490 623
rect 4295 598 4299 599
rect 4295 593 4299 594
rect 4431 598 4435 599
rect 4431 593 4435 594
rect 4479 598 4483 599
rect 4479 593 4483 594
rect 4599 598 4603 599
rect 4599 593 4603 594
rect 4695 598 4699 599
rect 4695 593 4699 594
rect 4799 598 4803 599
rect 4799 593 4803 594
rect 4935 598 4939 599
rect 4935 593 4939 594
rect 5023 598 5027 599
rect 5023 593 5027 594
rect 5191 598 5195 599
rect 5191 593 5195 594
rect 5255 598 5259 599
rect 5255 593 5259 594
rect 5447 598 5451 599
rect 5447 593 5451 594
rect 5487 598 5491 599
rect 5487 593 5491 594
rect 4296 569 4298 593
rect 4480 569 4482 593
rect 4696 569 4698 593
rect 4936 569 4938 593
rect 5192 569 5194 593
rect 5448 569 5450 593
rect 4294 568 4300 569
rect 4294 564 4295 568
rect 4299 564 4300 568
rect 4294 563 4300 564
rect 4478 568 4484 569
rect 4478 564 4479 568
rect 4483 564 4484 568
rect 4478 563 4484 564
rect 4694 568 4700 569
rect 4694 564 4695 568
rect 4699 564 4700 568
rect 4694 563 4700 564
rect 4934 568 4940 569
rect 4934 564 4935 568
rect 4939 564 4940 568
rect 4934 563 4940 564
rect 5190 568 5196 569
rect 5190 564 5191 568
rect 5195 564 5196 568
rect 5190 563 5196 564
rect 5446 568 5452 569
rect 5446 564 5447 568
rect 5451 564 5452 568
rect 5446 563 5452 564
rect 4266 553 4272 554
rect 4266 549 4267 553
rect 4271 549 4272 553
rect 4266 548 4272 549
rect 4450 553 4456 554
rect 4450 549 4451 553
rect 4455 549 4456 553
rect 4450 548 4456 549
rect 4666 553 4672 554
rect 4666 549 4667 553
rect 4671 549 4672 553
rect 4666 548 4672 549
rect 4906 553 4912 554
rect 4906 549 4907 553
rect 4911 549 4912 553
rect 4906 548 4912 549
rect 5162 553 5168 554
rect 5162 549 5163 553
rect 5167 549 5168 553
rect 5162 548 5168 549
rect 5418 553 5424 554
rect 5418 549 5419 553
rect 5423 549 5424 553
rect 5418 548 5424 549
rect 4218 511 4224 512
rect 4218 507 4219 511
rect 4223 507 4224 511
rect 4218 506 4224 507
rect 4268 475 4270 548
rect 4452 475 4454 548
rect 4466 543 4472 544
rect 4466 539 4467 543
rect 4471 539 4472 543
rect 4466 538 4472 539
rect 4468 512 4470 538
rect 4466 511 4472 512
rect 4466 507 4467 511
rect 4471 507 4472 511
rect 4466 506 4472 507
rect 4570 495 4576 496
rect 4570 491 4571 495
rect 4575 491 4576 495
rect 4570 490 4576 491
rect 3839 474 3843 475
rect 3839 469 3843 470
rect 3859 474 3863 475
rect 3859 469 3863 470
rect 3995 474 3999 475
rect 3995 469 3999 470
rect 4131 474 4135 475
rect 4131 469 4135 470
rect 4267 474 4271 475
rect 4267 469 4271 470
rect 4451 474 4455 475
rect 4451 469 4455 470
rect 3651 466 3655 467
rect 3651 461 3655 462
rect 3799 466 3803 467
rect 3799 461 3803 462
rect 3634 443 3640 444
rect 3634 439 3635 443
rect 3639 439 3640 443
rect 3634 438 3640 439
rect 3642 443 3648 444
rect 3642 439 3643 443
rect 3647 439 3648 443
rect 3642 438 3648 439
rect 3636 408 3638 438
rect 3634 407 3640 408
rect 3634 403 3635 407
rect 3639 403 3640 407
rect 3634 402 3640 403
rect 3652 400 3654 461
rect 3800 401 3802 461
rect 3840 409 3842 469
rect 3838 408 3844 409
rect 4452 408 4454 469
rect 4572 452 4574 490
rect 4668 475 4670 548
rect 4682 543 4688 544
rect 4682 539 4683 543
rect 4687 539 4688 543
rect 4682 538 4688 539
rect 4684 512 4686 538
rect 4682 511 4688 512
rect 4682 507 4683 511
rect 4687 507 4688 511
rect 4682 506 4688 507
rect 4908 475 4910 548
rect 4922 543 4928 544
rect 4922 539 4923 543
rect 4927 539 4928 543
rect 4922 538 4928 539
rect 4924 512 4926 538
rect 4922 511 4928 512
rect 4922 507 4923 511
rect 4927 507 4928 511
rect 4922 506 4928 507
rect 5164 475 5166 548
rect 5178 543 5184 544
rect 5178 539 5179 543
rect 5183 539 5184 543
rect 5178 538 5184 539
rect 5186 543 5192 544
rect 5186 539 5187 543
rect 5191 539 5192 543
rect 5186 538 5192 539
rect 5180 512 5182 538
rect 5178 511 5184 512
rect 5178 507 5179 511
rect 5183 507 5184 511
rect 5178 506 5184 507
rect 5188 496 5190 538
rect 5186 495 5192 496
rect 5186 491 5187 495
rect 5191 491 5192 495
rect 5186 490 5192 491
rect 5420 475 5422 548
rect 5548 544 5550 678
rect 5594 651 5600 652
rect 5594 647 5595 651
rect 5599 647 5600 651
rect 5594 646 5600 647
rect 5546 543 5552 544
rect 5546 539 5547 543
rect 5551 539 5552 543
rect 5546 538 5552 539
rect 5434 511 5440 512
rect 5434 507 5435 511
rect 5439 507 5440 511
rect 5434 506 5440 507
rect 4651 474 4655 475
rect 4651 469 4655 470
rect 4667 474 4671 475
rect 4667 469 4671 470
rect 4859 474 4863 475
rect 4859 469 4863 470
rect 4907 474 4911 475
rect 4907 469 4911 470
rect 5067 474 5071 475
rect 5067 469 5071 470
rect 5163 474 5167 475
rect 5163 469 5167 470
rect 5283 474 5287 475
rect 5283 469 5287 470
rect 5419 474 5423 475
rect 5419 469 5423 470
rect 4570 451 4576 452
rect 4570 447 4571 451
rect 4575 447 4576 451
rect 4570 446 4576 447
rect 4578 451 4584 452
rect 4578 447 4579 451
rect 4583 447 4584 451
rect 4578 446 4584 447
rect 4580 416 4582 446
rect 4578 415 4584 416
rect 4578 411 4579 415
rect 4583 411 4584 415
rect 4578 410 4584 411
rect 4652 408 4654 469
rect 4778 451 4784 452
rect 4778 447 4779 451
rect 4783 447 4784 451
rect 4778 446 4784 447
rect 4780 416 4782 446
rect 4778 415 4784 416
rect 4778 411 4779 415
rect 4783 411 4784 415
rect 4778 410 4784 411
rect 4860 408 4862 469
rect 4986 451 4992 452
rect 4986 447 4987 451
rect 4991 447 4992 451
rect 4986 446 4992 447
rect 4988 416 4990 446
rect 4986 415 4992 416
rect 4986 411 4987 415
rect 4991 411 4992 415
rect 4986 410 4992 411
rect 5034 415 5040 416
rect 5034 411 5035 415
rect 5039 411 5040 415
rect 5034 410 5040 411
rect 3838 404 3839 408
rect 3843 404 3844 408
rect 3838 403 3844 404
rect 4450 407 4456 408
rect 4450 403 4451 407
rect 4455 403 4456 407
rect 4450 402 4456 403
rect 4650 407 4656 408
rect 4650 403 4651 407
rect 4655 403 4656 407
rect 4650 402 4656 403
rect 4858 407 4864 408
rect 4858 403 4859 407
rect 4863 403 4864 407
rect 4858 402 4864 403
rect 3798 400 3804 401
rect 3482 399 3488 400
rect 3482 395 3483 399
rect 3487 395 3488 399
rect 3482 394 3488 395
rect 3650 399 3656 400
rect 3650 395 3651 399
rect 3655 395 3656 399
rect 3798 396 3799 400
rect 3803 396 3804 400
rect 3798 395 3804 396
rect 3650 394 3656 395
rect 4478 392 4484 393
rect 3838 391 3844 392
rect 3838 387 3839 391
rect 3843 387 3844 391
rect 4478 388 4479 392
rect 4483 388 4484 392
rect 4478 387 4484 388
rect 4678 392 4684 393
rect 4678 388 4679 392
rect 4683 388 4684 392
rect 4678 387 4684 388
rect 4886 392 4892 393
rect 4886 388 4887 392
rect 4891 388 4892 392
rect 4886 387 4892 388
rect 3838 386 3844 387
rect 3510 384 3516 385
rect 3510 380 3511 384
rect 3515 380 3516 384
rect 3510 379 3516 380
rect 3678 384 3684 385
rect 3678 380 3679 384
rect 3683 380 3684 384
rect 3678 379 3684 380
rect 3798 383 3804 384
rect 3798 379 3799 383
rect 3803 379 3804 383
rect 3512 331 3514 379
rect 3680 331 3682 379
rect 3798 378 3804 379
rect 3800 331 3802 378
rect 3840 359 3842 386
rect 4480 359 4482 387
rect 4680 359 4682 387
rect 4888 359 4890 387
rect 3839 358 3843 359
rect 3839 353 3843 354
rect 4479 358 4483 359
rect 4479 353 4483 354
rect 4679 358 4683 359
rect 4679 353 4683 354
rect 4751 358 4755 359
rect 4751 353 4755 354
rect 4887 358 4891 359
rect 4887 353 4891 354
rect 4911 358 4915 359
rect 4911 353 4915 354
rect 3511 330 3515 331
rect 3511 325 3515 326
rect 3543 330 3547 331
rect 3543 325 3547 326
rect 3679 330 3683 331
rect 3679 325 3683 326
rect 3799 330 3803 331
rect 3840 330 3842 353
rect 3799 325 3803 326
rect 3838 329 3844 330
rect 4752 329 4754 353
rect 4912 329 4914 353
rect 3838 325 3839 329
rect 3843 325 3844 329
rect 3544 301 3546 325
rect 3680 301 3682 325
rect 3800 302 3802 325
rect 3838 324 3844 325
rect 4750 328 4756 329
rect 4750 324 4751 328
rect 4755 324 4756 328
rect 4750 323 4756 324
rect 4910 328 4916 329
rect 4910 324 4911 328
rect 4915 324 4916 328
rect 4910 323 4916 324
rect 4722 313 4728 314
rect 3838 312 3844 313
rect 3838 308 3839 312
rect 3843 308 3844 312
rect 4722 309 4723 313
rect 4727 309 4728 313
rect 4722 308 4728 309
rect 4882 313 4888 314
rect 4882 309 4883 313
rect 4887 309 4888 313
rect 4882 308 4888 309
rect 3838 307 3844 308
rect 3798 301 3804 302
rect 3542 300 3548 301
rect 3542 296 3543 300
rect 3547 296 3548 300
rect 3542 295 3548 296
rect 3678 300 3684 301
rect 3678 296 3679 300
rect 3683 296 3684 300
rect 3798 297 3799 301
rect 3803 297 3804 301
rect 3798 296 3804 297
rect 3678 295 3684 296
rect 3514 285 3520 286
rect 3514 281 3515 285
rect 3519 281 3520 285
rect 3514 280 3520 281
rect 3650 285 3656 286
rect 3650 281 3651 285
rect 3655 281 3656 285
rect 3650 280 3656 281
rect 3798 284 3804 285
rect 3798 280 3799 284
rect 3803 280 3804 284
rect 3422 243 3428 244
rect 3422 239 3423 243
rect 3427 239 3428 243
rect 3422 238 3428 239
rect 3516 203 3518 280
rect 3530 275 3536 276
rect 3530 271 3531 275
rect 3535 271 3536 275
rect 3530 270 3536 271
rect 3532 244 3534 270
rect 3530 243 3536 244
rect 3530 239 3531 243
rect 3535 239 3536 243
rect 3530 238 3536 239
rect 3652 203 3654 280
rect 3798 279 3804 280
rect 3666 275 3672 276
rect 3666 271 3667 275
rect 3671 271 3672 275
rect 3666 270 3672 271
rect 3668 244 3670 270
rect 3666 243 3672 244
rect 3666 239 3667 243
rect 3671 239 3672 243
rect 3666 238 3672 239
rect 3800 203 3802 279
rect 3840 207 3842 307
rect 4724 207 4726 308
rect 4858 303 4864 304
rect 4858 299 4859 303
rect 4863 299 4864 303
rect 4858 298 4864 299
rect 4860 272 4862 298
rect 4858 271 4864 272
rect 4858 267 4859 271
rect 4863 267 4864 271
rect 4858 266 4864 267
rect 4884 207 4886 308
rect 5036 272 5038 410
rect 5068 408 5070 469
rect 5284 408 5286 469
rect 5436 416 5438 506
rect 5507 474 5511 475
rect 5507 469 5511 470
rect 5434 415 5440 416
rect 5434 411 5435 415
rect 5439 411 5440 415
rect 5434 410 5440 411
rect 5508 408 5510 469
rect 5596 448 5598 646
rect 5664 645 5666 705
rect 5662 644 5668 645
rect 5662 640 5663 644
rect 5667 640 5668 644
rect 5662 639 5668 640
rect 5662 627 5668 628
rect 5662 623 5663 627
rect 5667 623 5668 627
rect 5662 622 5668 623
rect 5664 599 5666 622
rect 5663 598 5667 599
rect 5663 593 5667 594
rect 5664 570 5666 593
rect 5662 569 5668 570
rect 5662 565 5663 569
rect 5667 565 5668 569
rect 5662 564 5668 565
rect 5662 552 5668 553
rect 5662 548 5663 552
rect 5667 548 5668 552
rect 5662 547 5668 548
rect 5664 475 5666 547
rect 5663 474 5667 475
rect 5663 469 5667 470
rect 5594 447 5600 448
rect 5594 443 5595 447
rect 5599 443 5600 447
rect 5594 442 5600 443
rect 5602 415 5608 416
rect 5602 411 5603 415
rect 5607 411 5608 415
rect 5602 410 5608 411
rect 5066 407 5072 408
rect 5066 403 5067 407
rect 5071 403 5072 407
rect 5066 402 5072 403
rect 5282 407 5288 408
rect 5282 403 5283 407
rect 5287 403 5288 407
rect 5282 402 5288 403
rect 5506 407 5512 408
rect 5506 403 5507 407
rect 5511 403 5512 407
rect 5506 402 5512 403
rect 5094 392 5100 393
rect 5094 388 5095 392
rect 5099 388 5100 392
rect 5094 387 5100 388
rect 5310 392 5316 393
rect 5310 388 5311 392
rect 5315 388 5316 392
rect 5310 387 5316 388
rect 5534 392 5540 393
rect 5534 388 5535 392
rect 5539 388 5540 392
rect 5534 387 5540 388
rect 5096 359 5098 387
rect 5312 359 5314 387
rect 5536 359 5538 387
rect 5071 358 5075 359
rect 5071 353 5075 354
rect 5095 358 5099 359
rect 5095 353 5099 354
rect 5231 358 5235 359
rect 5231 353 5235 354
rect 5311 358 5315 359
rect 5311 353 5315 354
rect 5399 358 5403 359
rect 5399 353 5403 354
rect 5535 358 5539 359
rect 5535 353 5539 354
rect 5543 358 5547 359
rect 5543 353 5547 354
rect 5072 329 5074 353
rect 5232 329 5234 353
rect 5400 329 5402 353
rect 5544 329 5546 353
rect 5070 328 5076 329
rect 5070 324 5071 328
rect 5075 324 5076 328
rect 5070 323 5076 324
rect 5230 328 5236 329
rect 5230 324 5231 328
rect 5235 324 5236 328
rect 5230 323 5236 324
rect 5398 328 5404 329
rect 5398 324 5399 328
rect 5403 324 5404 328
rect 5398 323 5404 324
rect 5542 328 5548 329
rect 5542 324 5543 328
rect 5547 324 5548 328
rect 5542 323 5548 324
rect 5042 313 5048 314
rect 5042 309 5043 313
rect 5047 309 5048 313
rect 5042 308 5048 309
rect 5202 313 5208 314
rect 5202 309 5203 313
rect 5207 309 5208 313
rect 5202 308 5208 309
rect 5370 313 5376 314
rect 5370 309 5371 313
rect 5375 309 5376 313
rect 5370 308 5376 309
rect 5514 313 5520 314
rect 5514 309 5515 313
rect 5519 309 5520 313
rect 5514 308 5520 309
rect 5034 271 5040 272
rect 5034 267 5035 271
rect 5039 267 5040 271
rect 5034 266 5040 267
rect 5044 207 5046 308
rect 5130 295 5136 296
rect 5130 291 5131 295
rect 5135 291 5136 295
rect 5130 290 5136 291
rect 5132 272 5134 290
rect 5130 271 5136 272
rect 5130 267 5131 271
rect 5135 267 5136 271
rect 5130 266 5136 267
rect 5204 207 5206 308
rect 5218 303 5224 304
rect 5218 299 5219 303
rect 5223 299 5224 303
rect 5218 298 5224 299
rect 5220 272 5222 298
rect 5218 271 5224 272
rect 5218 267 5219 271
rect 5223 267 5224 271
rect 5218 266 5224 267
rect 5372 207 5374 308
rect 5386 271 5392 272
rect 5386 267 5387 271
rect 5391 267 5392 271
rect 5386 266 5392 267
rect 3839 206 3843 207
rect 3243 202 3247 203
rect 3243 197 3247 198
rect 3355 202 3359 203
rect 3355 197 3359 198
rect 3379 202 3383 203
rect 3379 197 3383 198
rect 3491 202 3495 203
rect 3491 197 3495 198
rect 3515 202 3519 203
rect 3515 197 3519 198
rect 3627 202 3631 203
rect 3627 197 3631 198
rect 3651 202 3655 203
rect 3651 197 3655 198
rect 3799 202 3803 203
rect 3839 201 3843 202
rect 4291 206 4295 207
rect 4291 201 4295 202
rect 4427 206 4431 207
rect 4427 201 4431 202
rect 4563 206 4567 207
rect 4563 201 4567 202
rect 4699 206 4703 207
rect 4699 201 4703 202
rect 4723 206 4727 207
rect 4723 201 4727 202
rect 4835 206 4839 207
rect 4835 201 4839 202
rect 4883 206 4887 207
rect 4883 201 4887 202
rect 4971 206 4975 207
rect 4971 201 4975 202
rect 5043 206 5047 207
rect 5043 201 5047 202
rect 5107 206 5111 207
rect 5107 201 5111 202
rect 5203 206 5207 207
rect 5203 201 5207 202
rect 5243 206 5247 207
rect 5243 201 5247 202
rect 5371 206 5375 207
rect 5371 201 5375 202
rect 5379 206 5383 207
rect 5379 201 5383 202
rect 3799 197 3803 198
rect 3234 195 3240 196
rect 3234 191 3235 195
rect 3239 191 3240 195
rect 3234 190 3240 191
rect 3306 175 3312 176
rect 3306 171 3307 175
rect 3311 171 3312 175
rect 3306 170 3312 171
rect 3308 152 3310 170
rect 3306 151 3312 152
rect 3306 147 3307 151
rect 3311 147 3312 151
rect 3306 146 3312 147
rect 3356 136 3358 197
rect 3492 136 3494 197
rect 3628 136 3630 197
rect 3800 137 3802 197
rect 3840 141 3842 201
rect 3838 140 3844 141
rect 4292 140 4294 201
rect 4428 140 4430 201
rect 4564 140 4566 201
rect 4700 140 4702 201
rect 4826 183 4832 184
rect 4826 179 4827 183
rect 4831 179 4832 183
rect 4826 178 4832 179
rect 4828 148 4830 178
rect 4826 147 4832 148
rect 4826 143 4827 147
rect 4831 143 4832 147
rect 4826 142 4832 143
rect 4836 140 4838 201
rect 4972 140 4974 201
rect 5108 140 5110 201
rect 5244 140 5246 201
rect 5380 140 5382 201
rect 5388 148 5390 266
rect 5516 207 5518 308
rect 5604 272 5606 410
rect 5664 409 5666 469
rect 5662 408 5668 409
rect 5662 404 5663 408
rect 5667 404 5668 408
rect 5662 403 5668 404
rect 5662 391 5668 392
rect 5662 387 5663 391
rect 5667 387 5668 391
rect 5662 386 5668 387
rect 5664 359 5666 386
rect 5663 358 5667 359
rect 5663 353 5667 354
rect 5664 330 5666 353
rect 5662 329 5668 330
rect 5662 325 5663 329
rect 5667 325 5668 329
rect 5662 324 5668 325
rect 5662 312 5668 313
rect 5662 308 5663 312
rect 5667 308 5668 312
rect 5662 307 5668 308
rect 5618 303 5624 304
rect 5618 299 5619 303
rect 5623 299 5624 303
rect 5618 298 5624 299
rect 5602 271 5608 272
rect 5602 267 5603 271
rect 5607 267 5608 271
rect 5602 266 5608 267
rect 5515 206 5519 207
rect 5515 201 5519 202
rect 5466 179 5472 180
rect 5466 175 5467 179
rect 5471 175 5472 179
rect 5466 174 5472 175
rect 5468 148 5470 174
rect 5386 147 5392 148
rect 5386 143 5387 147
rect 5391 143 5392 147
rect 5386 142 5392 143
rect 5466 147 5472 148
rect 5466 143 5467 147
rect 5471 143 5472 147
rect 5466 142 5472 143
rect 5516 140 5518 201
rect 5620 184 5622 298
rect 5664 207 5666 307
rect 5663 206 5667 207
rect 5663 201 5667 202
rect 5618 183 5624 184
rect 5618 179 5619 183
rect 5623 179 5624 183
rect 5618 178 5624 179
rect 5664 141 5666 201
rect 5662 140 5668 141
rect 3798 136 3804 137
rect 1936 111 1938 134
rect 1974 132 1975 136
rect 1979 132 1980 136
rect 1974 131 1980 132
rect 1994 135 2000 136
rect 1994 131 1995 135
rect 1999 131 2000 135
rect 1994 130 2000 131
rect 2130 135 2136 136
rect 2130 131 2131 135
rect 2135 131 2136 135
rect 2130 130 2136 131
rect 2266 135 2272 136
rect 2266 131 2267 135
rect 2271 131 2272 135
rect 2266 130 2272 131
rect 2402 135 2408 136
rect 2402 131 2403 135
rect 2407 131 2408 135
rect 2402 130 2408 131
rect 2538 135 2544 136
rect 2538 131 2539 135
rect 2543 131 2544 135
rect 2538 130 2544 131
rect 2674 135 2680 136
rect 2674 131 2675 135
rect 2679 131 2680 135
rect 2674 130 2680 131
rect 2810 135 2816 136
rect 2810 131 2811 135
rect 2815 131 2816 135
rect 2810 130 2816 131
rect 2946 135 2952 136
rect 2946 131 2947 135
rect 2951 131 2952 135
rect 2946 130 2952 131
rect 3082 135 3088 136
rect 3082 131 3083 135
rect 3087 131 3088 135
rect 3082 130 3088 131
rect 3218 135 3224 136
rect 3218 131 3219 135
rect 3223 131 3224 135
rect 3218 130 3224 131
rect 3354 135 3360 136
rect 3354 131 3355 135
rect 3359 131 3360 135
rect 3354 130 3360 131
rect 3490 135 3496 136
rect 3490 131 3491 135
rect 3495 131 3496 135
rect 3490 130 3496 131
rect 3626 135 3632 136
rect 3626 131 3627 135
rect 3631 131 3632 135
rect 3798 132 3799 136
rect 3803 132 3804 136
rect 3838 136 3839 140
rect 3843 136 3844 140
rect 3838 135 3844 136
rect 4290 139 4296 140
rect 4290 135 4291 139
rect 4295 135 4296 139
rect 4290 134 4296 135
rect 4426 139 4432 140
rect 4426 135 4427 139
rect 4431 135 4432 139
rect 4426 134 4432 135
rect 4562 139 4568 140
rect 4562 135 4563 139
rect 4567 135 4568 139
rect 4562 134 4568 135
rect 4698 139 4704 140
rect 4698 135 4699 139
rect 4703 135 4704 139
rect 4698 134 4704 135
rect 4834 139 4840 140
rect 4834 135 4835 139
rect 4839 135 4840 139
rect 4834 134 4840 135
rect 4970 139 4976 140
rect 4970 135 4971 139
rect 4975 135 4976 139
rect 4970 134 4976 135
rect 5106 139 5112 140
rect 5106 135 5107 139
rect 5111 135 5112 139
rect 5106 134 5112 135
rect 5242 139 5248 140
rect 5242 135 5243 139
rect 5247 135 5248 139
rect 5242 134 5248 135
rect 5378 139 5384 140
rect 5378 135 5379 139
rect 5383 135 5384 139
rect 5378 134 5384 135
rect 5514 139 5520 140
rect 5514 135 5515 139
rect 5519 135 5520 139
rect 5662 136 5663 140
rect 5667 136 5668 140
rect 5662 135 5668 136
rect 5514 134 5520 135
rect 3798 131 3804 132
rect 3626 130 3632 131
rect 4318 124 4324 125
rect 3838 123 3844 124
rect 2022 120 2028 121
rect 1974 119 1980 120
rect 1974 115 1975 119
rect 1979 115 1980 119
rect 2022 116 2023 120
rect 2027 116 2028 120
rect 2022 115 2028 116
rect 2158 120 2164 121
rect 2158 116 2159 120
rect 2163 116 2164 120
rect 2158 115 2164 116
rect 2294 120 2300 121
rect 2294 116 2295 120
rect 2299 116 2300 120
rect 2294 115 2300 116
rect 2430 120 2436 121
rect 2430 116 2431 120
rect 2435 116 2436 120
rect 2430 115 2436 116
rect 2566 120 2572 121
rect 2566 116 2567 120
rect 2571 116 2572 120
rect 2566 115 2572 116
rect 2702 120 2708 121
rect 2702 116 2703 120
rect 2707 116 2708 120
rect 2702 115 2708 116
rect 2838 120 2844 121
rect 2838 116 2839 120
rect 2843 116 2844 120
rect 2838 115 2844 116
rect 2974 120 2980 121
rect 2974 116 2975 120
rect 2979 116 2980 120
rect 2974 115 2980 116
rect 3110 120 3116 121
rect 3110 116 3111 120
rect 3115 116 3116 120
rect 3110 115 3116 116
rect 3246 120 3252 121
rect 3246 116 3247 120
rect 3251 116 3252 120
rect 3246 115 3252 116
rect 3382 120 3388 121
rect 3382 116 3383 120
rect 3387 116 3388 120
rect 3382 115 3388 116
rect 3518 120 3524 121
rect 3518 116 3519 120
rect 3523 116 3524 120
rect 3518 115 3524 116
rect 3654 120 3660 121
rect 3654 116 3655 120
rect 3659 116 3660 120
rect 3654 115 3660 116
rect 3798 119 3804 120
rect 3798 115 3799 119
rect 3803 115 3804 119
rect 3838 119 3839 123
rect 3843 119 3844 123
rect 4318 120 4319 124
rect 4323 120 4324 124
rect 4318 119 4324 120
rect 4454 124 4460 125
rect 4454 120 4455 124
rect 4459 120 4460 124
rect 4454 119 4460 120
rect 4590 124 4596 125
rect 4590 120 4591 124
rect 4595 120 4596 124
rect 4590 119 4596 120
rect 4726 124 4732 125
rect 4726 120 4727 124
rect 4731 120 4732 124
rect 4726 119 4732 120
rect 4862 124 4868 125
rect 4862 120 4863 124
rect 4867 120 4868 124
rect 4862 119 4868 120
rect 4998 124 5004 125
rect 4998 120 4999 124
rect 5003 120 5004 124
rect 4998 119 5004 120
rect 5134 124 5140 125
rect 5134 120 5135 124
rect 5139 120 5140 124
rect 5134 119 5140 120
rect 5270 124 5276 125
rect 5270 120 5271 124
rect 5275 120 5276 124
rect 5270 119 5276 120
rect 5406 124 5412 125
rect 5406 120 5407 124
rect 5411 120 5412 124
rect 5406 119 5412 120
rect 5542 124 5548 125
rect 5542 120 5543 124
rect 5547 120 5548 124
rect 5542 119 5548 120
rect 5662 123 5668 124
rect 5662 119 5663 123
rect 5667 119 5668 123
rect 3838 118 3844 119
rect 1974 114 1980 115
rect 111 110 115 111
rect 111 105 115 106
rect 175 110 179 111
rect 175 105 179 106
rect 311 110 315 111
rect 311 105 315 106
rect 447 110 451 111
rect 447 105 451 106
rect 583 110 587 111
rect 583 105 587 106
rect 719 110 723 111
rect 719 105 723 106
rect 855 110 859 111
rect 855 105 859 106
rect 991 110 995 111
rect 991 105 995 106
rect 1127 110 1131 111
rect 1127 105 1131 106
rect 1935 110 1939 111
rect 1935 105 1939 106
rect 1976 91 1978 114
rect 2024 91 2026 115
rect 2160 91 2162 115
rect 2296 91 2298 115
rect 2432 91 2434 115
rect 2568 91 2570 115
rect 2704 91 2706 115
rect 2840 91 2842 115
rect 2976 91 2978 115
rect 3112 91 3114 115
rect 3248 91 3250 115
rect 3384 91 3386 115
rect 3520 91 3522 115
rect 3656 91 3658 115
rect 3798 114 3804 115
rect 3800 91 3802 114
rect 3840 95 3842 118
rect 4320 95 4322 119
rect 4456 95 4458 119
rect 4592 95 4594 119
rect 4728 95 4730 119
rect 4864 95 4866 119
rect 5000 95 5002 119
rect 5136 95 5138 119
rect 5272 95 5274 119
rect 5408 95 5410 119
rect 5544 95 5546 119
rect 5662 118 5668 119
rect 5664 95 5666 118
rect 3839 94 3843 95
rect 1975 90 1979 91
rect 1975 85 1979 86
rect 2023 90 2027 91
rect 2023 85 2027 86
rect 2159 90 2163 91
rect 2159 85 2163 86
rect 2295 90 2299 91
rect 2295 85 2299 86
rect 2431 90 2435 91
rect 2431 85 2435 86
rect 2567 90 2571 91
rect 2567 85 2571 86
rect 2703 90 2707 91
rect 2703 85 2707 86
rect 2839 90 2843 91
rect 2839 85 2843 86
rect 2975 90 2979 91
rect 2975 85 2979 86
rect 3111 90 3115 91
rect 3111 85 3115 86
rect 3247 90 3251 91
rect 3247 85 3251 86
rect 3383 90 3387 91
rect 3383 85 3387 86
rect 3519 90 3523 91
rect 3519 85 3523 86
rect 3655 90 3659 91
rect 3655 85 3659 86
rect 3799 90 3803 91
rect 3839 89 3843 90
rect 4319 94 4323 95
rect 4319 89 4323 90
rect 4455 94 4459 95
rect 4455 89 4459 90
rect 4591 94 4595 95
rect 4591 89 4595 90
rect 4727 94 4731 95
rect 4727 89 4731 90
rect 4863 94 4867 95
rect 4863 89 4867 90
rect 4999 94 5003 95
rect 4999 89 5003 90
rect 5135 94 5139 95
rect 5135 89 5139 90
rect 5271 94 5275 95
rect 5271 89 5275 90
rect 5407 94 5411 95
rect 5407 89 5411 90
rect 5543 94 5547 95
rect 5543 89 5547 90
rect 5663 94 5667 95
rect 5663 89 5667 90
rect 3799 85 3803 86
<< m4c >>
rect 111 5754 115 5758
rect 131 5754 135 5758
rect 267 5754 271 5758
rect 403 5754 407 5758
rect 1935 5754 1939 5758
rect 111 5642 115 5646
rect 159 5642 163 5646
rect 295 5642 299 5646
rect 343 5642 347 5646
rect 1975 5686 1979 5690
rect 1995 5686 1999 5690
rect 2171 5686 2175 5690
rect 2371 5686 2375 5690
rect 2563 5686 2567 5690
rect 2747 5686 2751 5690
rect 2931 5686 2935 5690
rect 3107 5686 3111 5690
rect 3275 5686 3279 5690
rect 3443 5686 3447 5690
rect 3619 5686 3623 5690
rect 3799 5686 3803 5690
rect 3839 5690 3843 5694
rect 4467 5690 4471 5694
rect 4603 5690 4607 5694
rect 4739 5690 4743 5694
rect 4875 5690 4879 5694
rect 5663 5690 5667 5694
rect 431 5642 435 5646
rect 535 5642 539 5646
rect 735 5642 739 5646
rect 943 5642 947 5646
rect 1159 5642 1163 5646
rect 1383 5642 1387 5646
rect 1607 5642 1611 5646
rect 1815 5642 1819 5646
rect 1935 5642 1939 5646
rect 111 5530 115 5534
rect 315 5530 319 5534
rect 507 5530 511 5534
rect 707 5530 711 5534
rect 875 5530 879 5534
rect 915 5530 919 5534
rect 1975 5574 1979 5578
rect 2023 5574 2027 5578
rect 2199 5574 2203 5578
rect 2375 5574 2379 5578
rect 2399 5574 2403 5578
rect 2591 5574 2595 5578
rect 2607 5574 2611 5578
rect 1011 5530 1015 5534
rect 1131 5530 1135 5534
rect 1147 5530 1151 5534
rect 1291 5530 1295 5534
rect 1355 5530 1359 5534
rect 1435 5530 1439 5534
rect 1579 5530 1583 5534
rect 1723 5530 1727 5534
rect 1787 5530 1791 5534
rect 111 5418 115 5422
rect 719 5418 723 5422
rect 855 5418 859 5422
rect 903 5418 907 5422
rect 991 5418 995 5422
rect 1039 5418 1043 5422
rect 1127 5418 1131 5422
rect 1175 5418 1179 5422
rect 1263 5418 1267 5422
rect 111 5306 115 5310
rect 691 5306 695 5310
rect 723 5306 727 5310
rect 1319 5418 1323 5422
rect 1399 5418 1403 5422
rect 1463 5418 1467 5422
rect 1535 5418 1539 5422
rect 827 5306 831 5310
rect 875 5306 879 5310
rect 963 5306 967 5310
rect 1027 5306 1031 5310
rect 1099 5306 1103 5310
rect 1187 5306 1191 5310
rect 1235 5306 1239 5310
rect 1355 5306 1359 5310
rect 1371 5306 1375 5310
rect 111 5194 115 5198
rect 447 5194 451 5198
rect 623 5194 627 5198
rect 751 5194 755 5198
rect 807 5194 811 5198
rect 903 5194 907 5198
rect 999 5194 1003 5198
rect 1055 5194 1059 5198
rect 1199 5194 1203 5198
rect 1215 5194 1219 5198
rect 111 5074 115 5078
rect 155 5074 159 5078
rect 379 5074 383 5078
rect 419 5074 423 5078
rect 595 5074 599 5078
rect 627 5074 631 5078
rect 111 4934 115 4938
rect 159 4934 163 4938
rect 183 4934 187 4938
rect 295 4934 299 4938
rect 407 4934 411 4938
rect 431 4934 435 4938
rect 111 4810 115 4814
rect 131 4810 135 4814
rect 1935 5530 1939 5534
rect 1975 5458 1979 5462
rect 2347 5458 2351 5462
rect 1607 5418 1611 5422
rect 1671 5418 1675 5422
rect 1751 5418 1755 5422
rect 1807 5418 1811 5422
rect 1935 5418 1939 5422
rect 1975 5346 1979 5350
rect 2319 5346 2323 5350
rect 1507 5306 1511 5310
rect 1523 5306 1527 5310
rect 1643 5306 1647 5310
rect 1779 5306 1783 5310
rect 1935 5306 1939 5310
rect 1383 5194 1387 5198
rect 1399 5194 1403 5198
rect 1551 5194 1555 5198
rect 1607 5194 1611 5198
rect 779 5074 783 5078
rect 899 5074 903 5078
rect 971 5074 975 5078
rect 1171 5074 1175 5078
rect 1195 5074 1199 5078
rect 1371 5074 1375 5078
rect 2775 5574 2779 5578
rect 2831 5574 2835 5578
rect 2959 5574 2963 5578
rect 3047 5574 3051 5578
rect 2451 5458 2455 5462
rect 2579 5458 2583 5462
rect 2699 5458 2703 5462
rect 2803 5458 2807 5462
rect 3135 5574 3139 5578
rect 3263 5574 3267 5578
rect 3303 5574 3307 5578
rect 3471 5574 3475 5578
rect 3479 5574 3483 5578
rect 3647 5574 3651 5578
rect 3679 5574 3683 5578
rect 2947 5458 2951 5462
rect 3019 5458 3023 5462
rect 3187 5458 3191 5462
rect 3235 5458 3239 5462
rect 3427 5458 3431 5462
rect 3451 5458 3455 5462
rect 2479 5346 2483 5350
rect 2519 5346 2523 5350
rect 2719 5346 2723 5350
rect 2727 5346 2731 5350
rect 2919 5346 2923 5350
rect 2975 5346 2979 5350
rect 1975 5230 1979 5234
rect 2275 5230 2279 5234
rect 2291 5230 2295 5234
rect 2475 5230 2479 5234
rect 2491 5230 2495 5234
rect 1815 5194 1819 5198
rect 1935 5194 1939 5198
rect 3799 5574 3803 5578
rect 3839 5578 3843 5582
rect 4431 5578 4435 5582
rect 4495 5578 4499 5582
rect 4567 5578 4571 5582
rect 4631 5578 4635 5582
rect 4703 5578 4707 5582
rect 4767 5578 4771 5582
rect 4839 5578 4843 5582
rect 4903 5578 4907 5582
rect 3839 5466 3843 5470
rect 4403 5466 4407 5470
rect 4427 5466 4431 5470
rect 4539 5466 4543 5470
rect 4587 5466 4591 5470
rect 3651 5458 3655 5462
rect 3799 5458 3803 5462
rect 3119 5346 3123 5350
rect 3215 5346 3219 5350
rect 3327 5346 3331 5350
rect 3455 5346 3459 5350
rect 3535 5346 3539 5350
rect 2683 5230 2687 5234
rect 2691 5230 2695 5234
rect 2891 5230 2895 5234
rect 1975 5102 1979 5106
rect 2119 5102 2123 5106
rect 2303 5102 2307 5106
rect 2327 5102 2331 5106
rect 1499 5074 1503 5078
rect 1579 5074 1583 5078
rect 1787 5074 1791 5078
rect 1935 5074 1939 5078
rect 2503 5102 2507 5106
rect 2535 5102 2539 5106
rect 2711 5102 2715 5106
rect 2751 5102 2755 5106
rect 3091 5230 3095 5234
rect 3099 5230 3103 5234
rect 3299 5230 3303 5234
rect 3307 5230 3311 5234
rect 2919 5102 2923 5106
rect 2975 5102 2979 5106
rect 1975 4982 1979 4986
rect 1995 4982 1999 4986
rect 2091 4982 2095 4986
rect 2131 4982 2135 4986
rect 2267 4982 2271 4986
rect 2299 4982 2303 4986
rect 2419 4982 2423 4986
rect 2507 4982 2511 4986
rect 2619 4982 2623 4986
rect 2723 4982 2727 4986
rect 567 4934 571 4938
rect 655 4934 659 4938
rect 703 4934 707 4938
rect 927 4934 931 4938
rect 1223 4934 1227 4938
rect 1527 4934 1531 4938
rect 1815 4934 1819 4938
rect 1935 4934 1939 4938
rect 3679 5346 3683 5350
rect 3799 5346 3803 5350
rect 3839 5346 3843 5350
rect 4431 5346 4435 5350
rect 4455 5346 4459 5350
rect 3507 5230 3511 5234
rect 3799 5230 3803 5234
rect 4675 5466 4679 5470
rect 4747 5466 4751 5470
rect 4811 5466 4815 5470
rect 4975 5578 4979 5582
rect 5111 5578 5115 5582
rect 5663 5578 5667 5582
rect 4907 5466 4911 5470
rect 4947 5466 4951 5470
rect 5075 5466 5079 5470
rect 5083 5466 5087 5470
rect 5663 5466 5667 5470
rect 4615 5346 4619 5350
rect 4775 5346 4779 5350
rect 4799 5346 4803 5350
rect 4935 5346 4939 5350
rect 4983 5346 4987 5350
rect 5103 5346 5107 5350
rect 5175 5346 5179 5350
rect 3839 5218 3843 5222
rect 4403 5218 4407 5222
rect 4435 5218 4439 5222
rect 4587 5218 4591 5222
rect 4595 5218 4599 5222
rect 3127 5102 3131 5106
rect 3207 5102 3211 5106
rect 3335 5102 3339 5106
rect 3799 5102 3803 5106
rect 3839 5098 3843 5102
rect 3887 5098 3891 5102
rect 4087 5098 4091 5102
rect 4327 5098 4331 5102
rect 2859 4982 2863 4986
rect 2947 4982 2951 4986
rect 3123 4982 3127 4986
rect 3179 4982 3183 4986
rect 1975 4862 1979 4866
rect 2023 4862 2027 4866
rect 2159 4862 2163 4866
rect 2295 4862 2299 4866
rect 2327 4862 2331 4866
rect 2447 4862 2451 4866
rect 2559 4862 2563 4866
rect 2647 4862 2651 4866
rect 2823 4862 2827 4866
rect 2887 4862 2891 4866
rect 267 4810 271 4814
rect 403 4810 407 4814
rect 539 4810 543 4814
rect 675 4810 679 4814
rect 1935 4810 1939 4814
rect 111 4694 115 4698
rect 159 4694 163 4698
rect 1975 4738 1979 4742
rect 2019 4738 2023 4742
rect 2195 4738 2199 4742
rect 2299 4738 2303 4742
rect 2371 4738 2375 4742
rect 295 4694 299 4698
rect 431 4694 435 4698
rect 567 4694 571 4698
rect 703 4694 707 4698
rect 1935 4694 1939 4698
rect 111 4570 115 4574
rect 131 4570 135 4574
rect 251 4570 255 4574
rect 267 4570 271 4574
rect 403 4570 407 4574
rect 443 4570 447 4574
rect 539 4570 543 4574
rect 651 4570 655 4574
rect 675 4570 679 4574
rect 111 4458 115 4462
rect 279 4458 283 4462
rect 471 4458 475 4462
rect 511 4458 515 4462
rect 1975 4622 1979 4626
rect 2023 4622 2027 4626
rect 2047 4622 2051 4626
rect 875 4570 879 4574
rect 1099 4570 1103 4574
rect 1331 4570 1335 4574
rect 1571 4570 1575 4574
rect 1787 4570 1791 4574
rect 1935 4570 1939 4574
rect 679 4458 683 4462
rect 687 4458 691 4462
rect 871 4458 875 4462
rect 903 4458 907 4462
rect 1071 4458 1075 4462
rect 1127 4458 1131 4462
rect 1279 4458 1283 4462
rect 1359 4458 1363 4462
rect 1495 4458 1499 4462
rect 111 4342 115 4346
rect 483 4342 487 4346
rect 659 4342 663 4346
rect 715 4342 719 4346
rect 843 4342 847 4346
rect 851 4342 855 4346
rect 987 4342 991 4346
rect 1043 4342 1047 4346
rect 1123 4342 1127 4346
rect 1251 4342 1255 4346
rect 1259 4342 1263 4346
rect 2531 4738 2535 4742
rect 2547 4738 2551 4742
rect 3395 4982 3399 4986
rect 3651 4982 3655 4986
rect 3799 4982 3803 4986
rect 3839 4986 3843 4990
rect 3859 4986 3863 4990
rect 3995 4986 3999 4990
rect 4059 4986 4063 4990
rect 3103 4862 3107 4866
rect 3151 4862 3155 4866
rect 3399 4862 3403 4866
rect 3423 4862 3427 4866
rect 3679 4862 3683 4866
rect 4131 4986 4135 4990
rect 5663 5346 5667 5350
rect 4755 5218 4759 5222
rect 4771 5218 4775 5222
rect 4915 5218 4919 5222
rect 4955 5218 4959 5222
rect 5067 5218 5071 5222
rect 5147 5218 5151 5222
rect 5219 5218 5223 5222
rect 5379 5218 5383 5222
rect 5515 5218 5519 5222
rect 5663 5218 5667 5222
rect 4463 5098 4467 5102
rect 4567 5098 4571 5102
rect 4623 5098 4627 5102
rect 4783 5098 4787 5102
rect 4815 5098 4819 5102
rect 4943 5098 4947 5102
rect 5063 5098 5067 5102
rect 5095 5098 5099 5102
rect 5247 5098 5251 5102
rect 5311 5098 5315 5102
rect 5407 5098 5411 5102
rect 5543 5098 5547 5102
rect 4267 4986 4271 4990
rect 4299 4986 4303 4990
rect 4403 4986 4407 4990
rect 4539 4986 4543 4990
rect 4675 4986 4679 4990
rect 4787 4986 4791 4990
rect 4811 4986 4815 4990
rect 4947 4986 4951 4990
rect 5035 4986 5039 4990
rect 5083 4986 5087 4990
rect 5227 4986 5231 4990
rect 5283 4986 5287 4990
rect 4875 4968 4879 4972
rect 5239 4968 5243 4972
rect 5663 5098 5667 5102
rect 5379 4986 5383 4990
rect 5515 4986 5519 4990
rect 5663 4986 5667 4990
rect 3799 4862 3803 4866
rect 3839 4798 3843 4802
rect 3887 4798 3891 4802
rect 4023 4798 4027 4802
rect 4071 4798 4075 4802
rect 4159 4798 4163 4802
rect 4295 4798 4299 4802
rect 4431 4798 4435 4802
rect 4535 4798 4539 4802
rect 4567 4798 4571 4802
rect 4703 4798 4707 4802
rect 4783 4798 4787 4802
rect 4839 4798 4843 4802
rect 4975 4798 4979 4802
rect 5039 4798 5043 4802
rect 5111 4798 5115 4802
rect 5255 4798 5259 4802
rect 5303 4798 5307 4802
rect 5407 4798 5411 4802
rect 5543 4798 5547 4802
rect 2723 4738 2727 4742
rect 2795 4738 2799 4742
rect 3075 4738 3079 4742
rect 3371 4738 3375 4742
rect 3651 4738 3655 4742
rect 3799 4738 3803 4742
rect 2223 4622 2227 4626
rect 2263 4622 2267 4626
rect 2399 4622 2403 4626
rect 2527 4622 2531 4626
rect 2575 4622 2579 4626
rect 2751 4622 2755 4626
rect 2775 4622 2779 4626
rect 1975 4498 1979 4502
rect 1995 4498 1999 4502
rect 2235 4498 2239 4502
rect 2267 4498 2271 4502
rect 2499 4498 2503 4502
rect 2515 4498 2519 4502
rect 1599 4458 1603 4462
rect 1719 4458 1723 4462
rect 1815 4458 1819 4462
rect 1935 4458 1939 4462
rect 1395 4342 1399 4346
rect 1467 4342 1471 4346
rect 1531 4342 1535 4346
rect 1667 4342 1671 4346
rect 1691 4342 1695 4346
rect 111 4222 115 4226
rect 727 4222 731 4226
rect 743 4222 747 4226
rect 863 4222 867 4226
rect 879 4222 883 4226
rect 999 4222 1003 4226
rect 1015 4222 1019 4226
rect 1135 4222 1139 4226
rect 1151 4222 1155 4226
rect 1271 4222 1275 4226
rect 1287 4222 1291 4226
rect 111 4110 115 4114
rect 563 4110 567 4114
rect 699 4110 703 4114
rect 835 4110 839 4114
rect 1407 4222 1411 4226
rect 1423 4222 1427 4226
rect 1543 4222 1547 4226
rect 1559 4222 1563 4226
rect 971 4110 975 4114
rect 1107 4110 1111 4114
rect 1243 4110 1247 4114
rect 1379 4110 1383 4114
rect 111 3998 115 4002
rect 159 3998 163 4002
rect 327 3998 331 4002
rect 535 3998 539 4002
rect 591 3998 595 4002
rect 727 3998 731 4002
rect 751 3998 755 4002
rect 863 3998 867 4002
rect 111 3886 115 3890
rect 131 3886 135 3890
rect 1975 4374 1979 4378
rect 2023 4374 2027 4378
rect 2199 4374 2203 4378
rect 2295 4374 2299 4378
rect 1935 4342 1939 4346
rect 1975 4258 1979 4262
rect 1995 4258 1999 4262
rect 1679 4222 1683 4226
rect 1695 4222 1699 4226
rect 1815 4222 1819 4226
rect 1935 4222 1939 4226
rect 1515 4110 1519 4114
rect 1651 4110 1655 4114
rect 967 3998 971 4002
rect 999 3998 1003 4002
rect 1135 3998 1139 4002
rect 1183 3998 1187 4002
rect 1271 3998 1275 4002
rect 1399 3998 1403 4002
rect 1407 3998 1411 4002
rect 299 3886 303 3890
rect 355 3886 359 3890
rect 507 3886 511 3890
rect 619 3886 623 3890
rect 723 3886 727 3890
rect 899 3886 903 3890
rect 939 3886 943 3890
rect 1155 3886 1159 3890
rect 1195 3886 1199 3890
rect 111 3762 115 3766
rect 159 3762 163 3766
rect 247 3762 251 3766
rect 383 3762 387 3766
rect 519 3762 523 3766
rect 647 3762 651 3766
rect 791 3762 795 3766
rect 111 3634 115 3638
rect 219 3634 223 3638
rect 491 3634 495 3638
rect 1543 3998 1547 4002
rect 1615 3998 1619 4002
rect 3839 4686 3843 4690
rect 3859 4686 3863 4690
rect 3995 4686 3999 4690
rect 4043 4686 4047 4690
rect 4131 4686 4135 4690
rect 3015 4622 3019 4626
rect 3247 4622 3251 4626
rect 3471 4622 3475 4626
rect 3679 4622 3683 4626
rect 2747 4498 2751 4502
rect 2971 4498 2975 4502
rect 2987 4498 2991 4502
rect 2399 4374 2403 4378
rect 2543 4374 2547 4378
rect 2591 4374 2595 4378
rect 2775 4374 2779 4378
rect 2171 4258 2175 4262
rect 2243 4258 2247 4262
rect 2371 4258 2375 4262
rect 2507 4258 2511 4262
rect 2563 4258 2567 4262
rect 3799 4622 3803 4626
rect 4267 4686 4271 4690
rect 4403 4686 4407 4690
rect 4507 4686 4511 4690
rect 4539 4686 4543 4690
rect 4675 4686 4679 4690
rect 4755 4686 4759 4690
rect 4819 4686 4823 4690
rect 4963 4686 4967 4690
rect 5011 4686 5015 4690
rect 5107 4686 5111 4690
rect 5243 4686 5247 4690
rect 5275 4686 5279 4690
rect 3839 4574 3843 4578
rect 3887 4574 3891 4578
rect 4023 4574 4027 4578
rect 4159 4574 4163 4578
rect 4295 4574 4299 4578
rect 4431 4574 4435 4578
rect 4567 4574 4571 4578
rect 3187 4498 3191 4502
rect 3219 4498 3223 4502
rect 3395 4498 3399 4502
rect 3443 4498 3447 4502
rect 3611 4498 3615 4502
rect 3651 4498 3655 4502
rect 3799 4498 3803 4502
rect 3075 4488 3079 4492
rect 3735 4488 3739 4492
rect 5663 4798 5667 4802
rect 5379 4686 5383 4690
rect 5515 4686 5519 4690
rect 5663 4686 5667 4690
rect 4671 4574 4675 4578
rect 4703 4574 4707 4578
rect 4807 4574 4811 4578
rect 4847 4574 4851 4578
rect 4943 4574 4947 4578
rect 4991 4574 4995 4578
rect 5079 4574 5083 4578
rect 5135 4574 5139 4578
rect 5271 4574 5275 4578
rect 5407 4574 5411 4578
rect 5543 4574 5547 4578
rect 5663 4574 5667 4578
rect 3839 4458 3843 4462
rect 4347 4458 4351 4462
rect 4483 4458 4487 4462
rect 4619 4458 4623 4462
rect 4643 4458 4647 4462
rect 4755 4458 4759 4462
rect 4779 4458 4783 4462
rect 4891 4458 4895 4462
rect 4915 4458 4919 4462
rect 5051 4458 5055 4462
rect 2951 4374 2955 4378
rect 2999 4374 3003 4378
rect 3135 4374 3139 4378
rect 3215 4374 3219 4378
rect 3319 4374 3323 4378
rect 3423 4374 3427 4378
rect 3639 4374 3643 4378
rect 3799 4374 3803 4378
rect 3839 4330 3843 4334
rect 4135 4330 4139 4334
rect 4271 4330 4275 4334
rect 4375 4330 4379 4334
rect 4407 4330 4411 4334
rect 2747 4258 2751 4262
rect 2763 4258 2767 4262
rect 2923 4258 2927 4262
rect 3019 4258 3023 4262
rect 3107 4258 3111 4262
rect 3283 4258 3287 4262
rect 3291 4258 3295 4262
rect 3799 4258 3803 4262
rect 1975 4134 1979 4138
rect 2023 4134 2027 4138
rect 2271 4134 2275 4138
rect 2535 4134 2539 4138
rect 2791 4134 2795 4138
rect 3047 4134 3051 4138
rect 3135 4134 3139 4138
rect 3271 4134 3275 4138
rect 3311 4134 3315 4138
rect 1787 4110 1791 4114
rect 1935 4110 1939 4114
rect 1679 3998 1683 4002
rect 1815 3998 1819 4002
rect 1935 3998 1939 4002
rect 1371 3886 1375 3890
rect 1499 3886 1503 3890
rect 1587 3886 1591 3890
rect 1787 3886 1791 3890
rect 3839 4206 3843 4210
rect 3971 4206 3975 4210
rect 4107 4206 4111 4210
rect 4059 4179 4063 4180
rect 4059 4176 4063 4179
rect 5663 4458 5667 4462
rect 4511 4330 4515 4334
rect 4543 4330 4547 4334
rect 4647 4330 4651 4334
rect 4679 4330 4683 4334
rect 4783 4330 4787 4334
rect 4919 4330 4923 4334
rect 5663 4330 5667 4334
rect 4243 4206 4247 4210
rect 4379 4206 4383 4210
rect 4515 4206 4519 4210
rect 4651 4206 4655 4210
rect 5663 4206 5667 4210
rect 3407 4134 3411 4138
rect 3543 4134 3547 4138
rect 3679 4134 3683 4138
rect 3799 4134 3803 4138
rect 3839 4070 3843 4074
rect 3887 4070 3891 4074
rect 3999 4070 4003 4074
rect 4023 4070 4027 4074
rect 4135 4070 4139 4074
rect 4159 4070 4163 4074
rect 4271 4070 4275 4074
rect 3839 3958 3843 3962
rect 3859 3958 3863 3962
rect 3995 3958 3999 3962
rect 1975 3930 1979 3934
rect 1995 3930 1999 3934
rect 2403 3930 2407 3934
rect 2827 3930 2831 3934
rect 3107 3930 3111 3934
rect 3243 3930 3247 3934
rect 3251 3930 3255 3934
rect 3379 3930 3383 3934
rect 3515 3930 3519 3934
rect 3651 3930 3655 3934
rect 1935 3886 1939 3890
rect 1975 3818 1979 3822
rect 2023 3818 2027 3822
rect 927 3762 931 3766
rect 1063 3762 1067 3766
rect 1223 3762 1227 3766
rect 1343 3762 1347 3766
rect 1527 3762 1531 3766
rect 1815 3762 1819 3766
rect 1935 3762 1939 3766
rect 635 3634 639 3638
rect 763 3634 767 3638
rect 779 3634 783 3638
rect 923 3634 927 3638
rect 1035 3634 1039 3638
rect 1067 3634 1071 3638
rect 111 3502 115 3506
rect 431 3502 435 3506
rect 519 3502 523 3506
rect 567 3502 571 3506
rect 663 3502 667 3506
rect 703 3502 707 3506
rect 807 3502 811 3506
rect 839 3502 843 3506
rect 111 3382 115 3386
rect 323 3382 327 3386
rect 403 3382 407 3386
rect 459 3382 463 3386
rect 539 3382 543 3386
rect 595 3382 599 3386
rect 675 3382 679 3386
rect 731 3382 735 3386
rect 811 3382 815 3386
rect 111 3262 115 3266
rect 159 3262 163 3266
rect 335 3262 339 3266
rect 351 3262 355 3266
rect 487 3262 491 3266
rect 543 3262 547 3266
rect 111 3134 115 3138
rect 131 3134 135 3138
rect 951 3502 955 3506
rect 975 3502 979 3506
rect 3799 3930 3803 3934
rect 4523 4176 4527 4180
rect 4295 4070 4299 4074
rect 4407 4070 4411 4074
rect 4431 4070 4435 4074
rect 4543 4070 4547 4074
rect 4567 4070 4571 4074
rect 4703 4070 4707 4074
rect 4839 4070 4843 4074
rect 5663 4070 5667 4074
rect 4131 3958 4135 3962
rect 4147 3958 4151 3962
rect 4267 3958 4271 3962
rect 4299 3958 4303 3962
rect 4403 3958 4407 3962
rect 4459 3958 4463 3962
rect 4539 3958 4543 3962
rect 4619 3958 4623 3962
rect 4675 3958 4679 3962
rect 4779 3958 4783 3962
rect 4811 3958 4815 3962
rect 5663 3958 5667 3962
rect 2175 3818 2179 3822
rect 2351 3818 2355 3822
rect 2431 3818 2435 3822
rect 2535 3818 2539 3822
rect 2719 3818 2723 3822
rect 2855 3818 2859 3822
rect 2895 3818 2899 3822
rect 3071 3818 3075 3822
rect 3247 3818 3251 3822
rect 3279 3818 3283 3822
rect 3423 3818 3427 3822
rect 3607 3818 3611 3822
rect 1975 3698 1979 3702
rect 1995 3698 1999 3702
rect 2011 3698 2015 3702
rect 2147 3698 2151 3702
rect 2291 3698 2295 3702
rect 2323 3698 2327 3702
rect 2435 3698 2439 3702
rect 2507 3698 2511 3702
rect 2579 3698 2583 3702
rect 2691 3698 2695 3702
rect 2723 3698 2727 3702
rect 2867 3698 2871 3702
rect 3011 3698 3015 3702
rect 3043 3698 3047 3702
rect 3155 3698 3159 3702
rect 3219 3698 3223 3702
rect 3299 3698 3303 3702
rect 3395 3698 3399 3702
rect 1211 3634 1215 3638
rect 1315 3634 1319 3638
rect 1935 3634 1939 3638
rect 1975 3578 1979 3582
rect 2039 3578 2043 3582
rect 2175 3578 2179 3582
rect 2239 3578 2243 3582
rect 2319 3578 2323 3582
rect 2375 3578 2379 3582
rect 2463 3578 2467 3582
rect 2511 3578 2515 3582
rect 1095 3502 1099 3506
rect 1239 3502 1243 3506
rect 1935 3502 1939 3506
rect 2607 3578 2611 3582
rect 2647 3578 2651 3582
rect 2751 3578 2755 3582
rect 2783 3578 2787 3582
rect 2895 3578 2899 3582
rect 2919 3578 2923 3582
rect 1975 3462 1979 3466
rect 2171 3462 2175 3466
rect 2211 3462 2215 3466
rect 2347 3462 2351 3466
rect 2483 3462 2487 3466
rect 2531 3462 2535 3466
rect 2619 3462 2623 3466
rect 2715 3462 2719 3466
rect 2755 3462 2759 3466
rect 3679 3818 3683 3822
rect 3799 3818 3803 3822
rect 3839 3818 3843 3822
rect 3887 3818 3891 3822
rect 4023 3818 4027 3822
rect 4175 3818 4179 3822
rect 4327 3818 4331 3822
rect 4487 3818 4491 3822
rect 4503 3818 4507 3822
rect 4639 3818 4643 3822
rect 4647 3818 4651 3822
rect 4775 3818 4779 3822
rect 3579 3698 3583 3702
rect 3799 3698 3803 3702
rect 3839 3686 3843 3690
rect 4019 3686 4023 3690
rect 4807 3818 4811 3822
rect 4911 3818 4915 3822
rect 5047 3818 5051 3822
rect 5663 3818 5667 3822
rect 4155 3686 4159 3690
rect 4291 3686 4295 3690
rect 4427 3686 4431 3690
rect 4475 3686 4479 3690
rect 4563 3686 4567 3690
rect 4611 3686 4615 3690
rect 4699 3686 4703 3690
rect 4747 3686 4751 3690
rect 4835 3686 4839 3690
rect 4883 3686 4887 3690
rect 4971 3686 4975 3690
rect 5019 3686 5023 3690
rect 5107 3686 5111 3690
rect 5243 3686 5247 3690
rect 5379 3686 5383 3690
rect 5515 3686 5519 3690
rect 5663 3686 5667 3690
rect 3039 3578 3043 3582
rect 3055 3578 3059 3582
rect 3183 3578 3187 3582
rect 3191 3578 3195 3582
rect 3327 3578 3331 3582
rect 3463 3578 3467 3582
rect 3799 3578 3803 3582
rect 2891 3462 2895 3466
rect 2907 3462 2911 3466
rect 3027 3462 3031 3466
rect 3099 3462 3103 3466
rect 3163 3462 3167 3466
rect 3291 3462 3295 3466
rect 3299 3462 3303 3466
rect 867 3382 871 3386
rect 947 3382 951 3386
rect 1935 3382 1939 3386
rect 623 3262 627 3266
rect 1975 3326 1979 3330
rect 2151 3326 2155 3330
rect 2199 3326 2203 3330
rect 2375 3326 2379 3330
rect 2399 3326 2403 3330
rect 2559 3326 2563 3330
rect 2687 3326 2691 3330
rect 2743 3326 2747 3330
rect 2935 3326 2939 3330
rect 3015 3326 3019 3330
rect 751 3262 755 3266
rect 759 3262 763 3266
rect 895 3262 899 3266
rect 959 3262 963 3266
rect 1935 3262 1939 3266
rect 307 3134 311 3138
rect 371 3134 375 3138
rect 515 3134 519 3138
rect 627 3134 631 3138
rect 723 3134 727 3138
rect 875 3134 879 3138
rect 931 3134 935 3138
rect 111 3022 115 3026
rect 159 3022 163 3026
rect 175 3022 179 3026
rect 399 3022 403 3026
rect 407 3022 411 3026
rect 623 3022 627 3026
rect 655 3022 659 3026
rect 111 2906 115 2910
rect 147 2906 151 2910
rect 379 2906 383 2910
rect 395 2906 399 2910
rect 1115 3134 1119 3138
rect 1347 3134 1351 3138
rect 1579 3134 1583 3138
rect 1787 3134 1791 3138
rect 823 3022 827 3026
rect 903 3022 907 3026
rect 1007 3022 1011 3026
rect 1143 3022 1147 3026
rect 1183 3022 1187 3026
rect 1351 3022 1355 3026
rect 1375 3022 1379 3026
rect 1975 3214 1979 3218
rect 1995 3214 1999 3218
rect 2123 3214 2127 3218
rect 2147 3214 2151 3218
rect 2347 3214 2351 3218
rect 2371 3214 2375 3218
rect 2555 3214 2559 3218
rect 2659 3214 2663 3218
rect 3839 3526 3843 3530
rect 4047 3526 4051 3530
rect 4183 3526 4187 3530
rect 4319 3526 4323 3530
rect 4455 3526 4459 3530
rect 4591 3526 4595 3530
rect 4727 3526 4731 3530
rect 4863 3526 4867 3530
rect 4999 3526 5003 3530
rect 5135 3526 5139 3530
rect 5271 3526 5275 3530
rect 5407 3526 5411 3530
rect 5543 3526 5547 3530
rect 3435 3462 3439 3466
rect 3483 3462 3487 3466
rect 3651 3462 3655 3466
rect 3799 3462 3803 3466
rect 5663 3526 5667 3530
rect 3839 3406 3843 3410
rect 3859 3406 3863 3410
rect 4099 3406 4103 3410
rect 4347 3406 4351 3410
rect 4587 3406 4591 3410
rect 4811 3406 4815 3410
rect 5027 3406 5031 3410
rect 5235 3406 5239 3410
rect 5379 3406 5383 3410
rect 5451 3406 5455 3410
rect 5515 3406 5519 3410
rect 3127 3326 3131 3330
rect 3319 3326 3323 3330
rect 3359 3326 3363 3330
rect 3511 3326 3515 3330
rect 3679 3326 3683 3330
rect 3799 3326 3803 3330
rect 3839 3294 3843 3298
rect 3887 3294 3891 3298
rect 4127 3294 4131 3298
rect 2771 3214 2775 3218
rect 2987 3214 2991 3218
rect 3211 3214 3215 3218
rect 3331 3214 3335 3218
rect 3443 3214 3447 3218
rect 3651 3214 3655 3218
rect 1935 3134 1939 3138
rect 1975 3102 1979 3106
rect 2023 3102 2027 3106
rect 2175 3102 2179 3106
rect 2375 3102 2379 3106
rect 2583 3102 2587 3106
rect 2647 3102 2651 3106
rect 2783 3102 2787 3106
rect 2799 3102 2803 3106
rect 1511 3022 1515 3026
rect 1607 3022 1611 3026
rect 1671 3022 1675 3026
rect 1815 3022 1819 3026
rect 1935 3022 1939 3026
rect 595 2906 599 2910
rect 787 2906 791 2910
rect 795 2906 799 2910
rect 111 2782 115 2786
rect 423 2782 427 2786
rect 623 2782 627 2786
rect 655 2782 659 2786
rect 1975 2990 1979 2994
rect 2619 2990 2623 2994
rect 2755 2990 2759 2994
rect 2803 2990 2807 2994
rect 2927 3102 2931 3106
rect 3015 3102 3019 3106
rect 3079 3102 3083 3106
rect 3239 3102 3243 3106
rect 3799 3214 3803 3218
rect 4375 3294 4379 3298
rect 4607 3294 4611 3298
rect 4615 3294 4619 3298
rect 3839 3166 3843 3170
rect 3859 3166 3863 3170
rect 4099 3166 4103 3170
rect 4347 3166 4351 3170
rect 4467 3166 4471 3170
rect 4579 3166 4583 3170
rect 4651 3166 4655 3170
rect 3399 3102 3403 3106
rect 3471 3102 3475 3106
rect 3567 3102 3571 3106
rect 3679 3102 3683 3106
rect 3799 3102 3803 3106
rect 4815 3294 4819 3298
rect 4839 3294 4843 3298
rect 5015 3294 5019 3298
rect 5055 3294 5059 3298
rect 5199 3294 5203 3298
rect 5263 3294 5267 3298
rect 5383 3294 5387 3298
rect 5479 3294 5483 3298
rect 5543 3294 5547 3298
rect 4787 3166 4791 3170
rect 4859 3166 4863 3170
rect 4987 3166 4991 3170
rect 5075 3166 5079 3170
rect 5171 3166 5175 3170
rect 5307 3166 5311 3170
rect 5355 3166 5359 3170
rect 2899 2990 2903 2994
rect 2939 2990 2943 2994
rect 3051 2990 3055 2994
rect 3075 2990 3079 2994
rect 3211 2990 3215 2994
rect 3347 2990 3351 2994
rect 3371 2990 3375 2994
rect 3483 2990 3487 2994
rect 3539 2990 3543 2994
rect 971 2906 975 2910
rect 979 2906 983 2910
rect 1147 2906 1151 2910
rect 1155 2906 1159 2910
rect 1315 2906 1319 2910
rect 1323 2906 1327 2910
rect 1483 2906 1487 2910
rect 1643 2906 1647 2910
rect 1787 2906 1791 2910
rect 1935 2906 1939 2910
rect 815 2782 819 2786
rect 975 2782 979 2786
rect 999 2782 1003 2786
rect 1143 2782 1147 2786
rect 1175 2782 1179 2786
rect 111 2670 115 2674
rect 627 2670 631 2674
rect 771 2670 775 2674
rect 787 2670 791 2674
rect 907 2670 911 2674
rect 947 2670 951 2674
rect 1311 2782 1315 2786
rect 1343 2782 1347 2786
rect 1479 2782 1483 2786
rect 1511 2782 1515 2786
rect 1671 2782 1675 2786
rect 1815 2782 1819 2786
rect 1975 2826 1979 2830
rect 2023 2826 2027 2830
rect 2167 2826 2171 2830
rect 2335 2826 2339 2830
rect 2495 2826 2499 2830
rect 2663 2826 2667 2830
rect 2831 2826 2835 2830
rect 2967 2826 2971 2830
rect 2999 2826 3003 2830
rect 1935 2782 1939 2786
rect 1043 2670 1047 2674
rect 1115 2670 1119 2674
rect 1179 2670 1183 2674
rect 1283 2670 1287 2674
rect 1315 2670 1319 2674
rect 1451 2670 1455 2674
rect 111 2542 115 2546
rect 551 2542 555 2546
rect 687 2542 691 2546
rect 799 2542 803 2546
rect 831 2542 835 2546
rect 935 2542 939 2546
rect 983 2542 987 2546
rect 1071 2542 1075 2546
rect 1135 2542 1139 2546
rect 1207 2542 1211 2546
rect 1295 2542 1299 2546
rect 1343 2542 1347 2546
rect 111 2418 115 2422
rect 131 2418 135 2422
rect 339 2418 343 2422
rect 523 2418 527 2422
rect 563 2418 567 2422
rect 659 2418 663 2422
rect 111 2302 115 2306
rect 159 2302 163 2306
rect 1975 2714 1979 2718
rect 1995 2714 1999 2718
rect 2139 2714 2143 2718
rect 2307 2714 2311 2718
rect 2379 2714 2383 2718
rect 2467 2714 2471 2718
rect 1587 2670 1591 2674
rect 1723 2670 1727 2674
rect 1935 2670 1939 2674
rect 1455 2542 1459 2546
rect 1479 2542 1483 2546
rect 1615 2542 1619 2546
rect 1751 2542 1755 2546
rect 1783 2542 1787 2546
rect 803 2418 807 2422
rect 955 2418 959 2422
rect 1043 2418 1047 2422
rect 1107 2418 1111 2422
rect 1267 2418 1271 2422
rect 1291 2418 1295 2422
rect 2515 2714 2519 2718
rect 2635 2714 2639 2718
rect 2659 2714 2663 2718
rect 1975 2598 1979 2602
rect 2407 2598 2411 2602
rect 2511 2598 2515 2602
rect 2543 2598 2547 2602
rect 1935 2542 1939 2546
rect 3839 3054 3843 3058
rect 4255 3054 4259 3058
rect 4455 3054 4459 3058
rect 4495 3054 4499 3058
rect 3799 2990 3803 2994
rect 3839 2918 3843 2922
rect 3995 2918 3999 2922
rect 4211 2918 4215 2922
rect 4227 2918 4231 2922
rect 4427 2918 4431 2922
rect 4443 2918 4447 2922
rect 3103 2826 3107 2830
rect 3167 2826 3171 2830
rect 3239 2826 3243 2830
rect 3375 2826 3379 2830
rect 3511 2826 3515 2830
rect 3799 2826 3803 2830
rect 3839 2802 3843 2806
rect 3919 2802 3923 2806
rect 2803 2714 2807 2718
rect 2947 2714 2951 2718
rect 2971 2714 2975 2718
rect 3091 2714 3095 2718
rect 3139 2714 3143 2718
rect 3235 2714 3239 2718
rect 3799 2714 3803 2718
rect 2647 2598 2651 2602
rect 2687 2598 2691 2602
rect 2783 2598 2787 2602
rect 2831 2598 2835 2602
rect 2919 2598 2923 2602
rect 2975 2598 2979 2602
rect 3055 2598 3059 2602
rect 3119 2598 3123 2602
rect 3191 2598 3195 2602
rect 3263 2598 3267 2602
rect 1975 2470 1979 2474
rect 2307 2470 2311 2474
rect 2483 2470 2487 2474
rect 2515 2470 2519 2474
rect 2619 2470 2623 2474
rect 2715 2470 2719 2474
rect 2755 2470 2759 2474
rect 1427 2418 1431 2422
rect 1547 2418 1551 2422
rect 1587 2418 1591 2422
rect 1755 2418 1759 2422
rect 1787 2418 1791 2422
rect 1935 2418 1939 2422
rect 319 2302 323 2306
rect 367 2302 371 2306
rect 551 2302 555 2306
rect 591 2302 595 2306
rect 831 2302 835 2306
rect 1071 2302 1075 2306
rect 1151 2302 1155 2306
rect 1319 2302 1323 2306
rect 1495 2302 1499 2306
rect 1575 2302 1579 2306
rect 1815 2302 1819 2306
rect 111 2166 115 2170
rect 131 2166 135 2170
rect 291 2166 295 2170
rect 483 2166 487 2170
rect 523 2166 527 2170
rect 691 2166 695 2170
rect 803 2166 807 2170
rect 915 2166 919 2170
rect 1123 2166 1127 2170
rect 1147 2166 1151 2170
rect 111 2050 115 2054
rect 263 2050 267 2054
rect 319 2050 323 2054
rect 399 2050 403 2054
rect 511 2050 515 2054
rect 535 2050 539 2054
rect 679 2050 683 2054
rect 719 2050 723 2054
rect 823 2050 827 2054
rect 943 2050 947 2054
rect 967 2050 971 2054
rect 111 1926 115 1930
rect 235 1926 239 1930
rect 371 1926 375 1930
rect 435 1926 439 1930
rect 507 1926 511 1930
rect 627 1926 631 1930
rect 651 1926 655 1930
rect 111 1802 115 1806
rect 223 1802 227 1806
rect 263 1802 267 1806
rect 795 1926 799 1930
rect 811 1926 815 1930
rect 1975 2350 1979 2354
rect 2223 2350 2227 2354
rect 1935 2302 1939 2306
rect 2891 2470 2895 2474
rect 2907 2470 2911 2474
rect 4671 3054 4675 3058
rect 4679 3054 4683 3058
rect 4887 3054 4891 3058
rect 4911 3054 4915 3058
rect 5103 3054 5107 3058
rect 5167 3054 5171 3058
rect 5335 3054 5339 3058
rect 5663 3406 5667 3410
rect 5663 3294 5667 3298
rect 5515 3166 5519 3170
rect 5663 3166 5667 3170
rect 5423 3054 5427 3058
rect 5543 3054 5547 3058
rect 4643 2918 4647 2922
rect 4699 2918 4703 2922
rect 4883 2918 4887 2922
rect 4971 2918 4975 2922
rect 5139 2918 5143 2922
rect 5251 2918 5255 2922
rect 5395 2918 5399 2922
rect 4023 2802 4027 2806
rect 4055 2802 4059 2806
rect 4191 2802 4195 2806
rect 4239 2802 4243 2806
rect 4327 2802 4331 2806
rect 4463 2802 4467 2806
rect 4471 2802 4475 2806
rect 4727 2802 4731 2806
rect 4999 2802 5003 2806
rect 5279 2802 5283 2806
rect 3839 2678 3843 2682
rect 3891 2678 3895 2682
rect 4027 2678 4031 2682
rect 4099 2678 4103 2682
rect 4163 2678 4167 2682
rect 4299 2678 4303 2682
rect 4435 2678 4439 2682
rect 4515 2678 4519 2682
rect 4755 2678 4759 2682
rect 5011 2678 5015 2682
rect 5275 2678 5279 2682
rect 3327 2598 3331 2602
rect 3463 2598 3467 2602
rect 3799 2598 3803 2602
rect 3839 2562 3843 2566
rect 4127 2562 4131 2566
rect 4327 2562 4331 2566
rect 4495 2562 4499 2566
rect 4543 2562 4547 2566
rect 4631 2562 4635 2566
rect 4767 2562 4771 2566
rect 4783 2562 4787 2566
rect 4903 2562 4907 2566
rect 3027 2470 3031 2474
rect 3099 2470 3103 2474
rect 3163 2470 3167 2474
rect 3283 2470 3287 2474
rect 3299 2470 3303 2474
rect 3435 2470 3439 2474
rect 3467 2470 3471 2474
rect 3651 2470 3655 2474
rect 3799 2470 3803 2474
rect 2335 2350 2339 2354
rect 2503 2350 2507 2354
rect 2543 2350 2547 2354
rect 2743 2350 2747 2354
rect 2767 2350 2771 2354
rect 2935 2350 2939 2354
rect 3007 2350 3011 2354
rect 3127 2350 3131 2354
rect 3239 2350 3243 2354
rect 3311 2350 3315 2354
rect 3471 2350 3475 2354
rect 3495 2350 3499 2354
rect 3679 2350 3683 2354
rect 1975 2238 1979 2242
rect 1995 2238 1999 2242
rect 2155 2238 2159 2242
rect 2195 2238 2199 2242
rect 2387 2238 2391 2242
rect 2475 2238 2479 2242
rect 3839 2434 3843 2438
rect 4467 2434 4471 2438
rect 4603 2434 4607 2438
rect 4699 2434 4703 2438
rect 4739 2434 4743 2438
rect 5515 2918 5519 2922
rect 5663 3054 5667 3058
rect 5663 2918 5667 2922
rect 5543 2802 5547 2806
rect 5515 2678 5519 2682
rect 5039 2562 5043 2566
rect 5303 2562 5307 2566
rect 4835 2434 4839 2438
rect 4875 2434 4879 2438
rect 4971 2434 4975 2438
rect 5011 2434 5015 2438
rect 5107 2434 5111 2438
rect 5243 2434 5247 2438
rect 5379 2434 5383 2438
rect 3799 2350 3803 2354
rect 3839 2310 3843 2314
rect 3887 2310 3891 2314
rect 4183 2310 4187 2314
rect 4495 2310 4499 2314
rect 4727 2310 4731 2314
rect 4791 2310 4795 2314
rect 4863 2310 4867 2314
rect 4999 2310 5003 2314
rect 5087 2310 5091 2314
rect 5135 2310 5139 2314
rect 5271 2310 5275 2314
rect 2667 2238 2671 2242
rect 2739 2238 2743 2242
rect 2979 2238 2983 2242
rect 2987 2238 2991 2242
rect 3211 2238 3215 2242
rect 3331 2238 3335 2242
rect 3443 2238 3447 2242
rect 3651 2238 3655 2242
rect 3799 2238 3803 2242
rect 3839 2194 3843 2198
rect 3859 2194 3863 2198
rect 1387 2166 1391 2170
rect 1467 2166 1471 2170
rect 1635 2166 1639 2170
rect 1787 2166 1791 2170
rect 1935 2166 1939 2170
rect 1111 2050 1115 2054
rect 1175 2050 1179 2054
rect 1255 2050 1259 2054
rect 1399 2050 1403 2054
rect 1415 2050 1419 2054
rect 1543 2050 1547 2054
rect 1663 2050 1667 2054
rect 1679 2050 1683 2054
rect 1815 2050 1819 2054
rect 1935 2050 1939 2054
rect 939 1926 943 1930
rect 987 1926 991 1930
rect 1083 1926 1087 1930
rect 1155 1926 1159 1930
rect 1227 1926 1231 1930
rect 1323 1926 1327 1930
rect 1371 1926 1375 1930
rect 1483 1926 1487 1930
rect 1515 1926 1519 1930
rect 1643 1926 1647 1930
rect 1651 1926 1655 1930
rect 463 1802 467 1806
rect 655 1802 659 1806
rect 695 1802 699 1806
rect 839 1802 843 1806
rect 927 1802 931 1806
rect 1015 1802 1019 1806
rect 1159 1802 1163 1806
rect 1183 1802 1187 1806
rect 1351 1802 1355 1806
rect 111 1678 115 1682
rect 131 1678 135 1682
rect 195 1678 199 1682
rect 363 1678 367 1682
rect 435 1678 439 1682
rect 111 1554 115 1558
rect 159 1554 163 1558
rect 619 1678 623 1682
rect 667 1678 671 1682
rect 875 1678 879 1682
rect 899 1678 903 1682
rect 1131 1678 1135 1682
rect 1139 1678 1143 1682
rect 327 1554 331 1558
rect 391 1554 395 1558
rect 511 1554 515 1558
rect 111 1430 115 1434
rect 131 1430 135 1434
rect 299 1430 303 1434
rect 111 1318 115 1322
rect 159 1318 163 1322
rect 3995 2194 3999 2198
rect 4131 2194 4135 2198
rect 4155 2194 4159 2198
rect 4267 2194 4271 2198
rect 4403 2194 4407 2198
rect 4467 2194 4471 2198
rect 4539 2194 4543 2198
rect 3839 2062 3843 2066
rect 3887 2062 3891 2066
rect 4023 2062 4027 2066
rect 4159 2062 4163 2066
rect 4295 2062 4299 2066
rect 4431 2062 4435 2066
rect 3839 1950 3843 1954
rect 3859 1950 3863 1954
rect 1787 1926 1791 1930
rect 1935 1926 1939 1930
rect 1975 1926 1979 1930
rect 2023 1926 2027 1930
rect 2183 1926 2187 1930
rect 2415 1926 2419 1930
rect 2695 1926 2699 1930
rect 3015 1926 3019 1930
rect 3135 1926 3139 1930
rect 3271 1926 3275 1930
rect 3359 1926 3363 1930
rect 3407 1926 3411 1930
rect 3543 1926 3547 1930
rect 3679 1926 3683 1930
rect 3799 1926 3803 1930
rect 1391 1802 1395 1806
rect 1511 1802 1515 1806
rect 1671 1802 1675 1806
rect 1815 1802 1819 1806
rect 1935 1802 1939 1806
rect 1975 1802 1979 1806
rect 1995 1802 1999 1806
rect 2131 1802 2135 1806
rect 2267 1802 2271 1806
rect 2419 1802 2423 1806
rect 2579 1802 2583 1806
rect 2739 1802 2743 1806
rect 2899 1802 2903 1806
rect 3051 1802 3055 1806
rect 3107 1802 3111 1806
rect 3203 1802 3207 1806
rect 3243 1802 3247 1806
rect 1363 1678 1367 1682
rect 1935 1678 1939 1682
rect 1975 1678 1979 1682
rect 2023 1678 2027 1682
rect 2159 1678 2163 1682
rect 2167 1678 2171 1682
rect 2295 1678 2299 1682
rect 2319 1678 2323 1682
rect 2447 1678 2451 1682
rect 2479 1678 2483 1682
rect 2607 1678 2611 1682
rect 2639 1678 2643 1682
rect 647 1554 651 1558
rect 695 1554 699 1558
rect 887 1554 891 1558
rect 903 1554 907 1558
rect 1079 1554 1083 1558
rect 1167 1554 1171 1558
rect 1935 1554 1939 1558
rect 1975 1554 1979 1558
rect 1995 1554 1999 1558
rect 395 1430 399 1434
rect 483 1430 487 1434
rect 667 1430 671 1434
rect 683 1430 687 1434
rect 3023 1784 3027 1788
rect 5663 2802 5667 2806
rect 5663 2678 5667 2682
rect 5543 2562 5547 2566
rect 5515 2434 5519 2438
rect 5663 2562 5667 2566
rect 5663 2434 5667 2438
rect 5383 2310 5387 2314
rect 5407 2310 5411 2314
rect 5543 2310 5547 2314
rect 4699 2194 4703 2198
rect 4763 2194 4767 2198
rect 4891 2194 4895 2198
rect 5059 2194 5063 2198
rect 5099 2194 5103 2198
rect 5315 2194 5319 2198
rect 5355 2194 5359 2198
rect 5515 2194 5519 2198
rect 4567 2062 4571 2066
rect 4719 2062 4723 2066
rect 4727 2062 4731 2066
rect 4895 2062 4899 2066
rect 4919 2062 4923 2066
rect 5087 2062 5091 2066
rect 5127 2062 5131 2066
rect 5279 2062 5283 2066
rect 5343 2062 5347 2066
rect 5479 2062 5483 2066
rect 5543 2062 5547 2066
rect 5663 2310 5667 2314
rect 5663 2194 5667 2198
rect 3995 1950 3999 1954
rect 4043 1950 4047 1954
rect 4131 1950 4135 1954
rect 4267 1950 4271 1954
rect 4283 1950 4287 1954
rect 4403 1950 4407 1954
rect 4539 1950 4543 1954
rect 4563 1950 4567 1954
rect 4691 1950 4695 1954
rect 4867 1950 4871 1954
rect 4875 1950 4879 1954
rect 5059 1950 5063 1954
rect 5203 1950 5207 1954
rect 5251 1950 5255 1954
rect 5451 1950 5455 1954
rect 3839 1838 3843 1842
rect 3887 1838 3891 1842
rect 4071 1838 4075 1842
rect 4311 1838 4315 1842
rect 4407 1838 4411 1842
rect 3355 1802 3359 1806
rect 3379 1802 3383 1806
rect 3515 1802 3519 1806
rect 3651 1802 3655 1806
rect 3799 1802 3803 1806
rect 2767 1678 2771 1682
rect 2791 1678 2795 1682
rect 2927 1678 2931 1682
rect 2943 1678 2947 1682
rect 3079 1678 3083 1682
rect 3103 1678 3107 1682
rect 3231 1678 3235 1682
rect 3263 1678 3267 1682
rect 3771 1784 3775 1788
rect 4543 1838 4547 1842
rect 4591 1838 4595 1842
rect 4679 1838 4683 1842
rect 4815 1838 4819 1842
rect 4903 1838 4907 1842
rect 4951 1838 4955 1842
rect 5231 1838 5235 1842
rect 3839 1710 3843 1714
rect 4379 1710 4383 1714
rect 4515 1710 4519 1714
rect 4563 1710 4567 1714
rect 4651 1710 4655 1714
rect 4699 1710 4703 1714
rect 4787 1710 4791 1714
rect 4835 1710 4839 1714
rect 4923 1710 4927 1714
rect 3383 1678 3387 1682
rect 3423 1678 3427 1682
rect 3543 1678 3547 1682
rect 3679 1678 3683 1682
rect 3799 1678 3803 1682
rect 3839 1582 3843 1586
rect 4591 1582 4595 1586
rect 2131 1554 2135 1558
rect 2139 1554 2143 1558
rect 2267 1554 2271 1558
rect 2291 1554 2295 1558
rect 2403 1554 2407 1558
rect 2451 1554 2455 1558
rect 2539 1554 2543 1558
rect 2611 1554 2615 1558
rect 2675 1554 2679 1558
rect 2763 1554 2767 1558
rect 2811 1554 2815 1558
rect 2915 1554 2919 1558
rect 2947 1554 2951 1558
rect 3075 1554 3079 1558
rect 3083 1554 3087 1558
rect 3219 1554 3223 1558
rect 3235 1554 3239 1558
rect 3355 1554 3359 1558
rect 3395 1554 3399 1558
rect 3491 1554 3495 1558
rect 3799 1554 3803 1558
rect 859 1430 863 1434
rect 971 1430 975 1434
rect 1051 1430 1055 1434
rect 1259 1430 1263 1434
rect 1935 1430 1939 1434
rect 1975 1430 1979 1434
rect 2023 1430 2027 1434
rect 2159 1430 2163 1434
rect 2167 1430 2171 1434
rect 423 1318 427 1322
rect 455 1318 459 1322
rect 711 1318 715 1322
rect 775 1318 779 1322
rect 999 1318 1003 1322
rect 1095 1318 1099 1322
rect 1287 1318 1291 1322
rect 111 1182 115 1186
rect 131 1182 135 1186
rect 331 1182 335 1186
rect 427 1182 431 1186
rect 111 1070 115 1074
rect 159 1070 163 1074
rect 263 1070 267 1074
rect 2295 1430 2299 1434
rect 2303 1430 2307 1434
rect 2431 1430 2435 1434
rect 2439 1430 2443 1434
rect 2567 1430 2571 1434
rect 2575 1430 2579 1434
rect 1423 1318 1427 1322
rect 1935 1318 1939 1322
rect 1975 1318 1979 1322
rect 2131 1318 2135 1322
rect 2139 1318 2143 1322
rect 2267 1318 2271 1322
rect 2275 1318 2279 1322
rect 2403 1318 2407 1322
rect 2411 1318 2415 1322
rect 2703 1430 2707 1434
rect 2711 1430 2715 1434
rect 2839 1430 2843 1434
rect 2847 1430 2851 1434
rect 2975 1430 2979 1434
rect 2983 1430 2987 1434
rect 3111 1430 3115 1434
rect 3119 1430 3123 1434
rect 3247 1430 3251 1434
rect 3255 1430 3259 1434
rect 3383 1430 3387 1434
rect 3519 1430 3523 1434
rect 3799 1430 3803 1434
rect 4971 1710 4975 1714
rect 5107 1710 5111 1714
rect 5243 1710 5247 1714
rect 5379 1710 5383 1714
rect 4727 1582 4731 1586
rect 4863 1582 4867 1586
rect 4999 1582 5003 1586
rect 5135 1582 5139 1586
rect 5271 1582 5275 1586
rect 5515 1950 5519 1954
rect 5663 2062 5667 2066
rect 5663 1950 5667 1954
rect 5543 1838 5547 1842
rect 5515 1710 5519 1714
rect 5663 1838 5667 1842
rect 5663 1710 5667 1714
rect 5407 1582 5411 1586
rect 5543 1582 5547 1586
rect 5663 1582 5667 1586
rect 3839 1398 3843 1402
rect 4563 1398 4567 1402
rect 4699 1398 4703 1402
rect 4811 1398 4815 1402
rect 4835 1398 4839 1402
rect 4947 1398 4951 1402
rect 4971 1398 4975 1402
rect 5083 1398 5087 1402
rect 5107 1398 5111 1402
rect 5219 1398 5223 1402
rect 5243 1398 5247 1402
rect 5355 1398 5359 1402
rect 5379 1398 5383 1402
rect 5491 1398 5495 1402
rect 5515 1398 5519 1402
rect 5663 1398 5667 1402
rect 2547 1318 2551 1322
rect 2555 1318 2559 1322
rect 2683 1318 2687 1322
rect 2715 1318 2719 1322
rect 2819 1318 2823 1322
rect 2891 1318 2895 1322
rect 2955 1318 2959 1322
rect 3075 1318 3079 1322
rect 3091 1318 3095 1322
rect 3227 1318 3231 1322
rect 3267 1318 3271 1322
rect 2499 1296 2503 1300
rect 2723 1296 2727 1300
rect 1975 1206 1979 1210
rect 2023 1206 2027 1210
rect 2159 1206 2163 1210
rect 2239 1206 2243 1210
rect 2295 1206 2299 1210
rect 2431 1206 2435 1210
rect 2479 1206 2483 1210
rect 2583 1206 2587 1210
rect 2719 1206 2723 1210
rect 2743 1206 2747 1210
rect 563 1182 567 1186
rect 747 1182 751 1186
rect 803 1182 807 1186
rect 1043 1182 1047 1186
rect 1067 1182 1071 1186
rect 1283 1182 1287 1186
rect 1395 1182 1399 1186
rect 1523 1182 1527 1186
rect 1771 1182 1775 1186
rect 1935 1182 1939 1186
rect 2919 1206 2923 1210
rect 2959 1206 2963 1210
rect 359 1070 363 1074
rect 439 1070 443 1074
rect 591 1070 595 1074
rect 615 1070 619 1074
rect 783 1070 787 1074
rect 831 1070 835 1074
rect 111 954 115 958
rect 227 954 231 958
rect 235 954 239 958
rect 379 954 383 958
rect 411 954 415 958
rect 111 826 115 830
rect 255 826 259 830
rect 539 954 543 958
rect 587 954 591 958
rect 951 1070 955 1074
rect 1071 1070 1075 1074
rect 1111 1070 1115 1074
rect 1271 1070 1275 1074
rect 1311 1070 1315 1074
rect 1431 1070 1435 1074
rect 1551 1070 1555 1074
rect 1591 1070 1595 1074
rect 1751 1070 1755 1074
rect 3467 1318 3471 1322
rect 3651 1318 3655 1322
rect 3799 1318 3803 1322
rect 3103 1206 3107 1210
rect 3207 1206 3211 1210
rect 3295 1206 3299 1210
rect 3455 1206 3459 1210
rect 3495 1206 3499 1210
rect 1799 1070 1803 1074
rect 1935 1070 1939 1074
rect 1975 1070 1979 1074
rect 1995 1070 1999 1074
rect 2211 1070 2215 1074
rect 2451 1070 2455 1074
rect 2691 1070 2695 1074
rect 2931 1070 2935 1074
rect 3091 1070 3095 1074
rect 3179 1070 3183 1074
rect 3243 1070 3247 1074
rect 715 954 719 958
rect 755 954 759 958
rect 891 954 895 958
rect 923 954 927 958
rect 1075 954 1079 958
rect 1083 954 1087 958
rect 1243 954 1247 958
rect 1259 954 1263 958
rect 1403 954 1407 958
rect 1443 954 1447 958
rect 1563 954 1567 958
rect 1627 954 1631 958
rect 1723 954 1727 958
rect 1787 954 1791 958
rect 1935 954 1939 958
rect 375 826 379 830
rect 407 826 411 830
rect 567 826 571 830
rect 655 826 659 830
rect 743 826 747 830
rect 919 826 923 830
rect 943 826 947 830
rect 1103 826 1107 830
rect 111 714 115 718
rect 131 714 135 718
rect 307 714 311 718
rect 347 714 351 718
rect 499 714 503 718
rect 627 714 631 718
rect 683 714 687 718
rect 859 714 863 718
rect 915 714 919 718
rect 111 602 115 606
rect 159 602 163 606
rect 335 602 339 606
rect 375 602 379 606
rect 111 490 115 494
rect 131 490 135 494
rect 1975 930 1979 934
rect 2047 930 2051 934
rect 2351 930 2355 934
rect 2647 930 2651 934
rect 2927 930 2931 934
rect 1239 826 1243 830
rect 1287 826 1291 830
rect 1471 826 1475 830
rect 1535 826 1539 830
rect 1655 826 1659 830
rect 1815 826 1819 830
rect 1935 826 1939 830
rect 1975 818 1979 822
rect 1995 818 1999 822
rect 2019 818 2023 822
rect 2251 818 2255 822
rect 2323 818 2327 822
rect 1027 714 1031 718
rect 1187 714 1191 718
rect 1211 714 1215 718
rect 1339 714 1343 718
rect 1491 714 1495 718
rect 1507 714 1511 718
rect 1651 714 1655 718
rect 1787 714 1791 718
rect 527 602 531 606
rect 599 602 603 606
rect 711 602 715 606
rect 807 602 811 606
rect 887 602 891 606
rect 347 490 351 494
rect 427 490 431 494
rect 571 490 575 494
rect 999 602 1003 606
rect 1055 602 1059 606
rect 1175 602 1179 606
rect 1215 602 1219 606
rect 2523 818 2527 822
rect 2619 818 2623 822
rect 3119 930 3123 934
rect 3207 930 3211 934
rect 3271 930 3275 934
rect 3679 1206 3683 1210
rect 3839 1282 3843 1286
rect 4735 1282 4739 1286
rect 4839 1282 4843 1286
rect 4879 1282 4883 1286
rect 3799 1206 3803 1210
rect 4975 1282 4979 1286
rect 5031 1282 5035 1286
rect 5111 1282 5115 1286
rect 5191 1282 5195 1286
rect 5247 1282 5251 1286
rect 3839 1162 3843 1166
rect 3859 1162 3863 1166
rect 4067 1162 4071 1166
rect 4299 1162 4303 1166
rect 4539 1162 4543 1166
rect 4707 1162 4711 1166
rect 4779 1162 4783 1166
rect 4851 1162 4855 1166
rect 3395 1070 3399 1074
rect 3427 1070 3431 1074
rect 3651 1070 3655 1074
rect 3799 1070 3803 1074
rect 3839 1050 3843 1054
rect 3887 1050 3891 1054
rect 4071 1050 4075 1054
rect 4095 1050 4099 1054
rect 3839 938 3843 942
rect 3859 938 3863 942
rect 3423 930 3427 934
rect 3495 930 3499 934
rect 3799 930 3803 934
rect 2771 818 2775 822
rect 2899 818 2903 822
rect 3003 818 3007 822
rect 3179 818 3183 822
rect 3227 818 3231 822
rect 3451 818 3455 822
rect 3467 818 3471 822
rect 1935 714 1939 718
rect 1343 602 1347 606
rect 1367 602 1371 606
rect 1511 602 1515 606
rect 1519 602 1523 606
rect 1671 602 1675 606
rect 1679 602 1683 606
rect 1815 602 1819 606
rect 1935 602 1939 606
rect 1975 574 1979 578
rect 2023 574 2027 578
rect 2279 574 2283 578
rect 2551 574 2555 578
rect 2799 574 2803 578
rect 3031 574 3035 578
rect 3255 574 3259 578
rect 763 490 767 494
rect 779 490 783 494
rect 971 490 975 494
rect 1107 490 1111 494
rect 1147 490 1151 494
rect 1315 490 1319 494
rect 1459 490 1463 494
rect 1483 490 1487 494
rect 1643 490 1647 494
rect 1787 490 1791 494
rect 111 362 115 366
rect 159 362 163 366
rect 239 362 243 366
rect 391 362 395 366
rect 455 362 459 366
rect 551 362 555 366
rect 111 218 115 222
rect 147 218 151 222
rect 211 218 215 222
rect 711 362 715 366
rect 791 362 795 366
rect 871 362 875 366
rect 1031 362 1035 366
rect 1135 362 1139 366
rect 1487 362 1491 366
rect 283 218 287 222
rect 363 218 367 222
rect 419 218 423 222
rect 523 218 527 222
rect 555 218 559 222
rect 683 218 687 222
rect 691 218 695 222
rect 1935 490 1939 494
rect 4279 1050 4283 1054
rect 4327 1050 4331 1054
rect 4511 1050 4515 1054
rect 4567 1050 4571 1054
rect 3971 938 3975 942
rect 4043 938 4047 942
rect 4179 938 4183 942
rect 4251 938 4255 942
rect 4403 938 4407 942
rect 4483 938 4487 942
rect 3839 826 3843 830
rect 3887 826 3891 830
rect 3999 826 4003 830
rect 4047 826 4051 830
rect 4207 826 4211 830
rect 3651 818 3655 822
rect 3799 818 3803 822
rect 3839 706 3843 710
rect 3859 706 3863 710
rect 5359 1282 5363 1286
rect 5383 1282 5387 1286
rect 5519 1282 5523 1286
rect 5527 1282 5531 1286
rect 5003 1162 5007 1166
rect 5027 1162 5031 1166
rect 5163 1162 5167 1166
rect 5283 1162 5287 1166
rect 5331 1162 5335 1166
rect 4759 1050 4763 1054
rect 4807 1050 4811 1054
rect 5023 1050 5027 1054
rect 5055 1050 5059 1054
rect 5295 1050 5299 1054
rect 5311 1050 5315 1054
rect 5663 1282 5667 1286
rect 5499 1162 5503 1166
rect 5515 1162 5519 1166
rect 5663 1162 5667 1166
rect 5543 1050 5547 1054
rect 4643 938 4647 942
rect 4731 938 4735 942
rect 4899 938 4903 942
rect 4995 938 4999 942
rect 5171 938 5175 942
rect 5267 938 5271 942
rect 4279 826 4283 830
rect 4431 826 4435 830
rect 5663 1050 5667 1054
rect 5443 938 5447 942
rect 5515 938 5519 942
rect 4559 826 4563 830
rect 4671 826 4675 830
rect 4879 826 4883 830
rect 4927 826 4931 830
rect 5199 826 5203 830
rect 5223 826 5227 830
rect 5471 826 5475 830
rect 5543 826 5547 830
rect 5663 938 5667 942
rect 5663 826 5667 830
rect 3995 706 3999 710
rect 4019 706 4023 710
rect 4131 706 4135 710
rect 4251 706 4255 710
rect 4267 706 4271 710
rect 4403 706 4407 710
rect 4531 706 4535 710
rect 4571 706 4575 710
rect 4771 706 4775 710
rect 4851 706 4855 710
rect 4995 706 4999 710
rect 5195 706 5199 710
rect 5227 706 5231 710
rect 5459 706 5463 710
rect 5515 706 5519 710
rect 5663 706 5667 710
rect 3839 594 3843 598
rect 3887 594 3891 598
rect 3311 574 3315 578
rect 3447 574 3451 578
rect 3479 574 3483 578
rect 3583 574 3587 578
rect 3679 574 3683 578
rect 3799 574 3803 578
rect 1975 462 1979 466
rect 1995 462 1999 466
rect 2155 462 2159 466
rect 2347 462 2351 466
rect 2539 462 2543 466
rect 2731 462 2735 466
rect 2923 462 2927 466
rect 3115 462 3119 466
rect 3283 462 3287 466
rect 3299 462 3303 466
rect 3419 462 3423 466
rect 3483 462 3487 466
rect 3555 462 3559 466
rect 1815 362 1819 366
rect 1935 362 1939 366
rect 1975 326 1979 330
rect 2023 326 2027 330
rect 2047 326 2051 330
rect 2183 326 2187 330
rect 827 218 831 222
rect 843 218 847 222
rect 963 218 967 222
rect 1003 218 1007 222
rect 1099 218 1103 222
rect 1935 218 1939 222
rect 1975 198 1979 202
rect 1995 198 1999 202
rect 2019 198 2023 202
rect 2319 326 2323 330
rect 2375 326 2379 330
rect 2455 326 2459 330
rect 2567 326 2571 330
rect 2591 326 2595 330
rect 2727 326 2731 330
rect 2759 326 2763 330
rect 2863 326 2867 330
rect 2951 326 2955 330
rect 2999 326 3003 330
rect 3135 326 3139 330
rect 3143 326 3147 330
rect 3271 326 3275 330
rect 3327 326 3331 330
rect 3407 326 3411 330
rect 2131 198 2135 202
rect 2155 198 2159 202
rect 2267 198 2271 202
rect 2291 198 2295 202
rect 2403 198 2407 202
rect 2427 198 2431 202
rect 2539 198 2543 202
rect 2563 198 2567 202
rect 2675 198 2679 202
rect 2699 198 2703 202
rect 2811 198 2815 202
rect 2835 198 2839 202
rect 2947 198 2951 202
rect 2971 198 2975 202
rect 3083 198 3087 202
rect 3107 198 3111 202
rect 3219 198 3223 202
rect 4023 594 4027 598
rect 4159 594 4163 598
rect 4295 594 4299 598
rect 4431 594 4435 598
rect 4479 594 4483 598
rect 4599 594 4603 598
rect 4695 594 4699 598
rect 4799 594 4803 598
rect 4935 594 4939 598
rect 5023 594 5027 598
rect 5191 594 5195 598
rect 5255 594 5259 598
rect 5447 594 5451 598
rect 5487 594 5491 598
rect 3839 470 3843 474
rect 3859 470 3863 474
rect 3995 470 3999 474
rect 4131 470 4135 474
rect 4267 470 4271 474
rect 4451 470 4455 474
rect 3651 462 3655 466
rect 3799 462 3803 466
rect 4651 470 4655 474
rect 4667 470 4671 474
rect 4859 470 4863 474
rect 4907 470 4911 474
rect 5067 470 5071 474
rect 5163 470 5167 474
rect 5283 470 5287 474
rect 5419 470 5423 474
rect 3839 354 3843 358
rect 4479 354 4483 358
rect 4679 354 4683 358
rect 4751 354 4755 358
rect 4887 354 4891 358
rect 4911 354 4915 358
rect 3511 326 3515 330
rect 3543 326 3547 330
rect 3679 326 3683 330
rect 3799 326 3803 330
rect 5507 470 5511 474
rect 5663 594 5667 598
rect 5663 470 5667 474
rect 5071 354 5075 358
rect 5095 354 5099 358
rect 5231 354 5235 358
rect 5311 354 5315 358
rect 5399 354 5403 358
rect 5535 354 5539 358
rect 5543 354 5547 358
rect 3243 198 3247 202
rect 3355 198 3359 202
rect 3379 198 3383 202
rect 3491 198 3495 202
rect 3515 198 3519 202
rect 3627 198 3631 202
rect 3651 198 3655 202
rect 3799 198 3803 202
rect 3839 202 3843 206
rect 4291 202 4295 206
rect 4427 202 4431 206
rect 4563 202 4567 206
rect 4699 202 4703 206
rect 4723 202 4727 206
rect 4835 202 4839 206
rect 4883 202 4887 206
rect 4971 202 4975 206
rect 5043 202 5047 206
rect 5107 202 5111 206
rect 5203 202 5207 206
rect 5243 202 5247 206
rect 5371 202 5375 206
rect 5379 202 5383 206
rect 5663 354 5667 358
rect 5515 202 5519 206
rect 5663 202 5667 206
rect 111 106 115 110
rect 175 106 179 110
rect 311 106 315 110
rect 447 106 451 110
rect 583 106 587 110
rect 719 106 723 110
rect 855 106 859 110
rect 991 106 995 110
rect 1127 106 1131 110
rect 1935 106 1939 110
rect 1975 86 1979 90
rect 2023 86 2027 90
rect 2159 86 2163 90
rect 2295 86 2299 90
rect 2431 86 2435 90
rect 2567 86 2571 90
rect 2703 86 2707 90
rect 2839 86 2843 90
rect 2975 86 2979 90
rect 3111 86 3115 90
rect 3247 86 3251 90
rect 3383 86 3387 90
rect 3519 86 3523 90
rect 3655 86 3659 90
rect 3799 86 3803 90
rect 3839 90 3843 94
rect 4319 90 4323 94
rect 4455 90 4459 94
rect 4591 90 4595 94
rect 4727 90 4731 94
rect 4863 90 4867 94
rect 4999 90 5003 94
rect 5135 90 5139 94
rect 5271 90 5275 94
rect 5407 90 5411 94
rect 5543 90 5547 94
rect 5663 90 5667 94
<< m4 >>
rect 96 5753 97 5759
rect 103 5758 1959 5759
rect 103 5754 111 5758
rect 115 5754 131 5758
rect 135 5754 267 5758
rect 271 5754 403 5758
rect 407 5754 1935 5758
rect 1939 5754 1959 5758
rect 103 5753 1959 5754
rect 1965 5753 1966 5759
rect 3822 5694 5714 5695
rect 3822 5691 3839 5694
rect 1958 5685 1959 5691
rect 1965 5690 3823 5691
rect 1965 5686 1975 5690
rect 1979 5686 1995 5690
rect 1999 5686 2171 5690
rect 2175 5686 2371 5690
rect 2375 5686 2563 5690
rect 2567 5686 2747 5690
rect 2751 5686 2931 5690
rect 2935 5686 3107 5690
rect 3111 5686 3275 5690
rect 3279 5686 3443 5690
rect 3447 5686 3619 5690
rect 3623 5686 3799 5690
rect 3803 5686 3823 5690
rect 1965 5685 3823 5686
rect 3829 5690 3839 5691
rect 3843 5690 4467 5694
rect 4471 5690 4603 5694
rect 4607 5690 4739 5694
rect 4743 5690 4875 5694
rect 4879 5690 5663 5694
rect 5667 5690 5714 5694
rect 3829 5689 5714 5690
rect 3829 5685 3830 5689
rect 84 5641 85 5647
rect 91 5646 1947 5647
rect 91 5642 111 5646
rect 115 5642 159 5646
rect 163 5642 295 5646
rect 299 5642 343 5646
rect 347 5642 431 5646
rect 435 5642 535 5646
rect 539 5642 735 5646
rect 739 5642 943 5646
rect 947 5642 1159 5646
rect 1163 5642 1383 5646
rect 1387 5642 1607 5646
rect 1611 5642 1815 5646
rect 1819 5642 1935 5646
rect 1939 5642 1947 5646
rect 91 5641 1947 5642
rect 1953 5641 1954 5647
rect 3810 5582 5702 5583
rect 3810 5579 3839 5582
rect 1946 5573 1947 5579
rect 1953 5578 3811 5579
rect 1953 5574 1975 5578
rect 1979 5574 2023 5578
rect 2027 5574 2199 5578
rect 2203 5574 2375 5578
rect 2379 5574 2399 5578
rect 2403 5574 2591 5578
rect 2595 5574 2607 5578
rect 2611 5574 2775 5578
rect 2779 5574 2831 5578
rect 2835 5574 2959 5578
rect 2963 5574 3047 5578
rect 3051 5574 3135 5578
rect 3139 5574 3263 5578
rect 3267 5574 3303 5578
rect 3307 5574 3471 5578
rect 3475 5574 3479 5578
rect 3483 5574 3647 5578
rect 3651 5574 3679 5578
rect 3683 5574 3799 5578
rect 3803 5574 3811 5578
rect 1953 5573 3811 5574
rect 3817 5578 3839 5579
rect 3843 5578 4431 5582
rect 4435 5578 4495 5582
rect 4499 5578 4567 5582
rect 4571 5578 4631 5582
rect 4635 5578 4703 5582
rect 4707 5578 4767 5582
rect 4771 5578 4839 5582
rect 4843 5578 4903 5582
rect 4907 5578 4975 5582
rect 4979 5578 5111 5582
rect 5115 5578 5663 5582
rect 5667 5578 5702 5582
rect 3817 5577 5702 5578
rect 3817 5573 3818 5577
rect 96 5529 97 5535
rect 103 5534 1959 5535
rect 103 5530 111 5534
rect 115 5530 315 5534
rect 319 5530 507 5534
rect 511 5530 707 5534
rect 711 5530 875 5534
rect 879 5530 915 5534
rect 919 5530 1011 5534
rect 1015 5530 1131 5534
rect 1135 5530 1147 5534
rect 1151 5530 1291 5534
rect 1295 5530 1355 5534
rect 1359 5530 1435 5534
rect 1439 5530 1579 5534
rect 1583 5530 1723 5534
rect 1727 5530 1787 5534
rect 1791 5530 1935 5534
rect 1939 5530 1959 5534
rect 103 5529 1959 5530
rect 1965 5529 1966 5535
rect 3822 5465 3823 5471
rect 3829 5470 5707 5471
rect 3829 5466 3839 5470
rect 3843 5466 4403 5470
rect 4407 5466 4427 5470
rect 4431 5466 4539 5470
rect 4543 5466 4587 5470
rect 4591 5466 4675 5470
rect 4679 5466 4747 5470
rect 4751 5466 4811 5470
rect 4815 5466 4907 5470
rect 4911 5466 4947 5470
rect 4951 5466 5075 5470
rect 5079 5466 5083 5470
rect 5087 5466 5663 5470
rect 5667 5466 5707 5470
rect 3829 5465 5707 5466
rect 5713 5465 5714 5471
rect 3822 5463 3830 5465
rect 1958 5457 1959 5463
rect 1965 5462 3823 5463
rect 1965 5458 1975 5462
rect 1979 5458 2347 5462
rect 2351 5458 2451 5462
rect 2455 5458 2579 5462
rect 2583 5458 2699 5462
rect 2703 5458 2803 5462
rect 2807 5458 2947 5462
rect 2951 5458 3019 5462
rect 3023 5458 3187 5462
rect 3191 5458 3235 5462
rect 3239 5458 3427 5462
rect 3431 5458 3451 5462
rect 3455 5458 3651 5462
rect 3655 5458 3799 5462
rect 3803 5458 3823 5462
rect 1965 5457 3823 5458
rect 3829 5457 3830 5463
rect 84 5417 85 5423
rect 91 5422 1947 5423
rect 91 5418 111 5422
rect 115 5418 719 5422
rect 723 5418 855 5422
rect 859 5418 903 5422
rect 907 5418 991 5422
rect 995 5418 1039 5422
rect 1043 5418 1127 5422
rect 1131 5418 1175 5422
rect 1179 5418 1263 5422
rect 1267 5418 1319 5422
rect 1323 5418 1399 5422
rect 1403 5418 1463 5422
rect 1467 5418 1535 5422
rect 1539 5418 1607 5422
rect 1611 5418 1671 5422
rect 1675 5418 1751 5422
rect 1755 5418 1807 5422
rect 1811 5418 1935 5422
rect 1939 5418 1947 5422
rect 91 5417 1947 5418
rect 1953 5417 1954 5423
rect 1946 5345 1947 5351
rect 1953 5350 3811 5351
rect 1953 5346 1975 5350
rect 1979 5346 2319 5350
rect 2323 5346 2479 5350
rect 2483 5346 2519 5350
rect 2523 5346 2719 5350
rect 2723 5346 2727 5350
rect 2731 5346 2919 5350
rect 2923 5346 2975 5350
rect 2979 5346 3119 5350
rect 3123 5346 3215 5350
rect 3219 5346 3327 5350
rect 3331 5346 3455 5350
rect 3459 5346 3535 5350
rect 3539 5346 3679 5350
rect 3683 5346 3799 5350
rect 3803 5346 3811 5350
rect 1953 5345 3811 5346
rect 3817 5350 5702 5351
rect 3817 5346 3839 5350
rect 3843 5346 4431 5350
rect 4435 5346 4455 5350
rect 4459 5346 4615 5350
rect 4619 5346 4775 5350
rect 4779 5346 4799 5350
rect 4803 5346 4935 5350
rect 4939 5346 4983 5350
rect 4987 5346 5103 5350
rect 5107 5346 5175 5350
rect 5179 5346 5663 5350
rect 5667 5346 5702 5350
rect 3817 5345 5702 5346
rect 96 5305 97 5311
rect 103 5310 1959 5311
rect 103 5306 111 5310
rect 115 5306 691 5310
rect 695 5306 723 5310
rect 727 5306 827 5310
rect 831 5306 875 5310
rect 879 5306 963 5310
rect 967 5306 1027 5310
rect 1031 5306 1099 5310
rect 1103 5306 1187 5310
rect 1191 5306 1235 5310
rect 1239 5306 1355 5310
rect 1359 5306 1371 5310
rect 1375 5306 1507 5310
rect 1511 5306 1523 5310
rect 1527 5306 1643 5310
rect 1647 5306 1779 5310
rect 1783 5306 1935 5310
rect 1939 5306 1959 5310
rect 103 5305 1959 5306
rect 1965 5305 1966 5311
rect 1958 5229 1959 5235
rect 1965 5234 3823 5235
rect 1965 5230 1975 5234
rect 1979 5230 2275 5234
rect 2279 5230 2291 5234
rect 2295 5230 2475 5234
rect 2479 5230 2491 5234
rect 2495 5230 2683 5234
rect 2687 5230 2691 5234
rect 2695 5230 2891 5234
rect 2895 5230 3091 5234
rect 3095 5230 3099 5234
rect 3103 5230 3299 5234
rect 3303 5230 3307 5234
rect 3311 5230 3507 5234
rect 3511 5230 3799 5234
rect 3803 5230 3823 5234
rect 1965 5229 3823 5230
rect 3829 5229 3830 5235
rect 3822 5217 3823 5223
rect 3829 5222 5707 5223
rect 3829 5218 3839 5222
rect 3843 5218 4403 5222
rect 4407 5218 4435 5222
rect 4439 5218 4587 5222
rect 4591 5218 4595 5222
rect 4599 5218 4755 5222
rect 4759 5218 4771 5222
rect 4775 5218 4915 5222
rect 4919 5218 4955 5222
rect 4959 5218 5067 5222
rect 5071 5218 5147 5222
rect 5151 5218 5219 5222
rect 5223 5218 5379 5222
rect 5383 5218 5515 5222
rect 5519 5218 5663 5222
rect 5667 5218 5707 5222
rect 3829 5217 5707 5218
rect 5713 5217 5714 5223
rect 84 5193 85 5199
rect 91 5198 1947 5199
rect 91 5194 111 5198
rect 115 5194 447 5198
rect 451 5194 623 5198
rect 627 5194 751 5198
rect 755 5194 807 5198
rect 811 5194 903 5198
rect 907 5194 999 5198
rect 1003 5194 1055 5198
rect 1059 5194 1199 5198
rect 1203 5194 1215 5198
rect 1219 5194 1383 5198
rect 1387 5194 1399 5198
rect 1403 5194 1551 5198
rect 1555 5194 1607 5198
rect 1611 5194 1815 5198
rect 1819 5194 1935 5198
rect 1939 5194 1947 5198
rect 91 5193 1947 5194
rect 1953 5193 1954 5199
rect 1946 5101 1947 5107
rect 1953 5106 3811 5107
rect 1953 5102 1975 5106
rect 1979 5102 2119 5106
rect 2123 5102 2303 5106
rect 2307 5102 2327 5106
rect 2331 5102 2503 5106
rect 2507 5102 2535 5106
rect 2539 5102 2711 5106
rect 2715 5102 2751 5106
rect 2755 5102 2919 5106
rect 2923 5102 2975 5106
rect 2979 5102 3127 5106
rect 3131 5102 3207 5106
rect 3211 5102 3335 5106
rect 3339 5102 3799 5106
rect 3803 5102 3811 5106
rect 1953 5101 3811 5102
rect 3817 5103 3818 5107
rect 3817 5102 5702 5103
rect 3817 5101 3839 5102
rect 3810 5098 3839 5101
rect 3843 5098 3887 5102
rect 3891 5098 4087 5102
rect 4091 5098 4327 5102
rect 4331 5098 4463 5102
rect 4467 5098 4567 5102
rect 4571 5098 4623 5102
rect 4627 5098 4783 5102
rect 4787 5098 4815 5102
rect 4819 5098 4943 5102
rect 4947 5098 5063 5102
rect 5067 5098 5095 5102
rect 5099 5098 5247 5102
rect 5251 5098 5311 5102
rect 5315 5098 5407 5102
rect 5411 5098 5543 5102
rect 5547 5098 5663 5102
rect 5667 5098 5702 5102
rect 3810 5097 5702 5098
rect 96 5073 97 5079
rect 103 5078 1959 5079
rect 103 5074 111 5078
rect 115 5074 155 5078
rect 159 5074 379 5078
rect 383 5074 419 5078
rect 423 5074 595 5078
rect 599 5074 627 5078
rect 631 5074 779 5078
rect 783 5074 899 5078
rect 903 5074 971 5078
rect 975 5074 1171 5078
rect 1175 5074 1195 5078
rect 1199 5074 1371 5078
rect 1375 5074 1499 5078
rect 1503 5074 1579 5078
rect 1583 5074 1787 5078
rect 1791 5074 1935 5078
rect 1939 5074 1959 5078
rect 103 5073 1959 5074
rect 1965 5073 1966 5079
rect 3822 4990 5714 4991
rect 3822 4987 3839 4990
rect 1958 4981 1959 4987
rect 1965 4986 3823 4987
rect 1965 4982 1975 4986
rect 1979 4982 1995 4986
rect 1999 4982 2091 4986
rect 2095 4982 2131 4986
rect 2135 4982 2267 4986
rect 2271 4982 2299 4986
rect 2303 4982 2419 4986
rect 2423 4982 2507 4986
rect 2511 4982 2619 4986
rect 2623 4982 2723 4986
rect 2727 4982 2859 4986
rect 2863 4982 2947 4986
rect 2951 4982 3123 4986
rect 3127 4982 3179 4986
rect 3183 4982 3395 4986
rect 3399 4982 3651 4986
rect 3655 4982 3799 4986
rect 3803 4982 3823 4986
rect 1965 4981 3823 4982
rect 3829 4986 3839 4987
rect 3843 4986 3859 4990
rect 3863 4986 3995 4990
rect 3999 4986 4059 4990
rect 4063 4986 4131 4990
rect 4135 4986 4267 4990
rect 4271 4986 4299 4990
rect 4303 4986 4403 4990
rect 4407 4986 4539 4990
rect 4543 4986 4675 4990
rect 4679 4986 4787 4990
rect 4791 4986 4811 4990
rect 4815 4986 4947 4990
rect 4951 4986 5035 4990
rect 5039 4986 5083 4990
rect 5087 4986 5227 4990
rect 5231 4986 5283 4990
rect 5287 4986 5379 4990
rect 5383 4986 5515 4990
rect 5519 4986 5663 4990
rect 5667 4986 5714 4990
rect 3829 4985 5714 4986
rect 3829 4981 3830 4985
rect 4874 4972 4880 4973
rect 5238 4972 5244 4973
rect 4874 4968 4875 4972
rect 4879 4968 5239 4972
rect 5243 4968 5244 4972
rect 4874 4967 4880 4968
rect 5238 4967 5244 4968
rect 84 4933 85 4939
rect 91 4938 1947 4939
rect 91 4934 111 4938
rect 115 4934 159 4938
rect 163 4934 183 4938
rect 187 4934 295 4938
rect 299 4934 407 4938
rect 411 4934 431 4938
rect 435 4934 567 4938
rect 571 4934 655 4938
rect 659 4934 703 4938
rect 707 4934 927 4938
rect 931 4934 1223 4938
rect 1227 4934 1527 4938
rect 1531 4934 1815 4938
rect 1819 4934 1935 4938
rect 1939 4934 1947 4938
rect 91 4933 1947 4934
rect 1953 4933 1954 4939
rect 1946 4861 1947 4867
rect 1953 4866 3811 4867
rect 1953 4862 1975 4866
rect 1979 4862 2023 4866
rect 2027 4862 2159 4866
rect 2163 4862 2295 4866
rect 2299 4862 2327 4866
rect 2331 4862 2447 4866
rect 2451 4862 2559 4866
rect 2563 4862 2647 4866
rect 2651 4862 2823 4866
rect 2827 4862 2887 4866
rect 2891 4862 3103 4866
rect 3107 4862 3151 4866
rect 3155 4862 3399 4866
rect 3403 4862 3423 4866
rect 3427 4862 3679 4866
rect 3683 4862 3799 4866
rect 3803 4862 3811 4866
rect 1953 4861 3811 4862
rect 3817 4861 3818 4867
rect 96 4809 97 4815
rect 103 4814 1959 4815
rect 103 4810 111 4814
rect 115 4810 131 4814
rect 135 4810 267 4814
rect 271 4810 403 4814
rect 407 4810 539 4814
rect 543 4810 675 4814
rect 679 4810 1935 4814
rect 1939 4810 1959 4814
rect 103 4809 1959 4810
rect 1965 4809 1966 4815
rect 3810 4797 3811 4803
rect 3817 4802 5695 4803
rect 3817 4798 3839 4802
rect 3843 4798 3887 4802
rect 3891 4798 4023 4802
rect 4027 4798 4071 4802
rect 4075 4798 4159 4802
rect 4163 4798 4295 4802
rect 4299 4798 4431 4802
rect 4435 4798 4535 4802
rect 4539 4798 4567 4802
rect 4571 4798 4703 4802
rect 4707 4798 4783 4802
rect 4787 4798 4839 4802
rect 4843 4798 4975 4802
rect 4979 4798 5039 4802
rect 5043 4798 5111 4802
rect 5115 4798 5255 4802
rect 5259 4798 5303 4802
rect 5307 4798 5407 4802
rect 5411 4798 5543 4802
rect 5547 4798 5663 4802
rect 5667 4798 5695 4802
rect 3817 4797 5695 4798
rect 5701 4797 5702 4803
rect 1958 4737 1959 4743
rect 1965 4742 3823 4743
rect 1965 4738 1975 4742
rect 1979 4738 2019 4742
rect 2023 4738 2195 4742
rect 2199 4738 2299 4742
rect 2303 4738 2371 4742
rect 2375 4738 2531 4742
rect 2535 4738 2547 4742
rect 2551 4738 2723 4742
rect 2727 4738 2795 4742
rect 2799 4738 3075 4742
rect 3079 4738 3371 4742
rect 3375 4738 3651 4742
rect 3655 4738 3799 4742
rect 3803 4738 3823 4742
rect 1965 4737 3823 4738
rect 3829 4737 3830 4743
rect 84 4693 85 4699
rect 91 4698 1947 4699
rect 91 4694 111 4698
rect 115 4694 159 4698
rect 163 4694 295 4698
rect 299 4694 431 4698
rect 435 4694 567 4698
rect 571 4694 703 4698
rect 707 4694 1935 4698
rect 1939 4694 1947 4698
rect 91 4693 1947 4694
rect 1953 4693 1954 4699
rect 3822 4685 3823 4691
rect 3829 4690 5707 4691
rect 3829 4686 3839 4690
rect 3843 4686 3859 4690
rect 3863 4686 3995 4690
rect 3999 4686 4043 4690
rect 4047 4686 4131 4690
rect 4135 4686 4267 4690
rect 4271 4686 4403 4690
rect 4407 4686 4507 4690
rect 4511 4686 4539 4690
rect 4543 4686 4675 4690
rect 4679 4686 4755 4690
rect 4759 4686 4819 4690
rect 4823 4686 4963 4690
rect 4967 4686 5011 4690
rect 5015 4686 5107 4690
rect 5111 4686 5243 4690
rect 5247 4686 5275 4690
rect 5279 4686 5379 4690
rect 5383 4686 5515 4690
rect 5519 4686 5663 4690
rect 5667 4686 5707 4690
rect 3829 4685 5707 4686
rect 5713 4685 5714 4691
rect 1946 4621 1947 4627
rect 1953 4626 3811 4627
rect 1953 4622 1975 4626
rect 1979 4622 2023 4626
rect 2027 4622 2047 4626
rect 2051 4622 2223 4626
rect 2227 4622 2263 4626
rect 2267 4622 2399 4626
rect 2403 4622 2527 4626
rect 2531 4622 2575 4626
rect 2579 4622 2751 4626
rect 2755 4622 2775 4626
rect 2779 4622 3015 4626
rect 3019 4622 3247 4626
rect 3251 4622 3471 4626
rect 3475 4622 3679 4626
rect 3683 4622 3799 4626
rect 3803 4622 3811 4626
rect 1953 4621 3811 4622
rect 3817 4621 3818 4627
rect 96 4569 97 4575
rect 103 4574 1959 4575
rect 103 4570 111 4574
rect 115 4570 131 4574
rect 135 4570 251 4574
rect 255 4570 267 4574
rect 271 4570 403 4574
rect 407 4570 443 4574
rect 447 4570 539 4574
rect 543 4570 651 4574
rect 655 4570 675 4574
rect 679 4570 875 4574
rect 879 4570 1099 4574
rect 1103 4570 1331 4574
rect 1335 4570 1571 4574
rect 1575 4570 1787 4574
rect 1791 4570 1935 4574
rect 1939 4570 1959 4574
rect 103 4569 1959 4570
rect 1965 4569 1966 4575
rect 3810 4573 3811 4579
rect 3817 4578 5695 4579
rect 3817 4574 3839 4578
rect 3843 4574 3887 4578
rect 3891 4574 4023 4578
rect 4027 4574 4159 4578
rect 4163 4574 4295 4578
rect 4299 4574 4431 4578
rect 4435 4574 4567 4578
rect 4571 4574 4671 4578
rect 4675 4574 4703 4578
rect 4707 4574 4807 4578
rect 4811 4574 4847 4578
rect 4851 4574 4943 4578
rect 4947 4574 4991 4578
rect 4995 4574 5079 4578
rect 5083 4574 5135 4578
rect 5139 4574 5271 4578
rect 5275 4574 5407 4578
rect 5411 4574 5543 4578
rect 5547 4574 5663 4578
rect 5667 4574 5695 4578
rect 3817 4573 5695 4574
rect 5701 4573 5702 4579
rect 1958 4497 1959 4503
rect 1965 4502 3823 4503
rect 1965 4498 1975 4502
rect 1979 4498 1995 4502
rect 1999 4498 2235 4502
rect 2239 4498 2267 4502
rect 2271 4498 2499 4502
rect 2503 4498 2515 4502
rect 2519 4498 2747 4502
rect 2751 4498 2971 4502
rect 2975 4498 2987 4502
rect 2991 4498 3187 4502
rect 3191 4498 3219 4502
rect 3223 4498 3395 4502
rect 3399 4498 3443 4502
rect 3447 4498 3611 4502
rect 3615 4498 3651 4502
rect 3655 4498 3799 4502
rect 3803 4498 3823 4502
rect 1965 4497 3823 4498
rect 3829 4497 3830 4503
rect 3074 4492 3080 4493
rect 3734 4492 3740 4493
rect 3074 4488 3075 4492
rect 3079 4488 3735 4492
rect 3739 4488 3740 4492
rect 3074 4487 3080 4488
rect 3734 4487 3740 4488
rect 84 4457 85 4463
rect 91 4462 1947 4463
rect 91 4458 111 4462
rect 115 4458 279 4462
rect 283 4458 471 4462
rect 475 4458 511 4462
rect 515 4458 679 4462
rect 683 4458 687 4462
rect 691 4458 871 4462
rect 875 4458 903 4462
rect 907 4458 1071 4462
rect 1075 4458 1127 4462
rect 1131 4458 1279 4462
rect 1283 4458 1359 4462
rect 1363 4458 1495 4462
rect 1499 4458 1599 4462
rect 1603 4458 1719 4462
rect 1723 4458 1815 4462
rect 1819 4458 1935 4462
rect 1939 4458 1947 4462
rect 91 4457 1947 4458
rect 1953 4457 1954 4463
rect 3822 4457 3823 4463
rect 3829 4462 5707 4463
rect 3829 4458 3839 4462
rect 3843 4458 4347 4462
rect 4351 4458 4483 4462
rect 4487 4458 4619 4462
rect 4623 4458 4643 4462
rect 4647 4458 4755 4462
rect 4759 4458 4779 4462
rect 4783 4458 4891 4462
rect 4895 4458 4915 4462
rect 4919 4458 5051 4462
rect 5055 4458 5663 4462
rect 5667 4458 5707 4462
rect 3829 4457 5707 4458
rect 5713 4457 5714 4463
rect 1946 4373 1947 4379
rect 1953 4378 3811 4379
rect 1953 4374 1975 4378
rect 1979 4374 2023 4378
rect 2027 4374 2199 4378
rect 2203 4374 2295 4378
rect 2299 4374 2399 4378
rect 2403 4374 2543 4378
rect 2547 4374 2591 4378
rect 2595 4374 2775 4378
rect 2779 4374 2951 4378
rect 2955 4374 2999 4378
rect 3003 4374 3135 4378
rect 3139 4374 3215 4378
rect 3219 4374 3319 4378
rect 3323 4374 3423 4378
rect 3427 4374 3639 4378
rect 3643 4374 3799 4378
rect 3803 4374 3811 4378
rect 1953 4373 3811 4374
rect 3817 4373 3818 4379
rect 96 4341 97 4347
rect 103 4346 1959 4347
rect 103 4342 111 4346
rect 115 4342 483 4346
rect 487 4342 659 4346
rect 663 4342 715 4346
rect 719 4342 843 4346
rect 847 4342 851 4346
rect 855 4342 987 4346
rect 991 4342 1043 4346
rect 1047 4342 1123 4346
rect 1127 4342 1251 4346
rect 1255 4342 1259 4346
rect 1263 4342 1395 4346
rect 1399 4342 1467 4346
rect 1471 4342 1531 4346
rect 1535 4342 1667 4346
rect 1671 4342 1691 4346
rect 1695 4342 1935 4346
rect 1939 4342 1959 4346
rect 103 4341 1959 4342
rect 1965 4341 1966 4347
rect 3810 4329 3811 4335
rect 3817 4334 5695 4335
rect 3817 4330 3839 4334
rect 3843 4330 4135 4334
rect 4139 4330 4271 4334
rect 4275 4330 4375 4334
rect 4379 4330 4407 4334
rect 4411 4330 4511 4334
rect 4515 4330 4543 4334
rect 4547 4330 4647 4334
rect 4651 4330 4679 4334
rect 4683 4330 4783 4334
rect 4787 4330 4919 4334
rect 4923 4330 5663 4334
rect 5667 4330 5695 4334
rect 3817 4329 5695 4330
rect 5701 4329 5702 4335
rect 1958 4257 1959 4263
rect 1965 4262 3823 4263
rect 1965 4258 1975 4262
rect 1979 4258 1995 4262
rect 1999 4258 2171 4262
rect 2175 4258 2243 4262
rect 2247 4258 2371 4262
rect 2375 4258 2507 4262
rect 2511 4258 2563 4262
rect 2567 4258 2747 4262
rect 2751 4258 2763 4262
rect 2767 4258 2923 4262
rect 2927 4258 3019 4262
rect 3023 4258 3107 4262
rect 3111 4258 3283 4262
rect 3287 4258 3291 4262
rect 3295 4258 3799 4262
rect 3803 4258 3823 4262
rect 1965 4257 3823 4258
rect 3829 4257 3830 4263
rect 84 4221 85 4227
rect 91 4226 1947 4227
rect 91 4222 111 4226
rect 115 4222 727 4226
rect 731 4222 743 4226
rect 747 4222 863 4226
rect 867 4222 879 4226
rect 883 4222 999 4226
rect 1003 4222 1015 4226
rect 1019 4222 1135 4226
rect 1139 4222 1151 4226
rect 1155 4222 1271 4226
rect 1275 4222 1287 4226
rect 1291 4222 1407 4226
rect 1411 4222 1423 4226
rect 1427 4222 1543 4226
rect 1547 4222 1559 4226
rect 1563 4222 1679 4226
rect 1683 4222 1695 4226
rect 1699 4222 1815 4226
rect 1819 4222 1935 4226
rect 1939 4222 1947 4226
rect 91 4221 1947 4222
rect 1953 4221 1954 4227
rect 3822 4205 3823 4211
rect 3829 4210 5707 4211
rect 3829 4206 3839 4210
rect 3843 4206 3971 4210
rect 3975 4206 4107 4210
rect 4111 4206 4243 4210
rect 4247 4206 4379 4210
rect 4383 4206 4515 4210
rect 4519 4206 4651 4210
rect 4655 4206 5663 4210
rect 5667 4206 5707 4210
rect 3829 4205 5707 4206
rect 5713 4205 5714 4211
rect 4058 4180 4064 4181
rect 4522 4180 4528 4181
rect 4058 4176 4059 4180
rect 4063 4176 4523 4180
rect 4527 4176 4528 4180
rect 4058 4175 4064 4176
rect 4522 4175 4528 4176
rect 1946 4133 1947 4139
rect 1953 4138 3811 4139
rect 1953 4134 1975 4138
rect 1979 4134 2023 4138
rect 2027 4134 2271 4138
rect 2275 4134 2535 4138
rect 2539 4134 2791 4138
rect 2795 4134 3047 4138
rect 3051 4134 3135 4138
rect 3139 4134 3271 4138
rect 3275 4134 3311 4138
rect 3315 4134 3407 4138
rect 3411 4134 3543 4138
rect 3547 4134 3679 4138
rect 3683 4134 3799 4138
rect 3803 4134 3811 4138
rect 1953 4133 3811 4134
rect 3817 4133 3818 4139
rect 96 4109 97 4115
rect 103 4114 1959 4115
rect 103 4110 111 4114
rect 115 4110 563 4114
rect 567 4110 699 4114
rect 703 4110 835 4114
rect 839 4110 971 4114
rect 975 4110 1107 4114
rect 1111 4110 1243 4114
rect 1247 4110 1379 4114
rect 1383 4110 1515 4114
rect 1519 4110 1651 4114
rect 1655 4110 1787 4114
rect 1791 4110 1935 4114
rect 1939 4110 1959 4114
rect 103 4109 1959 4110
rect 1965 4109 1966 4115
rect 3810 4069 3811 4075
rect 3817 4074 5695 4075
rect 3817 4070 3839 4074
rect 3843 4070 3887 4074
rect 3891 4070 3999 4074
rect 4003 4070 4023 4074
rect 4027 4070 4135 4074
rect 4139 4070 4159 4074
rect 4163 4070 4271 4074
rect 4275 4070 4295 4074
rect 4299 4070 4407 4074
rect 4411 4070 4431 4074
rect 4435 4070 4543 4074
rect 4547 4070 4567 4074
rect 4571 4070 4703 4074
rect 4707 4070 4839 4074
rect 4843 4070 5663 4074
rect 5667 4070 5695 4074
rect 3817 4069 5695 4070
rect 5701 4069 5702 4075
rect 84 3997 85 4003
rect 91 4002 1947 4003
rect 91 3998 111 4002
rect 115 3998 159 4002
rect 163 3998 327 4002
rect 331 3998 535 4002
rect 539 3998 591 4002
rect 595 3998 727 4002
rect 731 3998 751 4002
rect 755 3998 863 4002
rect 867 3998 967 4002
rect 971 3998 999 4002
rect 1003 3998 1135 4002
rect 1139 3998 1183 4002
rect 1187 3998 1271 4002
rect 1275 3998 1399 4002
rect 1403 3998 1407 4002
rect 1411 3998 1543 4002
rect 1547 3998 1615 4002
rect 1619 3998 1679 4002
rect 1683 3998 1815 4002
rect 1819 3998 1935 4002
rect 1939 3998 1947 4002
rect 91 3997 1947 3998
rect 1953 3997 1954 4003
rect 3822 3957 3823 3963
rect 3829 3962 5707 3963
rect 3829 3958 3839 3962
rect 3843 3958 3859 3962
rect 3863 3958 3995 3962
rect 3999 3958 4131 3962
rect 4135 3958 4147 3962
rect 4151 3958 4267 3962
rect 4271 3958 4299 3962
rect 4303 3958 4403 3962
rect 4407 3958 4459 3962
rect 4463 3958 4539 3962
rect 4543 3958 4619 3962
rect 4623 3958 4675 3962
rect 4679 3958 4779 3962
rect 4783 3958 4811 3962
rect 4815 3958 5663 3962
rect 5667 3958 5707 3962
rect 3829 3957 5707 3958
rect 5713 3957 5714 3963
rect 1958 3929 1959 3935
rect 1965 3934 3823 3935
rect 1965 3930 1975 3934
rect 1979 3930 1995 3934
rect 1999 3930 2403 3934
rect 2407 3930 2827 3934
rect 2831 3930 3107 3934
rect 3111 3930 3243 3934
rect 3247 3930 3251 3934
rect 3255 3930 3379 3934
rect 3383 3930 3515 3934
rect 3519 3930 3651 3934
rect 3655 3930 3799 3934
rect 3803 3930 3823 3934
rect 1965 3929 3823 3930
rect 3829 3929 3830 3935
rect 96 3885 97 3891
rect 103 3890 1959 3891
rect 103 3886 111 3890
rect 115 3886 131 3890
rect 135 3886 299 3890
rect 303 3886 355 3890
rect 359 3886 507 3890
rect 511 3886 619 3890
rect 623 3886 723 3890
rect 727 3886 899 3890
rect 903 3886 939 3890
rect 943 3886 1155 3890
rect 1159 3886 1195 3890
rect 1199 3886 1371 3890
rect 1375 3886 1499 3890
rect 1503 3886 1587 3890
rect 1591 3886 1787 3890
rect 1791 3886 1935 3890
rect 1939 3886 1959 3890
rect 103 3885 1959 3886
rect 1965 3885 1966 3891
rect 1946 3817 1947 3823
rect 1953 3822 3811 3823
rect 1953 3818 1975 3822
rect 1979 3818 2023 3822
rect 2027 3818 2175 3822
rect 2179 3818 2351 3822
rect 2355 3818 2431 3822
rect 2435 3818 2535 3822
rect 2539 3818 2719 3822
rect 2723 3818 2855 3822
rect 2859 3818 2895 3822
rect 2899 3818 3071 3822
rect 3075 3818 3247 3822
rect 3251 3818 3279 3822
rect 3283 3818 3423 3822
rect 3427 3818 3607 3822
rect 3611 3818 3679 3822
rect 3683 3818 3799 3822
rect 3803 3818 3811 3822
rect 1953 3817 3811 3818
rect 3817 3822 5702 3823
rect 3817 3818 3839 3822
rect 3843 3818 3887 3822
rect 3891 3818 4023 3822
rect 4027 3818 4175 3822
rect 4179 3818 4327 3822
rect 4331 3818 4487 3822
rect 4491 3818 4503 3822
rect 4507 3818 4639 3822
rect 4643 3818 4647 3822
rect 4651 3818 4775 3822
rect 4779 3818 4807 3822
rect 4811 3818 4911 3822
rect 4915 3818 5047 3822
rect 5051 3818 5663 3822
rect 5667 3818 5702 3822
rect 3817 3817 5702 3818
rect 84 3761 85 3767
rect 91 3766 1947 3767
rect 91 3762 111 3766
rect 115 3762 159 3766
rect 163 3762 247 3766
rect 251 3762 383 3766
rect 387 3762 519 3766
rect 523 3762 647 3766
rect 651 3762 791 3766
rect 795 3762 927 3766
rect 931 3762 1063 3766
rect 1067 3762 1223 3766
rect 1227 3762 1343 3766
rect 1347 3762 1527 3766
rect 1531 3762 1815 3766
rect 1819 3762 1935 3766
rect 1939 3762 1947 3766
rect 91 3761 1947 3762
rect 1953 3761 1954 3767
rect 1958 3697 1959 3703
rect 1965 3702 3823 3703
rect 1965 3698 1975 3702
rect 1979 3698 1995 3702
rect 1999 3698 2011 3702
rect 2015 3698 2147 3702
rect 2151 3698 2291 3702
rect 2295 3698 2323 3702
rect 2327 3698 2435 3702
rect 2439 3698 2507 3702
rect 2511 3698 2579 3702
rect 2583 3698 2691 3702
rect 2695 3698 2723 3702
rect 2727 3698 2867 3702
rect 2871 3698 3011 3702
rect 3015 3698 3043 3702
rect 3047 3698 3155 3702
rect 3159 3698 3219 3702
rect 3223 3698 3299 3702
rect 3303 3698 3395 3702
rect 3399 3698 3579 3702
rect 3583 3698 3799 3702
rect 3803 3698 3823 3702
rect 1965 3697 3823 3698
rect 3829 3697 3830 3703
rect 3822 3685 3823 3691
rect 3829 3690 5707 3691
rect 3829 3686 3839 3690
rect 3843 3686 4019 3690
rect 4023 3686 4155 3690
rect 4159 3686 4291 3690
rect 4295 3686 4427 3690
rect 4431 3686 4475 3690
rect 4479 3686 4563 3690
rect 4567 3686 4611 3690
rect 4615 3686 4699 3690
rect 4703 3686 4747 3690
rect 4751 3686 4835 3690
rect 4839 3686 4883 3690
rect 4887 3686 4971 3690
rect 4975 3686 5019 3690
rect 5023 3686 5107 3690
rect 5111 3686 5243 3690
rect 5247 3686 5379 3690
rect 5383 3686 5515 3690
rect 5519 3686 5663 3690
rect 5667 3686 5707 3690
rect 3829 3685 5707 3686
rect 5713 3685 5714 3691
rect 96 3633 97 3639
rect 103 3638 1959 3639
rect 103 3634 111 3638
rect 115 3634 219 3638
rect 223 3634 491 3638
rect 495 3634 635 3638
rect 639 3634 763 3638
rect 767 3634 779 3638
rect 783 3634 923 3638
rect 927 3634 1035 3638
rect 1039 3634 1067 3638
rect 1071 3634 1211 3638
rect 1215 3634 1315 3638
rect 1319 3634 1935 3638
rect 1939 3634 1959 3638
rect 103 3633 1959 3634
rect 1965 3633 1966 3639
rect 1946 3577 1947 3583
rect 1953 3582 3811 3583
rect 1953 3578 1975 3582
rect 1979 3578 2039 3582
rect 2043 3578 2175 3582
rect 2179 3578 2239 3582
rect 2243 3578 2319 3582
rect 2323 3578 2375 3582
rect 2379 3578 2463 3582
rect 2467 3578 2511 3582
rect 2515 3578 2607 3582
rect 2611 3578 2647 3582
rect 2651 3578 2751 3582
rect 2755 3578 2783 3582
rect 2787 3578 2895 3582
rect 2899 3578 2919 3582
rect 2923 3578 3039 3582
rect 3043 3578 3055 3582
rect 3059 3578 3183 3582
rect 3187 3578 3191 3582
rect 3195 3578 3327 3582
rect 3331 3578 3463 3582
rect 3467 3578 3799 3582
rect 3803 3578 3811 3582
rect 1953 3577 3811 3578
rect 3817 3577 3818 3583
rect 3810 3525 3811 3531
rect 3817 3530 5695 3531
rect 3817 3526 3839 3530
rect 3843 3526 4047 3530
rect 4051 3526 4183 3530
rect 4187 3526 4319 3530
rect 4323 3526 4455 3530
rect 4459 3526 4591 3530
rect 4595 3526 4727 3530
rect 4731 3526 4863 3530
rect 4867 3526 4999 3530
rect 5003 3526 5135 3530
rect 5139 3526 5271 3530
rect 5275 3526 5407 3530
rect 5411 3526 5543 3530
rect 5547 3526 5663 3530
rect 5667 3526 5695 3530
rect 3817 3525 5695 3526
rect 5701 3525 5702 3531
rect 84 3501 85 3507
rect 91 3506 1947 3507
rect 91 3502 111 3506
rect 115 3502 431 3506
rect 435 3502 519 3506
rect 523 3502 567 3506
rect 571 3502 663 3506
rect 667 3502 703 3506
rect 707 3502 807 3506
rect 811 3502 839 3506
rect 843 3502 951 3506
rect 955 3502 975 3506
rect 979 3502 1095 3506
rect 1099 3502 1239 3506
rect 1243 3502 1935 3506
rect 1939 3502 1947 3506
rect 91 3501 1947 3502
rect 1953 3501 1954 3507
rect 1958 3461 1959 3467
rect 1965 3466 3823 3467
rect 1965 3462 1975 3466
rect 1979 3462 2171 3466
rect 2175 3462 2211 3466
rect 2215 3462 2347 3466
rect 2351 3462 2483 3466
rect 2487 3462 2531 3466
rect 2535 3462 2619 3466
rect 2623 3462 2715 3466
rect 2719 3462 2755 3466
rect 2759 3462 2891 3466
rect 2895 3462 2907 3466
rect 2911 3462 3027 3466
rect 3031 3462 3099 3466
rect 3103 3462 3163 3466
rect 3167 3462 3291 3466
rect 3295 3462 3299 3466
rect 3303 3462 3435 3466
rect 3439 3462 3483 3466
rect 3487 3462 3651 3466
rect 3655 3462 3799 3466
rect 3803 3462 3823 3466
rect 1965 3461 3823 3462
rect 3829 3461 3830 3467
rect 3822 3405 3823 3411
rect 3829 3410 5707 3411
rect 3829 3406 3839 3410
rect 3843 3406 3859 3410
rect 3863 3406 4099 3410
rect 4103 3406 4347 3410
rect 4351 3406 4587 3410
rect 4591 3406 4811 3410
rect 4815 3406 5027 3410
rect 5031 3406 5235 3410
rect 5239 3406 5379 3410
rect 5383 3406 5451 3410
rect 5455 3406 5515 3410
rect 5519 3406 5663 3410
rect 5667 3406 5707 3410
rect 3829 3405 5707 3406
rect 5713 3405 5714 3411
rect 96 3381 97 3387
rect 103 3386 1959 3387
rect 103 3382 111 3386
rect 115 3382 323 3386
rect 327 3382 403 3386
rect 407 3382 459 3386
rect 463 3382 539 3386
rect 543 3382 595 3386
rect 599 3382 675 3386
rect 679 3382 731 3386
rect 735 3382 811 3386
rect 815 3382 867 3386
rect 871 3382 947 3386
rect 951 3382 1935 3386
rect 1939 3382 1959 3386
rect 103 3381 1959 3382
rect 1965 3381 1966 3387
rect 1946 3325 1947 3331
rect 1953 3330 3811 3331
rect 1953 3326 1975 3330
rect 1979 3326 2151 3330
rect 2155 3326 2199 3330
rect 2203 3326 2375 3330
rect 2379 3326 2399 3330
rect 2403 3326 2559 3330
rect 2563 3326 2687 3330
rect 2691 3326 2743 3330
rect 2747 3326 2935 3330
rect 2939 3326 3015 3330
rect 3019 3326 3127 3330
rect 3131 3326 3319 3330
rect 3323 3326 3359 3330
rect 3363 3326 3511 3330
rect 3515 3326 3679 3330
rect 3683 3326 3799 3330
rect 3803 3326 3811 3330
rect 1953 3325 3811 3326
rect 3817 3325 3818 3331
rect 3810 3293 3811 3299
rect 3817 3298 5695 3299
rect 3817 3294 3839 3298
rect 3843 3294 3887 3298
rect 3891 3294 4127 3298
rect 4131 3294 4375 3298
rect 4379 3294 4607 3298
rect 4611 3294 4615 3298
rect 4619 3294 4815 3298
rect 4819 3294 4839 3298
rect 4843 3294 5015 3298
rect 5019 3294 5055 3298
rect 5059 3294 5199 3298
rect 5203 3294 5263 3298
rect 5267 3294 5383 3298
rect 5387 3294 5479 3298
rect 5483 3294 5543 3298
rect 5547 3294 5663 3298
rect 5667 3294 5695 3298
rect 3817 3293 5695 3294
rect 5701 3293 5702 3299
rect 84 3261 85 3267
rect 91 3266 1947 3267
rect 91 3262 111 3266
rect 115 3262 159 3266
rect 163 3262 335 3266
rect 339 3262 351 3266
rect 355 3262 487 3266
rect 491 3262 543 3266
rect 547 3262 623 3266
rect 627 3262 751 3266
rect 755 3262 759 3266
rect 763 3262 895 3266
rect 899 3262 959 3266
rect 963 3262 1935 3266
rect 1939 3262 1947 3266
rect 91 3261 1947 3262
rect 1953 3261 1954 3267
rect 1958 3213 1959 3219
rect 1965 3218 3823 3219
rect 1965 3214 1975 3218
rect 1979 3214 1995 3218
rect 1999 3214 2123 3218
rect 2127 3214 2147 3218
rect 2151 3214 2347 3218
rect 2351 3214 2371 3218
rect 2375 3214 2555 3218
rect 2559 3214 2659 3218
rect 2663 3214 2771 3218
rect 2775 3214 2987 3218
rect 2991 3214 3211 3218
rect 3215 3214 3331 3218
rect 3335 3214 3443 3218
rect 3447 3214 3651 3218
rect 3655 3214 3799 3218
rect 3803 3214 3823 3218
rect 1965 3213 3823 3214
rect 3829 3213 3830 3219
rect 3822 3165 3823 3171
rect 3829 3170 5707 3171
rect 3829 3166 3839 3170
rect 3843 3166 3859 3170
rect 3863 3166 4099 3170
rect 4103 3166 4347 3170
rect 4351 3166 4467 3170
rect 4471 3166 4579 3170
rect 4583 3166 4651 3170
rect 4655 3166 4787 3170
rect 4791 3166 4859 3170
rect 4863 3166 4987 3170
rect 4991 3166 5075 3170
rect 5079 3166 5171 3170
rect 5175 3166 5307 3170
rect 5311 3166 5355 3170
rect 5359 3166 5515 3170
rect 5519 3166 5663 3170
rect 5667 3166 5707 3170
rect 3829 3165 5707 3166
rect 5713 3165 5714 3171
rect 96 3133 97 3139
rect 103 3138 1959 3139
rect 103 3134 111 3138
rect 115 3134 131 3138
rect 135 3134 307 3138
rect 311 3134 371 3138
rect 375 3134 515 3138
rect 519 3134 627 3138
rect 631 3134 723 3138
rect 727 3134 875 3138
rect 879 3134 931 3138
rect 935 3134 1115 3138
rect 1119 3134 1347 3138
rect 1351 3134 1579 3138
rect 1583 3134 1787 3138
rect 1791 3134 1935 3138
rect 1939 3134 1959 3138
rect 103 3133 1959 3134
rect 1965 3133 1966 3139
rect 1946 3101 1947 3107
rect 1953 3106 3811 3107
rect 1953 3102 1975 3106
rect 1979 3102 2023 3106
rect 2027 3102 2175 3106
rect 2179 3102 2375 3106
rect 2379 3102 2583 3106
rect 2587 3102 2647 3106
rect 2651 3102 2783 3106
rect 2787 3102 2799 3106
rect 2803 3102 2927 3106
rect 2931 3102 3015 3106
rect 3019 3102 3079 3106
rect 3083 3102 3239 3106
rect 3243 3102 3399 3106
rect 3403 3102 3471 3106
rect 3475 3102 3567 3106
rect 3571 3102 3679 3106
rect 3683 3102 3799 3106
rect 3803 3102 3811 3106
rect 1953 3101 3811 3102
rect 3817 3101 3818 3107
rect 3810 3053 3811 3059
rect 3817 3058 5695 3059
rect 3817 3054 3839 3058
rect 3843 3054 4255 3058
rect 4259 3054 4455 3058
rect 4459 3054 4495 3058
rect 4499 3054 4671 3058
rect 4675 3054 4679 3058
rect 4683 3054 4887 3058
rect 4891 3054 4911 3058
rect 4915 3054 5103 3058
rect 5107 3054 5167 3058
rect 5171 3054 5335 3058
rect 5339 3054 5423 3058
rect 5427 3054 5543 3058
rect 5547 3054 5663 3058
rect 5667 3054 5695 3058
rect 3817 3053 5695 3054
rect 5701 3053 5702 3059
rect 84 3021 85 3027
rect 91 3026 1947 3027
rect 91 3022 111 3026
rect 115 3022 159 3026
rect 163 3022 175 3026
rect 179 3022 399 3026
rect 403 3022 407 3026
rect 411 3022 623 3026
rect 627 3022 655 3026
rect 659 3022 823 3026
rect 827 3022 903 3026
rect 907 3022 1007 3026
rect 1011 3022 1143 3026
rect 1147 3022 1183 3026
rect 1187 3022 1351 3026
rect 1355 3022 1375 3026
rect 1379 3022 1511 3026
rect 1515 3022 1607 3026
rect 1611 3022 1671 3026
rect 1675 3022 1815 3026
rect 1819 3022 1935 3026
rect 1939 3022 1947 3026
rect 91 3021 1947 3022
rect 1953 3021 1954 3027
rect 1958 2989 1959 2995
rect 1965 2994 3823 2995
rect 1965 2990 1975 2994
rect 1979 2990 2619 2994
rect 2623 2990 2755 2994
rect 2759 2990 2803 2994
rect 2807 2990 2899 2994
rect 2903 2990 2939 2994
rect 2943 2990 3051 2994
rect 3055 2990 3075 2994
rect 3079 2990 3211 2994
rect 3215 2990 3347 2994
rect 3351 2990 3371 2994
rect 3375 2990 3483 2994
rect 3487 2990 3539 2994
rect 3543 2990 3799 2994
rect 3803 2990 3823 2994
rect 1965 2989 3823 2990
rect 3829 2989 3830 2995
rect 3822 2917 3823 2923
rect 3829 2922 5707 2923
rect 3829 2918 3839 2922
rect 3843 2918 3995 2922
rect 3999 2918 4211 2922
rect 4215 2918 4227 2922
rect 4231 2918 4427 2922
rect 4431 2918 4443 2922
rect 4447 2918 4643 2922
rect 4647 2918 4699 2922
rect 4703 2918 4883 2922
rect 4887 2918 4971 2922
rect 4975 2918 5139 2922
rect 5143 2918 5251 2922
rect 5255 2918 5395 2922
rect 5399 2918 5515 2922
rect 5519 2918 5663 2922
rect 5667 2918 5707 2922
rect 3829 2917 5707 2918
rect 5713 2917 5714 2923
rect 96 2905 97 2911
rect 103 2910 1959 2911
rect 103 2906 111 2910
rect 115 2906 147 2910
rect 151 2906 379 2910
rect 383 2906 395 2910
rect 399 2906 595 2910
rect 599 2906 787 2910
rect 791 2906 795 2910
rect 799 2906 971 2910
rect 975 2906 979 2910
rect 983 2906 1147 2910
rect 1151 2906 1155 2910
rect 1159 2906 1315 2910
rect 1319 2906 1323 2910
rect 1327 2906 1483 2910
rect 1487 2906 1643 2910
rect 1647 2906 1787 2910
rect 1791 2906 1935 2910
rect 1939 2906 1959 2910
rect 103 2905 1959 2906
rect 1965 2905 1966 2911
rect 1946 2825 1947 2831
rect 1953 2830 3811 2831
rect 1953 2826 1975 2830
rect 1979 2826 2023 2830
rect 2027 2826 2167 2830
rect 2171 2826 2335 2830
rect 2339 2826 2495 2830
rect 2499 2826 2663 2830
rect 2667 2826 2831 2830
rect 2835 2826 2967 2830
rect 2971 2826 2999 2830
rect 3003 2826 3103 2830
rect 3107 2826 3167 2830
rect 3171 2826 3239 2830
rect 3243 2826 3375 2830
rect 3379 2826 3511 2830
rect 3515 2826 3799 2830
rect 3803 2826 3811 2830
rect 1953 2825 3811 2826
rect 3817 2825 3818 2831
rect 3810 2801 3811 2807
rect 3817 2806 5695 2807
rect 3817 2802 3839 2806
rect 3843 2802 3919 2806
rect 3923 2802 4023 2806
rect 4027 2802 4055 2806
rect 4059 2802 4191 2806
rect 4195 2802 4239 2806
rect 4243 2802 4327 2806
rect 4331 2802 4463 2806
rect 4467 2802 4471 2806
rect 4475 2802 4727 2806
rect 4731 2802 4999 2806
rect 5003 2802 5279 2806
rect 5283 2802 5543 2806
rect 5547 2802 5663 2806
rect 5667 2802 5695 2806
rect 3817 2801 5695 2802
rect 5701 2801 5702 2807
rect 84 2781 85 2787
rect 91 2786 1947 2787
rect 91 2782 111 2786
rect 115 2782 423 2786
rect 427 2782 623 2786
rect 627 2782 655 2786
rect 659 2782 815 2786
rect 819 2782 975 2786
rect 979 2782 999 2786
rect 1003 2782 1143 2786
rect 1147 2782 1175 2786
rect 1179 2782 1311 2786
rect 1315 2782 1343 2786
rect 1347 2782 1479 2786
rect 1483 2782 1511 2786
rect 1515 2782 1671 2786
rect 1675 2782 1815 2786
rect 1819 2782 1935 2786
rect 1939 2782 1947 2786
rect 91 2781 1947 2782
rect 1953 2781 1954 2787
rect 1958 2713 1959 2719
rect 1965 2718 3823 2719
rect 1965 2714 1975 2718
rect 1979 2714 1995 2718
rect 1999 2714 2139 2718
rect 2143 2714 2307 2718
rect 2311 2714 2379 2718
rect 2383 2714 2467 2718
rect 2471 2714 2515 2718
rect 2519 2714 2635 2718
rect 2639 2714 2659 2718
rect 2663 2714 2803 2718
rect 2807 2714 2947 2718
rect 2951 2714 2971 2718
rect 2975 2714 3091 2718
rect 3095 2714 3139 2718
rect 3143 2714 3235 2718
rect 3239 2714 3799 2718
rect 3803 2714 3823 2718
rect 1965 2713 3823 2714
rect 3829 2713 3830 2719
rect 3822 2677 3823 2683
rect 3829 2682 5707 2683
rect 3829 2678 3839 2682
rect 3843 2678 3891 2682
rect 3895 2678 4027 2682
rect 4031 2678 4099 2682
rect 4103 2678 4163 2682
rect 4167 2678 4299 2682
rect 4303 2678 4435 2682
rect 4439 2678 4515 2682
rect 4519 2678 4755 2682
rect 4759 2678 5011 2682
rect 5015 2678 5275 2682
rect 5279 2678 5515 2682
rect 5519 2678 5663 2682
rect 5667 2678 5707 2682
rect 3829 2677 5707 2678
rect 5713 2677 5714 2683
rect 96 2669 97 2675
rect 103 2674 1959 2675
rect 103 2670 111 2674
rect 115 2670 627 2674
rect 631 2670 771 2674
rect 775 2670 787 2674
rect 791 2670 907 2674
rect 911 2670 947 2674
rect 951 2670 1043 2674
rect 1047 2670 1115 2674
rect 1119 2670 1179 2674
rect 1183 2670 1283 2674
rect 1287 2670 1315 2674
rect 1319 2670 1451 2674
rect 1455 2670 1587 2674
rect 1591 2670 1723 2674
rect 1727 2670 1935 2674
rect 1939 2670 1959 2674
rect 103 2669 1959 2670
rect 1965 2669 1966 2675
rect 1946 2597 1947 2603
rect 1953 2602 3811 2603
rect 1953 2598 1975 2602
rect 1979 2598 2407 2602
rect 2411 2598 2511 2602
rect 2515 2598 2543 2602
rect 2547 2598 2647 2602
rect 2651 2598 2687 2602
rect 2691 2598 2783 2602
rect 2787 2598 2831 2602
rect 2835 2598 2919 2602
rect 2923 2598 2975 2602
rect 2979 2598 3055 2602
rect 3059 2598 3119 2602
rect 3123 2598 3191 2602
rect 3195 2598 3263 2602
rect 3267 2598 3327 2602
rect 3331 2598 3463 2602
rect 3467 2598 3799 2602
rect 3803 2598 3811 2602
rect 1953 2597 3811 2598
rect 3817 2597 3818 2603
rect 3810 2561 3811 2567
rect 3817 2566 5695 2567
rect 3817 2562 3839 2566
rect 3843 2562 4127 2566
rect 4131 2562 4327 2566
rect 4331 2562 4495 2566
rect 4499 2562 4543 2566
rect 4547 2562 4631 2566
rect 4635 2562 4767 2566
rect 4771 2562 4783 2566
rect 4787 2562 4903 2566
rect 4907 2562 5039 2566
rect 5043 2562 5303 2566
rect 5307 2562 5543 2566
rect 5547 2562 5663 2566
rect 5667 2562 5695 2566
rect 3817 2561 5695 2562
rect 5701 2561 5702 2567
rect 84 2541 85 2547
rect 91 2546 1947 2547
rect 91 2542 111 2546
rect 115 2542 551 2546
rect 555 2542 687 2546
rect 691 2542 799 2546
rect 803 2542 831 2546
rect 835 2542 935 2546
rect 939 2542 983 2546
rect 987 2542 1071 2546
rect 1075 2542 1135 2546
rect 1139 2542 1207 2546
rect 1211 2542 1295 2546
rect 1299 2542 1343 2546
rect 1347 2542 1455 2546
rect 1459 2542 1479 2546
rect 1483 2542 1615 2546
rect 1619 2542 1751 2546
rect 1755 2542 1783 2546
rect 1787 2542 1935 2546
rect 1939 2542 1947 2546
rect 91 2541 1947 2542
rect 1953 2541 1954 2547
rect 1958 2469 1959 2475
rect 1965 2474 3823 2475
rect 1965 2470 1975 2474
rect 1979 2470 2307 2474
rect 2311 2470 2483 2474
rect 2487 2470 2515 2474
rect 2519 2470 2619 2474
rect 2623 2470 2715 2474
rect 2719 2470 2755 2474
rect 2759 2470 2891 2474
rect 2895 2470 2907 2474
rect 2911 2470 3027 2474
rect 3031 2470 3099 2474
rect 3103 2470 3163 2474
rect 3167 2470 3283 2474
rect 3287 2470 3299 2474
rect 3303 2470 3435 2474
rect 3439 2470 3467 2474
rect 3471 2470 3651 2474
rect 3655 2470 3799 2474
rect 3803 2470 3823 2474
rect 1965 2469 3823 2470
rect 3829 2469 3830 2475
rect 3822 2433 3823 2439
rect 3829 2438 5707 2439
rect 3829 2434 3839 2438
rect 3843 2434 4467 2438
rect 4471 2434 4603 2438
rect 4607 2434 4699 2438
rect 4703 2434 4739 2438
rect 4743 2434 4835 2438
rect 4839 2434 4875 2438
rect 4879 2434 4971 2438
rect 4975 2434 5011 2438
rect 5015 2434 5107 2438
rect 5111 2434 5243 2438
rect 5247 2434 5379 2438
rect 5383 2434 5515 2438
rect 5519 2434 5663 2438
rect 5667 2434 5707 2438
rect 3829 2433 5707 2434
rect 5713 2433 5714 2439
rect 96 2417 97 2423
rect 103 2422 1959 2423
rect 103 2418 111 2422
rect 115 2418 131 2422
rect 135 2418 339 2422
rect 343 2418 523 2422
rect 527 2418 563 2422
rect 567 2418 659 2422
rect 663 2418 803 2422
rect 807 2418 955 2422
rect 959 2418 1043 2422
rect 1047 2418 1107 2422
rect 1111 2418 1267 2422
rect 1271 2418 1291 2422
rect 1295 2418 1427 2422
rect 1431 2418 1547 2422
rect 1551 2418 1587 2422
rect 1591 2418 1755 2422
rect 1759 2418 1787 2422
rect 1791 2418 1935 2422
rect 1939 2418 1959 2422
rect 103 2417 1959 2418
rect 1965 2417 1966 2423
rect 1946 2349 1947 2355
rect 1953 2354 3811 2355
rect 1953 2350 1975 2354
rect 1979 2350 2223 2354
rect 2227 2350 2335 2354
rect 2339 2350 2503 2354
rect 2507 2350 2543 2354
rect 2547 2350 2743 2354
rect 2747 2350 2767 2354
rect 2771 2350 2935 2354
rect 2939 2350 3007 2354
rect 3011 2350 3127 2354
rect 3131 2350 3239 2354
rect 3243 2350 3311 2354
rect 3315 2350 3471 2354
rect 3475 2350 3495 2354
rect 3499 2350 3679 2354
rect 3683 2350 3799 2354
rect 3803 2350 3811 2354
rect 1953 2349 3811 2350
rect 3817 2349 3818 2355
rect 3810 2309 3811 2315
rect 3817 2314 5695 2315
rect 3817 2310 3839 2314
rect 3843 2310 3887 2314
rect 3891 2310 4183 2314
rect 4187 2310 4495 2314
rect 4499 2310 4727 2314
rect 4731 2310 4791 2314
rect 4795 2310 4863 2314
rect 4867 2310 4999 2314
rect 5003 2310 5087 2314
rect 5091 2310 5135 2314
rect 5139 2310 5271 2314
rect 5275 2310 5383 2314
rect 5387 2310 5407 2314
rect 5411 2310 5543 2314
rect 5547 2310 5663 2314
rect 5667 2310 5695 2314
rect 3817 2309 5695 2310
rect 5701 2309 5702 2315
rect 84 2301 85 2307
rect 91 2306 1947 2307
rect 91 2302 111 2306
rect 115 2302 159 2306
rect 163 2302 319 2306
rect 323 2302 367 2306
rect 371 2302 551 2306
rect 555 2302 591 2306
rect 595 2302 831 2306
rect 835 2302 1071 2306
rect 1075 2302 1151 2306
rect 1155 2302 1319 2306
rect 1323 2302 1495 2306
rect 1499 2302 1575 2306
rect 1579 2302 1815 2306
rect 1819 2302 1935 2306
rect 1939 2302 1947 2306
rect 91 2301 1947 2302
rect 1953 2301 1954 2307
rect 1958 2237 1959 2243
rect 1965 2242 3823 2243
rect 1965 2238 1975 2242
rect 1979 2238 1995 2242
rect 1999 2238 2155 2242
rect 2159 2238 2195 2242
rect 2199 2238 2387 2242
rect 2391 2238 2475 2242
rect 2479 2238 2667 2242
rect 2671 2238 2739 2242
rect 2743 2238 2979 2242
rect 2983 2238 2987 2242
rect 2991 2238 3211 2242
rect 3215 2238 3331 2242
rect 3335 2238 3443 2242
rect 3447 2238 3651 2242
rect 3655 2238 3799 2242
rect 3803 2238 3823 2242
rect 1965 2237 3823 2238
rect 3829 2237 3830 2243
rect 3822 2193 3823 2199
rect 3829 2198 5707 2199
rect 3829 2194 3839 2198
rect 3843 2194 3859 2198
rect 3863 2194 3995 2198
rect 3999 2194 4131 2198
rect 4135 2194 4155 2198
rect 4159 2194 4267 2198
rect 4271 2194 4403 2198
rect 4407 2194 4467 2198
rect 4471 2194 4539 2198
rect 4543 2194 4699 2198
rect 4703 2194 4763 2198
rect 4767 2194 4891 2198
rect 4895 2194 5059 2198
rect 5063 2194 5099 2198
rect 5103 2194 5315 2198
rect 5319 2194 5355 2198
rect 5359 2194 5515 2198
rect 5519 2194 5663 2198
rect 5667 2194 5707 2198
rect 3829 2193 5707 2194
rect 5713 2193 5714 2199
rect 96 2165 97 2171
rect 103 2170 1959 2171
rect 103 2166 111 2170
rect 115 2166 131 2170
rect 135 2166 291 2170
rect 295 2166 483 2170
rect 487 2166 523 2170
rect 527 2166 691 2170
rect 695 2166 803 2170
rect 807 2166 915 2170
rect 919 2166 1123 2170
rect 1127 2166 1147 2170
rect 1151 2166 1387 2170
rect 1391 2166 1467 2170
rect 1471 2166 1635 2170
rect 1639 2166 1787 2170
rect 1791 2166 1935 2170
rect 1939 2166 1959 2170
rect 103 2165 1959 2166
rect 1965 2165 1966 2171
rect 3810 2061 3811 2067
rect 3817 2066 5695 2067
rect 3817 2062 3839 2066
rect 3843 2062 3887 2066
rect 3891 2062 4023 2066
rect 4027 2062 4159 2066
rect 4163 2062 4295 2066
rect 4299 2062 4431 2066
rect 4435 2062 4567 2066
rect 4571 2062 4719 2066
rect 4723 2062 4727 2066
rect 4731 2062 4895 2066
rect 4899 2062 4919 2066
rect 4923 2062 5087 2066
rect 5091 2062 5127 2066
rect 5131 2062 5279 2066
rect 5283 2062 5343 2066
rect 5347 2062 5479 2066
rect 5483 2062 5543 2066
rect 5547 2062 5663 2066
rect 5667 2062 5695 2066
rect 3817 2061 5695 2062
rect 5701 2061 5702 2067
rect 84 2049 85 2055
rect 91 2054 1947 2055
rect 91 2050 111 2054
rect 115 2050 263 2054
rect 267 2050 319 2054
rect 323 2050 399 2054
rect 403 2050 511 2054
rect 515 2050 535 2054
rect 539 2050 679 2054
rect 683 2050 719 2054
rect 723 2050 823 2054
rect 827 2050 943 2054
rect 947 2050 967 2054
rect 971 2050 1111 2054
rect 1115 2050 1175 2054
rect 1179 2050 1255 2054
rect 1259 2050 1399 2054
rect 1403 2050 1415 2054
rect 1419 2050 1543 2054
rect 1547 2050 1663 2054
rect 1667 2050 1679 2054
rect 1683 2050 1815 2054
rect 1819 2050 1935 2054
rect 1939 2050 1947 2054
rect 91 2049 1947 2050
rect 1953 2049 1954 2055
rect 3822 1949 3823 1955
rect 3829 1954 5707 1955
rect 3829 1950 3839 1954
rect 3843 1950 3859 1954
rect 3863 1950 3995 1954
rect 3999 1950 4043 1954
rect 4047 1950 4131 1954
rect 4135 1950 4267 1954
rect 4271 1950 4283 1954
rect 4287 1950 4403 1954
rect 4407 1950 4539 1954
rect 4543 1950 4563 1954
rect 4567 1950 4691 1954
rect 4695 1950 4867 1954
rect 4871 1950 4875 1954
rect 4879 1950 5059 1954
rect 5063 1950 5203 1954
rect 5207 1950 5251 1954
rect 5255 1950 5451 1954
rect 5455 1950 5515 1954
rect 5519 1950 5663 1954
rect 5667 1950 5707 1954
rect 3829 1949 5707 1950
rect 5713 1949 5714 1955
rect 1946 1935 1947 1941
rect 1953 1935 1978 1941
rect 1972 1931 1978 1935
rect 96 1925 97 1931
rect 103 1930 1959 1931
rect 103 1926 111 1930
rect 115 1926 235 1930
rect 239 1926 371 1930
rect 375 1926 435 1930
rect 439 1926 507 1930
rect 511 1926 627 1930
rect 631 1926 651 1930
rect 655 1926 795 1930
rect 799 1926 811 1930
rect 815 1926 939 1930
rect 943 1926 987 1930
rect 991 1926 1083 1930
rect 1087 1926 1155 1930
rect 1159 1926 1227 1930
rect 1231 1926 1323 1930
rect 1327 1926 1371 1930
rect 1375 1926 1483 1930
rect 1487 1926 1515 1930
rect 1519 1926 1643 1930
rect 1647 1926 1651 1930
rect 1655 1926 1787 1930
rect 1791 1926 1935 1930
rect 1939 1926 1959 1930
rect 103 1925 1959 1926
rect 1965 1925 1966 1931
rect 1972 1930 3811 1931
rect 1972 1926 1975 1930
rect 1979 1926 2023 1930
rect 2027 1926 2183 1930
rect 2187 1926 2415 1930
rect 2419 1926 2695 1930
rect 2699 1926 3015 1930
rect 3019 1926 3135 1930
rect 3139 1926 3271 1930
rect 3275 1926 3359 1930
rect 3363 1926 3407 1930
rect 3411 1926 3543 1930
rect 3547 1926 3679 1930
rect 3683 1926 3799 1930
rect 3803 1926 3811 1930
rect 1972 1925 3811 1926
rect 3817 1925 3818 1931
rect 3810 1837 3811 1843
rect 3817 1842 5695 1843
rect 3817 1838 3839 1842
rect 3843 1838 3887 1842
rect 3891 1838 4071 1842
rect 4075 1838 4311 1842
rect 4315 1838 4407 1842
rect 4411 1838 4543 1842
rect 4547 1838 4591 1842
rect 4595 1838 4679 1842
rect 4683 1838 4815 1842
rect 4819 1838 4903 1842
rect 4907 1838 4951 1842
rect 4955 1838 5231 1842
rect 5235 1838 5543 1842
rect 5547 1838 5663 1842
rect 5667 1838 5695 1842
rect 3817 1837 5695 1838
rect 5701 1837 5702 1843
rect 84 1801 85 1807
rect 91 1806 1947 1807
rect 91 1802 111 1806
rect 115 1802 223 1806
rect 227 1802 263 1806
rect 267 1802 463 1806
rect 467 1802 655 1806
rect 659 1802 695 1806
rect 699 1802 839 1806
rect 843 1802 927 1806
rect 931 1802 1015 1806
rect 1019 1802 1159 1806
rect 1163 1802 1183 1806
rect 1187 1802 1351 1806
rect 1355 1802 1391 1806
rect 1395 1802 1511 1806
rect 1515 1802 1671 1806
rect 1675 1802 1815 1806
rect 1819 1802 1935 1806
rect 1939 1802 1947 1806
rect 91 1801 1947 1802
rect 1953 1801 1954 1807
rect 1958 1801 1959 1807
rect 1965 1806 3823 1807
rect 1965 1802 1975 1806
rect 1979 1802 1995 1806
rect 1999 1802 2131 1806
rect 2135 1802 2267 1806
rect 2271 1802 2419 1806
rect 2423 1802 2579 1806
rect 2583 1802 2739 1806
rect 2743 1802 2899 1806
rect 2903 1802 3051 1806
rect 3055 1802 3107 1806
rect 3111 1802 3203 1806
rect 3207 1802 3243 1806
rect 3247 1802 3355 1806
rect 3359 1802 3379 1806
rect 3383 1802 3515 1806
rect 3519 1802 3651 1806
rect 3655 1802 3799 1806
rect 3803 1802 3823 1806
rect 1965 1801 3823 1802
rect 3829 1801 3830 1807
rect 3022 1788 3028 1789
rect 3770 1788 3776 1789
rect 3022 1784 3023 1788
rect 3027 1784 3771 1788
rect 3775 1784 3776 1788
rect 3022 1783 3028 1784
rect 3770 1783 3776 1784
rect 3822 1709 3823 1715
rect 3829 1714 5707 1715
rect 3829 1710 3839 1714
rect 3843 1710 4379 1714
rect 4383 1710 4515 1714
rect 4519 1710 4563 1714
rect 4567 1710 4651 1714
rect 4655 1710 4699 1714
rect 4703 1710 4787 1714
rect 4791 1710 4835 1714
rect 4839 1710 4923 1714
rect 4927 1710 4971 1714
rect 4975 1710 5107 1714
rect 5111 1710 5243 1714
rect 5247 1710 5379 1714
rect 5383 1710 5515 1714
rect 5519 1710 5663 1714
rect 5667 1710 5707 1714
rect 3829 1709 5707 1710
rect 5713 1709 5714 1715
rect 1946 1687 1947 1693
rect 1953 1687 1978 1693
rect 1972 1683 1978 1687
rect 96 1677 97 1683
rect 103 1682 1959 1683
rect 103 1678 111 1682
rect 115 1678 131 1682
rect 135 1678 195 1682
rect 199 1678 363 1682
rect 367 1678 435 1682
rect 439 1678 619 1682
rect 623 1678 667 1682
rect 671 1678 875 1682
rect 879 1678 899 1682
rect 903 1678 1131 1682
rect 1135 1678 1139 1682
rect 1143 1678 1363 1682
rect 1367 1678 1935 1682
rect 1939 1678 1959 1682
rect 103 1677 1959 1678
rect 1965 1677 1966 1683
rect 1972 1682 3811 1683
rect 1972 1678 1975 1682
rect 1979 1678 2023 1682
rect 2027 1678 2159 1682
rect 2163 1678 2167 1682
rect 2171 1678 2295 1682
rect 2299 1678 2319 1682
rect 2323 1678 2447 1682
rect 2451 1678 2479 1682
rect 2483 1678 2607 1682
rect 2611 1678 2639 1682
rect 2643 1678 2767 1682
rect 2771 1678 2791 1682
rect 2795 1678 2927 1682
rect 2931 1678 2943 1682
rect 2947 1678 3079 1682
rect 3083 1678 3103 1682
rect 3107 1678 3231 1682
rect 3235 1678 3263 1682
rect 3267 1678 3383 1682
rect 3387 1678 3423 1682
rect 3427 1678 3543 1682
rect 3547 1678 3679 1682
rect 3683 1678 3799 1682
rect 3803 1678 3811 1682
rect 1972 1677 3811 1678
rect 3817 1677 3818 1683
rect 3810 1581 3811 1587
rect 3817 1586 5695 1587
rect 3817 1582 3839 1586
rect 3843 1582 4591 1586
rect 4595 1582 4727 1586
rect 4731 1582 4863 1586
rect 4867 1582 4999 1586
rect 5003 1582 5135 1586
rect 5139 1582 5271 1586
rect 5275 1582 5407 1586
rect 5411 1582 5543 1586
rect 5547 1582 5663 1586
rect 5667 1582 5695 1586
rect 3817 1581 5695 1582
rect 5701 1581 5702 1587
rect 84 1553 85 1559
rect 91 1558 1947 1559
rect 91 1554 111 1558
rect 115 1554 159 1558
rect 163 1554 327 1558
rect 331 1554 391 1558
rect 395 1554 511 1558
rect 515 1554 647 1558
rect 651 1554 695 1558
rect 699 1554 887 1558
rect 891 1554 903 1558
rect 907 1554 1079 1558
rect 1083 1554 1167 1558
rect 1171 1554 1935 1558
rect 1939 1554 1947 1558
rect 91 1553 1947 1554
rect 1953 1553 1954 1559
rect 1958 1553 1959 1559
rect 1965 1558 3823 1559
rect 1965 1554 1975 1558
rect 1979 1554 1995 1558
rect 1999 1554 2131 1558
rect 2135 1554 2139 1558
rect 2143 1554 2267 1558
rect 2271 1554 2291 1558
rect 2295 1554 2403 1558
rect 2407 1554 2451 1558
rect 2455 1554 2539 1558
rect 2543 1554 2611 1558
rect 2615 1554 2675 1558
rect 2679 1554 2763 1558
rect 2767 1554 2811 1558
rect 2815 1554 2915 1558
rect 2919 1554 2947 1558
rect 2951 1554 3075 1558
rect 3079 1554 3083 1558
rect 3087 1554 3219 1558
rect 3223 1554 3235 1558
rect 3239 1554 3355 1558
rect 3359 1554 3395 1558
rect 3399 1554 3491 1558
rect 3495 1554 3799 1558
rect 3803 1554 3823 1558
rect 1965 1553 3823 1554
rect 3829 1553 3830 1559
rect 1946 1439 1947 1445
rect 1953 1439 1978 1445
rect 1972 1435 1978 1439
rect 96 1429 97 1435
rect 103 1434 1959 1435
rect 103 1430 111 1434
rect 115 1430 131 1434
rect 135 1430 299 1434
rect 303 1430 395 1434
rect 399 1430 483 1434
rect 487 1430 667 1434
rect 671 1430 683 1434
rect 687 1430 859 1434
rect 863 1430 971 1434
rect 975 1430 1051 1434
rect 1055 1430 1259 1434
rect 1263 1430 1935 1434
rect 1939 1430 1959 1434
rect 103 1429 1959 1430
rect 1965 1429 1966 1435
rect 1972 1434 3811 1435
rect 1972 1430 1975 1434
rect 1979 1430 2023 1434
rect 2027 1430 2159 1434
rect 2163 1430 2167 1434
rect 2171 1430 2295 1434
rect 2299 1430 2303 1434
rect 2307 1430 2431 1434
rect 2435 1430 2439 1434
rect 2443 1430 2567 1434
rect 2571 1430 2575 1434
rect 2579 1430 2703 1434
rect 2707 1430 2711 1434
rect 2715 1430 2839 1434
rect 2843 1430 2847 1434
rect 2851 1430 2975 1434
rect 2979 1430 2983 1434
rect 2987 1430 3111 1434
rect 3115 1430 3119 1434
rect 3123 1430 3247 1434
rect 3251 1430 3255 1434
rect 3259 1430 3383 1434
rect 3387 1430 3519 1434
rect 3523 1430 3799 1434
rect 3803 1430 3811 1434
rect 1972 1429 3811 1430
rect 3817 1429 3818 1435
rect 3822 1397 3823 1403
rect 3829 1402 5707 1403
rect 3829 1398 3839 1402
rect 3843 1398 4563 1402
rect 4567 1398 4699 1402
rect 4703 1398 4811 1402
rect 4815 1398 4835 1402
rect 4839 1398 4947 1402
rect 4951 1398 4971 1402
rect 4975 1398 5083 1402
rect 5087 1398 5107 1402
rect 5111 1398 5219 1402
rect 5223 1398 5243 1402
rect 5247 1398 5355 1402
rect 5359 1398 5379 1402
rect 5383 1398 5491 1402
rect 5495 1398 5515 1402
rect 5519 1398 5663 1402
rect 5667 1398 5707 1402
rect 3829 1397 5707 1398
rect 5713 1397 5714 1403
rect 84 1317 85 1323
rect 91 1322 1947 1323
rect 91 1318 111 1322
rect 115 1318 159 1322
rect 163 1318 423 1322
rect 427 1318 455 1322
rect 459 1318 711 1322
rect 715 1318 775 1322
rect 779 1318 999 1322
rect 1003 1318 1095 1322
rect 1099 1318 1287 1322
rect 1291 1318 1423 1322
rect 1427 1318 1935 1322
rect 1939 1318 1947 1322
rect 91 1317 1947 1318
rect 1953 1317 1954 1323
rect 1958 1317 1959 1323
rect 1965 1322 3823 1323
rect 1965 1318 1975 1322
rect 1979 1318 2131 1322
rect 2135 1318 2139 1322
rect 2143 1318 2267 1322
rect 2271 1318 2275 1322
rect 2279 1318 2403 1322
rect 2407 1318 2411 1322
rect 2415 1318 2547 1322
rect 2551 1318 2555 1322
rect 2559 1318 2683 1322
rect 2687 1318 2715 1322
rect 2719 1318 2819 1322
rect 2823 1318 2891 1322
rect 2895 1318 2955 1322
rect 2959 1318 3075 1322
rect 3079 1318 3091 1322
rect 3095 1318 3227 1322
rect 3231 1318 3267 1322
rect 3271 1318 3467 1322
rect 3471 1318 3651 1322
rect 3655 1318 3799 1322
rect 3803 1318 3823 1322
rect 1965 1317 3823 1318
rect 3829 1317 3830 1323
rect 2498 1300 2504 1301
rect 2722 1300 2728 1301
rect 2498 1296 2499 1300
rect 2503 1296 2723 1300
rect 2727 1296 2728 1300
rect 2498 1295 2504 1296
rect 2722 1295 2728 1296
rect 3810 1281 3811 1287
rect 3817 1286 5695 1287
rect 3817 1282 3839 1286
rect 3843 1282 4735 1286
rect 4739 1282 4839 1286
rect 4843 1282 4879 1286
rect 4883 1282 4975 1286
rect 4979 1282 5031 1286
rect 5035 1282 5111 1286
rect 5115 1282 5191 1286
rect 5195 1282 5247 1286
rect 5251 1282 5359 1286
rect 5363 1282 5383 1286
rect 5387 1282 5519 1286
rect 5523 1282 5527 1286
rect 5531 1282 5663 1286
rect 5667 1282 5695 1286
rect 3817 1281 5695 1282
rect 5701 1281 5702 1287
rect 1946 1205 1947 1211
rect 1953 1210 3811 1211
rect 1953 1206 1975 1210
rect 1979 1206 2023 1210
rect 2027 1206 2159 1210
rect 2163 1206 2239 1210
rect 2243 1206 2295 1210
rect 2299 1206 2431 1210
rect 2435 1206 2479 1210
rect 2483 1206 2583 1210
rect 2587 1206 2719 1210
rect 2723 1206 2743 1210
rect 2747 1206 2919 1210
rect 2923 1206 2959 1210
rect 2963 1206 3103 1210
rect 3107 1206 3207 1210
rect 3211 1206 3295 1210
rect 3299 1206 3455 1210
rect 3459 1206 3495 1210
rect 3499 1206 3679 1210
rect 3683 1206 3799 1210
rect 3803 1206 3811 1210
rect 1953 1205 3811 1206
rect 3817 1205 3818 1211
rect 96 1181 97 1187
rect 103 1186 1959 1187
rect 103 1182 111 1186
rect 115 1182 131 1186
rect 135 1182 331 1186
rect 335 1182 427 1186
rect 431 1182 563 1186
rect 567 1182 747 1186
rect 751 1182 803 1186
rect 807 1182 1043 1186
rect 1047 1182 1067 1186
rect 1071 1182 1283 1186
rect 1287 1182 1395 1186
rect 1399 1182 1523 1186
rect 1527 1182 1771 1186
rect 1775 1182 1935 1186
rect 1939 1182 1959 1186
rect 103 1181 1959 1182
rect 1965 1181 1966 1187
rect 3822 1161 3823 1167
rect 3829 1166 5707 1167
rect 3829 1162 3839 1166
rect 3843 1162 3859 1166
rect 3863 1162 4067 1166
rect 4071 1162 4299 1166
rect 4303 1162 4539 1166
rect 4543 1162 4707 1166
rect 4711 1162 4779 1166
rect 4783 1162 4851 1166
rect 4855 1162 5003 1166
rect 5007 1162 5027 1166
rect 5031 1162 5163 1166
rect 5167 1162 5283 1166
rect 5287 1162 5331 1166
rect 5335 1162 5499 1166
rect 5503 1162 5515 1166
rect 5519 1162 5663 1166
rect 5667 1162 5707 1166
rect 3829 1161 5707 1162
rect 5713 1161 5714 1167
rect 84 1069 85 1075
rect 91 1074 1947 1075
rect 91 1070 111 1074
rect 115 1070 159 1074
rect 163 1070 263 1074
rect 267 1070 359 1074
rect 363 1070 439 1074
rect 443 1070 591 1074
rect 595 1070 615 1074
rect 619 1070 783 1074
rect 787 1070 831 1074
rect 835 1070 951 1074
rect 955 1070 1071 1074
rect 1075 1070 1111 1074
rect 1115 1070 1271 1074
rect 1275 1070 1311 1074
rect 1315 1070 1431 1074
rect 1435 1070 1551 1074
rect 1555 1070 1591 1074
rect 1595 1070 1751 1074
rect 1755 1070 1799 1074
rect 1803 1070 1935 1074
rect 1939 1070 1947 1074
rect 91 1069 1947 1070
rect 1953 1069 1954 1075
rect 1958 1069 1959 1075
rect 1965 1074 3823 1075
rect 1965 1070 1975 1074
rect 1979 1070 1995 1074
rect 1999 1070 2211 1074
rect 2215 1070 2451 1074
rect 2455 1070 2691 1074
rect 2695 1070 2931 1074
rect 2935 1070 3091 1074
rect 3095 1070 3179 1074
rect 3183 1070 3243 1074
rect 3247 1070 3395 1074
rect 3399 1070 3427 1074
rect 3431 1070 3651 1074
rect 3655 1070 3799 1074
rect 3803 1070 3823 1074
rect 1965 1069 3823 1070
rect 3829 1069 3830 1075
rect 3810 1049 3811 1055
rect 3817 1054 5695 1055
rect 3817 1050 3839 1054
rect 3843 1050 3887 1054
rect 3891 1050 4071 1054
rect 4075 1050 4095 1054
rect 4099 1050 4279 1054
rect 4283 1050 4327 1054
rect 4331 1050 4511 1054
rect 4515 1050 4567 1054
rect 4571 1050 4759 1054
rect 4763 1050 4807 1054
rect 4811 1050 5023 1054
rect 5027 1050 5055 1054
rect 5059 1050 5295 1054
rect 5299 1050 5311 1054
rect 5315 1050 5543 1054
rect 5547 1050 5663 1054
rect 5667 1050 5695 1054
rect 3817 1049 5695 1050
rect 5701 1049 5702 1055
rect 96 953 97 959
rect 103 958 1959 959
rect 103 954 111 958
rect 115 954 227 958
rect 231 954 235 958
rect 239 954 379 958
rect 383 954 411 958
rect 415 954 539 958
rect 543 954 587 958
rect 591 954 715 958
rect 719 954 755 958
rect 759 954 891 958
rect 895 954 923 958
rect 927 954 1075 958
rect 1079 954 1083 958
rect 1087 954 1243 958
rect 1247 954 1259 958
rect 1263 954 1403 958
rect 1407 954 1443 958
rect 1447 954 1563 958
rect 1567 954 1627 958
rect 1631 954 1723 958
rect 1727 954 1787 958
rect 1791 954 1935 958
rect 1939 954 1959 958
rect 103 953 1959 954
rect 1965 953 1966 959
rect 3822 937 3823 943
rect 3829 942 5707 943
rect 3829 938 3839 942
rect 3843 938 3859 942
rect 3863 938 3971 942
rect 3975 938 4043 942
rect 4047 938 4179 942
rect 4183 938 4251 942
rect 4255 938 4403 942
rect 4407 938 4483 942
rect 4487 938 4643 942
rect 4647 938 4731 942
rect 4735 938 4899 942
rect 4903 938 4995 942
rect 4999 938 5171 942
rect 5175 938 5267 942
rect 5271 938 5443 942
rect 5447 938 5515 942
rect 5519 938 5663 942
rect 5667 938 5707 942
rect 3829 937 5707 938
rect 5713 937 5714 943
rect 1946 929 1947 935
rect 1953 934 3811 935
rect 1953 930 1975 934
rect 1979 930 2047 934
rect 2051 930 2351 934
rect 2355 930 2647 934
rect 2651 930 2927 934
rect 2931 930 3119 934
rect 3123 930 3207 934
rect 3211 930 3271 934
rect 3275 930 3423 934
rect 3427 930 3495 934
rect 3499 930 3799 934
rect 3803 930 3811 934
rect 1953 929 3811 930
rect 3817 929 3818 935
rect 84 825 85 831
rect 91 830 1947 831
rect 91 826 111 830
rect 115 826 255 830
rect 259 826 375 830
rect 379 826 407 830
rect 411 826 567 830
rect 571 826 655 830
rect 659 826 743 830
rect 747 826 919 830
rect 923 826 943 830
rect 947 826 1103 830
rect 1107 826 1239 830
rect 1243 826 1287 830
rect 1291 826 1471 830
rect 1475 826 1535 830
rect 1539 826 1655 830
rect 1659 826 1815 830
rect 1819 826 1935 830
rect 1939 826 1947 830
rect 91 825 1947 826
rect 1953 825 1954 831
rect 3810 827 3811 833
rect 3817 831 3842 833
rect 3817 830 5695 831
rect 3817 827 3839 830
rect 3836 826 3839 827
rect 3843 826 3887 830
rect 3891 826 3999 830
rect 4003 826 4047 830
rect 4051 826 4207 830
rect 4211 826 4279 830
rect 4283 826 4431 830
rect 4435 826 4559 830
rect 4563 826 4671 830
rect 4675 826 4879 830
rect 4883 826 4927 830
rect 4931 826 5199 830
rect 5203 826 5223 830
rect 5227 826 5471 830
rect 5475 826 5543 830
rect 5547 826 5663 830
rect 5667 826 5695 830
rect 3836 825 5695 826
rect 5701 825 5702 831
rect 1958 817 1959 823
rect 1965 822 3823 823
rect 1965 818 1975 822
rect 1979 818 1995 822
rect 1999 818 2019 822
rect 2023 818 2251 822
rect 2255 818 2323 822
rect 2327 818 2523 822
rect 2527 818 2619 822
rect 2623 818 2771 822
rect 2775 818 2899 822
rect 2903 818 3003 822
rect 3007 818 3179 822
rect 3183 818 3227 822
rect 3231 818 3451 822
rect 3455 818 3467 822
rect 3471 818 3651 822
rect 3655 818 3799 822
rect 3803 818 3823 822
rect 1965 817 3823 818
rect 3829 817 3830 823
rect 96 713 97 719
rect 103 718 1959 719
rect 103 714 111 718
rect 115 714 131 718
rect 135 714 307 718
rect 311 714 347 718
rect 351 714 499 718
rect 503 714 627 718
rect 631 714 683 718
rect 687 714 859 718
rect 863 714 915 718
rect 919 714 1027 718
rect 1031 714 1187 718
rect 1191 714 1211 718
rect 1215 714 1339 718
rect 1343 714 1491 718
rect 1495 714 1507 718
rect 1511 714 1651 718
rect 1655 714 1787 718
rect 1791 714 1935 718
rect 1939 714 1959 718
rect 103 713 1959 714
rect 1965 713 1966 719
rect 3822 705 3823 711
rect 3829 710 5707 711
rect 3829 706 3839 710
rect 3843 706 3859 710
rect 3863 706 3995 710
rect 3999 706 4019 710
rect 4023 706 4131 710
rect 4135 706 4251 710
rect 4255 706 4267 710
rect 4271 706 4403 710
rect 4407 706 4531 710
rect 4535 706 4571 710
rect 4575 706 4771 710
rect 4775 706 4851 710
rect 4855 706 4995 710
rect 4999 706 5195 710
rect 5199 706 5227 710
rect 5231 706 5459 710
rect 5463 706 5515 710
rect 5519 706 5663 710
rect 5667 706 5707 710
rect 3829 705 5707 706
rect 5713 705 5714 711
rect 84 601 85 607
rect 91 606 1947 607
rect 91 602 111 606
rect 115 602 159 606
rect 163 602 335 606
rect 339 602 375 606
rect 379 602 527 606
rect 531 602 599 606
rect 603 602 711 606
rect 715 602 807 606
rect 811 602 887 606
rect 891 602 999 606
rect 1003 602 1055 606
rect 1059 602 1175 606
rect 1179 602 1215 606
rect 1219 602 1343 606
rect 1347 602 1367 606
rect 1371 602 1511 606
rect 1515 602 1519 606
rect 1523 602 1671 606
rect 1675 602 1679 606
rect 1683 602 1815 606
rect 1819 602 1935 606
rect 1939 602 1947 606
rect 91 601 1947 602
rect 1953 601 1954 607
rect 3810 593 3811 599
rect 3817 598 5695 599
rect 3817 594 3839 598
rect 3843 594 3887 598
rect 3891 594 4023 598
rect 4027 594 4159 598
rect 4163 594 4295 598
rect 4299 594 4431 598
rect 4435 594 4479 598
rect 4483 594 4599 598
rect 4603 594 4695 598
rect 4699 594 4799 598
rect 4803 594 4935 598
rect 4939 594 5023 598
rect 5027 594 5191 598
rect 5195 594 5255 598
rect 5259 594 5447 598
rect 5451 594 5487 598
rect 5491 594 5663 598
rect 5667 594 5695 598
rect 3817 593 5695 594
rect 5701 593 5702 599
rect 1946 573 1947 579
rect 1953 578 3811 579
rect 1953 574 1975 578
rect 1979 574 2023 578
rect 2027 574 2279 578
rect 2283 574 2551 578
rect 2555 574 2799 578
rect 2803 574 3031 578
rect 3035 574 3255 578
rect 3259 574 3311 578
rect 3315 574 3447 578
rect 3451 574 3479 578
rect 3483 574 3583 578
rect 3587 574 3679 578
rect 3683 574 3799 578
rect 3803 574 3811 578
rect 1953 573 3811 574
rect 3817 573 3818 579
rect 96 489 97 495
rect 103 494 1959 495
rect 103 490 111 494
rect 115 490 131 494
rect 135 490 347 494
rect 351 490 427 494
rect 431 490 571 494
rect 575 490 763 494
rect 767 490 779 494
rect 783 490 971 494
rect 975 490 1107 494
rect 1111 490 1147 494
rect 1151 490 1315 494
rect 1319 490 1459 494
rect 1463 490 1483 494
rect 1487 490 1643 494
rect 1647 490 1787 494
rect 1791 490 1935 494
rect 1939 490 1959 494
rect 103 489 1959 490
rect 1965 489 1966 495
rect 3822 469 3823 475
rect 3829 474 5707 475
rect 3829 470 3839 474
rect 3843 470 3859 474
rect 3863 470 3995 474
rect 3999 470 4131 474
rect 4135 470 4267 474
rect 4271 470 4451 474
rect 4455 470 4651 474
rect 4655 470 4667 474
rect 4671 470 4859 474
rect 4863 470 4907 474
rect 4911 470 5067 474
rect 5071 470 5163 474
rect 5167 470 5283 474
rect 5287 470 5419 474
rect 5423 470 5507 474
rect 5511 470 5663 474
rect 5667 470 5707 474
rect 3829 469 5707 470
rect 5713 469 5714 475
rect 3822 467 3830 469
rect 1958 461 1959 467
rect 1965 466 3823 467
rect 1965 462 1975 466
rect 1979 462 1995 466
rect 1999 462 2155 466
rect 2159 462 2347 466
rect 2351 462 2539 466
rect 2543 462 2731 466
rect 2735 462 2923 466
rect 2927 462 3115 466
rect 3119 462 3283 466
rect 3287 462 3299 466
rect 3303 462 3419 466
rect 3423 462 3483 466
rect 3487 462 3555 466
rect 3559 462 3651 466
rect 3655 462 3799 466
rect 3803 462 3823 466
rect 1965 461 3823 462
rect 3829 461 3830 467
rect 84 361 85 367
rect 91 366 1947 367
rect 91 362 111 366
rect 115 362 159 366
rect 163 362 239 366
rect 243 362 391 366
rect 395 362 455 366
rect 459 362 551 366
rect 555 362 711 366
rect 715 362 791 366
rect 795 362 871 366
rect 875 362 1031 366
rect 1035 362 1135 366
rect 1139 362 1487 366
rect 1491 362 1815 366
rect 1819 362 1935 366
rect 1939 362 1947 366
rect 91 361 1947 362
rect 1953 361 1954 367
rect 3810 353 3811 359
rect 3817 358 5695 359
rect 3817 354 3839 358
rect 3843 354 4479 358
rect 4483 354 4679 358
rect 4683 354 4751 358
rect 4755 354 4887 358
rect 4891 354 4911 358
rect 4915 354 5071 358
rect 5075 354 5095 358
rect 5099 354 5231 358
rect 5235 354 5311 358
rect 5315 354 5399 358
rect 5403 354 5535 358
rect 5539 354 5543 358
rect 5547 354 5663 358
rect 5667 354 5695 358
rect 3817 353 5695 354
rect 5701 353 5702 359
rect 1946 325 1947 331
rect 1953 330 3811 331
rect 1953 326 1975 330
rect 1979 326 2023 330
rect 2027 326 2047 330
rect 2051 326 2183 330
rect 2187 326 2319 330
rect 2323 326 2375 330
rect 2379 326 2455 330
rect 2459 326 2567 330
rect 2571 326 2591 330
rect 2595 326 2727 330
rect 2731 326 2759 330
rect 2763 326 2863 330
rect 2867 326 2951 330
rect 2955 326 2999 330
rect 3003 326 3135 330
rect 3139 326 3143 330
rect 3147 326 3271 330
rect 3275 326 3327 330
rect 3331 326 3407 330
rect 3411 326 3511 330
rect 3515 326 3543 330
rect 3547 326 3679 330
rect 3683 326 3799 330
rect 3803 326 3811 330
rect 1953 325 3811 326
rect 3817 325 3818 331
rect 96 217 97 223
rect 103 222 1959 223
rect 103 218 111 222
rect 115 218 147 222
rect 151 218 211 222
rect 215 218 283 222
rect 287 218 363 222
rect 367 218 419 222
rect 423 218 523 222
rect 527 218 555 222
rect 559 218 683 222
rect 687 218 691 222
rect 695 218 827 222
rect 831 218 843 222
rect 847 218 963 222
rect 967 218 1003 222
rect 1007 218 1099 222
rect 1103 218 1935 222
rect 1939 218 1959 222
rect 103 217 1959 218
rect 1965 217 1966 223
rect 3822 206 5714 207
rect 3822 203 3839 206
rect 1958 197 1959 203
rect 1965 202 3823 203
rect 1965 198 1975 202
rect 1979 198 1995 202
rect 1999 198 2019 202
rect 2023 198 2131 202
rect 2135 198 2155 202
rect 2159 198 2267 202
rect 2271 198 2291 202
rect 2295 198 2403 202
rect 2407 198 2427 202
rect 2431 198 2539 202
rect 2543 198 2563 202
rect 2567 198 2675 202
rect 2679 198 2699 202
rect 2703 198 2811 202
rect 2815 198 2835 202
rect 2839 198 2947 202
rect 2951 198 2971 202
rect 2975 198 3083 202
rect 3087 198 3107 202
rect 3111 198 3219 202
rect 3223 198 3243 202
rect 3247 198 3355 202
rect 3359 198 3379 202
rect 3383 198 3491 202
rect 3495 198 3515 202
rect 3519 198 3627 202
rect 3631 198 3651 202
rect 3655 198 3799 202
rect 3803 198 3823 202
rect 1965 197 3823 198
rect 3829 202 3839 203
rect 3843 202 4291 206
rect 4295 202 4427 206
rect 4431 202 4563 206
rect 4567 202 4699 206
rect 4703 202 4723 206
rect 4727 202 4835 206
rect 4839 202 4883 206
rect 4887 202 4971 206
rect 4975 202 5043 206
rect 5047 202 5107 206
rect 5111 202 5203 206
rect 5207 202 5243 206
rect 5247 202 5371 206
rect 5375 202 5379 206
rect 5383 202 5515 206
rect 5519 202 5663 206
rect 5667 202 5714 206
rect 3829 201 5714 202
rect 3829 197 3830 201
rect 84 105 85 111
rect 91 110 1947 111
rect 91 106 111 110
rect 115 106 175 110
rect 179 106 311 110
rect 315 106 447 110
rect 451 106 583 110
rect 587 106 719 110
rect 723 106 855 110
rect 859 106 991 110
rect 995 106 1127 110
rect 1131 106 1935 110
rect 1939 106 1947 110
rect 91 105 1947 106
rect 1953 105 1954 111
rect 3810 94 5702 95
rect 3810 91 3839 94
rect 1946 85 1947 91
rect 1953 90 3811 91
rect 1953 86 1975 90
rect 1979 86 2023 90
rect 2027 86 2159 90
rect 2163 86 2295 90
rect 2299 86 2431 90
rect 2435 86 2567 90
rect 2571 86 2703 90
rect 2707 86 2839 90
rect 2843 86 2975 90
rect 2979 86 3111 90
rect 3115 86 3247 90
rect 3251 86 3383 90
rect 3387 86 3519 90
rect 3523 86 3655 90
rect 3659 86 3799 90
rect 3803 86 3811 90
rect 1953 85 3811 86
rect 3817 90 3839 91
rect 3843 90 4319 94
rect 4323 90 4455 94
rect 4459 90 4591 94
rect 4595 90 4727 94
rect 4731 90 4863 94
rect 4867 90 4999 94
rect 5003 90 5135 94
rect 5139 90 5271 94
rect 5275 90 5407 94
rect 5411 90 5543 94
rect 5547 90 5663 94
rect 5667 90 5702 94
rect 3817 89 5702 90
rect 3817 85 3818 89
<< m5c >>
rect 97 5753 103 5759
rect 1959 5753 1965 5759
rect 1959 5685 1965 5691
rect 3823 5685 3829 5691
rect 85 5641 91 5647
rect 1947 5641 1953 5647
rect 1947 5573 1953 5579
rect 3811 5573 3817 5579
rect 97 5529 103 5535
rect 1959 5529 1965 5535
rect 3823 5465 3829 5471
rect 5707 5465 5713 5471
rect 1959 5457 1965 5463
rect 3823 5457 3829 5463
rect 85 5417 91 5423
rect 1947 5417 1953 5423
rect 1947 5345 1953 5351
rect 3811 5345 3817 5351
rect 97 5305 103 5311
rect 1959 5305 1965 5311
rect 1959 5229 1965 5235
rect 3823 5229 3829 5235
rect 3823 5217 3829 5223
rect 5707 5217 5713 5223
rect 85 5193 91 5199
rect 1947 5193 1953 5199
rect 1947 5101 1953 5107
rect 3811 5101 3817 5107
rect 97 5073 103 5079
rect 1959 5073 1965 5079
rect 1959 4981 1965 4987
rect 3823 4981 3829 4987
rect 85 4933 91 4939
rect 1947 4933 1953 4939
rect 1947 4861 1953 4867
rect 3811 4861 3817 4867
rect 97 4809 103 4815
rect 1959 4809 1965 4815
rect 3811 4797 3817 4803
rect 5695 4797 5701 4803
rect 1959 4737 1965 4743
rect 3823 4737 3829 4743
rect 85 4693 91 4699
rect 1947 4693 1953 4699
rect 3823 4685 3829 4691
rect 5707 4685 5713 4691
rect 1947 4621 1953 4627
rect 3811 4621 3817 4627
rect 97 4569 103 4575
rect 1959 4569 1965 4575
rect 3811 4573 3817 4579
rect 5695 4573 5701 4579
rect 1959 4497 1965 4503
rect 3823 4497 3829 4503
rect 85 4457 91 4463
rect 1947 4457 1953 4463
rect 3823 4457 3829 4463
rect 5707 4457 5713 4463
rect 1947 4373 1953 4379
rect 3811 4373 3817 4379
rect 97 4341 103 4347
rect 1959 4341 1965 4347
rect 3811 4329 3817 4335
rect 5695 4329 5701 4335
rect 1959 4257 1965 4263
rect 3823 4257 3829 4263
rect 85 4221 91 4227
rect 1947 4221 1953 4227
rect 3823 4205 3829 4211
rect 5707 4205 5713 4211
rect 1947 4133 1953 4139
rect 3811 4133 3817 4139
rect 97 4109 103 4115
rect 1959 4109 1965 4115
rect 3811 4069 3817 4075
rect 5695 4069 5701 4075
rect 85 3997 91 4003
rect 1947 3997 1953 4003
rect 3823 3957 3829 3963
rect 5707 3957 5713 3963
rect 1959 3929 1965 3935
rect 3823 3929 3829 3935
rect 97 3885 103 3891
rect 1959 3885 1965 3891
rect 1947 3817 1953 3823
rect 3811 3817 3817 3823
rect 85 3761 91 3767
rect 1947 3761 1953 3767
rect 1959 3697 1965 3703
rect 3823 3697 3829 3703
rect 3823 3685 3829 3691
rect 5707 3685 5713 3691
rect 97 3633 103 3639
rect 1959 3633 1965 3639
rect 1947 3577 1953 3583
rect 3811 3577 3817 3583
rect 3811 3525 3817 3531
rect 5695 3525 5701 3531
rect 85 3501 91 3507
rect 1947 3501 1953 3507
rect 1959 3461 1965 3467
rect 3823 3461 3829 3467
rect 3823 3405 3829 3411
rect 5707 3405 5713 3411
rect 97 3381 103 3387
rect 1959 3381 1965 3387
rect 1947 3325 1953 3331
rect 3811 3325 3817 3331
rect 3811 3293 3817 3299
rect 5695 3293 5701 3299
rect 85 3261 91 3267
rect 1947 3261 1953 3267
rect 1959 3213 1965 3219
rect 3823 3213 3829 3219
rect 3823 3165 3829 3171
rect 5707 3165 5713 3171
rect 97 3133 103 3139
rect 1959 3133 1965 3139
rect 1947 3101 1953 3107
rect 3811 3101 3817 3107
rect 3811 3053 3817 3059
rect 5695 3053 5701 3059
rect 85 3021 91 3027
rect 1947 3021 1953 3027
rect 1959 2989 1965 2995
rect 3823 2989 3829 2995
rect 3823 2917 3829 2923
rect 5707 2917 5713 2923
rect 97 2905 103 2911
rect 1959 2905 1965 2911
rect 1947 2825 1953 2831
rect 3811 2825 3817 2831
rect 3811 2801 3817 2807
rect 5695 2801 5701 2807
rect 85 2781 91 2787
rect 1947 2781 1953 2787
rect 1959 2713 1965 2719
rect 3823 2713 3829 2719
rect 3823 2677 3829 2683
rect 5707 2677 5713 2683
rect 97 2669 103 2675
rect 1959 2669 1965 2675
rect 1947 2597 1953 2603
rect 3811 2597 3817 2603
rect 3811 2561 3817 2567
rect 5695 2561 5701 2567
rect 85 2541 91 2547
rect 1947 2541 1953 2547
rect 1959 2469 1965 2475
rect 3823 2469 3829 2475
rect 3823 2433 3829 2439
rect 5707 2433 5713 2439
rect 97 2417 103 2423
rect 1959 2417 1965 2423
rect 1947 2349 1953 2355
rect 3811 2349 3817 2355
rect 3811 2309 3817 2315
rect 5695 2309 5701 2315
rect 85 2301 91 2307
rect 1947 2301 1953 2307
rect 1959 2237 1965 2243
rect 3823 2237 3829 2243
rect 3823 2193 3829 2199
rect 5707 2193 5713 2199
rect 97 2165 103 2171
rect 1959 2165 1965 2171
rect 3811 2061 3817 2067
rect 5695 2061 5701 2067
rect 85 2049 91 2055
rect 1947 2049 1953 2055
rect 3823 1949 3829 1955
rect 5707 1949 5713 1955
rect 1947 1935 1953 1941
rect 97 1925 103 1931
rect 1959 1925 1965 1931
rect 3811 1925 3817 1931
rect 3811 1837 3817 1843
rect 5695 1837 5701 1843
rect 85 1801 91 1807
rect 1947 1801 1953 1807
rect 1959 1801 1965 1807
rect 3823 1801 3829 1807
rect 3823 1709 3829 1715
rect 5707 1709 5713 1715
rect 1947 1687 1953 1693
rect 97 1677 103 1683
rect 1959 1677 1965 1683
rect 3811 1677 3817 1683
rect 3811 1581 3817 1587
rect 5695 1581 5701 1587
rect 85 1553 91 1559
rect 1947 1553 1953 1559
rect 1959 1553 1965 1559
rect 3823 1553 3829 1559
rect 1947 1439 1953 1445
rect 97 1429 103 1435
rect 1959 1429 1965 1435
rect 3811 1429 3817 1435
rect 3823 1397 3829 1403
rect 5707 1397 5713 1403
rect 85 1317 91 1323
rect 1947 1317 1953 1323
rect 1959 1317 1965 1323
rect 3823 1317 3829 1323
rect 3811 1281 3817 1287
rect 5695 1281 5701 1287
rect 1947 1205 1953 1211
rect 3811 1205 3817 1211
rect 97 1181 103 1187
rect 1959 1181 1965 1187
rect 3823 1161 3829 1167
rect 5707 1161 5713 1167
rect 85 1069 91 1075
rect 1947 1069 1953 1075
rect 1959 1069 1965 1075
rect 3823 1069 3829 1075
rect 3811 1049 3817 1055
rect 5695 1049 5701 1055
rect 97 953 103 959
rect 1959 953 1965 959
rect 3823 937 3829 943
rect 5707 937 5713 943
rect 1947 929 1953 935
rect 3811 929 3817 935
rect 85 825 91 831
rect 1947 825 1953 831
rect 3811 827 3817 833
rect 5695 825 5701 831
rect 1959 817 1965 823
rect 3823 817 3829 823
rect 97 713 103 719
rect 1959 713 1965 719
rect 3823 705 3829 711
rect 5707 705 5713 711
rect 85 601 91 607
rect 1947 601 1953 607
rect 3811 593 3817 599
rect 5695 593 5701 599
rect 1947 573 1953 579
rect 3811 573 3817 579
rect 97 489 103 495
rect 1959 489 1965 495
rect 3823 469 3829 475
rect 5707 469 5713 475
rect 1959 461 1965 467
rect 3823 461 3829 467
rect 85 361 91 367
rect 1947 361 1953 367
rect 3811 353 3817 359
rect 5695 353 5701 359
rect 1947 325 1953 331
rect 3811 325 3817 331
rect 97 217 103 223
rect 1959 217 1965 223
rect 1959 197 1965 203
rect 3823 197 3829 203
rect 85 105 91 111
rect 1947 105 1953 111
rect 1947 85 1953 91
rect 3811 85 3817 91
<< m5 >>
rect 84 5647 92 5760
rect 84 5641 85 5647
rect 91 5641 92 5647
rect 84 5423 92 5641
rect 84 5417 85 5423
rect 91 5417 92 5423
rect 84 5199 92 5417
rect 84 5193 85 5199
rect 91 5193 92 5199
rect 84 4939 92 5193
rect 84 4933 85 4939
rect 91 4933 92 4939
rect 84 4699 92 4933
rect 84 4693 85 4699
rect 91 4693 92 4699
rect 84 4463 92 4693
rect 84 4457 85 4463
rect 91 4457 92 4463
rect 84 4227 92 4457
rect 84 4221 85 4227
rect 91 4221 92 4227
rect 84 4003 92 4221
rect 84 3997 85 4003
rect 91 3997 92 4003
rect 84 3767 92 3997
rect 84 3761 85 3767
rect 91 3761 92 3767
rect 84 3507 92 3761
rect 84 3501 85 3507
rect 91 3501 92 3507
rect 84 3267 92 3501
rect 84 3261 85 3267
rect 91 3261 92 3267
rect 84 3027 92 3261
rect 84 3021 85 3027
rect 91 3021 92 3027
rect 84 2787 92 3021
rect 84 2781 85 2787
rect 91 2781 92 2787
rect 84 2547 92 2781
rect 84 2541 85 2547
rect 91 2541 92 2547
rect 84 2307 92 2541
rect 84 2301 85 2307
rect 91 2301 92 2307
rect 84 2055 92 2301
rect 84 2049 85 2055
rect 91 2049 92 2055
rect 84 1807 92 2049
rect 84 1801 85 1807
rect 91 1801 92 1807
rect 84 1559 92 1801
rect 84 1553 85 1559
rect 91 1553 92 1559
rect 84 1323 92 1553
rect 84 1317 85 1323
rect 91 1317 92 1323
rect 84 1075 92 1317
rect 84 1069 85 1075
rect 91 1069 92 1075
rect 84 831 92 1069
rect 84 825 85 831
rect 91 825 92 831
rect 84 607 92 825
rect 84 601 85 607
rect 91 601 92 607
rect 84 367 92 601
rect 84 361 85 367
rect 91 361 92 367
rect 84 111 92 361
rect 84 105 85 111
rect 91 105 92 111
rect 84 72 92 105
rect 96 5759 104 5760
rect 96 5753 97 5759
rect 103 5753 104 5759
rect 96 5535 104 5753
rect 96 5529 97 5535
rect 103 5529 104 5535
rect 96 5311 104 5529
rect 96 5305 97 5311
rect 103 5305 104 5311
rect 96 5079 104 5305
rect 96 5073 97 5079
rect 103 5073 104 5079
rect 96 4815 104 5073
rect 96 4809 97 4815
rect 103 4809 104 4815
rect 96 4575 104 4809
rect 96 4569 97 4575
rect 103 4569 104 4575
rect 96 4347 104 4569
rect 96 4341 97 4347
rect 103 4341 104 4347
rect 96 4115 104 4341
rect 96 4109 97 4115
rect 103 4109 104 4115
rect 96 3891 104 4109
rect 96 3885 97 3891
rect 103 3885 104 3891
rect 96 3639 104 3885
rect 96 3633 97 3639
rect 103 3633 104 3639
rect 96 3387 104 3633
rect 96 3381 97 3387
rect 103 3381 104 3387
rect 96 3139 104 3381
rect 96 3133 97 3139
rect 103 3133 104 3139
rect 96 2911 104 3133
rect 96 2905 97 2911
rect 103 2905 104 2911
rect 96 2675 104 2905
rect 96 2669 97 2675
rect 103 2669 104 2675
rect 96 2423 104 2669
rect 96 2417 97 2423
rect 103 2417 104 2423
rect 96 2171 104 2417
rect 96 2165 97 2171
rect 103 2165 104 2171
rect 96 1931 104 2165
rect 96 1925 97 1931
rect 103 1925 104 1931
rect 96 1683 104 1925
rect 96 1677 97 1683
rect 103 1677 104 1683
rect 96 1435 104 1677
rect 96 1429 97 1435
rect 103 1429 104 1435
rect 96 1187 104 1429
rect 96 1181 97 1187
rect 103 1181 104 1187
rect 96 959 104 1181
rect 96 953 97 959
rect 103 953 104 959
rect 96 719 104 953
rect 96 713 97 719
rect 103 713 104 719
rect 96 495 104 713
rect 96 489 97 495
rect 103 489 104 495
rect 96 223 104 489
rect 96 217 97 223
rect 103 217 104 223
rect 96 72 104 217
rect 1946 5647 1954 5760
rect 1946 5641 1947 5647
rect 1953 5641 1954 5647
rect 1946 5579 1954 5641
rect 1946 5573 1947 5579
rect 1953 5573 1954 5579
rect 1946 5423 1954 5573
rect 1946 5417 1947 5423
rect 1953 5417 1954 5423
rect 1946 5351 1954 5417
rect 1946 5345 1947 5351
rect 1953 5345 1954 5351
rect 1946 5199 1954 5345
rect 1946 5193 1947 5199
rect 1953 5193 1954 5199
rect 1946 5107 1954 5193
rect 1946 5101 1947 5107
rect 1953 5101 1954 5107
rect 1946 4939 1954 5101
rect 1946 4933 1947 4939
rect 1953 4933 1954 4939
rect 1946 4867 1954 4933
rect 1946 4861 1947 4867
rect 1953 4861 1954 4867
rect 1946 4699 1954 4861
rect 1946 4693 1947 4699
rect 1953 4693 1954 4699
rect 1946 4627 1954 4693
rect 1946 4621 1947 4627
rect 1953 4621 1954 4627
rect 1946 4463 1954 4621
rect 1946 4457 1947 4463
rect 1953 4457 1954 4463
rect 1946 4379 1954 4457
rect 1946 4373 1947 4379
rect 1953 4373 1954 4379
rect 1946 4227 1954 4373
rect 1946 4221 1947 4227
rect 1953 4221 1954 4227
rect 1946 4139 1954 4221
rect 1946 4133 1947 4139
rect 1953 4133 1954 4139
rect 1946 4003 1954 4133
rect 1946 3997 1947 4003
rect 1953 3997 1954 4003
rect 1946 3823 1954 3997
rect 1946 3817 1947 3823
rect 1953 3817 1954 3823
rect 1946 3767 1954 3817
rect 1946 3761 1947 3767
rect 1953 3761 1954 3767
rect 1946 3583 1954 3761
rect 1946 3577 1947 3583
rect 1953 3577 1954 3583
rect 1946 3507 1954 3577
rect 1946 3501 1947 3507
rect 1953 3501 1954 3507
rect 1946 3331 1954 3501
rect 1946 3325 1947 3331
rect 1953 3325 1954 3331
rect 1946 3267 1954 3325
rect 1946 3261 1947 3267
rect 1953 3261 1954 3267
rect 1946 3107 1954 3261
rect 1946 3101 1947 3107
rect 1953 3101 1954 3107
rect 1946 3027 1954 3101
rect 1946 3021 1947 3027
rect 1953 3021 1954 3027
rect 1946 2831 1954 3021
rect 1946 2825 1947 2831
rect 1953 2825 1954 2831
rect 1946 2787 1954 2825
rect 1946 2781 1947 2787
rect 1953 2781 1954 2787
rect 1946 2603 1954 2781
rect 1946 2597 1947 2603
rect 1953 2597 1954 2603
rect 1946 2547 1954 2597
rect 1946 2541 1947 2547
rect 1953 2541 1954 2547
rect 1946 2355 1954 2541
rect 1946 2349 1947 2355
rect 1953 2349 1954 2355
rect 1946 2307 1954 2349
rect 1946 2301 1947 2307
rect 1953 2301 1954 2307
rect 1946 2055 1954 2301
rect 1946 2049 1947 2055
rect 1953 2049 1954 2055
rect 1946 1941 1954 2049
rect 1946 1935 1947 1941
rect 1953 1935 1954 1941
rect 1946 1807 1954 1935
rect 1946 1801 1947 1807
rect 1953 1801 1954 1807
rect 1946 1693 1954 1801
rect 1946 1687 1947 1693
rect 1953 1687 1954 1693
rect 1946 1559 1954 1687
rect 1946 1553 1947 1559
rect 1953 1553 1954 1559
rect 1946 1445 1954 1553
rect 1946 1439 1947 1445
rect 1953 1439 1954 1445
rect 1946 1323 1954 1439
rect 1946 1317 1947 1323
rect 1953 1317 1954 1323
rect 1946 1211 1954 1317
rect 1946 1205 1947 1211
rect 1953 1205 1954 1211
rect 1946 1075 1954 1205
rect 1946 1069 1947 1075
rect 1953 1069 1954 1075
rect 1946 935 1954 1069
rect 1946 929 1947 935
rect 1953 929 1954 935
rect 1946 831 1954 929
rect 1946 825 1947 831
rect 1953 825 1954 831
rect 1946 607 1954 825
rect 1946 601 1947 607
rect 1953 601 1954 607
rect 1946 579 1954 601
rect 1946 573 1947 579
rect 1953 573 1954 579
rect 1946 367 1954 573
rect 1946 361 1947 367
rect 1953 361 1954 367
rect 1946 331 1954 361
rect 1946 325 1947 331
rect 1953 325 1954 331
rect 1946 111 1954 325
rect 1946 105 1947 111
rect 1953 105 1954 111
rect 1946 91 1954 105
rect 1946 85 1947 91
rect 1953 85 1954 91
rect 1946 72 1954 85
rect 1958 5759 1966 5760
rect 1958 5753 1959 5759
rect 1965 5753 1966 5759
rect 1958 5691 1966 5753
rect 1958 5685 1959 5691
rect 1965 5685 1966 5691
rect 1958 5535 1966 5685
rect 1958 5529 1959 5535
rect 1965 5529 1966 5535
rect 1958 5463 1966 5529
rect 1958 5457 1959 5463
rect 1965 5457 1966 5463
rect 1958 5311 1966 5457
rect 1958 5305 1959 5311
rect 1965 5305 1966 5311
rect 1958 5235 1966 5305
rect 1958 5229 1959 5235
rect 1965 5229 1966 5235
rect 1958 5079 1966 5229
rect 1958 5073 1959 5079
rect 1965 5073 1966 5079
rect 1958 4987 1966 5073
rect 1958 4981 1959 4987
rect 1965 4981 1966 4987
rect 1958 4815 1966 4981
rect 1958 4809 1959 4815
rect 1965 4809 1966 4815
rect 1958 4743 1966 4809
rect 1958 4737 1959 4743
rect 1965 4737 1966 4743
rect 1958 4575 1966 4737
rect 1958 4569 1959 4575
rect 1965 4569 1966 4575
rect 1958 4503 1966 4569
rect 1958 4497 1959 4503
rect 1965 4497 1966 4503
rect 1958 4347 1966 4497
rect 1958 4341 1959 4347
rect 1965 4341 1966 4347
rect 1958 4263 1966 4341
rect 1958 4257 1959 4263
rect 1965 4257 1966 4263
rect 1958 4115 1966 4257
rect 1958 4109 1959 4115
rect 1965 4109 1966 4115
rect 1958 3935 1966 4109
rect 1958 3929 1959 3935
rect 1965 3929 1966 3935
rect 1958 3891 1966 3929
rect 1958 3885 1959 3891
rect 1965 3885 1966 3891
rect 1958 3703 1966 3885
rect 1958 3697 1959 3703
rect 1965 3697 1966 3703
rect 1958 3639 1966 3697
rect 1958 3633 1959 3639
rect 1965 3633 1966 3639
rect 1958 3467 1966 3633
rect 1958 3461 1959 3467
rect 1965 3461 1966 3467
rect 1958 3387 1966 3461
rect 1958 3381 1959 3387
rect 1965 3381 1966 3387
rect 1958 3219 1966 3381
rect 1958 3213 1959 3219
rect 1965 3213 1966 3219
rect 1958 3139 1966 3213
rect 1958 3133 1959 3139
rect 1965 3133 1966 3139
rect 1958 2995 1966 3133
rect 1958 2989 1959 2995
rect 1965 2989 1966 2995
rect 1958 2911 1966 2989
rect 1958 2905 1959 2911
rect 1965 2905 1966 2911
rect 1958 2719 1966 2905
rect 1958 2713 1959 2719
rect 1965 2713 1966 2719
rect 1958 2675 1966 2713
rect 1958 2669 1959 2675
rect 1965 2669 1966 2675
rect 1958 2475 1966 2669
rect 1958 2469 1959 2475
rect 1965 2469 1966 2475
rect 1958 2423 1966 2469
rect 1958 2417 1959 2423
rect 1965 2417 1966 2423
rect 1958 2243 1966 2417
rect 1958 2237 1959 2243
rect 1965 2237 1966 2243
rect 1958 2171 1966 2237
rect 1958 2165 1959 2171
rect 1965 2165 1966 2171
rect 1958 1931 1966 2165
rect 1958 1925 1959 1931
rect 1965 1925 1966 1931
rect 1958 1807 1966 1925
rect 1958 1801 1959 1807
rect 1965 1801 1966 1807
rect 1958 1683 1966 1801
rect 1958 1677 1959 1683
rect 1965 1677 1966 1683
rect 1958 1559 1966 1677
rect 1958 1553 1959 1559
rect 1965 1553 1966 1559
rect 1958 1435 1966 1553
rect 1958 1429 1959 1435
rect 1965 1429 1966 1435
rect 1958 1323 1966 1429
rect 1958 1317 1959 1323
rect 1965 1317 1966 1323
rect 1958 1187 1966 1317
rect 1958 1181 1959 1187
rect 1965 1181 1966 1187
rect 1958 1075 1966 1181
rect 1958 1069 1959 1075
rect 1965 1069 1966 1075
rect 1958 959 1966 1069
rect 1958 953 1959 959
rect 1965 953 1966 959
rect 1958 823 1966 953
rect 1958 817 1959 823
rect 1965 817 1966 823
rect 1958 719 1966 817
rect 1958 713 1959 719
rect 1965 713 1966 719
rect 1958 495 1966 713
rect 1958 489 1959 495
rect 1965 489 1966 495
rect 1958 467 1966 489
rect 1958 461 1959 467
rect 1965 461 1966 467
rect 1958 223 1966 461
rect 1958 217 1959 223
rect 1965 217 1966 223
rect 1958 203 1966 217
rect 1958 197 1959 203
rect 1965 197 1966 203
rect 1958 72 1966 197
rect 3810 5579 3818 5760
rect 3810 5573 3811 5579
rect 3817 5573 3818 5579
rect 3810 5351 3818 5573
rect 3810 5345 3811 5351
rect 3817 5345 3818 5351
rect 3810 5107 3818 5345
rect 3810 5101 3811 5107
rect 3817 5101 3818 5107
rect 3810 4867 3818 5101
rect 3810 4861 3811 4867
rect 3817 4861 3818 4867
rect 3810 4803 3818 4861
rect 3810 4797 3811 4803
rect 3817 4797 3818 4803
rect 3810 4627 3818 4797
rect 3810 4621 3811 4627
rect 3817 4621 3818 4627
rect 3810 4579 3818 4621
rect 3810 4573 3811 4579
rect 3817 4573 3818 4579
rect 3810 4379 3818 4573
rect 3810 4373 3811 4379
rect 3817 4373 3818 4379
rect 3810 4335 3818 4373
rect 3810 4329 3811 4335
rect 3817 4329 3818 4335
rect 3810 4139 3818 4329
rect 3810 4133 3811 4139
rect 3817 4133 3818 4139
rect 3810 4075 3818 4133
rect 3810 4069 3811 4075
rect 3817 4069 3818 4075
rect 3810 3823 3818 4069
rect 3810 3817 3811 3823
rect 3817 3817 3818 3823
rect 3810 3583 3818 3817
rect 3810 3577 3811 3583
rect 3817 3577 3818 3583
rect 3810 3531 3818 3577
rect 3810 3525 3811 3531
rect 3817 3525 3818 3531
rect 3810 3331 3818 3525
rect 3810 3325 3811 3331
rect 3817 3325 3818 3331
rect 3810 3299 3818 3325
rect 3810 3293 3811 3299
rect 3817 3293 3818 3299
rect 3810 3107 3818 3293
rect 3810 3101 3811 3107
rect 3817 3101 3818 3107
rect 3810 3059 3818 3101
rect 3810 3053 3811 3059
rect 3817 3053 3818 3059
rect 3810 2831 3818 3053
rect 3810 2825 3811 2831
rect 3817 2825 3818 2831
rect 3810 2807 3818 2825
rect 3810 2801 3811 2807
rect 3817 2801 3818 2807
rect 3810 2603 3818 2801
rect 3810 2597 3811 2603
rect 3817 2597 3818 2603
rect 3810 2567 3818 2597
rect 3810 2561 3811 2567
rect 3817 2561 3818 2567
rect 3810 2355 3818 2561
rect 3810 2349 3811 2355
rect 3817 2349 3818 2355
rect 3810 2315 3818 2349
rect 3810 2309 3811 2315
rect 3817 2309 3818 2315
rect 3810 2067 3818 2309
rect 3810 2061 3811 2067
rect 3817 2061 3818 2067
rect 3810 1931 3818 2061
rect 3810 1925 3811 1931
rect 3817 1925 3818 1931
rect 3810 1843 3818 1925
rect 3810 1837 3811 1843
rect 3817 1837 3818 1843
rect 3810 1683 3818 1837
rect 3810 1677 3811 1683
rect 3817 1677 3818 1683
rect 3810 1587 3818 1677
rect 3810 1581 3811 1587
rect 3817 1581 3818 1587
rect 3810 1435 3818 1581
rect 3810 1429 3811 1435
rect 3817 1429 3818 1435
rect 3810 1287 3818 1429
rect 3810 1281 3811 1287
rect 3817 1281 3818 1287
rect 3810 1211 3818 1281
rect 3810 1205 3811 1211
rect 3817 1205 3818 1211
rect 3810 1055 3818 1205
rect 3810 1049 3811 1055
rect 3817 1049 3818 1055
rect 3810 935 3818 1049
rect 3810 929 3811 935
rect 3817 929 3818 935
rect 3810 833 3818 929
rect 3810 827 3811 833
rect 3817 827 3818 833
rect 3810 599 3818 827
rect 3810 593 3811 599
rect 3817 593 3818 599
rect 3810 579 3818 593
rect 3810 573 3811 579
rect 3817 573 3818 579
rect 3810 359 3818 573
rect 3810 353 3811 359
rect 3817 353 3818 359
rect 3810 331 3818 353
rect 3810 325 3811 331
rect 3817 325 3818 331
rect 3810 91 3818 325
rect 3810 85 3811 91
rect 3817 85 3818 91
rect 3810 72 3818 85
rect 3822 5691 3830 5760
rect 3822 5685 3823 5691
rect 3829 5685 3830 5691
rect 3822 5471 3830 5685
rect 3822 5465 3823 5471
rect 3829 5465 3830 5471
rect 3822 5463 3830 5465
rect 3822 5457 3823 5463
rect 3829 5457 3830 5463
rect 3822 5235 3830 5457
rect 3822 5229 3823 5235
rect 3829 5229 3830 5235
rect 3822 5223 3830 5229
rect 3822 5217 3823 5223
rect 3829 5217 3830 5223
rect 3822 4987 3830 5217
rect 3822 4981 3823 4987
rect 3829 4981 3830 4987
rect 3822 4743 3830 4981
rect 3822 4737 3823 4743
rect 3829 4737 3830 4743
rect 3822 4691 3830 4737
rect 3822 4685 3823 4691
rect 3829 4685 3830 4691
rect 3822 4503 3830 4685
rect 3822 4497 3823 4503
rect 3829 4497 3830 4503
rect 3822 4463 3830 4497
rect 3822 4457 3823 4463
rect 3829 4457 3830 4463
rect 3822 4263 3830 4457
rect 3822 4257 3823 4263
rect 3829 4257 3830 4263
rect 3822 4211 3830 4257
rect 3822 4205 3823 4211
rect 3829 4205 3830 4211
rect 3822 3963 3830 4205
rect 3822 3957 3823 3963
rect 3829 3957 3830 3963
rect 3822 3935 3830 3957
rect 3822 3929 3823 3935
rect 3829 3929 3830 3935
rect 3822 3703 3830 3929
rect 3822 3697 3823 3703
rect 3829 3697 3830 3703
rect 3822 3691 3830 3697
rect 3822 3685 3823 3691
rect 3829 3685 3830 3691
rect 3822 3467 3830 3685
rect 3822 3461 3823 3467
rect 3829 3461 3830 3467
rect 3822 3411 3830 3461
rect 3822 3405 3823 3411
rect 3829 3405 3830 3411
rect 3822 3219 3830 3405
rect 3822 3213 3823 3219
rect 3829 3213 3830 3219
rect 3822 3171 3830 3213
rect 3822 3165 3823 3171
rect 3829 3165 3830 3171
rect 3822 2995 3830 3165
rect 3822 2989 3823 2995
rect 3829 2989 3830 2995
rect 3822 2923 3830 2989
rect 3822 2917 3823 2923
rect 3829 2917 3830 2923
rect 3822 2719 3830 2917
rect 3822 2713 3823 2719
rect 3829 2713 3830 2719
rect 3822 2683 3830 2713
rect 3822 2677 3823 2683
rect 3829 2677 3830 2683
rect 3822 2475 3830 2677
rect 3822 2469 3823 2475
rect 3829 2469 3830 2475
rect 3822 2439 3830 2469
rect 3822 2433 3823 2439
rect 3829 2433 3830 2439
rect 3822 2243 3830 2433
rect 3822 2237 3823 2243
rect 3829 2237 3830 2243
rect 3822 2199 3830 2237
rect 3822 2193 3823 2199
rect 3829 2193 3830 2199
rect 3822 1955 3830 2193
rect 3822 1949 3823 1955
rect 3829 1949 3830 1955
rect 3822 1807 3830 1949
rect 3822 1801 3823 1807
rect 3829 1801 3830 1807
rect 3822 1715 3830 1801
rect 3822 1709 3823 1715
rect 3829 1709 3830 1715
rect 3822 1559 3830 1709
rect 3822 1553 3823 1559
rect 3829 1553 3830 1559
rect 3822 1403 3830 1553
rect 3822 1397 3823 1403
rect 3829 1397 3830 1403
rect 3822 1323 3830 1397
rect 3822 1317 3823 1323
rect 3829 1317 3830 1323
rect 3822 1167 3830 1317
rect 3822 1161 3823 1167
rect 3829 1161 3830 1167
rect 3822 1075 3830 1161
rect 3822 1069 3823 1075
rect 3829 1069 3830 1075
rect 3822 943 3830 1069
rect 3822 937 3823 943
rect 3829 937 3830 943
rect 3822 823 3830 937
rect 3822 817 3823 823
rect 3829 817 3830 823
rect 3822 711 3830 817
rect 3822 705 3823 711
rect 3829 705 3830 711
rect 3822 475 3830 705
rect 3822 469 3823 475
rect 3829 469 3830 475
rect 3822 467 3830 469
rect 3822 461 3823 467
rect 3829 461 3830 467
rect 3822 203 3830 461
rect 3822 197 3823 203
rect 3829 197 3830 203
rect 3822 72 3830 197
rect 5694 4803 5702 5760
rect 5694 4797 5695 4803
rect 5701 4797 5702 4803
rect 5694 4579 5702 4797
rect 5694 4573 5695 4579
rect 5701 4573 5702 4579
rect 5694 4335 5702 4573
rect 5694 4329 5695 4335
rect 5701 4329 5702 4335
rect 5694 4075 5702 4329
rect 5694 4069 5695 4075
rect 5701 4069 5702 4075
rect 5694 3531 5702 4069
rect 5694 3525 5695 3531
rect 5701 3525 5702 3531
rect 5694 3299 5702 3525
rect 5694 3293 5695 3299
rect 5701 3293 5702 3299
rect 5694 3059 5702 3293
rect 5694 3053 5695 3059
rect 5701 3053 5702 3059
rect 5694 2807 5702 3053
rect 5694 2801 5695 2807
rect 5701 2801 5702 2807
rect 5694 2567 5702 2801
rect 5694 2561 5695 2567
rect 5701 2561 5702 2567
rect 5694 2315 5702 2561
rect 5694 2309 5695 2315
rect 5701 2309 5702 2315
rect 5694 2067 5702 2309
rect 5694 2061 5695 2067
rect 5701 2061 5702 2067
rect 5694 1843 5702 2061
rect 5694 1837 5695 1843
rect 5701 1837 5702 1843
rect 5694 1587 5702 1837
rect 5694 1581 5695 1587
rect 5701 1581 5702 1587
rect 5694 1287 5702 1581
rect 5694 1281 5695 1287
rect 5701 1281 5702 1287
rect 5694 1055 5702 1281
rect 5694 1049 5695 1055
rect 5701 1049 5702 1055
rect 5694 831 5702 1049
rect 5694 825 5695 831
rect 5701 825 5702 831
rect 5694 599 5702 825
rect 5694 593 5695 599
rect 5701 593 5702 599
rect 5694 359 5702 593
rect 5694 353 5695 359
rect 5701 353 5702 359
rect 5694 72 5702 353
rect 5706 5471 5714 5760
rect 5706 5465 5707 5471
rect 5713 5465 5714 5471
rect 5706 5223 5714 5465
rect 5706 5217 5707 5223
rect 5713 5217 5714 5223
rect 5706 4691 5714 5217
rect 5706 4685 5707 4691
rect 5713 4685 5714 4691
rect 5706 4463 5714 4685
rect 5706 4457 5707 4463
rect 5713 4457 5714 4463
rect 5706 4211 5714 4457
rect 5706 4205 5707 4211
rect 5713 4205 5714 4211
rect 5706 3963 5714 4205
rect 5706 3957 5707 3963
rect 5713 3957 5714 3963
rect 5706 3691 5714 3957
rect 5706 3685 5707 3691
rect 5713 3685 5714 3691
rect 5706 3411 5714 3685
rect 5706 3405 5707 3411
rect 5713 3405 5714 3411
rect 5706 3171 5714 3405
rect 5706 3165 5707 3171
rect 5713 3165 5714 3171
rect 5706 2923 5714 3165
rect 5706 2917 5707 2923
rect 5713 2917 5714 2923
rect 5706 2683 5714 2917
rect 5706 2677 5707 2683
rect 5713 2677 5714 2683
rect 5706 2439 5714 2677
rect 5706 2433 5707 2439
rect 5713 2433 5714 2439
rect 5706 2199 5714 2433
rect 5706 2193 5707 2199
rect 5713 2193 5714 2199
rect 5706 1955 5714 2193
rect 5706 1949 5707 1955
rect 5713 1949 5714 1955
rect 5706 1715 5714 1949
rect 5706 1709 5707 1715
rect 5713 1709 5714 1715
rect 5706 1403 5714 1709
rect 5706 1397 5707 1403
rect 5713 1397 5714 1403
rect 5706 1167 5714 1397
rect 5706 1161 5707 1167
rect 5713 1161 5714 1167
rect 5706 943 5714 1161
rect 5706 937 5707 943
rect 5713 937 5714 943
rect 5706 711 5714 937
rect 5706 705 5707 711
rect 5713 705 5714 711
rect 5706 475 5714 705
rect 5706 469 5707 475
rect 5713 469 5714 475
rect 5706 72 5714 469
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__269
timestamp 1731220477
transform 1 0 5656 0 1 5604
box 7 3 12 24
use welltap_svt  __well_tap__268
timestamp 1731220477
transform 1 0 3832 0 1 5604
box 7 3 12 24
use welltap_svt  __well_tap__267
timestamp 1731220477
transform 1 0 5656 0 -1 5556
box 7 3 12 24
use welltap_svt  __well_tap__266
timestamp 1731220477
transform 1 0 3832 0 -1 5556
box 7 3 12 24
use welltap_svt  __well_tap__265
timestamp 1731220477
transform 1 0 5656 0 1 5380
box 7 3 12 24
use welltap_svt  __well_tap__264
timestamp 1731220477
transform 1 0 3832 0 1 5380
box 7 3 12 24
use welltap_svt  __well_tap__263
timestamp 1731220477
transform 1 0 5656 0 -1 5324
box 7 3 12 24
use welltap_svt  __well_tap__262
timestamp 1731220477
transform 1 0 3832 0 -1 5324
box 7 3 12 24
use welltap_svt  __well_tap__261
timestamp 1731220477
transform 1 0 5656 0 1 5132
box 7 3 12 24
use welltap_svt  __well_tap__260
timestamp 1731220477
transform 1 0 3832 0 1 5132
box 7 3 12 24
use welltap_svt  __well_tap__259
timestamp 1731220477
transform 1 0 5656 0 -1 5076
box 7 3 12 24
use welltap_svt  __well_tap__258
timestamp 1731220477
transform 1 0 3832 0 -1 5076
box 7 3 12 24
use welltap_svt  __well_tap__257
timestamp 1731220477
transform 1 0 5656 0 1 4900
box 7 3 12 24
use welltap_svt  __well_tap__256
timestamp 1731220477
transform 1 0 3832 0 1 4900
box 7 3 12 24
use welltap_svt  __well_tap__255
timestamp 1731220477
transform 1 0 5656 0 -1 4776
box 7 3 12 24
use welltap_svt  __well_tap__254
timestamp 1731220477
transform 1 0 3832 0 -1 4776
box 7 3 12 24
use welltap_svt  __well_tap__253
timestamp 1731220477
transform 1 0 5656 0 1 4600
box 7 3 12 24
use welltap_svt  __well_tap__252
timestamp 1731220477
transform 1 0 3832 0 1 4600
box 7 3 12 24
use welltap_svt  __well_tap__251
timestamp 1731220477
transform 1 0 5656 0 -1 4552
box 7 3 12 24
use welltap_svt  __well_tap__250
timestamp 1731220477
transform 1 0 3832 0 -1 4552
box 7 3 12 24
use welltap_svt  __well_tap__249
timestamp 1731220477
transform 1 0 5656 0 1 4372
box 7 3 12 24
use welltap_svt  __well_tap__248
timestamp 1731220477
transform 1 0 3832 0 1 4372
box 7 3 12 24
use welltap_svt  __well_tap__247
timestamp 1731220477
transform 1 0 5656 0 -1 4308
box 7 3 12 24
use welltap_svt  __well_tap__246
timestamp 1731220477
transform 1 0 3832 0 -1 4308
box 7 3 12 24
use welltap_svt  __well_tap__245
timestamp 1731220477
transform 1 0 5656 0 1 4120
box 7 3 12 24
use welltap_svt  __well_tap__244
timestamp 1731220477
transform 1 0 3832 0 1 4120
box 7 3 12 24
use welltap_svt  __well_tap__243
timestamp 1731220477
transform 1 0 5656 0 -1 4048
box 7 3 12 24
use welltap_svt  __well_tap__242
timestamp 1731220477
transform 1 0 3832 0 -1 4048
box 7 3 12 24
use welltap_svt  __well_tap__241
timestamp 1731220477
transform 1 0 5656 0 1 3872
box 7 3 12 24
use welltap_svt  __well_tap__240
timestamp 1731220477
transform 1 0 3832 0 1 3872
box 7 3 12 24
use welltap_svt  __well_tap__239
timestamp 1731220477
transform 1 0 5656 0 -1 3796
box 7 3 12 24
use welltap_svt  __well_tap__238
timestamp 1731220477
transform 1 0 3832 0 -1 3796
box 7 3 12 24
use welltap_svt  __well_tap__237
timestamp 1731220477
transform 1 0 5656 0 1 3600
box 7 3 12 24
use welltap_svt  __well_tap__236
timestamp 1731220477
transform 1 0 3832 0 1 3600
box 7 3 12 24
use welltap_svt  __well_tap__235
timestamp 1731220477
transform 1 0 5656 0 -1 3504
box 7 3 12 24
use welltap_svt  __well_tap__234
timestamp 1731220477
transform 1 0 3832 0 -1 3504
box 7 3 12 24
use welltap_svt  __well_tap__233
timestamp 1731220477
transform 1 0 5656 0 1 3320
box 7 3 12 24
use welltap_svt  __well_tap__232
timestamp 1731220477
transform 1 0 3832 0 1 3320
box 7 3 12 24
use welltap_svt  __well_tap__231
timestamp 1731220477
transform 1 0 5656 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__230
timestamp 1731220477
transform 1 0 3832 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__229
timestamp 1731220477
transform 1 0 5656 0 1 3080
box 7 3 12 24
use welltap_svt  __well_tap__228
timestamp 1731220477
transform 1 0 3832 0 1 3080
box 7 3 12 24
use welltap_svt  __well_tap__227
timestamp 1731220477
transform 1 0 5656 0 -1 3032
box 7 3 12 24
use welltap_svt  __well_tap__226
timestamp 1731220477
transform 1 0 3832 0 -1 3032
box 7 3 12 24
use welltap_svt  __well_tap__225
timestamp 1731220477
transform 1 0 5656 0 1 2832
box 7 3 12 24
use welltap_svt  __well_tap__224
timestamp 1731220477
transform 1 0 3832 0 1 2832
box 7 3 12 24
use welltap_svt  __well_tap__223
timestamp 1731220477
transform 1 0 5656 0 -1 2780
box 7 3 12 24
use welltap_svt  __well_tap__222
timestamp 1731220477
transform 1 0 3832 0 -1 2780
box 7 3 12 24
use welltap_svt  __well_tap__221
timestamp 1731220477
transform 1 0 5656 0 1 2592
box 7 3 12 24
use welltap_svt  __well_tap__220
timestamp 1731220477
transform 1 0 3832 0 1 2592
box 7 3 12 24
use welltap_svt  __well_tap__219
timestamp 1731220477
transform 1 0 5656 0 -1 2540
box 7 3 12 24
use welltap_svt  __well_tap__218
timestamp 1731220477
transform 1 0 3832 0 -1 2540
box 7 3 12 24
use welltap_svt  __well_tap__217
timestamp 1731220477
transform 1 0 5656 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__216
timestamp 1731220477
transform 1 0 3832 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__215
timestamp 1731220477
transform 1 0 5656 0 -1 2288
box 7 3 12 24
use welltap_svt  __well_tap__214
timestamp 1731220477
transform 1 0 3832 0 -1 2288
box 7 3 12 24
use welltap_svt  __well_tap__213
timestamp 1731220477
transform 1 0 5656 0 1 2108
box 7 3 12 24
use welltap_svt  __well_tap__212
timestamp 1731220477
transform 1 0 3832 0 1 2108
box 7 3 12 24
use welltap_svt  __well_tap__211
timestamp 1731220477
transform 1 0 5656 0 -1 2040
box 7 3 12 24
use welltap_svt  __well_tap__210
timestamp 1731220477
transform 1 0 3832 0 -1 2040
box 7 3 12 24
use welltap_svt  __well_tap__209
timestamp 1731220477
transform 1 0 5656 0 1 1864
box 7 3 12 24
use welltap_svt  __well_tap__208
timestamp 1731220477
transform 1 0 3832 0 1 1864
box 7 3 12 24
use welltap_svt  __well_tap__207
timestamp 1731220477
transform 1 0 5656 0 -1 1816
box 7 3 12 24
use welltap_svt  __well_tap__206
timestamp 1731220477
transform 1 0 3832 0 -1 1816
box 7 3 12 24
use welltap_svt  __well_tap__205
timestamp 1731220477
transform 1 0 5656 0 1 1624
box 7 3 12 24
use welltap_svt  __well_tap__204
timestamp 1731220477
transform 1 0 3832 0 1 1624
box 7 3 12 24
use welltap_svt  __well_tap__203
timestamp 1731220477
transform 1 0 5656 0 -1 1560
box 7 3 12 24
use welltap_svt  __well_tap__202
timestamp 1731220477
transform 1 0 3832 0 -1 1560
box 7 3 12 24
use welltap_svt  __well_tap__201
timestamp 1731220477
transform 1 0 5656 0 1 1312
box 7 3 12 24
use welltap_svt  __well_tap__200
timestamp 1731220477
transform 1 0 3832 0 1 1312
box 7 3 12 24
use welltap_svt  __well_tap__199
timestamp 1731220477
transform 1 0 5656 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__198
timestamp 1731220477
transform 1 0 3832 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__197
timestamp 1731220477
transform 1 0 5656 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__196
timestamp 1731220477
transform 1 0 3832 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__195
timestamp 1731220477
transform 1 0 5656 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220477
transform 1 0 3832 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220477
transform 1 0 5656 0 1 852
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220477
transform 1 0 3832 0 1 852
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220477
transform 1 0 5656 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220477
transform 1 0 3832 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220477
transform 1 0 5656 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220477
transform 1 0 3832 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220477
transform 1 0 5656 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220477
transform 1 0 3832 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220477
transform 1 0 5656 0 1 384
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220477
transform 1 0 3832 0 1 384
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220477
transform 1 0 5656 0 -1 332
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220477
transform 1 0 3832 0 -1 332
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220477
transform 1 0 5656 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220477
transform 1 0 3832 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220477
transform 1 0 3792 0 1 5600
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220477
transform 1 0 1968 0 1 5600
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220477
transform 1 0 3792 0 -1 5552
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220477
transform 1 0 1968 0 -1 5552
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220477
transform 1 0 3792 0 1 5372
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220477
transform 1 0 1968 0 1 5372
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220477
transform 1 0 3792 0 -1 5324
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220477
transform 1 0 1968 0 -1 5324
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220477
transform 1 0 3792 0 1 5144
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220477
transform 1 0 1968 0 1 5144
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220477
transform 1 0 3792 0 -1 5080
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220477
transform 1 0 1968 0 -1 5080
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220477
transform 1 0 3792 0 1 4896
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220477
transform 1 0 1968 0 1 4896
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220477
transform 1 0 3792 0 -1 4840
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220477
transform 1 0 1968 0 -1 4840
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220477
transform 1 0 3792 0 1 4652
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220477
transform 1 0 1968 0 1 4652
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220477
transform 1 0 3792 0 -1 4600
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220477
transform 1 0 1968 0 -1 4600
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220477
transform 1 0 3792 0 1 4412
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220477
transform 1 0 1968 0 1 4412
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220477
transform 1 0 3792 0 -1 4352
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220477
transform 1 0 1968 0 -1 4352
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220477
transform 1 0 3792 0 1 4172
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220477
transform 1 0 1968 0 1 4172
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220477
transform 1 0 3792 0 -1 4112
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220477
transform 1 0 1968 0 -1 4112
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220477
transform 1 0 3792 0 1 3844
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220477
transform 1 0 1968 0 1 3844
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220477
transform 1 0 3792 0 -1 3796
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220477
transform 1 0 1968 0 -1 3796
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220477
transform 1 0 3792 0 1 3612
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220477
transform 1 0 1968 0 1 3612
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220477
transform 1 0 3792 0 -1 3556
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220477
transform 1 0 1968 0 -1 3556
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220477
transform 1 0 3792 0 1 3376
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220477
transform 1 0 1968 0 1 3376
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220477
transform 1 0 3792 0 -1 3304
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220477
transform 1 0 1968 0 -1 3304
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220477
transform 1 0 3792 0 1 3128
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220477
transform 1 0 1968 0 1 3128
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220477
transform 1 0 3792 0 -1 3080
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220477
transform 1 0 1968 0 -1 3080
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220477
transform 1 0 3792 0 1 2904
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220477
transform 1 0 1968 0 1 2904
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220477
transform 1 0 3792 0 -1 2804
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220477
transform 1 0 1968 0 -1 2804
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220477
transform 1 0 3792 0 1 2628
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220477
transform 1 0 1968 0 1 2628
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220477
transform 1 0 3792 0 -1 2576
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220477
transform 1 0 1968 0 -1 2576
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220477
transform 1 0 3792 0 1 2384
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220477
transform 1 0 1968 0 1 2384
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220477
transform 1 0 3792 0 -1 2328
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220477
transform 1 0 1968 0 -1 2328
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220477
transform 1 0 3792 0 1 2152
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220477
transform 1 0 1968 0 1 2152
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220477
transform 1 0 3792 0 -1 1904
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220477
transform 1 0 1968 0 -1 1904
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220477
transform 1 0 3792 0 1 1716
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220477
transform 1 0 1968 0 1 1716
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220477
transform 1 0 3792 0 -1 1656
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220477
transform 1 0 1968 0 -1 1656
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220477
transform 1 0 3792 0 1 1468
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220477
transform 1 0 1968 0 1 1468
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220477
transform 1 0 3792 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220477
transform 1 0 1968 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220477
transform 1 0 3792 0 1 1232
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220477
transform 1 0 1968 0 1 1232
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220477
transform 1 0 3792 0 -1 1184
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220477
transform 1 0 1968 0 -1 1184
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220477
transform 1 0 3792 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220477
transform 1 0 1968 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220477
transform 1 0 3792 0 -1 908
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220477
transform 1 0 1968 0 -1 908
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220477
transform 1 0 3792 0 1 732
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220477
transform 1 0 1968 0 1 732
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220477
transform 1 0 3792 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220477
transform 1 0 1968 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220477
transform 1 0 3792 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220477
transform 1 0 1968 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220477
transform 1 0 3792 0 -1 304
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220477
transform 1 0 1968 0 -1 304
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220477
transform 1 0 3792 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220477
transform 1 0 1968 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220477
transform 1 0 1928 0 1 5668
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220477
transform 1 0 104 0 1 5668
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220477
transform 1 0 1928 0 -1 5620
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220477
transform 1 0 104 0 -1 5620
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220477
transform 1 0 1928 0 1 5444
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220477
transform 1 0 104 0 1 5444
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220477
transform 1 0 1928 0 -1 5396
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220477
transform 1 0 104 0 -1 5396
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220477
transform 1 0 1928 0 1 5220
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220477
transform 1 0 104 0 1 5220
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220477
transform 1 0 1928 0 -1 5172
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220477
transform 1 0 104 0 -1 5172
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220477
transform 1 0 1928 0 1 4988
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220477
transform 1 0 104 0 1 4988
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220477
transform 1 0 1928 0 -1 4912
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220477
transform 1 0 104 0 -1 4912
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220477
transform 1 0 1928 0 1 4724
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220477
transform 1 0 104 0 1 4724
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220477
transform 1 0 1928 0 -1 4672
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220477
transform 1 0 104 0 -1 4672
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220477
transform 1 0 1928 0 1 4484
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220477
transform 1 0 104 0 1 4484
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220477
transform 1 0 1928 0 -1 4436
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220477
transform 1 0 104 0 -1 4436
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220477
transform 1 0 1928 0 1 4256
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220477
transform 1 0 104 0 1 4256
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220477
transform 1 0 1928 0 -1 4200
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220477
transform 1 0 104 0 -1 4200
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220477
transform 1 0 1928 0 1 4024
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220477
transform 1 0 104 0 1 4024
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220477
transform 1 0 1928 0 -1 3976
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220477
transform 1 0 104 0 -1 3976
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220477
transform 1 0 1928 0 1 3800
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220477
transform 1 0 104 0 1 3800
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220477
transform 1 0 1928 0 -1 3740
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220477
transform 1 0 104 0 -1 3740
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220477
transform 1 0 1928 0 1 3548
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220477
transform 1 0 104 0 1 3548
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220477
transform 1 0 1928 0 -1 3480
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220477
transform 1 0 104 0 -1 3480
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220477
transform 1 0 1928 0 1 3296
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220477
transform 1 0 104 0 1 3296
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220477
transform 1 0 1928 0 -1 3240
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220477
transform 1 0 104 0 -1 3240
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220477
transform 1 0 1928 0 1 3048
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220477
transform 1 0 104 0 1 3048
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220477
transform 1 0 1928 0 -1 3000
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220477
transform 1 0 104 0 -1 3000
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220477
transform 1 0 1928 0 1 2820
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220477
transform 1 0 104 0 1 2820
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220477
transform 1 0 1928 0 -1 2760
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220477
transform 1 0 104 0 -1 2760
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220477
transform 1 0 1928 0 1 2584
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220477
transform 1 0 104 0 1 2584
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220477
transform 1 0 1928 0 -1 2520
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220477
transform 1 0 104 0 -1 2520
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220477
transform 1 0 1928 0 1 2332
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220477
transform 1 0 104 0 1 2332
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220477
transform 1 0 1928 0 -1 2280
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220477
transform 1 0 104 0 -1 2280
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220477
transform 1 0 1928 0 1 2080
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220477
transform 1 0 104 0 1 2080
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220477
transform 1 0 1928 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220477
transform 1 0 104 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220477
transform 1 0 1928 0 1 1840
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220477
transform 1 0 104 0 1 1840
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220477
transform 1 0 1928 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220477
transform 1 0 104 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220477
transform 1 0 1928 0 1 1592
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220477
transform 1 0 104 0 1 1592
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220477
transform 1 0 1928 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220477
transform 1 0 104 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220477
transform 1 0 1928 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220477
transform 1 0 104 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220477
transform 1 0 1928 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220477
transform 1 0 104 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220477
transform 1 0 1928 0 1 1096
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220477
transform 1 0 104 0 1 1096
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220477
transform 1 0 1928 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220477
transform 1 0 104 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220477
transform 1 0 1928 0 1 868
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220477
transform 1 0 104 0 1 868
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220477
transform 1 0 1928 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220477
transform 1 0 104 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220477
transform 1 0 1928 0 1 628
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220477
transform 1 0 104 0 1 628
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220477
transform 1 0 1928 0 -1 580
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220477
transform 1 0 104 0 -1 580
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220477
transform 1 0 1928 0 1 404
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220477
transform 1 0 104 0 1 404
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220477
transform 1 0 1928 0 -1 340
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220477
transform 1 0 104 0 -1 340
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220477
transform 1 0 1928 0 1 132
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220477
transform 1 0 104 0 1 132
box 7 3 12 24
use _0_0std_0_0cells_0_0FAX1  tst_5999_6
timestamp 1731220477
transform 1 0 5376 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5998_6
timestamp 1731220477
transform 1 0 5512 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5997_6
timestamp 1731220477
transform 1 0 5512 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5996_6
timestamp 1731220477
transform 1 0 5504 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5995_6
timestamp 1731220477
transform 1 0 5456 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5994_6
timestamp 1731220477
transform 1 0 5416 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5993_6
timestamp 1731220477
transform 1 0 5280 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5992_6
timestamp 1731220477
transform 1 0 5200 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5991_6
timestamp 1731220477
transform 1 0 5040 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5990_6
timestamp 1731220477
transform 1 0 5368 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5989_6
timestamp 1731220477
transform 1 0 5240 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5988_6
timestamp 1731220477
transform 1 0 5104 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5987_6
timestamp 1731220477
transform 1 0 4968 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5986_6
timestamp 1731220477
transform 1 0 4832 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5985_6
timestamp 1731220477
transform 1 0 4696 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5984_6
timestamp 1731220477
transform 1 0 4560 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5983_6
timestamp 1731220477
transform 1 0 4424 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5982_6
timestamp 1731220477
transform 1 0 4288 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5981_6
timestamp 1731220477
transform 1 0 4720 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5980_6
timestamp 1731220477
transform 1 0 4880 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5979_6
timestamp 1731220477
transform 1 0 5064 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5978_6
timestamp 1731220477
transform 1 0 4856 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5977_6
timestamp 1731220477
transform 1 0 4648 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5976_6
timestamp 1731220477
transform 1 0 4448 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5975_6
timestamp 1731220477
transform 1 0 5160 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5974_6
timestamp 1731220477
transform 1 0 4904 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5973_6
timestamp 1731220477
transform 1 0 4664 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5972_6
timestamp 1731220477
transform 1 0 4448 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5971_6
timestamp 1731220477
transform 1 0 4264 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5970_6
timestamp 1731220477
transform 1 0 5224 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5969_6
timestamp 1731220477
transform 1 0 4992 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5968_6
timestamp 1731220477
transform 1 0 4768 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5967_6
timestamp 1731220477
transform 1 0 4568 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5966_6
timestamp 1731220477
transform 1 0 4248 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5965_6
timestamp 1731220477
transform 1 0 3968 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5964_6
timestamp 1731220477
transform 1 0 3856 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5963_6
timestamp 1731220477
transform 1 0 4040 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5962_6
timestamp 1731220477
transform 1 0 4064 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5961_6
timestamp 1731220477
transform 1 0 3856 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5960_6
timestamp 1731220477
transform 1 0 3648 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5959_6
timestamp 1731220477
transform 1 0 3648 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5958_6
timestamp 1731220477
transform 1 0 3464 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5957_6
timestamp 1731220477
transform 1 0 3424 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5956_6
timestamp 1731220477
transform 1 0 3176 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5955_6
timestamp 1731220477
transform 1 0 3392 0 1 960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5954_6
timestamp 1731220477
transform 1 0 3240 0 1 960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5953_6
timestamp 1731220477
transform 1 0 3176 0 -1 932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5952_6
timestamp 1731220477
transform 1 0 3464 0 -1 932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5951_6
timestamp 1731220477
transform 1 0 3448 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5950_6
timestamp 1731220477
transform 1 0 3224 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5949_6
timestamp 1731220477
transform 1 0 3648 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5948_6
timestamp 1731220477
transform 1 0 3856 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5947_6
timestamp 1731220477
transform 1 0 3856 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5946_6
timestamp 1731220477
transform 1 0 3992 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5945_6
timestamp 1731220477
transform 1 0 4128 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5944_6
timestamp 1731220477
transform 1 0 4400 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5943_6
timestamp 1731220477
transform 1 0 4264 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5942_6
timestamp 1731220477
transform 1 0 4128 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5941_6
timestamp 1731220477
transform 1 0 3992 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5940_6
timestamp 1731220477
transform 1 0 3856 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5939_6
timestamp 1731220477
transform 1 0 4016 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5938_6
timestamp 1731220477
transform 1 0 5192 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5937_6
timestamp 1731220477
transform 1 0 4848 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5936_6
timestamp 1731220477
transform 1 0 4528 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5935_6
timestamp 1731220477
transform 1 0 4400 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5934_6
timestamp 1731220477
transform 1 0 4176 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5933_6
timestamp 1731220477
transform 1 0 4896 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5932_6
timestamp 1731220477
transform 1 0 4640 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5931_6
timestamp 1731220477
transform 1 0 4480 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5930_6
timestamp 1731220477
transform 1 0 4248 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5929_6
timestamp 1731220477
transform 1 0 4992 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5928_6
timestamp 1731220477
transform 1 0 4728 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5927_6
timestamp 1731220477
transform 1 0 4536 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5926_6
timestamp 1731220477
transform 1 0 4296 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5925_6
timestamp 1731220477
transform 1 0 5024 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5924_6
timestamp 1731220477
transform 1 0 4776 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5923_6
timestamp 1731220477
transform 1 0 4704 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5922_6
timestamp 1731220477
transform 1 0 5000 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5921_6
timestamp 1731220477
transform 1 0 4848 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5920_6
timestamp 1731220477
transform 1 0 4808 0 1 1288
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5919_6
timestamp 1731220477
transform 1 0 4944 0 1 1288
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5918_6
timestamp 1731220477
transform 1 0 5080 0 1 1288
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5917_6
timestamp 1731220477
transform 1 0 5216 0 1 1288
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5916_6
timestamp 1731220477
transform 1 0 5160 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5915_6
timestamp 1731220477
transform 1 0 5328 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5914_6
timestamp 1731220477
transform 1 0 5280 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5913_6
timestamp 1731220477
transform 1 0 5264 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5912_6
timestamp 1731220477
transform 1 0 5168 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5911_6
timestamp 1731220477
transform 1 0 5440 0 1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5910_6
timestamp 1731220477
transform 1 0 5512 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5909_6
timestamp 1731220477
transform 1 0 5512 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5908_6
timestamp 1731220477
transform 1 0 5512 0 1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5907_6
timestamp 1731220477
transform 1 0 5496 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5906_6
timestamp 1731220477
transform 1 0 5488 0 1 1288
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5905_6
timestamp 1731220477
transform 1 0 5352 0 1 1288
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5904_6
timestamp 1731220477
transform 1 0 5512 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5903_6
timestamp 1731220477
transform 1 0 5376 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5902_6
timestamp 1731220477
transform 1 0 5104 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5901_6
timestamp 1731220477
transform 1 0 4968 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5900_6
timestamp 1731220477
transform 1 0 5240 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5899_6
timestamp 1731220477
transform 1 0 5104 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5898_6
timestamp 1731220477
transform 1 0 4968 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5897_6
timestamp 1731220477
transform 1 0 4832 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5896_6
timestamp 1731220477
transform 1 0 4696 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5895_6
timestamp 1731220477
transform 1 0 4560 0 -1 1584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5894_6
timestamp 1731220477
transform 1 0 4560 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5893_6
timestamp 1731220477
transform 1 0 4696 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5892_6
timestamp 1731220477
transform 1 0 4832 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5891_6
timestamp 1731220477
transform 1 0 4920 0 -1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5890_6
timestamp 1731220477
transform 1 0 4784 0 -1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5889_6
timestamp 1731220477
transform 1 0 4648 0 -1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5888_6
timestamp 1731220477
transform 1 0 4512 0 -1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5887_6
timestamp 1731220477
transform 1 0 4376 0 -1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5886_6
timestamp 1731220477
transform 1 0 5200 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5885_6
timestamp 1731220477
transform 1 0 4872 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5884_6
timestamp 1731220477
transform 1 0 4560 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5883_6
timestamp 1731220477
transform 1 0 4280 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5882_6
timestamp 1731220477
transform 1 0 4040 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5881_6
timestamp 1731220477
transform 1 0 4536 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5880_6
timestamp 1731220477
transform 1 0 4688 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5879_6
timestamp 1731220477
transform 1 0 4864 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5878_6
timestamp 1731220477
transform 1 0 5056 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5877_6
timestamp 1731220477
transform 1 0 5248 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5876_6
timestamp 1731220477
transform 1 0 5312 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5875_6
timestamp 1731220477
transform 1 0 5096 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5874_6
timestamp 1731220477
transform 1 0 4888 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5873_6
timestamp 1731220477
transform 1 0 4696 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5872_6
timestamp 1731220477
transform 1 0 4536 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5871_6
timestamp 1731220477
transform 1 0 4464 0 -1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5870_6
timestamp 1731220477
transform 1 0 4152 0 -1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5869_6
timestamp 1731220477
transform 1 0 4760 0 -1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5868_6
timestamp 1731220477
transform 1 0 5056 0 -1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5867_6
timestamp 1731220477
transform 1 0 5352 0 -1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5866_6
timestamp 1731220477
transform 1 0 5240 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5865_6
timestamp 1731220477
transform 1 0 5104 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5864_6
timestamp 1731220477
transform 1 0 4968 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5863_6
timestamp 1731220477
transform 1 0 4832 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5862_6
timestamp 1731220477
transform 1 0 4696 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5861_6
timestamp 1731220477
transform 1 0 5008 0 -1 2564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5860_6
timestamp 1731220477
transform 1 0 4872 0 -1 2564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5859_6
timestamp 1731220477
transform 1 0 4736 0 -1 2564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5858_6
timestamp 1731220477
transform 1 0 4600 0 -1 2564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5857_6
timestamp 1731220477
transform 1 0 4464 0 -1 2564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5856_6
timestamp 1731220477
transform 1 0 5008 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5855_6
timestamp 1731220477
transform 1 0 4752 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5854_6
timestamp 1731220477
transform 1 0 4512 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5853_6
timestamp 1731220477
transform 1 0 4296 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5852_6
timestamp 1731220477
transform 1 0 4096 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5851_6
timestamp 1731220477
transform 1 0 4432 0 -1 2804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5850_6
timestamp 1731220477
transform 1 0 4296 0 -1 2804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5849_6
timestamp 1731220477
transform 1 0 4160 0 -1 2804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5848_6
timestamp 1731220477
transform 1 0 4024 0 -1 2804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5847_6
timestamp 1731220477
transform 1 0 3888 0 -1 2804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5846_6
timestamp 1731220477
transform 1 0 3992 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5845_6
timestamp 1731220477
transform 1 0 4208 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5844_6
timestamp 1731220477
transform 1 0 4968 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5843_6
timestamp 1731220477
transform 1 0 4696 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5842_6
timestamp 1731220477
transform 1 0 4440 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5841_6
timestamp 1731220477
transform 1 0 4424 0 -1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5840_6
timestamp 1731220477
transform 1 0 4224 0 -1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5839_6
timestamp 1731220477
transform 1 0 5136 0 -1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5838_6
timestamp 1731220477
transform 1 0 4880 0 -1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5837_6
timestamp 1731220477
transform 1 0 4640 0 -1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5836_6
timestamp 1731220477
transform 1 0 4464 0 1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5835_6
timestamp 1731220477
transform 1 0 4648 0 1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5834_6
timestamp 1731220477
transform 1 0 5304 0 1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5833_6
timestamp 1731220477
transform 1 0 5072 0 1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5832_6
timestamp 1731220477
transform 1 0 4856 0 1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5831_6
timestamp 1731220477
transform 1 0 4576 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5830_6
timestamp 1731220477
transform 1 0 4344 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5829_6
timestamp 1731220477
transform 1 0 4984 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5828_6
timestamp 1731220477
transform 1 0 4784 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5827_6
timestamp 1731220477
transform 1 0 4584 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5826_6
timestamp 1731220477
transform 1 0 4808 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5825_6
timestamp 1731220477
transform 1 0 5024 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5824_6
timestamp 1731220477
transform 1 0 5232 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5823_6
timestamp 1731220477
transform 1 0 5448 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5822_6
timestamp 1731220477
transform 1 0 5352 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5821_6
timestamp 1731220477
transform 1 0 5168 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5820_6
timestamp 1731220477
transform 1 0 5392 0 -1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5819_6
timestamp 1731220477
transform 1 0 5248 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5818_6
timestamp 1731220477
transform 1 0 5272 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5817_6
timestamp 1731220477
transform 1 0 5376 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5816_6
timestamp 1731220477
transform 1 0 5448 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5815_6
timestamp 1731220477
transform 1 0 5376 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5814_6
timestamp 1731220477
transform 1 0 5240 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5813_6
timestamp 1731220477
transform 1 0 5512 0 1 1600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5812_6
timestamp 1731220477
transform 1 0 5512 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5811_6
timestamp 1731220477
transform 1 0 5512 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5810_6
timestamp 1731220477
transform 1 0 5512 0 1 2324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5809_6
timestamp 1731220477
transform 1 0 5512 0 1 2568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5808_6
timestamp 1731220477
transform 1 0 5512 0 1 2808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5807_6
timestamp 1731220477
transform 1 0 5512 0 1 3056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5806_6
timestamp 1731220477
transform 1 0 5512 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5805_6
timestamp 1731220477
transform 1 0 5512 0 -1 3528
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5804_6
timestamp 1731220477
transform 1 0 5376 0 -1 3528
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5803_6
timestamp 1731220477
transform 1 0 5512 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5802_6
timestamp 1731220477
transform 1 0 5376 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5801_6
timestamp 1731220477
transform 1 0 5240 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5800_6
timestamp 1731220477
transform 1 0 5104 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5799_6
timestamp 1731220477
transform 1 0 4968 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5798_6
timestamp 1731220477
transform 1 0 4832 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5797_6
timestamp 1731220477
transform 1 0 4696 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5796_6
timestamp 1731220477
transform 1 0 4560 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5795_6
timestamp 1731220477
transform 1 0 4424 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5794_6
timestamp 1731220477
transform 1 0 4288 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5793_6
timestamp 1731220477
transform 1 0 4152 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5792_6
timestamp 1731220477
transform 1 0 4016 0 1 3576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5791_6
timestamp 1731220477
transform 1 0 5016 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5790_6
timestamp 1731220477
transform 1 0 4880 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5789_6
timestamp 1731220477
transform 1 0 4744 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5788_6
timestamp 1731220477
transform 1 0 4608 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5787_6
timestamp 1731220477
transform 1 0 4472 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5786_6
timestamp 1731220477
transform 1 0 4776 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5785_6
timestamp 1731220477
transform 1 0 4616 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5784_6
timestamp 1731220477
transform 1 0 4456 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5783_6
timestamp 1731220477
transform 1 0 4296 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5782_6
timestamp 1731220477
transform 1 0 4144 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5781_6
timestamp 1731220477
transform 1 0 4808 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5780_6
timestamp 1731220477
transform 1 0 4672 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5779_6
timestamp 1731220477
transform 1 0 4536 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5778_6
timestamp 1731220477
transform 1 0 4400 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5777_6
timestamp 1731220477
transform 1 0 4264 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5776_6
timestamp 1731220477
transform 1 0 4104 0 1 4096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5775_6
timestamp 1731220477
transform 1 0 3968 0 1 4096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5774_6
timestamp 1731220477
transform 1 0 4512 0 1 4096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5773_6
timestamp 1731220477
transform 1 0 4376 0 1 4096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5772_6
timestamp 1731220477
transform 1 0 4240 0 1 4096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5771_6
timestamp 1731220477
transform 1 0 4104 0 -1 4332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5770_6
timestamp 1731220477
transform 1 0 4240 0 -1 4332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5769_6
timestamp 1731220477
transform 1 0 4648 0 -1 4332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5768_6
timestamp 1731220477
transform 1 0 4512 0 -1 4332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5767_6
timestamp 1731220477
transform 1 0 4376 0 -1 4332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5766_6
timestamp 1731220477
transform 1 0 4344 0 1 4348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5765_6
timestamp 1731220477
transform 1 0 4480 0 1 4348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5764_6
timestamp 1731220477
transform 1 0 4616 0 1 4348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5763_6
timestamp 1731220477
transform 1 0 4752 0 1 4348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5762_6
timestamp 1731220477
transform 1 0 4888 0 1 4348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5761_6
timestamp 1731220477
transform 1 0 5048 0 -1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5760_6
timestamp 1731220477
transform 1 0 4912 0 -1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5759_6
timestamp 1731220477
transform 1 0 4776 0 -1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5758_6
timestamp 1731220477
transform 1 0 4640 0 -1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5757_6
timestamp 1731220477
transform 1 0 4400 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5756_6
timestamp 1731220477
transform 1 0 4264 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5755_6
timestamp 1731220477
transform 1 0 4128 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5754_6
timestamp 1731220477
transform 1 0 4536 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5753_6
timestamp 1731220477
transform 1 0 4672 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5752_6
timestamp 1731220477
transform 1 0 4816 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5751_6
timestamp 1731220477
transform 1 0 4960 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5750_6
timestamp 1731220477
transform 1 0 5104 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5749_6
timestamp 1731220477
transform 1 0 5240 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5748_6
timestamp 1731220477
transform 1 0 5512 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5747_6
timestamp 1731220477
transform 1 0 5376 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5746_6
timestamp 1731220477
transform 1 0 5272 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5745_6
timestamp 1731220477
transform 1 0 5008 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5744_6
timestamp 1731220477
transform 1 0 5512 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5743_6
timestamp 1731220477
transform 1 0 5512 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5742_6
timestamp 1731220477
transform 1 0 5376 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5741_6
timestamp 1731220477
transform 1 0 5280 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5740_6
timestamp 1731220477
transform 1 0 5032 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5739_6
timestamp 1731220477
transform 1 0 5512 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5738_6
timestamp 1731220477
transform 1 0 5512 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5737_6
timestamp 1731220477
transform 1 0 5376 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5736_6
timestamp 1731220477
transform 1 0 5216 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5735_6
timestamp 1731220477
transform 1 0 5064 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5734_6
timestamp 1731220477
transform 1 0 4912 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5733_6
timestamp 1731220477
transform 1 0 4752 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5732_6
timestamp 1731220477
transform 1 0 4592 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5731_6
timestamp 1731220477
transform 1 0 4768 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5730_6
timestamp 1731220477
transform 1 0 4952 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5729_6
timestamp 1731220477
transform 1 0 5144 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5728_6
timestamp 1731220477
transform 1 0 5072 0 1 5356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5727_6
timestamp 1731220477
transform 1 0 4904 0 1 5356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5726_6
timestamp 1731220477
transform 1 0 4744 0 1 5356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5725_6
timestamp 1731220477
transform 1 0 5080 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5724_6
timestamp 1731220477
transform 1 0 4944 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5723_6
timestamp 1731220477
transform 1 0 4808 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5722_6
timestamp 1731220477
transform 1 0 4672 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5721_6
timestamp 1731220477
transform 1 0 4872 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5720_6
timestamp 1731220477
transform 1 0 4736 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5719_6
timestamp 1731220477
transform 1 0 4600 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5718_6
timestamp 1731220477
transform 1 0 4464 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5717_6
timestamp 1731220477
transform 1 0 4400 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5716_6
timestamp 1731220477
transform 1 0 4536 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5715_6
timestamp 1731220477
transform 1 0 4584 0 1 5356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5714_6
timestamp 1731220477
transform 1 0 4424 0 1 5356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5713_6
timestamp 1731220477
transform 1 0 4400 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5712_6
timestamp 1731220477
transform 1 0 4584 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5711_6
timestamp 1731220477
transform 1 0 4432 0 1 5108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5710_6
timestamp 1731220477
transform 1 0 4296 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5709_6
timestamp 1731220477
transform 1 0 4536 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5708_6
timestamp 1731220477
transform 1 0 4784 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5707_6
timestamp 1731220477
transform 1 0 5224 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5706_6
timestamp 1731220477
transform 1 0 5080 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5705_6
timestamp 1731220477
transform 1 0 4944 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5704_6
timestamp 1731220477
transform 1 0 4808 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5703_6
timestamp 1731220477
transform 1 0 4672 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5702_6
timestamp 1731220477
transform 1 0 4536 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5701_6
timestamp 1731220477
transform 1 0 4400 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5700_6
timestamp 1731220477
transform 1 0 4264 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5699_6
timestamp 1731220477
transform 1 0 4128 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5698_6
timestamp 1731220477
transform 1 0 4056 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5697_6
timestamp 1731220477
transform 1 0 3856 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5696_6
timestamp 1731220477
transform 1 0 3992 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5695_6
timestamp 1731220477
transform 1 0 3856 0 1 4876
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5694_6
timestamp 1731220477
transform 1 0 3648 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5693_6
timestamp 1731220477
transform 1 0 3648 0 -1 4864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5692_6
timestamp 1731220477
transform 1 0 3856 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5691_6
timestamp 1731220477
transform 1 0 4040 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5690_6
timestamp 1731220477
transform 1 0 4752 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5689_6
timestamp 1731220477
transform 1 0 4504 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5688_6
timestamp 1731220477
transform 1 0 4264 0 -1 4800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5687_6
timestamp 1731220477
transform 1 0 3992 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5686_6
timestamp 1731220477
transform 1 0 3856 0 1 4576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5685_6
timestamp 1731220477
transform 1 0 3648 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5684_6
timestamp 1731220477
transform 1 0 3440 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5683_6
timestamp 1731220477
transform 1 0 3216 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5682_6
timestamp 1731220477
transform 1 0 2984 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5681_6
timestamp 1731220477
transform 1 0 3608 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5680_6
timestamp 1731220477
transform 1 0 3392 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5679_6
timestamp 1731220477
transform 1 0 3184 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5678_6
timestamp 1731220477
transform 1 0 2968 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5677_6
timestamp 1731220477
transform 1 0 2744 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5676_6
timestamp 1731220477
transform 1 0 3288 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5675_6
timestamp 1731220477
transform 1 0 3104 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5674_6
timestamp 1731220477
transform 1 0 2920 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5673_6
timestamp 1731220477
transform 1 0 2744 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5672_6
timestamp 1731220477
transform 1 0 2560 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5671_6
timestamp 1731220477
transform 1 0 2504 0 1 4148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5670_6
timestamp 1731220477
transform 1 0 2240 0 1 4148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5669_6
timestamp 1731220477
transform 1 0 2760 0 1 4148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5668_6
timestamp 1731220477
transform 1 0 3016 0 1 4148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5667_6
timestamp 1731220477
transform 1 0 3280 0 1 4148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5666_6
timestamp 1731220477
transform 1 0 3240 0 -1 4136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5665_6
timestamp 1731220477
transform 1 0 3104 0 -1 4136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5664_6
timestamp 1731220477
transform 1 0 3376 0 -1 4136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5663_6
timestamp 1731220477
transform 1 0 3512 0 -1 4136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5662_6
timestamp 1731220477
transform 1 0 3648 0 -1 4136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5661_6
timestamp 1731220477
transform 1 0 3856 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5660_6
timestamp 1731220477
transform 1 0 3992 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5659_6
timestamp 1731220477
transform 1 0 4128 0 -1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5658_6
timestamp 1731220477
transform 1 0 3992 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5657_6
timestamp 1731220477
transform 1 0 3856 0 1 3848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5656_6
timestamp 1731220477
transform 1 0 3648 0 1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5655_6
timestamp 1731220477
transform 1 0 3248 0 1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5654_6
timestamp 1731220477
transform 1 0 2824 0 1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5653_6
timestamp 1731220477
transform 1 0 2400 0 1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5652_6
timestamp 1731220477
transform 1 0 3576 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5651_6
timestamp 1731220477
transform 1 0 3392 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5650_6
timestamp 1731220477
transform 1 0 3216 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5649_6
timestamp 1731220477
transform 1 0 3040 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5648_6
timestamp 1731220477
transform 1 0 2864 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5647_6
timestamp 1731220477
transform 1 0 3296 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5646_6
timestamp 1731220477
transform 1 0 3152 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5645_6
timestamp 1731220477
transform 1 0 3008 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5644_6
timestamp 1731220477
transform 1 0 2864 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5643_6
timestamp 1731220477
transform 1 0 2720 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5642_6
timestamp 1731220477
transform 1 0 2888 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5641_6
timestamp 1731220477
transform 1 0 3024 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5640_6
timestamp 1731220477
transform 1 0 3160 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5639_6
timestamp 1731220477
transform 1 0 3432 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5638_6
timestamp 1731220477
transform 1 0 3296 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5637_6
timestamp 1731220477
transform 1 0 3288 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5636_6
timestamp 1731220477
transform 1 0 3096 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5635_6
timestamp 1731220477
transform 1 0 3480 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5634_6
timestamp 1731220477
transform 1 0 3648 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5633_6
timestamp 1731220477
transform 1 0 3856 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5632_6
timestamp 1731220477
transform 1 0 4096 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5631_6
timestamp 1731220477
transform 1 0 4344 0 1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5630_6
timestamp 1731220477
transform 1 0 4096 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5629_6
timestamp 1731220477
transform 1 0 3856 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5628_6
timestamp 1731220477
transform 1 0 3648 0 -1 3328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5627_6
timestamp 1731220477
transform 1 0 3648 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5626_6
timestamp 1731220477
transform 1 0 3440 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5625_6
timestamp 1731220477
transform 1 0 3208 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5624_6
timestamp 1731220477
transform 1 0 3368 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5623_6
timestamp 1731220477
transform 1 0 3536 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5622_6
timestamp 1731220477
transform 1 0 3480 0 1 2880
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5621_6
timestamp 1731220477
transform 1 0 3344 0 1 2880
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5620_6
timestamp 1731220477
transform 1 0 3208 0 1 2880
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5619_6
timestamp 1731220477
transform 1 0 3072 0 1 2880
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5618_6
timestamp 1731220477
transform 1 0 3208 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5617_6
timestamp 1731220477
transform 1 0 3048 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5616_6
timestamp 1731220477
transform 1 0 2896 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5615_6
timestamp 1731220477
transform 1 0 2768 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5614_6
timestamp 1731220477
transform 1 0 2552 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5613_6
timestamp 1731220477
transform 1 0 2656 0 -1 3328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5612_6
timestamp 1731220477
transform 1 0 2368 0 -1 3328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5611_6
timestamp 1731220477
transform 1 0 2120 0 -1 3328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5610_6
timestamp 1731220477
transform 1 0 2344 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5609_6
timestamp 1731220477
transform 1 0 2144 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5608_6
timestamp 1731220477
transform 1 0 1992 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5607_6
timestamp 1731220477
transform 1 0 1784 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5606_6
timestamp 1731220477
transform 1 0 1576 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5605_6
timestamp 1731220477
transform 1 0 1344 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5604_6
timestamp 1731220477
transform 1 0 1784 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5603_6
timestamp 1731220477
transform 1 0 1640 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5602_6
timestamp 1731220477
transform 1 0 1480 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5601_6
timestamp 1731220477
transform 1 0 1320 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5600_6
timestamp 1731220477
transform 1 0 1152 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5599_6
timestamp 1731220477
transform 1 0 1312 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5598_6
timestamp 1731220477
transform 1 0 1480 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5597_6
timestamp 1731220477
transform 1 0 1640 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5596_6
timestamp 1731220477
transform 1 0 1784 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5595_6
timestamp 1731220477
transform 1 0 1992 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5594_6
timestamp 1731220477
transform 1 0 2136 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5593_6
timestamp 1731220477
transform 1 0 2304 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5592_6
timestamp 1731220477
transform 1 0 2464 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5591_6
timestamp 1731220477
transform 1 0 2376 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5590_6
timestamp 1731220477
transform 1 0 2512 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5589_6
timestamp 1731220477
transform 1 0 2480 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5588_6
timestamp 1731220477
transform 1 0 2616 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5587_6
timestamp 1731220477
transform 1 0 2752 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5586_6
timestamp 1731220477
transform 1 0 2712 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5585_6
timestamp 1731220477
transform 1 0 2512 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5584_6
timestamp 1731220477
transform 1 0 2304 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5583_6
timestamp 1731220477
transform 1 0 2192 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5582_6
timestamp 1731220477
transform 1 0 2472 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5581_6
timestamp 1731220477
transform 1 0 3328 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5580_6
timestamp 1731220477
transform 1 0 2984 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5579_6
timestamp 1731220477
transform 1 0 2664 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5578_6
timestamp 1731220477
transform 1 0 2384 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5577_6
timestamp 1731220477
transform 1 0 2152 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5576_6
timestamp 1731220477
transform 1 0 1992 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5575_6
timestamp 1731220477
transform 1 0 1784 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5574_6
timestamp 1731220477
transform 1 0 1784 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5573_6
timestamp 1731220477
transform 1 0 1544 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5572_6
timestamp 1731220477
transform 1 0 1288 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5571_6
timestamp 1731220477
transform 1 0 1424 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5570_6
timestamp 1731220477
transform 1 0 1584 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5569_6
timestamp 1731220477
transform 1 0 1752 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5568_6
timestamp 1731220477
transform 1 0 1720 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5567_6
timestamp 1731220477
transform 1 0 1584 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5566_6
timestamp 1731220477
transform 1 0 1448 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5565_6
timestamp 1731220477
transform 1 0 1448 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5564_6
timestamp 1731220477
transform 1 0 1280 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5563_6
timestamp 1731220477
transform 1 0 1112 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5562_6
timestamp 1731220477
transform 1 0 1144 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5561_6
timestamp 1731220477
transform 1 0 968 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5560_6
timestamp 1731220477
transform 1 0 784 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5559_6
timestamp 1731220477
transform 1 0 976 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5558_6
timestamp 1731220477
transform 1 0 792 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5557_6
timestamp 1731220477
transform 1 0 592 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5556_6
timestamp 1731220477
transform 1 0 624 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5555_6
timestamp 1731220477
transform 1 0 872 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5554_6
timestamp 1731220477
transform 1 0 1112 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5553_6
timestamp 1731220477
transform 1 0 928 0 -1 3264
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5552_6
timestamp 1731220477
transform 1 0 720 0 -1 3264
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5551_6
timestamp 1731220477
transform 1 0 592 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5550_6
timestamp 1731220477
transform 1 0 864 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5549_6
timestamp 1731220477
transform 1 0 728 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5548_6
timestamp 1731220477
transform 1 0 672 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5547_6
timestamp 1731220477
transform 1 0 536 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5546_6
timestamp 1731220477
transform 1 0 400 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5545_6
timestamp 1731220477
transform 1 0 320 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5544_6
timestamp 1731220477
transform 1 0 456 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5543_6
timestamp 1731220477
transform 1 0 512 0 -1 3264
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5542_6
timestamp 1731220477
transform 1 0 304 0 -1 3264
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5541_6
timestamp 1731220477
transform 1 0 128 0 -1 3264
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5540_6
timestamp 1731220477
transform 1 0 128 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5539_6
timestamp 1731220477
transform 1 0 368 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5538_6
timestamp 1731220477
transform 1 0 144 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5537_6
timestamp 1731220477
transform 1 0 376 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5536_6
timestamp 1731220477
transform 1 0 392 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5535_6
timestamp 1731220477
transform 1 0 592 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5534_6
timestamp 1731220477
transform 1 0 624 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5533_6
timestamp 1731220477
transform 1 0 784 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5532_6
timestamp 1731220477
transform 1 0 944 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5531_6
timestamp 1731220477
transform 1 0 904 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5530_6
timestamp 1731220477
transform 1 0 768 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5529_6
timestamp 1731220477
transform 1 0 1040 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5528_6
timestamp 1731220477
transform 1 0 1176 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5527_6
timestamp 1731220477
transform 1 0 1312 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5526_6
timestamp 1731220477
transform 1 0 1264 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5525_6
timestamp 1731220477
transform 1 0 1104 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5524_6
timestamp 1731220477
transform 1 0 952 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5523_6
timestamp 1731220477
transform 1 0 800 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5522_6
timestamp 1731220477
transform 1 0 656 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5521_6
timestamp 1731220477
transform 1 0 520 0 -1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5520_6
timestamp 1731220477
transform 1 0 1040 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5519_6
timestamp 1731220477
transform 1 0 800 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5518_6
timestamp 1731220477
transform 1 0 560 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5517_6
timestamp 1731220477
transform 1 0 336 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5516_6
timestamp 1731220477
transform 1 0 128 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5515_6
timestamp 1731220477
transform 1 0 800 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5514_6
timestamp 1731220477
transform 1 0 520 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5513_6
timestamp 1731220477
transform 1 0 288 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5512_6
timestamp 1731220477
transform 1 0 128 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5511_6
timestamp 1731220477
transform 1 0 1120 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5510_6
timestamp 1731220477
transform 1 0 1464 0 -1 2304
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5509_6
timestamp 1731220477
transform 1 0 1144 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5508_6
timestamp 1731220477
transform 1 0 480 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5507_6
timestamp 1731220477
transform 1 0 288 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5506_6
timestamp 1731220477
transform 1 0 688 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5505_6
timestamp 1731220477
transform 1 0 912 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5504_6
timestamp 1731220477
transform 1 0 936 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5503_6
timestamp 1731220477
transform 1 0 792 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5502_6
timestamp 1731220477
transform 1 0 648 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5501_6
timestamp 1731220477
transform 1 0 504 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5500_6
timestamp 1731220477
transform 1 0 368 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5499_6
timestamp 1731220477
transform 1 0 232 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5498_6
timestamp 1731220477
transform 1 0 624 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5497_6
timestamp 1731220477
transform 1 0 432 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5496_6
timestamp 1731220477
transform 1 0 232 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5495_6
timestamp 1731220477
transform 1 0 192 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5494_6
timestamp 1731220477
transform 1 0 432 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5493_6
timestamp 1731220477
transform 1 0 360 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5492_6
timestamp 1731220477
transform 1 0 128 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5491_6
timestamp 1731220477
transform 1 0 128 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5490_6
timestamp 1731220477
transform 1 0 296 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5489_6
timestamp 1731220477
transform 1 0 392 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5488_6
timestamp 1731220477
transform 1 0 128 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5487_6
timestamp 1731220477
transform 1 0 128 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5486_6
timestamp 1731220477
transform 1 0 424 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5485_6
timestamp 1731220477
transform 1 0 560 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5484_6
timestamp 1731220477
transform 1 0 328 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5483_6
timestamp 1731220477
transform 1 0 128 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5482_6
timestamp 1731220477
transform 1 0 232 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5481_6
timestamp 1731220477
transform 1 0 408 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5480_6
timestamp 1731220477
transform 1 0 376 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5479_6
timestamp 1731220477
transform 1 0 224 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5478_6
timestamp 1731220477
transform 1 0 624 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5477_6
timestamp 1731220477
transform 1 0 344 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5476_6
timestamp 1731220477
transform 1 0 304 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5475_6
timestamp 1731220477
transform 1 0 128 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5474_6
timestamp 1731220477
transform 1 0 496 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5473_6
timestamp 1731220477
transform 1 0 344 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5472_6
timestamp 1731220477
transform 1 0 128 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5471_6
timestamp 1731220477
transform 1 0 128 0 1 380
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5470_6
timestamp 1731220477
transform 1 0 424 0 1 380
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5469_6
timestamp 1731220477
transform 1 0 520 0 -1 364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5468_6
timestamp 1731220477
transform 1 0 360 0 -1 364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5467_6
timestamp 1731220477
transform 1 0 208 0 -1 364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5466_6
timestamp 1731220477
transform 1 0 144 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5465_6
timestamp 1731220477
transform 1 0 280 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5464_6
timestamp 1731220477
transform 1 0 416 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5463_6
timestamp 1731220477
transform 1 0 552 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5462_6
timestamp 1731220477
transform 1 0 688 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5461_6
timestamp 1731220477
transform 1 0 1096 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5460_6
timestamp 1731220477
transform 1 0 960 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5459_6
timestamp 1731220477
transform 1 0 824 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5458_6
timestamp 1731220477
transform 1 0 680 0 -1 364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5457_6
timestamp 1731220477
transform 1 0 840 0 -1 364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5456_6
timestamp 1731220477
transform 1 0 1000 0 -1 364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5455_6
timestamp 1731220477
transform 1 0 1456 0 1 380
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5454_6
timestamp 1731220477
transform 1 0 1104 0 1 380
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5453_6
timestamp 1731220477
transform 1 0 760 0 1 380
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5452_6
timestamp 1731220477
transform 1 0 568 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5451_6
timestamp 1731220477
transform 1 0 776 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5450_6
timestamp 1731220477
transform 1 0 968 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5449_6
timestamp 1731220477
transform 1 0 856 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5448_6
timestamp 1731220477
transform 1 0 680 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5447_6
timestamp 1731220477
transform 1 0 1024 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5446_6
timestamp 1731220477
transform 1 0 912 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5445_6
timestamp 1731220477
transform 1 0 1208 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5444_6
timestamp 1731220477
transform 1 0 1072 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5443_6
timestamp 1731220477
transform 1 0 888 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5442_6
timestamp 1731220477
transform 1 0 712 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5441_6
timestamp 1731220477
transform 1 0 536 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5440_6
timestamp 1731220477
transform 1 0 584 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5439_6
timestamp 1731220477
transform 1 0 752 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5438_6
timestamp 1731220477
transform 1 0 920 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5437_6
timestamp 1731220477
transform 1 0 800 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5436_6
timestamp 1731220477
transform 1 0 1040 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5435_6
timestamp 1731220477
transform 1 0 1280 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5434_6
timestamp 1731220477
transform 1 0 1064 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5433_6
timestamp 1731220477
transform 1 0 744 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5432_6
timestamp 1731220477
transform 1 0 1392 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5431_6
timestamp 1731220477
transform 1 0 1256 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5430_6
timestamp 1731220477
transform 1 0 968 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5429_6
timestamp 1731220477
transform 1 0 680 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5428_6
timestamp 1731220477
transform 1 0 1048 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5427_6
timestamp 1731220477
transform 1 0 856 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5426_6
timestamp 1731220477
transform 1 0 664 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5425_6
timestamp 1731220477
transform 1 0 480 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5424_6
timestamp 1731220477
transform 1 0 616 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5423_6
timestamp 1731220477
transform 1 0 872 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5422_6
timestamp 1731220477
transform 1 0 1136 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5421_6
timestamp 1731220477
transform 1 0 1128 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5420_6
timestamp 1731220477
transform 1 0 896 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5419_6
timestamp 1731220477
transform 1 0 664 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5418_6
timestamp 1731220477
transform 1 0 1360 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5417_6
timestamp 1731220477
transform 1 0 1152 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5416_6
timestamp 1731220477
transform 1 0 984 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5415_6
timestamp 1731220477
transform 1 0 808 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5414_6
timestamp 1731220477
transform 1 0 1080 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5413_6
timestamp 1731220477
transform 1 0 1224 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5412_6
timestamp 1731220477
transform 1 0 1368 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5411_6
timestamp 1731220477
transform 1 0 1384 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5410_6
timestamp 1731220477
transform 1 0 1632 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5409_6
timestamp 1731220477
transform 1 0 1512 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5408_6
timestamp 1731220477
transform 1 0 1784 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5407_6
timestamp 1731220477
transform 1 0 1648 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5406_6
timestamp 1731220477
transform 1 0 1640 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5405_6
timestamp 1731220477
transform 1 0 1480 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5404_6
timestamp 1731220477
transform 1 0 1320 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5403_6
timestamp 1731220477
transform 1 0 1784 0 1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5402_6
timestamp 1731220477
transform 1 0 1992 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5401_6
timestamp 1731220477
transform 1 0 2128 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5400_6
timestamp 1731220477
transform 1 0 2264 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5399_6
timestamp 1731220477
transform 1 0 2416 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5398_6
timestamp 1731220477
transform 1 0 2576 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5397_6
timestamp 1731220477
transform 1 0 2736 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5396_6
timestamp 1731220477
transform 1 0 2608 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5395_6
timestamp 1731220477
transform 1 0 2448 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5394_6
timestamp 1731220477
transform 1 0 2288 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5393_6
timestamp 1731220477
transform 1 0 2136 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5392_6
timestamp 1731220477
transform 1 0 1992 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5391_6
timestamp 1731220477
transform 1 0 1992 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5390_6
timestamp 1731220477
transform 1 0 2128 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5389_6
timestamp 1731220477
transform 1 0 2264 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5388_6
timestamp 1731220477
transform 1 0 2136 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5387_6
timestamp 1731220477
transform 1 0 2272 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5386_6
timestamp 1731220477
transform 1 0 2408 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5385_6
timestamp 1731220477
transform 1 0 2712 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5384_6
timestamp 1731220477
transform 1 0 2552 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5383_6
timestamp 1731220477
transform 1 0 2400 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5382_6
timestamp 1731220477
transform 1 0 2264 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5381_6
timestamp 1731220477
transform 1 0 2128 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5380_6
timestamp 1731220477
transform 1 0 2688 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5379_6
timestamp 1731220477
transform 1 0 2448 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5378_6
timestamp 1731220477
transform 1 0 2208 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5377_6
timestamp 1731220477
transform 1 0 1992 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5376_6
timestamp 1731220477
transform 1 0 1768 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5375_6
timestamp 1731220477
transform 1 0 1520 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5374_6
timestamp 1731220477
transform 1 0 1720 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5373_6
timestamp 1731220477
transform 1 0 1560 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5372_6
timestamp 1731220477
transform 1 0 1400 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5371_6
timestamp 1731220477
transform 1 0 1240 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5370_6
timestamp 1731220477
transform 1 0 1080 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5369_6
timestamp 1731220477
transform 1 0 1256 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5368_6
timestamp 1731220477
transform 1 0 1440 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5367_6
timestamp 1731220477
transform 1 0 1624 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5366_6
timestamp 1731220477
transform 1 0 1784 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5365_6
timestamp 1731220477
transform 1 0 2016 0 -1 932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5364_6
timestamp 1731220477
transform 1 0 2320 0 -1 932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5363_6
timestamp 1731220477
transform 1 0 2520 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5362_6
timestamp 1731220477
transform 1 0 2248 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5361_6
timestamp 1731220477
transform 1 0 1992 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5360_6
timestamp 1731220477
transform 1 0 1784 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5359_6
timestamp 1731220477
transform 1 0 1504 0 -1 828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5358_6
timestamp 1731220477
transform 1 0 1784 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5357_6
timestamp 1731220477
transform 1 0 1648 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5356_6
timestamp 1731220477
transform 1 0 1488 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5355_6
timestamp 1731220477
transform 1 0 1336 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5354_6
timestamp 1731220477
transform 1 0 1184 0 1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5353_6
timestamp 1731220477
transform 1 0 1144 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5352_6
timestamp 1731220477
transform 1 0 1312 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5351_6
timestamp 1731220477
transform 1 0 1480 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5350_6
timestamp 1731220477
transform 1 0 1640 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5349_6
timestamp 1731220477
transform 1 0 1784 0 -1 604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5348_6
timestamp 1731220477
transform 1 0 1784 0 1 380
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5347_6
timestamp 1731220477
transform 1 0 1992 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5346_6
timestamp 1731220477
transform 1 0 2152 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5345_6
timestamp 1731220477
transform 1 0 2728 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5344_6
timestamp 1731220477
transform 1 0 2536 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5343_6
timestamp 1731220477
transform 1 0 2344 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5342_6
timestamp 1731220477
transform 1 0 2016 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5341_6
timestamp 1731220477
transform 1 0 1992 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5340_6
timestamp 1731220477
transform 1 0 2128 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5339_6
timestamp 1731220477
transform 1 0 2264 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5338_6
timestamp 1731220477
transform 1 0 2400 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5337_6
timestamp 1731220477
transform 1 0 2808 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5336_6
timestamp 1731220477
transform 1 0 2672 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5335_6
timestamp 1731220477
transform 1 0 2536 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5334_6
timestamp 1731220477
transform 1 0 2424 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5333_6
timestamp 1731220477
transform 1 0 2288 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5332_6
timestamp 1731220477
transform 1 0 2152 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5331_6
timestamp 1731220477
transform 1 0 2560 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5330_6
timestamp 1731220477
transform 1 0 2696 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5329_6
timestamp 1731220477
transform 1 0 2944 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5328_6
timestamp 1731220477
transform 1 0 3080 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5327_6
timestamp 1731220477
transform 1 0 3216 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5326_6
timestamp 1731220477
transform 1 0 3624 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5325_6
timestamp 1731220477
transform 1 0 3488 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5324_6
timestamp 1731220477
transform 1 0 3352 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5323_6
timestamp 1731220477
transform 1 0 3104 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5322_6
timestamp 1731220477
transform 1 0 2968 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5321_6
timestamp 1731220477
transform 1 0 2832 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5320_6
timestamp 1731220477
transform 1 0 3240 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5319_6
timestamp 1731220477
transform 1 0 3648 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5318_6
timestamp 1731220477
transform 1 0 3512 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5317_6
timestamp 1731220477
transform 1 0 3376 0 -1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5316_6
timestamp 1731220477
transform 1 0 3296 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5315_6
timestamp 1731220477
transform 1 0 3112 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5314_6
timestamp 1731220477
transform 1 0 2920 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5313_6
timestamp 1731220477
transform 1 0 3480 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5312_6
timestamp 1731220477
transform 1 0 3648 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5311_6
timestamp 1731220477
transform 1 0 3552 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5310_6
timestamp 1731220477
transform 1 0 3416 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5309_6
timestamp 1731220477
transform 1 0 3280 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5308_6
timestamp 1731220477
transform 1 0 3000 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5307_6
timestamp 1731220477
transform 1 0 2768 0 1 708
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5306_6
timestamp 1731220477
transform 1 0 2616 0 -1 932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5305_6
timestamp 1731220477
transform 1 0 2896 0 -1 932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5304_6
timestamp 1731220477
transform 1 0 3088 0 1 960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5303_6
timestamp 1731220477
transform 1 0 2928 0 -1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5302_6
timestamp 1731220477
transform 1 0 2888 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5301_6
timestamp 1731220477
transform 1 0 3072 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5300_6
timestamp 1731220477
transform 1 0 3264 0 1 1208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5299_6
timestamp 1731220477
transform 1 0 3224 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5298_6
timestamp 1731220477
transform 1 0 3088 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5297_6
timestamp 1731220477
transform 1 0 2952 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5296_6
timestamp 1731220477
transform 1 0 2816 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5295_6
timestamp 1731220477
transform 1 0 2680 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5294_6
timestamp 1731220477
transform 1 0 2544 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5293_6
timestamp 1731220477
transform 1 0 2536 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5292_6
timestamp 1731220477
transform 1 0 2400 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5291_6
timestamp 1731220477
transform 1 0 2672 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5290_6
timestamp 1731220477
transform 1 0 2808 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5289_6
timestamp 1731220477
transform 1 0 2944 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5288_6
timestamp 1731220477
transform 1 0 3080 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5287_6
timestamp 1731220477
transform 1 0 3488 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5286_6
timestamp 1731220477
transform 1 0 3352 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5285_6
timestamp 1731220477
transform 1 0 3216 0 1 1444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5284_6
timestamp 1731220477
transform 1 0 3072 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5283_6
timestamp 1731220477
transform 1 0 2912 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5282_6
timestamp 1731220477
transform 1 0 2760 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5281_6
timestamp 1731220477
transform 1 0 3392 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5280_6
timestamp 1731220477
transform 1 0 3232 0 -1 1680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5279_6
timestamp 1731220477
transform 1 0 3200 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5278_6
timestamp 1731220477
transform 1 0 3048 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5277_6
timestamp 1731220477
transform 1 0 2896 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5276_6
timestamp 1731220477
transform 1 0 3648 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5275_6
timestamp 1731220477
transform 1 0 3512 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5274_6
timestamp 1731220477
transform 1 0 3352 0 1 1692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5273_6
timestamp 1731220477
transform 1 0 3240 0 -1 1928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5272_6
timestamp 1731220477
transform 1 0 3104 0 -1 1928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5271_6
timestamp 1731220477
transform 1 0 3376 0 -1 1928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5270_6
timestamp 1731220477
transform 1 0 3512 0 -1 1928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5269_6
timestamp 1731220477
transform 1 0 3648 0 -1 1928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5268_6
timestamp 1731220477
transform 1 0 3856 0 1 1840
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5267_6
timestamp 1731220477
transform 1 0 3856 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5266_6
timestamp 1731220477
transform 1 0 3992 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5265_6
timestamp 1731220477
transform 1 0 4128 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5264_6
timestamp 1731220477
transform 1 0 4264 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5263_6
timestamp 1731220477
transform 1 0 4400 0 -1 2064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5262_6
timestamp 1731220477
transform 1 0 4400 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5261_6
timestamp 1731220477
transform 1 0 4264 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5260_6
timestamp 1731220477
transform 1 0 4128 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5259_6
timestamp 1731220477
transform 1 0 3992 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5258_6
timestamp 1731220477
transform 1 0 3856 0 1 2084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5257_6
timestamp 1731220477
transform 1 0 3856 0 -1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5256_6
timestamp 1731220477
transform 1 0 3648 0 1 2128
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5255_6
timestamp 1731220477
transform 1 0 3648 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5254_6
timestamp 1731220477
transform 1 0 3440 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5253_6
timestamp 1731220477
transform 1 0 3208 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5252_6
timestamp 1731220477
transform 1 0 2976 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5251_6
timestamp 1731220477
transform 1 0 2736 0 -1 2352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5250_6
timestamp 1731220477
transform 1 0 3648 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5249_6
timestamp 1731220477
transform 1 0 3464 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5248_6
timestamp 1731220477
transform 1 0 3280 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5247_6
timestamp 1731220477
transform 1 0 3096 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5246_6
timestamp 1731220477
transform 1 0 2904 0 1 2360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5245_6
timestamp 1731220477
transform 1 0 3432 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5244_6
timestamp 1731220477
transform 1 0 3296 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5243_6
timestamp 1731220477
transform 1 0 3160 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5242_6
timestamp 1731220477
transform 1 0 3024 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5241_6
timestamp 1731220477
transform 1 0 2888 0 -1 2600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5240_6
timestamp 1731220477
transform 1 0 3232 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5239_6
timestamp 1731220477
transform 1 0 3088 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5238_6
timestamp 1731220477
transform 1 0 2944 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5237_6
timestamp 1731220477
transform 1 0 2800 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5236_6
timestamp 1731220477
transform 1 0 2656 0 1 2604
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5235_6
timestamp 1731220477
transform 1 0 2632 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5234_6
timestamp 1731220477
transform 1 0 2800 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5233_6
timestamp 1731220477
transform 1 0 3136 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5232_6
timestamp 1731220477
transform 1 0 2968 0 -1 2828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5231_6
timestamp 1731220477
transform 1 0 2936 0 1 2880
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5230_6
timestamp 1731220477
transform 1 0 2800 0 1 2880
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5229_6
timestamp 1731220477
transform 1 0 2752 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5228_6
timestamp 1731220477
transform 1 0 2616 0 -1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5227_6
timestamp 1731220477
transform 1 0 2984 0 1 3104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5226_6
timestamp 1731220477
transform 1 0 3328 0 -1 3328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5225_6
timestamp 1731220477
transform 1 0 2984 0 -1 3328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5224_6
timestamp 1731220477
transform 1 0 2904 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5223_6
timestamp 1731220477
transform 1 0 2528 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5222_6
timestamp 1731220477
transform 1 0 2344 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5221_6
timestamp 1731220477
transform 1 0 2168 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5220_6
timestamp 1731220477
transform 1 0 2712 0 1 3352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5219_6
timestamp 1731220477
transform 1 0 2752 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5218_6
timestamp 1731220477
transform 1 0 2616 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5217_6
timestamp 1731220477
transform 1 0 2480 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5216_6
timestamp 1731220477
transform 1 0 2344 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5215_6
timestamp 1731220477
transform 1 0 2208 0 -1 3580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5214_6
timestamp 1731220477
transform 1 0 2576 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5213_6
timestamp 1731220477
transform 1 0 2432 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5212_6
timestamp 1731220477
transform 1 0 2288 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5211_6
timestamp 1731220477
transform 1 0 2144 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5210_6
timestamp 1731220477
transform 1 0 2008 0 1 3588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5209_6
timestamp 1731220477
transform 1 0 2688 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5208_6
timestamp 1731220477
transform 1 0 2504 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5207_6
timestamp 1731220477
transform 1 0 2320 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5206_6
timestamp 1731220477
transform 1 0 2144 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5205_6
timestamp 1731220477
transform 1 0 1992 0 -1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5204_6
timestamp 1731220477
transform 1 0 1992 0 1 3820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5203_6
timestamp 1731220477
transform 1 0 1784 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5202_6
timestamp 1731220477
transform 1 0 1784 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5201_6
timestamp 1731220477
transform 1 0 1584 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5200_6
timestamp 1731220477
transform 1 0 1512 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5199_6
timestamp 1731220477
transform 1 0 1648 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5198_6
timestamp 1731220477
transform 1 0 1784 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5197_6
timestamp 1731220477
transform 1 0 1648 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5196_6
timestamp 1731220477
transform 1 0 1784 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5195_6
timestamp 1731220477
transform 1 0 1992 0 1 4148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5194_6
timestamp 1731220477
transform 1 0 1992 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5193_6
timestamp 1731220477
transform 1 0 2168 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5192_6
timestamp 1731220477
transform 1 0 2368 0 -1 4376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5191_6
timestamp 1731220477
transform 1 0 2264 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5190_6
timestamp 1731220477
transform 1 0 2512 0 1 4388
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5189_6
timestamp 1731220477
transform 1 0 2496 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5188_6
timestamp 1731220477
transform 1 0 2232 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5187_6
timestamp 1731220477
transform 1 0 2744 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5186_6
timestamp 1731220477
transform 1 0 2720 0 1 4628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5185_6
timestamp 1731220477
transform 1 0 2544 0 1 4628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5184_6
timestamp 1731220477
transform 1 0 3072 0 -1 4864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5183_6
timestamp 1731220477
transform 1 0 3368 0 -1 4864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5182_6
timestamp 1731220477
transform 1 0 3392 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5181_6
timestamp 1731220477
transform 1 0 3176 0 -1 5104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5180_6
timestamp 1731220477
transform 1 0 2944 0 -1 5104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5179_6
timestamp 1731220477
transform 1 0 3096 0 1 5120
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5178_6
timestamp 1731220477
transform 1 0 3304 0 1 5120
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5177_6
timestamp 1731220477
transform 1 0 3296 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5176_6
timestamp 1731220477
transform 1 0 3088 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5175_6
timestamp 1731220477
transform 1 0 3504 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5174_6
timestamp 1731220477
transform 1 0 3424 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5173_6
timestamp 1731220477
transform 1 0 3184 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5172_6
timestamp 1731220477
transform 1 0 3648 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5171_6
timestamp 1731220477
transform 1 0 3448 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5170_6
timestamp 1731220477
transform 1 0 3232 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5169_6
timestamp 1731220477
transform 1 0 3648 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5168_6
timestamp 1731220477
transform 1 0 3616 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5167_6
timestamp 1731220477
transform 1 0 3440 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5166_6
timestamp 1731220477
transform 1 0 3272 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5165_6
timestamp 1731220477
transform 1 0 3104 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5164_6
timestamp 1731220477
transform 1 0 2928 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5163_6
timestamp 1731220477
transform 1 0 2744 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5162_6
timestamp 1731220477
transform 1 0 3016 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5161_6
timestamp 1731220477
transform 1 0 2800 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5160_6
timestamp 1731220477
transform 1 0 2696 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5159_6
timestamp 1731220477
transform 1 0 2944 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5158_6
timestamp 1731220477
transform 1 0 2888 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5157_6
timestamp 1731220477
transform 1 0 2888 0 1 5120
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5156_6
timestamp 1731220477
transform 1 0 2680 0 1 5120
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5155_6
timestamp 1731220477
transform 1 0 2720 0 -1 5104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5154_6
timestamp 1731220477
transform 1 0 3120 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5153_6
timestamp 1731220477
transform 1 0 2792 0 -1 4864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5152_6
timestamp 1731220477
transform 1 0 2528 0 -1 4864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5151_6
timestamp 1731220477
transform 1 0 2296 0 -1 4864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5150_6
timestamp 1731220477
transform 1 0 2368 0 1 4628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5149_6
timestamp 1731220477
transform 1 0 2192 0 1 4628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5148_6
timestamp 1731220477
transform 1 0 2016 0 1 4628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5147_6
timestamp 1731220477
transform 1 0 1992 0 -1 4624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5146_6
timestamp 1731220477
transform 1 0 1784 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5145_6
timestamp 1731220477
transform 1 0 1568 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5144_6
timestamp 1731220477
transform 1 0 1328 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5143_6
timestamp 1731220477
transform 1 0 1464 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5142_6
timestamp 1731220477
transform 1 0 1688 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5141_6
timestamp 1731220477
transform 1 0 1664 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5140_6
timestamp 1731220477
transform 1 0 1528 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5139_6
timestamp 1731220477
transform 1 0 1392 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5138_6
timestamp 1731220477
transform 1 0 1512 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5137_6
timestamp 1731220477
transform 1 0 1376 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5136_6
timestamp 1731220477
transform 1 0 1376 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5135_6
timestamp 1731220477
transform 1 0 1240 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5134_6
timestamp 1731220477
transform 1 0 1368 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5133_6
timestamp 1731220477
transform 1 0 1152 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5132_6
timestamp 1731220477
transform 1 0 1192 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5131_6
timestamp 1731220477
transform 1 0 1496 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5130_6
timestamp 1731220477
transform 1 0 1312 0 -1 3764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5129_6
timestamp 1731220477
transform 1 0 1032 0 -1 3764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5128_6
timestamp 1731220477
transform 1 0 1208 0 1 3524
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5127_6
timestamp 1731220477
transform 1 0 1064 0 1 3524
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5126_6
timestamp 1731220477
transform 1 0 920 0 1 3524
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5125_6
timestamp 1731220477
transform 1 0 944 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5124_6
timestamp 1731220477
transform 1 0 808 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5123_6
timestamp 1731220477
transform 1 0 776 0 1 3524
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5122_6
timestamp 1731220477
transform 1 0 632 0 1 3524
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5121_6
timestamp 1731220477
transform 1 0 488 0 1 3524
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5120_6
timestamp 1731220477
transform 1 0 488 0 -1 3764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5119_6
timestamp 1731220477
transform 1 0 216 0 -1 3764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5118_6
timestamp 1731220477
transform 1 0 760 0 -1 3764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5117_6
timestamp 1731220477
transform 1 0 896 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5116_6
timestamp 1731220477
transform 1 0 616 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5115_6
timestamp 1731220477
transform 1 0 352 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5114_6
timestamp 1731220477
transform 1 0 128 0 1 3776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5113_6
timestamp 1731220477
transform 1 0 128 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5112_6
timestamp 1731220477
transform 1 0 296 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5111_6
timestamp 1731220477
transform 1 0 504 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5110_6
timestamp 1731220477
transform 1 0 720 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5109_6
timestamp 1731220477
transform 1 0 936 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5108_6
timestamp 1731220477
transform 1 0 832 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5107_6
timestamp 1731220477
transform 1 0 696 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5106_6
timestamp 1731220477
transform 1 0 560 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5105_6
timestamp 1731220477
transform 1 0 1104 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5104_6
timestamp 1731220477
transform 1 0 968 0 1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5103_6
timestamp 1731220477
transform 1 0 832 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5102_6
timestamp 1731220477
transform 1 0 696 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5101_6
timestamp 1731220477
transform 1 0 968 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5100_6
timestamp 1731220477
transform 1 0 1104 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_599_6
timestamp 1731220477
transform 1 0 1240 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_598_6
timestamp 1731220477
transform 1 0 1256 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_597_6
timestamp 1731220477
transform 1 0 1120 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_596_6
timestamp 1731220477
transform 1 0 984 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_595_6
timestamp 1731220477
transform 1 0 848 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_594_6
timestamp 1731220477
transform 1 0 712 0 1 4232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_593_6
timestamp 1731220477
transform 1 0 1248 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_592_6
timestamp 1731220477
transform 1 0 1040 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_591_6
timestamp 1731220477
transform 1 0 840 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_590_6
timestamp 1731220477
transform 1 0 656 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_589_6
timestamp 1731220477
transform 1 0 480 0 -1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_588_6
timestamp 1731220477
transform 1 0 1096 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_587_6
timestamp 1731220477
transform 1 0 872 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_586_6
timestamp 1731220477
transform 1 0 648 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_585_6
timestamp 1731220477
transform 1 0 440 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_584_6
timestamp 1731220477
transform 1 0 248 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_583_6
timestamp 1731220477
transform 1 0 672 0 -1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_582_6
timestamp 1731220477
transform 1 0 536 0 -1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_581_6
timestamp 1731220477
transform 1 0 400 0 -1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_580_6
timestamp 1731220477
transform 1 0 264 0 -1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_579_6
timestamp 1731220477
transform 1 0 128 0 -1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_578_6
timestamp 1731220477
transform 1 0 672 0 1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_577_6
timestamp 1731220477
transform 1 0 536 0 1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_576_6
timestamp 1731220477
transform 1 0 400 0 1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_575_6
timestamp 1731220477
transform 1 0 264 0 1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_574_6
timestamp 1731220477
transform 1 0 128 0 1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_573_6
timestamp 1731220477
transform 1 0 128 0 -1 4936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_572_6
timestamp 1731220477
transform 1 0 264 0 -1 4936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_571_6
timestamp 1731220477
transform 1 0 672 0 -1 4936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_570_6
timestamp 1731220477
transform 1 0 536 0 -1 4936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_569_6
timestamp 1731220477
transform 1 0 400 0 -1 4936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_568_6
timestamp 1731220477
transform 1 0 376 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_567_6
timestamp 1731220477
transform 1 0 152 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_566_6
timestamp 1731220477
transform 1 0 1192 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_565_6
timestamp 1731220477
transform 1 0 896 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_564_6
timestamp 1731220477
transform 1 0 624 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_563_6
timestamp 1731220477
transform 1 0 592 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_562_6
timestamp 1731220477
transform 1 0 416 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_561_6
timestamp 1731220477
transform 1 0 776 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_560_6
timestamp 1731220477
transform 1 0 968 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_559_6
timestamp 1731220477
transform 1 0 1168 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_558_6
timestamp 1731220477
transform 1 0 1184 0 1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_557_6
timestamp 1731220477
transform 1 0 1024 0 1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_556_6
timestamp 1731220477
transform 1 0 872 0 1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_555_6
timestamp 1731220477
transform 1 0 720 0 1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_554_6
timestamp 1731220477
transform 1 0 688 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_553_6
timestamp 1731220477
transform 1 0 824 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_552_6
timestamp 1731220477
transform 1 0 960 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_551_6
timestamp 1731220477
transform 1 0 1096 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_550_6
timestamp 1731220477
transform 1 0 1776 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_549_6
timestamp 1731220477
transform 1 0 1640 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_548_6
timestamp 1731220477
transform 1 0 1504 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_547_6
timestamp 1731220477
transform 1 0 1432 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_546_6
timestamp 1731220477
transform 1 0 1288 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_545_6
timestamp 1731220477
transform 1 0 1720 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_544_6
timestamp 1731220477
transform 1 0 1576 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_543_6
timestamp 1731220477
transform 1 0 1352 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_542_6
timestamp 1731220477
transform 1 0 1576 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_541_6
timestamp 1731220477
transform 1 0 1784 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_540_6
timestamp 1731220477
transform 1 0 1992 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_539_6
timestamp 1731220477
transform 1 0 2168 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_538_6
timestamp 1731220477
transform 1 0 2368 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_537_6
timestamp 1731220477
transform 1 0 2560 0 1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_536_6
timestamp 1731220477
transform 1 0 2576 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_535_6
timestamp 1731220477
transform 1 0 2344 0 -1 5576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_534_6
timestamp 1731220477
transform 1 0 2448 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_533_6
timestamp 1731220477
transform 1 0 2288 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_532_6
timestamp 1731220477
transform 1 0 2688 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_531_6
timestamp 1731220477
transform 1 0 2488 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_530_6
timestamp 1731220477
transform 1 0 2472 0 1 5120
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_529_6
timestamp 1731220477
transform 1 0 2272 0 1 5120
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_528_6
timestamp 1731220477
transform 1 0 2088 0 -1 5104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_527_6
timestamp 1731220477
transform 1 0 2296 0 -1 5104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_526_6
timestamp 1731220477
transform 1 0 2504 0 -1 5104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_525_6
timestamp 1731220477
transform 1 0 2856 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_524_6
timestamp 1731220477
transform 1 0 2616 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_523_6
timestamp 1731220477
transform 1 0 2416 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_522_6
timestamp 1731220477
transform 1 0 2264 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_521_6
timestamp 1731220477
transform 1 0 2128 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_520_6
timestamp 1731220477
transform 1 0 1992 0 1 4872
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_519_6
timestamp 1731220477
transform 1 0 1784 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_518_6
timestamp 1731220477
transform 1 0 1496 0 1 4964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_517_6
timestamp 1731220477
transform 1 0 1368 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_516_6
timestamp 1731220477
transform 1 0 1784 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_515_6
timestamp 1731220477
transform 1 0 1576 0 -1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_514_6
timestamp 1731220477
transform 1 0 1520 0 1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_513_6
timestamp 1731220477
transform 1 0 1352 0 1 5196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_512_6
timestamp 1731220477
transform 1 0 1368 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_511_6
timestamp 1731220477
transform 1 0 1232 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_510_6
timestamp 1731220477
transform 1 0 1144 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_59_6
timestamp 1731220477
transform 1 0 1008 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_58_6
timestamp 1731220477
transform 1 0 872 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_57_6
timestamp 1731220477
transform 1 0 1128 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_56_6
timestamp 1731220477
transform 1 0 912 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_55_6
timestamp 1731220477
transform 1 0 704 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_54_6
timestamp 1731220477
transform 1 0 504 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_53_6
timestamp 1731220477
transform 1 0 312 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_52_6
timestamp 1731220477
transform 1 0 400 0 1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_51_6
timestamp 1731220477
transform 1 0 264 0 1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_50_6
timestamp 1731220477
transform 1 0 128 0 1 5644
box 3 5 132 108
<< end >>
