magic
tech sky130l
timestamp 1731220455
<< m2 >>
rect 110 5705 116 5706
rect 1934 5705 1940 5706
rect 110 5701 111 5705
rect 115 5701 116 5705
rect 110 5700 116 5701
rect 158 5704 164 5705
rect 158 5700 159 5704
rect 163 5700 164 5704
rect 158 5699 164 5700
rect 294 5704 300 5705
rect 294 5700 295 5704
rect 299 5700 300 5704
rect 294 5699 300 5700
rect 430 5704 436 5705
rect 430 5700 431 5704
rect 435 5700 436 5704
rect 430 5699 436 5700
rect 566 5704 572 5705
rect 566 5700 567 5704
rect 571 5700 572 5704
rect 566 5699 572 5700
rect 702 5704 708 5705
rect 702 5700 703 5704
rect 707 5700 708 5704
rect 702 5699 708 5700
rect 838 5704 844 5705
rect 838 5700 839 5704
rect 843 5700 844 5704
rect 838 5699 844 5700
rect 974 5704 980 5705
rect 974 5700 975 5704
rect 979 5700 980 5704
rect 1934 5701 1935 5705
rect 1939 5701 1940 5705
rect 1934 5700 1940 5701
rect 974 5699 980 5700
rect 130 5689 136 5690
rect 110 5688 116 5689
rect 110 5684 111 5688
rect 115 5684 116 5688
rect 130 5685 131 5689
rect 135 5685 136 5689
rect 130 5684 136 5685
rect 266 5689 272 5690
rect 266 5685 267 5689
rect 271 5685 272 5689
rect 266 5684 272 5685
rect 402 5689 408 5690
rect 402 5685 403 5689
rect 407 5685 408 5689
rect 402 5684 408 5685
rect 538 5689 544 5690
rect 538 5685 539 5689
rect 543 5685 544 5689
rect 538 5684 544 5685
rect 674 5689 680 5690
rect 674 5685 675 5689
rect 679 5685 680 5689
rect 674 5684 680 5685
rect 810 5689 816 5690
rect 810 5685 811 5689
rect 815 5685 816 5689
rect 810 5684 816 5685
rect 946 5689 952 5690
rect 946 5685 947 5689
rect 951 5685 952 5689
rect 946 5684 952 5685
rect 1934 5688 1940 5689
rect 1934 5684 1935 5688
rect 1939 5684 1940 5688
rect 110 5683 116 5684
rect 1934 5683 1940 5684
rect 1974 5645 1980 5646
rect 3798 5645 3804 5646
rect 1974 5641 1975 5645
rect 1979 5641 1980 5645
rect 1974 5640 1980 5641
rect 2102 5644 2108 5645
rect 2102 5640 2103 5644
rect 2107 5640 2108 5644
rect 2102 5639 2108 5640
rect 2238 5644 2244 5645
rect 2238 5640 2239 5644
rect 2243 5640 2244 5644
rect 2238 5639 2244 5640
rect 2374 5644 2380 5645
rect 2374 5640 2375 5644
rect 2379 5640 2380 5644
rect 2374 5639 2380 5640
rect 2510 5644 2516 5645
rect 2510 5640 2511 5644
rect 2515 5640 2516 5644
rect 2510 5639 2516 5640
rect 2646 5644 2652 5645
rect 2646 5640 2647 5644
rect 2651 5640 2652 5644
rect 2646 5639 2652 5640
rect 2782 5644 2788 5645
rect 2782 5640 2783 5644
rect 2787 5640 2788 5644
rect 2782 5639 2788 5640
rect 2918 5644 2924 5645
rect 2918 5640 2919 5644
rect 2923 5640 2924 5644
rect 2918 5639 2924 5640
rect 3054 5644 3060 5645
rect 3054 5640 3055 5644
rect 3059 5640 3060 5644
rect 3054 5639 3060 5640
rect 3190 5644 3196 5645
rect 3190 5640 3191 5644
rect 3195 5640 3196 5644
rect 3190 5639 3196 5640
rect 3326 5644 3332 5645
rect 3326 5640 3327 5644
rect 3331 5640 3332 5644
rect 3326 5639 3332 5640
rect 3462 5644 3468 5645
rect 3462 5640 3463 5644
rect 3467 5640 3468 5644
rect 3462 5639 3468 5640
rect 3598 5644 3604 5645
rect 3598 5640 3599 5644
rect 3603 5640 3604 5644
rect 3798 5641 3799 5645
rect 3803 5641 3804 5645
rect 3798 5640 3804 5641
rect 3598 5639 3604 5640
rect 2074 5629 2080 5630
rect 1974 5628 1980 5629
rect 1974 5624 1975 5628
rect 1979 5624 1980 5628
rect 2074 5625 2075 5629
rect 2079 5625 2080 5629
rect 2074 5624 2080 5625
rect 2210 5629 2216 5630
rect 2210 5625 2211 5629
rect 2215 5625 2216 5629
rect 2210 5624 2216 5625
rect 2346 5629 2352 5630
rect 2346 5625 2347 5629
rect 2351 5625 2352 5629
rect 2346 5624 2352 5625
rect 2482 5629 2488 5630
rect 2482 5625 2483 5629
rect 2487 5625 2488 5629
rect 2482 5624 2488 5625
rect 2618 5629 2624 5630
rect 2618 5625 2619 5629
rect 2623 5625 2624 5629
rect 2618 5624 2624 5625
rect 2754 5629 2760 5630
rect 2754 5625 2755 5629
rect 2759 5625 2760 5629
rect 2754 5624 2760 5625
rect 2890 5629 2896 5630
rect 2890 5625 2891 5629
rect 2895 5625 2896 5629
rect 2890 5624 2896 5625
rect 3026 5629 3032 5630
rect 3026 5625 3027 5629
rect 3031 5625 3032 5629
rect 3026 5624 3032 5625
rect 3162 5629 3168 5630
rect 3162 5625 3163 5629
rect 3167 5625 3168 5629
rect 3162 5624 3168 5625
rect 3298 5629 3304 5630
rect 3298 5625 3299 5629
rect 3303 5625 3304 5629
rect 3298 5624 3304 5625
rect 3434 5629 3440 5630
rect 3434 5625 3435 5629
rect 3439 5625 3440 5629
rect 3434 5624 3440 5625
rect 3570 5629 3576 5630
rect 3570 5625 3571 5629
rect 3575 5625 3576 5629
rect 3570 5624 3576 5625
rect 3798 5628 3804 5629
rect 3798 5624 3799 5628
rect 3803 5624 3804 5628
rect 1974 5623 1980 5624
rect 3798 5623 3804 5624
rect 3838 5544 3844 5545
rect 5662 5544 5668 5545
rect 110 5540 116 5541
rect 1934 5540 1940 5541
rect 110 5536 111 5540
rect 115 5536 116 5540
rect 110 5535 116 5536
rect 754 5539 760 5540
rect 754 5535 755 5539
rect 759 5535 760 5539
rect 754 5534 760 5535
rect 890 5539 896 5540
rect 890 5535 891 5539
rect 895 5535 896 5539
rect 890 5534 896 5535
rect 1026 5539 1032 5540
rect 1026 5535 1027 5539
rect 1031 5535 1032 5539
rect 1026 5534 1032 5535
rect 1162 5539 1168 5540
rect 1162 5535 1163 5539
rect 1167 5535 1168 5539
rect 1934 5536 1935 5540
rect 1939 5536 1940 5540
rect 3838 5540 3839 5544
rect 3843 5540 3844 5544
rect 3838 5539 3844 5540
rect 4242 5543 4248 5544
rect 4242 5539 4243 5543
rect 4247 5539 4248 5543
rect 4242 5538 4248 5539
rect 4378 5543 4384 5544
rect 4378 5539 4379 5543
rect 4383 5539 4384 5543
rect 4378 5538 4384 5539
rect 4514 5543 4520 5544
rect 4514 5539 4515 5543
rect 4519 5539 4520 5543
rect 4514 5538 4520 5539
rect 4650 5543 4656 5544
rect 4650 5539 4651 5543
rect 4655 5539 4656 5543
rect 4650 5538 4656 5539
rect 4786 5543 4792 5544
rect 4786 5539 4787 5543
rect 4791 5539 4792 5543
rect 4786 5538 4792 5539
rect 4922 5543 4928 5544
rect 4922 5539 4923 5543
rect 4927 5539 4928 5543
rect 4922 5538 4928 5539
rect 5058 5543 5064 5544
rect 5058 5539 5059 5543
rect 5063 5539 5064 5543
rect 5662 5540 5663 5544
rect 5667 5540 5668 5544
rect 5662 5539 5668 5540
rect 5058 5538 5064 5539
rect 1934 5535 1940 5536
rect 1162 5534 1168 5535
rect 4270 5528 4276 5529
rect 3838 5527 3844 5528
rect 782 5524 788 5525
rect 110 5523 116 5524
rect 110 5519 111 5523
rect 115 5519 116 5523
rect 782 5520 783 5524
rect 787 5520 788 5524
rect 782 5519 788 5520
rect 918 5524 924 5525
rect 918 5520 919 5524
rect 923 5520 924 5524
rect 918 5519 924 5520
rect 1054 5524 1060 5525
rect 1054 5520 1055 5524
rect 1059 5520 1060 5524
rect 1054 5519 1060 5520
rect 1190 5524 1196 5525
rect 1190 5520 1191 5524
rect 1195 5520 1196 5524
rect 1190 5519 1196 5520
rect 1934 5523 1940 5524
rect 1934 5519 1935 5523
rect 1939 5519 1940 5523
rect 3838 5523 3839 5527
rect 3843 5523 3844 5527
rect 4270 5524 4271 5528
rect 4275 5524 4276 5528
rect 4270 5523 4276 5524
rect 4406 5528 4412 5529
rect 4406 5524 4407 5528
rect 4411 5524 4412 5528
rect 4406 5523 4412 5524
rect 4542 5528 4548 5529
rect 4542 5524 4543 5528
rect 4547 5524 4548 5528
rect 4542 5523 4548 5524
rect 4678 5528 4684 5529
rect 4678 5524 4679 5528
rect 4683 5524 4684 5528
rect 4678 5523 4684 5524
rect 4814 5528 4820 5529
rect 4814 5524 4815 5528
rect 4819 5524 4820 5528
rect 4814 5523 4820 5524
rect 4950 5528 4956 5529
rect 4950 5524 4951 5528
rect 4955 5524 4956 5528
rect 4950 5523 4956 5524
rect 5086 5528 5092 5529
rect 5086 5524 5087 5528
rect 5091 5524 5092 5528
rect 5086 5523 5092 5524
rect 5662 5527 5668 5528
rect 5662 5523 5663 5527
rect 5667 5523 5668 5527
rect 3838 5522 3844 5523
rect 5662 5522 5668 5523
rect 110 5518 116 5519
rect 1934 5518 1940 5519
rect 1974 5496 1980 5497
rect 3798 5496 3804 5497
rect 1974 5492 1975 5496
rect 1979 5492 1980 5496
rect 1974 5491 1980 5492
rect 1994 5495 2000 5496
rect 1994 5491 1995 5495
rect 1999 5491 2000 5495
rect 1994 5490 2000 5491
rect 2130 5495 2136 5496
rect 2130 5491 2131 5495
rect 2135 5491 2136 5495
rect 2130 5490 2136 5491
rect 2266 5495 2272 5496
rect 2266 5491 2267 5495
rect 2271 5491 2272 5495
rect 2266 5490 2272 5491
rect 2402 5495 2408 5496
rect 2402 5491 2403 5495
rect 2407 5491 2408 5495
rect 2402 5490 2408 5491
rect 2554 5495 2560 5496
rect 2554 5491 2555 5495
rect 2559 5491 2560 5495
rect 2554 5490 2560 5491
rect 2706 5495 2712 5496
rect 2706 5491 2707 5495
rect 2711 5491 2712 5495
rect 2706 5490 2712 5491
rect 2858 5495 2864 5496
rect 2858 5491 2859 5495
rect 2863 5491 2864 5495
rect 2858 5490 2864 5491
rect 3010 5495 3016 5496
rect 3010 5491 3011 5495
rect 3015 5491 3016 5495
rect 3010 5490 3016 5491
rect 3162 5495 3168 5496
rect 3162 5491 3163 5495
rect 3167 5491 3168 5495
rect 3162 5490 3168 5491
rect 3322 5495 3328 5496
rect 3322 5491 3323 5495
rect 3327 5491 3328 5495
rect 3322 5490 3328 5491
rect 3482 5495 3488 5496
rect 3482 5491 3483 5495
rect 3487 5491 3488 5495
rect 3798 5492 3799 5496
rect 3803 5492 3804 5496
rect 3798 5491 3804 5492
rect 3482 5490 3488 5491
rect 2022 5480 2028 5481
rect 1974 5479 1980 5480
rect 1974 5475 1975 5479
rect 1979 5475 1980 5479
rect 2022 5476 2023 5480
rect 2027 5476 2028 5480
rect 2022 5475 2028 5476
rect 2158 5480 2164 5481
rect 2158 5476 2159 5480
rect 2163 5476 2164 5480
rect 2158 5475 2164 5476
rect 2294 5480 2300 5481
rect 2294 5476 2295 5480
rect 2299 5476 2300 5480
rect 2294 5475 2300 5476
rect 2430 5480 2436 5481
rect 2430 5476 2431 5480
rect 2435 5476 2436 5480
rect 2430 5475 2436 5476
rect 2582 5480 2588 5481
rect 2582 5476 2583 5480
rect 2587 5476 2588 5480
rect 2582 5475 2588 5476
rect 2734 5480 2740 5481
rect 2734 5476 2735 5480
rect 2739 5476 2740 5480
rect 2734 5475 2740 5476
rect 2886 5480 2892 5481
rect 2886 5476 2887 5480
rect 2891 5476 2892 5480
rect 2886 5475 2892 5476
rect 3038 5480 3044 5481
rect 3038 5476 3039 5480
rect 3043 5476 3044 5480
rect 3038 5475 3044 5476
rect 3190 5480 3196 5481
rect 3190 5476 3191 5480
rect 3195 5476 3196 5480
rect 3190 5475 3196 5476
rect 3350 5480 3356 5481
rect 3350 5476 3351 5480
rect 3355 5476 3356 5480
rect 3350 5475 3356 5476
rect 3510 5480 3516 5481
rect 3510 5476 3511 5480
rect 3515 5476 3516 5480
rect 3510 5475 3516 5476
rect 3798 5479 3804 5480
rect 3798 5475 3799 5479
rect 3803 5475 3804 5479
rect 1974 5474 1980 5475
rect 3798 5474 3804 5475
rect 3838 5469 3844 5470
rect 5662 5469 5668 5470
rect 3838 5465 3839 5469
rect 3843 5465 3844 5469
rect 3838 5464 3844 5465
rect 4454 5468 4460 5469
rect 4454 5464 4455 5468
rect 4459 5464 4460 5468
rect 4454 5463 4460 5464
rect 4590 5468 4596 5469
rect 4590 5464 4591 5468
rect 4595 5464 4596 5468
rect 4590 5463 4596 5464
rect 4726 5468 4732 5469
rect 4726 5464 4727 5468
rect 4731 5464 4732 5468
rect 4726 5463 4732 5464
rect 4862 5468 4868 5469
rect 4862 5464 4863 5468
rect 4867 5464 4868 5468
rect 5662 5465 5663 5469
rect 5667 5465 5668 5469
rect 5662 5464 5668 5465
rect 4862 5463 4868 5464
rect 110 5453 116 5454
rect 1934 5453 1940 5454
rect 4426 5453 4432 5454
rect 110 5449 111 5453
rect 115 5449 116 5453
rect 110 5448 116 5449
rect 862 5452 868 5453
rect 862 5448 863 5452
rect 867 5448 868 5452
rect 862 5447 868 5448
rect 998 5452 1004 5453
rect 998 5448 999 5452
rect 1003 5448 1004 5452
rect 998 5447 1004 5448
rect 1134 5452 1140 5453
rect 1134 5448 1135 5452
rect 1139 5448 1140 5452
rect 1134 5447 1140 5448
rect 1270 5452 1276 5453
rect 1270 5448 1271 5452
rect 1275 5448 1276 5452
rect 1270 5447 1276 5448
rect 1406 5452 1412 5453
rect 1406 5448 1407 5452
rect 1411 5448 1412 5452
rect 1406 5447 1412 5448
rect 1542 5452 1548 5453
rect 1542 5448 1543 5452
rect 1547 5448 1548 5452
rect 1542 5447 1548 5448
rect 1678 5452 1684 5453
rect 1678 5448 1679 5452
rect 1683 5448 1684 5452
rect 1678 5447 1684 5448
rect 1814 5452 1820 5453
rect 1814 5448 1815 5452
rect 1819 5448 1820 5452
rect 1934 5449 1935 5453
rect 1939 5449 1940 5453
rect 1934 5448 1940 5449
rect 3838 5452 3844 5453
rect 3838 5448 3839 5452
rect 3843 5448 3844 5452
rect 4426 5449 4427 5453
rect 4431 5449 4432 5453
rect 4426 5448 4432 5449
rect 4562 5453 4568 5454
rect 4562 5449 4563 5453
rect 4567 5449 4568 5453
rect 4562 5448 4568 5449
rect 4698 5453 4704 5454
rect 4698 5449 4699 5453
rect 4703 5449 4704 5453
rect 4698 5448 4704 5449
rect 4834 5453 4840 5454
rect 4834 5449 4835 5453
rect 4839 5449 4840 5453
rect 4834 5448 4840 5449
rect 5662 5452 5668 5453
rect 5662 5448 5663 5452
rect 5667 5448 5668 5452
rect 1814 5447 1820 5448
rect 3838 5447 3844 5448
rect 5662 5447 5668 5448
rect 834 5437 840 5438
rect 110 5436 116 5437
rect 110 5432 111 5436
rect 115 5432 116 5436
rect 834 5433 835 5437
rect 839 5433 840 5437
rect 834 5432 840 5433
rect 970 5437 976 5438
rect 970 5433 971 5437
rect 975 5433 976 5437
rect 970 5432 976 5433
rect 1106 5437 1112 5438
rect 1106 5433 1107 5437
rect 1111 5433 1112 5437
rect 1106 5432 1112 5433
rect 1242 5437 1248 5438
rect 1242 5433 1243 5437
rect 1247 5433 1248 5437
rect 1242 5432 1248 5433
rect 1378 5437 1384 5438
rect 1378 5433 1379 5437
rect 1383 5433 1384 5437
rect 1378 5432 1384 5433
rect 1514 5437 1520 5438
rect 1514 5433 1515 5437
rect 1519 5433 1520 5437
rect 1514 5432 1520 5433
rect 1650 5437 1656 5438
rect 1650 5433 1651 5437
rect 1655 5433 1656 5437
rect 1650 5432 1656 5433
rect 1786 5437 1792 5438
rect 1786 5433 1787 5437
rect 1791 5433 1792 5437
rect 1786 5432 1792 5433
rect 1934 5436 1940 5437
rect 1934 5432 1935 5436
rect 1939 5432 1940 5436
rect 110 5431 116 5432
rect 1934 5431 1940 5432
rect 1974 5409 1980 5410
rect 3798 5409 3804 5410
rect 1974 5405 1975 5409
rect 1979 5405 1980 5409
rect 1974 5404 1980 5405
rect 2830 5408 2836 5409
rect 2830 5404 2831 5408
rect 2835 5404 2836 5408
rect 2830 5403 2836 5404
rect 2966 5408 2972 5409
rect 2966 5404 2967 5408
rect 2971 5404 2972 5408
rect 2966 5403 2972 5404
rect 3102 5408 3108 5409
rect 3102 5404 3103 5408
rect 3107 5404 3108 5408
rect 3102 5403 3108 5404
rect 3238 5408 3244 5409
rect 3238 5404 3239 5408
rect 3243 5404 3244 5408
rect 3798 5405 3799 5409
rect 3803 5405 3804 5409
rect 3798 5404 3804 5405
rect 3238 5403 3244 5404
rect 2802 5393 2808 5394
rect 1974 5392 1980 5393
rect 1974 5388 1975 5392
rect 1979 5388 1980 5392
rect 2802 5389 2803 5393
rect 2807 5389 2808 5393
rect 2802 5388 2808 5389
rect 2938 5393 2944 5394
rect 2938 5389 2939 5393
rect 2943 5389 2944 5393
rect 2938 5388 2944 5389
rect 3074 5393 3080 5394
rect 3074 5389 3075 5393
rect 3079 5389 3080 5393
rect 3074 5388 3080 5389
rect 3210 5393 3216 5394
rect 3210 5389 3211 5393
rect 3215 5389 3216 5393
rect 3210 5388 3216 5389
rect 3798 5392 3804 5393
rect 3798 5388 3799 5392
rect 3803 5388 3804 5392
rect 1974 5387 1980 5388
rect 3798 5387 3804 5388
rect 3838 5320 3844 5321
rect 5662 5320 5668 5321
rect 3838 5316 3839 5320
rect 3843 5316 3844 5320
rect 3838 5315 3844 5316
rect 4282 5319 4288 5320
rect 4282 5315 4283 5319
rect 4287 5315 4288 5319
rect 4282 5314 4288 5315
rect 4482 5319 4488 5320
rect 4482 5315 4483 5319
rect 4487 5315 4488 5319
rect 4482 5314 4488 5315
rect 4698 5319 4704 5320
rect 4698 5315 4699 5319
rect 4703 5315 4704 5319
rect 4698 5314 4704 5315
rect 4930 5319 4936 5320
rect 4930 5315 4931 5319
rect 4935 5315 4936 5319
rect 4930 5314 4936 5315
rect 5170 5319 5176 5320
rect 5170 5315 5171 5319
rect 5175 5315 5176 5319
rect 5170 5314 5176 5315
rect 5418 5319 5424 5320
rect 5418 5315 5419 5319
rect 5423 5315 5424 5319
rect 5662 5316 5663 5320
rect 5667 5316 5668 5320
rect 5662 5315 5668 5316
rect 5418 5314 5424 5315
rect 110 5304 116 5305
rect 1934 5304 1940 5305
rect 4310 5304 4316 5305
rect 110 5300 111 5304
rect 115 5300 116 5304
rect 110 5299 116 5300
rect 426 5303 432 5304
rect 426 5299 427 5303
rect 431 5299 432 5303
rect 426 5298 432 5299
rect 562 5303 568 5304
rect 562 5299 563 5303
rect 567 5299 568 5303
rect 562 5298 568 5299
rect 698 5303 704 5304
rect 698 5299 699 5303
rect 703 5299 704 5303
rect 698 5298 704 5299
rect 834 5303 840 5304
rect 834 5299 835 5303
rect 839 5299 840 5303
rect 834 5298 840 5299
rect 970 5303 976 5304
rect 970 5299 971 5303
rect 975 5299 976 5303
rect 970 5298 976 5299
rect 1106 5303 1112 5304
rect 1106 5299 1107 5303
rect 1111 5299 1112 5303
rect 1106 5298 1112 5299
rect 1242 5303 1248 5304
rect 1242 5299 1243 5303
rect 1247 5299 1248 5303
rect 1242 5298 1248 5299
rect 1378 5303 1384 5304
rect 1378 5299 1379 5303
rect 1383 5299 1384 5303
rect 1378 5298 1384 5299
rect 1514 5303 1520 5304
rect 1514 5299 1515 5303
rect 1519 5299 1520 5303
rect 1514 5298 1520 5299
rect 1650 5303 1656 5304
rect 1650 5299 1651 5303
rect 1655 5299 1656 5303
rect 1650 5298 1656 5299
rect 1786 5303 1792 5304
rect 1786 5299 1787 5303
rect 1791 5299 1792 5303
rect 1934 5300 1935 5304
rect 1939 5300 1940 5304
rect 1934 5299 1940 5300
rect 3838 5303 3844 5304
rect 3838 5299 3839 5303
rect 3843 5299 3844 5303
rect 4310 5300 4311 5304
rect 4315 5300 4316 5304
rect 4310 5299 4316 5300
rect 4510 5304 4516 5305
rect 4510 5300 4511 5304
rect 4515 5300 4516 5304
rect 4510 5299 4516 5300
rect 4726 5304 4732 5305
rect 4726 5300 4727 5304
rect 4731 5300 4732 5304
rect 4726 5299 4732 5300
rect 4958 5304 4964 5305
rect 4958 5300 4959 5304
rect 4963 5300 4964 5304
rect 4958 5299 4964 5300
rect 5198 5304 5204 5305
rect 5198 5300 5199 5304
rect 5203 5300 5204 5304
rect 5198 5299 5204 5300
rect 5446 5304 5452 5305
rect 5446 5300 5447 5304
rect 5451 5300 5452 5304
rect 5446 5299 5452 5300
rect 5662 5303 5668 5304
rect 5662 5299 5663 5303
rect 5667 5299 5668 5303
rect 1786 5298 1792 5299
rect 3838 5298 3844 5299
rect 5662 5298 5668 5299
rect 454 5288 460 5289
rect 110 5287 116 5288
rect 110 5283 111 5287
rect 115 5283 116 5287
rect 454 5284 455 5288
rect 459 5284 460 5288
rect 454 5283 460 5284
rect 590 5288 596 5289
rect 590 5284 591 5288
rect 595 5284 596 5288
rect 590 5283 596 5284
rect 726 5288 732 5289
rect 726 5284 727 5288
rect 731 5284 732 5288
rect 726 5283 732 5284
rect 862 5288 868 5289
rect 862 5284 863 5288
rect 867 5284 868 5288
rect 862 5283 868 5284
rect 998 5288 1004 5289
rect 998 5284 999 5288
rect 1003 5284 1004 5288
rect 998 5283 1004 5284
rect 1134 5288 1140 5289
rect 1134 5284 1135 5288
rect 1139 5284 1140 5288
rect 1134 5283 1140 5284
rect 1270 5288 1276 5289
rect 1270 5284 1271 5288
rect 1275 5284 1276 5288
rect 1270 5283 1276 5284
rect 1406 5288 1412 5289
rect 1406 5284 1407 5288
rect 1411 5284 1412 5288
rect 1406 5283 1412 5284
rect 1542 5288 1548 5289
rect 1542 5284 1543 5288
rect 1547 5284 1548 5288
rect 1542 5283 1548 5284
rect 1678 5288 1684 5289
rect 1678 5284 1679 5288
rect 1683 5284 1684 5288
rect 1678 5283 1684 5284
rect 1814 5288 1820 5289
rect 1814 5284 1815 5288
rect 1819 5284 1820 5288
rect 1814 5283 1820 5284
rect 1934 5287 1940 5288
rect 1934 5283 1935 5287
rect 1939 5283 1940 5287
rect 110 5282 116 5283
rect 1934 5282 1940 5283
rect 110 5229 116 5230
rect 1934 5229 1940 5230
rect 110 5225 111 5229
rect 115 5225 116 5229
rect 110 5224 116 5225
rect 454 5228 460 5229
rect 454 5224 455 5228
rect 459 5224 460 5228
rect 454 5223 460 5224
rect 590 5228 596 5229
rect 590 5224 591 5228
rect 595 5224 596 5228
rect 590 5223 596 5224
rect 726 5228 732 5229
rect 726 5224 727 5228
rect 731 5224 732 5228
rect 726 5223 732 5224
rect 862 5228 868 5229
rect 862 5224 863 5228
rect 867 5224 868 5228
rect 862 5223 868 5224
rect 998 5228 1004 5229
rect 998 5224 999 5228
rect 1003 5224 1004 5228
rect 998 5223 1004 5224
rect 1134 5228 1140 5229
rect 1134 5224 1135 5228
rect 1139 5224 1140 5228
rect 1134 5223 1140 5224
rect 1270 5228 1276 5229
rect 1270 5224 1271 5228
rect 1275 5224 1276 5228
rect 1270 5223 1276 5224
rect 1406 5228 1412 5229
rect 1406 5224 1407 5228
rect 1411 5224 1412 5228
rect 1406 5223 1412 5224
rect 1542 5228 1548 5229
rect 1542 5224 1543 5228
rect 1547 5224 1548 5228
rect 1542 5223 1548 5224
rect 1678 5228 1684 5229
rect 1678 5224 1679 5228
rect 1683 5224 1684 5228
rect 1678 5223 1684 5224
rect 1814 5228 1820 5229
rect 1814 5224 1815 5228
rect 1819 5224 1820 5228
rect 1934 5225 1935 5229
rect 1939 5225 1940 5229
rect 1934 5224 1940 5225
rect 1974 5224 1980 5225
rect 3798 5224 3804 5225
rect 1814 5223 1820 5224
rect 1974 5220 1975 5224
rect 1979 5220 1980 5224
rect 1974 5219 1980 5220
rect 1994 5223 2000 5224
rect 1994 5219 1995 5223
rect 1999 5219 2000 5223
rect 1994 5218 2000 5219
rect 2218 5223 2224 5224
rect 2218 5219 2219 5223
rect 2223 5219 2224 5223
rect 2218 5218 2224 5219
rect 2466 5223 2472 5224
rect 2466 5219 2467 5223
rect 2471 5219 2472 5223
rect 2466 5218 2472 5219
rect 2714 5223 2720 5224
rect 2714 5219 2715 5223
rect 2719 5219 2720 5223
rect 2714 5218 2720 5219
rect 2970 5223 2976 5224
rect 2970 5219 2971 5223
rect 2975 5219 2976 5223
rect 3798 5220 3799 5224
rect 3803 5220 3804 5224
rect 3798 5219 3804 5220
rect 2970 5218 2976 5219
rect 3838 5217 3844 5218
rect 5662 5217 5668 5218
rect 426 5213 432 5214
rect 110 5212 116 5213
rect 110 5208 111 5212
rect 115 5208 116 5212
rect 426 5209 427 5213
rect 431 5209 432 5213
rect 426 5208 432 5209
rect 562 5213 568 5214
rect 562 5209 563 5213
rect 567 5209 568 5213
rect 562 5208 568 5209
rect 698 5213 704 5214
rect 698 5209 699 5213
rect 703 5209 704 5213
rect 698 5208 704 5209
rect 834 5213 840 5214
rect 834 5209 835 5213
rect 839 5209 840 5213
rect 834 5208 840 5209
rect 970 5213 976 5214
rect 970 5209 971 5213
rect 975 5209 976 5213
rect 970 5208 976 5209
rect 1106 5213 1112 5214
rect 1106 5209 1107 5213
rect 1111 5209 1112 5213
rect 1106 5208 1112 5209
rect 1242 5213 1248 5214
rect 1242 5209 1243 5213
rect 1247 5209 1248 5213
rect 1242 5208 1248 5209
rect 1378 5213 1384 5214
rect 1378 5209 1379 5213
rect 1383 5209 1384 5213
rect 1378 5208 1384 5209
rect 1514 5213 1520 5214
rect 1514 5209 1515 5213
rect 1519 5209 1520 5213
rect 1514 5208 1520 5209
rect 1650 5213 1656 5214
rect 1650 5209 1651 5213
rect 1655 5209 1656 5213
rect 1650 5208 1656 5209
rect 1786 5213 1792 5214
rect 3838 5213 3839 5217
rect 3843 5213 3844 5217
rect 1786 5209 1787 5213
rect 1791 5209 1792 5213
rect 1786 5208 1792 5209
rect 1934 5212 1940 5213
rect 3838 5212 3844 5213
rect 3886 5216 3892 5217
rect 3886 5212 3887 5216
rect 3891 5212 3892 5216
rect 1934 5208 1935 5212
rect 1939 5208 1940 5212
rect 3886 5211 3892 5212
rect 4022 5216 4028 5217
rect 4022 5212 4023 5216
rect 4027 5212 4028 5216
rect 4022 5211 4028 5212
rect 4158 5216 4164 5217
rect 4158 5212 4159 5216
rect 4163 5212 4164 5216
rect 4158 5211 4164 5212
rect 4294 5216 4300 5217
rect 4294 5212 4295 5216
rect 4299 5212 4300 5216
rect 4294 5211 4300 5212
rect 4430 5216 4436 5217
rect 4430 5212 4431 5216
rect 4435 5212 4436 5216
rect 4430 5211 4436 5212
rect 4566 5216 4572 5217
rect 4566 5212 4567 5216
rect 4571 5212 4572 5216
rect 4566 5211 4572 5212
rect 4702 5216 4708 5217
rect 4702 5212 4703 5216
rect 4707 5212 4708 5216
rect 4702 5211 4708 5212
rect 4838 5216 4844 5217
rect 4838 5212 4839 5216
rect 4843 5212 4844 5216
rect 4838 5211 4844 5212
rect 4990 5216 4996 5217
rect 4990 5212 4991 5216
rect 4995 5212 4996 5216
rect 4990 5211 4996 5212
rect 5150 5216 5156 5217
rect 5150 5212 5151 5216
rect 5155 5212 5156 5216
rect 5150 5211 5156 5212
rect 5318 5216 5324 5217
rect 5318 5212 5319 5216
rect 5323 5212 5324 5216
rect 5318 5211 5324 5212
rect 5494 5216 5500 5217
rect 5494 5212 5495 5216
rect 5499 5212 5500 5216
rect 5662 5213 5663 5217
rect 5667 5213 5668 5217
rect 5662 5212 5668 5213
rect 5494 5211 5500 5212
rect 2022 5208 2028 5209
rect 110 5207 116 5208
rect 1934 5207 1940 5208
rect 1974 5207 1980 5208
rect 1974 5203 1975 5207
rect 1979 5203 1980 5207
rect 2022 5204 2023 5208
rect 2027 5204 2028 5208
rect 2022 5203 2028 5204
rect 2246 5208 2252 5209
rect 2246 5204 2247 5208
rect 2251 5204 2252 5208
rect 2246 5203 2252 5204
rect 2494 5208 2500 5209
rect 2494 5204 2495 5208
rect 2499 5204 2500 5208
rect 2494 5203 2500 5204
rect 2742 5208 2748 5209
rect 2742 5204 2743 5208
rect 2747 5204 2748 5208
rect 2742 5203 2748 5204
rect 2998 5208 3004 5209
rect 2998 5204 2999 5208
rect 3003 5204 3004 5208
rect 2998 5203 3004 5204
rect 3798 5207 3804 5208
rect 3798 5203 3799 5207
rect 3803 5203 3804 5207
rect 1974 5202 1980 5203
rect 3798 5202 3804 5203
rect 3858 5201 3864 5202
rect 3838 5200 3844 5201
rect 3838 5196 3839 5200
rect 3843 5196 3844 5200
rect 3858 5197 3859 5201
rect 3863 5197 3864 5201
rect 3858 5196 3864 5197
rect 3994 5201 4000 5202
rect 3994 5197 3995 5201
rect 3999 5197 4000 5201
rect 3994 5196 4000 5197
rect 4130 5201 4136 5202
rect 4130 5197 4131 5201
rect 4135 5197 4136 5201
rect 4130 5196 4136 5197
rect 4266 5201 4272 5202
rect 4266 5197 4267 5201
rect 4271 5197 4272 5201
rect 4266 5196 4272 5197
rect 4402 5201 4408 5202
rect 4402 5197 4403 5201
rect 4407 5197 4408 5201
rect 4402 5196 4408 5197
rect 4538 5201 4544 5202
rect 4538 5197 4539 5201
rect 4543 5197 4544 5201
rect 4538 5196 4544 5197
rect 4674 5201 4680 5202
rect 4674 5197 4675 5201
rect 4679 5197 4680 5201
rect 4674 5196 4680 5197
rect 4810 5201 4816 5202
rect 4810 5197 4811 5201
rect 4815 5197 4816 5201
rect 4810 5196 4816 5197
rect 4962 5201 4968 5202
rect 4962 5197 4963 5201
rect 4967 5197 4968 5201
rect 4962 5196 4968 5197
rect 5122 5201 5128 5202
rect 5122 5197 5123 5201
rect 5127 5197 5128 5201
rect 5122 5196 5128 5197
rect 5290 5201 5296 5202
rect 5290 5197 5291 5201
rect 5295 5197 5296 5201
rect 5290 5196 5296 5197
rect 5466 5201 5472 5202
rect 5466 5197 5467 5201
rect 5471 5197 5472 5201
rect 5466 5196 5472 5197
rect 5662 5200 5668 5201
rect 5662 5196 5663 5200
rect 5667 5196 5668 5200
rect 3838 5195 3844 5196
rect 5662 5195 5668 5196
rect 1974 5145 1980 5146
rect 3798 5145 3804 5146
rect 1974 5141 1975 5145
rect 1979 5141 1980 5145
rect 1974 5140 1980 5141
rect 2022 5144 2028 5145
rect 2022 5140 2023 5144
rect 2027 5140 2028 5144
rect 2022 5139 2028 5140
rect 2158 5144 2164 5145
rect 2158 5140 2159 5144
rect 2163 5140 2164 5144
rect 2158 5139 2164 5140
rect 2294 5144 2300 5145
rect 2294 5140 2295 5144
rect 2299 5140 2300 5144
rect 2294 5139 2300 5140
rect 2430 5144 2436 5145
rect 2430 5140 2431 5144
rect 2435 5140 2436 5144
rect 2430 5139 2436 5140
rect 2566 5144 2572 5145
rect 2566 5140 2567 5144
rect 2571 5140 2572 5144
rect 2566 5139 2572 5140
rect 2702 5144 2708 5145
rect 2702 5140 2703 5144
rect 2707 5140 2708 5144
rect 2702 5139 2708 5140
rect 2838 5144 2844 5145
rect 2838 5140 2839 5144
rect 2843 5140 2844 5144
rect 2838 5139 2844 5140
rect 2974 5144 2980 5145
rect 2974 5140 2975 5144
rect 2979 5140 2980 5144
rect 2974 5139 2980 5140
rect 3110 5144 3116 5145
rect 3110 5140 3111 5144
rect 3115 5140 3116 5144
rect 3110 5139 3116 5140
rect 3246 5144 3252 5145
rect 3246 5140 3247 5144
rect 3251 5140 3252 5144
rect 3246 5139 3252 5140
rect 3390 5144 3396 5145
rect 3390 5140 3391 5144
rect 3395 5140 3396 5144
rect 3390 5139 3396 5140
rect 3542 5144 3548 5145
rect 3542 5140 3543 5144
rect 3547 5140 3548 5144
rect 3542 5139 3548 5140
rect 3678 5144 3684 5145
rect 3678 5140 3679 5144
rect 3683 5140 3684 5144
rect 3798 5141 3799 5145
rect 3803 5141 3804 5145
rect 3798 5140 3804 5141
rect 3678 5139 3684 5140
rect 1994 5129 2000 5130
rect 1974 5128 1980 5129
rect 1974 5124 1975 5128
rect 1979 5124 1980 5128
rect 1994 5125 1995 5129
rect 1999 5125 2000 5129
rect 1994 5124 2000 5125
rect 2130 5129 2136 5130
rect 2130 5125 2131 5129
rect 2135 5125 2136 5129
rect 2130 5124 2136 5125
rect 2266 5129 2272 5130
rect 2266 5125 2267 5129
rect 2271 5125 2272 5129
rect 2266 5124 2272 5125
rect 2402 5129 2408 5130
rect 2402 5125 2403 5129
rect 2407 5125 2408 5129
rect 2402 5124 2408 5125
rect 2538 5129 2544 5130
rect 2538 5125 2539 5129
rect 2543 5125 2544 5129
rect 2538 5124 2544 5125
rect 2674 5129 2680 5130
rect 2674 5125 2675 5129
rect 2679 5125 2680 5129
rect 2674 5124 2680 5125
rect 2810 5129 2816 5130
rect 2810 5125 2811 5129
rect 2815 5125 2816 5129
rect 2810 5124 2816 5125
rect 2946 5129 2952 5130
rect 2946 5125 2947 5129
rect 2951 5125 2952 5129
rect 2946 5124 2952 5125
rect 3082 5129 3088 5130
rect 3082 5125 3083 5129
rect 3087 5125 3088 5129
rect 3082 5124 3088 5125
rect 3218 5129 3224 5130
rect 3218 5125 3219 5129
rect 3223 5125 3224 5129
rect 3218 5124 3224 5125
rect 3362 5129 3368 5130
rect 3362 5125 3363 5129
rect 3367 5125 3368 5129
rect 3362 5124 3368 5125
rect 3514 5129 3520 5130
rect 3514 5125 3515 5129
rect 3519 5125 3520 5129
rect 3514 5124 3520 5125
rect 3650 5129 3656 5130
rect 3650 5125 3651 5129
rect 3655 5125 3656 5129
rect 3650 5124 3656 5125
rect 3798 5128 3804 5129
rect 3798 5124 3799 5128
rect 3803 5124 3804 5128
rect 1974 5123 1980 5124
rect 3798 5123 3804 5124
rect 3838 5068 3844 5069
rect 5662 5068 5668 5069
rect 110 5064 116 5065
rect 1934 5064 1940 5065
rect 110 5060 111 5064
rect 115 5060 116 5064
rect 110 5059 116 5060
rect 266 5063 272 5064
rect 266 5059 267 5063
rect 271 5059 272 5063
rect 266 5058 272 5059
rect 402 5063 408 5064
rect 402 5059 403 5063
rect 407 5059 408 5063
rect 402 5058 408 5059
rect 538 5063 544 5064
rect 538 5059 539 5063
rect 543 5059 544 5063
rect 538 5058 544 5059
rect 674 5063 680 5064
rect 674 5059 675 5063
rect 679 5059 680 5063
rect 674 5058 680 5059
rect 810 5063 816 5064
rect 810 5059 811 5063
rect 815 5059 816 5063
rect 810 5058 816 5059
rect 946 5063 952 5064
rect 946 5059 947 5063
rect 951 5059 952 5063
rect 1934 5060 1935 5064
rect 1939 5060 1940 5064
rect 3838 5064 3839 5068
rect 3843 5064 3844 5068
rect 3838 5063 3844 5064
rect 3978 5067 3984 5068
rect 3978 5063 3979 5067
rect 3983 5063 3984 5067
rect 3978 5062 3984 5063
rect 4274 5067 4280 5068
rect 4274 5063 4275 5067
rect 4279 5063 4280 5067
rect 4274 5062 4280 5063
rect 4578 5067 4584 5068
rect 4578 5063 4579 5067
rect 4583 5063 4584 5067
rect 4578 5062 4584 5063
rect 4882 5067 4888 5068
rect 4882 5063 4883 5067
rect 4887 5063 4888 5067
rect 4882 5062 4888 5063
rect 5194 5067 5200 5068
rect 5194 5063 5195 5067
rect 5199 5063 5200 5067
rect 5194 5062 5200 5063
rect 5514 5067 5520 5068
rect 5514 5063 5515 5067
rect 5519 5063 5520 5067
rect 5662 5064 5663 5068
rect 5667 5064 5668 5068
rect 5662 5063 5668 5064
rect 5514 5062 5520 5063
rect 1934 5059 1940 5060
rect 946 5058 952 5059
rect 4006 5052 4012 5053
rect 3838 5051 3844 5052
rect 294 5048 300 5049
rect 110 5047 116 5048
rect 110 5043 111 5047
rect 115 5043 116 5047
rect 294 5044 295 5048
rect 299 5044 300 5048
rect 294 5043 300 5044
rect 430 5048 436 5049
rect 430 5044 431 5048
rect 435 5044 436 5048
rect 430 5043 436 5044
rect 566 5048 572 5049
rect 566 5044 567 5048
rect 571 5044 572 5048
rect 566 5043 572 5044
rect 702 5048 708 5049
rect 702 5044 703 5048
rect 707 5044 708 5048
rect 702 5043 708 5044
rect 838 5048 844 5049
rect 838 5044 839 5048
rect 843 5044 844 5048
rect 838 5043 844 5044
rect 974 5048 980 5049
rect 974 5044 975 5048
rect 979 5044 980 5048
rect 974 5043 980 5044
rect 1934 5047 1940 5048
rect 1934 5043 1935 5047
rect 1939 5043 1940 5047
rect 3838 5047 3839 5051
rect 3843 5047 3844 5051
rect 4006 5048 4007 5052
rect 4011 5048 4012 5052
rect 4006 5047 4012 5048
rect 4302 5052 4308 5053
rect 4302 5048 4303 5052
rect 4307 5048 4308 5052
rect 4302 5047 4308 5048
rect 4606 5052 4612 5053
rect 4606 5048 4607 5052
rect 4611 5048 4612 5052
rect 4606 5047 4612 5048
rect 4910 5052 4916 5053
rect 4910 5048 4911 5052
rect 4915 5048 4916 5052
rect 4910 5047 4916 5048
rect 5222 5052 5228 5053
rect 5222 5048 5223 5052
rect 5227 5048 5228 5052
rect 5222 5047 5228 5048
rect 5542 5052 5548 5053
rect 5542 5048 5543 5052
rect 5547 5048 5548 5052
rect 5542 5047 5548 5048
rect 5662 5051 5668 5052
rect 5662 5047 5663 5051
rect 5667 5047 5668 5051
rect 3838 5046 3844 5047
rect 5662 5046 5668 5047
rect 110 5042 116 5043
rect 1934 5042 1940 5043
rect 1974 4996 1980 4997
rect 3798 4996 3804 4997
rect 1974 4992 1975 4996
rect 1979 4992 1980 4996
rect 1974 4991 1980 4992
rect 3106 4995 3112 4996
rect 3106 4991 3107 4995
rect 3111 4991 3112 4995
rect 3106 4990 3112 4991
rect 3242 4995 3248 4996
rect 3242 4991 3243 4995
rect 3247 4991 3248 4995
rect 3242 4990 3248 4991
rect 3378 4995 3384 4996
rect 3378 4991 3379 4995
rect 3383 4991 3384 4995
rect 3378 4990 3384 4991
rect 3514 4995 3520 4996
rect 3514 4991 3515 4995
rect 3519 4991 3520 4995
rect 3514 4990 3520 4991
rect 3650 4995 3656 4996
rect 3650 4991 3651 4995
rect 3655 4991 3656 4995
rect 3798 4992 3799 4996
rect 3803 4992 3804 4996
rect 3798 4991 3804 4992
rect 3650 4990 3656 4991
rect 3134 4980 3140 4981
rect 1974 4979 1980 4980
rect 110 4977 116 4978
rect 1934 4977 1940 4978
rect 110 4973 111 4977
rect 115 4973 116 4977
rect 110 4972 116 4973
rect 158 4976 164 4977
rect 158 4972 159 4976
rect 163 4972 164 4976
rect 158 4971 164 4972
rect 294 4976 300 4977
rect 294 4972 295 4976
rect 299 4972 300 4976
rect 294 4971 300 4972
rect 430 4976 436 4977
rect 430 4972 431 4976
rect 435 4972 436 4976
rect 430 4971 436 4972
rect 566 4976 572 4977
rect 566 4972 567 4976
rect 571 4972 572 4976
rect 566 4971 572 4972
rect 702 4976 708 4977
rect 702 4972 703 4976
rect 707 4972 708 4976
rect 1934 4973 1935 4977
rect 1939 4973 1940 4977
rect 1974 4975 1975 4979
rect 1979 4975 1980 4979
rect 3134 4976 3135 4980
rect 3139 4976 3140 4980
rect 3134 4975 3140 4976
rect 3270 4980 3276 4981
rect 3270 4976 3271 4980
rect 3275 4976 3276 4980
rect 3270 4975 3276 4976
rect 3406 4980 3412 4981
rect 3406 4976 3407 4980
rect 3411 4976 3412 4980
rect 3406 4975 3412 4976
rect 3542 4980 3548 4981
rect 3542 4976 3543 4980
rect 3547 4976 3548 4980
rect 3542 4975 3548 4976
rect 3678 4980 3684 4981
rect 3678 4976 3679 4980
rect 3683 4976 3684 4980
rect 3678 4975 3684 4976
rect 3798 4979 3804 4980
rect 3798 4975 3799 4979
rect 3803 4975 3804 4979
rect 1974 4974 1980 4975
rect 3798 4974 3804 4975
rect 3838 4977 3844 4978
rect 5662 4977 5668 4978
rect 1934 4972 1940 4973
rect 3838 4973 3839 4977
rect 3843 4973 3844 4977
rect 3838 4972 3844 4973
rect 4862 4976 4868 4977
rect 4862 4972 4863 4976
rect 4867 4972 4868 4976
rect 702 4971 708 4972
rect 4862 4971 4868 4972
rect 4998 4976 5004 4977
rect 4998 4972 4999 4976
rect 5003 4972 5004 4976
rect 4998 4971 5004 4972
rect 5134 4976 5140 4977
rect 5134 4972 5135 4976
rect 5139 4972 5140 4976
rect 5134 4971 5140 4972
rect 5270 4976 5276 4977
rect 5270 4972 5271 4976
rect 5275 4972 5276 4976
rect 5270 4971 5276 4972
rect 5406 4976 5412 4977
rect 5406 4972 5407 4976
rect 5411 4972 5412 4976
rect 5406 4971 5412 4972
rect 5542 4976 5548 4977
rect 5542 4972 5543 4976
rect 5547 4972 5548 4976
rect 5662 4973 5663 4977
rect 5667 4973 5668 4977
rect 5662 4972 5668 4973
rect 5542 4971 5548 4972
rect 130 4961 136 4962
rect 110 4960 116 4961
rect 110 4956 111 4960
rect 115 4956 116 4960
rect 130 4957 131 4961
rect 135 4957 136 4961
rect 130 4956 136 4957
rect 266 4961 272 4962
rect 266 4957 267 4961
rect 271 4957 272 4961
rect 266 4956 272 4957
rect 402 4961 408 4962
rect 402 4957 403 4961
rect 407 4957 408 4961
rect 402 4956 408 4957
rect 538 4961 544 4962
rect 538 4957 539 4961
rect 543 4957 544 4961
rect 538 4956 544 4957
rect 674 4961 680 4962
rect 4834 4961 4840 4962
rect 674 4957 675 4961
rect 679 4957 680 4961
rect 674 4956 680 4957
rect 1934 4960 1940 4961
rect 1934 4956 1935 4960
rect 1939 4956 1940 4960
rect 110 4955 116 4956
rect 1934 4955 1940 4956
rect 3838 4960 3844 4961
rect 3838 4956 3839 4960
rect 3843 4956 3844 4960
rect 4834 4957 4835 4961
rect 4839 4957 4840 4961
rect 4834 4956 4840 4957
rect 4970 4961 4976 4962
rect 4970 4957 4971 4961
rect 4975 4957 4976 4961
rect 4970 4956 4976 4957
rect 5106 4961 5112 4962
rect 5106 4957 5107 4961
rect 5111 4957 5112 4961
rect 5106 4956 5112 4957
rect 5242 4961 5248 4962
rect 5242 4957 5243 4961
rect 5247 4957 5248 4961
rect 5242 4956 5248 4957
rect 5378 4961 5384 4962
rect 5378 4957 5379 4961
rect 5383 4957 5384 4961
rect 5378 4956 5384 4957
rect 5514 4961 5520 4962
rect 5514 4957 5515 4961
rect 5519 4957 5520 4961
rect 5514 4956 5520 4957
rect 5662 4960 5668 4961
rect 5662 4956 5663 4960
rect 5667 4956 5668 4960
rect 3838 4955 3844 4956
rect 5662 4955 5668 4956
rect 1974 4913 1980 4914
rect 3798 4913 3804 4914
rect 1974 4909 1975 4913
rect 1979 4909 1980 4913
rect 1974 4908 1980 4909
rect 3134 4912 3140 4913
rect 3134 4908 3135 4912
rect 3139 4908 3140 4912
rect 3134 4907 3140 4908
rect 3270 4912 3276 4913
rect 3270 4908 3271 4912
rect 3275 4908 3276 4912
rect 3270 4907 3276 4908
rect 3406 4912 3412 4913
rect 3406 4908 3407 4912
rect 3411 4908 3412 4912
rect 3406 4907 3412 4908
rect 3542 4912 3548 4913
rect 3542 4908 3543 4912
rect 3547 4908 3548 4912
rect 3542 4907 3548 4908
rect 3678 4912 3684 4913
rect 3678 4908 3679 4912
rect 3683 4908 3684 4912
rect 3798 4909 3799 4913
rect 3803 4909 3804 4913
rect 3798 4908 3804 4909
rect 3678 4907 3684 4908
rect 3106 4897 3112 4898
rect 1974 4896 1980 4897
rect 1974 4892 1975 4896
rect 1979 4892 1980 4896
rect 3106 4893 3107 4897
rect 3111 4893 3112 4897
rect 3106 4892 3112 4893
rect 3242 4897 3248 4898
rect 3242 4893 3243 4897
rect 3247 4893 3248 4897
rect 3242 4892 3248 4893
rect 3378 4897 3384 4898
rect 3378 4893 3379 4897
rect 3383 4893 3384 4897
rect 3378 4892 3384 4893
rect 3514 4897 3520 4898
rect 3514 4893 3515 4897
rect 3519 4893 3520 4897
rect 3514 4892 3520 4893
rect 3650 4897 3656 4898
rect 3650 4893 3651 4897
rect 3655 4893 3656 4897
rect 3650 4892 3656 4893
rect 3798 4896 3804 4897
rect 3798 4892 3799 4896
rect 3803 4892 3804 4896
rect 1974 4891 1980 4892
rect 3798 4891 3804 4892
rect 110 4820 116 4821
rect 1934 4820 1940 4821
rect 110 4816 111 4820
rect 115 4816 116 4820
rect 110 4815 116 4816
rect 130 4819 136 4820
rect 130 4815 131 4819
rect 135 4815 136 4819
rect 130 4814 136 4815
rect 266 4819 272 4820
rect 266 4815 267 4819
rect 271 4815 272 4819
rect 266 4814 272 4815
rect 402 4819 408 4820
rect 402 4815 403 4819
rect 407 4815 408 4819
rect 402 4814 408 4815
rect 538 4819 544 4820
rect 538 4815 539 4819
rect 543 4815 544 4819
rect 538 4814 544 4815
rect 674 4819 680 4820
rect 674 4815 675 4819
rect 679 4815 680 4819
rect 1934 4816 1935 4820
rect 1939 4816 1940 4820
rect 1934 4815 1940 4816
rect 3838 4816 3844 4817
rect 5662 4816 5668 4817
rect 674 4814 680 4815
rect 3838 4812 3839 4816
rect 3843 4812 3844 4816
rect 3838 4811 3844 4812
rect 4482 4815 4488 4816
rect 4482 4811 4483 4815
rect 4487 4811 4488 4815
rect 4482 4810 4488 4811
rect 4674 4815 4680 4816
rect 4674 4811 4675 4815
rect 4679 4811 4680 4815
rect 4674 4810 4680 4811
rect 4874 4815 4880 4816
rect 4874 4811 4875 4815
rect 4879 4811 4880 4815
rect 4874 4810 4880 4811
rect 5090 4815 5096 4816
rect 5090 4811 5091 4815
rect 5095 4811 5096 4815
rect 5090 4810 5096 4811
rect 5314 4815 5320 4816
rect 5314 4811 5315 4815
rect 5319 4811 5320 4815
rect 5314 4810 5320 4811
rect 5514 4815 5520 4816
rect 5514 4811 5515 4815
rect 5519 4811 5520 4815
rect 5662 4812 5663 4816
rect 5667 4812 5668 4816
rect 5662 4811 5668 4812
rect 5514 4810 5520 4811
rect 158 4804 164 4805
rect 110 4803 116 4804
rect 110 4799 111 4803
rect 115 4799 116 4803
rect 158 4800 159 4804
rect 163 4800 164 4804
rect 158 4799 164 4800
rect 294 4804 300 4805
rect 294 4800 295 4804
rect 299 4800 300 4804
rect 294 4799 300 4800
rect 430 4804 436 4805
rect 430 4800 431 4804
rect 435 4800 436 4804
rect 430 4799 436 4800
rect 566 4804 572 4805
rect 566 4800 567 4804
rect 571 4800 572 4804
rect 566 4799 572 4800
rect 702 4804 708 4805
rect 702 4800 703 4804
rect 707 4800 708 4804
rect 702 4799 708 4800
rect 1934 4803 1940 4804
rect 1934 4799 1935 4803
rect 1939 4799 1940 4803
rect 4510 4800 4516 4801
rect 110 4798 116 4799
rect 1934 4798 1940 4799
rect 3838 4799 3844 4800
rect 3838 4795 3839 4799
rect 3843 4795 3844 4799
rect 4510 4796 4511 4800
rect 4515 4796 4516 4800
rect 4510 4795 4516 4796
rect 4702 4800 4708 4801
rect 4702 4796 4703 4800
rect 4707 4796 4708 4800
rect 4702 4795 4708 4796
rect 4902 4800 4908 4801
rect 4902 4796 4903 4800
rect 4907 4796 4908 4800
rect 4902 4795 4908 4796
rect 5118 4800 5124 4801
rect 5118 4796 5119 4800
rect 5123 4796 5124 4800
rect 5118 4795 5124 4796
rect 5342 4800 5348 4801
rect 5342 4796 5343 4800
rect 5347 4796 5348 4800
rect 5342 4795 5348 4796
rect 5542 4800 5548 4801
rect 5542 4796 5543 4800
rect 5547 4796 5548 4800
rect 5542 4795 5548 4796
rect 5662 4799 5668 4800
rect 5662 4795 5663 4799
rect 5667 4795 5668 4799
rect 3838 4794 3844 4795
rect 5662 4794 5668 4795
rect 110 4741 116 4742
rect 1934 4741 1940 4742
rect 110 4737 111 4741
rect 115 4737 116 4741
rect 110 4736 116 4737
rect 158 4740 164 4741
rect 158 4736 159 4740
rect 163 4736 164 4740
rect 158 4735 164 4736
rect 294 4740 300 4741
rect 294 4736 295 4740
rect 299 4736 300 4740
rect 294 4735 300 4736
rect 430 4740 436 4741
rect 430 4736 431 4740
rect 435 4736 436 4740
rect 430 4735 436 4736
rect 566 4740 572 4741
rect 566 4736 567 4740
rect 571 4736 572 4740
rect 566 4735 572 4736
rect 702 4740 708 4741
rect 702 4736 703 4740
rect 707 4736 708 4740
rect 1934 4737 1935 4741
rect 1939 4737 1940 4741
rect 1934 4736 1940 4737
rect 1974 4736 1980 4737
rect 3798 4736 3804 4737
rect 702 4735 708 4736
rect 1974 4732 1975 4736
rect 1979 4732 1980 4736
rect 1974 4731 1980 4732
rect 3106 4735 3112 4736
rect 3106 4731 3107 4735
rect 3111 4731 3112 4735
rect 3106 4730 3112 4731
rect 3242 4735 3248 4736
rect 3242 4731 3243 4735
rect 3247 4731 3248 4735
rect 3242 4730 3248 4731
rect 3378 4735 3384 4736
rect 3378 4731 3379 4735
rect 3383 4731 3384 4735
rect 3378 4730 3384 4731
rect 3514 4735 3520 4736
rect 3514 4731 3515 4735
rect 3519 4731 3520 4735
rect 3514 4730 3520 4731
rect 3650 4735 3656 4736
rect 3650 4731 3651 4735
rect 3655 4731 3656 4735
rect 3798 4732 3799 4736
rect 3803 4732 3804 4736
rect 3798 4731 3804 4732
rect 3650 4730 3656 4731
rect 130 4725 136 4726
rect 110 4724 116 4725
rect 110 4720 111 4724
rect 115 4720 116 4724
rect 130 4721 131 4725
rect 135 4721 136 4725
rect 130 4720 136 4721
rect 266 4725 272 4726
rect 266 4721 267 4725
rect 271 4721 272 4725
rect 266 4720 272 4721
rect 402 4725 408 4726
rect 402 4721 403 4725
rect 407 4721 408 4725
rect 402 4720 408 4721
rect 538 4725 544 4726
rect 538 4721 539 4725
rect 543 4721 544 4725
rect 538 4720 544 4721
rect 674 4725 680 4726
rect 674 4721 675 4725
rect 679 4721 680 4725
rect 674 4720 680 4721
rect 1934 4724 1940 4725
rect 1934 4720 1935 4724
rect 1939 4720 1940 4724
rect 3838 4721 3844 4722
rect 5662 4721 5668 4722
rect 3134 4720 3140 4721
rect 110 4719 116 4720
rect 1934 4719 1940 4720
rect 1974 4719 1980 4720
rect 1974 4715 1975 4719
rect 1979 4715 1980 4719
rect 3134 4716 3135 4720
rect 3139 4716 3140 4720
rect 3134 4715 3140 4716
rect 3270 4720 3276 4721
rect 3270 4716 3271 4720
rect 3275 4716 3276 4720
rect 3270 4715 3276 4716
rect 3406 4720 3412 4721
rect 3406 4716 3407 4720
rect 3411 4716 3412 4720
rect 3406 4715 3412 4716
rect 3542 4720 3548 4721
rect 3542 4716 3543 4720
rect 3547 4716 3548 4720
rect 3542 4715 3548 4716
rect 3678 4720 3684 4721
rect 3678 4716 3679 4720
rect 3683 4716 3684 4720
rect 3678 4715 3684 4716
rect 3798 4719 3804 4720
rect 3798 4715 3799 4719
rect 3803 4715 3804 4719
rect 3838 4717 3839 4721
rect 3843 4717 3844 4721
rect 3838 4716 3844 4717
rect 4118 4720 4124 4721
rect 4118 4716 4119 4720
rect 4123 4716 4124 4720
rect 4118 4715 4124 4716
rect 4374 4720 4380 4721
rect 4374 4716 4375 4720
rect 4379 4716 4380 4720
rect 4374 4715 4380 4716
rect 4646 4720 4652 4721
rect 4646 4716 4647 4720
rect 4651 4716 4652 4720
rect 4646 4715 4652 4716
rect 4942 4720 4948 4721
rect 4942 4716 4943 4720
rect 4947 4716 4948 4720
rect 4942 4715 4948 4716
rect 5254 4720 5260 4721
rect 5254 4716 5255 4720
rect 5259 4716 5260 4720
rect 5254 4715 5260 4716
rect 5542 4720 5548 4721
rect 5542 4716 5543 4720
rect 5547 4716 5548 4720
rect 5662 4717 5663 4721
rect 5667 4717 5668 4721
rect 5662 4716 5668 4717
rect 5542 4715 5548 4716
rect 1974 4714 1980 4715
rect 3798 4714 3804 4715
rect 4090 4705 4096 4706
rect 3838 4704 3844 4705
rect 3838 4700 3839 4704
rect 3843 4700 3844 4704
rect 4090 4701 4091 4705
rect 4095 4701 4096 4705
rect 4090 4700 4096 4701
rect 4346 4705 4352 4706
rect 4346 4701 4347 4705
rect 4351 4701 4352 4705
rect 4346 4700 4352 4701
rect 4618 4705 4624 4706
rect 4618 4701 4619 4705
rect 4623 4701 4624 4705
rect 4618 4700 4624 4701
rect 4914 4705 4920 4706
rect 4914 4701 4915 4705
rect 4919 4701 4920 4705
rect 4914 4700 4920 4701
rect 5226 4705 5232 4706
rect 5226 4701 5227 4705
rect 5231 4701 5232 4705
rect 5226 4700 5232 4701
rect 5514 4705 5520 4706
rect 5514 4701 5515 4705
rect 5519 4701 5520 4705
rect 5514 4700 5520 4701
rect 5662 4704 5668 4705
rect 5662 4700 5663 4704
rect 5667 4700 5668 4704
rect 3838 4699 3844 4700
rect 5662 4699 5668 4700
rect 1974 4621 1980 4622
rect 3798 4621 3804 4622
rect 1974 4617 1975 4621
rect 1979 4617 1980 4621
rect 1974 4616 1980 4617
rect 2022 4620 2028 4621
rect 2022 4616 2023 4620
rect 2027 4616 2028 4620
rect 2022 4615 2028 4616
rect 2158 4620 2164 4621
rect 2158 4616 2159 4620
rect 2163 4616 2164 4620
rect 2158 4615 2164 4616
rect 2310 4620 2316 4621
rect 2310 4616 2311 4620
rect 2315 4616 2316 4620
rect 2310 4615 2316 4616
rect 2478 4620 2484 4621
rect 2478 4616 2479 4620
rect 2483 4616 2484 4620
rect 2478 4615 2484 4616
rect 2654 4620 2660 4621
rect 2654 4616 2655 4620
rect 2659 4616 2660 4620
rect 2654 4615 2660 4616
rect 2830 4620 2836 4621
rect 2830 4616 2831 4620
rect 2835 4616 2836 4620
rect 2830 4615 2836 4616
rect 3006 4620 3012 4621
rect 3006 4616 3007 4620
rect 3011 4616 3012 4620
rect 3006 4615 3012 4616
rect 3182 4620 3188 4621
rect 3182 4616 3183 4620
rect 3187 4616 3188 4620
rect 3182 4615 3188 4616
rect 3350 4620 3356 4621
rect 3350 4616 3351 4620
rect 3355 4616 3356 4620
rect 3350 4615 3356 4616
rect 3526 4620 3532 4621
rect 3526 4616 3527 4620
rect 3531 4616 3532 4620
rect 3526 4615 3532 4616
rect 3678 4620 3684 4621
rect 3678 4616 3679 4620
rect 3683 4616 3684 4620
rect 3798 4617 3799 4621
rect 3803 4617 3804 4621
rect 3798 4616 3804 4617
rect 3678 4615 3684 4616
rect 1994 4605 2000 4606
rect 1974 4604 1980 4605
rect 1974 4600 1975 4604
rect 1979 4600 1980 4604
rect 1994 4601 1995 4605
rect 1999 4601 2000 4605
rect 1994 4600 2000 4601
rect 2130 4605 2136 4606
rect 2130 4601 2131 4605
rect 2135 4601 2136 4605
rect 2130 4600 2136 4601
rect 2282 4605 2288 4606
rect 2282 4601 2283 4605
rect 2287 4601 2288 4605
rect 2282 4600 2288 4601
rect 2450 4605 2456 4606
rect 2450 4601 2451 4605
rect 2455 4601 2456 4605
rect 2450 4600 2456 4601
rect 2626 4605 2632 4606
rect 2626 4601 2627 4605
rect 2631 4601 2632 4605
rect 2626 4600 2632 4601
rect 2802 4605 2808 4606
rect 2802 4601 2803 4605
rect 2807 4601 2808 4605
rect 2802 4600 2808 4601
rect 2978 4605 2984 4606
rect 2978 4601 2979 4605
rect 2983 4601 2984 4605
rect 2978 4600 2984 4601
rect 3154 4605 3160 4606
rect 3154 4601 3155 4605
rect 3159 4601 3160 4605
rect 3154 4600 3160 4601
rect 3322 4605 3328 4606
rect 3322 4601 3323 4605
rect 3327 4601 3328 4605
rect 3322 4600 3328 4601
rect 3498 4605 3504 4606
rect 3498 4601 3499 4605
rect 3503 4601 3504 4605
rect 3498 4600 3504 4601
rect 3650 4605 3656 4606
rect 3650 4601 3651 4605
rect 3655 4601 3656 4605
rect 3650 4600 3656 4601
rect 3798 4604 3804 4605
rect 3798 4600 3799 4604
rect 3803 4600 3804 4604
rect 1974 4599 1980 4600
rect 3798 4599 3804 4600
rect 110 4584 116 4585
rect 1934 4584 1940 4585
rect 110 4580 111 4584
rect 115 4580 116 4584
rect 110 4579 116 4580
rect 210 4583 216 4584
rect 210 4579 211 4583
rect 215 4579 216 4583
rect 210 4578 216 4579
rect 426 4583 432 4584
rect 426 4579 427 4583
rect 431 4579 432 4583
rect 426 4578 432 4579
rect 666 4583 672 4584
rect 666 4579 667 4583
rect 671 4579 672 4583
rect 666 4578 672 4579
rect 930 4583 936 4584
rect 930 4579 931 4583
rect 935 4579 936 4583
rect 930 4578 936 4579
rect 1218 4583 1224 4584
rect 1218 4579 1219 4583
rect 1223 4579 1224 4583
rect 1218 4578 1224 4579
rect 1514 4583 1520 4584
rect 1514 4579 1515 4583
rect 1519 4579 1520 4583
rect 1514 4578 1520 4579
rect 1786 4583 1792 4584
rect 1786 4579 1787 4583
rect 1791 4579 1792 4583
rect 1934 4580 1935 4584
rect 1939 4580 1940 4584
rect 1934 4579 1940 4580
rect 1786 4578 1792 4579
rect 238 4568 244 4569
rect 110 4567 116 4568
rect 110 4563 111 4567
rect 115 4563 116 4567
rect 238 4564 239 4568
rect 243 4564 244 4568
rect 238 4563 244 4564
rect 454 4568 460 4569
rect 454 4564 455 4568
rect 459 4564 460 4568
rect 454 4563 460 4564
rect 694 4568 700 4569
rect 694 4564 695 4568
rect 699 4564 700 4568
rect 694 4563 700 4564
rect 958 4568 964 4569
rect 958 4564 959 4568
rect 963 4564 964 4568
rect 958 4563 964 4564
rect 1246 4568 1252 4569
rect 1246 4564 1247 4568
rect 1251 4564 1252 4568
rect 1246 4563 1252 4564
rect 1542 4568 1548 4569
rect 1542 4564 1543 4568
rect 1547 4564 1548 4568
rect 1542 4563 1548 4564
rect 1814 4568 1820 4569
rect 1814 4564 1815 4568
rect 1819 4564 1820 4568
rect 1814 4563 1820 4564
rect 1934 4567 1940 4568
rect 1934 4563 1935 4567
rect 1939 4563 1940 4567
rect 110 4562 116 4563
rect 1934 4562 1940 4563
rect 3838 4552 3844 4553
rect 5662 4552 5668 4553
rect 3838 4548 3839 4552
rect 3843 4548 3844 4552
rect 3838 4547 3844 4548
rect 4034 4551 4040 4552
rect 4034 4547 4035 4551
rect 4039 4547 4040 4551
rect 4034 4546 4040 4547
rect 4330 4551 4336 4552
rect 4330 4547 4331 4551
rect 4335 4547 4336 4551
rect 4330 4546 4336 4547
rect 4626 4551 4632 4552
rect 4626 4547 4627 4551
rect 4631 4547 4632 4551
rect 4626 4546 4632 4547
rect 4930 4551 4936 4552
rect 4930 4547 4931 4551
rect 4935 4547 4936 4551
rect 4930 4546 4936 4547
rect 5234 4551 5240 4552
rect 5234 4547 5235 4551
rect 5239 4547 5240 4551
rect 5234 4546 5240 4547
rect 5514 4551 5520 4552
rect 5514 4547 5515 4551
rect 5519 4547 5520 4551
rect 5662 4548 5663 4552
rect 5667 4548 5668 4552
rect 5662 4547 5668 4548
rect 5514 4546 5520 4547
rect 4062 4536 4068 4537
rect 3838 4535 3844 4536
rect 3838 4531 3839 4535
rect 3843 4531 3844 4535
rect 4062 4532 4063 4536
rect 4067 4532 4068 4536
rect 4062 4531 4068 4532
rect 4358 4536 4364 4537
rect 4358 4532 4359 4536
rect 4363 4532 4364 4536
rect 4358 4531 4364 4532
rect 4654 4536 4660 4537
rect 4654 4532 4655 4536
rect 4659 4532 4660 4536
rect 4654 4531 4660 4532
rect 4958 4536 4964 4537
rect 4958 4532 4959 4536
rect 4963 4532 4964 4536
rect 4958 4531 4964 4532
rect 5262 4536 5268 4537
rect 5262 4532 5263 4536
rect 5267 4532 5268 4536
rect 5262 4531 5268 4532
rect 5542 4536 5548 4537
rect 5542 4532 5543 4536
rect 5547 4532 5548 4536
rect 5542 4531 5548 4532
rect 5662 4535 5668 4536
rect 5662 4531 5663 4535
rect 5667 4531 5668 4535
rect 3838 4530 3844 4531
rect 5662 4530 5668 4531
rect 110 4509 116 4510
rect 1934 4509 1940 4510
rect 110 4505 111 4509
rect 115 4505 116 4509
rect 110 4504 116 4505
rect 446 4508 452 4509
rect 446 4504 447 4508
rect 451 4504 452 4508
rect 446 4503 452 4504
rect 622 4508 628 4509
rect 622 4504 623 4508
rect 627 4504 628 4508
rect 622 4503 628 4504
rect 806 4508 812 4509
rect 806 4504 807 4508
rect 811 4504 812 4508
rect 806 4503 812 4504
rect 998 4508 1004 4509
rect 998 4504 999 4508
rect 1003 4504 1004 4508
rect 998 4503 1004 4504
rect 1198 4508 1204 4509
rect 1198 4504 1199 4508
rect 1203 4504 1204 4508
rect 1198 4503 1204 4504
rect 1406 4508 1412 4509
rect 1406 4504 1407 4508
rect 1411 4504 1412 4508
rect 1406 4503 1412 4504
rect 1622 4508 1628 4509
rect 1622 4504 1623 4508
rect 1627 4504 1628 4508
rect 1622 4503 1628 4504
rect 1814 4508 1820 4509
rect 1814 4504 1815 4508
rect 1819 4504 1820 4508
rect 1934 4505 1935 4509
rect 1939 4505 1940 4509
rect 1934 4504 1940 4505
rect 1814 4503 1820 4504
rect 418 4493 424 4494
rect 110 4492 116 4493
rect 110 4488 111 4492
rect 115 4488 116 4492
rect 418 4489 419 4493
rect 423 4489 424 4493
rect 418 4488 424 4489
rect 594 4493 600 4494
rect 594 4489 595 4493
rect 599 4489 600 4493
rect 594 4488 600 4489
rect 778 4493 784 4494
rect 778 4489 779 4493
rect 783 4489 784 4493
rect 778 4488 784 4489
rect 970 4493 976 4494
rect 970 4489 971 4493
rect 975 4489 976 4493
rect 970 4488 976 4489
rect 1170 4493 1176 4494
rect 1170 4489 1171 4493
rect 1175 4489 1176 4493
rect 1170 4488 1176 4489
rect 1378 4493 1384 4494
rect 1378 4489 1379 4493
rect 1383 4489 1384 4493
rect 1378 4488 1384 4489
rect 1594 4493 1600 4494
rect 1594 4489 1595 4493
rect 1599 4489 1600 4493
rect 1594 4488 1600 4489
rect 1786 4493 1792 4494
rect 1786 4489 1787 4493
rect 1791 4489 1792 4493
rect 1786 4488 1792 4489
rect 1934 4492 1940 4493
rect 1934 4488 1935 4492
rect 1939 4488 1940 4492
rect 110 4487 116 4488
rect 1934 4487 1940 4488
rect 1974 4472 1980 4473
rect 3798 4472 3804 4473
rect 1974 4468 1975 4472
rect 1979 4468 1980 4472
rect 1974 4467 1980 4468
rect 1994 4471 2000 4472
rect 1994 4467 1995 4471
rect 1999 4467 2000 4471
rect 1994 4466 2000 4467
rect 2226 4471 2232 4472
rect 2226 4467 2227 4471
rect 2231 4467 2232 4471
rect 2226 4466 2232 4467
rect 2458 4471 2464 4472
rect 2458 4467 2459 4471
rect 2463 4467 2464 4471
rect 2458 4466 2464 4467
rect 2690 4471 2696 4472
rect 2690 4467 2691 4471
rect 2695 4467 2696 4471
rect 2690 4466 2696 4467
rect 2914 4471 2920 4472
rect 2914 4467 2915 4471
rect 2919 4467 2920 4471
rect 2914 4466 2920 4467
rect 3130 4471 3136 4472
rect 3130 4467 3131 4471
rect 3135 4467 3136 4471
rect 3130 4466 3136 4467
rect 3354 4471 3360 4472
rect 3354 4467 3355 4471
rect 3359 4467 3360 4471
rect 3354 4466 3360 4467
rect 3578 4471 3584 4472
rect 3578 4467 3579 4471
rect 3583 4467 3584 4471
rect 3798 4468 3799 4472
rect 3803 4468 3804 4472
rect 3798 4467 3804 4468
rect 3578 4466 3584 4467
rect 3838 4461 3844 4462
rect 5662 4461 5668 4462
rect 3838 4457 3839 4461
rect 3843 4457 3844 4461
rect 2022 4456 2028 4457
rect 1974 4455 1980 4456
rect 1974 4451 1975 4455
rect 1979 4451 1980 4455
rect 2022 4452 2023 4456
rect 2027 4452 2028 4456
rect 2022 4451 2028 4452
rect 2254 4456 2260 4457
rect 2254 4452 2255 4456
rect 2259 4452 2260 4456
rect 2254 4451 2260 4452
rect 2486 4456 2492 4457
rect 2486 4452 2487 4456
rect 2491 4452 2492 4456
rect 2486 4451 2492 4452
rect 2718 4456 2724 4457
rect 2718 4452 2719 4456
rect 2723 4452 2724 4456
rect 2718 4451 2724 4452
rect 2942 4456 2948 4457
rect 2942 4452 2943 4456
rect 2947 4452 2948 4456
rect 2942 4451 2948 4452
rect 3158 4456 3164 4457
rect 3158 4452 3159 4456
rect 3163 4452 3164 4456
rect 3158 4451 3164 4452
rect 3382 4456 3388 4457
rect 3382 4452 3383 4456
rect 3387 4452 3388 4456
rect 3382 4451 3388 4452
rect 3606 4456 3612 4457
rect 3838 4456 3844 4457
rect 4310 4460 4316 4461
rect 4310 4456 4311 4460
rect 4315 4456 4316 4460
rect 3606 4452 3607 4456
rect 3611 4452 3612 4456
rect 3606 4451 3612 4452
rect 3798 4455 3804 4456
rect 4310 4455 4316 4456
rect 4534 4460 4540 4461
rect 4534 4456 4535 4460
rect 4539 4456 4540 4460
rect 4534 4455 4540 4456
rect 4774 4460 4780 4461
rect 4774 4456 4775 4460
rect 4779 4456 4780 4460
rect 4774 4455 4780 4456
rect 5022 4460 5028 4461
rect 5022 4456 5023 4460
rect 5027 4456 5028 4460
rect 5022 4455 5028 4456
rect 5278 4460 5284 4461
rect 5278 4456 5279 4460
rect 5283 4456 5284 4460
rect 5278 4455 5284 4456
rect 5542 4460 5548 4461
rect 5542 4456 5543 4460
rect 5547 4456 5548 4460
rect 5662 4457 5663 4461
rect 5667 4457 5668 4461
rect 5662 4456 5668 4457
rect 5542 4455 5548 4456
rect 3798 4451 3799 4455
rect 3803 4451 3804 4455
rect 1974 4450 1980 4451
rect 3798 4450 3804 4451
rect 4282 4445 4288 4446
rect 3838 4444 3844 4445
rect 3838 4440 3839 4444
rect 3843 4440 3844 4444
rect 4282 4441 4283 4445
rect 4287 4441 4288 4445
rect 4282 4440 4288 4441
rect 4506 4445 4512 4446
rect 4506 4441 4507 4445
rect 4511 4441 4512 4445
rect 4506 4440 4512 4441
rect 4746 4445 4752 4446
rect 4746 4441 4747 4445
rect 4751 4441 4752 4445
rect 4746 4440 4752 4441
rect 4994 4445 5000 4446
rect 4994 4441 4995 4445
rect 4999 4441 5000 4445
rect 4994 4440 5000 4441
rect 5250 4445 5256 4446
rect 5250 4441 5251 4445
rect 5255 4441 5256 4445
rect 5250 4440 5256 4441
rect 5514 4445 5520 4446
rect 5514 4441 5515 4445
rect 5519 4441 5520 4445
rect 5514 4440 5520 4441
rect 5662 4444 5668 4445
rect 5662 4440 5663 4444
rect 5667 4440 5668 4444
rect 3838 4439 3844 4440
rect 5662 4439 5668 4440
rect 1974 4393 1980 4394
rect 3798 4393 3804 4394
rect 1974 4389 1975 4393
rect 1979 4389 1980 4393
rect 1974 4388 1980 4389
rect 2118 4392 2124 4393
rect 2118 4388 2119 4392
rect 2123 4388 2124 4392
rect 2118 4387 2124 4388
rect 2342 4392 2348 4393
rect 2342 4388 2343 4392
rect 2347 4388 2348 4392
rect 2342 4387 2348 4388
rect 2566 4392 2572 4393
rect 2566 4388 2567 4392
rect 2571 4388 2572 4392
rect 2566 4387 2572 4388
rect 2782 4392 2788 4393
rect 2782 4388 2783 4392
rect 2787 4388 2788 4392
rect 2782 4387 2788 4388
rect 2990 4392 2996 4393
rect 2990 4388 2991 4392
rect 2995 4388 2996 4392
rect 2990 4387 2996 4388
rect 3198 4392 3204 4393
rect 3198 4388 3199 4392
rect 3203 4388 3204 4392
rect 3198 4387 3204 4388
rect 3406 4392 3412 4393
rect 3406 4388 3407 4392
rect 3411 4388 3412 4392
rect 3798 4389 3799 4393
rect 3803 4389 3804 4393
rect 3798 4388 3804 4389
rect 3406 4387 3412 4388
rect 2090 4377 2096 4378
rect 1974 4376 1980 4377
rect 1974 4372 1975 4376
rect 1979 4372 1980 4376
rect 2090 4373 2091 4377
rect 2095 4373 2096 4377
rect 2090 4372 2096 4373
rect 2314 4377 2320 4378
rect 2314 4373 2315 4377
rect 2319 4373 2320 4377
rect 2314 4372 2320 4373
rect 2538 4377 2544 4378
rect 2538 4373 2539 4377
rect 2543 4373 2544 4377
rect 2538 4372 2544 4373
rect 2754 4377 2760 4378
rect 2754 4373 2755 4377
rect 2759 4373 2760 4377
rect 2754 4372 2760 4373
rect 2962 4377 2968 4378
rect 2962 4373 2963 4377
rect 2967 4373 2968 4377
rect 2962 4372 2968 4373
rect 3170 4377 3176 4378
rect 3170 4373 3171 4377
rect 3175 4373 3176 4377
rect 3170 4372 3176 4373
rect 3378 4377 3384 4378
rect 3378 4373 3379 4377
rect 3383 4373 3384 4377
rect 3378 4372 3384 4373
rect 3798 4376 3804 4377
rect 3798 4372 3799 4376
rect 3803 4372 3804 4376
rect 1974 4371 1980 4372
rect 3798 4371 3804 4372
rect 110 4356 116 4357
rect 1934 4356 1940 4357
rect 110 4352 111 4356
rect 115 4352 116 4356
rect 110 4351 116 4352
rect 570 4355 576 4356
rect 570 4351 571 4355
rect 575 4351 576 4355
rect 570 4350 576 4351
rect 738 4355 744 4356
rect 738 4351 739 4355
rect 743 4351 744 4355
rect 738 4350 744 4351
rect 914 4355 920 4356
rect 914 4351 915 4355
rect 919 4351 920 4355
rect 914 4350 920 4351
rect 1106 4355 1112 4356
rect 1106 4351 1107 4355
rect 1111 4351 1112 4355
rect 1106 4350 1112 4351
rect 1298 4355 1304 4356
rect 1298 4351 1299 4355
rect 1303 4351 1304 4355
rect 1298 4350 1304 4351
rect 1498 4355 1504 4356
rect 1498 4351 1499 4355
rect 1503 4351 1504 4355
rect 1498 4350 1504 4351
rect 1706 4355 1712 4356
rect 1706 4351 1707 4355
rect 1711 4351 1712 4355
rect 1934 4352 1935 4356
rect 1939 4352 1940 4356
rect 1934 4351 1940 4352
rect 1706 4350 1712 4351
rect 598 4340 604 4341
rect 110 4339 116 4340
rect 110 4335 111 4339
rect 115 4335 116 4339
rect 598 4336 599 4340
rect 603 4336 604 4340
rect 598 4335 604 4336
rect 766 4340 772 4341
rect 766 4336 767 4340
rect 771 4336 772 4340
rect 766 4335 772 4336
rect 942 4340 948 4341
rect 942 4336 943 4340
rect 947 4336 948 4340
rect 942 4335 948 4336
rect 1134 4340 1140 4341
rect 1134 4336 1135 4340
rect 1139 4336 1140 4340
rect 1134 4335 1140 4336
rect 1326 4340 1332 4341
rect 1326 4336 1327 4340
rect 1331 4336 1332 4340
rect 1326 4335 1332 4336
rect 1526 4340 1532 4341
rect 1526 4336 1527 4340
rect 1531 4336 1532 4340
rect 1526 4335 1532 4336
rect 1734 4340 1740 4341
rect 1734 4336 1735 4340
rect 1739 4336 1740 4340
rect 1734 4335 1740 4336
rect 1934 4339 1940 4340
rect 1934 4335 1935 4339
rect 1939 4335 1940 4339
rect 110 4334 116 4335
rect 1934 4334 1940 4335
rect 3838 4292 3844 4293
rect 5662 4292 5668 4293
rect 3838 4288 3839 4292
rect 3843 4288 3844 4292
rect 3838 4287 3844 4288
rect 4514 4291 4520 4292
rect 4514 4287 4515 4291
rect 4519 4287 4520 4291
rect 4514 4286 4520 4287
rect 4690 4291 4696 4292
rect 4690 4287 4691 4291
rect 4695 4287 4696 4291
rect 4690 4286 4696 4287
rect 4874 4291 4880 4292
rect 4874 4287 4875 4291
rect 4879 4287 4880 4291
rect 4874 4286 4880 4287
rect 5066 4291 5072 4292
rect 5066 4287 5067 4291
rect 5071 4287 5072 4291
rect 5066 4286 5072 4287
rect 5266 4291 5272 4292
rect 5266 4287 5267 4291
rect 5271 4287 5272 4291
rect 5266 4286 5272 4287
rect 5466 4291 5472 4292
rect 5466 4287 5467 4291
rect 5471 4287 5472 4291
rect 5662 4288 5663 4292
rect 5667 4288 5668 4292
rect 5662 4287 5668 4288
rect 5466 4286 5472 4287
rect 110 4281 116 4282
rect 1934 4281 1940 4282
rect 110 4277 111 4281
rect 115 4277 116 4281
rect 110 4276 116 4277
rect 654 4280 660 4281
rect 654 4276 655 4280
rect 659 4276 660 4280
rect 654 4275 660 4276
rect 822 4280 828 4281
rect 822 4276 823 4280
rect 827 4276 828 4280
rect 822 4275 828 4276
rect 990 4280 996 4281
rect 990 4276 991 4280
rect 995 4276 996 4280
rect 990 4275 996 4276
rect 1166 4280 1172 4281
rect 1166 4276 1167 4280
rect 1171 4276 1172 4280
rect 1166 4275 1172 4276
rect 1342 4280 1348 4281
rect 1342 4276 1343 4280
rect 1347 4276 1348 4280
rect 1342 4275 1348 4276
rect 1518 4280 1524 4281
rect 1518 4276 1519 4280
rect 1523 4276 1524 4280
rect 1518 4275 1524 4276
rect 1702 4280 1708 4281
rect 1702 4276 1703 4280
rect 1707 4276 1708 4280
rect 1934 4277 1935 4281
rect 1939 4277 1940 4281
rect 1934 4276 1940 4277
rect 4542 4276 4548 4277
rect 1702 4275 1708 4276
rect 3838 4275 3844 4276
rect 3838 4271 3839 4275
rect 3843 4271 3844 4275
rect 4542 4272 4543 4276
rect 4547 4272 4548 4276
rect 4542 4271 4548 4272
rect 4718 4276 4724 4277
rect 4718 4272 4719 4276
rect 4723 4272 4724 4276
rect 4718 4271 4724 4272
rect 4902 4276 4908 4277
rect 4902 4272 4903 4276
rect 4907 4272 4908 4276
rect 4902 4271 4908 4272
rect 5094 4276 5100 4277
rect 5094 4272 5095 4276
rect 5099 4272 5100 4276
rect 5094 4271 5100 4272
rect 5294 4276 5300 4277
rect 5294 4272 5295 4276
rect 5299 4272 5300 4276
rect 5294 4271 5300 4272
rect 5494 4276 5500 4277
rect 5494 4272 5495 4276
rect 5499 4272 5500 4276
rect 5494 4271 5500 4272
rect 5662 4275 5668 4276
rect 5662 4271 5663 4275
rect 5667 4271 5668 4275
rect 3838 4270 3844 4271
rect 5662 4270 5668 4271
rect 626 4265 632 4266
rect 110 4264 116 4265
rect 110 4260 111 4264
rect 115 4260 116 4264
rect 626 4261 627 4265
rect 631 4261 632 4265
rect 626 4260 632 4261
rect 794 4265 800 4266
rect 794 4261 795 4265
rect 799 4261 800 4265
rect 794 4260 800 4261
rect 962 4265 968 4266
rect 962 4261 963 4265
rect 967 4261 968 4265
rect 962 4260 968 4261
rect 1138 4265 1144 4266
rect 1138 4261 1139 4265
rect 1143 4261 1144 4265
rect 1138 4260 1144 4261
rect 1314 4265 1320 4266
rect 1314 4261 1315 4265
rect 1319 4261 1320 4265
rect 1314 4260 1320 4261
rect 1490 4265 1496 4266
rect 1490 4261 1491 4265
rect 1495 4261 1496 4265
rect 1490 4260 1496 4261
rect 1674 4265 1680 4266
rect 1674 4261 1675 4265
rect 1679 4261 1680 4265
rect 1674 4260 1680 4261
rect 1934 4264 1940 4265
rect 1934 4260 1935 4264
rect 1939 4260 1940 4264
rect 110 4259 116 4260
rect 1934 4259 1940 4260
rect 1974 4236 1980 4237
rect 3798 4236 3804 4237
rect 1974 4232 1975 4236
rect 1979 4232 1980 4236
rect 1974 4231 1980 4232
rect 2018 4235 2024 4236
rect 2018 4231 2019 4235
rect 2023 4231 2024 4235
rect 2018 4230 2024 4231
rect 2242 4235 2248 4236
rect 2242 4231 2243 4235
rect 2247 4231 2248 4235
rect 2242 4230 2248 4231
rect 2458 4235 2464 4236
rect 2458 4231 2459 4235
rect 2463 4231 2464 4235
rect 2458 4230 2464 4231
rect 2666 4235 2672 4236
rect 2666 4231 2667 4235
rect 2671 4231 2672 4235
rect 2666 4230 2672 4231
rect 2874 4235 2880 4236
rect 2874 4231 2875 4235
rect 2879 4231 2880 4235
rect 2874 4230 2880 4231
rect 3082 4235 3088 4236
rect 3082 4231 3083 4235
rect 3087 4231 3088 4235
rect 3082 4230 3088 4231
rect 3290 4235 3296 4236
rect 3290 4231 3291 4235
rect 3295 4231 3296 4235
rect 3798 4232 3799 4236
rect 3803 4232 3804 4236
rect 3798 4231 3804 4232
rect 3290 4230 3296 4231
rect 2046 4220 2052 4221
rect 1974 4219 1980 4220
rect 1974 4215 1975 4219
rect 1979 4215 1980 4219
rect 2046 4216 2047 4220
rect 2051 4216 2052 4220
rect 2046 4215 2052 4216
rect 2270 4220 2276 4221
rect 2270 4216 2271 4220
rect 2275 4216 2276 4220
rect 2270 4215 2276 4216
rect 2486 4220 2492 4221
rect 2486 4216 2487 4220
rect 2491 4216 2492 4220
rect 2486 4215 2492 4216
rect 2694 4220 2700 4221
rect 2694 4216 2695 4220
rect 2699 4216 2700 4220
rect 2694 4215 2700 4216
rect 2902 4220 2908 4221
rect 2902 4216 2903 4220
rect 2907 4216 2908 4220
rect 2902 4215 2908 4216
rect 3110 4220 3116 4221
rect 3110 4216 3111 4220
rect 3115 4216 3116 4220
rect 3110 4215 3116 4216
rect 3318 4220 3324 4221
rect 3318 4216 3319 4220
rect 3323 4216 3324 4220
rect 3318 4215 3324 4216
rect 3798 4219 3804 4220
rect 3798 4215 3799 4219
rect 3803 4215 3804 4219
rect 1974 4214 1980 4215
rect 3798 4214 3804 4215
rect 3838 4197 3844 4198
rect 5662 4197 5668 4198
rect 3838 4193 3839 4197
rect 3843 4193 3844 4197
rect 3838 4192 3844 4193
rect 4814 4196 4820 4197
rect 4814 4192 4815 4196
rect 4819 4192 4820 4196
rect 4814 4191 4820 4192
rect 4950 4196 4956 4197
rect 4950 4192 4951 4196
rect 4955 4192 4956 4196
rect 4950 4191 4956 4192
rect 5086 4196 5092 4197
rect 5086 4192 5087 4196
rect 5091 4192 5092 4196
rect 5086 4191 5092 4192
rect 5222 4196 5228 4197
rect 5222 4192 5223 4196
rect 5227 4192 5228 4196
rect 5222 4191 5228 4192
rect 5358 4196 5364 4197
rect 5358 4192 5359 4196
rect 5363 4192 5364 4196
rect 5358 4191 5364 4192
rect 5494 4196 5500 4197
rect 5494 4192 5495 4196
rect 5499 4192 5500 4196
rect 5662 4193 5663 4197
rect 5667 4193 5668 4197
rect 5662 4192 5668 4193
rect 5494 4191 5500 4192
rect 4786 4181 4792 4182
rect 3838 4180 3844 4181
rect 3838 4176 3839 4180
rect 3843 4176 3844 4180
rect 4786 4177 4787 4181
rect 4791 4177 4792 4181
rect 4786 4176 4792 4177
rect 4922 4181 4928 4182
rect 4922 4177 4923 4181
rect 4927 4177 4928 4181
rect 4922 4176 4928 4177
rect 5058 4181 5064 4182
rect 5058 4177 5059 4181
rect 5063 4177 5064 4181
rect 5058 4176 5064 4177
rect 5194 4181 5200 4182
rect 5194 4177 5195 4181
rect 5199 4177 5200 4181
rect 5194 4176 5200 4177
rect 5330 4181 5336 4182
rect 5330 4177 5331 4181
rect 5335 4177 5336 4181
rect 5330 4176 5336 4177
rect 5466 4181 5472 4182
rect 5466 4177 5467 4181
rect 5471 4177 5472 4181
rect 5466 4176 5472 4177
rect 5662 4180 5668 4181
rect 5662 4176 5663 4180
rect 5667 4176 5668 4180
rect 3838 4175 3844 4176
rect 5662 4175 5668 4176
rect 1974 4157 1980 4158
rect 3798 4157 3804 4158
rect 1974 4153 1975 4157
rect 1979 4153 1980 4157
rect 1974 4152 1980 4153
rect 2022 4156 2028 4157
rect 2022 4152 2023 4156
rect 2027 4152 2028 4156
rect 2022 4151 2028 4152
rect 2286 4156 2292 4157
rect 2286 4152 2287 4156
rect 2291 4152 2292 4156
rect 2286 4151 2292 4152
rect 2550 4156 2556 4157
rect 2550 4152 2551 4156
rect 2555 4152 2556 4156
rect 2550 4151 2556 4152
rect 2798 4156 2804 4157
rect 2798 4152 2799 4156
rect 2803 4152 2804 4156
rect 2798 4151 2804 4152
rect 3038 4156 3044 4157
rect 3038 4152 3039 4156
rect 3043 4152 3044 4156
rect 3038 4151 3044 4152
rect 3278 4156 3284 4157
rect 3278 4152 3279 4156
rect 3283 4152 3284 4156
rect 3278 4151 3284 4152
rect 3518 4156 3524 4157
rect 3518 4152 3519 4156
rect 3523 4152 3524 4156
rect 3798 4153 3799 4157
rect 3803 4153 3804 4157
rect 3798 4152 3804 4153
rect 3518 4151 3524 4152
rect 1994 4141 2000 4142
rect 1974 4140 1980 4141
rect 1974 4136 1975 4140
rect 1979 4136 1980 4140
rect 1994 4137 1995 4141
rect 1999 4137 2000 4141
rect 1994 4136 2000 4137
rect 2258 4141 2264 4142
rect 2258 4137 2259 4141
rect 2263 4137 2264 4141
rect 2258 4136 2264 4137
rect 2522 4141 2528 4142
rect 2522 4137 2523 4141
rect 2527 4137 2528 4141
rect 2522 4136 2528 4137
rect 2770 4141 2776 4142
rect 2770 4137 2771 4141
rect 2775 4137 2776 4141
rect 2770 4136 2776 4137
rect 3010 4141 3016 4142
rect 3010 4137 3011 4141
rect 3015 4137 3016 4141
rect 3010 4136 3016 4137
rect 3250 4141 3256 4142
rect 3250 4137 3251 4141
rect 3255 4137 3256 4141
rect 3250 4136 3256 4137
rect 3490 4141 3496 4142
rect 3490 4137 3491 4141
rect 3495 4137 3496 4141
rect 3490 4136 3496 4137
rect 3798 4140 3804 4141
rect 3798 4136 3799 4140
rect 3803 4136 3804 4140
rect 1974 4135 1980 4136
rect 3798 4135 3804 4136
rect 110 4120 116 4121
rect 1934 4120 1940 4121
rect 110 4116 111 4120
rect 115 4116 116 4120
rect 110 4115 116 4116
rect 346 4119 352 4120
rect 346 4115 347 4119
rect 351 4115 352 4119
rect 346 4114 352 4115
rect 514 4119 520 4120
rect 514 4115 515 4119
rect 519 4115 520 4119
rect 514 4114 520 4115
rect 698 4119 704 4120
rect 698 4115 699 4119
rect 703 4115 704 4119
rect 698 4114 704 4115
rect 890 4119 896 4120
rect 890 4115 891 4119
rect 895 4115 896 4119
rect 890 4114 896 4115
rect 1098 4119 1104 4120
rect 1098 4115 1099 4119
rect 1103 4115 1104 4119
rect 1098 4114 1104 4115
rect 1314 4119 1320 4120
rect 1314 4115 1315 4119
rect 1319 4115 1320 4119
rect 1314 4114 1320 4115
rect 1530 4119 1536 4120
rect 1530 4115 1531 4119
rect 1535 4115 1536 4119
rect 1934 4116 1935 4120
rect 1939 4116 1940 4120
rect 1934 4115 1940 4116
rect 1530 4114 1536 4115
rect 374 4104 380 4105
rect 110 4103 116 4104
rect 110 4099 111 4103
rect 115 4099 116 4103
rect 374 4100 375 4104
rect 379 4100 380 4104
rect 374 4099 380 4100
rect 542 4104 548 4105
rect 542 4100 543 4104
rect 547 4100 548 4104
rect 542 4099 548 4100
rect 726 4104 732 4105
rect 726 4100 727 4104
rect 731 4100 732 4104
rect 726 4099 732 4100
rect 918 4104 924 4105
rect 918 4100 919 4104
rect 923 4100 924 4104
rect 918 4099 924 4100
rect 1126 4104 1132 4105
rect 1126 4100 1127 4104
rect 1131 4100 1132 4104
rect 1126 4099 1132 4100
rect 1342 4104 1348 4105
rect 1342 4100 1343 4104
rect 1347 4100 1348 4104
rect 1342 4099 1348 4100
rect 1558 4104 1564 4105
rect 1558 4100 1559 4104
rect 1563 4100 1564 4104
rect 1558 4099 1564 4100
rect 1934 4103 1940 4104
rect 1934 4099 1935 4103
rect 1939 4099 1940 4103
rect 110 4098 116 4099
rect 1934 4098 1940 4099
rect 3838 4044 3844 4045
rect 5662 4044 5668 4045
rect 3838 4040 3839 4044
rect 3843 4040 3844 4044
rect 3838 4039 3844 4040
rect 4938 4043 4944 4044
rect 4938 4039 4939 4043
rect 4943 4039 4944 4043
rect 4938 4038 4944 4039
rect 5074 4043 5080 4044
rect 5074 4039 5075 4043
rect 5079 4039 5080 4043
rect 5074 4038 5080 4039
rect 5210 4043 5216 4044
rect 5210 4039 5211 4043
rect 5215 4039 5216 4043
rect 5210 4038 5216 4039
rect 5346 4043 5352 4044
rect 5346 4039 5347 4043
rect 5351 4039 5352 4043
rect 5346 4038 5352 4039
rect 5482 4043 5488 4044
rect 5482 4039 5483 4043
rect 5487 4039 5488 4043
rect 5662 4040 5663 4044
rect 5667 4040 5668 4044
rect 5662 4039 5668 4040
rect 5482 4038 5488 4039
rect 110 4029 116 4030
rect 1934 4029 1940 4030
rect 110 4025 111 4029
rect 115 4025 116 4029
rect 110 4024 116 4025
rect 230 4028 236 4029
rect 230 4024 231 4028
rect 235 4024 236 4028
rect 230 4023 236 4024
rect 422 4028 428 4029
rect 422 4024 423 4028
rect 427 4024 428 4028
rect 422 4023 428 4024
rect 614 4028 620 4029
rect 614 4024 615 4028
rect 619 4024 620 4028
rect 614 4023 620 4024
rect 806 4028 812 4029
rect 806 4024 807 4028
rect 811 4024 812 4028
rect 806 4023 812 4024
rect 990 4028 996 4029
rect 990 4024 991 4028
rect 995 4024 996 4028
rect 990 4023 996 4024
rect 1166 4028 1172 4029
rect 1166 4024 1167 4028
rect 1171 4024 1172 4028
rect 1166 4023 1172 4024
rect 1334 4028 1340 4029
rect 1334 4024 1335 4028
rect 1339 4024 1340 4028
rect 1334 4023 1340 4024
rect 1502 4028 1508 4029
rect 1502 4024 1503 4028
rect 1507 4024 1508 4028
rect 1502 4023 1508 4024
rect 1670 4028 1676 4029
rect 1670 4024 1671 4028
rect 1675 4024 1676 4028
rect 1670 4023 1676 4024
rect 1814 4028 1820 4029
rect 1814 4024 1815 4028
rect 1819 4024 1820 4028
rect 1934 4025 1935 4029
rect 1939 4025 1940 4029
rect 4966 4028 4972 4029
rect 1934 4024 1940 4025
rect 3838 4027 3844 4028
rect 1814 4023 1820 4024
rect 3838 4023 3839 4027
rect 3843 4023 3844 4027
rect 4966 4024 4967 4028
rect 4971 4024 4972 4028
rect 4966 4023 4972 4024
rect 5102 4028 5108 4029
rect 5102 4024 5103 4028
rect 5107 4024 5108 4028
rect 5102 4023 5108 4024
rect 5238 4028 5244 4029
rect 5238 4024 5239 4028
rect 5243 4024 5244 4028
rect 5238 4023 5244 4024
rect 5374 4028 5380 4029
rect 5374 4024 5375 4028
rect 5379 4024 5380 4028
rect 5374 4023 5380 4024
rect 5510 4028 5516 4029
rect 5510 4024 5511 4028
rect 5515 4024 5516 4028
rect 5510 4023 5516 4024
rect 5662 4027 5668 4028
rect 5662 4023 5663 4027
rect 5667 4023 5668 4027
rect 3838 4022 3844 4023
rect 5662 4022 5668 4023
rect 202 4013 208 4014
rect 110 4012 116 4013
rect 110 4008 111 4012
rect 115 4008 116 4012
rect 202 4009 203 4013
rect 207 4009 208 4013
rect 202 4008 208 4009
rect 394 4013 400 4014
rect 394 4009 395 4013
rect 399 4009 400 4013
rect 394 4008 400 4009
rect 586 4013 592 4014
rect 586 4009 587 4013
rect 591 4009 592 4013
rect 586 4008 592 4009
rect 778 4013 784 4014
rect 778 4009 779 4013
rect 783 4009 784 4013
rect 778 4008 784 4009
rect 962 4013 968 4014
rect 962 4009 963 4013
rect 967 4009 968 4013
rect 962 4008 968 4009
rect 1138 4013 1144 4014
rect 1138 4009 1139 4013
rect 1143 4009 1144 4013
rect 1138 4008 1144 4009
rect 1306 4013 1312 4014
rect 1306 4009 1307 4013
rect 1311 4009 1312 4013
rect 1306 4008 1312 4009
rect 1474 4013 1480 4014
rect 1474 4009 1475 4013
rect 1479 4009 1480 4013
rect 1474 4008 1480 4009
rect 1642 4013 1648 4014
rect 1642 4009 1643 4013
rect 1647 4009 1648 4013
rect 1642 4008 1648 4009
rect 1786 4013 1792 4014
rect 1786 4009 1787 4013
rect 1791 4009 1792 4013
rect 1786 4008 1792 4009
rect 1934 4012 1940 4013
rect 1934 4008 1935 4012
rect 1939 4008 1940 4012
rect 110 4007 116 4008
rect 1934 4007 1940 4008
rect 1974 4008 1980 4009
rect 3798 4008 3804 4009
rect 1974 4004 1975 4008
rect 1979 4004 1980 4008
rect 1974 4003 1980 4004
rect 1994 4007 2000 4008
rect 1994 4003 1995 4007
rect 1999 4003 2000 4007
rect 1994 4002 2000 4003
rect 2282 4007 2288 4008
rect 2282 4003 2283 4007
rect 2287 4003 2288 4007
rect 2282 4002 2288 4003
rect 2586 4007 2592 4008
rect 2586 4003 2587 4007
rect 2591 4003 2592 4007
rect 2586 4002 2592 4003
rect 2874 4007 2880 4008
rect 2874 4003 2875 4007
rect 2879 4003 2880 4007
rect 2874 4002 2880 4003
rect 3162 4007 3168 4008
rect 3162 4003 3163 4007
rect 3167 4003 3168 4007
rect 3162 4002 3168 4003
rect 3450 4007 3456 4008
rect 3450 4003 3451 4007
rect 3455 4003 3456 4007
rect 3798 4004 3799 4008
rect 3803 4004 3804 4008
rect 3798 4003 3804 4004
rect 3450 4002 3456 4003
rect 2022 3992 2028 3993
rect 1974 3991 1980 3992
rect 1974 3987 1975 3991
rect 1979 3987 1980 3991
rect 2022 3988 2023 3992
rect 2027 3988 2028 3992
rect 2022 3987 2028 3988
rect 2310 3992 2316 3993
rect 2310 3988 2311 3992
rect 2315 3988 2316 3992
rect 2310 3987 2316 3988
rect 2614 3992 2620 3993
rect 2614 3988 2615 3992
rect 2619 3988 2620 3992
rect 2614 3987 2620 3988
rect 2902 3992 2908 3993
rect 2902 3988 2903 3992
rect 2907 3988 2908 3992
rect 2902 3987 2908 3988
rect 3190 3992 3196 3993
rect 3190 3988 3191 3992
rect 3195 3988 3196 3992
rect 3190 3987 3196 3988
rect 3478 3992 3484 3993
rect 3478 3988 3479 3992
rect 3483 3988 3484 3992
rect 3478 3987 3484 3988
rect 3798 3991 3804 3992
rect 3798 3987 3799 3991
rect 3803 3987 3804 3991
rect 1974 3986 1980 3987
rect 3798 3986 3804 3987
rect 3838 3961 3844 3962
rect 5662 3961 5668 3962
rect 3838 3957 3839 3961
rect 3843 3957 3844 3961
rect 3838 3956 3844 3957
rect 4830 3960 4836 3961
rect 4830 3956 4831 3960
rect 4835 3956 4836 3960
rect 4830 3955 4836 3956
rect 4966 3960 4972 3961
rect 4966 3956 4967 3960
rect 4971 3956 4972 3960
rect 4966 3955 4972 3956
rect 5110 3960 5116 3961
rect 5110 3956 5111 3960
rect 5115 3956 5116 3960
rect 5110 3955 5116 3956
rect 5254 3960 5260 3961
rect 5254 3956 5255 3960
rect 5259 3956 5260 3960
rect 5254 3955 5260 3956
rect 5406 3960 5412 3961
rect 5406 3956 5407 3960
rect 5411 3956 5412 3960
rect 5406 3955 5412 3956
rect 5542 3960 5548 3961
rect 5542 3956 5543 3960
rect 5547 3956 5548 3960
rect 5662 3957 5663 3961
rect 5667 3957 5668 3961
rect 5662 3956 5668 3957
rect 5542 3955 5548 3956
rect 4802 3945 4808 3946
rect 3838 3944 3844 3945
rect 3838 3940 3839 3944
rect 3843 3940 3844 3944
rect 4802 3941 4803 3945
rect 4807 3941 4808 3945
rect 4802 3940 4808 3941
rect 4938 3945 4944 3946
rect 4938 3941 4939 3945
rect 4943 3941 4944 3945
rect 4938 3940 4944 3941
rect 5082 3945 5088 3946
rect 5082 3941 5083 3945
rect 5087 3941 5088 3945
rect 5082 3940 5088 3941
rect 5226 3945 5232 3946
rect 5226 3941 5227 3945
rect 5231 3941 5232 3945
rect 5226 3940 5232 3941
rect 5378 3945 5384 3946
rect 5378 3941 5379 3945
rect 5383 3941 5384 3945
rect 5378 3940 5384 3941
rect 5514 3945 5520 3946
rect 5514 3941 5515 3945
rect 5519 3941 5520 3945
rect 5514 3940 5520 3941
rect 5662 3944 5668 3945
rect 5662 3940 5663 3944
rect 5667 3940 5668 3944
rect 3838 3939 3844 3940
rect 5662 3939 5668 3940
rect 1974 3913 1980 3914
rect 3798 3913 3804 3914
rect 1974 3909 1975 3913
rect 1979 3909 1980 3913
rect 1974 3908 1980 3909
rect 2670 3912 2676 3913
rect 2670 3908 2671 3912
rect 2675 3908 2676 3912
rect 2670 3907 2676 3908
rect 2806 3912 2812 3913
rect 2806 3908 2807 3912
rect 2811 3908 2812 3912
rect 2806 3907 2812 3908
rect 2942 3912 2948 3913
rect 2942 3908 2943 3912
rect 2947 3908 2948 3912
rect 2942 3907 2948 3908
rect 3078 3912 3084 3913
rect 3078 3908 3079 3912
rect 3083 3908 3084 3912
rect 3078 3907 3084 3908
rect 3214 3912 3220 3913
rect 3214 3908 3215 3912
rect 3219 3908 3220 3912
rect 3798 3909 3799 3913
rect 3803 3909 3804 3913
rect 3798 3908 3804 3909
rect 3214 3907 3220 3908
rect 2642 3897 2648 3898
rect 1974 3896 1980 3897
rect 1974 3892 1975 3896
rect 1979 3892 1980 3896
rect 2642 3893 2643 3897
rect 2647 3893 2648 3897
rect 2642 3892 2648 3893
rect 2778 3897 2784 3898
rect 2778 3893 2779 3897
rect 2783 3893 2784 3897
rect 2778 3892 2784 3893
rect 2914 3897 2920 3898
rect 2914 3893 2915 3897
rect 2919 3893 2920 3897
rect 2914 3892 2920 3893
rect 3050 3897 3056 3898
rect 3050 3893 3051 3897
rect 3055 3893 3056 3897
rect 3050 3892 3056 3893
rect 3186 3897 3192 3898
rect 3186 3893 3187 3897
rect 3191 3893 3192 3897
rect 3186 3892 3192 3893
rect 3798 3896 3804 3897
rect 3798 3892 3799 3896
rect 3803 3892 3804 3896
rect 1974 3891 1980 3892
rect 3798 3891 3804 3892
rect 110 3880 116 3881
rect 1934 3880 1940 3881
rect 110 3876 111 3880
rect 115 3876 116 3880
rect 110 3875 116 3876
rect 250 3879 256 3880
rect 250 3875 251 3879
rect 255 3875 256 3879
rect 250 3874 256 3875
rect 450 3879 456 3880
rect 450 3875 451 3879
rect 455 3875 456 3879
rect 450 3874 456 3875
rect 642 3879 648 3880
rect 642 3875 643 3879
rect 647 3875 648 3879
rect 642 3874 648 3875
rect 826 3879 832 3880
rect 826 3875 827 3879
rect 831 3875 832 3879
rect 826 3874 832 3875
rect 1002 3879 1008 3880
rect 1002 3875 1003 3879
rect 1007 3875 1008 3879
rect 1002 3874 1008 3875
rect 1170 3879 1176 3880
rect 1170 3875 1171 3879
rect 1175 3875 1176 3879
rect 1170 3874 1176 3875
rect 1330 3879 1336 3880
rect 1330 3875 1331 3879
rect 1335 3875 1336 3879
rect 1330 3874 1336 3875
rect 1490 3879 1496 3880
rect 1490 3875 1491 3879
rect 1495 3875 1496 3879
rect 1490 3874 1496 3875
rect 1650 3879 1656 3880
rect 1650 3875 1651 3879
rect 1655 3875 1656 3879
rect 1650 3874 1656 3875
rect 1786 3879 1792 3880
rect 1786 3875 1787 3879
rect 1791 3875 1792 3879
rect 1934 3876 1935 3880
rect 1939 3876 1940 3880
rect 1934 3875 1940 3876
rect 1786 3874 1792 3875
rect 278 3864 284 3865
rect 110 3863 116 3864
rect 110 3859 111 3863
rect 115 3859 116 3863
rect 278 3860 279 3864
rect 283 3860 284 3864
rect 278 3859 284 3860
rect 478 3864 484 3865
rect 478 3860 479 3864
rect 483 3860 484 3864
rect 478 3859 484 3860
rect 670 3864 676 3865
rect 670 3860 671 3864
rect 675 3860 676 3864
rect 670 3859 676 3860
rect 854 3864 860 3865
rect 854 3860 855 3864
rect 859 3860 860 3864
rect 854 3859 860 3860
rect 1030 3864 1036 3865
rect 1030 3860 1031 3864
rect 1035 3860 1036 3864
rect 1030 3859 1036 3860
rect 1198 3864 1204 3865
rect 1198 3860 1199 3864
rect 1203 3860 1204 3864
rect 1198 3859 1204 3860
rect 1358 3864 1364 3865
rect 1358 3860 1359 3864
rect 1363 3860 1364 3864
rect 1358 3859 1364 3860
rect 1518 3864 1524 3865
rect 1518 3860 1519 3864
rect 1523 3860 1524 3864
rect 1518 3859 1524 3860
rect 1678 3864 1684 3865
rect 1678 3860 1679 3864
rect 1683 3860 1684 3864
rect 1678 3859 1684 3860
rect 1814 3864 1820 3865
rect 1814 3860 1815 3864
rect 1819 3860 1820 3864
rect 1814 3859 1820 3860
rect 1934 3863 1940 3864
rect 1934 3859 1935 3863
rect 1939 3859 1940 3863
rect 110 3858 116 3859
rect 1934 3858 1940 3859
rect 110 3805 116 3806
rect 1934 3805 1940 3806
rect 110 3801 111 3805
rect 115 3801 116 3805
rect 110 3800 116 3801
rect 310 3804 316 3805
rect 310 3800 311 3804
rect 315 3800 316 3804
rect 310 3799 316 3800
rect 510 3804 516 3805
rect 510 3800 511 3804
rect 515 3800 516 3804
rect 510 3799 516 3800
rect 734 3804 740 3805
rect 734 3800 735 3804
rect 739 3800 740 3804
rect 734 3799 740 3800
rect 990 3804 996 3805
rect 990 3800 991 3804
rect 995 3800 996 3804
rect 990 3799 996 3800
rect 1262 3804 1268 3805
rect 1262 3800 1263 3804
rect 1267 3800 1268 3804
rect 1262 3799 1268 3800
rect 1550 3804 1556 3805
rect 1550 3800 1551 3804
rect 1555 3800 1556 3804
rect 1550 3799 1556 3800
rect 1814 3804 1820 3805
rect 1814 3800 1815 3804
rect 1819 3800 1820 3804
rect 1934 3801 1935 3805
rect 1939 3801 1940 3805
rect 1934 3800 1940 3801
rect 1814 3799 1820 3800
rect 3838 3792 3844 3793
rect 5662 3792 5668 3793
rect 282 3789 288 3790
rect 110 3788 116 3789
rect 110 3784 111 3788
rect 115 3784 116 3788
rect 282 3785 283 3789
rect 287 3785 288 3789
rect 282 3784 288 3785
rect 482 3789 488 3790
rect 482 3785 483 3789
rect 487 3785 488 3789
rect 482 3784 488 3785
rect 706 3789 712 3790
rect 706 3785 707 3789
rect 711 3785 712 3789
rect 706 3784 712 3785
rect 962 3789 968 3790
rect 962 3785 963 3789
rect 967 3785 968 3789
rect 962 3784 968 3785
rect 1234 3789 1240 3790
rect 1234 3785 1235 3789
rect 1239 3785 1240 3789
rect 1234 3784 1240 3785
rect 1522 3789 1528 3790
rect 1522 3785 1523 3789
rect 1527 3785 1528 3789
rect 1522 3784 1528 3785
rect 1786 3789 1792 3790
rect 1786 3785 1787 3789
rect 1791 3785 1792 3789
rect 1786 3784 1792 3785
rect 1934 3788 1940 3789
rect 1934 3784 1935 3788
rect 1939 3784 1940 3788
rect 3838 3788 3839 3792
rect 3843 3788 3844 3792
rect 3838 3787 3844 3788
rect 4498 3791 4504 3792
rect 4498 3787 4499 3791
rect 4503 3787 4504 3791
rect 4498 3786 4504 3787
rect 4674 3791 4680 3792
rect 4674 3787 4675 3791
rect 4679 3787 4680 3791
rect 4674 3786 4680 3787
rect 4874 3791 4880 3792
rect 4874 3787 4875 3791
rect 4879 3787 4880 3791
rect 4874 3786 4880 3787
rect 5090 3791 5096 3792
rect 5090 3787 5091 3791
rect 5095 3787 5096 3791
rect 5090 3786 5096 3787
rect 5314 3791 5320 3792
rect 5314 3787 5315 3791
rect 5319 3787 5320 3791
rect 5314 3786 5320 3787
rect 5514 3791 5520 3792
rect 5514 3787 5515 3791
rect 5519 3787 5520 3791
rect 5662 3788 5663 3792
rect 5667 3788 5668 3792
rect 5662 3787 5668 3788
rect 5514 3786 5520 3787
rect 110 3783 116 3784
rect 1934 3783 1940 3784
rect 4526 3776 4532 3777
rect 3838 3775 3844 3776
rect 3838 3771 3839 3775
rect 3843 3771 3844 3775
rect 4526 3772 4527 3776
rect 4531 3772 4532 3776
rect 4526 3771 4532 3772
rect 4702 3776 4708 3777
rect 4702 3772 4703 3776
rect 4707 3772 4708 3776
rect 4702 3771 4708 3772
rect 4902 3776 4908 3777
rect 4902 3772 4903 3776
rect 4907 3772 4908 3776
rect 4902 3771 4908 3772
rect 5118 3776 5124 3777
rect 5118 3772 5119 3776
rect 5123 3772 5124 3776
rect 5118 3771 5124 3772
rect 5342 3776 5348 3777
rect 5342 3772 5343 3776
rect 5347 3772 5348 3776
rect 5342 3771 5348 3772
rect 5542 3776 5548 3777
rect 5542 3772 5543 3776
rect 5547 3772 5548 3776
rect 5542 3771 5548 3772
rect 5662 3775 5668 3776
rect 5662 3771 5663 3775
rect 5667 3771 5668 3775
rect 3838 3770 3844 3771
rect 5662 3770 5668 3771
rect 1974 3752 1980 3753
rect 3798 3752 3804 3753
rect 1974 3748 1975 3752
rect 1979 3748 1980 3752
rect 1974 3747 1980 3748
rect 1994 3751 2000 3752
rect 1994 3747 1995 3751
rect 1999 3747 2000 3751
rect 1994 3746 2000 3747
rect 2130 3751 2136 3752
rect 2130 3747 2131 3751
rect 2135 3747 2136 3751
rect 2130 3746 2136 3747
rect 2282 3751 2288 3752
rect 2282 3747 2283 3751
rect 2287 3747 2288 3751
rect 2282 3746 2288 3747
rect 2442 3751 2448 3752
rect 2442 3747 2443 3751
rect 2447 3747 2448 3751
rect 2442 3746 2448 3747
rect 2602 3751 2608 3752
rect 2602 3747 2603 3751
rect 2607 3747 2608 3751
rect 2602 3746 2608 3747
rect 2762 3751 2768 3752
rect 2762 3747 2763 3751
rect 2767 3747 2768 3751
rect 2762 3746 2768 3747
rect 2922 3751 2928 3752
rect 2922 3747 2923 3751
rect 2927 3747 2928 3751
rect 2922 3746 2928 3747
rect 3082 3751 3088 3752
rect 3082 3747 3083 3751
rect 3087 3747 3088 3751
rect 3082 3746 3088 3747
rect 3242 3751 3248 3752
rect 3242 3747 3243 3751
rect 3247 3747 3248 3751
rect 3242 3746 3248 3747
rect 3410 3751 3416 3752
rect 3410 3747 3411 3751
rect 3415 3747 3416 3751
rect 3798 3748 3799 3752
rect 3803 3748 3804 3752
rect 3798 3747 3804 3748
rect 3410 3746 3416 3747
rect 2022 3736 2028 3737
rect 1974 3735 1980 3736
rect 1974 3731 1975 3735
rect 1979 3731 1980 3735
rect 2022 3732 2023 3736
rect 2027 3732 2028 3736
rect 2022 3731 2028 3732
rect 2158 3736 2164 3737
rect 2158 3732 2159 3736
rect 2163 3732 2164 3736
rect 2158 3731 2164 3732
rect 2310 3736 2316 3737
rect 2310 3732 2311 3736
rect 2315 3732 2316 3736
rect 2310 3731 2316 3732
rect 2470 3736 2476 3737
rect 2470 3732 2471 3736
rect 2475 3732 2476 3736
rect 2470 3731 2476 3732
rect 2630 3736 2636 3737
rect 2630 3732 2631 3736
rect 2635 3732 2636 3736
rect 2630 3731 2636 3732
rect 2790 3736 2796 3737
rect 2790 3732 2791 3736
rect 2795 3732 2796 3736
rect 2790 3731 2796 3732
rect 2950 3736 2956 3737
rect 2950 3732 2951 3736
rect 2955 3732 2956 3736
rect 2950 3731 2956 3732
rect 3110 3736 3116 3737
rect 3110 3732 3111 3736
rect 3115 3732 3116 3736
rect 3110 3731 3116 3732
rect 3270 3736 3276 3737
rect 3270 3732 3271 3736
rect 3275 3732 3276 3736
rect 3270 3731 3276 3732
rect 3438 3736 3444 3737
rect 3438 3732 3439 3736
rect 3443 3732 3444 3736
rect 3438 3731 3444 3732
rect 3798 3735 3804 3736
rect 3798 3731 3799 3735
rect 3803 3731 3804 3735
rect 1974 3730 1980 3731
rect 3798 3730 3804 3731
rect 3838 3693 3844 3694
rect 5662 3693 5668 3694
rect 3838 3689 3839 3693
rect 3843 3689 3844 3693
rect 3838 3688 3844 3689
rect 4270 3692 4276 3693
rect 4270 3688 4271 3692
rect 4275 3688 4276 3692
rect 4270 3687 4276 3688
rect 4470 3692 4476 3693
rect 4470 3688 4471 3692
rect 4475 3688 4476 3692
rect 4470 3687 4476 3688
rect 4694 3692 4700 3693
rect 4694 3688 4695 3692
rect 4699 3688 4700 3692
rect 4694 3687 4700 3688
rect 4934 3692 4940 3693
rect 4934 3688 4935 3692
rect 4939 3688 4940 3692
rect 4934 3687 4940 3688
rect 5190 3692 5196 3693
rect 5190 3688 5191 3692
rect 5195 3688 5196 3692
rect 5190 3687 5196 3688
rect 5446 3692 5452 3693
rect 5446 3688 5447 3692
rect 5451 3688 5452 3692
rect 5662 3689 5663 3693
rect 5667 3689 5668 3693
rect 5662 3688 5668 3689
rect 5446 3687 5452 3688
rect 4242 3677 4248 3678
rect 3838 3676 3844 3677
rect 3838 3672 3839 3676
rect 3843 3672 3844 3676
rect 4242 3673 4243 3677
rect 4247 3673 4248 3677
rect 4242 3672 4248 3673
rect 4442 3677 4448 3678
rect 4442 3673 4443 3677
rect 4447 3673 4448 3677
rect 4442 3672 4448 3673
rect 4666 3677 4672 3678
rect 4666 3673 4667 3677
rect 4671 3673 4672 3677
rect 4666 3672 4672 3673
rect 4906 3677 4912 3678
rect 4906 3673 4907 3677
rect 4911 3673 4912 3677
rect 4906 3672 4912 3673
rect 5162 3677 5168 3678
rect 5162 3673 5163 3677
rect 5167 3673 5168 3677
rect 5162 3672 5168 3673
rect 5418 3677 5424 3678
rect 5418 3673 5419 3677
rect 5423 3673 5424 3677
rect 5418 3672 5424 3673
rect 5662 3676 5668 3677
rect 5662 3672 5663 3676
rect 5667 3672 5668 3676
rect 3838 3671 3844 3672
rect 5662 3671 5668 3672
rect 1974 3669 1980 3670
rect 3798 3669 3804 3670
rect 1974 3665 1975 3669
rect 1979 3665 1980 3669
rect 1974 3664 1980 3665
rect 2046 3668 2052 3669
rect 2046 3664 2047 3668
rect 2051 3664 2052 3668
rect 2046 3663 2052 3664
rect 2222 3668 2228 3669
rect 2222 3664 2223 3668
rect 2227 3664 2228 3668
rect 2222 3663 2228 3664
rect 2406 3668 2412 3669
rect 2406 3664 2407 3668
rect 2411 3664 2412 3668
rect 2406 3663 2412 3664
rect 2590 3668 2596 3669
rect 2590 3664 2591 3668
rect 2595 3664 2596 3668
rect 2590 3663 2596 3664
rect 2782 3668 2788 3669
rect 2782 3664 2783 3668
rect 2787 3664 2788 3668
rect 2782 3663 2788 3664
rect 2966 3668 2972 3669
rect 2966 3664 2967 3668
rect 2971 3664 2972 3668
rect 2966 3663 2972 3664
rect 3150 3668 3156 3669
rect 3150 3664 3151 3668
rect 3155 3664 3156 3668
rect 3150 3663 3156 3664
rect 3334 3668 3340 3669
rect 3334 3664 3335 3668
rect 3339 3664 3340 3668
rect 3334 3663 3340 3664
rect 3518 3668 3524 3669
rect 3518 3664 3519 3668
rect 3523 3664 3524 3668
rect 3518 3663 3524 3664
rect 3678 3668 3684 3669
rect 3678 3664 3679 3668
rect 3683 3664 3684 3668
rect 3798 3665 3799 3669
rect 3803 3665 3804 3669
rect 3798 3664 3804 3665
rect 3678 3663 3684 3664
rect 2018 3653 2024 3654
rect 1974 3652 1980 3653
rect 1974 3648 1975 3652
rect 1979 3648 1980 3652
rect 2018 3649 2019 3653
rect 2023 3649 2024 3653
rect 2018 3648 2024 3649
rect 2194 3653 2200 3654
rect 2194 3649 2195 3653
rect 2199 3649 2200 3653
rect 2194 3648 2200 3649
rect 2378 3653 2384 3654
rect 2378 3649 2379 3653
rect 2383 3649 2384 3653
rect 2378 3648 2384 3649
rect 2562 3653 2568 3654
rect 2562 3649 2563 3653
rect 2567 3649 2568 3653
rect 2562 3648 2568 3649
rect 2754 3653 2760 3654
rect 2754 3649 2755 3653
rect 2759 3649 2760 3653
rect 2754 3648 2760 3649
rect 2938 3653 2944 3654
rect 2938 3649 2939 3653
rect 2943 3649 2944 3653
rect 2938 3648 2944 3649
rect 3122 3653 3128 3654
rect 3122 3649 3123 3653
rect 3127 3649 3128 3653
rect 3122 3648 3128 3649
rect 3306 3653 3312 3654
rect 3306 3649 3307 3653
rect 3311 3649 3312 3653
rect 3306 3648 3312 3649
rect 3490 3653 3496 3654
rect 3490 3649 3491 3653
rect 3495 3649 3496 3653
rect 3490 3648 3496 3649
rect 3650 3653 3656 3654
rect 3650 3649 3651 3653
rect 3655 3649 3656 3653
rect 3650 3648 3656 3649
rect 3798 3652 3804 3653
rect 3798 3648 3799 3652
rect 3803 3648 3804 3652
rect 1974 3647 1980 3648
rect 3798 3647 3804 3648
rect 110 3632 116 3633
rect 1934 3632 1940 3633
rect 110 3628 111 3632
rect 115 3628 116 3632
rect 110 3627 116 3628
rect 154 3631 160 3632
rect 154 3627 155 3631
rect 159 3627 160 3631
rect 154 3626 160 3627
rect 290 3631 296 3632
rect 290 3627 291 3631
rect 295 3627 296 3631
rect 290 3626 296 3627
rect 426 3631 432 3632
rect 426 3627 427 3631
rect 431 3627 432 3631
rect 426 3626 432 3627
rect 562 3631 568 3632
rect 562 3627 563 3631
rect 567 3627 568 3631
rect 562 3626 568 3627
rect 698 3631 704 3632
rect 698 3627 699 3631
rect 703 3627 704 3631
rect 698 3626 704 3627
rect 834 3631 840 3632
rect 834 3627 835 3631
rect 839 3627 840 3631
rect 834 3626 840 3627
rect 970 3631 976 3632
rect 970 3627 971 3631
rect 975 3627 976 3631
rect 970 3626 976 3627
rect 1106 3631 1112 3632
rect 1106 3627 1107 3631
rect 1111 3627 1112 3631
rect 1106 3626 1112 3627
rect 1242 3631 1248 3632
rect 1242 3627 1243 3631
rect 1247 3627 1248 3631
rect 1242 3626 1248 3627
rect 1378 3631 1384 3632
rect 1378 3627 1379 3631
rect 1383 3627 1384 3631
rect 1378 3626 1384 3627
rect 1514 3631 1520 3632
rect 1514 3627 1515 3631
rect 1519 3627 1520 3631
rect 1934 3628 1935 3632
rect 1939 3628 1940 3632
rect 1934 3627 1940 3628
rect 1514 3626 1520 3627
rect 182 3616 188 3617
rect 110 3615 116 3616
rect 110 3611 111 3615
rect 115 3611 116 3615
rect 182 3612 183 3616
rect 187 3612 188 3616
rect 182 3611 188 3612
rect 318 3616 324 3617
rect 318 3612 319 3616
rect 323 3612 324 3616
rect 318 3611 324 3612
rect 454 3616 460 3617
rect 454 3612 455 3616
rect 459 3612 460 3616
rect 454 3611 460 3612
rect 590 3616 596 3617
rect 590 3612 591 3616
rect 595 3612 596 3616
rect 590 3611 596 3612
rect 726 3616 732 3617
rect 726 3612 727 3616
rect 731 3612 732 3616
rect 726 3611 732 3612
rect 862 3616 868 3617
rect 862 3612 863 3616
rect 867 3612 868 3616
rect 862 3611 868 3612
rect 998 3616 1004 3617
rect 998 3612 999 3616
rect 1003 3612 1004 3616
rect 998 3611 1004 3612
rect 1134 3616 1140 3617
rect 1134 3612 1135 3616
rect 1139 3612 1140 3616
rect 1134 3611 1140 3612
rect 1270 3616 1276 3617
rect 1270 3612 1271 3616
rect 1275 3612 1276 3616
rect 1270 3611 1276 3612
rect 1406 3616 1412 3617
rect 1406 3612 1407 3616
rect 1411 3612 1412 3616
rect 1406 3611 1412 3612
rect 1542 3616 1548 3617
rect 1542 3612 1543 3616
rect 1547 3612 1548 3616
rect 1542 3611 1548 3612
rect 1934 3615 1940 3616
rect 1934 3611 1935 3615
rect 1939 3611 1940 3615
rect 110 3610 116 3611
rect 1934 3610 1940 3611
rect 3838 3540 3844 3541
rect 5662 3540 5668 3541
rect 3838 3536 3839 3540
rect 3843 3536 3844 3540
rect 3838 3535 3844 3536
rect 3858 3539 3864 3540
rect 3858 3535 3859 3539
rect 3863 3535 3864 3539
rect 3858 3534 3864 3535
rect 3994 3539 4000 3540
rect 3994 3535 3995 3539
rect 3999 3535 4000 3539
rect 3994 3534 4000 3535
rect 4130 3539 4136 3540
rect 4130 3535 4131 3539
rect 4135 3535 4136 3539
rect 4130 3534 4136 3535
rect 4266 3539 4272 3540
rect 4266 3535 4267 3539
rect 4271 3535 4272 3539
rect 4266 3534 4272 3535
rect 4402 3539 4408 3540
rect 4402 3535 4403 3539
rect 4407 3535 4408 3539
rect 4402 3534 4408 3535
rect 4538 3539 4544 3540
rect 4538 3535 4539 3539
rect 4543 3535 4544 3539
rect 4538 3534 4544 3535
rect 4674 3539 4680 3540
rect 4674 3535 4675 3539
rect 4679 3535 4680 3539
rect 4674 3534 4680 3535
rect 4810 3539 4816 3540
rect 4810 3535 4811 3539
rect 4815 3535 4816 3539
rect 4810 3534 4816 3535
rect 4946 3539 4952 3540
rect 4946 3535 4947 3539
rect 4951 3535 4952 3539
rect 5662 3536 5663 3540
rect 5667 3536 5668 3540
rect 5662 3535 5668 3536
rect 4946 3534 4952 3535
rect 3886 3524 3892 3525
rect 3838 3523 3844 3524
rect 3838 3519 3839 3523
rect 3843 3519 3844 3523
rect 3886 3520 3887 3524
rect 3891 3520 3892 3524
rect 3886 3519 3892 3520
rect 4022 3524 4028 3525
rect 4022 3520 4023 3524
rect 4027 3520 4028 3524
rect 4022 3519 4028 3520
rect 4158 3524 4164 3525
rect 4158 3520 4159 3524
rect 4163 3520 4164 3524
rect 4158 3519 4164 3520
rect 4294 3524 4300 3525
rect 4294 3520 4295 3524
rect 4299 3520 4300 3524
rect 4294 3519 4300 3520
rect 4430 3524 4436 3525
rect 4430 3520 4431 3524
rect 4435 3520 4436 3524
rect 4430 3519 4436 3520
rect 4566 3524 4572 3525
rect 4566 3520 4567 3524
rect 4571 3520 4572 3524
rect 4566 3519 4572 3520
rect 4702 3524 4708 3525
rect 4702 3520 4703 3524
rect 4707 3520 4708 3524
rect 4702 3519 4708 3520
rect 4838 3524 4844 3525
rect 4838 3520 4839 3524
rect 4843 3520 4844 3524
rect 4838 3519 4844 3520
rect 4974 3524 4980 3525
rect 4974 3520 4975 3524
rect 4979 3520 4980 3524
rect 4974 3519 4980 3520
rect 5662 3523 5668 3524
rect 5662 3519 5663 3523
rect 5667 3519 5668 3523
rect 3838 3518 3844 3519
rect 5662 3518 5668 3519
rect 1974 3508 1980 3509
rect 3798 3508 3804 3509
rect 1974 3504 1975 3508
rect 1979 3504 1980 3508
rect 1974 3503 1980 3504
rect 2306 3507 2312 3508
rect 2306 3503 2307 3507
rect 2311 3503 2312 3507
rect 2306 3502 2312 3503
rect 2442 3507 2448 3508
rect 2442 3503 2443 3507
rect 2447 3503 2448 3507
rect 2442 3502 2448 3503
rect 2578 3507 2584 3508
rect 2578 3503 2579 3507
rect 2583 3503 2584 3507
rect 2578 3502 2584 3503
rect 2714 3507 2720 3508
rect 2714 3503 2715 3507
rect 2719 3503 2720 3507
rect 3798 3504 3799 3508
rect 3803 3504 3804 3508
rect 3798 3503 3804 3504
rect 2714 3502 2720 3503
rect 2334 3492 2340 3493
rect 1974 3491 1980 3492
rect 1974 3487 1975 3491
rect 1979 3487 1980 3491
rect 2334 3488 2335 3492
rect 2339 3488 2340 3492
rect 2334 3487 2340 3488
rect 2470 3492 2476 3493
rect 2470 3488 2471 3492
rect 2475 3488 2476 3492
rect 2470 3487 2476 3488
rect 2606 3492 2612 3493
rect 2606 3488 2607 3492
rect 2611 3488 2612 3492
rect 2606 3487 2612 3488
rect 2742 3492 2748 3493
rect 2742 3488 2743 3492
rect 2747 3488 2748 3492
rect 2742 3487 2748 3488
rect 3798 3491 3804 3492
rect 3798 3487 3799 3491
rect 3803 3487 3804 3491
rect 1974 3486 1980 3487
rect 3798 3486 3804 3487
rect 3838 3465 3844 3466
rect 5662 3465 5668 3466
rect 3838 3461 3839 3465
rect 3843 3461 3844 3465
rect 3838 3460 3844 3461
rect 3886 3464 3892 3465
rect 3886 3460 3887 3464
rect 3891 3460 3892 3464
rect 3886 3459 3892 3460
rect 4022 3464 4028 3465
rect 4022 3460 4023 3464
rect 4027 3460 4028 3464
rect 4022 3459 4028 3460
rect 4158 3464 4164 3465
rect 4158 3460 4159 3464
rect 4163 3460 4164 3464
rect 4158 3459 4164 3460
rect 4294 3464 4300 3465
rect 4294 3460 4295 3464
rect 4299 3460 4300 3464
rect 4294 3459 4300 3460
rect 4430 3464 4436 3465
rect 4430 3460 4431 3464
rect 4435 3460 4436 3464
rect 4430 3459 4436 3460
rect 4566 3464 4572 3465
rect 4566 3460 4567 3464
rect 4571 3460 4572 3464
rect 4566 3459 4572 3460
rect 4702 3464 4708 3465
rect 4702 3460 4703 3464
rect 4707 3460 4708 3464
rect 4702 3459 4708 3460
rect 4838 3464 4844 3465
rect 4838 3460 4839 3464
rect 4843 3460 4844 3464
rect 4838 3459 4844 3460
rect 4974 3464 4980 3465
rect 4974 3460 4975 3464
rect 4979 3460 4980 3464
rect 4974 3459 4980 3460
rect 5110 3464 5116 3465
rect 5110 3460 5111 3464
rect 5115 3460 5116 3464
rect 5110 3459 5116 3460
rect 5246 3464 5252 3465
rect 5246 3460 5247 3464
rect 5251 3460 5252 3464
rect 5246 3459 5252 3460
rect 5382 3464 5388 3465
rect 5382 3460 5383 3464
rect 5387 3460 5388 3464
rect 5382 3459 5388 3460
rect 5518 3464 5524 3465
rect 5518 3460 5519 3464
rect 5523 3460 5524 3464
rect 5662 3461 5663 3465
rect 5667 3461 5668 3465
rect 5662 3460 5668 3461
rect 5518 3459 5524 3460
rect 3858 3449 3864 3450
rect 3838 3448 3844 3449
rect 3838 3444 3839 3448
rect 3843 3444 3844 3448
rect 3858 3445 3859 3449
rect 3863 3445 3864 3449
rect 3858 3444 3864 3445
rect 3994 3449 4000 3450
rect 3994 3445 3995 3449
rect 3999 3445 4000 3449
rect 3994 3444 4000 3445
rect 4130 3449 4136 3450
rect 4130 3445 4131 3449
rect 4135 3445 4136 3449
rect 4130 3444 4136 3445
rect 4266 3449 4272 3450
rect 4266 3445 4267 3449
rect 4271 3445 4272 3449
rect 4266 3444 4272 3445
rect 4402 3449 4408 3450
rect 4402 3445 4403 3449
rect 4407 3445 4408 3449
rect 4402 3444 4408 3445
rect 4538 3449 4544 3450
rect 4538 3445 4539 3449
rect 4543 3445 4544 3449
rect 4538 3444 4544 3445
rect 4674 3449 4680 3450
rect 4674 3445 4675 3449
rect 4679 3445 4680 3449
rect 4674 3444 4680 3445
rect 4810 3449 4816 3450
rect 4810 3445 4811 3449
rect 4815 3445 4816 3449
rect 4810 3444 4816 3445
rect 4946 3449 4952 3450
rect 4946 3445 4947 3449
rect 4951 3445 4952 3449
rect 4946 3444 4952 3445
rect 5082 3449 5088 3450
rect 5082 3445 5083 3449
rect 5087 3445 5088 3449
rect 5082 3444 5088 3445
rect 5218 3449 5224 3450
rect 5218 3445 5219 3449
rect 5223 3445 5224 3449
rect 5218 3444 5224 3445
rect 5354 3449 5360 3450
rect 5354 3445 5355 3449
rect 5359 3445 5360 3449
rect 5354 3444 5360 3445
rect 5490 3449 5496 3450
rect 5490 3445 5491 3449
rect 5495 3445 5496 3449
rect 5490 3444 5496 3445
rect 5662 3448 5668 3449
rect 5662 3444 5663 3448
rect 5667 3444 5668 3448
rect 3838 3443 3844 3444
rect 5662 3443 5668 3444
rect 1974 3397 1980 3398
rect 3798 3397 3804 3398
rect 1974 3393 1975 3397
rect 1979 3393 1980 3397
rect 1974 3392 1980 3393
rect 2166 3396 2172 3397
rect 2166 3392 2167 3396
rect 2171 3392 2172 3396
rect 2166 3391 2172 3392
rect 2302 3396 2308 3397
rect 2302 3392 2303 3396
rect 2307 3392 2308 3396
rect 2302 3391 2308 3392
rect 2438 3396 2444 3397
rect 2438 3392 2439 3396
rect 2443 3392 2444 3396
rect 2438 3391 2444 3392
rect 2574 3396 2580 3397
rect 2574 3392 2575 3396
rect 2579 3392 2580 3396
rect 2574 3391 2580 3392
rect 2710 3396 2716 3397
rect 2710 3392 2711 3396
rect 2715 3392 2716 3396
rect 2710 3391 2716 3392
rect 2846 3396 2852 3397
rect 2846 3392 2847 3396
rect 2851 3392 2852 3396
rect 2846 3391 2852 3392
rect 2982 3396 2988 3397
rect 2982 3392 2983 3396
rect 2987 3392 2988 3396
rect 3798 3393 3799 3397
rect 3803 3393 3804 3397
rect 3798 3392 3804 3393
rect 2982 3391 2988 3392
rect 2138 3381 2144 3382
rect 1974 3380 1980 3381
rect 1974 3376 1975 3380
rect 1979 3376 1980 3380
rect 2138 3377 2139 3381
rect 2143 3377 2144 3381
rect 2138 3376 2144 3377
rect 2274 3381 2280 3382
rect 2274 3377 2275 3381
rect 2279 3377 2280 3381
rect 2274 3376 2280 3377
rect 2410 3381 2416 3382
rect 2410 3377 2411 3381
rect 2415 3377 2416 3381
rect 2410 3376 2416 3377
rect 2546 3381 2552 3382
rect 2546 3377 2547 3381
rect 2551 3377 2552 3381
rect 2546 3376 2552 3377
rect 2682 3381 2688 3382
rect 2682 3377 2683 3381
rect 2687 3377 2688 3381
rect 2682 3376 2688 3377
rect 2818 3381 2824 3382
rect 2818 3377 2819 3381
rect 2823 3377 2824 3381
rect 2818 3376 2824 3377
rect 2954 3381 2960 3382
rect 2954 3377 2955 3381
rect 2959 3377 2960 3381
rect 2954 3376 2960 3377
rect 3798 3380 3804 3381
rect 3798 3376 3799 3380
rect 3803 3376 3804 3380
rect 1974 3375 1980 3376
rect 3798 3375 3804 3376
rect 3838 3308 3844 3309
rect 5662 3308 5668 3309
rect 3838 3304 3839 3308
rect 3843 3304 3844 3308
rect 3838 3303 3844 3304
rect 3858 3307 3864 3308
rect 3858 3303 3859 3307
rect 3863 3303 3864 3307
rect 3858 3302 3864 3303
rect 3994 3307 4000 3308
rect 3994 3303 3995 3307
rect 3999 3303 4000 3307
rect 3994 3302 4000 3303
rect 4154 3307 4160 3308
rect 4154 3303 4155 3307
rect 4159 3303 4160 3307
rect 4154 3302 4160 3303
rect 4314 3307 4320 3308
rect 4314 3303 4315 3307
rect 4319 3303 4320 3307
rect 4314 3302 4320 3303
rect 4466 3307 4472 3308
rect 4466 3303 4467 3307
rect 4471 3303 4472 3307
rect 4466 3302 4472 3303
rect 4626 3307 4632 3308
rect 4626 3303 4627 3307
rect 4631 3303 4632 3307
rect 4626 3302 4632 3303
rect 4786 3307 4792 3308
rect 4786 3303 4787 3307
rect 4791 3303 4792 3307
rect 4786 3302 4792 3303
rect 4946 3307 4952 3308
rect 4946 3303 4947 3307
rect 4951 3303 4952 3307
rect 5662 3304 5663 3308
rect 5667 3304 5668 3308
rect 5662 3303 5668 3304
rect 4946 3302 4952 3303
rect 3886 3292 3892 3293
rect 3838 3291 3844 3292
rect 3838 3287 3839 3291
rect 3843 3287 3844 3291
rect 3886 3288 3887 3292
rect 3891 3288 3892 3292
rect 3886 3287 3892 3288
rect 4022 3292 4028 3293
rect 4022 3288 4023 3292
rect 4027 3288 4028 3292
rect 4022 3287 4028 3288
rect 4182 3292 4188 3293
rect 4182 3288 4183 3292
rect 4187 3288 4188 3292
rect 4182 3287 4188 3288
rect 4342 3292 4348 3293
rect 4342 3288 4343 3292
rect 4347 3288 4348 3292
rect 4342 3287 4348 3288
rect 4494 3292 4500 3293
rect 4494 3288 4495 3292
rect 4499 3288 4500 3292
rect 4494 3287 4500 3288
rect 4654 3292 4660 3293
rect 4654 3288 4655 3292
rect 4659 3288 4660 3292
rect 4654 3287 4660 3288
rect 4814 3292 4820 3293
rect 4814 3288 4815 3292
rect 4819 3288 4820 3292
rect 4814 3287 4820 3288
rect 4974 3292 4980 3293
rect 4974 3288 4975 3292
rect 4979 3288 4980 3292
rect 4974 3287 4980 3288
rect 5662 3291 5668 3292
rect 5662 3287 5663 3291
rect 5667 3287 5668 3291
rect 3838 3286 3844 3287
rect 5662 3286 5668 3287
rect 110 3269 116 3270
rect 1934 3269 1940 3270
rect 110 3265 111 3269
rect 115 3265 116 3269
rect 110 3264 116 3265
rect 158 3268 164 3269
rect 158 3264 159 3268
rect 163 3264 164 3268
rect 158 3263 164 3264
rect 294 3268 300 3269
rect 294 3264 295 3268
rect 299 3264 300 3268
rect 294 3263 300 3264
rect 430 3268 436 3269
rect 430 3264 431 3268
rect 435 3264 436 3268
rect 430 3263 436 3264
rect 566 3268 572 3269
rect 566 3264 567 3268
rect 571 3264 572 3268
rect 566 3263 572 3264
rect 702 3268 708 3269
rect 702 3264 703 3268
rect 707 3264 708 3268
rect 702 3263 708 3264
rect 838 3268 844 3269
rect 838 3264 839 3268
rect 843 3264 844 3268
rect 838 3263 844 3264
rect 974 3268 980 3269
rect 974 3264 975 3268
rect 979 3264 980 3268
rect 974 3263 980 3264
rect 1110 3268 1116 3269
rect 1110 3264 1111 3268
rect 1115 3264 1116 3268
rect 1110 3263 1116 3264
rect 1246 3268 1252 3269
rect 1246 3264 1247 3268
rect 1251 3264 1252 3268
rect 1246 3263 1252 3264
rect 1382 3268 1388 3269
rect 1382 3264 1383 3268
rect 1387 3264 1388 3268
rect 1382 3263 1388 3264
rect 1518 3268 1524 3269
rect 1518 3264 1519 3268
rect 1523 3264 1524 3268
rect 1934 3265 1935 3269
rect 1939 3265 1940 3269
rect 1934 3264 1940 3265
rect 1518 3263 1524 3264
rect 130 3253 136 3254
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 130 3249 131 3253
rect 135 3249 136 3253
rect 130 3248 136 3249
rect 266 3253 272 3254
rect 266 3249 267 3253
rect 271 3249 272 3253
rect 266 3248 272 3249
rect 402 3253 408 3254
rect 402 3249 403 3253
rect 407 3249 408 3253
rect 402 3248 408 3249
rect 538 3253 544 3254
rect 538 3249 539 3253
rect 543 3249 544 3253
rect 538 3248 544 3249
rect 674 3253 680 3254
rect 674 3249 675 3253
rect 679 3249 680 3253
rect 674 3248 680 3249
rect 810 3253 816 3254
rect 810 3249 811 3253
rect 815 3249 816 3253
rect 810 3248 816 3249
rect 946 3253 952 3254
rect 946 3249 947 3253
rect 951 3249 952 3253
rect 946 3248 952 3249
rect 1082 3253 1088 3254
rect 1082 3249 1083 3253
rect 1087 3249 1088 3253
rect 1082 3248 1088 3249
rect 1218 3253 1224 3254
rect 1218 3249 1219 3253
rect 1223 3249 1224 3253
rect 1218 3248 1224 3249
rect 1354 3253 1360 3254
rect 1354 3249 1355 3253
rect 1359 3249 1360 3253
rect 1354 3248 1360 3249
rect 1490 3253 1496 3254
rect 1490 3249 1491 3253
rect 1495 3249 1496 3253
rect 1490 3248 1496 3249
rect 1934 3252 1940 3253
rect 1934 3248 1935 3252
rect 1939 3248 1940 3252
rect 110 3247 116 3248
rect 1934 3247 1940 3248
rect 1974 3248 1980 3249
rect 3798 3248 3804 3249
rect 1974 3244 1975 3248
rect 1979 3244 1980 3248
rect 1974 3243 1980 3244
rect 2058 3247 2064 3248
rect 2058 3243 2059 3247
rect 2063 3243 2064 3247
rect 2058 3242 2064 3243
rect 2202 3247 2208 3248
rect 2202 3243 2203 3247
rect 2207 3243 2208 3247
rect 2202 3242 2208 3243
rect 2362 3247 2368 3248
rect 2362 3243 2363 3247
rect 2367 3243 2368 3247
rect 2362 3242 2368 3243
rect 2538 3247 2544 3248
rect 2538 3243 2539 3247
rect 2543 3243 2544 3247
rect 2538 3242 2544 3243
rect 2738 3247 2744 3248
rect 2738 3243 2739 3247
rect 2743 3243 2744 3247
rect 2738 3242 2744 3243
rect 2954 3247 2960 3248
rect 2954 3243 2955 3247
rect 2959 3243 2960 3247
rect 2954 3242 2960 3243
rect 3186 3247 3192 3248
rect 3186 3243 3187 3247
rect 3191 3243 3192 3247
rect 3186 3242 3192 3243
rect 3426 3247 3432 3248
rect 3426 3243 3427 3247
rect 3431 3243 3432 3247
rect 3426 3242 3432 3243
rect 3650 3247 3656 3248
rect 3650 3243 3651 3247
rect 3655 3243 3656 3247
rect 3798 3244 3799 3248
rect 3803 3244 3804 3248
rect 3798 3243 3804 3244
rect 3650 3242 3656 3243
rect 2086 3232 2092 3233
rect 1974 3231 1980 3232
rect 1974 3227 1975 3231
rect 1979 3227 1980 3231
rect 2086 3228 2087 3232
rect 2091 3228 2092 3232
rect 2086 3227 2092 3228
rect 2230 3232 2236 3233
rect 2230 3228 2231 3232
rect 2235 3228 2236 3232
rect 2230 3227 2236 3228
rect 2390 3232 2396 3233
rect 2390 3228 2391 3232
rect 2395 3228 2396 3232
rect 2390 3227 2396 3228
rect 2566 3232 2572 3233
rect 2566 3228 2567 3232
rect 2571 3228 2572 3232
rect 2566 3227 2572 3228
rect 2766 3232 2772 3233
rect 2766 3228 2767 3232
rect 2771 3228 2772 3232
rect 2766 3227 2772 3228
rect 2982 3232 2988 3233
rect 2982 3228 2983 3232
rect 2987 3228 2988 3232
rect 2982 3227 2988 3228
rect 3214 3232 3220 3233
rect 3214 3228 3215 3232
rect 3219 3228 3220 3232
rect 3214 3227 3220 3228
rect 3454 3232 3460 3233
rect 3454 3228 3455 3232
rect 3459 3228 3460 3232
rect 3454 3227 3460 3228
rect 3678 3232 3684 3233
rect 3678 3228 3679 3232
rect 3683 3228 3684 3232
rect 3678 3227 3684 3228
rect 3798 3231 3804 3232
rect 3798 3227 3799 3231
rect 3803 3227 3804 3231
rect 1974 3226 1980 3227
rect 3798 3226 3804 3227
rect 3838 3221 3844 3222
rect 5662 3221 5668 3222
rect 3838 3217 3839 3221
rect 3843 3217 3844 3221
rect 3838 3216 3844 3217
rect 4806 3220 4812 3221
rect 4806 3216 4807 3220
rect 4811 3216 4812 3220
rect 4806 3215 4812 3216
rect 4942 3220 4948 3221
rect 4942 3216 4943 3220
rect 4947 3216 4948 3220
rect 4942 3215 4948 3216
rect 5078 3220 5084 3221
rect 5078 3216 5079 3220
rect 5083 3216 5084 3220
rect 5078 3215 5084 3216
rect 5214 3220 5220 3221
rect 5214 3216 5215 3220
rect 5219 3216 5220 3220
rect 5214 3215 5220 3216
rect 5350 3220 5356 3221
rect 5350 3216 5351 3220
rect 5355 3216 5356 3220
rect 5662 3217 5663 3221
rect 5667 3217 5668 3221
rect 5662 3216 5668 3217
rect 5350 3215 5356 3216
rect 4778 3205 4784 3206
rect 3838 3204 3844 3205
rect 3838 3200 3839 3204
rect 3843 3200 3844 3204
rect 4778 3201 4779 3205
rect 4783 3201 4784 3205
rect 4778 3200 4784 3201
rect 4914 3205 4920 3206
rect 4914 3201 4915 3205
rect 4919 3201 4920 3205
rect 4914 3200 4920 3201
rect 5050 3205 5056 3206
rect 5050 3201 5051 3205
rect 5055 3201 5056 3205
rect 5050 3200 5056 3201
rect 5186 3205 5192 3206
rect 5186 3201 5187 3205
rect 5191 3201 5192 3205
rect 5186 3200 5192 3201
rect 5322 3205 5328 3206
rect 5322 3201 5323 3205
rect 5327 3201 5328 3205
rect 5322 3200 5328 3201
rect 5662 3204 5668 3205
rect 5662 3200 5663 3204
rect 5667 3200 5668 3204
rect 3838 3199 3844 3200
rect 5662 3199 5668 3200
rect 1974 3169 1980 3170
rect 3798 3169 3804 3170
rect 1974 3165 1975 3169
rect 1979 3165 1980 3169
rect 1974 3164 1980 3165
rect 2022 3168 2028 3169
rect 2022 3164 2023 3168
rect 2027 3164 2028 3168
rect 2022 3163 2028 3164
rect 2158 3168 2164 3169
rect 2158 3164 2159 3168
rect 2163 3164 2164 3168
rect 2158 3163 2164 3164
rect 2302 3168 2308 3169
rect 2302 3164 2303 3168
rect 2307 3164 2308 3168
rect 2302 3163 2308 3164
rect 2454 3168 2460 3169
rect 2454 3164 2455 3168
rect 2459 3164 2460 3168
rect 2454 3163 2460 3164
rect 2614 3168 2620 3169
rect 2614 3164 2615 3168
rect 2619 3164 2620 3168
rect 2614 3163 2620 3164
rect 2782 3168 2788 3169
rect 2782 3164 2783 3168
rect 2787 3164 2788 3168
rect 2782 3163 2788 3164
rect 2950 3168 2956 3169
rect 2950 3164 2951 3168
rect 2955 3164 2956 3168
rect 2950 3163 2956 3164
rect 3126 3168 3132 3169
rect 3126 3164 3127 3168
rect 3131 3164 3132 3168
rect 3126 3163 3132 3164
rect 3310 3168 3316 3169
rect 3310 3164 3311 3168
rect 3315 3164 3316 3168
rect 3310 3163 3316 3164
rect 3502 3168 3508 3169
rect 3502 3164 3503 3168
rect 3507 3164 3508 3168
rect 3502 3163 3508 3164
rect 3678 3168 3684 3169
rect 3678 3164 3679 3168
rect 3683 3164 3684 3168
rect 3798 3165 3799 3169
rect 3803 3165 3804 3169
rect 3798 3164 3804 3165
rect 3678 3163 3684 3164
rect 1994 3153 2000 3154
rect 1974 3152 1980 3153
rect 1974 3148 1975 3152
rect 1979 3148 1980 3152
rect 1994 3149 1995 3153
rect 1999 3149 2000 3153
rect 1994 3148 2000 3149
rect 2130 3153 2136 3154
rect 2130 3149 2131 3153
rect 2135 3149 2136 3153
rect 2130 3148 2136 3149
rect 2274 3153 2280 3154
rect 2274 3149 2275 3153
rect 2279 3149 2280 3153
rect 2274 3148 2280 3149
rect 2426 3153 2432 3154
rect 2426 3149 2427 3153
rect 2431 3149 2432 3153
rect 2426 3148 2432 3149
rect 2586 3153 2592 3154
rect 2586 3149 2587 3153
rect 2591 3149 2592 3153
rect 2586 3148 2592 3149
rect 2754 3153 2760 3154
rect 2754 3149 2755 3153
rect 2759 3149 2760 3153
rect 2754 3148 2760 3149
rect 2922 3153 2928 3154
rect 2922 3149 2923 3153
rect 2927 3149 2928 3153
rect 2922 3148 2928 3149
rect 3098 3153 3104 3154
rect 3098 3149 3099 3153
rect 3103 3149 3104 3153
rect 3098 3148 3104 3149
rect 3282 3153 3288 3154
rect 3282 3149 3283 3153
rect 3287 3149 3288 3153
rect 3282 3148 3288 3149
rect 3474 3153 3480 3154
rect 3474 3149 3475 3153
rect 3479 3149 3480 3153
rect 3474 3148 3480 3149
rect 3650 3153 3656 3154
rect 3650 3149 3651 3153
rect 3655 3149 3656 3153
rect 3650 3148 3656 3149
rect 3798 3152 3804 3153
rect 3798 3148 3799 3152
rect 3803 3148 3804 3152
rect 1974 3147 1980 3148
rect 3798 3147 3804 3148
rect 110 3092 116 3093
rect 1934 3092 1940 3093
rect 110 3088 111 3092
rect 115 3088 116 3092
rect 110 3087 116 3088
rect 290 3091 296 3092
rect 290 3087 291 3091
rect 295 3087 296 3091
rect 290 3086 296 3087
rect 458 3091 464 3092
rect 458 3087 459 3091
rect 463 3087 464 3091
rect 458 3086 464 3087
rect 626 3091 632 3092
rect 626 3087 627 3091
rect 631 3087 632 3091
rect 626 3086 632 3087
rect 810 3091 816 3092
rect 810 3087 811 3091
rect 815 3087 816 3091
rect 810 3086 816 3087
rect 994 3091 1000 3092
rect 994 3087 995 3091
rect 999 3087 1000 3091
rect 994 3086 1000 3087
rect 1186 3091 1192 3092
rect 1186 3087 1187 3091
rect 1191 3087 1192 3091
rect 1186 3086 1192 3087
rect 1386 3091 1392 3092
rect 1386 3087 1387 3091
rect 1391 3087 1392 3091
rect 1386 3086 1392 3087
rect 1594 3091 1600 3092
rect 1594 3087 1595 3091
rect 1599 3087 1600 3091
rect 1594 3086 1600 3087
rect 1786 3091 1792 3092
rect 1786 3087 1787 3091
rect 1791 3087 1792 3091
rect 1934 3088 1935 3092
rect 1939 3088 1940 3092
rect 1934 3087 1940 3088
rect 1786 3086 1792 3087
rect 318 3076 324 3077
rect 110 3075 116 3076
rect 110 3071 111 3075
rect 115 3071 116 3075
rect 318 3072 319 3076
rect 323 3072 324 3076
rect 318 3071 324 3072
rect 486 3076 492 3077
rect 486 3072 487 3076
rect 491 3072 492 3076
rect 486 3071 492 3072
rect 654 3076 660 3077
rect 654 3072 655 3076
rect 659 3072 660 3076
rect 654 3071 660 3072
rect 838 3076 844 3077
rect 838 3072 839 3076
rect 843 3072 844 3076
rect 838 3071 844 3072
rect 1022 3076 1028 3077
rect 1022 3072 1023 3076
rect 1027 3072 1028 3076
rect 1022 3071 1028 3072
rect 1214 3076 1220 3077
rect 1214 3072 1215 3076
rect 1219 3072 1220 3076
rect 1214 3071 1220 3072
rect 1414 3076 1420 3077
rect 1414 3072 1415 3076
rect 1419 3072 1420 3076
rect 1414 3071 1420 3072
rect 1622 3076 1628 3077
rect 1622 3072 1623 3076
rect 1627 3072 1628 3076
rect 1622 3071 1628 3072
rect 1814 3076 1820 3077
rect 1814 3072 1815 3076
rect 1819 3072 1820 3076
rect 1814 3071 1820 3072
rect 1934 3075 1940 3076
rect 1934 3071 1935 3075
rect 1939 3071 1940 3075
rect 110 3070 116 3071
rect 1934 3070 1940 3071
rect 3838 3068 3844 3069
rect 5662 3068 5668 3069
rect 3838 3064 3839 3068
rect 3843 3064 3844 3068
rect 3838 3063 3844 3064
rect 4698 3067 4704 3068
rect 4698 3063 4699 3067
rect 4703 3063 4704 3067
rect 4698 3062 4704 3063
rect 4834 3067 4840 3068
rect 4834 3063 4835 3067
rect 4839 3063 4840 3067
rect 4834 3062 4840 3063
rect 4970 3067 4976 3068
rect 4970 3063 4971 3067
rect 4975 3063 4976 3067
rect 4970 3062 4976 3063
rect 5106 3067 5112 3068
rect 5106 3063 5107 3067
rect 5111 3063 5112 3067
rect 5106 3062 5112 3063
rect 5242 3067 5248 3068
rect 5242 3063 5243 3067
rect 5247 3063 5248 3067
rect 5242 3062 5248 3063
rect 5378 3067 5384 3068
rect 5378 3063 5379 3067
rect 5383 3063 5384 3067
rect 5378 3062 5384 3063
rect 5514 3067 5520 3068
rect 5514 3063 5515 3067
rect 5519 3063 5520 3067
rect 5662 3064 5663 3068
rect 5667 3064 5668 3068
rect 5662 3063 5668 3064
rect 5514 3062 5520 3063
rect 4726 3052 4732 3053
rect 3838 3051 3844 3052
rect 3838 3047 3839 3051
rect 3843 3047 3844 3051
rect 4726 3048 4727 3052
rect 4731 3048 4732 3052
rect 4726 3047 4732 3048
rect 4862 3052 4868 3053
rect 4862 3048 4863 3052
rect 4867 3048 4868 3052
rect 4862 3047 4868 3048
rect 4998 3052 5004 3053
rect 4998 3048 4999 3052
rect 5003 3048 5004 3052
rect 4998 3047 5004 3048
rect 5134 3052 5140 3053
rect 5134 3048 5135 3052
rect 5139 3048 5140 3052
rect 5134 3047 5140 3048
rect 5270 3052 5276 3053
rect 5270 3048 5271 3052
rect 5275 3048 5276 3052
rect 5270 3047 5276 3048
rect 5406 3052 5412 3053
rect 5406 3048 5407 3052
rect 5411 3048 5412 3052
rect 5406 3047 5412 3048
rect 5542 3052 5548 3053
rect 5542 3048 5543 3052
rect 5547 3048 5548 3052
rect 5542 3047 5548 3048
rect 5662 3051 5668 3052
rect 5662 3047 5663 3051
rect 5667 3047 5668 3051
rect 3838 3046 3844 3047
rect 5662 3046 5668 3047
rect 110 3017 116 3018
rect 1934 3017 1940 3018
rect 110 3013 111 3017
rect 115 3013 116 3017
rect 110 3012 116 3013
rect 326 3016 332 3017
rect 326 3012 327 3016
rect 331 3012 332 3016
rect 326 3011 332 3012
rect 486 3016 492 3017
rect 486 3012 487 3016
rect 491 3012 492 3016
rect 486 3011 492 3012
rect 646 3016 652 3017
rect 646 3012 647 3016
rect 651 3012 652 3016
rect 646 3011 652 3012
rect 806 3016 812 3017
rect 806 3012 807 3016
rect 811 3012 812 3016
rect 806 3011 812 3012
rect 958 3016 964 3017
rect 958 3012 959 3016
rect 963 3012 964 3016
rect 958 3011 964 3012
rect 1102 3016 1108 3017
rect 1102 3012 1103 3016
rect 1107 3012 1108 3016
rect 1102 3011 1108 3012
rect 1246 3016 1252 3017
rect 1246 3012 1247 3016
rect 1251 3012 1252 3016
rect 1246 3011 1252 3012
rect 1390 3016 1396 3017
rect 1390 3012 1391 3016
rect 1395 3012 1396 3016
rect 1390 3011 1396 3012
rect 1534 3016 1540 3017
rect 1534 3012 1535 3016
rect 1539 3012 1540 3016
rect 1534 3011 1540 3012
rect 1678 3016 1684 3017
rect 1678 3012 1679 3016
rect 1683 3012 1684 3016
rect 1678 3011 1684 3012
rect 1814 3016 1820 3017
rect 1814 3012 1815 3016
rect 1819 3012 1820 3016
rect 1934 3013 1935 3017
rect 1939 3013 1940 3017
rect 1934 3012 1940 3013
rect 1814 3011 1820 3012
rect 298 3001 304 3002
rect 110 3000 116 3001
rect 110 2996 111 3000
rect 115 2996 116 3000
rect 298 2997 299 3001
rect 303 2997 304 3001
rect 298 2996 304 2997
rect 458 3001 464 3002
rect 458 2997 459 3001
rect 463 2997 464 3001
rect 458 2996 464 2997
rect 618 3001 624 3002
rect 618 2997 619 3001
rect 623 2997 624 3001
rect 618 2996 624 2997
rect 778 3001 784 3002
rect 778 2997 779 3001
rect 783 2997 784 3001
rect 778 2996 784 2997
rect 930 3001 936 3002
rect 930 2997 931 3001
rect 935 2997 936 3001
rect 930 2996 936 2997
rect 1074 3001 1080 3002
rect 1074 2997 1075 3001
rect 1079 2997 1080 3001
rect 1074 2996 1080 2997
rect 1218 3001 1224 3002
rect 1218 2997 1219 3001
rect 1223 2997 1224 3001
rect 1218 2996 1224 2997
rect 1362 3001 1368 3002
rect 1362 2997 1363 3001
rect 1367 2997 1368 3001
rect 1362 2996 1368 2997
rect 1506 3001 1512 3002
rect 1506 2997 1507 3001
rect 1511 2997 1512 3001
rect 1506 2996 1512 2997
rect 1650 3001 1656 3002
rect 1650 2997 1651 3001
rect 1655 2997 1656 3001
rect 1650 2996 1656 2997
rect 1786 3001 1792 3002
rect 1786 2997 1787 3001
rect 1791 2997 1792 3001
rect 1786 2996 1792 2997
rect 1934 3000 1940 3001
rect 1934 2996 1935 3000
rect 1939 2996 1940 3000
rect 110 2995 116 2996
rect 1934 2995 1940 2996
rect 1974 3000 1980 3001
rect 3798 3000 3804 3001
rect 1974 2996 1975 3000
rect 1979 2996 1980 3000
rect 1974 2995 1980 2996
rect 2810 2999 2816 3000
rect 2810 2995 2811 2999
rect 2815 2995 2816 2999
rect 2810 2994 2816 2995
rect 3002 2999 3008 3000
rect 3002 2995 3003 2999
rect 3007 2995 3008 2999
rect 3002 2994 3008 2995
rect 3202 2999 3208 3000
rect 3202 2995 3203 2999
rect 3207 2995 3208 2999
rect 3202 2994 3208 2995
rect 3402 2999 3408 3000
rect 3402 2995 3403 2999
rect 3407 2995 3408 2999
rect 3402 2994 3408 2995
rect 3602 2999 3608 3000
rect 3602 2995 3603 2999
rect 3607 2995 3608 2999
rect 3798 2996 3799 3000
rect 3803 2996 3804 3000
rect 3798 2995 3804 2996
rect 3602 2994 3608 2995
rect 3838 2993 3844 2994
rect 5662 2993 5668 2994
rect 3838 2989 3839 2993
rect 3843 2989 3844 2993
rect 3838 2988 3844 2989
rect 4366 2992 4372 2993
rect 4366 2988 4367 2992
rect 4371 2988 4372 2992
rect 4366 2987 4372 2988
rect 4566 2992 4572 2993
rect 4566 2988 4567 2992
rect 4571 2988 4572 2992
rect 4566 2987 4572 2988
rect 4782 2992 4788 2993
rect 4782 2988 4783 2992
rect 4787 2988 4788 2992
rect 4782 2987 4788 2988
rect 5022 2992 5028 2993
rect 5022 2988 5023 2992
rect 5027 2988 5028 2992
rect 5022 2987 5028 2988
rect 5278 2992 5284 2993
rect 5278 2988 5279 2992
rect 5283 2988 5284 2992
rect 5278 2987 5284 2988
rect 5534 2992 5540 2993
rect 5534 2988 5535 2992
rect 5539 2988 5540 2992
rect 5662 2989 5663 2993
rect 5667 2989 5668 2993
rect 5662 2988 5668 2989
rect 5534 2987 5540 2988
rect 2838 2984 2844 2985
rect 1974 2983 1980 2984
rect 1974 2979 1975 2983
rect 1979 2979 1980 2983
rect 2838 2980 2839 2984
rect 2843 2980 2844 2984
rect 2838 2979 2844 2980
rect 3030 2984 3036 2985
rect 3030 2980 3031 2984
rect 3035 2980 3036 2984
rect 3030 2979 3036 2980
rect 3230 2984 3236 2985
rect 3230 2980 3231 2984
rect 3235 2980 3236 2984
rect 3230 2979 3236 2980
rect 3430 2984 3436 2985
rect 3430 2980 3431 2984
rect 3435 2980 3436 2984
rect 3430 2979 3436 2980
rect 3630 2984 3636 2985
rect 3630 2980 3631 2984
rect 3635 2980 3636 2984
rect 3630 2979 3636 2980
rect 3798 2983 3804 2984
rect 3798 2979 3799 2983
rect 3803 2979 3804 2983
rect 1974 2978 1980 2979
rect 3798 2978 3804 2979
rect 4338 2977 4344 2978
rect 3838 2976 3844 2977
rect 3838 2972 3839 2976
rect 3843 2972 3844 2976
rect 4338 2973 4339 2977
rect 4343 2973 4344 2977
rect 4338 2972 4344 2973
rect 4538 2977 4544 2978
rect 4538 2973 4539 2977
rect 4543 2973 4544 2977
rect 4538 2972 4544 2973
rect 4754 2977 4760 2978
rect 4754 2973 4755 2977
rect 4759 2973 4760 2977
rect 4754 2972 4760 2973
rect 4994 2977 5000 2978
rect 4994 2973 4995 2977
rect 4999 2973 5000 2977
rect 4994 2972 5000 2973
rect 5250 2977 5256 2978
rect 5250 2973 5251 2977
rect 5255 2973 5256 2977
rect 5250 2972 5256 2973
rect 5506 2977 5512 2978
rect 5506 2973 5507 2977
rect 5511 2973 5512 2977
rect 5506 2972 5512 2973
rect 5662 2976 5668 2977
rect 5662 2972 5663 2976
rect 5667 2972 5668 2976
rect 3838 2971 3844 2972
rect 5662 2971 5668 2972
rect 1974 2917 1980 2918
rect 3798 2917 3804 2918
rect 1974 2913 1975 2917
rect 1979 2913 1980 2917
rect 1974 2912 1980 2913
rect 2846 2916 2852 2917
rect 2846 2912 2847 2916
rect 2851 2912 2852 2916
rect 2846 2911 2852 2912
rect 2982 2916 2988 2917
rect 2982 2912 2983 2916
rect 2987 2912 2988 2916
rect 2982 2911 2988 2912
rect 3118 2916 3124 2917
rect 3118 2912 3119 2916
rect 3123 2912 3124 2916
rect 3118 2911 3124 2912
rect 3254 2916 3260 2917
rect 3254 2912 3255 2916
rect 3259 2912 3260 2916
rect 3254 2911 3260 2912
rect 3390 2916 3396 2917
rect 3390 2912 3391 2916
rect 3395 2912 3396 2916
rect 3390 2911 3396 2912
rect 3526 2916 3532 2917
rect 3526 2912 3527 2916
rect 3531 2912 3532 2916
rect 3526 2911 3532 2912
rect 3670 2916 3676 2917
rect 3670 2912 3671 2916
rect 3675 2912 3676 2916
rect 3798 2913 3799 2917
rect 3803 2913 3804 2917
rect 3798 2912 3804 2913
rect 3670 2911 3676 2912
rect 2818 2901 2824 2902
rect 1974 2900 1980 2901
rect 1974 2896 1975 2900
rect 1979 2896 1980 2900
rect 2818 2897 2819 2901
rect 2823 2897 2824 2901
rect 2818 2896 2824 2897
rect 2954 2901 2960 2902
rect 2954 2897 2955 2901
rect 2959 2897 2960 2901
rect 2954 2896 2960 2897
rect 3090 2901 3096 2902
rect 3090 2897 3091 2901
rect 3095 2897 3096 2901
rect 3090 2896 3096 2897
rect 3226 2901 3232 2902
rect 3226 2897 3227 2901
rect 3231 2897 3232 2901
rect 3226 2896 3232 2897
rect 3362 2901 3368 2902
rect 3362 2897 3363 2901
rect 3367 2897 3368 2901
rect 3362 2896 3368 2897
rect 3498 2901 3504 2902
rect 3498 2897 3499 2901
rect 3503 2897 3504 2901
rect 3498 2896 3504 2897
rect 3642 2901 3648 2902
rect 3642 2897 3643 2901
rect 3647 2897 3648 2901
rect 3642 2896 3648 2897
rect 3798 2900 3804 2901
rect 3798 2896 3799 2900
rect 3803 2896 3804 2900
rect 1974 2895 1980 2896
rect 3798 2895 3804 2896
rect 110 2868 116 2869
rect 1934 2868 1940 2869
rect 110 2864 111 2868
rect 115 2864 116 2868
rect 110 2863 116 2864
rect 154 2867 160 2868
rect 154 2863 155 2867
rect 159 2863 160 2867
rect 154 2862 160 2863
rect 378 2867 384 2868
rect 378 2863 379 2867
rect 383 2863 384 2867
rect 378 2862 384 2863
rect 594 2867 600 2868
rect 594 2863 595 2867
rect 599 2863 600 2867
rect 594 2862 600 2863
rect 810 2867 816 2868
rect 810 2863 811 2867
rect 815 2863 816 2867
rect 810 2862 816 2863
rect 1018 2867 1024 2868
rect 1018 2863 1019 2867
rect 1023 2863 1024 2867
rect 1018 2862 1024 2863
rect 1218 2867 1224 2868
rect 1218 2863 1219 2867
rect 1223 2863 1224 2867
rect 1218 2862 1224 2863
rect 1410 2867 1416 2868
rect 1410 2863 1411 2867
rect 1415 2863 1416 2867
rect 1410 2862 1416 2863
rect 1610 2867 1616 2868
rect 1610 2863 1611 2867
rect 1615 2863 1616 2867
rect 1610 2862 1616 2863
rect 1786 2867 1792 2868
rect 1786 2863 1787 2867
rect 1791 2863 1792 2867
rect 1934 2864 1935 2868
rect 1939 2864 1940 2868
rect 1934 2863 1940 2864
rect 1786 2862 1792 2863
rect 182 2852 188 2853
rect 110 2851 116 2852
rect 110 2847 111 2851
rect 115 2847 116 2851
rect 182 2848 183 2852
rect 187 2848 188 2852
rect 182 2847 188 2848
rect 406 2852 412 2853
rect 406 2848 407 2852
rect 411 2848 412 2852
rect 406 2847 412 2848
rect 622 2852 628 2853
rect 622 2848 623 2852
rect 627 2848 628 2852
rect 622 2847 628 2848
rect 838 2852 844 2853
rect 838 2848 839 2852
rect 843 2848 844 2852
rect 838 2847 844 2848
rect 1046 2852 1052 2853
rect 1046 2848 1047 2852
rect 1051 2848 1052 2852
rect 1046 2847 1052 2848
rect 1246 2852 1252 2853
rect 1246 2848 1247 2852
rect 1251 2848 1252 2852
rect 1246 2847 1252 2848
rect 1438 2852 1444 2853
rect 1438 2848 1439 2852
rect 1443 2848 1444 2852
rect 1438 2847 1444 2848
rect 1638 2852 1644 2853
rect 1638 2848 1639 2852
rect 1643 2848 1644 2852
rect 1638 2847 1644 2848
rect 1814 2852 1820 2853
rect 1814 2848 1815 2852
rect 1819 2848 1820 2852
rect 1814 2847 1820 2848
rect 1934 2851 1940 2852
rect 1934 2847 1935 2851
rect 1939 2847 1940 2851
rect 110 2846 116 2847
rect 1934 2846 1940 2847
rect 3838 2844 3844 2845
rect 5662 2844 5668 2845
rect 3838 2840 3839 2844
rect 3843 2840 3844 2844
rect 3838 2839 3844 2840
rect 4034 2843 4040 2844
rect 4034 2839 4035 2843
rect 4039 2839 4040 2843
rect 4034 2838 4040 2839
rect 4314 2843 4320 2844
rect 4314 2839 4315 2843
rect 4319 2839 4320 2843
rect 4314 2838 4320 2839
rect 4602 2843 4608 2844
rect 4602 2839 4603 2843
rect 4607 2839 4608 2843
rect 4602 2838 4608 2839
rect 4906 2843 4912 2844
rect 4906 2839 4907 2843
rect 4911 2839 4912 2843
rect 4906 2838 4912 2839
rect 5218 2843 5224 2844
rect 5218 2839 5219 2843
rect 5223 2839 5224 2843
rect 5218 2838 5224 2839
rect 5514 2843 5520 2844
rect 5514 2839 5515 2843
rect 5519 2839 5520 2843
rect 5662 2840 5663 2844
rect 5667 2840 5668 2844
rect 5662 2839 5668 2840
rect 5514 2838 5520 2839
rect 4062 2828 4068 2829
rect 3838 2827 3844 2828
rect 3838 2823 3839 2827
rect 3843 2823 3844 2827
rect 4062 2824 4063 2828
rect 4067 2824 4068 2828
rect 4062 2823 4068 2824
rect 4342 2828 4348 2829
rect 4342 2824 4343 2828
rect 4347 2824 4348 2828
rect 4342 2823 4348 2824
rect 4630 2828 4636 2829
rect 4630 2824 4631 2828
rect 4635 2824 4636 2828
rect 4630 2823 4636 2824
rect 4934 2828 4940 2829
rect 4934 2824 4935 2828
rect 4939 2824 4940 2828
rect 4934 2823 4940 2824
rect 5246 2828 5252 2829
rect 5246 2824 5247 2828
rect 5251 2824 5252 2828
rect 5246 2823 5252 2824
rect 5542 2828 5548 2829
rect 5542 2824 5543 2828
rect 5547 2824 5548 2828
rect 5542 2823 5548 2824
rect 5662 2827 5668 2828
rect 5662 2823 5663 2827
rect 5667 2823 5668 2827
rect 3838 2822 3844 2823
rect 5662 2822 5668 2823
rect 1974 2768 1980 2769
rect 3798 2768 3804 2769
rect 1974 2764 1975 2768
rect 1979 2764 1980 2768
rect 1974 2763 1980 2764
rect 2010 2767 2016 2768
rect 2010 2763 2011 2767
rect 2015 2763 2016 2767
rect 2010 2762 2016 2763
rect 2250 2767 2256 2768
rect 2250 2763 2251 2767
rect 2255 2763 2256 2767
rect 2250 2762 2256 2763
rect 2490 2767 2496 2768
rect 2490 2763 2491 2767
rect 2495 2763 2496 2767
rect 2490 2762 2496 2763
rect 2730 2767 2736 2768
rect 2730 2763 2731 2767
rect 2735 2763 2736 2767
rect 2730 2762 2736 2763
rect 2970 2767 2976 2768
rect 2970 2763 2971 2767
rect 2975 2763 2976 2767
rect 3798 2764 3799 2768
rect 3803 2764 3804 2768
rect 3798 2763 3804 2764
rect 2970 2762 2976 2763
rect 110 2761 116 2762
rect 1934 2761 1940 2762
rect 110 2757 111 2761
rect 115 2757 116 2761
rect 110 2756 116 2757
rect 286 2760 292 2761
rect 286 2756 287 2760
rect 291 2756 292 2760
rect 286 2755 292 2756
rect 422 2760 428 2761
rect 422 2756 423 2760
rect 427 2756 428 2760
rect 422 2755 428 2756
rect 558 2760 564 2761
rect 558 2756 559 2760
rect 563 2756 564 2760
rect 558 2755 564 2756
rect 694 2760 700 2761
rect 694 2756 695 2760
rect 699 2756 700 2760
rect 694 2755 700 2756
rect 830 2760 836 2761
rect 830 2756 831 2760
rect 835 2756 836 2760
rect 1934 2757 1935 2761
rect 1939 2757 1940 2761
rect 1934 2756 1940 2757
rect 3838 2761 3844 2762
rect 5662 2761 5668 2762
rect 3838 2757 3839 2761
rect 3843 2757 3844 2761
rect 3838 2756 3844 2757
rect 3966 2760 3972 2761
rect 3966 2756 3967 2760
rect 3971 2756 3972 2760
rect 830 2755 836 2756
rect 3966 2755 3972 2756
rect 4254 2760 4260 2761
rect 4254 2756 4255 2760
rect 4259 2756 4260 2760
rect 4254 2755 4260 2756
rect 4566 2760 4572 2761
rect 4566 2756 4567 2760
rect 4571 2756 4572 2760
rect 4566 2755 4572 2756
rect 4894 2760 4900 2761
rect 4894 2756 4895 2760
rect 4899 2756 4900 2760
rect 4894 2755 4900 2756
rect 5230 2760 5236 2761
rect 5230 2756 5231 2760
rect 5235 2756 5236 2760
rect 5230 2755 5236 2756
rect 5542 2760 5548 2761
rect 5542 2756 5543 2760
rect 5547 2756 5548 2760
rect 5662 2757 5663 2761
rect 5667 2757 5668 2761
rect 5662 2756 5668 2757
rect 5542 2755 5548 2756
rect 2038 2752 2044 2753
rect 1974 2751 1980 2752
rect 1974 2747 1975 2751
rect 1979 2747 1980 2751
rect 2038 2748 2039 2752
rect 2043 2748 2044 2752
rect 2038 2747 2044 2748
rect 2278 2752 2284 2753
rect 2278 2748 2279 2752
rect 2283 2748 2284 2752
rect 2278 2747 2284 2748
rect 2518 2752 2524 2753
rect 2518 2748 2519 2752
rect 2523 2748 2524 2752
rect 2518 2747 2524 2748
rect 2758 2752 2764 2753
rect 2758 2748 2759 2752
rect 2763 2748 2764 2752
rect 2758 2747 2764 2748
rect 2998 2752 3004 2753
rect 2998 2748 2999 2752
rect 3003 2748 3004 2752
rect 2998 2747 3004 2748
rect 3798 2751 3804 2752
rect 3798 2747 3799 2751
rect 3803 2747 3804 2751
rect 1974 2746 1980 2747
rect 3798 2746 3804 2747
rect 258 2745 264 2746
rect 110 2744 116 2745
rect 110 2740 111 2744
rect 115 2740 116 2744
rect 258 2741 259 2745
rect 263 2741 264 2745
rect 258 2740 264 2741
rect 394 2745 400 2746
rect 394 2741 395 2745
rect 399 2741 400 2745
rect 394 2740 400 2741
rect 530 2745 536 2746
rect 530 2741 531 2745
rect 535 2741 536 2745
rect 530 2740 536 2741
rect 666 2745 672 2746
rect 666 2741 667 2745
rect 671 2741 672 2745
rect 666 2740 672 2741
rect 802 2745 808 2746
rect 3938 2745 3944 2746
rect 802 2741 803 2745
rect 807 2741 808 2745
rect 802 2740 808 2741
rect 1934 2744 1940 2745
rect 1934 2740 1935 2744
rect 1939 2740 1940 2744
rect 110 2739 116 2740
rect 1934 2739 1940 2740
rect 3838 2744 3844 2745
rect 3838 2740 3839 2744
rect 3843 2740 3844 2744
rect 3938 2741 3939 2745
rect 3943 2741 3944 2745
rect 3938 2740 3944 2741
rect 4226 2745 4232 2746
rect 4226 2741 4227 2745
rect 4231 2741 4232 2745
rect 4226 2740 4232 2741
rect 4538 2745 4544 2746
rect 4538 2741 4539 2745
rect 4543 2741 4544 2745
rect 4538 2740 4544 2741
rect 4866 2745 4872 2746
rect 4866 2741 4867 2745
rect 4871 2741 4872 2745
rect 4866 2740 4872 2741
rect 5202 2745 5208 2746
rect 5202 2741 5203 2745
rect 5207 2741 5208 2745
rect 5202 2740 5208 2741
rect 5514 2745 5520 2746
rect 5514 2741 5515 2745
rect 5519 2741 5520 2745
rect 5514 2740 5520 2741
rect 5662 2744 5668 2745
rect 5662 2740 5663 2744
rect 5667 2740 5668 2744
rect 3838 2739 3844 2740
rect 5662 2739 5668 2740
rect 1974 2693 1980 2694
rect 3798 2693 3804 2694
rect 1974 2689 1975 2693
rect 1979 2689 1980 2693
rect 1974 2688 1980 2689
rect 2022 2692 2028 2693
rect 2022 2688 2023 2692
rect 2027 2688 2028 2692
rect 2022 2687 2028 2688
rect 2158 2692 2164 2693
rect 2158 2688 2159 2692
rect 2163 2688 2164 2692
rect 2158 2687 2164 2688
rect 2294 2692 2300 2693
rect 2294 2688 2295 2692
rect 2299 2688 2300 2692
rect 2294 2687 2300 2688
rect 2430 2692 2436 2693
rect 2430 2688 2431 2692
rect 2435 2688 2436 2692
rect 2430 2687 2436 2688
rect 2566 2692 2572 2693
rect 2566 2688 2567 2692
rect 2571 2688 2572 2692
rect 2566 2687 2572 2688
rect 2702 2692 2708 2693
rect 2702 2688 2703 2692
rect 2707 2688 2708 2692
rect 2702 2687 2708 2688
rect 2838 2692 2844 2693
rect 2838 2688 2839 2692
rect 2843 2688 2844 2692
rect 2838 2687 2844 2688
rect 2974 2692 2980 2693
rect 2974 2688 2975 2692
rect 2979 2688 2980 2692
rect 2974 2687 2980 2688
rect 3110 2692 3116 2693
rect 3110 2688 3111 2692
rect 3115 2688 3116 2692
rect 3110 2687 3116 2688
rect 3246 2692 3252 2693
rect 3246 2688 3247 2692
rect 3251 2688 3252 2692
rect 3246 2687 3252 2688
rect 3382 2692 3388 2693
rect 3382 2688 3383 2692
rect 3387 2688 3388 2692
rect 3798 2689 3799 2693
rect 3803 2689 3804 2693
rect 3798 2688 3804 2689
rect 3382 2687 3388 2688
rect 1994 2677 2000 2678
rect 1974 2676 1980 2677
rect 1974 2672 1975 2676
rect 1979 2672 1980 2676
rect 1994 2673 1995 2677
rect 1999 2673 2000 2677
rect 1994 2672 2000 2673
rect 2130 2677 2136 2678
rect 2130 2673 2131 2677
rect 2135 2673 2136 2677
rect 2130 2672 2136 2673
rect 2266 2677 2272 2678
rect 2266 2673 2267 2677
rect 2271 2673 2272 2677
rect 2266 2672 2272 2673
rect 2402 2677 2408 2678
rect 2402 2673 2403 2677
rect 2407 2673 2408 2677
rect 2402 2672 2408 2673
rect 2538 2677 2544 2678
rect 2538 2673 2539 2677
rect 2543 2673 2544 2677
rect 2538 2672 2544 2673
rect 2674 2677 2680 2678
rect 2674 2673 2675 2677
rect 2679 2673 2680 2677
rect 2674 2672 2680 2673
rect 2810 2677 2816 2678
rect 2810 2673 2811 2677
rect 2815 2673 2816 2677
rect 2810 2672 2816 2673
rect 2946 2677 2952 2678
rect 2946 2673 2947 2677
rect 2951 2673 2952 2677
rect 2946 2672 2952 2673
rect 3082 2677 3088 2678
rect 3082 2673 3083 2677
rect 3087 2673 3088 2677
rect 3082 2672 3088 2673
rect 3218 2677 3224 2678
rect 3218 2673 3219 2677
rect 3223 2673 3224 2677
rect 3218 2672 3224 2673
rect 3354 2677 3360 2678
rect 3354 2673 3355 2677
rect 3359 2673 3360 2677
rect 3354 2672 3360 2673
rect 3798 2676 3804 2677
rect 3798 2672 3799 2676
rect 3803 2672 3804 2676
rect 1974 2671 1980 2672
rect 3798 2671 3804 2672
rect 3838 2608 3844 2609
rect 5662 2608 5668 2609
rect 3838 2604 3839 2608
rect 3843 2604 3844 2608
rect 3838 2603 3844 2604
rect 4026 2607 4032 2608
rect 4026 2603 4027 2607
rect 4031 2603 4032 2607
rect 4026 2602 4032 2603
rect 4274 2607 4280 2608
rect 4274 2603 4275 2607
rect 4279 2603 4280 2607
rect 4274 2602 4280 2603
rect 4554 2607 4560 2608
rect 4554 2603 4555 2607
rect 4559 2603 4560 2607
rect 4554 2602 4560 2603
rect 4866 2607 4872 2608
rect 4866 2603 4867 2607
rect 4871 2603 4872 2607
rect 4866 2602 4872 2603
rect 5202 2607 5208 2608
rect 5202 2603 5203 2607
rect 5207 2603 5208 2607
rect 5202 2602 5208 2603
rect 5514 2607 5520 2608
rect 5514 2603 5515 2607
rect 5519 2603 5520 2607
rect 5662 2604 5663 2608
rect 5667 2604 5668 2608
rect 5662 2603 5668 2604
rect 5514 2602 5520 2603
rect 110 2592 116 2593
rect 1934 2592 1940 2593
rect 4054 2592 4060 2593
rect 110 2588 111 2592
rect 115 2588 116 2592
rect 110 2587 116 2588
rect 538 2591 544 2592
rect 538 2587 539 2591
rect 543 2587 544 2591
rect 538 2586 544 2587
rect 698 2591 704 2592
rect 698 2587 699 2591
rect 703 2587 704 2591
rect 698 2586 704 2587
rect 882 2591 888 2592
rect 882 2587 883 2591
rect 887 2587 888 2591
rect 882 2586 888 2587
rect 1090 2591 1096 2592
rect 1090 2587 1091 2591
rect 1095 2587 1096 2591
rect 1090 2586 1096 2587
rect 1322 2591 1328 2592
rect 1322 2587 1323 2591
rect 1327 2587 1328 2591
rect 1322 2586 1328 2587
rect 1562 2591 1568 2592
rect 1562 2587 1563 2591
rect 1567 2587 1568 2591
rect 1562 2586 1568 2587
rect 1786 2591 1792 2592
rect 1786 2587 1787 2591
rect 1791 2587 1792 2591
rect 1934 2588 1935 2592
rect 1939 2588 1940 2592
rect 1934 2587 1940 2588
rect 3838 2591 3844 2592
rect 3838 2587 3839 2591
rect 3843 2587 3844 2591
rect 4054 2588 4055 2592
rect 4059 2588 4060 2592
rect 4054 2587 4060 2588
rect 4302 2592 4308 2593
rect 4302 2588 4303 2592
rect 4307 2588 4308 2592
rect 4302 2587 4308 2588
rect 4582 2592 4588 2593
rect 4582 2588 4583 2592
rect 4587 2588 4588 2592
rect 4582 2587 4588 2588
rect 4894 2592 4900 2593
rect 4894 2588 4895 2592
rect 4899 2588 4900 2592
rect 4894 2587 4900 2588
rect 5230 2592 5236 2593
rect 5230 2588 5231 2592
rect 5235 2588 5236 2592
rect 5230 2587 5236 2588
rect 5542 2592 5548 2593
rect 5542 2588 5543 2592
rect 5547 2588 5548 2592
rect 5542 2587 5548 2588
rect 5662 2591 5668 2592
rect 5662 2587 5663 2591
rect 5667 2587 5668 2591
rect 1786 2586 1792 2587
rect 3838 2586 3844 2587
rect 5662 2586 5668 2587
rect 566 2576 572 2577
rect 110 2575 116 2576
rect 110 2571 111 2575
rect 115 2571 116 2575
rect 566 2572 567 2576
rect 571 2572 572 2576
rect 566 2571 572 2572
rect 726 2576 732 2577
rect 726 2572 727 2576
rect 731 2572 732 2576
rect 726 2571 732 2572
rect 910 2576 916 2577
rect 910 2572 911 2576
rect 915 2572 916 2576
rect 910 2571 916 2572
rect 1118 2576 1124 2577
rect 1118 2572 1119 2576
rect 1123 2572 1124 2576
rect 1118 2571 1124 2572
rect 1350 2576 1356 2577
rect 1350 2572 1351 2576
rect 1355 2572 1356 2576
rect 1350 2571 1356 2572
rect 1590 2576 1596 2577
rect 1590 2572 1591 2576
rect 1595 2572 1596 2576
rect 1590 2571 1596 2572
rect 1814 2576 1820 2577
rect 1814 2572 1815 2576
rect 1819 2572 1820 2576
rect 1814 2571 1820 2572
rect 1934 2575 1940 2576
rect 1934 2571 1935 2575
rect 1939 2571 1940 2575
rect 110 2570 116 2571
rect 1934 2570 1940 2571
rect 1974 2544 1980 2545
rect 3798 2544 3804 2545
rect 1974 2540 1975 2544
rect 1979 2540 1980 2544
rect 1974 2539 1980 2540
rect 1994 2543 2000 2544
rect 1994 2539 1995 2543
rect 1999 2539 2000 2543
rect 1994 2538 2000 2539
rect 2202 2543 2208 2544
rect 2202 2539 2203 2543
rect 2207 2539 2208 2543
rect 2202 2538 2208 2539
rect 2418 2543 2424 2544
rect 2418 2539 2419 2543
rect 2423 2539 2424 2543
rect 2418 2538 2424 2539
rect 2626 2543 2632 2544
rect 2626 2539 2627 2543
rect 2631 2539 2632 2543
rect 2626 2538 2632 2539
rect 2826 2543 2832 2544
rect 2826 2539 2827 2543
rect 2831 2539 2832 2543
rect 2826 2538 2832 2539
rect 3018 2543 3024 2544
rect 3018 2539 3019 2543
rect 3023 2539 3024 2543
rect 3018 2538 3024 2539
rect 3210 2543 3216 2544
rect 3210 2539 3211 2543
rect 3215 2539 3216 2543
rect 3210 2538 3216 2539
rect 3402 2543 3408 2544
rect 3402 2539 3403 2543
rect 3407 2539 3408 2543
rect 3798 2540 3799 2544
rect 3803 2540 3804 2544
rect 3798 2539 3804 2540
rect 3402 2538 3408 2539
rect 3838 2529 3844 2530
rect 5662 2529 5668 2530
rect 2022 2528 2028 2529
rect 1974 2527 1980 2528
rect 1974 2523 1975 2527
rect 1979 2523 1980 2527
rect 2022 2524 2023 2528
rect 2027 2524 2028 2528
rect 2022 2523 2028 2524
rect 2230 2528 2236 2529
rect 2230 2524 2231 2528
rect 2235 2524 2236 2528
rect 2230 2523 2236 2524
rect 2446 2528 2452 2529
rect 2446 2524 2447 2528
rect 2451 2524 2452 2528
rect 2446 2523 2452 2524
rect 2654 2528 2660 2529
rect 2654 2524 2655 2528
rect 2659 2524 2660 2528
rect 2654 2523 2660 2524
rect 2854 2528 2860 2529
rect 2854 2524 2855 2528
rect 2859 2524 2860 2528
rect 2854 2523 2860 2524
rect 3046 2528 3052 2529
rect 3046 2524 3047 2528
rect 3051 2524 3052 2528
rect 3046 2523 3052 2524
rect 3238 2528 3244 2529
rect 3238 2524 3239 2528
rect 3243 2524 3244 2528
rect 3238 2523 3244 2524
rect 3430 2528 3436 2529
rect 3430 2524 3431 2528
rect 3435 2524 3436 2528
rect 3430 2523 3436 2524
rect 3798 2527 3804 2528
rect 3798 2523 3799 2527
rect 3803 2523 3804 2527
rect 3838 2525 3839 2529
rect 3843 2525 3844 2529
rect 3838 2524 3844 2525
rect 4334 2528 4340 2529
rect 4334 2524 4335 2528
rect 4339 2524 4340 2528
rect 4334 2523 4340 2524
rect 4558 2528 4564 2529
rect 4558 2524 4559 2528
rect 4563 2524 4564 2528
rect 4558 2523 4564 2524
rect 4798 2528 4804 2529
rect 4798 2524 4799 2528
rect 4803 2524 4804 2528
rect 4798 2523 4804 2524
rect 5046 2528 5052 2529
rect 5046 2524 5047 2528
rect 5051 2524 5052 2528
rect 5046 2523 5052 2524
rect 5302 2528 5308 2529
rect 5302 2524 5303 2528
rect 5307 2524 5308 2528
rect 5302 2523 5308 2524
rect 5542 2528 5548 2529
rect 5542 2524 5543 2528
rect 5547 2524 5548 2528
rect 5662 2525 5663 2529
rect 5667 2525 5668 2529
rect 5662 2524 5668 2525
rect 5542 2523 5548 2524
rect 1974 2522 1980 2523
rect 3798 2522 3804 2523
rect 4306 2513 4312 2514
rect 3838 2512 3844 2513
rect 3838 2508 3839 2512
rect 3843 2508 3844 2512
rect 4306 2509 4307 2513
rect 4311 2509 4312 2513
rect 4306 2508 4312 2509
rect 4530 2513 4536 2514
rect 4530 2509 4531 2513
rect 4535 2509 4536 2513
rect 4530 2508 4536 2509
rect 4770 2513 4776 2514
rect 4770 2509 4771 2513
rect 4775 2509 4776 2513
rect 4770 2508 4776 2509
rect 5018 2513 5024 2514
rect 5018 2509 5019 2513
rect 5023 2509 5024 2513
rect 5018 2508 5024 2509
rect 5274 2513 5280 2514
rect 5274 2509 5275 2513
rect 5279 2509 5280 2513
rect 5274 2508 5280 2509
rect 5514 2513 5520 2514
rect 5514 2509 5515 2513
rect 5519 2509 5520 2513
rect 5514 2508 5520 2509
rect 5662 2512 5668 2513
rect 5662 2508 5663 2512
rect 5667 2508 5668 2512
rect 3838 2507 3844 2508
rect 5662 2507 5668 2508
rect 110 2505 116 2506
rect 1934 2505 1940 2506
rect 110 2501 111 2505
rect 115 2501 116 2505
rect 110 2500 116 2501
rect 694 2504 700 2505
rect 694 2500 695 2504
rect 699 2500 700 2504
rect 694 2499 700 2500
rect 846 2504 852 2505
rect 846 2500 847 2504
rect 851 2500 852 2504
rect 846 2499 852 2500
rect 998 2504 1004 2505
rect 998 2500 999 2504
rect 1003 2500 1004 2504
rect 998 2499 1004 2500
rect 1158 2504 1164 2505
rect 1158 2500 1159 2504
rect 1163 2500 1164 2504
rect 1158 2499 1164 2500
rect 1326 2504 1332 2505
rect 1326 2500 1327 2504
rect 1331 2500 1332 2504
rect 1326 2499 1332 2500
rect 1494 2504 1500 2505
rect 1494 2500 1495 2504
rect 1499 2500 1500 2504
rect 1494 2499 1500 2500
rect 1662 2504 1668 2505
rect 1662 2500 1663 2504
rect 1667 2500 1668 2504
rect 1662 2499 1668 2500
rect 1814 2504 1820 2505
rect 1814 2500 1815 2504
rect 1819 2500 1820 2504
rect 1934 2501 1935 2505
rect 1939 2501 1940 2505
rect 1934 2500 1940 2501
rect 1814 2499 1820 2500
rect 666 2489 672 2490
rect 110 2488 116 2489
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 666 2485 667 2489
rect 671 2485 672 2489
rect 666 2484 672 2485
rect 818 2489 824 2490
rect 818 2485 819 2489
rect 823 2485 824 2489
rect 818 2484 824 2485
rect 970 2489 976 2490
rect 970 2485 971 2489
rect 975 2485 976 2489
rect 970 2484 976 2485
rect 1130 2489 1136 2490
rect 1130 2485 1131 2489
rect 1135 2485 1136 2489
rect 1130 2484 1136 2485
rect 1298 2489 1304 2490
rect 1298 2485 1299 2489
rect 1303 2485 1304 2489
rect 1298 2484 1304 2485
rect 1466 2489 1472 2490
rect 1466 2485 1467 2489
rect 1471 2485 1472 2489
rect 1466 2484 1472 2485
rect 1634 2489 1640 2490
rect 1634 2485 1635 2489
rect 1639 2485 1640 2489
rect 1634 2484 1640 2485
rect 1786 2489 1792 2490
rect 1786 2485 1787 2489
rect 1791 2485 1792 2489
rect 1786 2484 1792 2485
rect 1934 2488 1940 2489
rect 1934 2484 1935 2488
rect 1939 2484 1940 2488
rect 110 2483 116 2484
rect 1934 2483 1940 2484
rect 1974 2461 1980 2462
rect 3798 2461 3804 2462
rect 1974 2457 1975 2461
rect 1979 2457 1980 2461
rect 1974 2456 1980 2457
rect 2318 2460 2324 2461
rect 2318 2456 2319 2460
rect 2323 2456 2324 2460
rect 2318 2455 2324 2456
rect 2566 2460 2572 2461
rect 2566 2456 2567 2460
rect 2571 2456 2572 2460
rect 2566 2455 2572 2456
rect 2798 2460 2804 2461
rect 2798 2456 2799 2460
rect 2803 2456 2804 2460
rect 2798 2455 2804 2456
rect 3022 2460 3028 2461
rect 3022 2456 3023 2460
rect 3027 2456 3028 2460
rect 3022 2455 3028 2456
rect 3238 2460 3244 2461
rect 3238 2456 3239 2460
rect 3243 2456 3244 2460
rect 3238 2455 3244 2456
rect 3454 2460 3460 2461
rect 3454 2456 3455 2460
rect 3459 2456 3460 2460
rect 3454 2455 3460 2456
rect 3670 2460 3676 2461
rect 3670 2456 3671 2460
rect 3675 2456 3676 2460
rect 3798 2457 3799 2461
rect 3803 2457 3804 2461
rect 3798 2456 3804 2457
rect 3670 2455 3676 2456
rect 2290 2445 2296 2446
rect 1974 2444 1980 2445
rect 1974 2440 1975 2444
rect 1979 2440 1980 2444
rect 2290 2441 2291 2445
rect 2295 2441 2296 2445
rect 2290 2440 2296 2441
rect 2538 2445 2544 2446
rect 2538 2441 2539 2445
rect 2543 2441 2544 2445
rect 2538 2440 2544 2441
rect 2770 2445 2776 2446
rect 2770 2441 2771 2445
rect 2775 2441 2776 2445
rect 2770 2440 2776 2441
rect 2994 2445 3000 2446
rect 2994 2441 2995 2445
rect 2999 2441 3000 2445
rect 2994 2440 3000 2441
rect 3210 2445 3216 2446
rect 3210 2441 3211 2445
rect 3215 2441 3216 2445
rect 3210 2440 3216 2441
rect 3426 2445 3432 2446
rect 3426 2441 3427 2445
rect 3431 2441 3432 2445
rect 3426 2440 3432 2441
rect 3642 2445 3648 2446
rect 3642 2441 3643 2445
rect 3647 2441 3648 2445
rect 3642 2440 3648 2441
rect 3798 2444 3804 2445
rect 3798 2440 3799 2444
rect 3803 2440 3804 2444
rect 1974 2439 1980 2440
rect 3798 2439 3804 2440
rect 3838 2364 3844 2365
rect 5662 2364 5668 2365
rect 3838 2360 3839 2364
rect 3843 2360 3844 2364
rect 3838 2359 3844 2360
rect 4490 2363 4496 2364
rect 4490 2359 4491 2363
rect 4495 2359 4496 2363
rect 4490 2358 4496 2359
rect 4634 2363 4640 2364
rect 4634 2359 4635 2363
rect 4639 2359 4640 2363
rect 4634 2358 4640 2359
rect 4794 2363 4800 2364
rect 4794 2359 4795 2363
rect 4799 2359 4800 2363
rect 4794 2358 4800 2359
rect 4962 2363 4968 2364
rect 4962 2359 4963 2363
rect 4967 2359 4968 2363
rect 4962 2358 4968 2359
rect 5138 2363 5144 2364
rect 5138 2359 5139 2363
rect 5143 2359 5144 2363
rect 5138 2358 5144 2359
rect 5322 2363 5328 2364
rect 5322 2359 5323 2363
rect 5327 2359 5328 2363
rect 5322 2358 5328 2359
rect 5514 2363 5520 2364
rect 5514 2359 5515 2363
rect 5519 2359 5520 2363
rect 5662 2360 5663 2364
rect 5667 2360 5668 2364
rect 5662 2359 5668 2360
rect 5514 2358 5520 2359
rect 110 2348 116 2349
rect 1934 2348 1940 2349
rect 4518 2348 4524 2349
rect 110 2344 111 2348
rect 115 2344 116 2348
rect 110 2343 116 2344
rect 354 2347 360 2348
rect 354 2343 355 2347
rect 359 2343 360 2347
rect 354 2342 360 2343
rect 506 2347 512 2348
rect 506 2343 507 2347
rect 511 2343 512 2347
rect 506 2342 512 2343
rect 674 2347 680 2348
rect 674 2343 675 2347
rect 679 2343 680 2347
rect 674 2342 680 2343
rect 858 2347 864 2348
rect 858 2343 859 2347
rect 863 2343 864 2347
rect 858 2342 864 2343
rect 1058 2347 1064 2348
rect 1058 2343 1059 2347
rect 1063 2343 1064 2347
rect 1058 2342 1064 2343
rect 1266 2347 1272 2348
rect 1266 2343 1267 2347
rect 1271 2343 1272 2347
rect 1266 2342 1272 2343
rect 1482 2347 1488 2348
rect 1482 2343 1483 2347
rect 1487 2343 1488 2347
rect 1482 2342 1488 2343
rect 1698 2347 1704 2348
rect 1698 2343 1699 2347
rect 1703 2343 1704 2347
rect 1934 2344 1935 2348
rect 1939 2344 1940 2348
rect 1934 2343 1940 2344
rect 3838 2347 3844 2348
rect 3838 2343 3839 2347
rect 3843 2343 3844 2347
rect 4518 2344 4519 2348
rect 4523 2344 4524 2348
rect 4518 2343 4524 2344
rect 4662 2348 4668 2349
rect 4662 2344 4663 2348
rect 4667 2344 4668 2348
rect 4662 2343 4668 2344
rect 4822 2348 4828 2349
rect 4822 2344 4823 2348
rect 4827 2344 4828 2348
rect 4822 2343 4828 2344
rect 4990 2348 4996 2349
rect 4990 2344 4991 2348
rect 4995 2344 4996 2348
rect 4990 2343 4996 2344
rect 5166 2348 5172 2349
rect 5166 2344 5167 2348
rect 5171 2344 5172 2348
rect 5166 2343 5172 2344
rect 5350 2348 5356 2349
rect 5350 2344 5351 2348
rect 5355 2344 5356 2348
rect 5350 2343 5356 2344
rect 5542 2348 5548 2349
rect 5542 2344 5543 2348
rect 5547 2344 5548 2348
rect 5542 2343 5548 2344
rect 5662 2347 5668 2348
rect 5662 2343 5663 2347
rect 5667 2343 5668 2347
rect 1698 2342 1704 2343
rect 3838 2342 3844 2343
rect 5662 2342 5668 2343
rect 382 2332 388 2333
rect 110 2331 116 2332
rect 110 2327 111 2331
rect 115 2327 116 2331
rect 382 2328 383 2332
rect 387 2328 388 2332
rect 382 2327 388 2328
rect 534 2332 540 2333
rect 534 2328 535 2332
rect 539 2328 540 2332
rect 534 2327 540 2328
rect 702 2332 708 2333
rect 702 2328 703 2332
rect 707 2328 708 2332
rect 702 2327 708 2328
rect 886 2332 892 2333
rect 886 2328 887 2332
rect 891 2328 892 2332
rect 886 2327 892 2328
rect 1086 2332 1092 2333
rect 1086 2328 1087 2332
rect 1091 2328 1092 2332
rect 1086 2327 1092 2328
rect 1294 2332 1300 2333
rect 1294 2328 1295 2332
rect 1299 2328 1300 2332
rect 1294 2327 1300 2328
rect 1510 2332 1516 2333
rect 1510 2328 1511 2332
rect 1515 2328 1516 2332
rect 1510 2327 1516 2328
rect 1726 2332 1732 2333
rect 1726 2328 1727 2332
rect 1731 2328 1732 2332
rect 1726 2327 1732 2328
rect 1934 2331 1940 2332
rect 1934 2327 1935 2331
rect 1939 2327 1940 2331
rect 110 2326 116 2327
rect 1934 2326 1940 2327
rect 1974 2304 1980 2305
rect 3798 2304 3804 2305
rect 1974 2300 1975 2304
rect 1979 2300 1980 2304
rect 1974 2299 1980 2300
rect 2330 2303 2336 2304
rect 2330 2299 2331 2303
rect 2335 2299 2336 2303
rect 2330 2298 2336 2299
rect 2538 2303 2544 2304
rect 2538 2299 2539 2303
rect 2543 2299 2544 2303
rect 2538 2298 2544 2299
rect 2738 2303 2744 2304
rect 2738 2299 2739 2303
rect 2743 2299 2744 2303
rect 2738 2298 2744 2299
rect 2930 2303 2936 2304
rect 2930 2299 2931 2303
rect 2935 2299 2936 2303
rect 2930 2298 2936 2299
rect 3122 2303 3128 2304
rect 3122 2299 3123 2303
rect 3127 2299 3128 2303
rect 3122 2298 3128 2299
rect 3306 2303 3312 2304
rect 3306 2299 3307 2303
rect 3311 2299 3312 2303
rect 3306 2298 3312 2299
rect 3490 2303 3496 2304
rect 3490 2299 3491 2303
rect 3495 2299 3496 2303
rect 3490 2298 3496 2299
rect 3650 2303 3656 2304
rect 3650 2299 3651 2303
rect 3655 2299 3656 2303
rect 3798 2300 3799 2304
rect 3803 2300 3804 2304
rect 3798 2299 3804 2300
rect 3650 2298 3656 2299
rect 2358 2288 2364 2289
rect 1974 2287 1980 2288
rect 1974 2283 1975 2287
rect 1979 2283 1980 2287
rect 2358 2284 2359 2288
rect 2363 2284 2364 2288
rect 2358 2283 2364 2284
rect 2566 2288 2572 2289
rect 2566 2284 2567 2288
rect 2571 2284 2572 2288
rect 2566 2283 2572 2284
rect 2766 2288 2772 2289
rect 2766 2284 2767 2288
rect 2771 2284 2772 2288
rect 2766 2283 2772 2284
rect 2958 2288 2964 2289
rect 2958 2284 2959 2288
rect 2963 2284 2964 2288
rect 2958 2283 2964 2284
rect 3150 2288 3156 2289
rect 3150 2284 3151 2288
rect 3155 2284 3156 2288
rect 3150 2283 3156 2284
rect 3334 2288 3340 2289
rect 3334 2284 3335 2288
rect 3339 2284 3340 2288
rect 3334 2283 3340 2284
rect 3518 2288 3524 2289
rect 3518 2284 3519 2288
rect 3523 2284 3524 2288
rect 3518 2283 3524 2284
rect 3678 2288 3684 2289
rect 3678 2284 3679 2288
rect 3683 2284 3684 2288
rect 3678 2283 3684 2284
rect 3798 2287 3804 2288
rect 3798 2283 3799 2287
rect 3803 2283 3804 2287
rect 1974 2282 1980 2283
rect 3798 2282 3804 2283
rect 3838 2269 3844 2270
rect 5662 2269 5668 2270
rect 110 2265 116 2266
rect 1934 2265 1940 2266
rect 110 2261 111 2265
rect 115 2261 116 2265
rect 110 2260 116 2261
rect 158 2264 164 2265
rect 158 2260 159 2264
rect 163 2260 164 2264
rect 158 2259 164 2260
rect 334 2264 340 2265
rect 334 2260 335 2264
rect 339 2260 340 2264
rect 334 2259 340 2260
rect 542 2264 548 2265
rect 542 2260 543 2264
rect 547 2260 548 2264
rect 542 2259 548 2260
rect 758 2264 764 2265
rect 758 2260 759 2264
rect 763 2260 764 2264
rect 758 2259 764 2260
rect 974 2264 980 2265
rect 974 2260 975 2264
rect 979 2260 980 2264
rect 974 2259 980 2260
rect 1198 2264 1204 2265
rect 1198 2260 1199 2264
rect 1203 2260 1204 2264
rect 1198 2259 1204 2260
rect 1430 2264 1436 2265
rect 1430 2260 1431 2264
rect 1435 2260 1436 2264
rect 1430 2259 1436 2260
rect 1670 2264 1676 2265
rect 1670 2260 1671 2264
rect 1675 2260 1676 2264
rect 1934 2261 1935 2265
rect 1939 2261 1940 2265
rect 3838 2265 3839 2269
rect 3843 2265 3844 2269
rect 3838 2264 3844 2265
rect 3886 2268 3892 2269
rect 3886 2264 3887 2268
rect 3891 2264 3892 2268
rect 3886 2263 3892 2264
rect 4070 2268 4076 2269
rect 4070 2264 4071 2268
rect 4075 2264 4076 2268
rect 4070 2263 4076 2264
rect 4270 2268 4276 2269
rect 4270 2264 4271 2268
rect 4275 2264 4276 2268
rect 4270 2263 4276 2264
rect 4462 2268 4468 2269
rect 4462 2264 4463 2268
rect 4467 2264 4468 2268
rect 4462 2263 4468 2264
rect 4654 2268 4660 2269
rect 4654 2264 4655 2268
rect 4659 2264 4660 2268
rect 4654 2263 4660 2264
rect 4838 2268 4844 2269
rect 4838 2264 4839 2268
rect 4843 2264 4844 2268
rect 4838 2263 4844 2264
rect 5014 2268 5020 2269
rect 5014 2264 5015 2268
rect 5019 2264 5020 2268
rect 5014 2263 5020 2264
rect 5182 2268 5188 2269
rect 5182 2264 5183 2268
rect 5187 2264 5188 2268
rect 5182 2263 5188 2264
rect 5358 2268 5364 2269
rect 5358 2264 5359 2268
rect 5363 2264 5364 2268
rect 5358 2263 5364 2264
rect 5534 2268 5540 2269
rect 5534 2264 5535 2268
rect 5539 2264 5540 2268
rect 5662 2265 5663 2269
rect 5667 2265 5668 2269
rect 5662 2264 5668 2265
rect 5534 2263 5540 2264
rect 1934 2260 1940 2261
rect 1670 2259 1676 2260
rect 3858 2253 3864 2254
rect 3838 2252 3844 2253
rect 130 2249 136 2250
rect 110 2248 116 2249
rect 110 2244 111 2248
rect 115 2244 116 2248
rect 130 2245 131 2249
rect 135 2245 136 2249
rect 130 2244 136 2245
rect 306 2249 312 2250
rect 306 2245 307 2249
rect 311 2245 312 2249
rect 306 2244 312 2245
rect 514 2249 520 2250
rect 514 2245 515 2249
rect 519 2245 520 2249
rect 514 2244 520 2245
rect 730 2249 736 2250
rect 730 2245 731 2249
rect 735 2245 736 2249
rect 730 2244 736 2245
rect 946 2249 952 2250
rect 946 2245 947 2249
rect 951 2245 952 2249
rect 946 2244 952 2245
rect 1170 2249 1176 2250
rect 1170 2245 1171 2249
rect 1175 2245 1176 2249
rect 1170 2244 1176 2245
rect 1402 2249 1408 2250
rect 1402 2245 1403 2249
rect 1407 2245 1408 2249
rect 1402 2244 1408 2245
rect 1642 2249 1648 2250
rect 1642 2245 1643 2249
rect 1647 2245 1648 2249
rect 1642 2244 1648 2245
rect 1934 2248 1940 2249
rect 1934 2244 1935 2248
rect 1939 2244 1940 2248
rect 3838 2248 3839 2252
rect 3843 2248 3844 2252
rect 3858 2249 3859 2253
rect 3863 2249 3864 2253
rect 3858 2248 3864 2249
rect 4042 2253 4048 2254
rect 4042 2249 4043 2253
rect 4047 2249 4048 2253
rect 4042 2248 4048 2249
rect 4242 2253 4248 2254
rect 4242 2249 4243 2253
rect 4247 2249 4248 2253
rect 4242 2248 4248 2249
rect 4434 2253 4440 2254
rect 4434 2249 4435 2253
rect 4439 2249 4440 2253
rect 4434 2248 4440 2249
rect 4626 2253 4632 2254
rect 4626 2249 4627 2253
rect 4631 2249 4632 2253
rect 4626 2248 4632 2249
rect 4810 2253 4816 2254
rect 4810 2249 4811 2253
rect 4815 2249 4816 2253
rect 4810 2248 4816 2249
rect 4986 2253 4992 2254
rect 4986 2249 4987 2253
rect 4991 2249 4992 2253
rect 4986 2248 4992 2249
rect 5154 2253 5160 2254
rect 5154 2249 5155 2253
rect 5159 2249 5160 2253
rect 5154 2248 5160 2249
rect 5330 2253 5336 2254
rect 5330 2249 5331 2253
rect 5335 2249 5336 2253
rect 5330 2248 5336 2249
rect 5506 2253 5512 2254
rect 5506 2249 5507 2253
rect 5511 2249 5512 2253
rect 5506 2248 5512 2249
rect 5662 2252 5668 2253
rect 5662 2248 5663 2252
rect 5667 2248 5668 2252
rect 3838 2247 3844 2248
rect 5662 2247 5668 2248
rect 110 2243 116 2244
rect 1934 2243 1940 2244
rect 1974 2201 1980 2202
rect 3798 2201 3804 2202
rect 1974 2197 1975 2201
rect 1979 2197 1980 2201
rect 1974 2196 1980 2197
rect 2462 2200 2468 2201
rect 2462 2196 2463 2200
rect 2467 2196 2468 2200
rect 2462 2195 2468 2196
rect 2598 2200 2604 2201
rect 2598 2196 2599 2200
rect 2603 2196 2604 2200
rect 2598 2195 2604 2196
rect 2734 2200 2740 2201
rect 2734 2196 2735 2200
rect 2739 2196 2740 2200
rect 3798 2197 3799 2201
rect 3803 2197 3804 2201
rect 3798 2196 3804 2197
rect 2734 2195 2740 2196
rect 2434 2185 2440 2186
rect 1974 2184 1980 2185
rect 1974 2180 1975 2184
rect 1979 2180 1980 2184
rect 2434 2181 2435 2185
rect 2439 2181 2440 2185
rect 2434 2180 2440 2181
rect 2570 2185 2576 2186
rect 2570 2181 2571 2185
rect 2575 2181 2576 2185
rect 2570 2180 2576 2181
rect 2706 2185 2712 2186
rect 2706 2181 2707 2185
rect 2711 2181 2712 2185
rect 2706 2180 2712 2181
rect 3798 2184 3804 2185
rect 3798 2180 3799 2184
rect 3803 2180 3804 2184
rect 1974 2179 1980 2180
rect 3798 2179 3804 2180
rect 3838 2120 3844 2121
rect 5662 2120 5668 2121
rect 3838 2116 3839 2120
rect 3843 2116 3844 2120
rect 3838 2115 3844 2116
rect 3858 2119 3864 2120
rect 3858 2115 3859 2119
rect 3863 2115 3864 2119
rect 3858 2114 3864 2115
rect 4042 2119 4048 2120
rect 4042 2115 4043 2119
rect 4047 2115 4048 2119
rect 4042 2114 4048 2115
rect 4250 2119 4256 2120
rect 4250 2115 4251 2119
rect 4255 2115 4256 2119
rect 4250 2114 4256 2115
rect 4458 2119 4464 2120
rect 4458 2115 4459 2119
rect 4463 2115 4464 2119
rect 4458 2114 4464 2115
rect 4658 2119 4664 2120
rect 4658 2115 4659 2119
rect 4663 2115 4664 2119
rect 4658 2114 4664 2115
rect 4850 2119 4856 2120
rect 4850 2115 4851 2119
rect 4855 2115 4856 2119
rect 4850 2114 4856 2115
rect 5034 2119 5040 2120
rect 5034 2115 5035 2119
rect 5039 2115 5040 2119
rect 5034 2114 5040 2115
rect 5218 2119 5224 2120
rect 5218 2115 5219 2119
rect 5223 2115 5224 2119
rect 5218 2114 5224 2115
rect 5410 2119 5416 2120
rect 5410 2115 5411 2119
rect 5415 2115 5416 2119
rect 5662 2116 5663 2120
rect 5667 2116 5668 2120
rect 5662 2115 5668 2116
rect 5410 2114 5416 2115
rect 3886 2104 3892 2105
rect 3838 2103 3844 2104
rect 3838 2099 3839 2103
rect 3843 2099 3844 2103
rect 3886 2100 3887 2104
rect 3891 2100 3892 2104
rect 3886 2099 3892 2100
rect 4070 2104 4076 2105
rect 4070 2100 4071 2104
rect 4075 2100 4076 2104
rect 4070 2099 4076 2100
rect 4278 2104 4284 2105
rect 4278 2100 4279 2104
rect 4283 2100 4284 2104
rect 4278 2099 4284 2100
rect 4486 2104 4492 2105
rect 4486 2100 4487 2104
rect 4491 2100 4492 2104
rect 4486 2099 4492 2100
rect 4686 2104 4692 2105
rect 4686 2100 4687 2104
rect 4691 2100 4692 2104
rect 4686 2099 4692 2100
rect 4878 2104 4884 2105
rect 4878 2100 4879 2104
rect 4883 2100 4884 2104
rect 4878 2099 4884 2100
rect 5062 2104 5068 2105
rect 5062 2100 5063 2104
rect 5067 2100 5068 2104
rect 5062 2099 5068 2100
rect 5246 2104 5252 2105
rect 5246 2100 5247 2104
rect 5251 2100 5252 2104
rect 5246 2099 5252 2100
rect 5438 2104 5444 2105
rect 5438 2100 5439 2104
rect 5443 2100 5444 2104
rect 5438 2099 5444 2100
rect 5662 2103 5668 2104
rect 5662 2099 5663 2103
rect 5667 2099 5668 2103
rect 3838 2098 3844 2099
rect 5662 2098 5668 2099
rect 110 2096 116 2097
rect 1934 2096 1940 2097
rect 110 2092 111 2096
rect 115 2092 116 2096
rect 110 2091 116 2092
rect 130 2095 136 2096
rect 130 2091 131 2095
rect 135 2091 136 2095
rect 130 2090 136 2091
rect 298 2095 304 2096
rect 298 2091 299 2095
rect 303 2091 304 2095
rect 298 2090 304 2091
rect 498 2095 504 2096
rect 498 2091 499 2095
rect 503 2091 504 2095
rect 498 2090 504 2091
rect 714 2095 720 2096
rect 714 2091 715 2095
rect 719 2091 720 2095
rect 714 2090 720 2091
rect 930 2095 936 2096
rect 930 2091 931 2095
rect 935 2091 936 2095
rect 930 2090 936 2091
rect 1154 2095 1160 2096
rect 1154 2091 1155 2095
rect 1159 2091 1160 2095
rect 1154 2090 1160 2091
rect 1386 2095 1392 2096
rect 1386 2091 1387 2095
rect 1391 2091 1392 2095
rect 1386 2090 1392 2091
rect 1626 2095 1632 2096
rect 1626 2091 1627 2095
rect 1631 2091 1632 2095
rect 1934 2092 1935 2096
rect 1939 2092 1940 2096
rect 1934 2091 1940 2092
rect 1626 2090 1632 2091
rect 158 2080 164 2081
rect 110 2079 116 2080
rect 110 2075 111 2079
rect 115 2075 116 2079
rect 158 2076 159 2080
rect 163 2076 164 2080
rect 158 2075 164 2076
rect 326 2080 332 2081
rect 326 2076 327 2080
rect 331 2076 332 2080
rect 326 2075 332 2076
rect 526 2080 532 2081
rect 526 2076 527 2080
rect 531 2076 532 2080
rect 526 2075 532 2076
rect 742 2080 748 2081
rect 742 2076 743 2080
rect 747 2076 748 2080
rect 742 2075 748 2076
rect 958 2080 964 2081
rect 958 2076 959 2080
rect 963 2076 964 2080
rect 958 2075 964 2076
rect 1182 2080 1188 2081
rect 1182 2076 1183 2080
rect 1187 2076 1188 2080
rect 1182 2075 1188 2076
rect 1414 2080 1420 2081
rect 1414 2076 1415 2080
rect 1419 2076 1420 2080
rect 1414 2075 1420 2076
rect 1654 2080 1660 2081
rect 1654 2076 1655 2080
rect 1659 2076 1660 2080
rect 1654 2075 1660 2076
rect 1934 2079 1940 2080
rect 1934 2075 1935 2079
rect 1939 2075 1940 2079
rect 110 2074 116 2075
rect 1934 2074 1940 2075
rect 3838 2025 3844 2026
rect 5662 2025 5668 2026
rect 3838 2021 3839 2025
rect 3843 2021 3844 2025
rect 1974 2020 1980 2021
rect 3798 2020 3804 2021
rect 3838 2020 3844 2021
rect 4286 2024 4292 2025
rect 4286 2020 4287 2024
rect 4291 2020 4292 2024
rect 1974 2016 1975 2020
rect 1979 2016 1980 2020
rect 1974 2015 1980 2016
rect 2418 2019 2424 2020
rect 2418 2015 2419 2019
rect 2423 2015 2424 2019
rect 2418 2014 2424 2015
rect 2610 2019 2616 2020
rect 2610 2015 2611 2019
rect 2615 2015 2616 2019
rect 2610 2014 2616 2015
rect 2794 2019 2800 2020
rect 2794 2015 2795 2019
rect 2799 2015 2800 2019
rect 2794 2014 2800 2015
rect 2978 2019 2984 2020
rect 2978 2015 2979 2019
rect 2983 2015 2984 2019
rect 2978 2014 2984 2015
rect 3154 2019 3160 2020
rect 3154 2015 3155 2019
rect 3159 2015 3160 2019
rect 3154 2014 3160 2015
rect 3322 2019 3328 2020
rect 3322 2015 3323 2019
rect 3327 2015 3328 2019
rect 3322 2014 3328 2015
rect 3498 2019 3504 2020
rect 3498 2015 3499 2019
rect 3503 2015 3504 2019
rect 3498 2014 3504 2015
rect 3650 2019 3656 2020
rect 3650 2015 3651 2019
rect 3655 2015 3656 2019
rect 3798 2016 3799 2020
rect 3803 2016 3804 2020
rect 4286 2019 4292 2020
rect 4422 2024 4428 2025
rect 4422 2020 4423 2024
rect 4427 2020 4428 2024
rect 4422 2019 4428 2020
rect 4558 2024 4564 2025
rect 4558 2020 4559 2024
rect 4563 2020 4564 2024
rect 4558 2019 4564 2020
rect 4694 2024 4700 2025
rect 4694 2020 4695 2024
rect 4699 2020 4700 2024
rect 4694 2019 4700 2020
rect 4838 2024 4844 2025
rect 4838 2020 4839 2024
rect 4843 2020 4844 2024
rect 5662 2021 5663 2025
rect 5667 2021 5668 2025
rect 5662 2020 5668 2021
rect 4838 2019 4844 2020
rect 3798 2015 3804 2016
rect 3650 2014 3656 2015
rect 110 2013 116 2014
rect 1934 2013 1940 2014
rect 110 2009 111 2013
rect 115 2009 116 2013
rect 110 2008 116 2009
rect 158 2012 164 2013
rect 158 2008 159 2012
rect 163 2008 164 2012
rect 158 2007 164 2008
rect 342 2012 348 2013
rect 342 2008 343 2012
rect 347 2008 348 2012
rect 342 2007 348 2008
rect 566 2012 572 2013
rect 566 2008 567 2012
rect 571 2008 572 2012
rect 566 2007 572 2008
rect 806 2012 812 2013
rect 806 2008 807 2012
rect 811 2008 812 2012
rect 806 2007 812 2008
rect 1062 2012 1068 2013
rect 1062 2008 1063 2012
rect 1067 2008 1068 2012
rect 1062 2007 1068 2008
rect 1334 2012 1340 2013
rect 1334 2008 1335 2012
rect 1339 2008 1340 2012
rect 1334 2007 1340 2008
rect 1606 2012 1612 2013
rect 1606 2008 1607 2012
rect 1611 2008 1612 2012
rect 1934 2009 1935 2013
rect 1939 2009 1940 2013
rect 4258 2009 4264 2010
rect 1934 2008 1940 2009
rect 3838 2008 3844 2009
rect 1606 2007 1612 2008
rect 2446 2004 2452 2005
rect 1974 2003 1980 2004
rect 1974 1999 1975 2003
rect 1979 1999 1980 2003
rect 2446 2000 2447 2004
rect 2451 2000 2452 2004
rect 2446 1999 2452 2000
rect 2638 2004 2644 2005
rect 2638 2000 2639 2004
rect 2643 2000 2644 2004
rect 2638 1999 2644 2000
rect 2822 2004 2828 2005
rect 2822 2000 2823 2004
rect 2827 2000 2828 2004
rect 2822 1999 2828 2000
rect 3006 2004 3012 2005
rect 3006 2000 3007 2004
rect 3011 2000 3012 2004
rect 3006 1999 3012 2000
rect 3182 2004 3188 2005
rect 3182 2000 3183 2004
rect 3187 2000 3188 2004
rect 3182 1999 3188 2000
rect 3350 2004 3356 2005
rect 3350 2000 3351 2004
rect 3355 2000 3356 2004
rect 3350 1999 3356 2000
rect 3526 2004 3532 2005
rect 3526 2000 3527 2004
rect 3531 2000 3532 2004
rect 3526 1999 3532 2000
rect 3678 2004 3684 2005
rect 3838 2004 3839 2008
rect 3843 2004 3844 2008
rect 4258 2005 4259 2009
rect 4263 2005 4264 2009
rect 4258 2004 4264 2005
rect 4394 2009 4400 2010
rect 4394 2005 4395 2009
rect 4399 2005 4400 2009
rect 4394 2004 4400 2005
rect 4530 2009 4536 2010
rect 4530 2005 4531 2009
rect 4535 2005 4536 2009
rect 4530 2004 4536 2005
rect 4666 2009 4672 2010
rect 4666 2005 4667 2009
rect 4671 2005 4672 2009
rect 4666 2004 4672 2005
rect 4810 2009 4816 2010
rect 4810 2005 4811 2009
rect 4815 2005 4816 2009
rect 4810 2004 4816 2005
rect 5662 2008 5668 2009
rect 5662 2004 5663 2008
rect 5667 2004 5668 2008
rect 3678 2000 3679 2004
rect 3683 2000 3684 2004
rect 3678 1999 3684 2000
rect 3798 2003 3804 2004
rect 3838 2003 3844 2004
rect 5662 2003 5668 2004
rect 3798 1999 3799 2003
rect 3803 1999 3804 2003
rect 1974 1998 1980 1999
rect 3798 1998 3804 1999
rect 130 1997 136 1998
rect 110 1996 116 1997
rect 110 1992 111 1996
rect 115 1992 116 1996
rect 130 1993 131 1997
rect 135 1993 136 1997
rect 130 1992 136 1993
rect 314 1997 320 1998
rect 314 1993 315 1997
rect 319 1993 320 1997
rect 314 1992 320 1993
rect 538 1997 544 1998
rect 538 1993 539 1997
rect 543 1993 544 1997
rect 538 1992 544 1993
rect 778 1997 784 1998
rect 778 1993 779 1997
rect 783 1993 784 1997
rect 778 1992 784 1993
rect 1034 1997 1040 1998
rect 1034 1993 1035 1997
rect 1039 1993 1040 1997
rect 1034 1992 1040 1993
rect 1306 1997 1312 1998
rect 1306 1993 1307 1997
rect 1311 1993 1312 1997
rect 1306 1992 1312 1993
rect 1578 1997 1584 1998
rect 1578 1993 1579 1997
rect 1583 1993 1584 1997
rect 1578 1992 1584 1993
rect 1934 1996 1940 1997
rect 1934 1992 1935 1996
rect 1939 1992 1940 1996
rect 110 1991 116 1992
rect 1934 1991 1940 1992
rect 1974 1933 1980 1934
rect 3798 1933 3804 1934
rect 1974 1929 1975 1933
rect 1979 1929 1980 1933
rect 1974 1928 1980 1929
rect 2358 1932 2364 1933
rect 2358 1928 2359 1932
rect 2363 1928 2364 1932
rect 2358 1927 2364 1928
rect 2494 1932 2500 1933
rect 2494 1928 2495 1932
rect 2499 1928 2500 1932
rect 2494 1927 2500 1928
rect 2630 1932 2636 1933
rect 2630 1928 2631 1932
rect 2635 1928 2636 1932
rect 2630 1927 2636 1928
rect 2766 1932 2772 1933
rect 2766 1928 2767 1932
rect 2771 1928 2772 1932
rect 2766 1927 2772 1928
rect 2902 1932 2908 1933
rect 2902 1928 2903 1932
rect 2907 1928 2908 1932
rect 2902 1927 2908 1928
rect 3038 1932 3044 1933
rect 3038 1928 3039 1932
rect 3043 1928 3044 1932
rect 3038 1927 3044 1928
rect 3174 1932 3180 1933
rect 3174 1928 3175 1932
rect 3179 1928 3180 1932
rect 3174 1927 3180 1928
rect 3318 1932 3324 1933
rect 3318 1928 3319 1932
rect 3323 1928 3324 1932
rect 3798 1929 3799 1933
rect 3803 1929 3804 1933
rect 3798 1928 3804 1929
rect 3318 1927 3324 1928
rect 2330 1917 2336 1918
rect 1974 1916 1980 1917
rect 1974 1912 1975 1916
rect 1979 1912 1980 1916
rect 2330 1913 2331 1917
rect 2335 1913 2336 1917
rect 2330 1912 2336 1913
rect 2466 1917 2472 1918
rect 2466 1913 2467 1917
rect 2471 1913 2472 1917
rect 2466 1912 2472 1913
rect 2602 1917 2608 1918
rect 2602 1913 2603 1917
rect 2607 1913 2608 1917
rect 2602 1912 2608 1913
rect 2738 1917 2744 1918
rect 2738 1913 2739 1917
rect 2743 1913 2744 1917
rect 2738 1912 2744 1913
rect 2874 1917 2880 1918
rect 2874 1913 2875 1917
rect 2879 1913 2880 1917
rect 2874 1912 2880 1913
rect 3010 1917 3016 1918
rect 3010 1913 3011 1917
rect 3015 1913 3016 1917
rect 3010 1912 3016 1913
rect 3146 1917 3152 1918
rect 3146 1913 3147 1917
rect 3151 1913 3152 1917
rect 3146 1912 3152 1913
rect 3290 1917 3296 1918
rect 3290 1913 3291 1917
rect 3295 1913 3296 1917
rect 3290 1912 3296 1913
rect 3798 1916 3804 1917
rect 3798 1912 3799 1916
rect 3803 1912 3804 1916
rect 1974 1911 1980 1912
rect 3798 1911 3804 1912
rect 110 1860 116 1861
rect 1934 1860 1940 1861
rect 110 1856 111 1860
rect 115 1856 116 1860
rect 110 1855 116 1856
rect 330 1859 336 1860
rect 330 1855 331 1859
rect 335 1855 336 1859
rect 330 1854 336 1855
rect 498 1859 504 1860
rect 498 1855 499 1859
rect 503 1855 504 1859
rect 498 1854 504 1855
rect 666 1859 672 1860
rect 666 1855 667 1859
rect 671 1855 672 1859
rect 666 1854 672 1855
rect 842 1859 848 1860
rect 842 1855 843 1859
rect 847 1855 848 1859
rect 842 1854 848 1855
rect 1026 1859 1032 1860
rect 1026 1855 1027 1859
rect 1031 1855 1032 1859
rect 1026 1854 1032 1855
rect 1218 1859 1224 1860
rect 1218 1855 1219 1859
rect 1223 1855 1224 1859
rect 1218 1854 1224 1855
rect 1410 1859 1416 1860
rect 1410 1855 1411 1859
rect 1415 1855 1416 1859
rect 1410 1854 1416 1855
rect 1602 1859 1608 1860
rect 1602 1855 1603 1859
rect 1607 1855 1608 1859
rect 1934 1856 1935 1860
rect 1939 1856 1940 1860
rect 1934 1855 1940 1856
rect 3838 1856 3844 1857
rect 5662 1856 5668 1857
rect 1602 1854 1608 1855
rect 3838 1852 3839 1856
rect 3843 1852 3844 1856
rect 3838 1851 3844 1852
rect 3954 1855 3960 1856
rect 3954 1851 3955 1855
rect 3959 1851 3960 1855
rect 3954 1850 3960 1851
rect 4194 1855 4200 1856
rect 4194 1851 4195 1855
rect 4199 1851 4200 1855
rect 4194 1850 4200 1851
rect 4466 1855 4472 1856
rect 4466 1851 4467 1855
rect 4471 1851 4472 1855
rect 4466 1850 4472 1851
rect 4770 1855 4776 1856
rect 4770 1851 4771 1855
rect 4775 1851 4776 1855
rect 4770 1850 4776 1851
rect 5090 1855 5096 1856
rect 5090 1851 5091 1855
rect 5095 1851 5096 1855
rect 5090 1850 5096 1851
rect 5410 1855 5416 1856
rect 5410 1851 5411 1855
rect 5415 1851 5416 1855
rect 5662 1852 5663 1856
rect 5667 1852 5668 1856
rect 5662 1851 5668 1852
rect 5410 1850 5416 1851
rect 358 1844 364 1845
rect 110 1843 116 1844
rect 110 1839 111 1843
rect 115 1839 116 1843
rect 358 1840 359 1844
rect 363 1840 364 1844
rect 358 1839 364 1840
rect 526 1844 532 1845
rect 526 1840 527 1844
rect 531 1840 532 1844
rect 526 1839 532 1840
rect 694 1844 700 1845
rect 694 1840 695 1844
rect 699 1840 700 1844
rect 694 1839 700 1840
rect 870 1844 876 1845
rect 870 1840 871 1844
rect 875 1840 876 1844
rect 870 1839 876 1840
rect 1054 1844 1060 1845
rect 1054 1840 1055 1844
rect 1059 1840 1060 1844
rect 1054 1839 1060 1840
rect 1246 1844 1252 1845
rect 1246 1840 1247 1844
rect 1251 1840 1252 1844
rect 1246 1839 1252 1840
rect 1438 1844 1444 1845
rect 1438 1840 1439 1844
rect 1443 1840 1444 1844
rect 1438 1839 1444 1840
rect 1630 1844 1636 1845
rect 1630 1840 1631 1844
rect 1635 1840 1636 1844
rect 1630 1839 1636 1840
rect 1934 1843 1940 1844
rect 1934 1839 1935 1843
rect 1939 1839 1940 1843
rect 3982 1840 3988 1841
rect 110 1838 116 1839
rect 1934 1838 1940 1839
rect 3838 1839 3844 1840
rect 3838 1835 3839 1839
rect 3843 1835 3844 1839
rect 3982 1836 3983 1840
rect 3987 1836 3988 1840
rect 3982 1835 3988 1836
rect 4222 1840 4228 1841
rect 4222 1836 4223 1840
rect 4227 1836 4228 1840
rect 4222 1835 4228 1836
rect 4494 1840 4500 1841
rect 4494 1836 4495 1840
rect 4499 1836 4500 1840
rect 4494 1835 4500 1836
rect 4798 1840 4804 1841
rect 4798 1836 4799 1840
rect 4803 1836 4804 1840
rect 4798 1835 4804 1836
rect 5118 1840 5124 1841
rect 5118 1836 5119 1840
rect 5123 1836 5124 1840
rect 5118 1835 5124 1836
rect 5438 1840 5444 1841
rect 5438 1836 5439 1840
rect 5443 1836 5444 1840
rect 5438 1835 5444 1836
rect 5662 1839 5668 1840
rect 5662 1835 5663 1839
rect 5667 1835 5668 1839
rect 3838 1834 3844 1835
rect 5662 1834 5668 1835
rect 1974 1784 1980 1785
rect 3798 1784 3804 1785
rect 1974 1780 1975 1784
rect 1979 1780 1980 1784
rect 1974 1779 1980 1780
rect 2210 1783 2216 1784
rect 2210 1779 2211 1783
rect 2215 1779 2216 1783
rect 2210 1778 2216 1779
rect 2354 1783 2360 1784
rect 2354 1779 2355 1783
rect 2359 1779 2360 1783
rect 2354 1778 2360 1779
rect 2498 1783 2504 1784
rect 2498 1779 2499 1783
rect 2503 1779 2504 1783
rect 2498 1778 2504 1779
rect 2642 1783 2648 1784
rect 2642 1779 2643 1783
rect 2647 1779 2648 1783
rect 2642 1778 2648 1779
rect 2786 1783 2792 1784
rect 2786 1779 2787 1783
rect 2791 1779 2792 1783
rect 2786 1778 2792 1779
rect 2930 1783 2936 1784
rect 2930 1779 2931 1783
rect 2935 1779 2936 1783
rect 2930 1778 2936 1779
rect 3082 1783 3088 1784
rect 3082 1779 3083 1783
rect 3087 1779 3088 1783
rect 3798 1780 3799 1784
rect 3803 1780 3804 1784
rect 3798 1779 3804 1780
rect 3838 1781 3844 1782
rect 5662 1781 5668 1782
rect 3082 1778 3088 1779
rect 3838 1777 3839 1781
rect 3843 1777 3844 1781
rect 3838 1776 3844 1777
rect 4366 1780 4372 1781
rect 4366 1776 4367 1780
rect 4371 1776 4372 1780
rect 4366 1775 4372 1776
rect 4574 1780 4580 1781
rect 4574 1776 4575 1780
rect 4579 1776 4580 1780
rect 4574 1775 4580 1776
rect 4782 1780 4788 1781
rect 4782 1776 4783 1780
rect 4787 1776 4788 1780
rect 4782 1775 4788 1776
rect 4982 1780 4988 1781
rect 4982 1776 4983 1780
rect 4987 1776 4988 1780
rect 4982 1775 4988 1776
rect 5174 1780 5180 1781
rect 5174 1776 5175 1780
rect 5179 1776 5180 1780
rect 5174 1775 5180 1776
rect 5366 1780 5372 1781
rect 5366 1776 5367 1780
rect 5371 1776 5372 1780
rect 5366 1775 5372 1776
rect 5542 1780 5548 1781
rect 5542 1776 5543 1780
rect 5547 1776 5548 1780
rect 5662 1777 5663 1781
rect 5667 1777 5668 1781
rect 5662 1776 5668 1777
rect 5542 1775 5548 1776
rect 110 1773 116 1774
rect 1934 1773 1940 1774
rect 110 1769 111 1773
rect 115 1769 116 1773
rect 110 1768 116 1769
rect 534 1772 540 1773
rect 534 1768 535 1772
rect 539 1768 540 1772
rect 534 1767 540 1768
rect 694 1772 700 1773
rect 694 1768 695 1772
rect 699 1768 700 1772
rect 694 1767 700 1768
rect 854 1772 860 1773
rect 854 1768 855 1772
rect 859 1768 860 1772
rect 854 1767 860 1768
rect 1014 1772 1020 1773
rect 1014 1768 1015 1772
rect 1019 1768 1020 1772
rect 1014 1767 1020 1768
rect 1182 1772 1188 1773
rect 1182 1768 1183 1772
rect 1187 1768 1188 1772
rect 1182 1767 1188 1768
rect 1350 1772 1356 1773
rect 1350 1768 1351 1772
rect 1355 1768 1356 1772
rect 1350 1767 1356 1768
rect 1518 1772 1524 1773
rect 1518 1768 1519 1772
rect 1523 1768 1524 1772
rect 1934 1769 1935 1773
rect 1939 1769 1940 1773
rect 1934 1768 1940 1769
rect 2238 1768 2244 1769
rect 1518 1767 1524 1768
rect 1974 1767 1980 1768
rect 1974 1763 1975 1767
rect 1979 1763 1980 1767
rect 2238 1764 2239 1768
rect 2243 1764 2244 1768
rect 2238 1763 2244 1764
rect 2382 1768 2388 1769
rect 2382 1764 2383 1768
rect 2387 1764 2388 1768
rect 2382 1763 2388 1764
rect 2526 1768 2532 1769
rect 2526 1764 2527 1768
rect 2531 1764 2532 1768
rect 2526 1763 2532 1764
rect 2670 1768 2676 1769
rect 2670 1764 2671 1768
rect 2675 1764 2676 1768
rect 2670 1763 2676 1764
rect 2814 1768 2820 1769
rect 2814 1764 2815 1768
rect 2819 1764 2820 1768
rect 2814 1763 2820 1764
rect 2958 1768 2964 1769
rect 2958 1764 2959 1768
rect 2963 1764 2964 1768
rect 2958 1763 2964 1764
rect 3110 1768 3116 1769
rect 3110 1764 3111 1768
rect 3115 1764 3116 1768
rect 3110 1763 3116 1764
rect 3798 1767 3804 1768
rect 3798 1763 3799 1767
rect 3803 1763 3804 1767
rect 4338 1765 4344 1766
rect 1974 1762 1980 1763
rect 3798 1762 3804 1763
rect 3838 1764 3844 1765
rect 3838 1760 3839 1764
rect 3843 1760 3844 1764
rect 4338 1761 4339 1765
rect 4343 1761 4344 1765
rect 4338 1760 4344 1761
rect 4546 1765 4552 1766
rect 4546 1761 4547 1765
rect 4551 1761 4552 1765
rect 4546 1760 4552 1761
rect 4754 1765 4760 1766
rect 4754 1761 4755 1765
rect 4759 1761 4760 1765
rect 4754 1760 4760 1761
rect 4954 1765 4960 1766
rect 4954 1761 4955 1765
rect 4959 1761 4960 1765
rect 4954 1760 4960 1761
rect 5146 1765 5152 1766
rect 5146 1761 5147 1765
rect 5151 1761 5152 1765
rect 5146 1760 5152 1761
rect 5338 1765 5344 1766
rect 5338 1761 5339 1765
rect 5343 1761 5344 1765
rect 5338 1760 5344 1761
rect 5514 1765 5520 1766
rect 5514 1761 5515 1765
rect 5519 1761 5520 1765
rect 5514 1760 5520 1761
rect 5662 1764 5668 1765
rect 5662 1760 5663 1764
rect 5667 1760 5668 1764
rect 3838 1759 3844 1760
rect 5662 1759 5668 1760
rect 506 1757 512 1758
rect 110 1756 116 1757
rect 110 1752 111 1756
rect 115 1752 116 1756
rect 506 1753 507 1757
rect 511 1753 512 1757
rect 506 1752 512 1753
rect 666 1757 672 1758
rect 666 1753 667 1757
rect 671 1753 672 1757
rect 666 1752 672 1753
rect 826 1757 832 1758
rect 826 1753 827 1757
rect 831 1753 832 1757
rect 826 1752 832 1753
rect 986 1757 992 1758
rect 986 1753 987 1757
rect 991 1753 992 1757
rect 986 1752 992 1753
rect 1154 1757 1160 1758
rect 1154 1753 1155 1757
rect 1159 1753 1160 1757
rect 1154 1752 1160 1753
rect 1322 1757 1328 1758
rect 1322 1753 1323 1757
rect 1327 1753 1328 1757
rect 1322 1752 1328 1753
rect 1490 1757 1496 1758
rect 1490 1753 1491 1757
rect 1495 1753 1496 1757
rect 1490 1752 1496 1753
rect 1934 1756 1940 1757
rect 1934 1752 1935 1756
rect 1939 1752 1940 1756
rect 110 1751 116 1752
rect 1934 1751 1940 1752
rect 1974 1709 1980 1710
rect 3798 1709 3804 1710
rect 1974 1705 1975 1709
rect 1979 1705 1980 1709
rect 1974 1704 1980 1705
rect 2022 1708 2028 1709
rect 2022 1704 2023 1708
rect 2027 1704 2028 1708
rect 2022 1703 2028 1704
rect 2214 1708 2220 1709
rect 2214 1704 2215 1708
rect 2219 1704 2220 1708
rect 2214 1703 2220 1704
rect 2406 1708 2412 1709
rect 2406 1704 2407 1708
rect 2411 1704 2412 1708
rect 2406 1703 2412 1704
rect 2598 1708 2604 1709
rect 2598 1704 2599 1708
rect 2603 1704 2604 1708
rect 2598 1703 2604 1704
rect 2790 1708 2796 1709
rect 2790 1704 2791 1708
rect 2795 1704 2796 1708
rect 2790 1703 2796 1704
rect 2974 1708 2980 1709
rect 2974 1704 2975 1708
rect 2979 1704 2980 1708
rect 2974 1703 2980 1704
rect 3150 1708 3156 1709
rect 3150 1704 3151 1708
rect 3155 1704 3156 1708
rect 3150 1703 3156 1704
rect 3334 1708 3340 1709
rect 3334 1704 3335 1708
rect 3339 1704 3340 1708
rect 3334 1703 3340 1704
rect 3518 1708 3524 1709
rect 3518 1704 3519 1708
rect 3523 1704 3524 1708
rect 3798 1705 3799 1709
rect 3803 1705 3804 1709
rect 3798 1704 3804 1705
rect 3518 1703 3524 1704
rect 1994 1693 2000 1694
rect 1974 1692 1980 1693
rect 1974 1688 1975 1692
rect 1979 1688 1980 1692
rect 1994 1689 1995 1693
rect 1999 1689 2000 1693
rect 1994 1688 2000 1689
rect 2186 1693 2192 1694
rect 2186 1689 2187 1693
rect 2191 1689 2192 1693
rect 2186 1688 2192 1689
rect 2378 1693 2384 1694
rect 2378 1689 2379 1693
rect 2383 1689 2384 1693
rect 2378 1688 2384 1689
rect 2570 1693 2576 1694
rect 2570 1689 2571 1693
rect 2575 1689 2576 1693
rect 2570 1688 2576 1689
rect 2762 1693 2768 1694
rect 2762 1689 2763 1693
rect 2767 1689 2768 1693
rect 2762 1688 2768 1689
rect 2946 1693 2952 1694
rect 2946 1689 2947 1693
rect 2951 1689 2952 1693
rect 2946 1688 2952 1689
rect 3122 1693 3128 1694
rect 3122 1689 3123 1693
rect 3127 1689 3128 1693
rect 3122 1688 3128 1689
rect 3306 1693 3312 1694
rect 3306 1689 3307 1693
rect 3311 1689 3312 1693
rect 3306 1688 3312 1689
rect 3490 1693 3496 1694
rect 3490 1689 3491 1693
rect 3495 1689 3496 1693
rect 3490 1688 3496 1689
rect 3798 1692 3804 1693
rect 3798 1688 3799 1692
rect 3803 1688 3804 1692
rect 1974 1687 1980 1688
rect 3798 1687 3804 1688
rect 3838 1616 3844 1617
rect 5662 1616 5668 1617
rect 3838 1612 3839 1616
rect 3843 1612 3844 1616
rect 3838 1611 3844 1612
rect 4602 1615 4608 1616
rect 4602 1611 4603 1615
rect 4607 1611 4608 1615
rect 4602 1610 4608 1611
rect 4786 1615 4792 1616
rect 4786 1611 4787 1615
rect 4791 1611 4792 1615
rect 4786 1610 4792 1611
rect 4970 1615 4976 1616
rect 4970 1611 4971 1615
rect 4975 1611 4976 1615
rect 4970 1610 4976 1611
rect 5154 1615 5160 1616
rect 5154 1611 5155 1615
rect 5159 1611 5160 1615
rect 5154 1610 5160 1611
rect 5338 1615 5344 1616
rect 5338 1611 5339 1615
rect 5343 1611 5344 1615
rect 5338 1610 5344 1611
rect 5514 1615 5520 1616
rect 5514 1611 5515 1615
rect 5519 1611 5520 1615
rect 5662 1612 5663 1616
rect 5667 1612 5668 1616
rect 5662 1611 5668 1612
rect 5514 1610 5520 1611
rect 110 1608 116 1609
rect 1934 1608 1940 1609
rect 110 1604 111 1608
rect 115 1604 116 1608
rect 110 1603 116 1604
rect 426 1607 432 1608
rect 426 1603 427 1607
rect 431 1603 432 1607
rect 426 1602 432 1603
rect 610 1607 616 1608
rect 610 1603 611 1607
rect 615 1603 616 1607
rect 610 1602 616 1603
rect 802 1607 808 1608
rect 802 1603 803 1607
rect 807 1603 808 1607
rect 802 1602 808 1603
rect 994 1607 1000 1608
rect 994 1603 995 1607
rect 999 1603 1000 1607
rect 994 1602 1000 1603
rect 1186 1607 1192 1608
rect 1186 1603 1187 1607
rect 1191 1603 1192 1607
rect 1186 1602 1192 1603
rect 1378 1607 1384 1608
rect 1378 1603 1379 1607
rect 1383 1603 1384 1607
rect 1934 1604 1935 1608
rect 1939 1604 1940 1608
rect 1934 1603 1940 1604
rect 1378 1602 1384 1603
rect 4630 1600 4636 1601
rect 3838 1599 3844 1600
rect 3838 1595 3839 1599
rect 3843 1595 3844 1599
rect 4630 1596 4631 1600
rect 4635 1596 4636 1600
rect 4630 1595 4636 1596
rect 4814 1600 4820 1601
rect 4814 1596 4815 1600
rect 4819 1596 4820 1600
rect 4814 1595 4820 1596
rect 4998 1600 5004 1601
rect 4998 1596 4999 1600
rect 5003 1596 5004 1600
rect 4998 1595 5004 1596
rect 5182 1600 5188 1601
rect 5182 1596 5183 1600
rect 5187 1596 5188 1600
rect 5182 1595 5188 1596
rect 5366 1600 5372 1601
rect 5366 1596 5367 1600
rect 5371 1596 5372 1600
rect 5366 1595 5372 1596
rect 5542 1600 5548 1601
rect 5542 1596 5543 1600
rect 5547 1596 5548 1600
rect 5542 1595 5548 1596
rect 5662 1599 5668 1600
rect 5662 1595 5663 1599
rect 5667 1595 5668 1599
rect 3838 1594 3844 1595
rect 5662 1594 5668 1595
rect 454 1592 460 1593
rect 110 1591 116 1592
rect 110 1587 111 1591
rect 115 1587 116 1591
rect 454 1588 455 1592
rect 459 1588 460 1592
rect 454 1587 460 1588
rect 638 1592 644 1593
rect 638 1588 639 1592
rect 643 1588 644 1592
rect 638 1587 644 1588
rect 830 1592 836 1593
rect 830 1588 831 1592
rect 835 1588 836 1592
rect 830 1587 836 1588
rect 1022 1592 1028 1593
rect 1022 1588 1023 1592
rect 1027 1588 1028 1592
rect 1022 1587 1028 1588
rect 1214 1592 1220 1593
rect 1214 1588 1215 1592
rect 1219 1588 1220 1592
rect 1214 1587 1220 1588
rect 1406 1592 1412 1593
rect 1406 1588 1407 1592
rect 1411 1588 1412 1592
rect 1406 1587 1412 1588
rect 1934 1591 1940 1592
rect 1934 1587 1935 1591
rect 1939 1587 1940 1591
rect 110 1586 116 1587
rect 1934 1586 1940 1587
rect 1974 1560 1980 1561
rect 3798 1560 3804 1561
rect 1974 1556 1975 1560
rect 1979 1556 1980 1560
rect 1974 1555 1980 1556
rect 1994 1559 2000 1560
rect 1994 1555 1995 1559
rect 1999 1555 2000 1559
rect 1994 1554 2000 1555
rect 2162 1559 2168 1560
rect 2162 1555 2163 1559
rect 2167 1555 2168 1559
rect 2162 1554 2168 1555
rect 2370 1559 2376 1560
rect 2370 1555 2371 1559
rect 2375 1555 2376 1559
rect 2370 1554 2376 1555
rect 2586 1559 2592 1560
rect 2586 1555 2587 1559
rect 2591 1555 2592 1559
rect 2586 1554 2592 1555
rect 2802 1559 2808 1560
rect 2802 1555 2803 1559
rect 2807 1555 2808 1559
rect 2802 1554 2808 1555
rect 3018 1559 3024 1560
rect 3018 1555 3019 1559
rect 3023 1555 3024 1559
rect 3018 1554 3024 1555
rect 3234 1559 3240 1560
rect 3234 1555 3235 1559
rect 3239 1555 3240 1559
rect 3234 1554 3240 1555
rect 3450 1559 3456 1560
rect 3450 1555 3451 1559
rect 3455 1555 3456 1559
rect 3450 1554 3456 1555
rect 3650 1559 3656 1560
rect 3650 1555 3651 1559
rect 3655 1555 3656 1559
rect 3798 1556 3799 1560
rect 3803 1556 3804 1560
rect 3798 1555 3804 1556
rect 3650 1554 3656 1555
rect 2022 1544 2028 1545
rect 1974 1543 1980 1544
rect 1974 1539 1975 1543
rect 1979 1539 1980 1543
rect 2022 1540 2023 1544
rect 2027 1540 2028 1544
rect 2022 1539 2028 1540
rect 2190 1544 2196 1545
rect 2190 1540 2191 1544
rect 2195 1540 2196 1544
rect 2190 1539 2196 1540
rect 2398 1544 2404 1545
rect 2398 1540 2399 1544
rect 2403 1540 2404 1544
rect 2398 1539 2404 1540
rect 2614 1544 2620 1545
rect 2614 1540 2615 1544
rect 2619 1540 2620 1544
rect 2614 1539 2620 1540
rect 2830 1544 2836 1545
rect 2830 1540 2831 1544
rect 2835 1540 2836 1544
rect 2830 1539 2836 1540
rect 3046 1544 3052 1545
rect 3046 1540 3047 1544
rect 3051 1540 3052 1544
rect 3046 1539 3052 1540
rect 3262 1544 3268 1545
rect 3262 1540 3263 1544
rect 3267 1540 3268 1544
rect 3262 1539 3268 1540
rect 3478 1544 3484 1545
rect 3478 1540 3479 1544
rect 3483 1540 3484 1544
rect 3478 1539 3484 1540
rect 3678 1544 3684 1545
rect 3678 1540 3679 1544
rect 3683 1540 3684 1544
rect 3678 1539 3684 1540
rect 3798 1543 3804 1544
rect 3798 1539 3799 1543
rect 3803 1539 3804 1543
rect 1974 1538 1980 1539
rect 3798 1538 3804 1539
rect 110 1525 116 1526
rect 1934 1525 1940 1526
rect 110 1521 111 1525
rect 115 1521 116 1525
rect 110 1520 116 1521
rect 358 1524 364 1525
rect 358 1520 359 1524
rect 363 1520 364 1524
rect 358 1519 364 1520
rect 630 1524 636 1525
rect 630 1520 631 1524
rect 635 1520 636 1524
rect 630 1519 636 1520
rect 886 1524 892 1525
rect 886 1520 887 1524
rect 891 1520 892 1524
rect 886 1519 892 1520
rect 1134 1524 1140 1525
rect 1134 1520 1135 1524
rect 1139 1520 1140 1524
rect 1134 1519 1140 1520
rect 1366 1524 1372 1525
rect 1366 1520 1367 1524
rect 1371 1520 1372 1524
rect 1366 1519 1372 1520
rect 1598 1524 1604 1525
rect 1598 1520 1599 1524
rect 1603 1520 1604 1524
rect 1598 1519 1604 1520
rect 1814 1524 1820 1525
rect 1814 1520 1815 1524
rect 1819 1520 1820 1524
rect 1934 1521 1935 1525
rect 1939 1521 1940 1525
rect 1934 1520 1940 1521
rect 3838 1525 3844 1526
rect 5662 1525 5668 1526
rect 3838 1521 3839 1525
rect 3843 1521 3844 1525
rect 3838 1520 3844 1521
rect 3886 1524 3892 1525
rect 3886 1520 3887 1524
rect 3891 1520 3892 1524
rect 1814 1519 1820 1520
rect 3886 1519 3892 1520
rect 4030 1524 4036 1525
rect 4030 1520 4031 1524
rect 4035 1520 4036 1524
rect 4030 1519 4036 1520
rect 4198 1524 4204 1525
rect 4198 1520 4199 1524
rect 4203 1520 4204 1524
rect 4198 1519 4204 1520
rect 4366 1524 4372 1525
rect 4366 1520 4367 1524
rect 4371 1520 4372 1524
rect 4366 1519 4372 1520
rect 4526 1524 4532 1525
rect 4526 1520 4527 1524
rect 4531 1520 4532 1524
rect 4526 1519 4532 1520
rect 4694 1524 4700 1525
rect 4694 1520 4695 1524
rect 4699 1520 4700 1524
rect 4694 1519 4700 1520
rect 4862 1524 4868 1525
rect 4862 1520 4863 1524
rect 4867 1520 4868 1524
rect 4862 1519 4868 1520
rect 5030 1524 5036 1525
rect 5030 1520 5031 1524
rect 5035 1520 5036 1524
rect 5030 1519 5036 1520
rect 5206 1524 5212 1525
rect 5206 1520 5207 1524
rect 5211 1520 5212 1524
rect 5206 1519 5212 1520
rect 5382 1524 5388 1525
rect 5382 1520 5383 1524
rect 5387 1520 5388 1524
rect 5382 1519 5388 1520
rect 5542 1524 5548 1525
rect 5542 1520 5543 1524
rect 5547 1520 5548 1524
rect 5662 1521 5663 1525
rect 5667 1521 5668 1525
rect 5662 1520 5668 1521
rect 5542 1519 5548 1520
rect 330 1509 336 1510
rect 110 1508 116 1509
rect 110 1504 111 1508
rect 115 1504 116 1508
rect 330 1505 331 1509
rect 335 1505 336 1509
rect 330 1504 336 1505
rect 602 1509 608 1510
rect 602 1505 603 1509
rect 607 1505 608 1509
rect 602 1504 608 1505
rect 858 1509 864 1510
rect 858 1505 859 1509
rect 863 1505 864 1509
rect 858 1504 864 1505
rect 1106 1509 1112 1510
rect 1106 1505 1107 1509
rect 1111 1505 1112 1509
rect 1106 1504 1112 1505
rect 1338 1509 1344 1510
rect 1338 1505 1339 1509
rect 1343 1505 1344 1509
rect 1338 1504 1344 1505
rect 1570 1509 1576 1510
rect 1570 1505 1571 1509
rect 1575 1505 1576 1509
rect 1570 1504 1576 1505
rect 1786 1509 1792 1510
rect 3858 1509 3864 1510
rect 1786 1505 1787 1509
rect 1791 1505 1792 1509
rect 1786 1504 1792 1505
rect 1934 1508 1940 1509
rect 1934 1504 1935 1508
rect 1939 1504 1940 1508
rect 110 1503 116 1504
rect 1934 1503 1940 1504
rect 3838 1508 3844 1509
rect 3838 1504 3839 1508
rect 3843 1504 3844 1508
rect 3858 1505 3859 1509
rect 3863 1505 3864 1509
rect 3858 1504 3864 1505
rect 4002 1509 4008 1510
rect 4002 1505 4003 1509
rect 4007 1505 4008 1509
rect 4002 1504 4008 1505
rect 4170 1509 4176 1510
rect 4170 1505 4171 1509
rect 4175 1505 4176 1509
rect 4170 1504 4176 1505
rect 4338 1509 4344 1510
rect 4338 1505 4339 1509
rect 4343 1505 4344 1509
rect 4338 1504 4344 1505
rect 4498 1509 4504 1510
rect 4498 1505 4499 1509
rect 4503 1505 4504 1509
rect 4498 1504 4504 1505
rect 4666 1509 4672 1510
rect 4666 1505 4667 1509
rect 4671 1505 4672 1509
rect 4666 1504 4672 1505
rect 4834 1509 4840 1510
rect 4834 1505 4835 1509
rect 4839 1505 4840 1509
rect 4834 1504 4840 1505
rect 5002 1509 5008 1510
rect 5002 1505 5003 1509
rect 5007 1505 5008 1509
rect 5002 1504 5008 1505
rect 5178 1509 5184 1510
rect 5178 1505 5179 1509
rect 5183 1505 5184 1509
rect 5178 1504 5184 1505
rect 5354 1509 5360 1510
rect 5354 1505 5355 1509
rect 5359 1505 5360 1509
rect 5354 1504 5360 1505
rect 5514 1509 5520 1510
rect 5514 1505 5515 1509
rect 5519 1505 5520 1509
rect 5514 1504 5520 1505
rect 5662 1508 5668 1509
rect 5662 1504 5663 1508
rect 5667 1504 5668 1508
rect 3838 1503 3844 1504
rect 5662 1503 5668 1504
rect 110 1376 116 1377
rect 1934 1376 1940 1377
rect 110 1372 111 1376
rect 115 1372 116 1376
rect 110 1371 116 1372
rect 130 1375 136 1376
rect 130 1371 131 1375
rect 135 1371 136 1375
rect 130 1370 136 1371
rect 306 1375 312 1376
rect 306 1371 307 1375
rect 311 1371 312 1375
rect 306 1370 312 1371
rect 498 1375 504 1376
rect 498 1371 499 1375
rect 503 1371 504 1375
rect 498 1370 504 1371
rect 682 1375 688 1376
rect 682 1371 683 1375
rect 687 1371 688 1375
rect 682 1370 688 1371
rect 858 1375 864 1376
rect 858 1371 859 1375
rect 863 1371 864 1375
rect 858 1370 864 1371
rect 1026 1375 1032 1376
rect 1026 1371 1027 1375
rect 1031 1371 1032 1375
rect 1026 1370 1032 1371
rect 1186 1375 1192 1376
rect 1186 1371 1187 1375
rect 1191 1371 1192 1375
rect 1186 1370 1192 1371
rect 1338 1375 1344 1376
rect 1338 1371 1339 1375
rect 1343 1371 1344 1375
rect 1338 1370 1344 1371
rect 1490 1375 1496 1376
rect 1490 1371 1491 1375
rect 1495 1371 1496 1375
rect 1490 1370 1496 1371
rect 1650 1375 1656 1376
rect 1650 1371 1651 1375
rect 1655 1371 1656 1375
rect 1650 1370 1656 1371
rect 1786 1375 1792 1376
rect 1786 1371 1787 1375
rect 1791 1371 1792 1375
rect 1934 1372 1935 1376
rect 1939 1372 1940 1376
rect 1934 1371 1940 1372
rect 3838 1372 3844 1373
rect 5662 1372 5668 1373
rect 1786 1370 1792 1371
rect 3838 1368 3839 1372
rect 3843 1368 3844 1372
rect 3838 1367 3844 1368
rect 3858 1371 3864 1372
rect 3858 1367 3859 1371
rect 3863 1367 3864 1371
rect 3858 1366 3864 1367
rect 4002 1371 4008 1372
rect 4002 1367 4003 1371
rect 4007 1367 4008 1371
rect 4002 1366 4008 1367
rect 4178 1371 4184 1372
rect 4178 1367 4179 1371
rect 4183 1367 4184 1371
rect 4178 1366 4184 1367
rect 4354 1371 4360 1372
rect 4354 1367 4355 1371
rect 4359 1367 4360 1371
rect 4354 1366 4360 1367
rect 4530 1371 4536 1372
rect 4530 1367 4531 1371
rect 4535 1367 4536 1371
rect 4530 1366 4536 1367
rect 4706 1371 4712 1372
rect 4706 1367 4707 1371
rect 4711 1367 4712 1371
rect 4706 1366 4712 1367
rect 4874 1371 4880 1372
rect 4874 1367 4875 1371
rect 4879 1367 4880 1371
rect 4874 1366 4880 1367
rect 5042 1371 5048 1372
rect 5042 1367 5043 1371
rect 5047 1367 5048 1371
rect 5042 1366 5048 1367
rect 5202 1371 5208 1372
rect 5202 1367 5203 1371
rect 5207 1367 5208 1371
rect 5202 1366 5208 1367
rect 5370 1371 5376 1372
rect 5370 1367 5371 1371
rect 5375 1367 5376 1371
rect 5370 1366 5376 1367
rect 5514 1371 5520 1372
rect 5514 1367 5515 1371
rect 5519 1367 5520 1371
rect 5662 1368 5663 1372
rect 5667 1368 5668 1372
rect 5662 1367 5668 1368
rect 5514 1366 5520 1367
rect 158 1360 164 1361
rect 110 1359 116 1360
rect 110 1355 111 1359
rect 115 1355 116 1359
rect 158 1356 159 1360
rect 163 1356 164 1360
rect 158 1355 164 1356
rect 334 1360 340 1361
rect 334 1356 335 1360
rect 339 1356 340 1360
rect 334 1355 340 1356
rect 526 1360 532 1361
rect 526 1356 527 1360
rect 531 1356 532 1360
rect 526 1355 532 1356
rect 710 1360 716 1361
rect 710 1356 711 1360
rect 715 1356 716 1360
rect 710 1355 716 1356
rect 886 1360 892 1361
rect 886 1356 887 1360
rect 891 1356 892 1360
rect 886 1355 892 1356
rect 1054 1360 1060 1361
rect 1054 1356 1055 1360
rect 1059 1356 1060 1360
rect 1054 1355 1060 1356
rect 1214 1360 1220 1361
rect 1214 1356 1215 1360
rect 1219 1356 1220 1360
rect 1214 1355 1220 1356
rect 1366 1360 1372 1361
rect 1366 1356 1367 1360
rect 1371 1356 1372 1360
rect 1366 1355 1372 1356
rect 1518 1360 1524 1361
rect 1518 1356 1519 1360
rect 1523 1356 1524 1360
rect 1518 1355 1524 1356
rect 1678 1360 1684 1361
rect 1678 1356 1679 1360
rect 1683 1356 1684 1360
rect 1678 1355 1684 1356
rect 1814 1360 1820 1361
rect 1814 1356 1815 1360
rect 1819 1356 1820 1360
rect 1814 1355 1820 1356
rect 1934 1359 1940 1360
rect 1934 1355 1935 1359
rect 1939 1355 1940 1359
rect 3886 1356 3892 1357
rect 110 1354 116 1355
rect 1934 1354 1940 1355
rect 3838 1355 3844 1356
rect 3838 1351 3839 1355
rect 3843 1351 3844 1355
rect 3886 1352 3887 1356
rect 3891 1352 3892 1356
rect 3886 1351 3892 1352
rect 4030 1356 4036 1357
rect 4030 1352 4031 1356
rect 4035 1352 4036 1356
rect 4030 1351 4036 1352
rect 4206 1356 4212 1357
rect 4206 1352 4207 1356
rect 4211 1352 4212 1356
rect 4206 1351 4212 1352
rect 4382 1356 4388 1357
rect 4382 1352 4383 1356
rect 4387 1352 4388 1356
rect 4382 1351 4388 1352
rect 4558 1356 4564 1357
rect 4558 1352 4559 1356
rect 4563 1352 4564 1356
rect 4558 1351 4564 1352
rect 4734 1356 4740 1357
rect 4734 1352 4735 1356
rect 4739 1352 4740 1356
rect 4734 1351 4740 1352
rect 4902 1356 4908 1357
rect 4902 1352 4903 1356
rect 4907 1352 4908 1356
rect 4902 1351 4908 1352
rect 5070 1356 5076 1357
rect 5070 1352 5071 1356
rect 5075 1352 5076 1356
rect 5070 1351 5076 1352
rect 5230 1356 5236 1357
rect 5230 1352 5231 1356
rect 5235 1352 5236 1356
rect 5230 1351 5236 1352
rect 5398 1356 5404 1357
rect 5398 1352 5399 1356
rect 5403 1352 5404 1356
rect 5398 1351 5404 1352
rect 5542 1356 5548 1357
rect 5542 1352 5543 1356
rect 5547 1352 5548 1356
rect 5542 1351 5548 1352
rect 5662 1355 5668 1356
rect 5662 1351 5663 1355
rect 5667 1351 5668 1355
rect 3838 1350 3844 1351
rect 5662 1350 5668 1351
rect 3838 1297 3844 1298
rect 5662 1297 5668 1298
rect 110 1293 116 1294
rect 1934 1293 1940 1294
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 158 1292 164 1293
rect 158 1288 159 1292
rect 163 1288 164 1292
rect 158 1287 164 1288
rect 374 1292 380 1293
rect 374 1288 375 1292
rect 379 1288 380 1292
rect 374 1287 380 1288
rect 598 1292 604 1293
rect 598 1288 599 1292
rect 603 1288 604 1292
rect 598 1287 604 1288
rect 806 1292 812 1293
rect 806 1288 807 1292
rect 811 1288 812 1292
rect 806 1287 812 1288
rect 998 1292 1004 1293
rect 998 1288 999 1292
rect 1003 1288 1004 1292
rect 998 1287 1004 1288
rect 1174 1292 1180 1293
rect 1174 1288 1175 1292
rect 1179 1288 1180 1292
rect 1174 1287 1180 1288
rect 1342 1292 1348 1293
rect 1342 1288 1343 1292
rect 1347 1288 1348 1292
rect 1342 1287 1348 1288
rect 1510 1292 1516 1293
rect 1510 1288 1511 1292
rect 1515 1288 1516 1292
rect 1510 1287 1516 1288
rect 1670 1292 1676 1293
rect 1670 1288 1671 1292
rect 1675 1288 1676 1292
rect 1670 1287 1676 1288
rect 1814 1292 1820 1293
rect 1814 1288 1815 1292
rect 1819 1288 1820 1292
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 3838 1293 3839 1297
rect 3843 1293 3844 1297
rect 3838 1292 3844 1293
rect 3886 1296 3892 1297
rect 3886 1292 3887 1296
rect 3891 1292 3892 1296
rect 3886 1291 3892 1292
rect 4174 1296 4180 1297
rect 4174 1292 4175 1296
rect 4179 1292 4180 1296
rect 4174 1291 4180 1292
rect 4470 1296 4476 1297
rect 4470 1292 4471 1296
rect 4475 1292 4476 1296
rect 4470 1291 4476 1292
rect 4750 1296 4756 1297
rect 4750 1292 4751 1296
rect 4755 1292 4756 1296
rect 4750 1291 4756 1292
rect 5022 1296 5028 1297
rect 5022 1292 5023 1296
rect 5027 1292 5028 1296
rect 5022 1291 5028 1292
rect 5286 1296 5292 1297
rect 5286 1292 5287 1296
rect 5291 1292 5292 1296
rect 5286 1291 5292 1292
rect 5542 1296 5548 1297
rect 5542 1292 5543 1296
rect 5547 1292 5548 1296
rect 5662 1293 5663 1297
rect 5667 1293 5668 1297
rect 5662 1292 5668 1293
rect 5542 1291 5548 1292
rect 1934 1288 1940 1289
rect 1814 1287 1820 1288
rect 1974 1281 1980 1282
rect 3798 1281 3804 1282
rect 3858 1281 3864 1282
rect 130 1277 136 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 130 1273 131 1277
rect 135 1273 136 1277
rect 130 1272 136 1273
rect 346 1277 352 1278
rect 346 1273 347 1277
rect 351 1273 352 1277
rect 346 1272 352 1273
rect 570 1277 576 1278
rect 570 1273 571 1277
rect 575 1273 576 1277
rect 570 1272 576 1273
rect 778 1277 784 1278
rect 778 1273 779 1277
rect 783 1273 784 1277
rect 778 1272 784 1273
rect 970 1277 976 1278
rect 970 1273 971 1277
rect 975 1273 976 1277
rect 970 1272 976 1273
rect 1146 1277 1152 1278
rect 1146 1273 1147 1277
rect 1151 1273 1152 1277
rect 1146 1272 1152 1273
rect 1314 1277 1320 1278
rect 1314 1273 1315 1277
rect 1319 1273 1320 1277
rect 1314 1272 1320 1273
rect 1482 1277 1488 1278
rect 1482 1273 1483 1277
rect 1487 1273 1488 1277
rect 1482 1272 1488 1273
rect 1642 1277 1648 1278
rect 1642 1273 1643 1277
rect 1647 1273 1648 1277
rect 1642 1272 1648 1273
rect 1786 1277 1792 1278
rect 1974 1277 1975 1281
rect 1979 1277 1980 1281
rect 1786 1273 1787 1277
rect 1791 1273 1792 1277
rect 1786 1272 1792 1273
rect 1934 1276 1940 1277
rect 1974 1276 1980 1277
rect 3270 1280 3276 1281
rect 3270 1276 3271 1280
rect 3275 1276 3276 1280
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 3270 1275 3276 1276
rect 3406 1280 3412 1281
rect 3406 1276 3407 1280
rect 3411 1276 3412 1280
rect 3406 1275 3412 1276
rect 3542 1280 3548 1281
rect 3542 1276 3543 1280
rect 3547 1276 3548 1280
rect 3542 1275 3548 1276
rect 3678 1280 3684 1281
rect 3678 1276 3679 1280
rect 3683 1276 3684 1280
rect 3798 1277 3799 1281
rect 3803 1277 3804 1281
rect 3798 1276 3804 1277
rect 3838 1280 3844 1281
rect 3838 1276 3839 1280
rect 3843 1276 3844 1280
rect 3858 1277 3859 1281
rect 3863 1277 3864 1281
rect 3858 1276 3864 1277
rect 4146 1281 4152 1282
rect 4146 1277 4147 1281
rect 4151 1277 4152 1281
rect 4146 1276 4152 1277
rect 4442 1281 4448 1282
rect 4442 1277 4443 1281
rect 4447 1277 4448 1281
rect 4442 1276 4448 1277
rect 4722 1281 4728 1282
rect 4722 1277 4723 1281
rect 4727 1277 4728 1281
rect 4722 1276 4728 1277
rect 4994 1281 5000 1282
rect 4994 1277 4995 1281
rect 4999 1277 5000 1281
rect 4994 1276 5000 1277
rect 5258 1281 5264 1282
rect 5258 1277 5259 1281
rect 5263 1277 5264 1281
rect 5258 1276 5264 1277
rect 5514 1281 5520 1282
rect 5514 1277 5515 1281
rect 5519 1277 5520 1281
rect 5514 1276 5520 1277
rect 5662 1280 5668 1281
rect 5662 1276 5663 1280
rect 5667 1276 5668 1280
rect 3678 1275 3684 1276
rect 3838 1275 3844 1276
rect 5662 1275 5668 1276
rect 110 1271 116 1272
rect 1934 1271 1940 1272
rect 3242 1265 3248 1266
rect 1974 1264 1980 1265
rect 1974 1260 1975 1264
rect 1979 1260 1980 1264
rect 3242 1261 3243 1265
rect 3247 1261 3248 1265
rect 3242 1260 3248 1261
rect 3378 1265 3384 1266
rect 3378 1261 3379 1265
rect 3383 1261 3384 1265
rect 3378 1260 3384 1261
rect 3514 1265 3520 1266
rect 3514 1261 3515 1265
rect 3519 1261 3520 1265
rect 3514 1260 3520 1261
rect 3650 1265 3656 1266
rect 3650 1261 3651 1265
rect 3655 1261 3656 1265
rect 3650 1260 3656 1261
rect 3798 1264 3804 1265
rect 3798 1260 3799 1264
rect 3803 1260 3804 1264
rect 1974 1259 1980 1260
rect 3798 1259 3804 1260
rect 110 1144 116 1145
rect 1934 1144 1940 1145
rect 110 1140 111 1144
rect 115 1140 116 1144
rect 110 1139 116 1140
rect 130 1143 136 1144
rect 130 1139 131 1143
rect 135 1139 136 1143
rect 130 1138 136 1139
rect 346 1143 352 1144
rect 346 1139 347 1143
rect 351 1139 352 1143
rect 346 1138 352 1139
rect 562 1143 568 1144
rect 562 1139 563 1143
rect 567 1139 568 1143
rect 562 1138 568 1139
rect 778 1143 784 1144
rect 778 1139 779 1143
rect 783 1139 784 1143
rect 778 1138 784 1139
rect 986 1143 992 1144
rect 986 1139 987 1143
rect 991 1139 992 1143
rect 986 1138 992 1139
rect 1194 1143 1200 1144
rect 1194 1139 1195 1143
rect 1199 1139 1200 1143
rect 1194 1138 1200 1139
rect 1394 1143 1400 1144
rect 1394 1139 1395 1143
rect 1399 1139 1400 1143
rect 1394 1138 1400 1139
rect 1602 1143 1608 1144
rect 1602 1139 1603 1143
rect 1607 1139 1608 1143
rect 1602 1138 1608 1139
rect 1786 1143 1792 1144
rect 1786 1139 1787 1143
rect 1791 1139 1792 1143
rect 1934 1140 1935 1144
rect 1939 1140 1940 1144
rect 1934 1139 1940 1140
rect 1786 1138 1792 1139
rect 3838 1136 3844 1137
rect 5662 1136 5668 1137
rect 3838 1132 3839 1136
rect 3843 1132 3844 1136
rect 3838 1131 3844 1132
rect 4426 1135 4432 1136
rect 4426 1131 4427 1135
rect 4431 1131 4432 1135
rect 4426 1130 4432 1131
rect 4562 1135 4568 1136
rect 4562 1131 4563 1135
rect 4567 1131 4568 1135
rect 4562 1130 4568 1131
rect 4698 1135 4704 1136
rect 4698 1131 4699 1135
rect 4703 1131 4704 1135
rect 4698 1130 4704 1131
rect 4834 1135 4840 1136
rect 4834 1131 4835 1135
rect 4839 1131 4840 1135
rect 4834 1130 4840 1131
rect 4970 1135 4976 1136
rect 4970 1131 4971 1135
rect 4975 1131 4976 1135
rect 4970 1130 4976 1131
rect 5106 1135 5112 1136
rect 5106 1131 5107 1135
rect 5111 1131 5112 1135
rect 5106 1130 5112 1131
rect 5242 1135 5248 1136
rect 5242 1131 5243 1135
rect 5247 1131 5248 1135
rect 5242 1130 5248 1131
rect 5378 1135 5384 1136
rect 5378 1131 5379 1135
rect 5383 1131 5384 1135
rect 5378 1130 5384 1131
rect 5514 1135 5520 1136
rect 5514 1131 5515 1135
rect 5519 1131 5520 1135
rect 5662 1132 5663 1136
rect 5667 1132 5668 1136
rect 5662 1131 5668 1132
rect 5514 1130 5520 1131
rect 158 1128 164 1129
rect 110 1127 116 1128
rect 110 1123 111 1127
rect 115 1123 116 1127
rect 158 1124 159 1128
rect 163 1124 164 1128
rect 158 1123 164 1124
rect 374 1128 380 1129
rect 374 1124 375 1128
rect 379 1124 380 1128
rect 374 1123 380 1124
rect 590 1128 596 1129
rect 590 1124 591 1128
rect 595 1124 596 1128
rect 590 1123 596 1124
rect 806 1128 812 1129
rect 806 1124 807 1128
rect 811 1124 812 1128
rect 806 1123 812 1124
rect 1014 1128 1020 1129
rect 1014 1124 1015 1128
rect 1019 1124 1020 1128
rect 1014 1123 1020 1124
rect 1222 1128 1228 1129
rect 1222 1124 1223 1128
rect 1227 1124 1228 1128
rect 1222 1123 1228 1124
rect 1422 1128 1428 1129
rect 1422 1124 1423 1128
rect 1427 1124 1428 1128
rect 1422 1123 1428 1124
rect 1630 1128 1636 1129
rect 1630 1124 1631 1128
rect 1635 1124 1636 1128
rect 1630 1123 1636 1124
rect 1814 1128 1820 1129
rect 1814 1124 1815 1128
rect 1819 1124 1820 1128
rect 1814 1123 1820 1124
rect 1934 1127 1940 1128
rect 1934 1123 1935 1127
rect 1939 1123 1940 1127
rect 110 1122 116 1123
rect 1934 1122 1940 1123
rect 1974 1120 1980 1121
rect 3798 1120 3804 1121
rect 4454 1120 4460 1121
rect 1974 1116 1975 1120
rect 1979 1116 1980 1120
rect 1974 1115 1980 1116
rect 1994 1119 2000 1120
rect 1994 1115 1995 1119
rect 1999 1115 2000 1119
rect 1994 1114 2000 1115
rect 2226 1119 2232 1120
rect 2226 1115 2227 1119
rect 2231 1115 2232 1119
rect 2226 1114 2232 1115
rect 2466 1119 2472 1120
rect 2466 1115 2467 1119
rect 2471 1115 2472 1119
rect 2466 1114 2472 1115
rect 2690 1119 2696 1120
rect 2690 1115 2691 1119
rect 2695 1115 2696 1119
rect 2690 1114 2696 1115
rect 2906 1119 2912 1120
rect 2906 1115 2907 1119
rect 2911 1115 2912 1119
rect 2906 1114 2912 1115
rect 3106 1119 3112 1120
rect 3106 1115 3107 1119
rect 3111 1115 3112 1119
rect 3106 1114 3112 1115
rect 3298 1119 3304 1120
rect 3298 1115 3299 1119
rect 3303 1115 3304 1119
rect 3298 1114 3304 1115
rect 3482 1119 3488 1120
rect 3482 1115 3483 1119
rect 3487 1115 3488 1119
rect 3482 1114 3488 1115
rect 3650 1119 3656 1120
rect 3650 1115 3651 1119
rect 3655 1115 3656 1119
rect 3798 1116 3799 1120
rect 3803 1116 3804 1120
rect 3798 1115 3804 1116
rect 3838 1119 3844 1120
rect 3838 1115 3839 1119
rect 3843 1115 3844 1119
rect 4454 1116 4455 1120
rect 4459 1116 4460 1120
rect 4454 1115 4460 1116
rect 4590 1120 4596 1121
rect 4590 1116 4591 1120
rect 4595 1116 4596 1120
rect 4590 1115 4596 1116
rect 4726 1120 4732 1121
rect 4726 1116 4727 1120
rect 4731 1116 4732 1120
rect 4726 1115 4732 1116
rect 4862 1120 4868 1121
rect 4862 1116 4863 1120
rect 4867 1116 4868 1120
rect 4862 1115 4868 1116
rect 4998 1120 5004 1121
rect 4998 1116 4999 1120
rect 5003 1116 5004 1120
rect 4998 1115 5004 1116
rect 5134 1120 5140 1121
rect 5134 1116 5135 1120
rect 5139 1116 5140 1120
rect 5134 1115 5140 1116
rect 5270 1120 5276 1121
rect 5270 1116 5271 1120
rect 5275 1116 5276 1120
rect 5270 1115 5276 1116
rect 5406 1120 5412 1121
rect 5406 1116 5407 1120
rect 5411 1116 5412 1120
rect 5406 1115 5412 1116
rect 5542 1120 5548 1121
rect 5542 1116 5543 1120
rect 5547 1116 5548 1120
rect 5542 1115 5548 1116
rect 5662 1119 5668 1120
rect 5662 1115 5663 1119
rect 5667 1115 5668 1119
rect 3650 1114 3656 1115
rect 3838 1114 3844 1115
rect 5662 1114 5668 1115
rect 2022 1104 2028 1105
rect 1974 1103 1980 1104
rect 1974 1099 1975 1103
rect 1979 1099 1980 1103
rect 2022 1100 2023 1104
rect 2027 1100 2028 1104
rect 2022 1099 2028 1100
rect 2254 1104 2260 1105
rect 2254 1100 2255 1104
rect 2259 1100 2260 1104
rect 2254 1099 2260 1100
rect 2494 1104 2500 1105
rect 2494 1100 2495 1104
rect 2499 1100 2500 1104
rect 2494 1099 2500 1100
rect 2718 1104 2724 1105
rect 2718 1100 2719 1104
rect 2723 1100 2724 1104
rect 2718 1099 2724 1100
rect 2934 1104 2940 1105
rect 2934 1100 2935 1104
rect 2939 1100 2940 1104
rect 2934 1099 2940 1100
rect 3134 1104 3140 1105
rect 3134 1100 3135 1104
rect 3139 1100 3140 1104
rect 3134 1099 3140 1100
rect 3326 1104 3332 1105
rect 3326 1100 3327 1104
rect 3331 1100 3332 1104
rect 3326 1099 3332 1100
rect 3510 1104 3516 1105
rect 3510 1100 3511 1104
rect 3515 1100 3516 1104
rect 3510 1099 3516 1100
rect 3678 1104 3684 1105
rect 3678 1100 3679 1104
rect 3683 1100 3684 1104
rect 3678 1099 3684 1100
rect 3798 1103 3804 1104
rect 3798 1099 3799 1103
rect 3803 1099 3804 1103
rect 1974 1098 1980 1099
rect 3798 1098 3804 1099
rect 110 1045 116 1046
rect 1934 1045 1940 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 470 1044 476 1045
rect 470 1040 471 1044
rect 475 1040 476 1044
rect 470 1039 476 1040
rect 606 1044 612 1045
rect 606 1040 607 1044
rect 611 1040 612 1044
rect 606 1039 612 1040
rect 742 1044 748 1045
rect 742 1040 743 1044
rect 747 1040 748 1044
rect 742 1039 748 1040
rect 886 1044 892 1045
rect 886 1040 887 1044
rect 891 1040 892 1044
rect 886 1039 892 1040
rect 1030 1044 1036 1045
rect 1030 1040 1031 1044
rect 1035 1040 1036 1044
rect 1934 1041 1935 1045
rect 1939 1041 1940 1045
rect 1934 1040 1940 1041
rect 1974 1045 1980 1046
rect 3798 1045 3804 1046
rect 1974 1041 1975 1045
rect 1979 1041 1980 1045
rect 1974 1040 1980 1041
rect 2182 1044 2188 1045
rect 2182 1040 2183 1044
rect 2187 1040 2188 1044
rect 1030 1039 1036 1040
rect 2182 1039 2188 1040
rect 2318 1044 2324 1045
rect 2318 1040 2319 1044
rect 2323 1040 2324 1044
rect 2318 1039 2324 1040
rect 2454 1044 2460 1045
rect 2454 1040 2455 1044
rect 2459 1040 2460 1044
rect 2454 1039 2460 1040
rect 2598 1044 2604 1045
rect 2598 1040 2599 1044
rect 2603 1040 2604 1044
rect 2598 1039 2604 1040
rect 2742 1044 2748 1045
rect 2742 1040 2743 1044
rect 2747 1040 2748 1044
rect 2742 1039 2748 1040
rect 2886 1044 2892 1045
rect 2886 1040 2887 1044
rect 2891 1040 2892 1044
rect 2886 1039 2892 1040
rect 3030 1044 3036 1045
rect 3030 1040 3031 1044
rect 3035 1040 3036 1044
rect 3030 1039 3036 1040
rect 3174 1044 3180 1045
rect 3174 1040 3175 1044
rect 3179 1040 3180 1044
rect 3174 1039 3180 1040
rect 3318 1044 3324 1045
rect 3318 1040 3319 1044
rect 3323 1040 3324 1044
rect 3318 1039 3324 1040
rect 3462 1044 3468 1045
rect 3462 1040 3463 1044
rect 3467 1040 3468 1044
rect 3798 1041 3799 1045
rect 3803 1041 3804 1045
rect 3798 1040 3804 1041
rect 3838 1045 3844 1046
rect 5662 1045 5668 1046
rect 3838 1041 3839 1045
rect 3843 1041 3844 1045
rect 3838 1040 3844 1041
rect 4366 1044 4372 1045
rect 4366 1040 4367 1044
rect 4371 1040 4372 1044
rect 3462 1039 3468 1040
rect 4366 1039 4372 1040
rect 4502 1044 4508 1045
rect 4502 1040 4503 1044
rect 4507 1040 4508 1044
rect 4502 1039 4508 1040
rect 4638 1044 4644 1045
rect 4638 1040 4639 1044
rect 4643 1040 4644 1044
rect 4638 1039 4644 1040
rect 4774 1044 4780 1045
rect 4774 1040 4775 1044
rect 4779 1040 4780 1044
rect 4774 1039 4780 1040
rect 4910 1044 4916 1045
rect 4910 1040 4911 1044
rect 4915 1040 4916 1044
rect 5662 1041 5663 1045
rect 5667 1041 5668 1045
rect 5662 1040 5668 1041
rect 4910 1039 4916 1040
rect 442 1029 448 1030
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 442 1025 443 1029
rect 447 1025 448 1029
rect 442 1024 448 1025
rect 578 1029 584 1030
rect 578 1025 579 1029
rect 583 1025 584 1029
rect 578 1024 584 1025
rect 714 1029 720 1030
rect 714 1025 715 1029
rect 719 1025 720 1029
rect 714 1024 720 1025
rect 858 1029 864 1030
rect 858 1025 859 1029
rect 863 1025 864 1029
rect 858 1024 864 1025
rect 1002 1029 1008 1030
rect 2154 1029 2160 1030
rect 1002 1025 1003 1029
rect 1007 1025 1008 1029
rect 1002 1024 1008 1025
rect 1934 1028 1940 1029
rect 1934 1024 1935 1028
rect 1939 1024 1940 1028
rect 110 1023 116 1024
rect 1934 1023 1940 1024
rect 1974 1028 1980 1029
rect 1974 1024 1975 1028
rect 1979 1024 1980 1028
rect 2154 1025 2155 1029
rect 2159 1025 2160 1029
rect 2154 1024 2160 1025
rect 2290 1029 2296 1030
rect 2290 1025 2291 1029
rect 2295 1025 2296 1029
rect 2290 1024 2296 1025
rect 2426 1029 2432 1030
rect 2426 1025 2427 1029
rect 2431 1025 2432 1029
rect 2426 1024 2432 1025
rect 2570 1029 2576 1030
rect 2570 1025 2571 1029
rect 2575 1025 2576 1029
rect 2570 1024 2576 1025
rect 2714 1029 2720 1030
rect 2714 1025 2715 1029
rect 2719 1025 2720 1029
rect 2714 1024 2720 1025
rect 2858 1029 2864 1030
rect 2858 1025 2859 1029
rect 2863 1025 2864 1029
rect 2858 1024 2864 1025
rect 3002 1029 3008 1030
rect 3002 1025 3003 1029
rect 3007 1025 3008 1029
rect 3002 1024 3008 1025
rect 3146 1029 3152 1030
rect 3146 1025 3147 1029
rect 3151 1025 3152 1029
rect 3146 1024 3152 1025
rect 3290 1029 3296 1030
rect 3290 1025 3291 1029
rect 3295 1025 3296 1029
rect 3290 1024 3296 1025
rect 3434 1029 3440 1030
rect 4338 1029 4344 1030
rect 3434 1025 3435 1029
rect 3439 1025 3440 1029
rect 3434 1024 3440 1025
rect 3798 1028 3804 1029
rect 3798 1024 3799 1028
rect 3803 1024 3804 1028
rect 1974 1023 1980 1024
rect 3798 1023 3804 1024
rect 3838 1028 3844 1029
rect 3838 1024 3839 1028
rect 3843 1024 3844 1028
rect 4338 1025 4339 1029
rect 4343 1025 4344 1029
rect 4338 1024 4344 1025
rect 4474 1029 4480 1030
rect 4474 1025 4475 1029
rect 4479 1025 4480 1029
rect 4474 1024 4480 1025
rect 4610 1029 4616 1030
rect 4610 1025 4611 1029
rect 4615 1025 4616 1029
rect 4610 1024 4616 1025
rect 4746 1029 4752 1030
rect 4746 1025 4747 1029
rect 4751 1025 4752 1029
rect 4746 1024 4752 1025
rect 4882 1029 4888 1030
rect 4882 1025 4883 1029
rect 4887 1025 4888 1029
rect 4882 1024 4888 1025
rect 5662 1028 5668 1029
rect 5662 1024 5663 1028
rect 5667 1024 5668 1028
rect 3838 1023 3844 1024
rect 5662 1023 5668 1024
rect 110 884 116 885
rect 1934 884 1940 885
rect 110 880 111 884
rect 115 880 116 884
rect 110 879 116 880
rect 258 883 264 884
rect 258 879 259 883
rect 263 879 264 883
rect 258 878 264 879
rect 394 883 400 884
rect 394 879 395 883
rect 399 879 400 883
rect 394 878 400 879
rect 530 883 536 884
rect 530 879 531 883
rect 535 879 536 883
rect 530 878 536 879
rect 666 883 672 884
rect 666 879 667 883
rect 671 879 672 883
rect 666 878 672 879
rect 802 883 808 884
rect 802 879 803 883
rect 807 879 808 883
rect 802 878 808 879
rect 938 883 944 884
rect 938 879 939 883
rect 943 879 944 883
rect 1934 880 1935 884
rect 1939 880 1940 884
rect 1934 879 1940 880
rect 1974 884 1980 885
rect 3798 884 3804 885
rect 1974 880 1975 884
rect 1979 880 1980 884
rect 1974 879 1980 880
rect 1994 883 2000 884
rect 1994 879 1995 883
rect 1999 879 2000 883
rect 938 878 944 879
rect 1994 878 2000 879
rect 2130 883 2136 884
rect 2130 879 2131 883
rect 2135 879 2136 883
rect 2130 878 2136 879
rect 2266 883 2272 884
rect 2266 879 2267 883
rect 2271 879 2272 883
rect 2266 878 2272 879
rect 2402 883 2408 884
rect 2402 879 2403 883
rect 2407 879 2408 883
rect 2402 878 2408 879
rect 2538 883 2544 884
rect 2538 879 2539 883
rect 2543 879 2544 883
rect 2538 878 2544 879
rect 2674 883 2680 884
rect 2674 879 2675 883
rect 2679 879 2680 883
rect 2674 878 2680 879
rect 2810 883 2816 884
rect 2810 879 2811 883
rect 2815 879 2816 883
rect 2810 878 2816 879
rect 2946 883 2952 884
rect 2946 879 2947 883
rect 2951 879 2952 883
rect 2946 878 2952 879
rect 3082 883 3088 884
rect 3082 879 3083 883
rect 3087 879 3088 883
rect 3082 878 3088 879
rect 3218 883 3224 884
rect 3218 879 3219 883
rect 3223 879 3224 883
rect 3218 878 3224 879
rect 3354 883 3360 884
rect 3354 879 3355 883
rect 3359 879 3360 883
rect 3354 878 3360 879
rect 3490 883 3496 884
rect 3490 879 3491 883
rect 3495 879 3496 883
rect 3798 880 3799 884
rect 3803 880 3804 884
rect 3798 879 3804 880
rect 3838 884 3844 885
rect 5662 884 5668 885
rect 3838 880 3839 884
rect 3843 880 3844 884
rect 3838 879 3844 880
rect 4018 883 4024 884
rect 4018 879 4019 883
rect 4023 879 4024 883
rect 3490 878 3496 879
rect 4018 878 4024 879
rect 4154 883 4160 884
rect 4154 879 4155 883
rect 4159 879 4160 883
rect 4154 878 4160 879
rect 4290 883 4296 884
rect 4290 879 4291 883
rect 4295 879 4296 883
rect 4290 878 4296 879
rect 4426 883 4432 884
rect 4426 879 4427 883
rect 4431 879 4432 883
rect 4426 878 4432 879
rect 4562 883 4568 884
rect 4562 879 4563 883
rect 4567 879 4568 883
rect 4562 878 4568 879
rect 4698 883 4704 884
rect 4698 879 4699 883
rect 4703 879 4704 883
rect 5662 880 5663 884
rect 5667 880 5668 884
rect 5662 879 5668 880
rect 4698 878 4704 879
rect 286 868 292 869
rect 110 867 116 868
rect 110 863 111 867
rect 115 863 116 867
rect 286 864 287 868
rect 291 864 292 868
rect 286 863 292 864
rect 422 868 428 869
rect 422 864 423 868
rect 427 864 428 868
rect 422 863 428 864
rect 558 868 564 869
rect 558 864 559 868
rect 563 864 564 868
rect 558 863 564 864
rect 694 868 700 869
rect 694 864 695 868
rect 699 864 700 868
rect 694 863 700 864
rect 830 868 836 869
rect 830 864 831 868
rect 835 864 836 868
rect 830 863 836 864
rect 966 868 972 869
rect 2022 868 2028 869
rect 966 864 967 868
rect 971 864 972 868
rect 966 863 972 864
rect 1934 867 1940 868
rect 1934 863 1935 867
rect 1939 863 1940 867
rect 110 862 116 863
rect 1934 862 1940 863
rect 1974 867 1980 868
rect 1974 863 1975 867
rect 1979 863 1980 867
rect 2022 864 2023 868
rect 2027 864 2028 868
rect 2022 863 2028 864
rect 2158 868 2164 869
rect 2158 864 2159 868
rect 2163 864 2164 868
rect 2158 863 2164 864
rect 2294 868 2300 869
rect 2294 864 2295 868
rect 2299 864 2300 868
rect 2294 863 2300 864
rect 2430 868 2436 869
rect 2430 864 2431 868
rect 2435 864 2436 868
rect 2430 863 2436 864
rect 2566 868 2572 869
rect 2566 864 2567 868
rect 2571 864 2572 868
rect 2566 863 2572 864
rect 2702 868 2708 869
rect 2702 864 2703 868
rect 2707 864 2708 868
rect 2702 863 2708 864
rect 2838 868 2844 869
rect 2838 864 2839 868
rect 2843 864 2844 868
rect 2838 863 2844 864
rect 2974 868 2980 869
rect 2974 864 2975 868
rect 2979 864 2980 868
rect 2974 863 2980 864
rect 3110 868 3116 869
rect 3110 864 3111 868
rect 3115 864 3116 868
rect 3110 863 3116 864
rect 3246 868 3252 869
rect 3246 864 3247 868
rect 3251 864 3252 868
rect 3246 863 3252 864
rect 3382 868 3388 869
rect 3382 864 3383 868
rect 3387 864 3388 868
rect 3382 863 3388 864
rect 3518 868 3524 869
rect 4046 868 4052 869
rect 3518 864 3519 868
rect 3523 864 3524 868
rect 3518 863 3524 864
rect 3798 867 3804 868
rect 3798 863 3799 867
rect 3803 863 3804 867
rect 1974 862 1980 863
rect 3798 862 3804 863
rect 3838 867 3844 868
rect 3838 863 3839 867
rect 3843 863 3844 867
rect 4046 864 4047 868
rect 4051 864 4052 868
rect 4046 863 4052 864
rect 4182 868 4188 869
rect 4182 864 4183 868
rect 4187 864 4188 868
rect 4182 863 4188 864
rect 4318 868 4324 869
rect 4318 864 4319 868
rect 4323 864 4324 868
rect 4318 863 4324 864
rect 4454 868 4460 869
rect 4454 864 4455 868
rect 4459 864 4460 868
rect 4454 863 4460 864
rect 4590 868 4596 869
rect 4590 864 4591 868
rect 4595 864 4596 868
rect 4590 863 4596 864
rect 4726 868 4732 869
rect 4726 864 4727 868
rect 4731 864 4732 868
rect 4726 863 4732 864
rect 5662 867 5668 868
rect 5662 863 5663 867
rect 5667 863 5668 867
rect 3838 862 3844 863
rect 5662 862 5668 863
rect 1974 809 1980 810
rect 3798 809 3804 810
rect 1974 805 1975 809
rect 1979 805 1980 809
rect 1974 804 1980 805
rect 2022 808 2028 809
rect 2022 804 2023 808
rect 2027 804 2028 808
rect 2022 803 2028 804
rect 2166 808 2172 809
rect 2166 804 2167 808
rect 2171 804 2172 808
rect 2166 803 2172 804
rect 2334 808 2340 809
rect 2334 804 2335 808
rect 2339 804 2340 808
rect 2334 803 2340 804
rect 2494 808 2500 809
rect 2494 804 2495 808
rect 2499 804 2500 808
rect 2494 803 2500 804
rect 2654 808 2660 809
rect 2654 804 2655 808
rect 2659 804 2660 808
rect 2654 803 2660 804
rect 2822 808 2828 809
rect 2822 804 2823 808
rect 2827 804 2828 808
rect 2822 803 2828 804
rect 2990 808 2996 809
rect 2990 804 2991 808
rect 2995 804 2996 808
rect 3798 805 3799 809
rect 3803 805 3804 809
rect 3798 804 3804 805
rect 2990 803 2996 804
rect 110 797 116 798
rect 1934 797 1940 798
rect 110 793 111 797
rect 115 793 116 797
rect 110 792 116 793
rect 238 796 244 797
rect 238 792 239 796
rect 243 792 244 796
rect 238 791 244 792
rect 438 796 444 797
rect 438 792 439 796
rect 443 792 444 796
rect 438 791 444 792
rect 646 796 652 797
rect 646 792 647 796
rect 651 792 652 796
rect 646 791 652 792
rect 854 796 860 797
rect 854 792 855 796
rect 859 792 860 796
rect 854 791 860 792
rect 1062 796 1068 797
rect 1062 792 1063 796
rect 1067 792 1068 796
rect 1934 793 1935 797
rect 1939 793 1940 797
rect 1994 793 2000 794
rect 1934 792 1940 793
rect 1974 792 1980 793
rect 1062 791 1068 792
rect 1974 788 1975 792
rect 1979 788 1980 792
rect 1994 789 1995 793
rect 1999 789 2000 793
rect 1994 788 2000 789
rect 2138 793 2144 794
rect 2138 789 2139 793
rect 2143 789 2144 793
rect 2138 788 2144 789
rect 2306 793 2312 794
rect 2306 789 2307 793
rect 2311 789 2312 793
rect 2306 788 2312 789
rect 2466 793 2472 794
rect 2466 789 2467 793
rect 2471 789 2472 793
rect 2466 788 2472 789
rect 2626 793 2632 794
rect 2626 789 2627 793
rect 2631 789 2632 793
rect 2626 788 2632 789
rect 2794 793 2800 794
rect 2794 789 2795 793
rect 2799 789 2800 793
rect 2794 788 2800 789
rect 2962 793 2968 794
rect 3838 793 3844 794
rect 5662 793 5668 794
rect 2962 789 2963 793
rect 2967 789 2968 793
rect 2962 788 2968 789
rect 3798 792 3804 793
rect 3798 788 3799 792
rect 3803 788 3804 792
rect 3838 789 3839 793
rect 3843 789 3844 793
rect 3838 788 3844 789
rect 3886 792 3892 793
rect 3886 788 3887 792
rect 3891 788 3892 792
rect 1974 787 1980 788
rect 3798 787 3804 788
rect 3886 787 3892 788
rect 4022 792 4028 793
rect 4022 788 4023 792
rect 4027 788 4028 792
rect 4022 787 4028 788
rect 4158 792 4164 793
rect 4158 788 4159 792
rect 4163 788 4164 792
rect 4158 787 4164 788
rect 4294 792 4300 793
rect 4294 788 4295 792
rect 4299 788 4300 792
rect 4294 787 4300 788
rect 4430 792 4436 793
rect 4430 788 4431 792
rect 4435 788 4436 792
rect 4430 787 4436 788
rect 4566 792 4572 793
rect 4566 788 4567 792
rect 4571 788 4572 792
rect 4566 787 4572 788
rect 4702 792 4708 793
rect 4702 788 4703 792
rect 4707 788 4708 792
rect 4702 787 4708 788
rect 4838 792 4844 793
rect 4838 788 4839 792
rect 4843 788 4844 792
rect 5662 789 5663 793
rect 5667 789 5668 793
rect 5662 788 5668 789
rect 4838 787 4844 788
rect 210 781 216 782
rect 110 780 116 781
rect 110 776 111 780
rect 115 776 116 780
rect 210 777 211 781
rect 215 777 216 781
rect 210 776 216 777
rect 410 781 416 782
rect 410 777 411 781
rect 415 777 416 781
rect 410 776 416 777
rect 618 781 624 782
rect 618 777 619 781
rect 623 777 624 781
rect 618 776 624 777
rect 826 781 832 782
rect 826 777 827 781
rect 831 777 832 781
rect 826 776 832 777
rect 1034 781 1040 782
rect 1034 777 1035 781
rect 1039 777 1040 781
rect 1034 776 1040 777
rect 1934 780 1940 781
rect 1934 776 1935 780
rect 1939 776 1940 780
rect 3858 777 3864 778
rect 110 775 116 776
rect 1934 775 1940 776
rect 3838 776 3844 777
rect 3838 772 3839 776
rect 3843 772 3844 776
rect 3858 773 3859 777
rect 3863 773 3864 777
rect 3858 772 3864 773
rect 3994 777 4000 778
rect 3994 773 3995 777
rect 3999 773 4000 777
rect 3994 772 4000 773
rect 4130 777 4136 778
rect 4130 773 4131 777
rect 4135 773 4136 777
rect 4130 772 4136 773
rect 4266 777 4272 778
rect 4266 773 4267 777
rect 4271 773 4272 777
rect 4266 772 4272 773
rect 4402 777 4408 778
rect 4402 773 4403 777
rect 4407 773 4408 777
rect 4402 772 4408 773
rect 4538 777 4544 778
rect 4538 773 4539 777
rect 4543 773 4544 777
rect 4538 772 4544 773
rect 4674 777 4680 778
rect 4674 773 4675 777
rect 4679 773 4680 777
rect 4674 772 4680 773
rect 4810 777 4816 778
rect 4810 773 4811 777
rect 4815 773 4816 777
rect 4810 772 4816 773
rect 5662 776 5668 777
rect 5662 772 5663 776
rect 5667 772 5668 776
rect 3838 771 3844 772
rect 5662 771 5668 772
rect 3838 644 3844 645
rect 5662 644 5668 645
rect 3838 640 3839 644
rect 3843 640 3844 644
rect 3838 639 3844 640
rect 3858 643 3864 644
rect 3858 639 3859 643
rect 3863 639 3864 643
rect 3858 638 3864 639
rect 3994 643 4000 644
rect 3994 639 3995 643
rect 3999 639 4000 643
rect 3994 638 4000 639
rect 4130 643 4136 644
rect 4130 639 4131 643
rect 4135 639 4136 643
rect 4130 638 4136 639
rect 4266 643 4272 644
rect 4266 639 4267 643
rect 4271 639 4272 643
rect 4266 638 4272 639
rect 4402 643 4408 644
rect 4402 639 4403 643
rect 4407 639 4408 643
rect 4402 638 4408 639
rect 4538 643 4544 644
rect 4538 639 4539 643
rect 4543 639 4544 643
rect 4538 638 4544 639
rect 4674 643 4680 644
rect 4674 639 4675 643
rect 4679 639 4680 643
rect 4674 638 4680 639
rect 4810 643 4816 644
rect 4810 639 4811 643
rect 4815 639 4816 643
rect 4810 638 4816 639
rect 4946 643 4952 644
rect 4946 639 4947 643
rect 4951 639 4952 643
rect 4946 638 4952 639
rect 5082 643 5088 644
rect 5082 639 5083 643
rect 5087 639 5088 643
rect 5662 640 5663 644
rect 5667 640 5668 644
rect 5662 639 5668 640
rect 5082 638 5088 639
rect 1974 632 1980 633
rect 3798 632 3804 633
rect 110 628 116 629
rect 1934 628 1940 629
rect 110 624 111 628
rect 115 624 116 628
rect 110 623 116 624
rect 130 627 136 628
rect 130 623 131 627
rect 135 623 136 627
rect 130 622 136 623
rect 346 627 352 628
rect 346 623 347 627
rect 351 623 352 627
rect 346 622 352 623
rect 586 627 592 628
rect 586 623 587 627
rect 591 623 592 627
rect 586 622 592 623
rect 826 627 832 628
rect 826 623 827 627
rect 831 623 832 627
rect 826 622 832 623
rect 1066 627 1072 628
rect 1066 623 1067 627
rect 1071 623 1072 627
rect 1066 622 1072 623
rect 1314 627 1320 628
rect 1314 623 1315 627
rect 1319 623 1320 627
rect 1314 622 1320 623
rect 1562 627 1568 628
rect 1562 623 1563 627
rect 1567 623 1568 627
rect 1562 622 1568 623
rect 1786 627 1792 628
rect 1786 623 1787 627
rect 1791 623 1792 627
rect 1934 624 1935 628
rect 1939 624 1940 628
rect 1974 628 1975 632
rect 1979 628 1980 632
rect 1974 627 1980 628
rect 1994 631 2000 632
rect 1994 627 1995 631
rect 1999 627 2000 631
rect 1994 626 2000 627
rect 2298 631 2304 632
rect 2298 627 2299 631
rect 2303 627 2304 631
rect 2298 626 2304 627
rect 2634 631 2640 632
rect 2634 627 2635 631
rect 2639 627 2640 631
rect 2634 626 2640 627
rect 2978 631 2984 632
rect 2978 627 2979 631
rect 2983 627 2984 631
rect 2978 626 2984 627
rect 3322 631 3328 632
rect 3322 627 3323 631
rect 3327 627 3328 631
rect 3322 626 3328 627
rect 3650 631 3656 632
rect 3650 627 3651 631
rect 3655 627 3656 631
rect 3798 628 3799 632
rect 3803 628 3804 632
rect 3886 628 3892 629
rect 3798 627 3804 628
rect 3838 627 3844 628
rect 3650 626 3656 627
rect 1934 623 1940 624
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3886 624 3887 628
rect 3891 624 3892 628
rect 3886 623 3892 624
rect 4022 628 4028 629
rect 4022 624 4023 628
rect 4027 624 4028 628
rect 4022 623 4028 624
rect 4158 628 4164 629
rect 4158 624 4159 628
rect 4163 624 4164 628
rect 4158 623 4164 624
rect 4294 628 4300 629
rect 4294 624 4295 628
rect 4299 624 4300 628
rect 4294 623 4300 624
rect 4430 628 4436 629
rect 4430 624 4431 628
rect 4435 624 4436 628
rect 4430 623 4436 624
rect 4566 628 4572 629
rect 4566 624 4567 628
rect 4571 624 4572 628
rect 4566 623 4572 624
rect 4702 628 4708 629
rect 4702 624 4703 628
rect 4707 624 4708 628
rect 4702 623 4708 624
rect 4838 628 4844 629
rect 4838 624 4839 628
rect 4843 624 4844 628
rect 4838 623 4844 624
rect 4974 628 4980 629
rect 4974 624 4975 628
rect 4979 624 4980 628
rect 4974 623 4980 624
rect 5110 628 5116 629
rect 5110 624 5111 628
rect 5115 624 5116 628
rect 5110 623 5116 624
rect 5662 627 5668 628
rect 5662 623 5663 627
rect 5667 623 5668 627
rect 1786 622 1792 623
rect 3838 622 3844 623
rect 5662 622 5668 623
rect 2022 616 2028 617
rect 1974 615 1980 616
rect 158 612 164 613
rect 110 611 116 612
rect 110 607 111 611
rect 115 607 116 611
rect 158 608 159 612
rect 163 608 164 612
rect 158 607 164 608
rect 374 612 380 613
rect 374 608 375 612
rect 379 608 380 612
rect 374 607 380 608
rect 614 612 620 613
rect 614 608 615 612
rect 619 608 620 612
rect 614 607 620 608
rect 854 612 860 613
rect 854 608 855 612
rect 859 608 860 612
rect 854 607 860 608
rect 1094 612 1100 613
rect 1094 608 1095 612
rect 1099 608 1100 612
rect 1094 607 1100 608
rect 1342 612 1348 613
rect 1342 608 1343 612
rect 1347 608 1348 612
rect 1342 607 1348 608
rect 1590 612 1596 613
rect 1590 608 1591 612
rect 1595 608 1596 612
rect 1590 607 1596 608
rect 1814 612 1820 613
rect 1814 608 1815 612
rect 1819 608 1820 612
rect 1814 607 1820 608
rect 1934 611 1940 612
rect 1934 607 1935 611
rect 1939 607 1940 611
rect 1974 611 1975 615
rect 1979 611 1980 615
rect 2022 612 2023 616
rect 2027 612 2028 616
rect 2022 611 2028 612
rect 2326 616 2332 617
rect 2326 612 2327 616
rect 2331 612 2332 616
rect 2326 611 2332 612
rect 2662 616 2668 617
rect 2662 612 2663 616
rect 2667 612 2668 616
rect 2662 611 2668 612
rect 3006 616 3012 617
rect 3006 612 3007 616
rect 3011 612 3012 616
rect 3006 611 3012 612
rect 3350 616 3356 617
rect 3350 612 3351 616
rect 3355 612 3356 616
rect 3350 611 3356 612
rect 3678 616 3684 617
rect 3678 612 3679 616
rect 3683 612 3684 616
rect 3678 611 3684 612
rect 3798 615 3804 616
rect 3798 611 3799 615
rect 3803 611 3804 615
rect 1974 610 1980 611
rect 3798 610 3804 611
rect 110 606 116 607
rect 1934 606 1940 607
rect 1974 557 1980 558
rect 3798 557 3804 558
rect 1974 553 1975 557
rect 1979 553 1980 557
rect 1974 552 1980 553
rect 2334 556 2340 557
rect 2334 552 2335 556
rect 2339 552 2340 556
rect 2334 551 2340 552
rect 2526 556 2532 557
rect 2526 552 2527 556
rect 2531 552 2532 556
rect 2526 551 2532 552
rect 2710 556 2716 557
rect 2710 552 2711 556
rect 2715 552 2716 556
rect 2710 551 2716 552
rect 2886 556 2892 557
rect 2886 552 2887 556
rect 2891 552 2892 556
rect 2886 551 2892 552
rect 3062 556 3068 557
rect 3062 552 3063 556
rect 3067 552 3068 556
rect 3062 551 3068 552
rect 3230 556 3236 557
rect 3230 552 3231 556
rect 3235 552 3236 556
rect 3230 551 3236 552
rect 3406 556 3412 557
rect 3406 552 3407 556
rect 3411 552 3412 556
rect 3406 551 3412 552
rect 3582 556 3588 557
rect 3582 552 3583 556
rect 3587 552 3588 556
rect 3798 553 3799 557
rect 3803 553 3804 557
rect 3798 552 3804 553
rect 3582 551 3588 552
rect 110 549 116 550
rect 1934 549 1940 550
rect 110 545 111 549
rect 115 545 116 549
rect 110 544 116 545
rect 158 548 164 549
rect 158 544 159 548
rect 163 544 164 548
rect 158 543 164 544
rect 406 548 412 549
rect 406 544 407 548
rect 411 544 412 548
rect 406 543 412 544
rect 670 548 676 549
rect 670 544 671 548
rect 675 544 676 548
rect 670 543 676 544
rect 934 548 940 549
rect 934 544 935 548
rect 939 544 940 548
rect 934 543 940 544
rect 1190 548 1196 549
rect 1190 544 1191 548
rect 1195 544 1196 548
rect 1190 543 1196 544
rect 1446 548 1452 549
rect 1446 544 1447 548
rect 1451 544 1452 548
rect 1446 543 1452 544
rect 1710 548 1716 549
rect 1710 544 1711 548
rect 1715 544 1716 548
rect 1934 545 1935 549
rect 1939 545 1940 549
rect 1934 544 1940 545
rect 3838 549 3844 550
rect 5662 549 5668 550
rect 3838 545 3839 549
rect 3843 545 3844 549
rect 3838 544 3844 545
rect 4046 548 4052 549
rect 4046 544 4047 548
rect 4051 544 4052 548
rect 1710 543 1716 544
rect 4046 543 4052 544
rect 4206 548 4212 549
rect 4206 544 4207 548
rect 4211 544 4212 548
rect 4206 543 4212 544
rect 4366 548 4372 549
rect 4366 544 4367 548
rect 4371 544 4372 548
rect 4366 543 4372 544
rect 4526 548 4532 549
rect 4526 544 4527 548
rect 4531 544 4532 548
rect 4526 543 4532 544
rect 4686 548 4692 549
rect 4686 544 4687 548
rect 4691 544 4692 548
rect 5662 545 5663 549
rect 5667 545 5668 549
rect 5662 544 5668 545
rect 4686 543 4692 544
rect 2306 541 2312 542
rect 1974 540 1980 541
rect 1974 536 1975 540
rect 1979 536 1980 540
rect 2306 537 2307 541
rect 2311 537 2312 541
rect 2306 536 2312 537
rect 2498 541 2504 542
rect 2498 537 2499 541
rect 2503 537 2504 541
rect 2498 536 2504 537
rect 2682 541 2688 542
rect 2682 537 2683 541
rect 2687 537 2688 541
rect 2682 536 2688 537
rect 2858 541 2864 542
rect 2858 537 2859 541
rect 2863 537 2864 541
rect 2858 536 2864 537
rect 3034 541 3040 542
rect 3034 537 3035 541
rect 3039 537 3040 541
rect 3034 536 3040 537
rect 3202 541 3208 542
rect 3202 537 3203 541
rect 3207 537 3208 541
rect 3202 536 3208 537
rect 3378 541 3384 542
rect 3378 537 3379 541
rect 3383 537 3384 541
rect 3378 536 3384 537
rect 3554 541 3560 542
rect 3554 537 3555 541
rect 3559 537 3560 541
rect 3554 536 3560 537
rect 3798 540 3804 541
rect 3798 536 3799 540
rect 3803 536 3804 540
rect 1974 535 1980 536
rect 3798 535 3804 536
rect 130 533 136 534
rect 110 532 116 533
rect 110 528 111 532
rect 115 528 116 532
rect 130 529 131 533
rect 135 529 136 533
rect 130 528 136 529
rect 378 533 384 534
rect 378 529 379 533
rect 383 529 384 533
rect 378 528 384 529
rect 642 533 648 534
rect 642 529 643 533
rect 647 529 648 533
rect 642 528 648 529
rect 906 533 912 534
rect 906 529 907 533
rect 911 529 912 533
rect 906 528 912 529
rect 1162 533 1168 534
rect 1162 529 1163 533
rect 1167 529 1168 533
rect 1162 528 1168 529
rect 1418 533 1424 534
rect 1418 529 1419 533
rect 1423 529 1424 533
rect 1418 528 1424 529
rect 1682 533 1688 534
rect 4018 533 4024 534
rect 1682 529 1683 533
rect 1687 529 1688 533
rect 1682 528 1688 529
rect 1934 532 1940 533
rect 1934 528 1935 532
rect 1939 528 1940 532
rect 110 527 116 528
rect 1934 527 1940 528
rect 3838 532 3844 533
rect 3838 528 3839 532
rect 3843 528 3844 532
rect 4018 529 4019 533
rect 4023 529 4024 533
rect 4018 528 4024 529
rect 4178 533 4184 534
rect 4178 529 4179 533
rect 4183 529 4184 533
rect 4178 528 4184 529
rect 4338 533 4344 534
rect 4338 529 4339 533
rect 4343 529 4344 533
rect 4338 528 4344 529
rect 4498 533 4504 534
rect 4498 529 4499 533
rect 4503 529 4504 533
rect 4498 528 4504 529
rect 4658 533 4664 534
rect 4658 529 4659 533
rect 4663 529 4664 533
rect 4658 528 4664 529
rect 5662 532 5668 533
rect 5662 528 5663 532
rect 5667 528 5668 532
rect 3838 527 3844 528
rect 5662 527 5668 528
rect 1974 408 1980 409
rect 3798 408 3804 409
rect 1974 404 1975 408
rect 1979 404 1980 408
rect 1974 403 1980 404
rect 2170 407 2176 408
rect 2170 403 2171 407
rect 2175 403 2176 407
rect 2170 402 2176 403
rect 2314 407 2320 408
rect 2314 403 2315 407
rect 2319 403 2320 407
rect 2314 402 2320 403
rect 2458 407 2464 408
rect 2458 403 2459 407
rect 2463 403 2464 407
rect 2458 402 2464 403
rect 2602 407 2608 408
rect 2602 403 2603 407
rect 2607 403 2608 407
rect 2602 402 2608 403
rect 2746 407 2752 408
rect 2746 403 2747 407
rect 2751 403 2752 407
rect 2746 402 2752 403
rect 2890 407 2896 408
rect 2890 403 2891 407
rect 2895 403 2896 407
rect 2890 402 2896 403
rect 3034 407 3040 408
rect 3034 403 3035 407
rect 3039 403 3040 407
rect 3798 404 3799 408
rect 3803 404 3804 408
rect 3798 403 3804 404
rect 3034 402 3040 403
rect 110 400 116 401
rect 1934 400 1940 401
rect 110 396 111 400
rect 115 396 116 400
rect 110 395 116 396
rect 194 399 200 400
rect 194 395 195 399
rect 199 395 200 399
rect 194 394 200 395
rect 426 399 432 400
rect 426 395 427 399
rect 431 395 432 399
rect 426 394 432 395
rect 658 399 664 400
rect 658 395 659 399
rect 663 395 664 399
rect 658 394 664 395
rect 882 399 888 400
rect 882 395 883 399
rect 887 395 888 399
rect 882 394 888 395
rect 1098 399 1104 400
rect 1098 395 1099 399
rect 1103 395 1104 399
rect 1098 394 1104 395
rect 1322 399 1328 400
rect 1322 395 1323 399
rect 1327 395 1328 399
rect 1322 394 1328 395
rect 1546 399 1552 400
rect 1546 395 1547 399
rect 1551 395 1552 399
rect 1934 396 1935 400
rect 1939 396 1940 400
rect 1934 395 1940 396
rect 1546 394 1552 395
rect 2198 392 2204 393
rect 1974 391 1980 392
rect 1974 387 1975 391
rect 1979 387 1980 391
rect 2198 388 2199 392
rect 2203 388 2204 392
rect 2198 387 2204 388
rect 2342 392 2348 393
rect 2342 388 2343 392
rect 2347 388 2348 392
rect 2342 387 2348 388
rect 2486 392 2492 393
rect 2486 388 2487 392
rect 2491 388 2492 392
rect 2486 387 2492 388
rect 2630 392 2636 393
rect 2630 388 2631 392
rect 2635 388 2636 392
rect 2630 387 2636 388
rect 2774 392 2780 393
rect 2774 388 2775 392
rect 2779 388 2780 392
rect 2774 387 2780 388
rect 2918 392 2924 393
rect 2918 388 2919 392
rect 2923 388 2924 392
rect 2918 387 2924 388
rect 3062 392 3068 393
rect 3838 392 3844 393
rect 5662 392 5668 393
rect 3062 388 3063 392
rect 3067 388 3068 392
rect 3062 387 3068 388
rect 3798 391 3804 392
rect 3798 387 3799 391
rect 3803 387 3804 391
rect 3838 388 3839 392
rect 3843 388 3844 392
rect 3838 387 3844 388
rect 3930 391 3936 392
rect 3930 387 3931 391
rect 3935 387 3936 391
rect 1974 386 1980 387
rect 3798 386 3804 387
rect 3930 386 3936 387
rect 4130 391 4136 392
rect 4130 387 4131 391
rect 4135 387 4136 391
rect 4130 386 4136 387
rect 4330 391 4336 392
rect 4330 387 4331 391
rect 4335 387 4336 391
rect 4330 386 4336 387
rect 4522 391 4528 392
rect 4522 387 4523 391
rect 4527 387 4528 391
rect 4522 386 4528 387
rect 4722 391 4728 392
rect 4722 387 4723 391
rect 4727 387 4728 391
rect 4722 386 4728 387
rect 4922 391 4928 392
rect 4922 387 4923 391
rect 4927 387 4928 391
rect 5662 388 5663 392
rect 5667 388 5668 392
rect 5662 387 5668 388
rect 4922 386 4928 387
rect 222 384 228 385
rect 110 383 116 384
rect 110 379 111 383
rect 115 379 116 383
rect 222 380 223 384
rect 227 380 228 384
rect 222 379 228 380
rect 454 384 460 385
rect 454 380 455 384
rect 459 380 460 384
rect 454 379 460 380
rect 686 384 692 385
rect 686 380 687 384
rect 691 380 692 384
rect 686 379 692 380
rect 910 384 916 385
rect 910 380 911 384
rect 915 380 916 384
rect 910 379 916 380
rect 1126 384 1132 385
rect 1126 380 1127 384
rect 1131 380 1132 384
rect 1126 379 1132 380
rect 1350 384 1356 385
rect 1350 380 1351 384
rect 1355 380 1356 384
rect 1350 379 1356 380
rect 1574 384 1580 385
rect 1574 380 1575 384
rect 1579 380 1580 384
rect 1574 379 1580 380
rect 1934 383 1940 384
rect 1934 379 1935 383
rect 1939 379 1940 383
rect 110 378 116 379
rect 1934 378 1940 379
rect 3958 376 3964 377
rect 3838 375 3844 376
rect 3838 371 3839 375
rect 3843 371 3844 375
rect 3958 372 3959 376
rect 3963 372 3964 376
rect 3958 371 3964 372
rect 4158 376 4164 377
rect 4158 372 4159 376
rect 4163 372 4164 376
rect 4158 371 4164 372
rect 4358 376 4364 377
rect 4358 372 4359 376
rect 4363 372 4364 376
rect 4358 371 4364 372
rect 4550 376 4556 377
rect 4550 372 4551 376
rect 4555 372 4556 376
rect 4550 371 4556 372
rect 4750 376 4756 377
rect 4750 372 4751 376
rect 4755 372 4756 376
rect 4750 371 4756 372
rect 4950 376 4956 377
rect 4950 372 4951 376
rect 4955 372 4956 376
rect 4950 371 4956 372
rect 5662 375 5668 376
rect 5662 371 5663 375
rect 5667 371 5668 375
rect 3838 370 3844 371
rect 5662 370 5668 371
rect 1974 329 1980 330
rect 3798 329 3804 330
rect 1974 325 1975 329
rect 1979 325 1980 329
rect 1974 324 1980 325
rect 2022 328 2028 329
rect 2022 324 2023 328
rect 2027 324 2028 328
rect 2022 323 2028 324
rect 2174 328 2180 329
rect 2174 324 2175 328
rect 2179 324 2180 328
rect 2174 323 2180 324
rect 2366 328 2372 329
rect 2366 324 2367 328
rect 2371 324 2372 328
rect 2366 323 2372 324
rect 2590 328 2596 329
rect 2590 324 2591 328
rect 2595 324 2596 328
rect 2590 323 2596 324
rect 2846 328 2852 329
rect 2846 324 2847 328
rect 2851 324 2852 328
rect 2846 323 2852 324
rect 3118 328 3124 329
rect 3118 324 3119 328
rect 3123 324 3124 328
rect 3118 323 3124 324
rect 3406 328 3412 329
rect 3406 324 3407 328
rect 3411 324 3412 328
rect 3406 323 3412 324
rect 3678 328 3684 329
rect 3678 324 3679 328
rect 3683 324 3684 328
rect 3798 325 3799 329
rect 3803 325 3804 329
rect 3798 324 3804 325
rect 3678 323 3684 324
rect 110 317 116 318
rect 1934 317 1940 318
rect 110 313 111 317
rect 115 313 116 317
rect 110 312 116 313
rect 350 316 356 317
rect 350 312 351 316
rect 355 312 356 316
rect 350 311 356 312
rect 574 316 580 317
rect 574 312 575 316
rect 579 312 580 316
rect 574 311 580 312
rect 798 316 804 317
rect 798 312 799 316
rect 803 312 804 316
rect 798 311 804 312
rect 1014 316 1020 317
rect 1014 312 1015 316
rect 1019 312 1020 316
rect 1014 311 1020 312
rect 1230 316 1236 317
rect 1230 312 1231 316
rect 1235 312 1236 316
rect 1230 311 1236 312
rect 1454 316 1460 317
rect 1454 312 1455 316
rect 1459 312 1460 316
rect 1934 313 1935 317
rect 1939 313 1940 317
rect 3838 317 3844 318
rect 5662 317 5668 318
rect 1994 313 2000 314
rect 1934 312 1940 313
rect 1974 312 1980 313
rect 1454 311 1460 312
rect 1974 308 1975 312
rect 1979 308 1980 312
rect 1994 309 1995 313
rect 1999 309 2000 313
rect 1994 308 2000 309
rect 2146 313 2152 314
rect 2146 309 2147 313
rect 2151 309 2152 313
rect 2146 308 2152 309
rect 2338 313 2344 314
rect 2338 309 2339 313
rect 2343 309 2344 313
rect 2338 308 2344 309
rect 2562 313 2568 314
rect 2562 309 2563 313
rect 2567 309 2568 313
rect 2562 308 2568 309
rect 2818 313 2824 314
rect 2818 309 2819 313
rect 2823 309 2824 313
rect 2818 308 2824 309
rect 3090 313 3096 314
rect 3090 309 3091 313
rect 3095 309 3096 313
rect 3090 308 3096 309
rect 3378 313 3384 314
rect 3378 309 3379 313
rect 3383 309 3384 313
rect 3378 308 3384 309
rect 3650 313 3656 314
rect 3838 313 3839 317
rect 3843 313 3844 317
rect 3650 309 3651 313
rect 3655 309 3656 313
rect 3650 308 3656 309
rect 3798 312 3804 313
rect 3838 312 3844 313
rect 3886 316 3892 317
rect 3886 312 3887 316
rect 3891 312 3892 316
rect 3798 308 3799 312
rect 3803 308 3804 312
rect 3886 311 3892 312
rect 4134 316 4140 317
rect 4134 312 4135 316
rect 4139 312 4140 316
rect 4134 311 4140 312
rect 4382 316 4388 317
rect 4382 312 4383 316
rect 4387 312 4388 316
rect 4382 311 4388 312
rect 4614 316 4620 317
rect 4614 312 4615 316
rect 4619 312 4620 316
rect 4614 311 4620 312
rect 4822 316 4828 317
rect 4822 312 4823 316
rect 4827 312 4828 316
rect 4822 311 4828 312
rect 5014 316 5020 317
rect 5014 312 5015 316
rect 5019 312 5020 316
rect 5014 311 5020 312
rect 5198 316 5204 317
rect 5198 312 5199 316
rect 5203 312 5204 316
rect 5198 311 5204 312
rect 5382 316 5388 317
rect 5382 312 5383 316
rect 5387 312 5388 316
rect 5382 311 5388 312
rect 5542 316 5548 317
rect 5542 312 5543 316
rect 5547 312 5548 316
rect 5662 313 5663 317
rect 5667 313 5668 317
rect 5662 312 5668 313
rect 5542 311 5548 312
rect 1974 307 1980 308
rect 3798 307 3804 308
rect 322 301 328 302
rect 110 300 116 301
rect 110 296 111 300
rect 115 296 116 300
rect 322 297 323 301
rect 327 297 328 301
rect 322 296 328 297
rect 546 301 552 302
rect 546 297 547 301
rect 551 297 552 301
rect 546 296 552 297
rect 770 301 776 302
rect 770 297 771 301
rect 775 297 776 301
rect 770 296 776 297
rect 986 301 992 302
rect 986 297 987 301
rect 991 297 992 301
rect 986 296 992 297
rect 1202 301 1208 302
rect 1202 297 1203 301
rect 1207 297 1208 301
rect 1202 296 1208 297
rect 1426 301 1432 302
rect 3858 301 3864 302
rect 1426 297 1427 301
rect 1431 297 1432 301
rect 1426 296 1432 297
rect 1934 300 1940 301
rect 1934 296 1935 300
rect 1939 296 1940 300
rect 110 295 116 296
rect 1934 295 1940 296
rect 3838 300 3844 301
rect 3838 296 3839 300
rect 3843 296 3844 300
rect 3858 297 3859 301
rect 3863 297 3864 301
rect 3858 296 3864 297
rect 4106 301 4112 302
rect 4106 297 4107 301
rect 4111 297 4112 301
rect 4106 296 4112 297
rect 4354 301 4360 302
rect 4354 297 4355 301
rect 4359 297 4360 301
rect 4354 296 4360 297
rect 4586 301 4592 302
rect 4586 297 4587 301
rect 4591 297 4592 301
rect 4586 296 4592 297
rect 4794 301 4800 302
rect 4794 297 4795 301
rect 4799 297 4800 301
rect 4794 296 4800 297
rect 4986 301 4992 302
rect 4986 297 4987 301
rect 4991 297 4992 301
rect 4986 296 4992 297
rect 5170 301 5176 302
rect 5170 297 5171 301
rect 5175 297 5176 301
rect 5170 296 5176 297
rect 5354 301 5360 302
rect 5354 297 5355 301
rect 5359 297 5360 301
rect 5354 296 5360 297
rect 5514 301 5520 302
rect 5514 297 5515 301
rect 5519 297 5520 301
rect 5514 296 5520 297
rect 5662 300 5668 301
rect 5662 296 5663 300
rect 5667 296 5668 300
rect 3838 295 3844 296
rect 5662 295 5668 296
rect 3838 156 3844 157
rect 5662 156 5668 157
rect 1974 152 1980 153
rect 3798 152 3804 153
rect 1974 148 1975 152
rect 1979 148 1980 152
rect 1974 147 1980 148
rect 1994 151 2000 152
rect 1994 147 1995 151
rect 1999 147 2000 151
rect 1994 146 2000 147
rect 2170 151 2176 152
rect 2170 147 2171 151
rect 2175 147 2176 151
rect 2170 146 2176 147
rect 2362 151 2368 152
rect 2362 147 2363 151
rect 2367 147 2368 151
rect 2362 146 2368 147
rect 2546 151 2552 152
rect 2546 147 2547 151
rect 2551 147 2552 151
rect 2546 146 2552 147
rect 2722 151 2728 152
rect 2722 147 2723 151
rect 2727 147 2728 151
rect 2722 146 2728 147
rect 2890 151 2896 152
rect 2890 147 2891 151
rect 2895 147 2896 151
rect 2890 146 2896 147
rect 3050 151 3056 152
rect 3050 147 3051 151
rect 3055 147 3056 151
rect 3050 146 3056 147
rect 3202 151 3208 152
rect 3202 147 3203 151
rect 3207 147 3208 151
rect 3202 146 3208 147
rect 3354 151 3360 152
rect 3354 147 3355 151
rect 3359 147 3360 151
rect 3354 146 3360 147
rect 3514 151 3520 152
rect 3514 147 3515 151
rect 3519 147 3520 151
rect 3514 146 3520 147
rect 3650 151 3656 152
rect 3650 147 3651 151
rect 3655 147 3656 151
rect 3798 148 3799 152
rect 3803 148 3804 152
rect 3838 152 3839 156
rect 3843 152 3844 156
rect 3838 151 3844 152
rect 4290 155 4296 156
rect 4290 151 4291 155
rect 4295 151 4296 155
rect 4290 150 4296 151
rect 4426 155 4432 156
rect 4426 151 4427 155
rect 4431 151 4432 155
rect 4426 150 4432 151
rect 4562 155 4568 156
rect 4562 151 4563 155
rect 4567 151 4568 155
rect 4562 150 4568 151
rect 4698 155 4704 156
rect 4698 151 4699 155
rect 4703 151 4704 155
rect 4698 150 4704 151
rect 4834 155 4840 156
rect 4834 151 4835 155
rect 4839 151 4840 155
rect 4834 150 4840 151
rect 4970 155 4976 156
rect 4970 151 4971 155
rect 4975 151 4976 155
rect 4970 150 4976 151
rect 5106 155 5112 156
rect 5106 151 5107 155
rect 5111 151 5112 155
rect 5106 150 5112 151
rect 5242 155 5248 156
rect 5242 151 5243 155
rect 5247 151 5248 155
rect 5242 150 5248 151
rect 5378 155 5384 156
rect 5378 151 5379 155
rect 5383 151 5384 155
rect 5378 150 5384 151
rect 5514 155 5520 156
rect 5514 151 5515 155
rect 5519 151 5520 155
rect 5662 152 5663 156
rect 5667 152 5668 156
rect 5662 151 5668 152
rect 5514 150 5520 151
rect 3798 147 3804 148
rect 3650 146 3656 147
rect 4318 140 4324 141
rect 3838 139 3844 140
rect 2022 136 2028 137
rect 1974 135 1980 136
rect 110 132 116 133
rect 1934 132 1940 133
rect 110 128 111 132
rect 115 128 116 132
rect 110 127 116 128
rect 130 131 136 132
rect 130 127 131 131
rect 135 127 136 131
rect 130 126 136 127
rect 266 131 272 132
rect 266 127 267 131
rect 271 127 272 131
rect 266 126 272 127
rect 402 131 408 132
rect 402 127 403 131
rect 407 127 408 131
rect 402 126 408 127
rect 538 131 544 132
rect 538 127 539 131
rect 543 127 544 131
rect 538 126 544 127
rect 674 131 680 132
rect 674 127 675 131
rect 679 127 680 131
rect 674 126 680 127
rect 810 131 816 132
rect 810 127 811 131
rect 815 127 816 131
rect 810 126 816 127
rect 946 131 952 132
rect 946 127 947 131
rect 951 127 952 131
rect 946 126 952 127
rect 1082 131 1088 132
rect 1082 127 1083 131
rect 1087 127 1088 131
rect 1082 126 1088 127
rect 1226 131 1232 132
rect 1226 127 1227 131
rect 1231 127 1232 131
rect 1226 126 1232 127
rect 1370 131 1376 132
rect 1370 127 1371 131
rect 1375 127 1376 131
rect 1370 126 1376 127
rect 1514 131 1520 132
rect 1514 127 1515 131
rect 1519 127 1520 131
rect 1514 126 1520 127
rect 1650 131 1656 132
rect 1650 127 1651 131
rect 1655 127 1656 131
rect 1650 126 1656 127
rect 1786 131 1792 132
rect 1786 127 1787 131
rect 1791 127 1792 131
rect 1934 128 1935 132
rect 1939 128 1940 132
rect 1974 131 1975 135
rect 1979 131 1980 135
rect 2022 132 2023 136
rect 2027 132 2028 136
rect 2022 131 2028 132
rect 2198 136 2204 137
rect 2198 132 2199 136
rect 2203 132 2204 136
rect 2198 131 2204 132
rect 2390 136 2396 137
rect 2390 132 2391 136
rect 2395 132 2396 136
rect 2390 131 2396 132
rect 2574 136 2580 137
rect 2574 132 2575 136
rect 2579 132 2580 136
rect 2574 131 2580 132
rect 2750 136 2756 137
rect 2750 132 2751 136
rect 2755 132 2756 136
rect 2750 131 2756 132
rect 2918 136 2924 137
rect 2918 132 2919 136
rect 2923 132 2924 136
rect 2918 131 2924 132
rect 3078 136 3084 137
rect 3078 132 3079 136
rect 3083 132 3084 136
rect 3078 131 3084 132
rect 3230 136 3236 137
rect 3230 132 3231 136
rect 3235 132 3236 136
rect 3230 131 3236 132
rect 3382 136 3388 137
rect 3382 132 3383 136
rect 3387 132 3388 136
rect 3382 131 3388 132
rect 3542 136 3548 137
rect 3542 132 3543 136
rect 3547 132 3548 136
rect 3542 131 3548 132
rect 3678 136 3684 137
rect 3678 132 3679 136
rect 3683 132 3684 136
rect 3678 131 3684 132
rect 3798 135 3804 136
rect 3798 131 3799 135
rect 3803 131 3804 135
rect 3838 135 3839 139
rect 3843 135 3844 139
rect 4318 136 4319 140
rect 4323 136 4324 140
rect 4318 135 4324 136
rect 4454 140 4460 141
rect 4454 136 4455 140
rect 4459 136 4460 140
rect 4454 135 4460 136
rect 4590 140 4596 141
rect 4590 136 4591 140
rect 4595 136 4596 140
rect 4590 135 4596 136
rect 4726 140 4732 141
rect 4726 136 4727 140
rect 4731 136 4732 140
rect 4726 135 4732 136
rect 4862 140 4868 141
rect 4862 136 4863 140
rect 4867 136 4868 140
rect 4862 135 4868 136
rect 4998 140 5004 141
rect 4998 136 4999 140
rect 5003 136 5004 140
rect 4998 135 5004 136
rect 5134 140 5140 141
rect 5134 136 5135 140
rect 5139 136 5140 140
rect 5134 135 5140 136
rect 5270 140 5276 141
rect 5270 136 5271 140
rect 5275 136 5276 140
rect 5270 135 5276 136
rect 5406 140 5412 141
rect 5406 136 5407 140
rect 5411 136 5412 140
rect 5406 135 5412 136
rect 5542 140 5548 141
rect 5542 136 5543 140
rect 5547 136 5548 140
rect 5542 135 5548 136
rect 5662 139 5668 140
rect 5662 135 5663 139
rect 5667 135 5668 139
rect 3838 134 3844 135
rect 5662 134 5668 135
rect 1974 130 1980 131
rect 3798 130 3804 131
rect 1934 127 1940 128
rect 1786 126 1792 127
rect 158 116 164 117
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 158 112 159 116
rect 163 112 164 116
rect 158 111 164 112
rect 294 116 300 117
rect 294 112 295 116
rect 299 112 300 116
rect 294 111 300 112
rect 430 116 436 117
rect 430 112 431 116
rect 435 112 436 116
rect 430 111 436 112
rect 566 116 572 117
rect 566 112 567 116
rect 571 112 572 116
rect 566 111 572 112
rect 702 116 708 117
rect 702 112 703 116
rect 707 112 708 116
rect 702 111 708 112
rect 838 116 844 117
rect 838 112 839 116
rect 843 112 844 116
rect 838 111 844 112
rect 974 116 980 117
rect 974 112 975 116
rect 979 112 980 116
rect 974 111 980 112
rect 1110 116 1116 117
rect 1110 112 1111 116
rect 1115 112 1116 116
rect 1110 111 1116 112
rect 1254 116 1260 117
rect 1254 112 1255 116
rect 1259 112 1260 116
rect 1254 111 1260 112
rect 1398 116 1404 117
rect 1398 112 1399 116
rect 1403 112 1404 116
rect 1398 111 1404 112
rect 1542 116 1548 117
rect 1542 112 1543 116
rect 1547 112 1548 116
rect 1542 111 1548 112
rect 1678 116 1684 117
rect 1678 112 1679 116
rect 1683 112 1684 116
rect 1678 111 1684 112
rect 1814 116 1820 117
rect 1814 112 1815 116
rect 1819 112 1820 116
rect 1814 111 1820 112
rect 1934 115 1940 116
rect 1934 111 1935 115
rect 1939 111 1940 115
rect 110 110 116 111
rect 1934 110 1940 111
<< m3c >>
rect 111 5701 115 5705
rect 159 5700 163 5704
rect 295 5700 299 5704
rect 431 5700 435 5704
rect 567 5700 571 5704
rect 703 5700 707 5704
rect 839 5700 843 5704
rect 975 5700 979 5704
rect 1935 5701 1939 5705
rect 111 5684 115 5688
rect 131 5685 135 5689
rect 267 5685 271 5689
rect 403 5685 407 5689
rect 539 5685 543 5689
rect 675 5685 679 5689
rect 811 5685 815 5689
rect 947 5685 951 5689
rect 1935 5684 1939 5688
rect 1975 5641 1979 5645
rect 2103 5640 2107 5644
rect 2239 5640 2243 5644
rect 2375 5640 2379 5644
rect 2511 5640 2515 5644
rect 2647 5640 2651 5644
rect 2783 5640 2787 5644
rect 2919 5640 2923 5644
rect 3055 5640 3059 5644
rect 3191 5640 3195 5644
rect 3327 5640 3331 5644
rect 3463 5640 3467 5644
rect 3599 5640 3603 5644
rect 3799 5641 3803 5645
rect 1975 5624 1979 5628
rect 2075 5625 2079 5629
rect 2211 5625 2215 5629
rect 2347 5625 2351 5629
rect 2483 5625 2487 5629
rect 2619 5625 2623 5629
rect 2755 5625 2759 5629
rect 2891 5625 2895 5629
rect 3027 5625 3031 5629
rect 3163 5625 3167 5629
rect 3299 5625 3303 5629
rect 3435 5625 3439 5629
rect 3571 5625 3575 5629
rect 3799 5624 3803 5628
rect 111 5536 115 5540
rect 755 5535 759 5539
rect 891 5535 895 5539
rect 1027 5535 1031 5539
rect 1163 5535 1167 5539
rect 1935 5536 1939 5540
rect 3839 5540 3843 5544
rect 4243 5539 4247 5543
rect 4379 5539 4383 5543
rect 4515 5539 4519 5543
rect 4651 5539 4655 5543
rect 4787 5539 4791 5543
rect 4923 5539 4927 5543
rect 5059 5539 5063 5543
rect 5663 5540 5667 5544
rect 111 5519 115 5523
rect 783 5520 787 5524
rect 919 5520 923 5524
rect 1055 5520 1059 5524
rect 1191 5520 1195 5524
rect 1935 5519 1939 5523
rect 3839 5523 3843 5527
rect 4271 5524 4275 5528
rect 4407 5524 4411 5528
rect 4543 5524 4547 5528
rect 4679 5524 4683 5528
rect 4815 5524 4819 5528
rect 4951 5524 4955 5528
rect 5087 5524 5091 5528
rect 5663 5523 5667 5527
rect 1975 5492 1979 5496
rect 1995 5491 1999 5495
rect 2131 5491 2135 5495
rect 2267 5491 2271 5495
rect 2403 5491 2407 5495
rect 2555 5491 2559 5495
rect 2707 5491 2711 5495
rect 2859 5491 2863 5495
rect 3011 5491 3015 5495
rect 3163 5491 3167 5495
rect 3323 5491 3327 5495
rect 3483 5491 3487 5495
rect 3799 5492 3803 5496
rect 1975 5475 1979 5479
rect 2023 5476 2027 5480
rect 2159 5476 2163 5480
rect 2295 5476 2299 5480
rect 2431 5476 2435 5480
rect 2583 5476 2587 5480
rect 2735 5476 2739 5480
rect 2887 5476 2891 5480
rect 3039 5476 3043 5480
rect 3191 5476 3195 5480
rect 3351 5476 3355 5480
rect 3511 5476 3515 5480
rect 3799 5475 3803 5479
rect 3839 5465 3843 5469
rect 4455 5464 4459 5468
rect 4591 5464 4595 5468
rect 4727 5464 4731 5468
rect 4863 5464 4867 5468
rect 5663 5465 5667 5469
rect 111 5449 115 5453
rect 863 5448 867 5452
rect 999 5448 1003 5452
rect 1135 5448 1139 5452
rect 1271 5448 1275 5452
rect 1407 5448 1411 5452
rect 1543 5448 1547 5452
rect 1679 5448 1683 5452
rect 1815 5448 1819 5452
rect 1935 5449 1939 5453
rect 3839 5448 3843 5452
rect 4427 5449 4431 5453
rect 4563 5449 4567 5453
rect 4699 5449 4703 5453
rect 4835 5449 4839 5453
rect 5663 5448 5667 5452
rect 111 5432 115 5436
rect 835 5433 839 5437
rect 971 5433 975 5437
rect 1107 5433 1111 5437
rect 1243 5433 1247 5437
rect 1379 5433 1383 5437
rect 1515 5433 1519 5437
rect 1651 5433 1655 5437
rect 1787 5433 1791 5437
rect 1935 5432 1939 5436
rect 1975 5405 1979 5409
rect 2831 5404 2835 5408
rect 2967 5404 2971 5408
rect 3103 5404 3107 5408
rect 3239 5404 3243 5408
rect 3799 5405 3803 5409
rect 1975 5388 1979 5392
rect 2803 5389 2807 5393
rect 2939 5389 2943 5393
rect 3075 5389 3079 5393
rect 3211 5389 3215 5393
rect 3799 5388 3803 5392
rect 3839 5316 3843 5320
rect 4283 5315 4287 5319
rect 4483 5315 4487 5319
rect 4699 5315 4703 5319
rect 4931 5315 4935 5319
rect 5171 5315 5175 5319
rect 5419 5315 5423 5319
rect 5663 5316 5667 5320
rect 111 5300 115 5304
rect 427 5299 431 5303
rect 563 5299 567 5303
rect 699 5299 703 5303
rect 835 5299 839 5303
rect 971 5299 975 5303
rect 1107 5299 1111 5303
rect 1243 5299 1247 5303
rect 1379 5299 1383 5303
rect 1515 5299 1519 5303
rect 1651 5299 1655 5303
rect 1787 5299 1791 5303
rect 1935 5300 1939 5304
rect 3839 5299 3843 5303
rect 4311 5300 4315 5304
rect 4511 5300 4515 5304
rect 4727 5300 4731 5304
rect 4959 5300 4963 5304
rect 5199 5300 5203 5304
rect 5447 5300 5451 5304
rect 5663 5299 5667 5303
rect 111 5283 115 5287
rect 455 5284 459 5288
rect 591 5284 595 5288
rect 727 5284 731 5288
rect 863 5284 867 5288
rect 999 5284 1003 5288
rect 1135 5284 1139 5288
rect 1271 5284 1275 5288
rect 1407 5284 1411 5288
rect 1543 5284 1547 5288
rect 1679 5284 1683 5288
rect 1815 5284 1819 5288
rect 1935 5283 1939 5287
rect 111 5225 115 5229
rect 455 5224 459 5228
rect 591 5224 595 5228
rect 727 5224 731 5228
rect 863 5224 867 5228
rect 999 5224 1003 5228
rect 1135 5224 1139 5228
rect 1271 5224 1275 5228
rect 1407 5224 1411 5228
rect 1543 5224 1547 5228
rect 1679 5224 1683 5228
rect 1815 5224 1819 5228
rect 1935 5225 1939 5229
rect 1975 5220 1979 5224
rect 1995 5219 1999 5223
rect 2219 5219 2223 5223
rect 2467 5219 2471 5223
rect 2715 5219 2719 5223
rect 2971 5219 2975 5223
rect 3799 5220 3803 5224
rect 111 5208 115 5212
rect 427 5209 431 5213
rect 563 5209 567 5213
rect 699 5209 703 5213
rect 835 5209 839 5213
rect 971 5209 975 5213
rect 1107 5209 1111 5213
rect 1243 5209 1247 5213
rect 1379 5209 1383 5213
rect 1515 5209 1519 5213
rect 1651 5209 1655 5213
rect 3839 5213 3843 5217
rect 1787 5209 1791 5213
rect 3887 5212 3891 5216
rect 1935 5208 1939 5212
rect 4023 5212 4027 5216
rect 4159 5212 4163 5216
rect 4295 5212 4299 5216
rect 4431 5212 4435 5216
rect 4567 5212 4571 5216
rect 4703 5212 4707 5216
rect 4839 5212 4843 5216
rect 4991 5212 4995 5216
rect 5151 5212 5155 5216
rect 5319 5212 5323 5216
rect 5495 5212 5499 5216
rect 5663 5213 5667 5217
rect 1975 5203 1979 5207
rect 2023 5204 2027 5208
rect 2247 5204 2251 5208
rect 2495 5204 2499 5208
rect 2743 5204 2747 5208
rect 2999 5204 3003 5208
rect 3799 5203 3803 5207
rect 3839 5196 3843 5200
rect 3859 5197 3863 5201
rect 3995 5197 3999 5201
rect 4131 5197 4135 5201
rect 4267 5197 4271 5201
rect 4403 5197 4407 5201
rect 4539 5197 4543 5201
rect 4675 5197 4679 5201
rect 4811 5197 4815 5201
rect 4963 5197 4967 5201
rect 5123 5197 5127 5201
rect 5291 5197 5295 5201
rect 5467 5197 5471 5201
rect 5663 5196 5667 5200
rect 1975 5141 1979 5145
rect 2023 5140 2027 5144
rect 2159 5140 2163 5144
rect 2295 5140 2299 5144
rect 2431 5140 2435 5144
rect 2567 5140 2571 5144
rect 2703 5140 2707 5144
rect 2839 5140 2843 5144
rect 2975 5140 2979 5144
rect 3111 5140 3115 5144
rect 3247 5140 3251 5144
rect 3391 5140 3395 5144
rect 3543 5140 3547 5144
rect 3679 5140 3683 5144
rect 3799 5141 3803 5145
rect 1975 5124 1979 5128
rect 1995 5125 1999 5129
rect 2131 5125 2135 5129
rect 2267 5125 2271 5129
rect 2403 5125 2407 5129
rect 2539 5125 2543 5129
rect 2675 5125 2679 5129
rect 2811 5125 2815 5129
rect 2947 5125 2951 5129
rect 3083 5125 3087 5129
rect 3219 5125 3223 5129
rect 3363 5125 3367 5129
rect 3515 5125 3519 5129
rect 3651 5125 3655 5129
rect 3799 5124 3803 5128
rect 111 5060 115 5064
rect 267 5059 271 5063
rect 403 5059 407 5063
rect 539 5059 543 5063
rect 675 5059 679 5063
rect 811 5059 815 5063
rect 947 5059 951 5063
rect 1935 5060 1939 5064
rect 3839 5064 3843 5068
rect 3979 5063 3983 5067
rect 4275 5063 4279 5067
rect 4579 5063 4583 5067
rect 4883 5063 4887 5067
rect 5195 5063 5199 5067
rect 5515 5063 5519 5067
rect 5663 5064 5667 5068
rect 111 5043 115 5047
rect 295 5044 299 5048
rect 431 5044 435 5048
rect 567 5044 571 5048
rect 703 5044 707 5048
rect 839 5044 843 5048
rect 975 5044 979 5048
rect 1935 5043 1939 5047
rect 3839 5047 3843 5051
rect 4007 5048 4011 5052
rect 4303 5048 4307 5052
rect 4607 5048 4611 5052
rect 4911 5048 4915 5052
rect 5223 5048 5227 5052
rect 5543 5048 5547 5052
rect 5663 5047 5667 5051
rect 1975 4992 1979 4996
rect 3107 4991 3111 4995
rect 3243 4991 3247 4995
rect 3379 4991 3383 4995
rect 3515 4991 3519 4995
rect 3651 4991 3655 4995
rect 3799 4992 3803 4996
rect 111 4973 115 4977
rect 159 4972 163 4976
rect 295 4972 299 4976
rect 431 4972 435 4976
rect 567 4972 571 4976
rect 703 4972 707 4976
rect 1935 4973 1939 4977
rect 1975 4975 1979 4979
rect 3135 4976 3139 4980
rect 3271 4976 3275 4980
rect 3407 4976 3411 4980
rect 3543 4976 3547 4980
rect 3679 4976 3683 4980
rect 3799 4975 3803 4979
rect 3839 4973 3843 4977
rect 4863 4972 4867 4976
rect 4999 4972 5003 4976
rect 5135 4972 5139 4976
rect 5271 4972 5275 4976
rect 5407 4972 5411 4976
rect 5543 4972 5547 4976
rect 5663 4973 5667 4977
rect 111 4956 115 4960
rect 131 4957 135 4961
rect 267 4957 271 4961
rect 403 4957 407 4961
rect 539 4957 543 4961
rect 675 4957 679 4961
rect 1935 4956 1939 4960
rect 3839 4956 3843 4960
rect 4835 4957 4839 4961
rect 4971 4957 4975 4961
rect 5107 4957 5111 4961
rect 5243 4957 5247 4961
rect 5379 4957 5383 4961
rect 5515 4957 5519 4961
rect 5663 4956 5667 4960
rect 1975 4909 1979 4913
rect 3135 4908 3139 4912
rect 3271 4908 3275 4912
rect 3407 4908 3411 4912
rect 3543 4908 3547 4912
rect 3679 4908 3683 4912
rect 3799 4909 3803 4913
rect 1975 4892 1979 4896
rect 3107 4893 3111 4897
rect 3243 4893 3247 4897
rect 3379 4893 3383 4897
rect 3515 4893 3519 4897
rect 3651 4893 3655 4897
rect 3799 4892 3803 4896
rect 111 4816 115 4820
rect 131 4815 135 4819
rect 267 4815 271 4819
rect 403 4815 407 4819
rect 539 4815 543 4819
rect 675 4815 679 4819
rect 1935 4816 1939 4820
rect 3839 4812 3843 4816
rect 4483 4811 4487 4815
rect 4675 4811 4679 4815
rect 4875 4811 4879 4815
rect 5091 4811 5095 4815
rect 5315 4811 5319 4815
rect 5515 4811 5519 4815
rect 5663 4812 5667 4816
rect 111 4799 115 4803
rect 159 4800 163 4804
rect 295 4800 299 4804
rect 431 4800 435 4804
rect 567 4800 571 4804
rect 703 4800 707 4804
rect 1935 4799 1939 4803
rect 3839 4795 3843 4799
rect 4511 4796 4515 4800
rect 4703 4796 4707 4800
rect 4903 4796 4907 4800
rect 5119 4796 5123 4800
rect 5343 4796 5347 4800
rect 5543 4796 5547 4800
rect 5663 4795 5667 4799
rect 111 4737 115 4741
rect 159 4736 163 4740
rect 295 4736 299 4740
rect 431 4736 435 4740
rect 567 4736 571 4740
rect 703 4736 707 4740
rect 1935 4737 1939 4741
rect 1975 4732 1979 4736
rect 3107 4731 3111 4735
rect 3243 4731 3247 4735
rect 3379 4731 3383 4735
rect 3515 4731 3519 4735
rect 3651 4731 3655 4735
rect 3799 4732 3803 4736
rect 111 4720 115 4724
rect 131 4721 135 4725
rect 267 4721 271 4725
rect 403 4721 407 4725
rect 539 4721 543 4725
rect 675 4721 679 4725
rect 1935 4720 1939 4724
rect 1975 4715 1979 4719
rect 3135 4716 3139 4720
rect 3271 4716 3275 4720
rect 3407 4716 3411 4720
rect 3543 4716 3547 4720
rect 3679 4716 3683 4720
rect 3799 4715 3803 4719
rect 3839 4717 3843 4721
rect 4119 4716 4123 4720
rect 4375 4716 4379 4720
rect 4647 4716 4651 4720
rect 4943 4716 4947 4720
rect 5255 4716 5259 4720
rect 5543 4716 5547 4720
rect 5663 4717 5667 4721
rect 3839 4700 3843 4704
rect 4091 4701 4095 4705
rect 4347 4701 4351 4705
rect 4619 4701 4623 4705
rect 4915 4701 4919 4705
rect 5227 4701 5231 4705
rect 5515 4701 5519 4705
rect 5663 4700 5667 4704
rect 1975 4617 1979 4621
rect 2023 4616 2027 4620
rect 2159 4616 2163 4620
rect 2311 4616 2315 4620
rect 2479 4616 2483 4620
rect 2655 4616 2659 4620
rect 2831 4616 2835 4620
rect 3007 4616 3011 4620
rect 3183 4616 3187 4620
rect 3351 4616 3355 4620
rect 3527 4616 3531 4620
rect 3679 4616 3683 4620
rect 3799 4617 3803 4621
rect 1975 4600 1979 4604
rect 1995 4601 1999 4605
rect 2131 4601 2135 4605
rect 2283 4601 2287 4605
rect 2451 4601 2455 4605
rect 2627 4601 2631 4605
rect 2803 4601 2807 4605
rect 2979 4601 2983 4605
rect 3155 4601 3159 4605
rect 3323 4601 3327 4605
rect 3499 4601 3503 4605
rect 3651 4601 3655 4605
rect 3799 4600 3803 4604
rect 111 4580 115 4584
rect 211 4579 215 4583
rect 427 4579 431 4583
rect 667 4579 671 4583
rect 931 4579 935 4583
rect 1219 4579 1223 4583
rect 1515 4579 1519 4583
rect 1787 4579 1791 4583
rect 1935 4580 1939 4584
rect 111 4563 115 4567
rect 239 4564 243 4568
rect 455 4564 459 4568
rect 695 4564 699 4568
rect 959 4564 963 4568
rect 1247 4564 1251 4568
rect 1543 4564 1547 4568
rect 1815 4564 1819 4568
rect 1935 4563 1939 4567
rect 3839 4548 3843 4552
rect 4035 4547 4039 4551
rect 4331 4547 4335 4551
rect 4627 4547 4631 4551
rect 4931 4547 4935 4551
rect 5235 4547 5239 4551
rect 5515 4547 5519 4551
rect 5663 4548 5667 4552
rect 3839 4531 3843 4535
rect 4063 4532 4067 4536
rect 4359 4532 4363 4536
rect 4655 4532 4659 4536
rect 4959 4532 4963 4536
rect 5263 4532 5267 4536
rect 5543 4532 5547 4536
rect 5663 4531 5667 4535
rect 111 4505 115 4509
rect 447 4504 451 4508
rect 623 4504 627 4508
rect 807 4504 811 4508
rect 999 4504 1003 4508
rect 1199 4504 1203 4508
rect 1407 4504 1411 4508
rect 1623 4504 1627 4508
rect 1815 4504 1819 4508
rect 1935 4505 1939 4509
rect 111 4488 115 4492
rect 419 4489 423 4493
rect 595 4489 599 4493
rect 779 4489 783 4493
rect 971 4489 975 4493
rect 1171 4489 1175 4493
rect 1379 4489 1383 4493
rect 1595 4489 1599 4493
rect 1787 4489 1791 4493
rect 1935 4488 1939 4492
rect 1975 4468 1979 4472
rect 1995 4467 1999 4471
rect 2227 4467 2231 4471
rect 2459 4467 2463 4471
rect 2691 4467 2695 4471
rect 2915 4467 2919 4471
rect 3131 4467 3135 4471
rect 3355 4467 3359 4471
rect 3579 4467 3583 4471
rect 3799 4468 3803 4472
rect 3839 4457 3843 4461
rect 1975 4451 1979 4455
rect 2023 4452 2027 4456
rect 2255 4452 2259 4456
rect 2487 4452 2491 4456
rect 2719 4452 2723 4456
rect 2943 4452 2947 4456
rect 3159 4452 3163 4456
rect 3383 4452 3387 4456
rect 4311 4456 4315 4460
rect 3607 4452 3611 4456
rect 4535 4456 4539 4460
rect 4775 4456 4779 4460
rect 5023 4456 5027 4460
rect 5279 4456 5283 4460
rect 5543 4456 5547 4460
rect 5663 4457 5667 4461
rect 3799 4451 3803 4455
rect 3839 4440 3843 4444
rect 4283 4441 4287 4445
rect 4507 4441 4511 4445
rect 4747 4441 4751 4445
rect 4995 4441 4999 4445
rect 5251 4441 5255 4445
rect 5515 4441 5519 4445
rect 5663 4440 5667 4444
rect 1975 4389 1979 4393
rect 2119 4388 2123 4392
rect 2343 4388 2347 4392
rect 2567 4388 2571 4392
rect 2783 4388 2787 4392
rect 2991 4388 2995 4392
rect 3199 4388 3203 4392
rect 3407 4388 3411 4392
rect 3799 4389 3803 4393
rect 1975 4372 1979 4376
rect 2091 4373 2095 4377
rect 2315 4373 2319 4377
rect 2539 4373 2543 4377
rect 2755 4373 2759 4377
rect 2963 4373 2967 4377
rect 3171 4373 3175 4377
rect 3379 4373 3383 4377
rect 3799 4372 3803 4376
rect 111 4352 115 4356
rect 571 4351 575 4355
rect 739 4351 743 4355
rect 915 4351 919 4355
rect 1107 4351 1111 4355
rect 1299 4351 1303 4355
rect 1499 4351 1503 4355
rect 1707 4351 1711 4355
rect 1935 4352 1939 4356
rect 111 4335 115 4339
rect 599 4336 603 4340
rect 767 4336 771 4340
rect 943 4336 947 4340
rect 1135 4336 1139 4340
rect 1327 4336 1331 4340
rect 1527 4336 1531 4340
rect 1735 4336 1739 4340
rect 1935 4335 1939 4339
rect 3839 4288 3843 4292
rect 4515 4287 4519 4291
rect 4691 4287 4695 4291
rect 4875 4287 4879 4291
rect 5067 4287 5071 4291
rect 5267 4287 5271 4291
rect 5467 4287 5471 4291
rect 5663 4288 5667 4292
rect 111 4277 115 4281
rect 655 4276 659 4280
rect 823 4276 827 4280
rect 991 4276 995 4280
rect 1167 4276 1171 4280
rect 1343 4276 1347 4280
rect 1519 4276 1523 4280
rect 1703 4276 1707 4280
rect 1935 4277 1939 4281
rect 3839 4271 3843 4275
rect 4543 4272 4547 4276
rect 4719 4272 4723 4276
rect 4903 4272 4907 4276
rect 5095 4272 5099 4276
rect 5295 4272 5299 4276
rect 5495 4272 5499 4276
rect 5663 4271 5667 4275
rect 111 4260 115 4264
rect 627 4261 631 4265
rect 795 4261 799 4265
rect 963 4261 967 4265
rect 1139 4261 1143 4265
rect 1315 4261 1319 4265
rect 1491 4261 1495 4265
rect 1675 4261 1679 4265
rect 1935 4260 1939 4264
rect 1975 4232 1979 4236
rect 2019 4231 2023 4235
rect 2243 4231 2247 4235
rect 2459 4231 2463 4235
rect 2667 4231 2671 4235
rect 2875 4231 2879 4235
rect 3083 4231 3087 4235
rect 3291 4231 3295 4235
rect 3799 4232 3803 4236
rect 1975 4215 1979 4219
rect 2047 4216 2051 4220
rect 2271 4216 2275 4220
rect 2487 4216 2491 4220
rect 2695 4216 2699 4220
rect 2903 4216 2907 4220
rect 3111 4216 3115 4220
rect 3319 4216 3323 4220
rect 3799 4215 3803 4219
rect 3839 4193 3843 4197
rect 4815 4192 4819 4196
rect 4951 4192 4955 4196
rect 5087 4192 5091 4196
rect 5223 4192 5227 4196
rect 5359 4192 5363 4196
rect 5495 4192 5499 4196
rect 5663 4193 5667 4197
rect 3839 4176 3843 4180
rect 4787 4177 4791 4181
rect 4923 4177 4927 4181
rect 5059 4177 5063 4181
rect 5195 4177 5199 4181
rect 5331 4177 5335 4181
rect 5467 4177 5471 4181
rect 5663 4176 5667 4180
rect 1975 4153 1979 4157
rect 2023 4152 2027 4156
rect 2287 4152 2291 4156
rect 2551 4152 2555 4156
rect 2799 4152 2803 4156
rect 3039 4152 3043 4156
rect 3279 4152 3283 4156
rect 3519 4152 3523 4156
rect 3799 4153 3803 4157
rect 1975 4136 1979 4140
rect 1995 4137 1999 4141
rect 2259 4137 2263 4141
rect 2523 4137 2527 4141
rect 2771 4137 2775 4141
rect 3011 4137 3015 4141
rect 3251 4137 3255 4141
rect 3491 4137 3495 4141
rect 3799 4136 3803 4140
rect 111 4116 115 4120
rect 347 4115 351 4119
rect 515 4115 519 4119
rect 699 4115 703 4119
rect 891 4115 895 4119
rect 1099 4115 1103 4119
rect 1315 4115 1319 4119
rect 1531 4115 1535 4119
rect 1935 4116 1939 4120
rect 111 4099 115 4103
rect 375 4100 379 4104
rect 543 4100 547 4104
rect 727 4100 731 4104
rect 919 4100 923 4104
rect 1127 4100 1131 4104
rect 1343 4100 1347 4104
rect 1559 4100 1563 4104
rect 1935 4099 1939 4103
rect 3839 4040 3843 4044
rect 4939 4039 4943 4043
rect 5075 4039 5079 4043
rect 5211 4039 5215 4043
rect 5347 4039 5351 4043
rect 5483 4039 5487 4043
rect 5663 4040 5667 4044
rect 111 4025 115 4029
rect 231 4024 235 4028
rect 423 4024 427 4028
rect 615 4024 619 4028
rect 807 4024 811 4028
rect 991 4024 995 4028
rect 1167 4024 1171 4028
rect 1335 4024 1339 4028
rect 1503 4024 1507 4028
rect 1671 4024 1675 4028
rect 1815 4024 1819 4028
rect 1935 4025 1939 4029
rect 3839 4023 3843 4027
rect 4967 4024 4971 4028
rect 5103 4024 5107 4028
rect 5239 4024 5243 4028
rect 5375 4024 5379 4028
rect 5511 4024 5515 4028
rect 5663 4023 5667 4027
rect 111 4008 115 4012
rect 203 4009 207 4013
rect 395 4009 399 4013
rect 587 4009 591 4013
rect 779 4009 783 4013
rect 963 4009 967 4013
rect 1139 4009 1143 4013
rect 1307 4009 1311 4013
rect 1475 4009 1479 4013
rect 1643 4009 1647 4013
rect 1787 4009 1791 4013
rect 1935 4008 1939 4012
rect 1975 4004 1979 4008
rect 1995 4003 1999 4007
rect 2283 4003 2287 4007
rect 2587 4003 2591 4007
rect 2875 4003 2879 4007
rect 3163 4003 3167 4007
rect 3451 4003 3455 4007
rect 3799 4004 3803 4008
rect 1975 3987 1979 3991
rect 2023 3988 2027 3992
rect 2311 3988 2315 3992
rect 2615 3988 2619 3992
rect 2903 3988 2907 3992
rect 3191 3988 3195 3992
rect 3479 3988 3483 3992
rect 3799 3987 3803 3991
rect 3839 3957 3843 3961
rect 4831 3956 4835 3960
rect 4967 3956 4971 3960
rect 5111 3956 5115 3960
rect 5255 3956 5259 3960
rect 5407 3956 5411 3960
rect 5543 3956 5547 3960
rect 5663 3957 5667 3961
rect 3839 3940 3843 3944
rect 4803 3941 4807 3945
rect 4939 3941 4943 3945
rect 5083 3941 5087 3945
rect 5227 3941 5231 3945
rect 5379 3941 5383 3945
rect 5515 3941 5519 3945
rect 5663 3940 5667 3944
rect 1975 3909 1979 3913
rect 2671 3908 2675 3912
rect 2807 3908 2811 3912
rect 2943 3908 2947 3912
rect 3079 3908 3083 3912
rect 3215 3908 3219 3912
rect 3799 3909 3803 3913
rect 1975 3892 1979 3896
rect 2643 3893 2647 3897
rect 2779 3893 2783 3897
rect 2915 3893 2919 3897
rect 3051 3893 3055 3897
rect 3187 3893 3191 3897
rect 3799 3892 3803 3896
rect 111 3876 115 3880
rect 251 3875 255 3879
rect 451 3875 455 3879
rect 643 3875 647 3879
rect 827 3875 831 3879
rect 1003 3875 1007 3879
rect 1171 3875 1175 3879
rect 1331 3875 1335 3879
rect 1491 3875 1495 3879
rect 1651 3875 1655 3879
rect 1787 3875 1791 3879
rect 1935 3876 1939 3880
rect 111 3859 115 3863
rect 279 3860 283 3864
rect 479 3860 483 3864
rect 671 3860 675 3864
rect 855 3860 859 3864
rect 1031 3860 1035 3864
rect 1199 3860 1203 3864
rect 1359 3860 1363 3864
rect 1519 3860 1523 3864
rect 1679 3860 1683 3864
rect 1815 3860 1819 3864
rect 1935 3859 1939 3863
rect 111 3801 115 3805
rect 311 3800 315 3804
rect 511 3800 515 3804
rect 735 3800 739 3804
rect 991 3800 995 3804
rect 1263 3800 1267 3804
rect 1551 3800 1555 3804
rect 1815 3800 1819 3804
rect 1935 3801 1939 3805
rect 111 3784 115 3788
rect 283 3785 287 3789
rect 483 3785 487 3789
rect 707 3785 711 3789
rect 963 3785 967 3789
rect 1235 3785 1239 3789
rect 1523 3785 1527 3789
rect 1787 3785 1791 3789
rect 1935 3784 1939 3788
rect 3839 3788 3843 3792
rect 4499 3787 4503 3791
rect 4675 3787 4679 3791
rect 4875 3787 4879 3791
rect 5091 3787 5095 3791
rect 5315 3787 5319 3791
rect 5515 3787 5519 3791
rect 5663 3788 5667 3792
rect 3839 3771 3843 3775
rect 4527 3772 4531 3776
rect 4703 3772 4707 3776
rect 4903 3772 4907 3776
rect 5119 3772 5123 3776
rect 5343 3772 5347 3776
rect 5543 3772 5547 3776
rect 5663 3771 5667 3775
rect 1975 3748 1979 3752
rect 1995 3747 1999 3751
rect 2131 3747 2135 3751
rect 2283 3747 2287 3751
rect 2443 3747 2447 3751
rect 2603 3747 2607 3751
rect 2763 3747 2767 3751
rect 2923 3747 2927 3751
rect 3083 3747 3087 3751
rect 3243 3747 3247 3751
rect 3411 3747 3415 3751
rect 3799 3748 3803 3752
rect 1975 3731 1979 3735
rect 2023 3732 2027 3736
rect 2159 3732 2163 3736
rect 2311 3732 2315 3736
rect 2471 3732 2475 3736
rect 2631 3732 2635 3736
rect 2791 3732 2795 3736
rect 2951 3732 2955 3736
rect 3111 3732 3115 3736
rect 3271 3732 3275 3736
rect 3439 3732 3443 3736
rect 3799 3731 3803 3735
rect 3839 3689 3843 3693
rect 4271 3688 4275 3692
rect 4471 3688 4475 3692
rect 4695 3688 4699 3692
rect 4935 3688 4939 3692
rect 5191 3688 5195 3692
rect 5447 3688 5451 3692
rect 5663 3689 5667 3693
rect 3839 3672 3843 3676
rect 4243 3673 4247 3677
rect 4443 3673 4447 3677
rect 4667 3673 4671 3677
rect 4907 3673 4911 3677
rect 5163 3673 5167 3677
rect 5419 3673 5423 3677
rect 5663 3672 5667 3676
rect 1975 3665 1979 3669
rect 2047 3664 2051 3668
rect 2223 3664 2227 3668
rect 2407 3664 2411 3668
rect 2591 3664 2595 3668
rect 2783 3664 2787 3668
rect 2967 3664 2971 3668
rect 3151 3664 3155 3668
rect 3335 3664 3339 3668
rect 3519 3664 3523 3668
rect 3679 3664 3683 3668
rect 3799 3665 3803 3669
rect 1975 3648 1979 3652
rect 2019 3649 2023 3653
rect 2195 3649 2199 3653
rect 2379 3649 2383 3653
rect 2563 3649 2567 3653
rect 2755 3649 2759 3653
rect 2939 3649 2943 3653
rect 3123 3649 3127 3653
rect 3307 3649 3311 3653
rect 3491 3649 3495 3653
rect 3651 3649 3655 3653
rect 3799 3648 3803 3652
rect 111 3628 115 3632
rect 155 3627 159 3631
rect 291 3627 295 3631
rect 427 3627 431 3631
rect 563 3627 567 3631
rect 699 3627 703 3631
rect 835 3627 839 3631
rect 971 3627 975 3631
rect 1107 3627 1111 3631
rect 1243 3627 1247 3631
rect 1379 3627 1383 3631
rect 1515 3627 1519 3631
rect 1935 3628 1939 3632
rect 111 3611 115 3615
rect 183 3612 187 3616
rect 319 3612 323 3616
rect 455 3612 459 3616
rect 591 3612 595 3616
rect 727 3612 731 3616
rect 863 3612 867 3616
rect 999 3612 1003 3616
rect 1135 3612 1139 3616
rect 1271 3612 1275 3616
rect 1407 3612 1411 3616
rect 1543 3612 1547 3616
rect 1935 3611 1939 3615
rect 3839 3536 3843 3540
rect 3859 3535 3863 3539
rect 3995 3535 3999 3539
rect 4131 3535 4135 3539
rect 4267 3535 4271 3539
rect 4403 3535 4407 3539
rect 4539 3535 4543 3539
rect 4675 3535 4679 3539
rect 4811 3535 4815 3539
rect 4947 3535 4951 3539
rect 5663 3536 5667 3540
rect 3839 3519 3843 3523
rect 3887 3520 3891 3524
rect 4023 3520 4027 3524
rect 4159 3520 4163 3524
rect 4295 3520 4299 3524
rect 4431 3520 4435 3524
rect 4567 3520 4571 3524
rect 4703 3520 4707 3524
rect 4839 3520 4843 3524
rect 4975 3520 4979 3524
rect 5663 3519 5667 3523
rect 1975 3504 1979 3508
rect 2307 3503 2311 3507
rect 2443 3503 2447 3507
rect 2579 3503 2583 3507
rect 2715 3503 2719 3507
rect 3799 3504 3803 3508
rect 1975 3487 1979 3491
rect 2335 3488 2339 3492
rect 2471 3488 2475 3492
rect 2607 3488 2611 3492
rect 2743 3488 2747 3492
rect 3799 3487 3803 3491
rect 3839 3461 3843 3465
rect 3887 3460 3891 3464
rect 4023 3460 4027 3464
rect 4159 3460 4163 3464
rect 4295 3460 4299 3464
rect 4431 3460 4435 3464
rect 4567 3460 4571 3464
rect 4703 3460 4707 3464
rect 4839 3460 4843 3464
rect 4975 3460 4979 3464
rect 5111 3460 5115 3464
rect 5247 3460 5251 3464
rect 5383 3460 5387 3464
rect 5519 3460 5523 3464
rect 5663 3461 5667 3465
rect 3839 3444 3843 3448
rect 3859 3445 3863 3449
rect 3995 3445 3999 3449
rect 4131 3445 4135 3449
rect 4267 3445 4271 3449
rect 4403 3445 4407 3449
rect 4539 3445 4543 3449
rect 4675 3445 4679 3449
rect 4811 3445 4815 3449
rect 4947 3445 4951 3449
rect 5083 3445 5087 3449
rect 5219 3445 5223 3449
rect 5355 3445 5359 3449
rect 5491 3445 5495 3449
rect 5663 3444 5667 3448
rect 1975 3393 1979 3397
rect 2167 3392 2171 3396
rect 2303 3392 2307 3396
rect 2439 3392 2443 3396
rect 2575 3392 2579 3396
rect 2711 3392 2715 3396
rect 2847 3392 2851 3396
rect 2983 3392 2987 3396
rect 3799 3393 3803 3397
rect 1975 3376 1979 3380
rect 2139 3377 2143 3381
rect 2275 3377 2279 3381
rect 2411 3377 2415 3381
rect 2547 3377 2551 3381
rect 2683 3377 2687 3381
rect 2819 3377 2823 3381
rect 2955 3377 2959 3381
rect 3799 3376 3803 3380
rect 3839 3304 3843 3308
rect 3859 3303 3863 3307
rect 3995 3303 3999 3307
rect 4155 3303 4159 3307
rect 4315 3303 4319 3307
rect 4467 3303 4471 3307
rect 4627 3303 4631 3307
rect 4787 3303 4791 3307
rect 4947 3303 4951 3307
rect 5663 3304 5667 3308
rect 3839 3287 3843 3291
rect 3887 3288 3891 3292
rect 4023 3288 4027 3292
rect 4183 3288 4187 3292
rect 4343 3288 4347 3292
rect 4495 3288 4499 3292
rect 4655 3288 4659 3292
rect 4815 3288 4819 3292
rect 4975 3288 4979 3292
rect 5663 3287 5667 3291
rect 111 3265 115 3269
rect 159 3264 163 3268
rect 295 3264 299 3268
rect 431 3264 435 3268
rect 567 3264 571 3268
rect 703 3264 707 3268
rect 839 3264 843 3268
rect 975 3264 979 3268
rect 1111 3264 1115 3268
rect 1247 3264 1251 3268
rect 1383 3264 1387 3268
rect 1519 3264 1523 3268
rect 1935 3265 1939 3269
rect 111 3248 115 3252
rect 131 3249 135 3253
rect 267 3249 271 3253
rect 403 3249 407 3253
rect 539 3249 543 3253
rect 675 3249 679 3253
rect 811 3249 815 3253
rect 947 3249 951 3253
rect 1083 3249 1087 3253
rect 1219 3249 1223 3253
rect 1355 3249 1359 3253
rect 1491 3249 1495 3253
rect 1935 3248 1939 3252
rect 1975 3244 1979 3248
rect 2059 3243 2063 3247
rect 2203 3243 2207 3247
rect 2363 3243 2367 3247
rect 2539 3243 2543 3247
rect 2739 3243 2743 3247
rect 2955 3243 2959 3247
rect 3187 3243 3191 3247
rect 3427 3243 3431 3247
rect 3651 3243 3655 3247
rect 3799 3244 3803 3248
rect 1975 3227 1979 3231
rect 2087 3228 2091 3232
rect 2231 3228 2235 3232
rect 2391 3228 2395 3232
rect 2567 3228 2571 3232
rect 2767 3228 2771 3232
rect 2983 3228 2987 3232
rect 3215 3228 3219 3232
rect 3455 3228 3459 3232
rect 3679 3228 3683 3232
rect 3799 3227 3803 3231
rect 3839 3217 3843 3221
rect 4807 3216 4811 3220
rect 4943 3216 4947 3220
rect 5079 3216 5083 3220
rect 5215 3216 5219 3220
rect 5351 3216 5355 3220
rect 5663 3217 5667 3221
rect 3839 3200 3843 3204
rect 4779 3201 4783 3205
rect 4915 3201 4919 3205
rect 5051 3201 5055 3205
rect 5187 3201 5191 3205
rect 5323 3201 5327 3205
rect 5663 3200 5667 3204
rect 1975 3165 1979 3169
rect 2023 3164 2027 3168
rect 2159 3164 2163 3168
rect 2303 3164 2307 3168
rect 2455 3164 2459 3168
rect 2615 3164 2619 3168
rect 2783 3164 2787 3168
rect 2951 3164 2955 3168
rect 3127 3164 3131 3168
rect 3311 3164 3315 3168
rect 3503 3164 3507 3168
rect 3679 3164 3683 3168
rect 3799 3165 3803 3169
rect 1975 3148 1979 3152
rect 1995 3149 1999 3153
rect 2131 3149 2135 3153
rect 2275 3149 2279 3153
rect 2427 3149 2431 3153
rect 2587 3149 2591 3153
rect 2755 3149 2759 3153
rect 2923 3149 2927 3153
rect 3099 3149 3103 3153
rect 3283 3149 3287 3153
rect 3475 3149 3479 3153
rect 3651 3149 3655 3153
rect 3799 3148 3803 3152
rect 111 3088 115 3092
rect 291 3087 295 3091
rect 459 3087 463 3091
rect 627 3087 631 3091
rect 811 3087 815 3091
rect 995 3087 999 3091
rect 1187 3087 1191 3091
rect 1387 3087 1391 3091
rect 1595 3087 1599 3091
rect 1787 3087 1791 3091
rect 1935 3088 1939 3092
rect 111 3071 115 3075
rect 319 3072 323 3076
rect 487 3072 491 3076
rect 655 3072 659 3076
rect 839 3072 843 3076
rect 1023 3072 1027 3076
rect 1215 3072 1219 3076
rect 1415 3072 1419 3076
rect 1623 3072 1627 3076
rect 1815 3072 1819 3076
rect 1935 3071 1939 3075
rect 3839 3064 3843 3068
rect 4699 3063 4703 3067
rect 4835 3063 4839 3067
rect 4971 3063 4975 3067
rect 5107 3063 5111 3067
rect 5243 3063 5247 3067
rect 5379 3063 5383 3067
rect 5515 3063 5519 3067
rect 5663 3064 5667 3068
rect 3839 3047 3843 3051
rect 4727 3048 4731 3052
rect 4863 3048 4867 3052
rect 4999 3048 5003 3052
rect 5135 3048 5139 3052
rect 5271 3048 5275 3052
rect 5407 3048 5411 3052
rect 5543 3048 5547 3052
rect 5663 3047 5667 3051
rect 111 3013 115 3017
rect 327 3012 331 3016
rect 487 3012 491 3016
rect 647 3012 651 3016
rect 807 3012 811 3016
rect 959 3012 963 3016
rect 1103 3012 1107 3016
rect 1247 3012 1251 3016
rect 1391 3012 1395 3016
rect 1535 3012 1539 3016
rect 1679 3012 1683 3016
rect 1815 3012 1819 3016
rect 1935 3013 1939 3017
rect 111 2996 115 3000
rect 299 2997 303 3001
rect 459 2997 463 3001
rect 619 2997 623 3001
rect 779 2997 783 3001
rect 931 2997 935 3001
rect 1075 2997 1079 3001
rect 1219 2997 1223 3001
rect 1363 2997 1367 3001
rect 1507 2997 1511 3001
rect 1651 2997 1655 3001
rect 1787 2997 1791 3001
rect 1935 2996 1939 3000
rect 1975 2996 1979 3000
rect 2811 2995 2815 2999
rect 3003 2995 3007 2999
rect 3203 2995 3207 2999
rect 3403 2995 3407 2999
rect 3603 2995 3607 2999
rect 3799 2996 3803 3000
rect 3839 2989 3843 2993
rect 4367 2988 4371 2992
rect 4567 2988 4571 2992
rect 4783 2988 4787 2992
rect 5023 2988 5027 2992
rect 5279 2988 5283 2992
rect 5535 2988 5539 2992
rect 5663 2989 5667 2993
rect 1975 2979 1979 2983
rect 2839 2980 2843 2984
rect 3031 2980 3035 2984
rect 3231 2980 3235 2984
rect 3431 2980 3435 2984
rect 3631 2980 3635 2984
rect 3799 2979 3803 2983
rect 3839 2972 3843 2976
rect 4339 2973 4343 2977
rect 4539 2973 4543 2977
rect 4755 2973 4759 2977
rect 4995 2973 4999 2977
rect 5251 2973 5255 2977
rect 5507 2973 5511 2977
rect 5663 2972 5667 2976
rect 1975 2913 1979 2917
rect 2847 2912 2851 2916
rect 2983 2912 2987 2916
rect 3119 2912 3123 2916
rect 3255 2912 3259 2916
rect 3391 2912 3395 2916
rect 3527 2912 3531 2916
rect 3671 2912 3675 2916
rect 3799 2913 3803 2917
rect 1975 2896 1979 2900
rect 2819 2897 2823 2901
rect 2955 2897 2959 2901
rect 3091 2897 3095 2901
rect 3227 2897 3231 2901
rect 3363 2897 3367 2901
rect 3499 2897 3503 2901
rect 3643 2897 3647 2901
rect 3799 2896 3803 2900
rect 111 2864 115 2868
rect 155 2863 159 2867
rect 379 2863 383 2867
rect 595 2863 599 2867
rect 811 2863 815 2867
rect 1019 2863 1023 2867
rect 1219 2863 1223 2867
rect 1411 2863 1415 2867
rect 1611 2863 1615 2867
rect 1787 2863 1791 2867
rect 1935 2864 1939 2868
rect 111 2847 115 2851
rect 183 2848 187 2852
rect 407 2848 411 2852
rect 623 2848 627 2852
rect 839 2848 843 2852
rect 1047 2848 1051 2852
rect 1247 2848 1251 2852
rect 1439 2848 1443 2852
rect 1639 2848 1643 2852
rect 1815 2848 1819 2852
rect 1935 2847 1939 2851
rect 3839 2840 3843 2844
rect 4035 2839 4039 2843
rect 4315 2839 4319 2843
rect 4603 2839 4607 2843
rect 4907 2839 4911 2843
rect 5219 2839 5223 2843
rect 5515 2839 5519 2843
rect 5663 2840 5667 2844
rect 3839 2823 3843 2827
rect 4063 2824 4067 2828
rect 4343 2824 4347 2828
rect 4631 2824 4635 2828
rect 4935 2824 4939 2828
rect 5247 2824 5251 2828
rect 5543 2824 5547 2828
rect 5663 2823 5667 2827
rect 1975 2764 1979 2768
rect 2011 2763 2015 2767
rect 2251 2763 2255 2767
rect 2491 2763 2495 2767
rect 2731 2763 2735 2767
rect 2971 2763 2975 2767
rect 3799 2764 3803 2768
rect 111 2757 115 2761
rect 287 2756 291 2760
rect 423 2756 427 2760
rect 559 2756 563 2760
rect 695 2756 699 2760
rect 831 2756 835 2760
rect 1935 2757 1939 2761
rect 3839 2757 3843 2761
rect 3967 2756 3971 2760
rect 4255 2756 4259 2760
rect 4567 2756 4571 2760
rect 4895 2756 4899 2760
rect 5231 2756 5235 2760
rect 5543 2756 5547 2760
rect 5663 2757 5667 2761
rect 1975 2747 1979 2751
rect 2039 2748 2043 2752
rect 2279 2748 2283 2752
rect 2519 2748 2523 2752
rect 2759 2748 2763 2752
rect 2999 2748 3003 2752
rect 3799 2747 3803 2751
rect 111 2740 115 2744
rect 259 2741 263 2745
rect 395 2741 399 2745
rect 531 2741 535 2745
rect 667 2741 671 2745
rect 803 2741 807 2745
rect 1935 2740 1939 2744
rect 3839 2740 3843 2744
rect 3939 2741 3943 2745
rect 4227 2741 4231 2745
rect 4539 2741 4543 2745
rect 4867 2741 4871 2745
rect 5203 2741 5207 2745
rect 5515 2741 5519 2745
rect 5663 2740 5667 2744
rect 1975 2689 1979 2693
rect 2023 2688 2027 2692
rect 2159 2688 2163 2692
rect 2295 2688 2299 2692
rect 2431 2688 2435 2692
rect 2567 2688 2571 2692
rect 2703 2688 2707 2692
rect 2839 2688 2843 2692
rect 2975 2688 2979 2692
rect 3111 2688 3115 2692
rect 3247 2688 3251 2692
rect 3383 2688 3387 2692
rect 3799 2689 3803 2693
rect 1975 2672 1979 2676
rect 1995 2673 1999 2677
rect 2131 2673 2135 2677
rect 2267 2673 2271 2677
rect 2403 2673 2407 2677
rect 2539 2673 2543 2677
rect 2675 2673 2679 2677
rect 2811 2673 2815 2677
rect 2947 2673 2951 2677
rect 3083 2673 3087 2677
rect 3219 2673 3223 2677
rect 3355 2673 3359 2677
rect 3799 2672 3803 2676
rect 3839 2604 3843 2608
rect 4027 2603 4031 2607
rect 4275 2603 4279 2607
rect 4555 2603 4559 2607
rect 4867 2603 4871 2607
rect 5203 2603 5207 2607
rect 5515 2603 5519 2607
rect 5663 2604 5667 2608
rect 111 2588 115 2592
rect 539 2587 543 2591
rect 699 2587 703 2591
rect 883 2587 887 2591
rect 1091 2587 1095 2591
rect 1323 2587 1327 2591
rect 1563 2587 1567 2591
rect 1787 2587 1791 2591
rect 1935 2588 1939 2592
rect 3839 2587 3843 2591
rect 4055 2588 4059 2592
rect 4303 2588 4307 2592
rect 4583 2588 4587 2592
rect 4895 2588 4899 2592
rect 5231 2588 5235 2592
rect 5543 2588 5547 2592
rect 5663 2587 5667 2591
rect 111 2571 115 2575
rect 567 2572 571 2576
rect 727 2572 731 2576
rect 911 2572 915 2576
rect 1119 2572 1123 2576
rect 1351 2572 1355 2576
rect 1591 2572 1595 2576
rect 1815 2572 1819 2576
rect 1935 2571 1939 2575
rect 1975 2540 1979 2544
rect 1995 2539 1999 2543
rect 2203 2539 2207 2543
rect 2419 2539 2423 2543
rect 2627 2539 2631 2543
rect 2827 2539 2831 2543
rect 3019 2539 3023 2543
rect 3211 2539 3215 2543
rect 3403 2539 3407 2543
rect 3799 2540 3803 2544
rect 1975 2523 1979 2527
rect 2023 2524 2027 2528
rect 2231 2524 2235 2528
rect 2447 2524 2451 2528
rect 2655 2524 2659 2528
rect 2855 2524 2859 2528
rect 3047 2524 3051 2528
rect 3239 2524 3243 2528
rect 3431 2524 3435 2528
rect 3799 2523 3803 2527
rect 3839 2525 3843 2529
rect 4335 2524 4339 2528
rect 4559 2524 4563 2528
rect 4799 2524 4803 2528
rect 5047 2524 5051 2528
rect 5303 2524 5307 2528
rect 5543 2524 5547 2528
rect 5663 2525 5667 2529
rect 3839 2508 3843 2512
rect 4307 2509 4311 2513
rect 4531 2509 4535 2513
rect 4771 2509 4775 2513
rect 5019 2509 5023 2513
rect 5275 2509 5279 2513
rect 5515 2509 5519 2513
rect 5663 2508 5667 2512
rect 111 2501 115 2505
rect 695 2500 699 2504
rect 847 2500 851 2504
rect 999 2500 1003 2504
rect 1159 2500 1163 2504
rect 1327 2500 1331 2504
rect 1495 2500 1499 2504
rect 1663 2500 1667 2504
rect 1815 2500 1819 2504
rect 1935 2501 1939 2505
rect 111 2484 115 2488
rect 667 2485 671 2489
rect 819 2485 823 2489
rect 971 2485 975 2489
rect 1131 2485 1135 2489
rect 1299 2485 1303 2489
rect 1467 2485 1471 2489
rect 1635 2485 1639 2489
rect 1787 2485 1791 2489
rect 1935 2484 1939 2488
rect 1975 2457 1979 2461
rect 2319 2456 2323 2460
rect 2567 2456 2571 2460
rect 2799 2456 2803 2460
rect 3023 2456 3027 2460
rect 3239 2456 3243 2460
rect 3455 2456 3459 2460
rect 3671 2456 3675 2460
rect 3799 2457 3803 2461
rect 1975 2440 1979 2444
rect 2291 2441 2295 2445
rect 2539 2441 2543 2445
rect 2771 2441 2775 2445
rect 2995 2441 2999 2445
rect 3211 2441 3215 2445
rect 3427 2441 3431 2445
rect 3643 2441 3647 2445
rect 3799 2440 3803 2444
rect 3839 2360 3843 2364
rect 4491 2359 4495 2363
rect 4635 2359 4639 2363
rect 4795 2359 4799 2363
rect 4963 2359 4967 2363
rect 5139 2359 5143 2363
rect 5323 2359 5327 2363
rect 5515 2359 5519 2363
rect 5663 2360 5667 2364
rect 111 2344 115 2348
rect 355 2343 359 2347
rect 507 2343 511 2347
rect 675 2343 679 2347
rect 859 2343 863 2347
rect 1059 2343 1063 2347
rect 1267 2343 1271 2347
rect 1483 2343 1487 2347
rect 1699 2343 1703 2347
rect 1935 2344 1939 2348
rect 3839 2343 3843 2347
rect 4519 2344 4523 2348
rect 4663 2344 4667 2348
rect 4823 2344 4827 2348
rect 4991 2344 4995 2348
rect 5167 2344 5171 2348
rect 5351 2344 5355 2348
rect 5543 2344 5547 2348
rect 5663 2343 5667 2347
rect 111 2327 115 2331
rect 383 2328 387 2332
rect 535 2328 539 2332
rect 703 2328 707 2332
rect 887 2328 891 2332
rect 1087 2328 1091 2332
rect 1295 2328 1299 2332
rect 1511 2328 1515 2332
rect 1727 2328 1731 2332
rect 1935 2327 1939 2331
rect 1975 2300 1979 2304
rect 2331 2299 2335 2303
rect 2539 2299 2543 2303
rect 2739 2299 2743 2303
rect 2931 2299 2935 2303
rect 3123 2299 3127 2303
rect 3307 2299 3311 2303
rect 3491 2299 3495 2303
rect 3651 2299 3655 2303
rect 3799 2300 3803 2304
rect 1975 2283 1979 2287
rect 2359 2284 2363 2288
rect 2567 2284 2571 2288
rect 2767 2284 2771 2288
rect 2959 2284 2963 2288
rect 3151 2284 3155 2288
rect 3335 2284 3339 2288
rect 3519 2284 3523 2288
rect 3679 2284 3683 2288
rect 3799 2283 3803 2287
rect 111 2261 115 2265
rect 159 2260 163 2264
rect 335 2260 339 2264
rect 543 2260 547 2264
rect 759 2260 763 2264
rect 975 2260 979 2264
rect 1199 2260 1203 2264
rect 1431 2260 1435 2264
rect 1671 2260 1675 2264
rect 1935 2261 1939 2265
rect 3839 2265 3843 2269
rect 3887 2264 3891 2268
rect 4071 2264 4075 2268
rect 4271 2264 4275 2268
rect 4463 2264 4467 2268
rect 4655 2264 4659 2268
rect 4839 2264 4843 2268
rect 5015 2264 5019 2268
rect 5183 2264 5187 2268
rect 5359 2264 5363 2268
rect 5535 2264 5539 2268
rect 5663 2265 5667 2269
rect 111 2244 115 2248
rect 131 2245 135 2249
rect 307 2245 311 2249
rect 515 2245 519 2249
rect 731 2245 735 2249
rect 947 2245 951 2249
rect 1171 2245 1175 2249
rect 1403 2245 1407 2249
rect 1643 2245 1647 2249
rect 1935 2244 1939 2248
rect 3839 2248 3843 2252
rect 3859 2249 3863 2253
rect 4043 2249 4047 2253
rect 4243 2249 4247 2253
rect 4435 2249 4439 2253
rect 4627 2249 4631 2253
rect 4811 2249 4815 2253
rect 4987 2249 4991 2253
rect 5155 2249 5159 2253
rect 5331 2249 5335 2253
rect 5507 2249 5511 2253
rect 5663 2248 5667 2252
rect 1975 2197 1979 2201
rect 2463 2196 2467 2200
rect 2599 2196 2603 2200
rect 2735 2196 2739 2200
rect 3799 2197 3803 2201
rect 1975 2180 1979 2184
rect 2435 2181 2439 2185
rect 2571 2181 2575 2185
rect 2707 2181 2711 2185
rect 3799 2180 3803 2184
rect 3839 2116 3843 2120
rect 3859 2115 3863 2119
rect 4043 2115 4047 2119
rect 4251 2115 4255 2119
rect 4459 2115 4463 2119
rect 4659 2115 4663 2119
rect 4851 2115 4855 2119
rect 5035 2115 5039 2119
rect 5219 2115 5223 2119
rect 5411 2115 5415 2119
rect 5663 2116 5667 2120
rect 3839 2099 3843 2103
rect 3887 2100 3891 2104
rect 4071 2100 4075 2104
rect 4279 2100 4283 2104
rect 4487 2100 4491 2104
rect 4687 2100 4691 2104
rect 4879 2100 4883 2104
rect 5063 2100 5067 2104
rect 5247 2100 5251 2104
rect 5439 2100 5443 2104
rect 5663 2099 5667 2103
rect 111 2092 115 2096
rect 131 2091 135 2095
rect 299 2091 303 2095
rect 499 2091 503 2095
rect 715 2091 719 2095
rect 931 2091 935 2095
rect 1155 2091 1159 2095
rect 1387 2091 1391 2095
rect 1627 2091 1631 2095
rect 1935 2092 1939 2096
rect 111 2075 115 2079
rect 159 2076 163 2080
rect 327 2076 331 2080
rect 527 2076 531 2080
rect 743 2076 747 2080
rect 959 2076 963 2080
rect 1183 2076 1187 2080
rect 1415 2076 1419 2080
rect 1655 2076 1659 2080
rect 1935 2075 1939 2079
rect 3839 2021 3843 2025
rect 4287 2020 4291 2024
rect 1975 2016 1979 2020
rect 2419 2015 2423 2019
rect 2611 2015 2615 2019
rect 2795 2015 2799 2019
rect 2979 2015 2983 2019
rect 3155 2015 3159 2019
rect 3323 2015 3327 2019
rect 3499 2015 3503 2019
rect 3651 2015 3655 2019
rect 3799 2016 3803 2020
rect 4423 2020 4427 2024
rect 4559 2020 4563 2024
rect 4695 2020 4699 2024
rect 4839 2020 4843 2024
rect 5663 2021 5667 2025
rect 111 2009 115 2013
rect 159 2008 163 2012
rect 343 2008 347 2012
rect 567 2008 571 2012
rect 807 2008 811 2012
rect 1063 2008 1067 2012
rect 1335 2008 1339 2012
rect 1607 2008 1611 2012
rect 1935 2009 1939 2013
rect 1975 1999 1979 2003
rect 2447 2000 2451 2004
rect 2639 2000 2643 2004
rect 2823 2000 2827 2004
rect 3007 2000 3011 2004
rect 3183 2000 3187 2004
rect 3351 2000 3355 2004
rect 3527 2000 3531 2004
rect 3839 2004 3843 2008
rect 4259 2005 4263 2009
rect 4395 2005 4399 2009
rect 4531 2005 4535 2009
rect 4667 2005 4671 2009
rect 4811 2005 4815 2009
rect 5663 2004 5667 2008
rect 3679 2000 3683 2004
rect 3799 1999 3803 2003
rect 111 1992 115 1996
rect 131 1993 135 1997
rect 315 1993 319 1997
rect 539 1993 543 1997
rect 779 1993 783 1997
rect 1035 1993 1039 1997
rect 1307 1993 1311 1997
rect 1579 1993 1583 1997
rect 1935 1992 1939 1996
rect 1975 1929 1979 1933
rect 2359 1928 2363 1932
rect 2495 1928 2499 1932
rect 2631 1928 2635 1932
rect 2767 1928 2771 1932
rect 2903 1928 2907 1932
rect 3039 1928 3043 1932
rect 3175 1928 3179 1932
rect 3319 1928 3323 1932
rect 3799 1929 3803 1933
rect 1975 1912 1979 1916
rect 2331 1913 2335 1917
rect 2467 1913 2471 1917
rect 2603 1913 2607 1917
rect 2739 1913 2743 1917
rect 2875 1913 2879 1917
rect 3011 1913 3015 1917
rect 3147 1913 3151 1917
rect 3291 1913 3295 1917
rect 3799 1912 3803 1916
rect 111 1856 115 1860
rect 331 1855 335 1859
rect 499 1855 503 1859
rect 667 1855 671 1859
rect 843 1855 847 1859
rect 1027 1855 1031 1859
rect 1219 1855 1223 1859
rect 1411 1855 1415 1859
rect 1603 1855 1607 1859
rect 1935 1856 1939 1860
rect 3839 1852 3843 1856
rect 3955 1851 3959 1855
rect 4195 1851 4199 1855
rect 4467 1851 4471 1855
rect 4771 1851 4775 1855
rect 5091 1851 5095 1855
rect 5411 1851 5415 1855
rect 5663 1852 5667 1856
rect 111 1839 115 1843
rect 359 1840 363 1844
rect 527 1840 531 1844
rect 695 1840 699 1844
rect 871 1840 875 1844
rect 1055 1840 1059 1844
rect 1247 1840 1251 1844
rect 1439 1840 1443 1844
rect 1631 1840 1635 1844
rect 1935 1839 1939 1843
rect 3839 1835 3843 1839
rect 3983 1836 3987 1840
rect 4223 1836 4227 1840
rect 4495 1836 4499 1840
rect 4799 1836 4803 1840
rect 5119 1836 5123 1840
rect 5439 1836 5443 1840
rect 5663 1835 5667 1839
rect 1975 1780 1979 1784
rect 2211 1779 2215 1783
rect 2355 1779 2359 1783
rect 2499 1779 2503 1783
rect 2643 1779 2647 1783
rect 2787 1779 2791 1783
rect 2931 1779 2935 1783
rect 3083 1779 3087 1783
rect 3799 1780 3803 1784
rect 3839 1777 3843 1781
rect 4367 1776 4371 1780
rect 4575 1776 4579 1780
rect 4783 1776 4787 1780
rect 4983 1776 4987 1780
rect 5175 1776 5179 1780
rect 5367 1776 5371 1780
rect 5543 1776 5547 1780
rect 5663 1777 5667 1781
rect 111 1769 115 1773
rect 535 1768 539 1772
rect 695 1768 699 1772
rect 855 1768 859 1772
rect 1015 1768 1019 1772
rect 1183 1768 1187 1772
rect 1351 1768 1355 1772
rect 1519 1768 1523 1772
rect 1935 1769 1939 1773
rect 1975 1763 1979 1767
rect 2239 1764 2243 1768
rect 2383 1764 2387 1768
rect 2527 1764 2531 1768
rect 2671 1764 2675 1768
rect 2815 1764 2819 1768
rect 2959 1764 2963 1768
rect 3111 1764 3115 1768
rect 3799 1763 3803 1767
rect 3839 1760 3843 1764
rect 4339 1761 4343 1765
rect 4547 1761 4551 1765
rect 4755 1761 4759 1765
rect 4955 1761 4959 1765
rect 5147 1761 5151 1765
rect 5339 1761 5343 1765
rect 5515 1761 5519 1765
rect 5663 1760 5667 1764
rect 111 1752 115 1756
rect 507 1753 511 1757
rect 667 1753 671 1757
rect 827 1753 831 1757
rect 987 1753 991 1757
rect 1155 1753 1159 1757
rect 1323 1753 1327 1757
rect 1491 1753 1495 1757
rect 1935 1752 1939 1756
rect 1975 1705 1979 1709
rect 2023 1704 2027 1708
rect 2215 1704 2219 1708
rect 2407 1704 2411 1708
rect 2599 1704 2603 1708
rect 2791 1704 2795 1708
rect 2975 1704 2979 1708
rect 3151 1704 3155 1708
rect 3335 1704 3339 1708
rect 3519 1704 3523 1708
rect 3799 1705 3803 1709
rect 1975 1688 1979 1692
rect 1995 1689 1999 1693
rect 2187 1689 2191 1693
rect 2379 1689 2383 1693
rect 2571 1689 2575 1693
rect 2763 1689 2767 1693
rect 2947 1689 2951 1693
rect 3123 1689 3127 1693
rect 3307 1689 3311 1693
rect 3491 1689 3495 1693
rect 3799 1688 3803 1692
rect 3839 1612 3843 1616
rect 4603 1611 4607 1615
rect 4787 1611 4791 1615
rect 4971 1611 4975 1615
rect 5155 1611 5159 1615
rect 5339 1611 5343 1615
rect 5515 1611 5519 1615
rect 5663 1612 5667 1616
rect 111 1604 115 1608
rect 427 1603 431 1607
rect 611 1603 615 1607
rect 803 1603 807 1607
rect 995 1603 999 1607
rect 1187 1603 1191 1607
rect 1379 1603 1383 1607
rect 1935 1604 1939 1608
rect 3839 1595 3843 1599
rect 4631 1596 4635 1600
rect 4815 1596 4819 1600
rect 4999 1596 5003 1600
rect 5183 1596 5187 1600
rect 5367 1596 5371 1600
rect 5543 1596 5547 1600
rect 5663 1595 5667 1599
rect 111 1587 115 1591
rect 455 1588 459 1592
rect 639 1588 643 1592
rect 831 1588 835 1592
rect 1023 1588 1027 1592
rect 1215 1588 1219 1592
rect 1407 1588 1411 1592
rect 1935 1587 1939 1591
rect 1975 1556 1979 1560
rect 1995 1555 1999 1559
rect 2163 1555 2167 1559
rect 2371 1555 2375 1559
rect 2587 1555 2591 1559
rect 2803 1555 2807 1559
rect 3019 1555 3023 1559
rect 3235 1555 3239 1559
rect 3451 1555 3455 1559
rect 3651 1555 3655 1559
rect 3799 1556 3803 1560
rect 1975 1539 1979 1543
rect 2023 1540 2027 1544
rect 2191 1540 2195 1544
rect 2399 1540 2403 1544
rect 2615 1540 2619 1544
rect 2831 1540 2835 1544
rect 3047 1540 3051 1544
rect 3263 1540 3267 1544
rect 3479 1540 3483 1544
rect 3679 1540 3683 1544
rect 3799 1539 3803 1543
rect 111 1521 115 1525
rect 359 1520 363 1524
rect 631 1520 635 1524
rect 887 1520 891 1524
rect 1135 1520 1139 1524
rect 1367 1520 1371 1524
rect 1599 1520 1603 1524
rect 1815 1520 1819 1524
rect 1935 1521 1939 1525
rect 3839 1521 3843 1525
rect 3887 1520 3891 1524
rect 4031 1520 4035 1524
rect 4199 1520 4203 1524
rect 4367 1520 4371 1524
rect 4527 1520 4531 1524
rect 4695 1520 4699 1524
rect 4863 1520 4867 1524
rect 5031 1520 5035 1524
rect 5207 1520 5211 1524
rect 5383 1520 5387 1524
rect 5543 1520 5547 1524
rect 5663 1521 5667 1525
rect 111 1504 115 1508
rect 331 1505 335 1509
rect 603 1505 607 1509
rect 859 1505 863 1509
rect 1107 1505 1111 1509
rect 1339 1505 1343 1509
rect 1571 1505 1575 1509
rect 1787 1505 1791 1509
rect 1935 1504 1939 1508
rect 3839 1504 3843 1508
rect 3859 1505 3863 1509
rect 4003 1505 4007 1509
rect 4171 1505 4175 1509
rect 4339 1505 4343 1509
rect 4499 1505 4503 1509
rect 4667 1505 4671 1509
rect 4835 1505 4839 1509
rect 5003 1505 5007 1509
rect 5179 1505 5183 1509
rect 5355 1505 5359 1509
rect 5515 1505 5519 1509
rect 5663 1504 5667 1508
rect 111 1372 115 1376
rect 131 1371 135 1375
rect 307 1371 311 1375
rect 499 1371 503 1375
rect 683 1371 687 1375
rect 859 1371 863 1375
rect 1027 1371 1031 1375
rect 1187 1371 1191 1375
rect 1339 1371 1343 1375
rect 1491 1371 1495 1375
rect 1651 1371 1655 1375
rect 1787 1371 1791 1375
rect 1935 1372 1939 1376
rect 3839 1368 3843 1372
rect 3859 1367 3863 1371
rect 4003 1367 4007 1371
rect 4179 1367 4183 1371
rect 4355 1367 4359 1371
rect 4531 1367 4535 1371
rect 4707 1367 4711 1371
rect 4875 1367 4879 1371
rect 5043 1367 5047 1371
rect 5203 1367 5207 1371
rect 5371 1367 5375 1371
rect 5515 1367 5519 1371
rect 5663 1368 5667 1372
rect 111 1355 115 1359
rect 159 1356 163 1360
rect 335 1356 339 1360
rect 527 1356 531 1360
rect 711 1356 715 1360
rect 887 1356 891 1360
rect 1055 1356 1059 1360
rect 1215 1356 1219 1360
rect 1367 1356 1371 1360
rect 1519 1356 1523 1360
rect 1679 1356 1683 1360
rect 1815 1356 1819 1360
rect 1935 1355 1939 1359
rect 3839 1351 3843 1355
rect 3887 1352 3891 1356
rect 4031 1352 4035 1356
rect 4207 1352 4211 1356
rect 4383 1352 4387 1356
rect 4559 1352 4563 1356
rect 4735 1352 4739 1356
rect 4903 1352 4907 1356
rect 5071 1352 5075 1356
rect 5231 1352 5235 1356
rect 5399 1352 5403 1356
rect 5543 1352 5547 1356
rect 5663 1351 5667 1355
rect 111 1289 115 1293
rect 159 1288 163 1292
rect 375 1288 379 1292
rect 599 1288 603 1292
rect 807 1288 811 1292
rect 999 1288 1003 1292
rect 1175 1288 1179 1292
rect 1343 1288 1347 1292
rect 1511 1288 1515 1292
rect 1671 1288 1675 1292
rect 1815 1288 1819 1292
rect 1935 1289 1939 1293
rect 3839 1293 3843 1297
rect 3887 1292 3891 1296
rect 4175 1292 4179 1296
rect 4471 1292 4475 1296
rect 4751 1292 4755 1296
rect 5023 1292 5027 1296
rect 5287 1292 5291 1296
rect 5543 1292 5547 1296
rect 5663 1293 5667 1297
rect 111 1272 115 1276
rect 131 1273 135 1277
rect 347 1273 351 1277
rect 571 1273 575 1277
rect 779 1273 783 1277
rect 971 1273 975 1277
rect 1147 1273 1151 1277
rect 1315 1273 1319 1277
rect 1483 1273 1487 1277
rect 1643 1273 1647 1277
rect 1975 1277 1979 1281
rect 1787 1273 1791 1277
rect 3271 1276 3275 1280
rect 1935 1272 1939 1276
rect 3407 1276 3411 1280
rect 3543 1276 3547 1280
rect 3679 1276 3683 1280
rect 3799 1277 3803 1281
rect 3839 1276 3843 1280
rect 3859 1277 3863 1281
rect 4147 1277 4151 1281
rect 4443 1277 4447 1281
rect 4723 1277 4727 1281
rect 4995 1277 4999 1281
rect 5259 1277 5263 1281
rect 5515 1277 5519 1281
rect 5663 1276 5667 1280
rect 1975 1260 1979 1264
rect 3243 1261 3247 1265
rect 3379 1261 3383 1265
rect 3515 1261 3519 1265
rect 3651 1261 3655 1265
rect 3799 1260 3803 1264
rect 111 1140 115 1144
rect 131 1139 135 1143
rect 347 1139 351 1143
rect 563 1139 567 1143
rect 779 1139 783 1143
rect 987 1139 991 1143
rect 1195 1139 1199 1143
rect 1395 1139 1399 1143
rect 1603 1139 1607 1143
rect 1787 1139 1791 1143
rect 1935 1140 1939 1144
rect 3839 1132 3843 1136
rect 4427 1131 4431 1135
rect 4563 1131 4567 1135
rect 4699 1131 4703 1135
rect 4835 1131 4839 1135
rect 4971 1131 4975 1135
rect 5107 1131 5111 1135
rect 5243 1131 5247 1135
rect 5379 1131 5383 1135
rect 5515 1131 5519 1135
rect 5663 1132 5667 1136
rect 111 1123 115 1127
rect 159 1124 163 1128
rect 375 1124 379 1128
rect 591 1124 595 1128
rect 807 1124 811 1128
rect 1015 1124 1019 1128
rect 1223 1124 1227 1128
rect 1423 1124 1427 1128
rect 1631 1124 1635 1128
rect 1815 1124 1819 1128
rect 1935 1123 1939 1127
rect 1975 1116 1979 1120
rect 1995 1115 1999 1119
rect 2227 1115 2231 1119
rect 2467 1115 2471 1119
rect 2691 1115 2695 1119
rect 2907 1115 2911 1119
rect 3107 1115 3111 1119
rect 3299 1115 3303 1119
rect 3483 1115 3487 1119
rect 3651 1115 3655 1119
rect 3799 1116 3803 1120
rect 3839 1115 3843 1119
rect 4455 1116 4459 1120
rect 4591 1116 4595 1120
rect 4727 1116 4731 1120
rect 4863 1116 4867 1120
rect 4999 1116 5003 1120
rect 5135 1116 5139 1120
rect 5271 1116 5275 1120
rect 5407 1116 5411 1120
rect 5543 1116 5547 1120
rect 5663 1115 5667 1119
rect 1975 1099 1979 1103
rect 2023 1100 2027 1104
rect 2255 1100 2259 1104
rect 2495 1100 2499 1104
rect 2719 1100 2723 1104
rect 2935 1100 2939 1104
rect 3135 1100 3139 1104
rect 3327 1100 3331 1104
rect 3511 1100 3515 1104
rect 3679 1100 3683 1104
rect 3799 1099 3803 1103
rect 111 1041 115 1045
rect 471 1040 475 1044
rect 607 1040 611 1044
rect 743 1040 747 1044
rect 887 1040 891 1044
rect 1031 1040 1035 1044
rect 1935 1041 1939 1045
rect 1975 1041 1979 1045
rect 2183 1040 2187 1044
rect 2319 1040 2323 1044
rect 2455 1040 2459 1044
rect 2599 1040 2603 1044
rect 2743 1040 2747 1044
rect 2887 1040 2891 1044
rect 3031 1040 3035 1044
rect 3175 1040 3179 1044
rect 3319 1040 3323 1044
rect 3463 1040 3467 1044
rect 3799 1041 3803 1045
rect 3839 1041 3843 1045
rect 4367 1040 4371 1044
rect 4503 1040 4507 1044
rect 4639 1040 4643 1044
rect 4775 1040 4779 1044
rect 4911 1040 4915 1044
rect 5663 1041 5667 1045
rect 111 1024 115 1028
rect 443 1025 447 1029
rect 579 1025 583 1029
rect 715 1025 719 1029
rect 859 1025 863 1029
rect 1003 1025 1007 1029
rect 1935 1024 1939 1028
rect 1975 1024 1979 1028
rect 2155 1025 2159 1029
rect 2291 1025 2295 1029
rect 2427 1025 2431 1029
rect 2571 1025 2575 1029
rect 2715 1025 2719 1029
rect 2859 1025 2863 1029
rect 3003 1025 3007 1029
rect 3147 1025 3151 1029
rect 3291 1025 3295 1029
rect 3435 1025 3439 1029
rect 3799 1024 3803 1028
rect 3839 1024 3843 1028
rect 4339 1025 4343 1029
rect 4475 1025 4479 1029
rect 4611 1025 4615 1029
rect 4747 1025 4751 1029
rect 4883 1025 4887 1029
rect 5663 1024 5667 1028
rect 111 880 115 884
rect 259 879 263 883
rect 395 879 399 883
rect 531 879 535 883
rect 667 879 671 883
rect 803 879 807 883
rect 939 879 943 883
rect 1935 880 1939 884
rect 1975 880 1979 884
rect 1995 879 1999 883
rect 2131 879 2135 883
rect 2267 879 2271 883
rect 2403 879 2407 883
rect 2539 879 2543 883
rect 2675 879 2679 883
rect 2811 879 2815 883
rect 2947 879 2951 883
rect 3083 879 3087 883
rect 3219 879 3223 883
rect 3355 879 3359 883
rect 3491 879 3495 883
rect 3799 880 3803 884
rect 3839 880 3843 884
rect 4019 879 4023 883
rect 4155 879 4159 883
rect 4291 879 4295 883
rect 4427 879 4431 883
rect 4563 879 4567 883
rect 4699 879 4703 883
rect 5663 880 5667 884
rect 111 863 115 867
rect 287 864 291 868
rect 423 864 427 868
rect 559 864 563 868
rect 695 864 699 868
rect 831 864 835 868
rect 967 864 971 868
rect 1935 863 1939 867
rect 1975 863 1979 867
rect 2023 864 2027 868
rect 2159 864 2163 868
rect 2295 864 2299 868
rect 2431 864 2435 868
rect 2567 864 2571 868
rect 2703 864 2707 868
rect 2839 864 2843 868
rect 2975 864 2979 868
rect 3111 864 3115 868
rect 3247 864 3251 868
rect 3383 864 3387 868
rect 3519 864 3523 868
rect 3799 863 3803 867
rect 3839 863 3843 867
rect 4047 864 4051 868
rect 4183 864 4187 868
rect 4319 864 4323 868
rect 4455 864 4459 868
rect 4591 864 4595 868
rect 4727 864 4731 868
rect 5663 863 5667 867
rect 1975 805 1979 809
rect 2023 804 2027 808
rect 2167 804 2171 808
rect 2335 804 2339 808
rect 2495 804 2499 808
rect 2655 804 2659 808
rect 2823 804 2827 808
rect 2991 804 2995 808
rect 3799 805 3803 809
rect 111 793 115 797
rect 239 792 243 796
rect 439 792 443 796
rect 647 792 651 796
rect 855 792 859 796
rect 1063 792 1067 796
rect 1935 793 1939 797
rect 1975 788 1979 792
rect 1995 789 1999 793
rect 2139 789 2143 793
rect 2307 789 2311 793
rect 2467 789 2471 793
rect 2627 789 2631 793
rect 2795 789 2799 793
rect 2963 789 2967 793
rect 3799 788 3803 792
rect 3839 789 3843 793
rect 3887 788 3891 792
rect 4023 788 4027 792
rect 4159 788 4163 792
rect 4295 788 4299 792
rect 4431 788 4435 792
rect 4567 788 4571 792
rect 4703 788 4707 792
rect 4839 788 4843 792
rect 5663 789 5667 793
rect 111 776 115 780
rect 211 777 215 781
rect 411 777 415 781
rect 619 777 623 781
rect 827 777 831 781
rect 1035 777 1039 781
rect 1935 776 1939 780
rect 3839 772 3843 776
rect 3859 773 3863 777
rect 3995 773 3999 777
rect 4131 773 4135 777
rect 4267 773 4271 777
rect 4403 773 4407 777
rect 4539 773 4543 777
rect 4675 773 4679 777
rect 4811 773 4815 777
rect 5663 772 5667 776
rect 3839 640 3843 644
rect 3859 639 3863 643
rect 3995 639 3999 643
rect 4131 639 4135 643
rect 4267 639 4271 643
rect 4403 639 4407 643
rect 4539 639 4543 643
rect 4675 639 4679 643
rect 4811 639 4815 643
rect 4947 639 4951 643
rect 5083 639 5087 643
rect 5663 640 5667 644
rect 111 624 115 628
rect 131 623 135 627
rect 347 623 351 627
rect 587 623 591 627
rect 827 623 831 627
rect 1067 623 1071 627
rect 1315 623 1319 627
rect 1563 623 1567 627
rect 1787 623 1791 627
rect 1935 624 1939 628
rect 1975 628 1979 632
rect 1995 627 1999 631
rect 2299 627 2303 631
rect 2635 627 2639 631
rect 2979 627 2983 631
rect 3323 627 3327 631
rect 3651 627 3655 631
rect 3799 628 3803 632
rect 3839 623 3843 627
rect 3887 624 3891 628
rect 4023 624 4027 628
rect 4159 624 4163 628
rect 4295 624 4299 628
rect 4431 624 4435 628
rect 4567 624 4571 628
rect 4703 624 4707 628
rect 4839 624 4843 628
rect 4975 624 4979 628
rect 5111 624 5115 628
rect 5663 623 5667 627
rect 111 607 115 611
rect 159 608 163 612
rect 375 608 379 612
rect 615 608 619 612
rect 855 608 859 612
rect 1095 608 1099 612
rect 1343 608 1347 612
rect 1591 608 1595 612
rect 1815 608 1819 612
rect 1935 607 1939 611
rect 1975 611 1979 615
rect 2023 612 2027 616
rect 2327 612 2331 616
rect 2663 612 2667 616
rect 3007 612 3011 616
rect 3351 612 3355 616
rect 3679 612 3683 616
rect 3799 611 3803 615
rect 1975 553 1979 557
rect 2335 552 2339 556
rect 2527 552 2531 556
rect 2711 552 2715 556
rect 2887 552 2891 556
rect 3063 552 3067 556
rect 3231 552 3235 556
rect 3407 552 3411 556
rect 3583 552 3587 556
rect 3799 553 3803 557
rect 111 545 115 549
rect 159 544 163 548
rect 407 544 411 548
rect 671 544 675 548
rect 935 544 939 548
rect 1191 544 1195 548
rect 1447 544 1451 548
rect 1711 544 1715 548
rect 1935 545 1939 549
rect 3839 545 3843 549
rect 4047 544 4051 548
rect 4207 544 4211 548
rect 4367 544 4371 548
rect 4527 544 4531 548
rect 4687 544 4691 548
rect 5663 545 5667 549
rect 1975 536 1979 540
rect 2307 537 2311 541
rect 2499 537 2503 541
rect 2683 537 2687 541
rect 2859 537 2863 541
rect 3035 537 3039 541
rect 3203 537 3207 541
rect 3379 537 3383 541
rect 3555 537 3559 541
rect 3799 536 3803 540
rect 111 528 115 532
rect 131 529 135 533
rect 379 529 383 533
rect 643 529 647 533
rect 907 529 911 533
rect 1163 529 1167 533
rect 1419 529 1423 533
rect 1683 529 1687 533
rect 1935 528 1939 532
rect 3839 528 3843 532
rect 4019 529 4023 533
rect 4179 529 4183 533
rect 4339 529 4343 533
rect 4499 529 4503 533
rect 4659 529 4663 533
rect 5663 528 5667 532
rect 1975 404 1979 408
rect 2171 403 2175 407
rect 2315 403 2319 407
rect 2459 403 2463 407
rect 2603 403 2607 407
rect 2747 403 2751 407
rect 2891 403 2895 407
rect 3035 403 3039 407
rect 3799 404 3803 408
rect 111 396 115 400
rect 195 395 199 399
rect 427 395 431 399
rect 659 395 663 399
rect 883 395 887 399
rect 1099 395 1103 399
rect 1323 395 1327 399
rect 1547 395 1551 399
rect 1935 396 1939 400
rect 1975 387 1979 391
rect 2199 388 2203 392
rect 2343 388 2347 392
rect 2487 388 2491 392
rect 2631 388 2635 392
rect 2775 388 2779 392
rect 2919 388 2923 392
rect 3063 388 3067 392
rect 3799 387 3803 391
rect 3839 388 3843 392
rect 3931 387 3935 391
rect 4131 387 4135 391
rect 4331 387 4335 391
rect 4523 387 4527 391
rect 4723 387 4727 391
rect 4923 387 4927 391
rect 5663 388 5667 392
rect 111 379 115 383
rect 223 380 227 384
rect 455 380 459 384
rect 687 380 691 384
rect 911 380 915 384
rect 1127 380 1131 384
rect 1351 380 1355 384
rect 1575 380 1579 384
rect 1935 379 1939 383
rect 3839 371 3843 375
rect 3959 372 3963 376
rect 4159 372 4163 376
rect 4359 372 4363 376
rect 4551 372 4555 376
rect 4751 372 4755 376
rect 4951 372 4955 376
rect 5663 371 5667 375
rect 1975 325 1979 329
rect 2023 324 2027 328
rect 2175 324 2179 328
rect 2367 324 2371 328
rect 2591 324 2595 328
rect 2847 324 2851 328
rect 3119 324 3123 328
rect 3407 324 3411 328
rect 3679 324 3683 328
rect 3799 325 3803 329
rect 111 313 115 317
rect 351 312 355 316
rect 575 312 579 316
rect 799 312 803 316
rect 1015 312 1019 316
rect 1231 312 1235 316
rect 1455 312 1459 316
rect 1935 313 1939 317
rect 1975 308 1979 312
rect 1995 309 1999 313
rect 2147 309 2151 313
rect 2339 309 2343 313
rect 2563 309 2567 313
rect 2819 309 2823 313
rect 3091 309 3095 313
rect 3379 309 3383 313
rect 3839 313 3843 317
rect 3651 309 3655 313
rect 3887 312 3891 316
rect 3799 308 3803 312
rect 4135 312 4139 316
rect 4383 312 4387 316
rect 4615 312 4619 316
rect 4823 312 4827 316
rect 5015 312 5019 316
rect 5199 312 5203 316
rect 5383 312 5387 316
rect 5543 312 5547 316
rect 5663 313 5667 317
rect 111 296 115 300
rect 323 297 327 301
rect 547 297 551 301
rect 771 297 775 301
rect 987 297 991 301
rect 1203 297 1207 301
rect 1427 297 1431 301
rect 1935 296 1939 300
rect 3839 296 3843 300
rect 3859 297 3863 301
rect 4107 297 4111 301
rect 4355 297 4359 301
rect 4587 297 4591 301
rect 4795 297 4799 301
rect 4987 297 4991 301
rect 5171 297 5175 301
rect 5355 297 5359 301
rect 5515 297 5519 301
rect 5663 296 5667 300
rect 1975 148 1979 152
rect 1995 147 1999 151
rect 2171 147 2175 151
rect 2363 147 2367 151
rect 2547 147 2551 151
rect 2723 147 2727 151
rect 2891 147 2895 151
rect 3051 147 3055 151
rect 3203 147 3207 151
rect 3355 147 3359 151
rect 3515 147 3519 151
rect 3651 147 3655 151
rect 3799 148 3803 152
rect 3839 152 3843 156
rect 4291 151 4295 155
rect 4427 151 4431 155
rect 4563 151 4567 155
rect 4699 151 4703 155
rect 4835 151 4839 155
rect 4971 151 4975 155
rect 5107 151 5111 155
rect 5243 151 5247 155
rect 5379 151 5383 155
rect 5515 151 5519 155
rect 5663 152 5667 156
rect 111 128 115 132
rect 131 127 135 131
rect 267 127 271 131
rect 403 127 407 131
rect 539 127 543 131
rect 675 127 679 131
rect 811 127 815 131
rect 947 127 951 131
rect 1083 127 1087 131
rect 1227 127 1231 131
rect 1371 127 1375 131
rect 1515 127 1519 131
rect 1651 127 1655 131
rect 1787 127 1791 131
rect 1935 128 1939 132
rect 1975 131 1979 135
rect 2023 132 2027 136
rect 2199 132 2203 136
rect 2391 132 2395 136
rect 2575 132 2579 136
rect 2751 132 2755 136
rect 2919 132 2923 136
rect 3079 132 3083 136
rect 3231 132 3235 136
rect 3383 132 3387 136
rect 3543 132 3547 136
rect 3679 132 3683 136
rect 3799 131 3803 135
rect 3839 135 3843 139
rect 4319 136 4323 140
rect 4455 136 4459 140
rect 4591 136 4595 140
rect 4727 136 4731 140
rect 4863 136 4867 140
rect 4999 136 5003 140
rect 5135 136 5139 140
rect 5271 136 5275 140
rect 5407 136 5411 140
rect 5543 136 5547 140
rect 5663 135 5667 139
rect 111 111 115 115
rect 159 112 163 116
rect 295 112 299 116
rect 431 112 435 116
rect 567 112 571 116
rect 703 112 707 116
rect 839 112 843 116
rect 975 112 979 116
rect 1111 112 1115 116
rect 1255 112 1259 116
rect 1399 112 1403 116
rect 1543 112 1547 116
rect 1679 112 1683 116
rect 1815 112 1819 116
rect 1935 111 1939 115
<< m3 >>
rect 111 5734 115 5735
rect 111 5729 115 5730
rect 159 5734 163 5735
rect 159 5729 163 5730
rect 295 5734 299 5735
rect 295 5729 299 5730
rect 431 5734 435 5735
rect 431 5729 435 5730
rect 567 5734 571 5735
rect 567 5729 571 5730
rect 703 5734 707 5735
rect 703 5729 707 5730
rect 839 5734 843 5735
rect 839 5729 843 5730
rect 975 5734 979 5735
rect 975 5729 979 5730
rect 1935 5734 1939 5735
rect 1935 5729 1939 5730
rect 112 5706 114 5729
rect 110 5705 116 5706
rect 160 5705 162 5729
rect 296 5705 298 5729
rect 432 5705 434 5729
rect 568 5705 570 5729
rect 704 5705 706 5729
rect 840 5705 842 5729
rect 976 5705 978 5729
rect 1936 5706 1938 5729
rect 1934 5705 1940 5706
rect 110 5701 111 5705
rect 115 5701 116 5705
rect 110 5700 116 5701
rect 158 5704 164 5705
rect 158 5700 159 5704
rect 163 5700 164 5704
rect 158 5699 164 5700
rect 294 5704 300 5705
rect 294 5700 295 5704
rect 299 5700 300 5704
rect 294 5699 300 5700
rect 430 5704 436 5705
rect 430 5700 431 5704
rect 435 5700 436 5704
rect 430 5699 436 5700
rect 566 5704 572 5705
rect 566 5700 567 5704
rect 571 5700 572 5704
rect 566 5699 572 5700
rect 702 5704 708 5705
rect 702 5700 703 5704
rect 707 5700 708 5704
rect 702 5699 708 5700
rect 838 5704 844 5705
rect 838 5700 839 5704
rect 843 5700 844 5704
rect 838 5699 844 5700
rect 974 5704 980 5705
rect 974 5700 975 5704
rect 979 5700 980 5704
rect 1934 5701 1935 5705
rect 1939 5701 1940 5705
rect 1934 5700 1940 5701
rect 974 5699 980 5700
rect 130 5689 136 5690
rect 110 5688 116 5689
rect 110 5684 111 5688
rect 115 5684 116 5688
rect 130 5685 131 5689
rect 135 5685 136 5689
rect 130 5684 136 5685
rect 266 5689 272 5690
rect 266 5685 267 5689
rect 271 5685 272 5689
rect 266 5684 272 5685
rect 402 5689 408 5690
rect 402 5685 403 5689
rect 407 5685 408 5689
rect 402 5684 408 5685
rect 538 5689 544 5690
rect 538 5685 539 5689
rect 543 5685 544 5689
rect 538 5684 544 5685
rect 674 5689 680 5690
rect 674 5685 675 5689
rect 679 5685 680 5689
rect 674 5684 680 5685
rect 810 5689 816 5690
rect 810 5685 811 5689
rect 815 5685 816 5689
rect 810 5684 816 5685
rect 946 5689 952 5690
rect 946 5685 947 5689
rect 951 5685 952 5689
rect 946 5684 952 5685
rect 1934 5688 1940 5689
rect 1934 5684 1935 5688
rect 1939 5684 1940 5688
rect 110 5683 116 5684
rect 112 5607 114 5683
rect 132 5607 134 5684
rect 268 5607 270 5684
rect 404 5607 406 5684
rect 540 5607 542 5684
rect 676 5607 678 5684
rect 812 5607 814 5684
rect 948 5607 950 5684
rect 1934 5683 1940 5684
rect 1936 5607 1938 5683
rect 1975 5674 1979 5675
rect 1975 5669 1979 5670
rect 2103 5674 2107 5675
rect 2103 5669 2107 5670
rect 2239 5674 2243 5675
rect 2239 5669 2243 5670
rect 2375 5674 2379 5675
rect 2375 5669 2379 5670
rect 2511 5674 2515 5675
rect 2511 5669 2515 5670
rect 2647 5674 2651 5675
rect 2647 5669 2651 5670
rect 2783 5674 2787 5675
rect 2783 5669 2787 5670
rect 2919 5674 2923 5675
rect 2919 5669 2923 5670
rect 3055 5674 3059 5675
rect 3055 5669 3059 5670
rect 3191 5674 3195 5675
rect 3191 5669 3195 5670
rect 3327 5674 3331 5675
rect 3327 5669 3331 5670
rect 3463 5674 3467 5675
rect 3463 5669 3467 5670
rect 3599 5674 3603 5675
rect 3599 5669 3603 5670
rect 3799 5674 3803 5675
rect 3799 5669 3803 5670
rect 1976 5646 1978 5669
rect 1974 5645 1980 5646
rect 2104 5645 2106 5669
rect 2240 5645 2242 5669
rect 2376 5645 2378 5669
rect 2512 5645 2514 5669
rect 2648 5645 2650 5669
rect 2784 5645 2786 5669
rect 2920 5645 2922 5669
rect 3056 5645 3058 5669
rect 3192 5645 3194 5669
rect 3328 5645 3330 5669
rect 3464 5645 3466 5669
rect 3600 5645 3602 5669
rect 3800 5646 3802 5669
rect 3798 5645 3804 5646
rect 1974 5641 1975 5645
rect 1979 5641 1980 5645
rect 1974 5640 1980 5641
rect 2102 5644 2108 5645
rect 2102 5640 2103 5644
rect 2107 5640 2108 5644
rect 2102 5639 2108 5640
rect 2238 5644 2244 5645
rect 2238 5640 2239 5644
rect 2243 5640 2244 5644
rect 2238 5639 2244 5640
rect 2374 5644 2380 5645
rect 2374 5640 2375 5644
rect 2379 5640 2380 5644
rect 2374 5639 2380 5640
rect 2510 5644 2516 5645
rect 2510 5640 2511 5644
rect 2515 5640 2516 5644
rect 2510 5639 2516 5640
rect 2646 5644 2652 5645
rect 2646 5640 2647 5644
rect 2651 5640 2652 5644
rect 2646 5639 2652 5640
rect 2782 5644 2788 5645
rect 2782 5640 2783 5644
rect 2787 5640 2788 5644
rect 2782 5639 2788 5640
rect 2918 5644 2924 5645
rect 2918 5640 2919 5644
rect 2923 5640 2924 5644
rect 2918 5639 2924 5640
rect 3054 5644 3060 5645
rect 3054 5640 3055 5644
rect 3059 5640 3060 5644
rect 3054 5639 3060 5640
rect 3190 5644 3196 5645
rect 3190 5640 3191 5644
rect 3195 5640 3196 5644
rect 3190 5639 3196 5640
rect 3326 5644 3332 5645
rect 3326 5640 3327 5644
rect 3331 5640 3332 5644
rect 3326 5639 3332 5640
rect 3462 5644 3468 5645
rect 3462 5640 3463 5644
rect 3467 5640 3468 5644
rect 3462 5639 3468 5640
rect 3598 5644 3604 5645
rect 3598 5640 3599 5644
rect 3603 5640 3604 5644
rect 3798 5641 3799 5645
rect 3803 5641 3804 5645
rect 3798 5640 3804 5641
rect 3598 5639 3604 5640
rect 2074 5629 2080 5630
rect 1974 5628 1980 5629
rect 1974 5624 1975 5628
rect 1979 5624 1980 5628
rect 2074 5625 2075 5629
rect 2079 5625 2080 5629
rect 2074 5624 2080 5625
rect 2210 5629 2216 5630
rect 2210 5625 2211 5629
rect 2215 5625 2216 5629
rect 2210 5624 2216 5625
rect 2346 5629 2352 5630
rect 2346 5625 2347 5629
rect 2351 5625 2352 5629
rect 2346 5624 2352 5625
rect 2482 5629 2488 5630
rect 2482 5625 2483 5629
rect 2487 5625 2488 5629
rect 2482 5624 2488 5625
rect 2618 5629 2624 5630
rect 2618 5625 2619 5629
rect 2623 5625 2624 5629
rect 2618 5624 2624 5625
rect 2754 5629 2760 5630
rect 2754 5625 2755 5629
rect 2759 5625 2760 5629
rect 2754 5624 2760 5625
rect 2890 5629 2896 5630
rect 2890 5625 2891 5629
rect 2895 5625 2896 5629
rect 2890 5624 2896 5625
rect 3026 5629 3032 5630
rect 3026 5625 3027 5629
rect 3031 5625 3032 5629
rect 3026 5624 3032 5625
rect 3162 5629 3168 5630
rect 3162 5625 3163 5629
rect 3167 5625 3168 5629
rect 3162 5624 3168 5625
rect 3298 5629 3304 5630
rect 3298 5625 3299 5629
rect 3303 5625 3304 5629
rect 3298 5624 3304 5625
rect 3434 5629 3440 5630
rect 3434 5625 3435 5629
rect 3439 5625 3440 5629
rect 3434 5624 3440 5625
rect 3570 5629 3576 5630
rect 3570 5625 3571 5629
rect 3575 5625 3576 5629
rect 3570 5624 3576 5625
rect 3798 5628 3804 5629
rect 3798 5624 3799 5628
rect 3803 5624 3804 5628
rect 1974 5623 1980 5624
rect 111 5606 115 5607
rect 111 5601 115 5602
rect 131 5606 135 5607
rect 131 5601 135 5602
rect 267 5606 271 5607
rect 267 5601 271 5602
rect 403 5606 407 5607
rect 403 5601 407 5602
rect 539 5606 543 5607
rect 539 5601 543 5602
rect 675 5606 679 5607
rect 675 5601 679 5602
rect 755 5606 759 5607
rect 755 5601 759 5602
rect 811 5606 815 5607
rect 811 5601 815 5602
rect 891 5606 895 5607
rect 891 5601 895 5602
rect 947 5606 951 5607
rect 947 5601 951 5602
rect 1027 5606 1031 5607
rect 1027 5601 1031 5602
rect 1163 5606 1167 5607
rect 1163 5601 1167 5602
rect 1935 5606 1939 5607
rect 1935 5601 1939 5602
rect 112 5541 114 5601
rect 110 5540 116 5541
rect 756 5540 758 5601
rect 892 5540 894 5601
rect 1028 5540 1030 5601
rect 1164 5540 1166 5601
rect 1936 5541 1938 5601
rect 1976 5563 1978 5623
rect 2076 5563 2078 5624
rect 2212 5563 2214 5624
rect 2348 5563 2350 5624
rect 2484 5563 2486 5624
rect 2620 5563 2622 5624
rect 2756 5563 2758 5624
rect 2892 5563 2894 5624
rect 3028 5563 3030 5624
rect 3164 5563 3166 5624
rect 3300 5563 3302 5624
rect 3436 5563 3438 5624
rect 3572 5563 3574 5624
rect 3798 5623 3804 5624
rect 3800 5563 3802 5623
rect 3839 5610 3843 5611
rect 3839 5605 3843 5606
rect 4243 5610 4247 5611
rect 4243 5605 4247 5606
rect 4379 5610 4383 5611
rect 4379 5605 4383 5606
rect 4515 5610 4519 5611
rect 4515 5605 4519 5606
rect 4651 5610 4655 5611
rect 4651 5605 4655 5606
rect 4787 5610 4791 5611
rect 4787 5605 4791 5606
rect 4923 5610 4927 5611
rect 4923 5605 4927 5606
rect 5059 5610 5063 5611
rect 5059 5605 5063 5606
rect 5663 5610 5667 5611
rect 5663 5605 5667 5606
rect 1975 5562 1979 5563
rect 1975 5557 1979 5558
rect 1995 5562 1999 5563
rect 1995 5557 1999 5558
rect 2075 5562 2079 5563
rect 2075 5557 2079 5558
rect 2131 5562 2135 5563
rect 2131 5557 2135 5558
rect 2211 5562 2215 5563
rect 2211 5557 2215 5558
rect 2267 5562 2271 5563
rect 2267 5557 2271 5558
rect 2347 5562 2351 5563
rect 2347 5557 2351 5558
rect 2403 5562 2407 5563
rect 2403 5557 2407 5558
rect 2483 5562 2487 5563
rect 2483 5557 2487 5558
rect 2555 5562 2559 5563
rect 2555 5557 2559 5558
rect 2619 5562 2623 5563
rect 2619 5557 2623 5558
rect 2707 5562 2711 5563
rect 2707 5557 2711 5558
rect 2755 5562 2759 5563
rect 2755 5557 2759 5558
rect 2859 5562 2863 5563
rect 2859 5557 2863 5558
rect 2891 5562 2895 5563
rect 2891 5557 2895 5558
rect 3011 5562 3015 5563
rect 3011 5557 3015 5558
rect 3027 5562 3031 5563
rect 3027 5557 3031 5558
rect 3163 5562 3167 5563
rect 3163 5557 3167 5558
rect 3299 5562 3303 5563
rect 3299 5557 3303 5558
rect 3323 5562 3327 5563
rect 3323 5557 3327 5558
rect 3435 5562 3439 5563
rect 3435 5557 3439 5558
rect 3483 5562 3487 5563
rect 3483 5557 3487 5558
rect 3571 5562 3575 5563
rect 3571 5557 3575 5558
rect 3799 5562 3803 5563
rect 3799 5557 3803 5558
rect 1934 5540 1940 5541
rect 110 5536 111 5540
rect 115 5536 116 5540
rect 110 5535 116 5536
rect 754 5539 760 5540
rect 754 5535 755 5539
rect 759 5535 760 5539
rect 754 5534 760 5535
rect 890 5539 896 5540
rect 890 5535 891 5539
rect 895 5535 896 5539
rect 890 5534 896 5535
rect 1026 5539 1032 5540
rect 1026 5535 1027 5539
rect 1031 5535 1032 5539
rect 1026 5534 1032 5535
rect 1162 5539 1168 5540
rect 1162 5535 1163 5539
rect 1167 5535 1168 5539
rect 1934 5536 1935 5540
rect 1939 5536 1940 5540
rect 1934 5535 1940 5536
rect 1162 5534 1168 5535
rect 782 5524 788 5525
rect 110 5523 116 5524
rect 110 5519 111 5523
rect 115 5519 116 5523
rect 782 5520 783 5524
rect 787 5520 788 5524
rect 782 5519 788 5520
rect 918 5524 924 5525
rect 918 5520 919 5524
rect 923 5520 924 5524
rect 918 5519 924 5520
rect 1054 5524 1060 5525
rect 1054 5520 1055 5524
rect 1059 5520 1060 5524
rect 1054 5519 1060 5520
rect 1190 5524 1196 5525
rect 1190 5520 1191 5524
rect 1195 5520 1196 5524
rect 1190 5519 1196 5520
rect 1934 5523 1940 5524
rect 1934 5519 1935 5523
rect 1939 5519 1940 5523
rect 110 5518 116 5519
rect 112 5483 114 5518
rect 784 5483 786 5519
rect 920 5483 922 5519
rect 1056 5483 1058 5519
rect 1192 5483 1194 5519
rect 1934 5518 1940 5519
rect 1936 5483 1938 5518
rect 1976 5497 1978 5557
rect 1974 5496 1980 5497
rect 1996 5496 1998 5557
rect 2132 5496 2134 5557
rect 2268 5496 2270 5557
rect 2404 5496 2406 5557
rect 2556 5496 2558 5557
rect 2708 5496 2710 5557
rect 2860 5496 2862 5557
rect 3012 5496 3014 5557
rect 3164 5496 3166 5557
rect 3324 5496 3326 5557
rect 3484 5496 3486 5557
rect 3800 5497 3802 5557
rect 3840 5545 3842 5605
rect 3838 5544 3844 5545
rect 4244 5544 4246 5605
rect 4380 5544 4382 5605
rect 4516 5544 4518 5605
rect 4652 5544 4654 5605
rect 4788 5544 4790 5605
rect 4924 5544 4926 5605
rect 5060 5544 5062 5605
rect 5664 5545 5666 5605
rect 5662 5544 5668 5545
rect 3838 5540 3839 5544
rect 3843 5540 3844 5544
rect 3838 5539 3844 5540
rect 4242 5543 4248 5544
rect 4242 5539 4243 5543
rect 4247 5539 4248 5543
rect 4242 5538 4248 5539
rect 4378 5543 4384 5544
rect 4378 5539 4379 5543
rect 4383 5539 4384 5543
rect 4378 5538 4384 5539
rect 4514 5543 4520 5544
rect 4514 5539 4515 5543
rect 4519 5539 4520 5543
rect 4514 5538 4520 5539
rect 4650 5543 4656 5544
rect 4650 5539 4651 5543
rect 4655 5539 4656 5543
rect 4650 5538 4656 5539
rect 4786 5543 4792 5544
rect 4786 5539 4787 5543
rect 4791 5539 4792 5543
rect 4786 5538 4792 5539
rect 4922 5543 4928 5544
rect 4922 5539 4923 5543
rect 4927 5539 4928 5543
rect 4922 5538 4928 5539
rect 5058 5543 5064 5544
rect 5058 5539 5059 5543
rect 5063 5539 5064 5543
rect 5662 5540 5663 5544
rect 5667 5540 5668 5544
rect 5662 5539 5668 5540
rect 5058 5538 5064 5539
rect 4270 5528 4276 5529
rect 3838 5527 3844 5528
rect 3838 5523 3839 5527
rect 3843 5523 3844 5527
rect 4270 5524 4271 5528
rect 4275 5524 4276 5528
rect 4270 5523 4276 5524
rect 4406 5528 4412 5529
rect 4406 5524 4407 5528
rect 4411 5524 4412 5528
rect 4406 5523 4412 5524
rect 4542 5528 4548 5529
rect 4542 5524 4543 5528
rect 4547 5524 4548 5528
rect 4542 5523 4548 5524
rect 4678 5528 4684 5529
rect 4678 5524 4679 5528
rect 4683 5524 4684 5528
rect 4678 5523 4684 5524
rect 4814 5528 4820 5529
rect 4814 5524 4815 5528
rect 4819 5524 4820 5528
rect 4814 5523 4820 5524
rect 4950 5528 4956 5529
rect 4950 5524 4951 5528
rect 4955 5524 4956 5528
rect 4950 5523 4956 5524
rect 5086 5528 5092 5529
rect 5086 5524 5087 5528
rect 5091 5524 5092 5528
rect 5086 5523 5092 5524
rect 5662 5527 5668 5528
rect 5662 5523 5663 5527
rect 5667 5523 5668 5527
rect 3838 5522 3844 5523
rect 3840 5499 3842 5522
rect 4272 5499 4274 5523
rect 4408 5499 4410 5523
rect 4544 5499 4546 5523
rect 4680 5499 4682 5523
rect 4816 5499 4818 5523
rect 4952 5499 4954 5523
rect 5088 5499 5090 5523
rect 5662 5522 5668 5523
rect 5664 5499 5666 5522
rect 3839 5498 3843 5499
rect 3798 5496 3804 5497
rect 1974 5492 1975 5496
rect 1979 5492 1980 5496
rect 1974 5491 1980 5492
rect 1994 5495 2000 5496
rect 1994 5491 1995 5495
rect 1999 5491 2000 5495
rect 1994 5490 2000 5491
rect 2130 5495 2136 5496
rect 2130 5491 2131 5495
rect 2135 5491 2136 5495
rect 2130 5490 2136 5491
rect 2266 5495 2272 5496
rect 2266 5491 2267 5495
rect 2271 5491 2272 5495
rect 2266 5490 2272 5491
rect 2402 5495 2408 5496
rect 2402 5491 2403 5495
rect 2407 5491 2408 5495
rect 2402 5490 2408 5491
rect 2554 5495 2560 5496
rect 2554 5491 2555 5495
rect 2559 5491 2560 5495
rect 2554 5490 2560 5491
rect 2706 5495 2712 5496
rect 2706 5491 2707 5495
rect 2711 5491 2712 5495
rect 2706 5490 2712 5491
rect 2858 5495 2864 5496
rect 2858 5491 2859 5495
rect 2863 5491 2864 5495
rect 2858 5490 2864 5491
rect 3010 5495 3016 5496
rect 3010 5491 3011 5495
rect 3015 5491 3016 5495
rect 3010 5490 3016 5491
rect 3162 5495 3168 5496
rect 3162 5491 3163 5495
rect 3167 5491 3168 5495
rect 3162 5490 3168 5491
rect 3322 5495 3328 5496
rect 3322 5491 3323 5495
rect 3327 5491 3328 5495
rect 3322 5490 3328 5491
rect 3482 5495 3488 5496
rect 3482 5491 3483 5495
rect 3487 5491 3488 5495
rect 3798 5492 3799 5496
rect 3803 5492 3804 5496
rect 3839 5493 3843 5494
rect 4271 5498 4275 5499
rect 4271 5493 4275 5494
rect 4407 5498 4411 5499
rect 4407 5493 4411 5494
rect 4455 5498 4459 5499
rect 4455 5493 4459 5494
rect 4543 5498 4547 5499
rect 4543 5493 4547 5494
rect 4591 5498 4595 5499
rect 4591 5493 4595 5494
rect 4679 5498 4683 5499
rect 4679 5493 4683 5494
rect 4727 5498 4731 5499
rect 4727 5493 4731 5494
rect 4815 5498 4819 5499
rect 4815 5493 4819 5494
rect 4863 5498 4867 5499
rect 4863 5493 4867 5494
rect 4951 5498 4955 5499
rect 4951 5493 4955 5494
rect 5087 5498 5091 5499
rect 5087 5493 5091 5494
rect 5663 5498 5667 5499
rect 5663 5493 5667 5494
rect 3798 5491 3804 5492
rect 3482 5490 3488 5491
rect 111 5482 115 5483
rect 111 5477 115 5478
rect 783 5482 787 5483
rect 783 5477 787 5478
rect 863 5482 867 5483
rect 863 5477 867 5478
rect 919 5482 923 5483
rect 919 5477 923 5478
rect 999 5482 1003 5483
rect 999 5477 1003 5478
rect 1055 5482 1059 5483
rect 1055 5477 1059 5478
rect 1135 5482 1139 5483
rect 1135 5477 1139 5478
rect 1191 5482 1195 5483
rect 1191 5477 1195 5478
rect 1271 5482 1275 5483
rect 1271 5477 1275 5478
rect 1407 5482 1411 5483
rect 1407 5477 1411 5478
rect 1543 5482 1547 5483
rect 1543 5477 1547 5478
rect 1679 5482 1683 5483
rect 1679 5477 1683 5478
rect 1815 5482 1819 5483
rect 1815 5477 1819 5478
rect 1935 5482 1939 5483
rect 2022 5480 2028 5481
rect 1935 5477 1939 5478
rect 1974 5479 1980 5480
rect 112 5454 114 5477
rect 110 5453 116 5454
rect 864 5453 866 5477
rect 1000 5453 1002 5477
rect 1136 5453 1138 5477
rect 1272 5453 1274 5477
rect 1408 5453 1410 5477
rect 1544 5453 1546 5477
rect 1680 5453 1682 5477
rect 1816 5453 1818 5477
rect 1936 5454 1938 5477
rect 1974 5475 1975 5479
rect 1979 5475 1980 5479
rect 2022 5476 2023 5480
rect 2027 5476 2028 5480
rect 2022 5475 2028 5476
rect 2158 5480 2164 5481
rect 2158 5476 2159 5480
rect 2163 5476 2164 5480
rect 2158 5475 2164 5476
rect 2294 5480 2300 5481
rect 2294 5476 2295 5480
rect 2299 5476 2300 5480
rect 2294 5475 2300 5476
rect 2430 5480 2436 5481
rect 2430 5476 2431 5480
rect 2435 5476 2436 5480
rect 2430 5475 2436 5476
rect 2582 5480 2588 5481
rect 2582 5476 2583 5480
rect 2587 5476 2588 5480
rect 2582 5475 2588 5476
rect 2734 5480 2740 5481
rect 2734 5476 2735 5480
rect 2739 5476 2740 5480
rect 2734 5475 2740 5476
rect 2886 5480 2892 5481
rect 2886 5476 2887 5480
rect 2891 5476 2892 5480
rect 2886 5475 2892 5476
rect 3038 5480 3044 5481
rect 3038 5476 3039 5480
rect 3043 5476 3044 5480
rect 3038 5475 3044 5476
rect 3190 5480 3196 5481
rect 3190 5476 3191 5480
rect 3195 5476 3196 5480
rect 3190 5475 3196 5476
rect 3350 5480 3356 5481
rect 3350 5476 3351 5480
rect 3355 5476 3356 5480
rect 3350 5475 3356 5476
rect 3510 5480 3516 5481
rect 3510 5476 3511 5480
rect 3515 5476 3516 5480
rect 3510 5475 3516 5476
rect 3798 5479 3804 5480
rect 3798 5475 3799 5479
rect 3803 5475 3804 5479
rect 1974 5474 1980 5475
rect 1934 5453 1940 5454
rect 110 5449 111 5453
rect 115 5449 116 5453
rect 110 5448 116 5449
rect 862 5452 868 5453
rect 862 5448 863 5452
rect 867 5448 868 5452
rect 862 5447 868 5448
rect 998 5452 1004 5453
rect 998 5448 999 5452
rect 1003 5448 1004 5452
rect 998 5447 1004 5448
rect 1134 5452 1140 5453
rect 1134 5448 1135 5452
rect 1139 5448 1140 5452
rect 1134 5447 1140 5448
rect 1270 5452 1276 5453
rect 1270 5448 1271 5452
rect 1275 5448 1276 5452
rect 1270 5447 1276 5448
rect 1406 5452 1412 5453
rect 1406 5448 1407 5452
rect 1411 5448 1412 5452
rect 1406 5447 1412 5448
rect 1542 5452 1548 5453
rect 1542 5448 1543 5452
rect 1547 5448 1548 5452
rect 1542 5447 1548 5448
rect 1678 5452 1684 5453
rect 1678 5448 1679 5452
rect 1683 5448 1684 5452
rect 1678 5447 1684 5448
rect 1814 5452 1820 5453
rect 1814 5448 1815 5452
rect 1819 5448 1820 5452
rect 1934 5449 1935 5453
rect 1939 5449 1940 5453
rect 1934 5448 1940 5449
rect 1814 5447 1820 5448
rect 1976 5439 1978 5474
rect 2024 5439 2026 5475
rect 2160 5439 2162 5475
rect 2296 5439 2298 5475
rect 2432 5439 2434 5475
rect 2584 5439 2586 5475
rect 2736 5439 2738 5475
rect 2888 5439 2890 5475
rect 3040 5439 3042 5475
rect 3192 5439 3194 5475
rect 3352 5439 3354 5475
rect 3512 5439 3514 5475
rect 3798 5474 3804 5475
rect 3800 5439 3802 5474
rect 3840 5470 3842 5493
rect 3838 5469 3844 5470
rect 4456 5469 4458 5493
rect 4592 5469 4594 5493
rect 4728 5469 4730 5493
rect 4864 5469 4866 5493
rect 5664 5470 5666 5493
rect 5662 5469 5668 5470
rect 3838 5465 3839 5469
rect 3843 5465 3844 5469
rect 3838 5464 3844 5465
rect 4454 5468 4460 5469
rect 4454 5464 4455 5468
rect 4459 5464 4460 5468
rect 4454 5463 4460 5464
rect 4590 5468 4596 5469
rect 4590 5464 4591 5468
rect 4595 5464 4596 5468
rect 4590 5463 4596 5464
rect 4726 5468 4732 5469
rect 4726 5464 4727 5468
rect 4731 5464 4732 5468
rect 4726 5463 4732 5464
rect 4862 5468 4868 5469
rect 4862 5464 4863 5468
rect 4867 5464 4868 5468
rect 5662 5465 5663 5469
rect 5667 5465 5668 5469
rect 5662 5464 5668 5465
rect 4862 5463 4868 5464
rect 4426 5453 4432 5454
rect 3838 5452 3844 5453
rect 3838 5448 3839 5452
rect 3843 5448 3844 5452
rect 4426 5449 4427 5453
rect 4431 5449 4432 5453
rect 4426 5448 4432 5449
rect 4562 5453 4568 5454
rect 4562 5449 4563 5453
rect 4567 5449 4568 5453
rect 4562 5448 4568 5449
rect 4698 5453 4704 5454
rect 4698 5449 4699 5453
rect 4703 5449 4704 5453
rect 4698 5448 4704 5449
rect 4834 5453 4840 5454
rect 4834 5449 4835 5453
rect 4839 5449 4840 5453
rect 4834 5448 4840 5449
rect 5662 5452 5668 5453
rect 5662 5448 5663 5452
rect 5667 5448 5668 5452
rect 3838 5447 3844 5448
rect 1975 5438 1979 5439
rect 834 5437 840 5438
rect 110 5436 116 5437
rect 110 5432 111 5436
rect 115 5432 116 5436
rect 834 5433 835 5437
rect 839 5433 840 5437
rect 834 5432 840 5433
rect 970 5437 976 5438
rect 970 5433 971 5437
rect 975 5433 976 5437
rect 970 5432 976 5433
rect 1106 5437 1112 5438
rect 1106 5433 1107 5437
rect 1111 5433 1112 5437
rect 1106 5432 1112 5433
rect 1242 5437 1248 5438
rect 1242 5433 1243 5437
rect 1247 5433 1248 5437
rect 1242 5432 1248 5433
rect 1378 5437 1384 5438
rect 1378 5433 1379 5437
rect 1383 5433 1384 5437
rect 1378 5432 1384 5433
rect 1514 5437 1520 5438
rect 1514 5433 1515 5437
rect 1519 5433 1520 5437
rect 1514 5432 1520 5433
rect 1650 5437 1656 5438
rect 1650 5433 1651 5437
rect 1655 5433 1656 5437
rect 1650 5432 1656 5433
rect 1786 5437 1792 5438
rect 1786 5433 1787 5437
rect 1791 5433 1792 5437
rect 1786 5432 1792 5433
rect 1934 5436 1940 5437
rect 1934 5432 1935 5436
rect 1939 5432 1940 5436
rect 1975 5433 1979 5434
rect 2023 5438 2027 5439
rect 2023 5433 2027 5434
rect 2159 5438 2163 5439
rect 2159 5433 2163 5434
rect 2295 5438 2299 5439
rect 2295 5433 2299 5434
rect 2431 5438 2435 5439
rect 2431 5433 2435 5434
rect 2583 5438 2587 5439
rect 2583 5433 2587 5434
rect 2735 5438 2739 5439
rect 2735 5433 2739 5434
rect 2831 5438 2835 5439
rect 2831 5433 2835 5434
rect 2887 5438 2891 5439
rect 2887 5433 2891 5434
rect 2967 5438 2971 5439
rect 2967 5433 2971 5434
rect 3039 5438 3043 5439
rect 3039 5433 3043 5434
rect 3103 5438 3107 5439
rect 3103 5433 3107 5434
rect 3191 5438 3195 5439
rect 3191 5433 3195 5434
rect 3239 5438 3243 5439
rect 3239 5433 3243 5434
rect 3351 5438 3355 5439
rect 3351 5433 3355 5434
rect 3511 5438 3515 5439
rect 3511 5433 3515 5434
rect 3799 5438 3803 5439
rect 3799 5433 3803 5434
rect 110 5431 116 5432
rect 112 5371 114 5431
rect 836 5371 838 5432
rect 972 5371 974 5432
rect 1108 5371 1110 5432
rect 1244 5371 1246 5432
rect 1380 5371 1382 5432
rect 1516 5371 1518 5432
rect 1652 5371 1654 5432
rect 1788 5371 1790 5432
rect 1934 5431 1940 5432
rect 1936 5371 1938 5431
rect 1976 5410 1978 5433
rect 1974 5409 1980 5410
rect 2832 5409 2834 5433
rect 2968 5409 2970 5433
rect 3104 5409 3106 5433
rect 3240 5409 3242 5433
rect 3800 5410 3802 5433
rect 3798 5409 3804 5410
rect 1974 5405 1975 5409
rect 1979 5405 1980 5409
rect 1974 5404 1980 5405
rect 2830 5408 2836 5409
rect 2830 5404 2831 5408
rect 2835 5404 2836 5408
rect 2830 5403 2836 5404
rect 2966 5408 2972 5409
rect 2966 5404 2967 5408
rect 2971 5404 2972 5408
rect 2966 5403 2972 5404
rect 3102 5408 3108 5409
rect 3102 5404 3103 5408
rect 3107 5404 3108 5408
rect 3102 5403 3108 5404
rect 3238 5408 3244 5409
rect 3238 5404 3239 5408
rect 3243 5404 3244 5408
rect 3798 5405 3799 5409
rect 3803 5405 3804 5409
rect 3798 5404 3804 5405
rect 3238 5403 3244 5404
rect 2802 5393 2808 5394
rect 1974 5392 1980 5393
rect 1974 5388 1975 5392
rect 1979 5388 1980 5392
rect 2802 5389 2803 5393
rect 2807 5389 2808 5393
rect 2802 5388 2808 5389
rect 2938 5393 2944 5394
rect 2938 5389 2939 5393
rect 2943 5389 2944 5393
rect 2938 5388 2944 5389
rect 3074 5393 3080 5394
rect 3074 5389 3075 5393
rect 3079 5389 3080 5393
rect 3074 5388 3080 5389
rect 3210 5393 3216 5394
rect 3210 5389 3211 5393
rect 3215 5389 3216 5393
rect 3210 5388 3216 5389
rect 3798 5392 3804 5393
rect 3798 5388 3799 5392
rect 3803 5388 3804 5392
rect 1974 5387 1980 5388
rect 111 5370 115 5371
rect 111 5365 115 5366
rect 427 5370 431 5371
rect 427 5365 431 5366
rect 563 5370 567 5371
rect 563 5365 567 5366
rect 699 5370 703 5371
rect 699 5365 703 5366
rect 835 5370 839 5371
rect 835 5365 839 5366
rect 971 5370 975 5371
rect 971 5365 975 5366
rect 1107 5370 1111 5371
rect 1107 5365 1111 5366
rect 1243 5370 1247 5371
rect 1243 5365 1247 5366
rect 1379 5370 1383 5371
rect 1379 5365 1383 5366
rect 1515 5370 1519 5371
rect 1515 5365 1519 5366
rect 1651 5370 1655 5371
rect 1651 5365 1655 5366
rect 1787 5370 1791 5371
rect 1787 5365 1791 5366
rect 1935 5370 1939 5371
rect 1935 5365 1939 5366
rect 112 5305 114 5365
rect 110 5304 116 5305
rect 428 5304 430 5365
rect 564 5304 566 5365
rect 700 5304 702 5365
rect 836 5304 838 5365
rect 972 5304 974 5365
rect 1108 5304 1110 5365
rect 1244 5304 1246 5365
rect 1380 5304 1382 5365
rect 1516 5304 1518 5365
rect 1652 5304 1654 5365
rect 1788 5304 1790 5365
rect 1936 5305 1938 5365
rect 1934 5304 1940 5305
rect 110 5300 111 5304
rect 115 5300 116 5304
rect 110 5299 116 5300
rect 426 5303 432 5304
rect 426 5299 427 5303
rect 431 5299 432 5303
rect 426 5298 432 5299
rect 562 5303 568 5304
rect 562 5299 563 5303
rect 567 5299 568 5303
rect 562 5298 568 5299
rect 698 5303 704 5304
rect 698 5299 699 5303
rect 703 5299 704 5303
rect 698 5298 704 5299
rect 834 5303 840 5304
rect 834 5299 835 5303
rect 839 5299 840 5303
rect 834 5298 840 5299
rect 970 5303 976 5304
rect 970 5299 971 5303
rect 975 5299 976 5303
rect 970 5298 976 5299
rect 1106 5303 1112 5304
rect 1106 5299 1107 5303
rect 1111 5299 1112 5303
rect 1106 5298 1112 5299
rect 1242 5303 1248 5304
rect 1242 5299 1243 5303
rect 1247 5299 1248 5303
rect 1242 5298 1248 5299
rect 1378 5303 1384 5304
rect 1378 5299 1379 5303
rect 1383 5299 1384 5303
rect 1378 5298 1384 5299
rect 1514 5303 1520 5304
rect 1514 5299 1515 5303
rect 1519 5299 1520 5303
rect 1514 5298 1520 5299
rect 1650 5303 1656 5304
rect 1650 5299 1651 5303
rect 1655 5299 1656 5303
rect 1650 5298 1656 5299
rect 1786 5303 1792 5304
rect 1786 5299 1787 5303
rect 1791 5299 1792 5303
rect 1934 5300 1935 5304
rect 1939 5300 1940 5304
rect 1934 5299 1940 5300
rect 1786 5298 1792 5299
rect 1976 5291 1978 5387
rect 2804 5291 2806 5388
rect 2940 5291 2942 5388
rect 3076 5291 3078 5388
rect 3212 5291 3214 5388
rect 3798 5387 3804 5388
rect 3840 5387 3842 5447
rect 4428 5387 4430 5448
rect 4564 5387 4566 5448
rect 4700 5387 4702 5448
rect 4836 5387 4838 5448
rect 5662 5447 5668 5448
rect 5664 5387 5666 5447
rect 3800 5291 3802 5387
rect 3839 5386 3843 5387
rect 3839 5381 3843 5382
rect 4283 5386 4287 5387
rect 4283 5381 4287 5382
rect 4427 5386 4431 5387
rect 4427 5381 4431 5382
rect 4483 5386 4487 5387
rect 4483 5381 4487 5382
rect 4563 5386 4567 5387
rect 4563 5381 4567 5382
rect 4699 5386 4703 5387
rect 4699 5381 4703 5382
rect 4835 5386 4839 5387
rect 4835 5381 4839 5382
rect 4931 5386 4935 5387
rect 4931 5381 4935 5382
rect 5171 5386 5175 5387
rect 5171 5381 5175 5382
rect 5419 5386 5423 5387
rect 5419 5381 5423 5382
rect 5663 5386 5667 5387
rect 5663 5381 5667 5382
rect 3840 5321 3842 5381
rect 3838 5320 3844 5321
rect 4284 5320 4286 5381
rect 4484 5320 4486 5381
rect 4700 5320 4702 5381
rect 4932 5320 4934 5381
rect 5172 5320 5174 5381
rect 5420 5320 5422 5381
rect 5664 5321 5666 5381
rect 5662 5320 5668 5321
rect 3838 5316 3839 5320
rect 3843 5316 3844 5320
rect 3838 5315 3844 5316
rect 4282 5319 4288 5320
rect 4282 5315 4283 5319
rect 4287 5315 4288 5319
rect 4282 5314 4288 5315
rect 4482 5319 4488 5320
rect 4482 5315 4483 5319
rect 4487 5315 4488 5319
rect 4482 5314 4488 5315
rect 4698 5319 4704 5320
rect 4698 5315 4699 5319
rect 4703 5315 4704 5319
rect 4698 5314 4704 5315
rect 4930 5319 4936 5320
rect 4930 5315 4931 5319
rect 4935 5315 4936 5319
rect 4930 5314 4936 5315
rect 5170 5319 5176 5320
rect 5170 5315 5171 5319
rect 5175 5315 5176 5319
rect 5170 5314 5176 5315
rect 5418 5319 5424 5320
rect 5418 5315 5419 5319
rect 5423 5315 5424 5319
rect 5662 5316 5663 5320
rect 5667 5316 5668 5320
rect 5662 5315 5668 5316
rect 5418 5314 5424 5315
rect 4310 5304 4316 5305
rect 3838 5303 3844 5304
rect 3838 5299 3839 5303
rect 3843 5299 3844 5303
rect 4310 5300 4311 5304
rect 4315 5300 4316 5304
rect 4310 5299 4316 5300
rect 4510 5304 4516 5305
rect 4510 5300 4511 5304
rect 4515 5300 4516 5304
rect 4510 5299 4516 5300
rect 4726 5304 4732 5305
rect 4726 5300 4727 5304
rect 4731 5300 4732 5304
rect 4726 5299 4732 5300
rect 4958 5304 4964 5305
rect 4958 5300 4959 5304
rect 4963 5300 4964 5304
rect 4958 5299 4964 5300
rect 5198 5304 5204 5305
rect 5198 5300 5199 5304
rect 5203 5300 5204 5304
rect 5198 5299 5204 5300
rect 5446 5304 5452 5305
rect 5446 5300 5447 5304
rect 5451 5300 5452 5304
rect 5446 5299 5452 5300
rect 5662 5303 5668 5304
rect 5662 5299 5663 5303
rect 5667 5299 5668 5303
rect 3838 5298 3844 5299
rect 1975 5290 1979 5291
rect 454 5288 460 5289
rect 110 5287 116 5288
rect 110 5283 111 5287
rect 115 5283 116 5287
rect 454 5284 455 5288
rect 459 5284 460 5288
rect 454 5283 460 5284
rect 590 5288 596 5289
rect 590 5284 591 5288
rect 595 5284 596 5288
rect 590 5283 596 5284
rect 726 5288 732 5289
rect 726 5284 727 5288
rect 731 5284 732 5288
rect 726 5283 732 5284
rect 862 5288 868 5289
rect 862 5284 863 5288
rect 867 5284 868 5288
rect 862 5283 868 5284
rect 998 5288 1004 5289
rect 998 5284 999 5288
rect 1003 5284 1004 5288
rect 998 5283 1004 5284
rect 1134 5288 1140 5289
rect 1134 5284 1135 5288
rect 1139 5284 1140 5288
rect 1134 5283 1140 5284
rect 1270 5288 1276 5289
rect 1270 5284 1271 5288
rect 1275 5284 1276 5288
rect 1270 5283 1276 5284
rect 1406 5288 1412 5289
rect 1406 5284 1407 5288
rect 1411 5284 1412 5288
rect 1406 5283 1412 5284
rect 1542 5288 1548 5289
rect 1542 5284 1543 5288
rect 1547 5284 1548 5288
rect 1542 5283 1548 5284
rect 1678 5288 1684 5289
rect 1678 5284 1679 5288
rect 1683 5284 1684 5288
rect 1678 5283 1684 5284
rect 1814 5288 1820 5289
rect 1814 5284 1815 5288
rect 1819 5284 1820 5288
rect 1814 5283 1820 5284
rect 1934 5287 1940 5288
rect 1934 5283 1935 5287
rect 1939 5283 1940 5287
rect 1975 5285 1979 5286
rect 1995 5290 1999 5291
rect 1995 5285 1999 5286
rect 2219 5290 2223 5291
rect 2219 5285 2223 5286
rect 2467 5290 2471 5291
rect 2467 5285 2471 5286
rect 2715 5290 2719 5291
rect 2715 5285 2719 5286
rect 2803 5290 2807 5291
rect 2803 5285 2807 5286
rect 2939 5290 2943 5291
rect 2939 5285 2943 5286
rect 2971 5290 2975 5291
rect 2971 5285 2975 5286
rect 3075 5290 3079 5291
rect 3075 5285 3079 5286
rect 3211 5290 3215 5291
rect 3211 5285 3215 5286
rect 3799 5290 3803 5291
rect 3799 5285 3803 5286
rect 110 5282 116 5283
rect 112 5259 114 5282
rect 456 5259 458 5283
rect 592 5259 594 5283
rect 728 5259 730 5283
rect 864 5259 866 5283
rect 1000 5259 1002 5283
rect 1136 5259 1138 5283
rect 1272 5259 1274 5283
rect 1408 5259 1410 5283
rect 1544 5259 1546 5283
rect 1680 5259 1682 5283
rect 1816 5259 1818 5283
rect 1934 5282 1940 5283
rect 1936 5259 1938 5282
rect 111 5258 115 5259
rect 111 5253 115 5254
rect 455 5258 459 5259
rect 455 5253 459 5254
rect 591 5258 595 5259
rect 591 5253 595 5254
rect 727 5258 731 5259
rect 727 5253 731 5254
rect 863 5258 867 5259
rect 863 5253 867 5254
rect 999 5258 1003 5259
rect 999 5253 1003 5254
rect 1135 5258 1139 5259
rect 1135 5253 1139 5254
rect 1271 5258 1275 5259
rect 1271 5253 1275 5254
rect 1407 5258 1411 5259
rect 1407 5253 1411 5254
rect 1543 5258 1547 5259
rect 1543 5253 1547 5254
rect 1679 5258 1683 5259
rect 1679 5253 1683 5254
rect 1815 5258 1819 5259
rect 1815 5253 1819 5254
rect 1935 5258 1939 5259
rect 1935 5253 1939 5254
rect 112 5230 114 5253
rect 110 5229 116 5230
rect 456 5229 458 5253
rect 592 5229 594 5253
rect 728 5229 730 5253
rect 864 5229 866 5253
rect 1000 5229 1002 5253
rect 1136 5229 1138 5253
rect 1272 5229 1274 5253
rect 1408 5229 1410 5253
rect 1544 5229 1546 5253
rect 1680 5229 1682 5253
rect 1816 5229 1818 5253
rect 1936 5230 1938 5253
rect 1934 5229 1940 5230
rect 110 5225 111 5229
rect 115 5225 116 5229
rect 110 5224 116 5225
rect 454 5228 460 5229
rect 454 5224 455 5228
rect 459 5224 460 5228
rect 454 5223 460 5224
rect 590 5228 596 5229
rect 590 5224 591 5228
rect 595 5224 596 5228
rect 590 5223 596 5224
rect 726 5228 732 5229
rect 726 5224 727 5228
rect 731 5224 732 5228
rect 726 5223 732 5224
rect 862 5228 868 5229
rect 862 5224 863 5228
rect 867 5224 868 5228
rect 862 5223 868 5224
rect 998 5228 1004 5229
rect 998 5224 999 5228
rect 1003 5224 1004 5228
rect 998 5223 1004 5224
rect 1134 5228 1140 5229
rect 1134 5224 1135 5228
rect 1139 5224 1140 5228
rect 1134 5223 1140 5224
rect 1270 5228 1276 5229
rect 1270 5224 1271 5228
rect 1275 5224 1276 5228
rect 1270 5223 1276 5224
rect 1406 5228 1412 5229
rect 1406 5224 1407 5228
rect 1411 5224 1412 5228
rect 1406 5223 1412 5224
rect 1542 5228 1548 5229
rect 1542 5224 1543 5228
rect 1547 5224 1548 5228
rect 1542 5223 1548 5224
rect 1678 5228 1684 5229
rect 1678 5224 1679 5228
rect 1683 5224 1684 5228
rect 1678 5223 1684 5224
rect 1814 5228 1820 5229
rect 1814 5224 1815 5228
rect 1819 5224 1820 5228
rect 1934 5225 1935 5229
rect 1939 5225 1940 5229
rect 1976 5225 1978 5285
rect 1934 5224 1940 5225
rect 1974 5224 1980 5225
rect 1996 5224 1998 5285
rect 2220 5224 2222 5285
rect 2468 5224 2470 5285
rect 2716 5224 2718 5285
rect 2972 5224 2974 5285
rect 3800 5225 3802 5285
rect 3840 5247 3842 5298
rect 4312 5247 4314 5299
rect 4512 5247 4514 5299
rect 4728 5247 4730 5299
rect 4960 5247 4962 5299
rect 5200 5247 5202 5299
rect 5448 5247 5450 5299
rect 5662 5298 5668 5299
rect 5664 5247 5666 5298
rect 3839 5246 3843 5247
rect 3839 5241 3843 5242
rect 3887 5246 3891 5247
rect 3887 5241 3891 5242
rect 4023 5246 4027 5247
rect 4023 5241 4027 5242
rect 4159 5246 4163 5247
rect 4159 5241 4163 5242
rect 4295 5246 4299 5247
rect 4295 5241 4299 5242
rect 4311 5246 4315 5247
rect 4311 5241 4315 5242
rect 4431 5246 4435 5247
rect 4431 5241 4435 5242
rect 4511 5246 4515 5247
rect 4511 5241 4515 5242
rect 4567 5246 4571 5247
rect 4567 5241 4571 5242
rect 4703 5246 4707 5247
rect 4703 5241 4707 5242
rect 4727 5246 4731 5247
rect 4727 5241 4731 5242
rect 4839 5246 4843 5247
rect 4839 5241 4843 5242
rect 4959 5246 4963 5247
rect 4959 5241 4963 5242
rect 4991 5246 4995 5247
rect 4991 5241 4995 5242
rect 5151 5246 5155 5247
rect 5151 5241 5155 5242
rect 5199 5246 5203 5247
rect 5199 5241 5203 5242
rect 5319 5246 5323 5247
rect 5319 5241 5323 5242
rect 5447 5246 5451 5247
rect 5447 5241 5451 5242
rect 5495 5246 5499 5247
rect 5495 5241 5499 5242
rect 5663 5246 5667 5247
rect 5663 5241 5667 5242
rect 3798 5224 3804 5225
rect 1814 5223 1820 5224
rect 1974 5220 1975 5224
rect 1979 5220 1980 5224
rect 1974 5219 1980 5220
rect 1994 5223 2000 5224
rect 1994 5219 1995 5223
rect 1999 5219 2000 5223
rect 1994 5218 2000 5219
rect 2218 5223 2224 5224
rect 2218 5219 2219 5223
rect 2223 5219 2224 5223
rect 2218 5218 2224 5219
rect 2466 5223 2472 5224
rect 2466 5219 2467 5223
rect 2471 5219 2472 5223
rect 2466 5218 2472 5219
rect 2714 5223 2720 5224
rect 2714 5219 2715 5223
rect 2719 5219 2720 5223
rect 2714 5218 2720 5219
rect 2970 5223 2976 5224
rect 2970 5219 2971 5223
rect 2975 5219 2976 5223
rect 3798 5220 3799 5224
rect 3803 5220 3804 5224
rect 3798 5219 3804 5220
rect 2970 5218 2976 5219
rect 3840 5218 3842 5241
rect 3838 5217 3844 5218
rect 3888 5217 3890 5241
rect 4024 5217 4026 5241
rect 4160 5217 4162 5241
rect 4296 5217 4298 5241
rect 4432 5217 4434 5241
rect 4568 5217 4570 5241
rect 4704 5217 4706 5241
rect 4840 5217 4842 5241
rect 4992 5217 4994 5241
rect 5152 5217 5154 5241
rect 5320 5217 5322 5241
rect 5496 5217 5498 5241
rect 5664 5218 5666 5241
rect 5662 5217 5668 5218
rect 426 5213 432 5214
rect 110 5212 116 5213
rect 110 5208 111 5212
rect 115 5208 116 5212
rect 426 5209 427 5213
rect 431 5209 432 5213
rect 426 5208 432 5209
rect 562 5213 568 5214
rect 562 5209 563 5213
rect 567 5209 568 5213
rect 562 5208 568 5209
rect 698 5213 704 5214
rect 698 5209 699 5213
rect 703 5209 704 5213
rect 698 5208 704 5209
rect 834 5213 840 5214
rect 834 5209 835 5213
rect 839 5209 840 5213
rect 834 5208 840 5209
rect 970 5213 976 5214
rect 970 5209 971 5213
rect 975 5209 976 5213
rect 970 5208 976 5209
rect 1106 5213 1112 5214
rect 1106 5209 1107 5213
rect 1111 5209 1112 5213
rect 1106 5208 1112 5209
rect 1242 5213 1248 5214
rect 1242 5209 1243 5213
rect 1247 5209 1248 5213
rect 1242 5208 1248 5209
rect 1378 5213 1384 5214
rect 1378 5209 1379 5213
rect 1383 5209 1384 5213
rect 1378 5208 1384 5209
rect 1514 5213 1520 5214
rect 1514 5209 1515 5213
rect 1519 5209 1520 5213
rect 1514 5208 1520 5209
rect 1650 5213 1656 5214
rect 1650 5209 1651 5213
rect 1655 5209 1656 5213
rect 1650 5208 1656 5209
rect 1786 5213 1792 5214
rect 3838 5213 3839 5217
rect 3843 5213 3844 5217
rect 1786 5209 1787 5213
rect 1791 5209 1792 5213
rect 1786 5208 1792 5209
rect 1934 5212 1940 5213
rect 3838 5212 3844 5213
rect 3886 5216 3892 5217
rect 3886 5212 3887 5216
rect 3891 5212 3892 5216
rect 1934 5208 1935 5212
rect 1939 5208 1940 5212
rect 3886 5211 3892 5212
rect 4022 5216 4028 5217
rect 4022 5212 4023 5216
rect 4027 5212 4028 5216
rect 4022 5211 4028 5212
rect 4158 5216 4164 5217
rect 4158 5212 4159 5216
rect 4163 5212 4164 5216
rect 4158 5211 4164 5212
rect 4294 5216 4300 5217
rect 4294 5212 4295 5216
rect 4299 5212 4300 5216
rect 4294 5211 4300 5212
rect 4430 5216 4436 5217
rect 4430 5212 4431 5216
rect 4435 5212 4436 5216
rect 4430 5211 4436 5212
rect 4566 5216 4572 5217
rect 4566 5212 4567 5216
rect 4571 5212 4572 5216
rect 4566 5211 4572 5212
rect 4702 5216 4708 5217
rect 4702 5212 4703 5216
rect 4707 5212 4708 5216
rect 4702 5211 4708 5212
rect 4838 5216 4844 5217
rect 4838 5212 4839 5216
rect 4843 5212 4844 5216
rect 4838 5211 4844 5212
rect 4990 5216 4996 5217
rect 4990 5212 4991 5216
rect 4995 5212 4996 5216
rect 4990 5211 4996 5212
rect 5150 5216 5156 5217
rect 5150 5212 5151 5216
rect 5155 5212 5156 5216
rect 5150 5211 5156 5212
rect 5318 5216 5324 5217
rect 5318 5212 5319 5216
rect 5323 5212 5324 5216
rect 5318 5211 5324 5212
rect 5494 5216 5500 5217
rect 5494 5212 5495 5216
rect 5499 5212 5500 5216
rect 5662 5213 5663 5217
rect 5667 5213 5668 5217
rect 5662 5212 5668 5213
rect 5494 5211 5500 5212
rect 2022 5208 2028 5209
rect 110 5207 116 5208
rect 112 5131 114 5207
rect 428 5131 430 5208
rect 564 5131 566 5208
rect 700 5131 702 5208
rect 836 5131 838 5208
rect 972 5131 974 5208
rect 1108 5131 1110 5208
rect 1244 5131 1246 5208
rect 1380 5131 1382 5208
rect 1516 5131 1518 5208
rect 1652 5131 1654 5208
rect 1788 5131 1790 5208
rect 1934 5207 1940 5208
rect 1974 5207 1980 5208
rect 1936 5131 1938 5207
rect 1974 5203 1975 5207
rect 1979 5203 1980 5207
rect 2022 5204 2023 5208
rect 2027 5204 2028 5208
rect 2022 5203 2028 5204
rect 2246 5208 2252 5209
rect 2246 5204 2247 5208
rect 2251 5204 2252 5208
rect 2246 5203 2252 5204
rect 2494 5208 2500 5209
rect 2494 5204 2495 5208
rect 2499 5204 2500 5208
rect 2494 5203 2500 5204
rect 2742 5208 2748 5209
rect 2742 5204 2743 5208
rect 2747 5204 2748 5208
rect 2742 5203 2748 5204
rect 2998 5208 3004 5209
rect 2998 5204 2999 5208
rect 3003 5204 3004 5208
rect 2998 5203 3004 5204
rect 3798 5207 3804 5208
rect 3798 5203 3799 5207
rect 3803 5203 3804 5207
rect 1974 5202 1980 5203
rect 1976 5175 1978 5202
rect 2024 5175 2026 5203
rect 2248 5175 2250 5203
rect 2496 5175 2498 5203
rect 2744 5175 2746 5203
rect 3000 5175 3002 5203
rect 3798 5202 3804 5203
rect 3800 5175 3802 5202
rect 3858 5201 3864 5202
rect 3838 5200 3844 5201
rect 3838 5196 3839 5200
rect 3843 5196 3844 5200
rect 3858 5197 3859 5201
rect 3863 5197 3864 5201
rect 3858 5196 3864 5197
rect 3994 5201 4000 5202
rect 3994 5197 3995 5201
rect 3999 5197 4000 5201
rect 3994 5196 4000 5197
rect 4130 5201 4136 5202
rect 4130 5197 4131 5201
rect 4135 5197 4136 5201
rect 4130 5196 4136 5197
rect 4266 5201 4272 5202
rect 4266 5197 4267 5201
rect 4271 5197 4272 5201
rect 4266 5196 4272 5197
rect 4402 5201 4408 5202
rect 4402 5197 4403 5201
rect 4407 5197 4408 5201
rect 4402 5196 4408 5197
rect 4538 5201 4544 5202
rect 4538 5197 4539 5201
rect 4543 5197 4544 5201
rect 4538 5196 4544 5197
rect 4674 5201 4680 5202
rect 4674 5197 4675 5201
rect 4679 5197 4680 5201
rect 4674 5196 4680 5197
rect 4810 5201 4816 5202
rect 4810 5197 4811 5201
rect 4815 5197 4816 5201
rect 4810 5196 4816 5197
rect 4962 5201 4968 5202
rect 4962 5197 4963 5201
rect 4967 5197 4968 5201
rect 4962 5196 4968 5197
rect 5122 5201 5128 5202
rect 5122 5197 5123 5201
rect 5127 5197 5128 5201
rect 5122 5196 5128 5197
rect 5290 5201 5296 5202
rect 5290 5197 5291 5201
rect 5295 5197 5296 5201
rect 5290 5196 5296 5197
rect 5466 5201 5472 5202
rect 5466 5197 5467 5201
rect 5471 5197 5472 5201
rect 5466 5196 5472 5197
rect 5662 5200 5668 5201
rect 5662 5196 5663 5200
rect 5667 5196 5668 5200
rect 3838 5195 3844 5196
rect 1975 5174 1979 5175
rect 1975 5169 1979 5170
rect 2023 5174 2027 5175
rect 2023 5169 2027 5170
rect 2159 5174 2163 5175
rect 2159 5169 2163 5170
rect 2247 5174 2251 5175
rect 2247 5169 2251 5170
rect 2295 5174 2299 5175
rect 2295 5169 2299 5170
rect 2431 5174 2435 5175
rect 2431 5169 2435 5170
rect 2495 5174 2499 5175
rect 2495 5169 2499 5170
rect 2567 5174 2571 5175
rect 2567 5169 2571 5170
rect 2703 5174 2707 5175
rect 2703 5169 2707 5170
rect 2743 5174 2747 5175
rect 2743 5169 2747 5170
rect 2839 5174 2843 5175
rect 2839 5169 2843 5170
rect 2975 5174 2979 5175
rect 2975 5169 2979 5170
rect 2999 5174 3003 5175
rect 2999 5169 3003 5170
rect 3111 5174 3115 5175
rect 3111 5169 3115 5170
rect 3247 5174 3251 5175
rect 3247 5169 3251 5170
rect 3391 5174 3395 5175
rect 3391 5169 3395 5170
rect 3543 5174 3547 5175
rect 3543 5169 3547 5170
rect 3679 5174 3683 5175
rect 3679 5169 3683 5170
rect 3799 5174 3803 5175
rect 3799 5169 3803 5170
rect 1976 5146 1978 5169
rect 1974 5145 1980 5146
rect 2024 5145 2026 5169
rect 2160 5145 2162 5169
rect 2296 5145 2298 5169
rect 2432 5145 2434 5169
rect 2568 5145 2570 5169
rect 2704 5145 2706 5169
rect 2840 5145 2842 5169
rect 2976 5145 2978 5169
rect 3112 5145 3114 5169
rect 3248 5145 3250 5169
rect 3392 5145 3394 5169
rect 3544 5145 3546 5169
rect 3680 5145 3682 5169
rect 3800 5146 3802 5169
rect 3798 5145 3804 5146
rect 1974 5141 1975 5145
rect 1979 5141 1980 5145
rect 1974 5140 1980 5141
rect 2022 5144 2028 5145
rect 2022 5140 2023 5144
rect 2027 5140 2028 5144
rect 2022 5139 2028 5140
rect 2158 5144 2164 5145
rect 2158 5140 2159 5144
rect 2163 5140 2164 5144
rect 2158 5139 2164 5140
rect 2294 5144 2300 5145
rect 2294 5140 2295 5144
rect 2299 5140 2300 5144
rect 2294 5139 2300 5140
rect 2430 5144 2436 5145
rect 2430 5140 2431 5144
rect 2435 5140 2436 5144
rect 2430 5139 2436 5140
rect 2566 5144 2572 5145
rect 2566 5140 2567 5144
rect 2571 5140 2572 5144
rect 2566 5139 2572 5140
rect 2702 5144 2708 5145
rect 2702 5140 2703 5144
rect 2707 5140 2708 5144
rect 2702 5139 2708 5140
rect 2838 5144 2844 5145
rect 2838 5140 2839 5144
rect 2843 5140 2844 5144
rect 2838 5139 2844 5140
rect 2974 5144 2980 5145
rect 2974 5140 2975 5144
rect 2979 5140 2980 5144
rect 2974 5139 2980 5140
rect 3110 5144 3116 5145
rect 3110 5140 3111 5144
rect 3115 5140 3116 5144
rect 3110 5139 3116 5140
rect 3246 5144 3252 5145
rect 3246 5140 3247 5144
rect 3251 5140 3252 5144
rect 3246 5139 3252 5140
rect 3390 5144 3396 5145
rect 3390 5140 3391 5144
rect 3395 5140 3396 5144
rect 3390 5139 3396 5140
rect 3542 5144 3548 5145
rect 3542 5140 3543 5144
rect 3547 5140 3548 5144
rect 3542 5139 3548 5140
rect 3678 5144 3684 5145
rect 3678 5140 3679 5144
rect 3683 5140 3684 5144
rect 3798 5141 3799 5145
rect 3803 5141 3804 5145
rect 3798 5140 3804 5141
rect 3678 5139 3684 5140
rect 3840 5135 3842 5195
rect 3860 5135 3862 5196
rect 3996 5135 3998 5196
rect 4132 5135 4134 5196
rect 4268 5135 4270 5196
rect 4404 5135 4406 5196
rect 4540 5135 4542 5196
rect 4676 5135 4678 5196
rect 4812 5135 4814 5196
rect 4964 5135 4966 5196
rect 5124 5135 5126 5196
rect 5292 5135 5294 5196
rect 5468 5135 5470 5196
rect 5662 5195 5668 5196
rect 5664 5135 5666 5195
rect 3839 5134 3843 5135
rect 111 5130 115 5131
rect 111 5125 115 5126
rect 267 5130 271 5131
rect 267 5125 271 5126
rect 403 5130 407 5131
rect 403 5125 407 5126
rect 427 5130 431 5131
rect 427 5125 431 5126
rect 539 5130 543 5131
rect 539 5125 543 5126
rect 563 5130 567 5131
rect 563 5125 567 5126
rect 675 5130 679 5131
rect 675 5125 679 5126
rect 699 5130 703 5131
rect 699 5125 703 5126
rect 811 5130 815 5131
rect 811 5125 815 5126
rect 835 5130 839 5131
rect 835 5125 839 5126
rect 947 5130 951 5131
rect 947 5125 951 5126
rect 971 5130 975 5131
rect 971 5125 975 5126
rect 1107 5130 1111 5131
rect 1107 5125 1111 5126
rect 1243 5130 1247 5131
rect 1243 5125 1247 5126
rect 1379 5130 1383 5131
rect 1379 5125 1383 5126
rect 1515 5130 1519 5131
rect 1515 5125 1519 5126
rect 1651 5130 1655 5131
rect 1651 5125 1655 5126
rect 1787 5130 1791 5131
rect 1787 5125 1791 5126
rect 1935 5130 1939 5131
rect 1994 5129 2000 5130
rect 1935 5125 1939 5126
rect 1974 5128 1980 5129
rect 112 5065 114 5125
rect 110 5064 116 5065
rect 268 5064 270 5125
rect 404 5064 406 5125
rect 540 5064 542 5125
rect 676 5064 678 5125
rect 812 5064 814 5125
rect 948 5064 950 5125
rect 1936 5065 1938 5125
rect 1974 5124 1975 5128
rect 1979 5124 1980 5128
rect 1994 5125 1995 5129
rect 1999 5125 2000 5129
rect 1994 5124 2000 5125
rect 2130 5129 2136 5130
rect 2130 5125 2131 5129
rect 2135 5125 2136 5129
rect 2130 5124 2136 5125
rect 2266 5129 2272 5130
rect 2266 5125 2267 5129
rect 2271 5125 2272 5129
rect 2266 5124 2272 5125
rect 2402 5129 2408 5130
rect 2402 5125 2403 5129
rect 2407 5125 2408 5129
rect 2402 5124 2408 5125
rect 2538 5129 2544 5130
rect 2538 5125 2539 5129
rect 2543 5125 2544 5129
rect 2538 5124 2544 5125
rect 2674 5129 2680 5130
rect 2674 5125 2675 5129
rect 2679 5125 2680 5129
rect 2674 5124 2680 5125
rect 2810 5129 2816 5130
rect 2810 5125 2811 5129
rect 2815 5125 2816 5129
rect 2810 5124 2816 5125
rect 2946 5129 2952 5130
rect 2946 5125 2947 5129
rect 2951 5125 2952 5129
rect 2946 5124 2952 5125
rect 3082 5129 3088 5130
rect 3082 5125 3083 5129
rect 3087 5125 3088 5129
rect 3082 5124 3088 5125
rect 3218 5129 3224 5130
rect 3218 5125 3219 5129
rect 3223 5125 3224 5129
rect 3218 5124 3224 5125
rect 3362 5129 3368 5130
rect 3362 5125 3363 5129
rect 3367 5125 3368 5129
rect 3362 5124 3368 5125
rect 3514 5129 3520 5130
rect 3514 5125 3515 5129
rect 3519 5125 3520 5129
rect 3514 5124 3520 5125
rect 3650 5129 3656 5130
rect 3839 5129 3843 5130
rect 3859 5134 3863 5135
rect 3859 5129 3863 5130
rect 3979 5134 3983 5135
rect 3979 5129 3983 5130
rect 3995 5134 3999 5135
rect 3995 5129 3999 5130
rect 4131 5134 4135 5135
rect 4131 5129 4135 5130
rect 4267 5134 4271 5135
rect 4267 5129 4271 5130
rect 4275 5134 4279 5135
rect 4275 5129 4279 5130
rect 4403 5134 4407 5135
rect 4403 5129 4407 5130
rect 4539 5134 4543 5135
rect 4539 5129 4543 5130
rect 4579 5134 4583 5135
rect 4579 5129 4583 5130
rect 4675 5134 4679 5135
rect 4675 5129 4679 5130
rect 4811 5134 4815 5135
rect 4811 5129 4815 5130
rect 4883 5134 4887 5135
rect 4883 5129 4887 5130
rect 4963 5134 4967 5135
rect 4963 5129 4967 5130
rect 5123 5134 5127 5135
rect 5123 5129 5127 5130
rect 5195 5134 5199 5135
rect 5195 5129 5199 5130
rect 5291 5134 5295 5135
rect 5291 5129 5295 5130
rect 5467 5134 5471 5135
rect 5467 5129 5471 5130
rect 5515 5134 5519 5135
rect 5515 5129 5519 5130
rect 5663 5134 5667 5135
rect 5663 5129 5667 5130
rect 3650 5125 3651 5129
rect 3655 5125 3656 5129
rect 3650 5124 3656 5125
rect 3798 5128 3804 5129
rect 3798 5124 3799 5128
rect 3803 5124 3804 5128
rect 1974 5123 1980 5124
rect 1934 5064 1940 5065
rect 110 5060 111 5064
rect 115 5060 116 5064
rect 110 5059 116 5060
rect 266 5063 272 5064
rect 266 5059 267 5063
rect 271 5059 272 5063
rect 266 5058 272 5059
rect 402 5063 408 5064
rect 402 5059 403 5063
rect 407 5059 408 5063
rect 402 5058 408 5059
rect 538 5063 544 5064
rect 538 5059 539 5063
rect 543 5059 544 5063
rect 538 5058 544 5059
rect 674 5063 680 5064
rect 674 5059 675 5063
rect 679 5059 680 5063
rect 674 5058 680 5059
rect 810 5063 816 5064
rect 810 5059 811 5063
rect 815 5059 816 5063
rect 810 5058 816 5059
rect 946 5063 952 5064
rect 946 5059 947 5063
rect 951 5059 952 5063
rect 1934 5060 1935 5064
rect 1939 5060 1940 5064
rect 1976 5063 1978 5123
rect 1996 5063 1998 5124
rect 2132 5063 2134 5124
rect 2268 5063 2270 5124
rect 2404 5063 2406 5124
rect 2540 5063 2542 5124
rect 2676 5063 2678 5124
rect 2812 5063 2814 5124
rect 2948 5063 2950 5124
rect 3084 5063 3086 5124
rect 3220 5063 3222 5124
rect 3364 5063 3366 5124
rect 3516 5063 3518 5124
rect 3652 5063 3654 5124
rect 3798 5123 3804 5124
rect 3800 5063 3802 5123
rect 3840 5069 3842 5129
rect 3838 5068 3844 5069
rect 3980 5068 3982 5129
rect 4276 5068 4278 5129
rect 4580 5068 4582 5129
rect 4884 5068 4886 5129
rect 5196 5068 5198 5129
rect 5516 5068 5518 5129
rect 5664 5069 5666 5129
rect 5662 5068 5668 5069
rect 3838 5064 3839 5068
rect 3843 5064 3844 5068
rect 3838 5063 3844 5064
rect 3978 5067 3984 5068
rect 3978 5063 3979 5067
rect 3983 5063 3984 5067
rect 1934 5059 1940 5060
rect 1975 5062 1979 5063
rect 946 5058 952 5059
rect 1975 5057 1979 5058
rect 1995 5062 1999 5063
rect 1995 5057 1999 5058
rect 2131 5062 2135 5063
rect 2131 5057 2135 5058
rect 2267 5062 2271 5063
rect 2267 5057 2271 5058
rect 2403 5062 2407 5063
rect 2403 5057 2407 5058
rect 2539 5062 2543 5063
rect 2539 5057 2543 5058
rect 2675 5062 2679 5063
rect 2675 5057 2679 5058
rect 2811 5062 2815 5063
rect 2811 5057 2815 5058
rect 2947 5062 2951 5063
rect 2947 5057 2951 5058
rect 3083 5062 3087 5063
rect 3083 5057 3087 5058
rect 3107 5062 3111 5063
rect 3107 5057 3111 5058
rect 3219 5062 3223 5063
rect 3219 5057 3223 5058
rect 3243 5062 3247 5063
rect 3243 5057 3247 5058
rect 3363 5062 3367 5063
rect 3363 5057 3367 5058
rect 3379 5062 3383 5063
rect 3379 5057 3383 5058
rect 3515 5062 3519 5063
rect 3515 5057 3519 5058
rect 3651 5062 3655 5063
rect 3651 5057 3655 5058
rect 3799 5062 3803 5063
rect 3978 5062 3984 5063
rect 4274 5067 4280 5068
rect 4274 5063 4275 5067
rect 4279 5063 4280 5067
rect 4274 5062 4280 5063
rect 4578 5067 4584 5068
rect 4578 5063 4579 5067
rect 4583 5063 4584 5067
rect 4578 5062 4584 5063
rect 4882 5067 4888 5068
rect 4882 5063 4883 5067
rect 4887 5063 4888 5067
rect 4882 5062 4888 5063
rect 5194 5067 5200 5068
rect 5194 5063 5195 5067
rect 5199 5063 5200 5067
rect 5194 5062 5200 5063
rect 5514 5067 5520 5068
rect 5514 5063 5515 5067
rect 5519 5063 5520 5067
rect 5662 5064 5663 5068
rect 5667 5064 5668 5068
rect 5662 5063 5668 5064
rect 5514 5062 5520 5063
rect 3799 5057 3803 5058
rect 294 5048 300 5049
rect 110 5047 116 5048
rect 110 5043 111 5047
rect 115 5043 116 5047
rect 294 5044 295 5048
rect 299 5044 300 5048
rect 294 5043 300 5044
rect 430 5048 436 5049
rect 430 5044 431 5048
rect 435 5044 436 5048
rect 430 5043 436 5044
rect 566 5048 572 5049
rect 566 5044 567 5048
rect 571 5044 572 5048
rect 566 5043 572 5044
rect 702 5048 708 5049
rect 702 5044 703 5048
rect 707 5044 708 5048
rect 702 5043 708 5044
rect 838 5048 844 5049
rect 838 5044 839 5048
rect 843 5044 844 5048
rect 838 5043 844 5044
rect 974 5048 980 5049
rect 974 5044 975 5048
rect 979 5044 980 5048
rect 974 5043 980 5044
rect 1934 5047 1940 5048
rect 1934 5043 1935 5047
rect 1939 5043 1940 5047
rect 110 5042 116 5043
rect 112 5007 114 5042
rect 296 5007 298 5043
rect 432 5007 434 5043
rect 568 5007 570 5043
rect 704 5007 706 5043
rect 840 5007 842 5043
rect 976 5007 978 5043
rect 1934 5042 1940 5043
rect 1936 5007 1938 5042
rect 111 5006 115 5007
rect 111 5001 115 5002
rect 159 5006 163 5007
rect 159 5001 163 5002
rect 295 5006 299 5007
rect 295 5001 299 5002
rect 431 5006 435 5007
rect 431 5001 435 5002
rect 567 5006 571 5007
rect 567 5001 571 5002
rect 703 5006 707 5007
rect 703 5001 707 5002
rect 839 5006 843 5007
rect 839 5001 843 5002
rect 975 5006 979 5007
rect 975 5001 979 5002
rect 1935 5006 1939 5007
rect 1935 5001 1939 5002
rect 112 4978 114 5001
rect 110 4977 116 4978
rect 160 4977 162 5001
rect 296 4977 298 5001
rect 432 4977 434 5001
rect 568 4977 570 5001
rect 704 4977 706 5001
rect 1936 4978 1938 5001
rect 1976 4997 1978 5057
rect 1974 4996 1980 4997
rect 3108 4996 3110 5057
rect 3244 4996 3246 5057
rect 3380 4996 3382 5057
rect 3516 4996 3518 5057
rect 3652 4996 3654 5057
rect 3800 4997 3802 5057
rect 4006 5052 4012 5053
rect 3838 5051 3844 5052
rect 3838 5047 3839 5051
rect 3843 5047 3844 5051
rect 4006 5048 4007 5052
rect 4011 5048 4012 5052
rect 4006 5047 4012 5048
rect 4302 5052 4308 5053
rect 4302 5048 4303 5052
rect 4307 5048 4308 5052
rect 4302 5047 4308 5048
rect 4606 5052 4612 5053
rect 4606 5048 4607 5052
rect 4611 5048 4612 5052
rect 4606 5047 4612 5048
rect 4910 5052 4916 5053
rect 4910 5048 4911 5052
rect 4915 5048 4916 5052
rect 4910 5047 4916 5048
rect 5222 5052 5228 5053
rect 5222 5048 5223 5052
rect 5227 5048 5228 5052
rect 5222 5047 5228 5048
rect 5542 5052 5548 5053
rect 5542 5048 5543 5052
rect 5547 5048 5548 5052
rect 5542 5047 5548 5048
rect 5662 5051 5668 5052
rect 5662 5047 5663 5051
rect 5667 5047 5668 5051
rect 3838 5046 3844 5047
rect 3840 5007 3842 5046
rect 4008 5007 4010 5047
rect 4304 5007 4306 5047
rect 4608 5007 4610 5047
rect 4912 5007 4914 5047
rect 5224 5007 5226 5047
rect 5544 5007 5546 5047
rect 5662 5046 5668 5047
rect 5664 5007 5666 5046
rect 3839 5006 3843 5007
rect 3839 5001 3843 5002
rect 4007 5006 4011 5007
rect 4007 5001 4011 5002
rect 4303 5006 4307 5007
rect 4303 5001 4307 5002
rect 4607 5006 4611 5007
rect 4607 5001 4611 5002
rect 4863 5006 4867 5007
rect 4863 5001 4867 5002
rect 4911 5006 4915 5007
rect 4911 5001 4915 5002
rect 4999 5006 5003 5007
rect 4999 5001 5003 5002
rect 5135 5006 5139 5007
rect 5135 5001 5139 5002
rect 5223 5006 5227 5007
rect 5223 5001 5227 5002
rect 5271 5006 5275 5007
rect 5271 5001 5275 5002
rect 5407 5006 5411 5007
rect 5407 5001 5411 5002
rect 5543 5006 5547 5007
rect 5543 5001 5547 5002
rect 5663 5006 5667 5007
rect 5663 5001 5667 5002
rect 3798 4996 3804 4997
rect 1974 4992 1975 4996
rect 1979 4992 1980 4996
rect 1974 4991 1980 4992
rect 3106 4995 3112 4996
rect 3106 4991 3107 4995
rect 3111 4991 3112 4995
rect 3106 4990 3112 4991
rect 3242 4995 3248 4996
rect 3242 4991 3243 4995
rect 3247 4991 3248 4995
rect 3242 4990 3248 4991
rect 3378 4995 3384 4996
rect 3378 4991 3379 4995
rect 3383 4991 3384 4995
rect 3378 4990 3384 4991
rect 3514 4995 3520 4996
rect 3514 4991 3515 4995
rect 3519 4991 3520 4995
rect 3514 4990 3520 4991
rect 3650 4995 3656 4996
rect 3650 4991 3651 4995
rect 3655 4991 3656 4995
rect 3798 4992 3799 4996
rect 3803 4992 3804 4996
rect 3798 4991 3804 4992
rect 3650 4990 3656 4991
rect 3134 4980 3140 4981
rect 1974 4979 1980 4980
rect 1934 4977 1940 4978
rect 110 4973 111 4977
rect 115 4973 116 4977
rect 110 4972 116 4973
rect 158 4976 164 4977
rect 158 4972 159 4976
rect 163 4972 164 4976
rect 158 4971 164 4972
rect 294 4976 300 4977
rect 294 4972 295 4976
rect 299 4972 300 4976
rect 294 4971 300 4972
rect 430 4976 436 4977
rect 430 4972 431 4976
rect 435 4972 436 4976
rect 430 4971 436 4972
rect 566 4976 572 4977
rect 566 4972 567 4976
rect 571 4972 572 4976
rect 566 4971 572 4972
rect 702 4976 708 4977
rect 702 4972 703 4976
rect 707 4972 708 4976
rect 1934 4973 1935 4977
rect 1939 4973 1940 4977
rect 1974 4975 1975 4979
rect 1979 4975 1980 4979
rect 3134 4976 3135 4980
rect 3139 4976 3140 4980
rect 3134 4975 3140 4976
rect 3270 4980 3276 4981
rect 3270 4976 3271 4980
rect 3275 4976 3276 4980
rect 3270 4975 3276 4976
rect 3406 4980 3412 4981
rect 3406 4976 3407 4980
rect 3411 4976 3412 4980
rect 3406 4975 3412 4976
rect 3542 4980 3548 4981
rect 3542 4976 3543 4980
rect 3547 4976 3548 4980
rect 3542 4975 3548 4976
rect 3678 4980 3684 4981
rect 3678 4976 3679 4980
rect 3683 4976 3684 4980
rect 3678 4975 3684 4976
rect 3798 4979 3804 4980
rect 3798 4975 3799 4979
rect 3803 4975 3804 4979
rect 3840 4978 3842 5001
rect 1974 4974 1980 4975
rect 1934 4972 1940 4973
rect 702 4971 708 4972
rect 130 4961 136 4962
rect 110 4960 116 4961
rect 110 4956 111 4960
rect 115 4956 116 4960
rect 130 4957 131 4961
rect 135 4957 136 4961
rect 130 4956 136 4957
rect 266 4961 272 4962
rect 266 4957 267 4961
rect 271 4957 272 4961
rect 266 4956 272 4957
rect 402 4961 408 4962
rect 402 4957 403 4961
rect 407 4957 408 4961
rect 402 4956 408 4957
rect 538 4961 544 4962
rect 538 4957 539 4961
rect 543 4957 544 4961
rect 538 4956 544 4957
rect 674 4961 680 4962
rect 674 4957 675 4961
rect 679 4957 680 4961
rect 674 4956 680 4957
rect 1934 4960 1940 4961
rect 1934 4956 1935 4960
rect 1939 4956 1940 4960
rect 110 4955 116 4956
rect 112 4887 114 4955
rect 132 4887 134 4956
rect 268 4887 270 4956
rect 404 4887 406 4956
rect 540 4887 542 4956
rect 676 4887 678 4956
rect 1934 4955 1940 4956
rect 1936 4887 1938 4955
rect 1976 4943 1978 4974
rect 3136 4943 3138 4975
rect 3272 4943 3274 4975
rect 3408 4943 3410 4975
rect 3544 4943 3546 4975
rect 3680 4943 3682 4975
rect 3798 4974 3804 4975
rect 3838 4977 3844 4978
rect 4864 4977 4866 5001
rect 5000 4977 5002 5001
rect 5136 4977 5138 5001
rect 5272 4977 5274 5001
rect 5408 4977 5410 5001
rect 5544 4977 5546 5001
rect 5664 4978 5666 5001
rect 5662 4977 5668 4978
rect 3800 4943 3802 4974
rect 3838 4973 3839 4977
rect 3843 4973 3844 4977
rect 3838 4972 3844 4973
rect 4862 4976 4868 4977
rect 4862 4972 4863 4976
rect 4867 4972 4868 4976
rect 4862 4971 4868 4972
rect 4998 4976 5004 4977
rect 4998 4972 4999 4976
rect 5003 4972 5004 4976
rect 4998 4971 5004 4972
rect 5134 4976 5140 4977
rect 5134 4972 5135 4976
rect 5139 4972 5140 4976
rect 5134 4971 5140 4972
rect 5270 4976 5276 4977
rect 5270 4972 5271 4976
rect 5275 4972 5276 4976
rect 5270 4971 5276 4972
rect 5406 4976 5412 4977
rect 5406 4972 5407 4976
rect 5411 4972 5412 4976
rect 5406 4971 5412 4972
rect 5542 4976 5548 4977
rect 5542 4972 5543 4976
rect 5547 4972 5548 4976
rect 5662 4973 5663 4977
rect 5667 4973 5668 4977
rect 5662 4972 5668 4973
rect 5542 4971 5548 4972
rect 4834 4961 4840 4962
rect 3838 4960 3844 4961
rect 3838 4956 3839 4960
rect 3843 4956 3844 4960
rect 4834 4957 4835 4961
rect 4839 4957 4840 4961
rect 4834 4956 4840 4957
rect 4970 4961 4976 4962
rect 4970 4957 4971 4961
rect 4975 4957 4976 4961
rect 4970 4956 4976 4957
rect 5106 4961 5112 4962
rect 5106 4957 5107 4961
rect 5111 4957 5112 4961
rect 5106 4956 5112 4957
rect 5242 4961 5248 4962
rect 5242 4957 5243 4961
rect 5247 4957 5248 4961
rect 5242 4956 5248 4957
rect 5378 4961 5384 4962
rect 5378 4957 5379 4961
rect 5383 4957 5384 4961
rect 5378 4956 5384 4957
rect 5514 4961 5520 4962
rect 5514 4957 5515 4961
rect 5519 4957 5520 4961
rect 5514 4956 5520 4957
rect 5662 4960 5668 4961
rect 5662 4956 5663 4960
rect 5667 4956 5668 4960
rect 3838 4955 3844 4956
rect 1975 4942 1979 4943
rect 1975 4937 1979 4938
rect 3135 4942 3139 4943
rect 3135 4937 3139 4938
rect 3271 4942 3275 4943
rect 3271 4937 3275 4938
rect 3407 4942 3411 4943
rect 3407 4937 3411 4938
rect 3543 4942 3547 4943
rect 3543 4937 3547 4938
rect 3679 4942 3683 4943
rect 3679 4937 3683 4938
rect 3799 4942 3803 4943
rect 3799 4937 3803 4938
rect 1976 4914 1978 4937
rect 1974 4913 1980 4914
rect 3136 4913 3138 4937
rect 3272 4913 3274 4937
rect 3408 4913 3410 4937
rect 3544 4913 3546 4937
rect 3680 4913 3682 4937
rect 3800 4914 3802 4937
rect 3798 4913 3804 4914
rect 1974 4909 1975 4913
rect 1979 4909 1980 4913
rect 1974 4908 1980 4909
rect 3134 4912 3140 4913
rect 3134 4908 3135 4912
rect 3139 4908 3140 4912
rect 3134 4907 3140 4908
rect 3270 4912 3276 4913
rect 3270 4908 3271 4912
rect 3275 4908 3276 4912
rect 3270 4907 3276 4908
rect 3406 4912 3412 4913
rect 3406 4908 3407 4912
rect 3411 4908 3412 4912
rect 3406 4907 3412 4908
rect 3542 4912 3548 4913
rect 3542 4908 3543 4912
rect 3547 4908 3548 4912
rect 3542 4907 3548 4908
rect 3678 4912 3684 4913
rect 3678 4908 3679 4912
rect 3683 4908 3684 4912
rect 3798 4909 3799 4913
rect 3803 4909 3804 4913
rect 3798 4908 3804 4909
rect 3678 4907 3684 4908
rect 3106 4897 3112 4898
rect 1974 4896 1980 4897
rect 1974 4892 1975 4896
rect 1979 4892 1980 4896
rect 3106 4893 3107 4897
rect 3111 4893 3112 4897
rect 3106 4892 3112 4893
rect 3242 4897 3248 4898
rect 3242 4893 3243 4897
rect 3247 4893 3248 4897
rect 3242 4892 3248 4893
rect 3378 4897 3384 4898
rect 3378 4893 3379 4897
rect 3383 4893 3384 4897
rect 3378 4892 3384 4893
rect 3514 4897 3520 4898
rect 3514 4893 3515 4897
rect 3519 4893 3520 4897
rect 3514 4892 3520 4893
rect 3650 4897 3656 4898
rect 3650 4893 3651 4897
rect 3655 4893 3656 4897
rect 3650 4892 3656 4893
rect 3798 4896 3804 4897
rect 3798 4892 3799 4896
rect 3803 4892 3804 4896
rect 1974 4891 1980 4892
rect 111 4886 115 4887
rect 111 4881 115 4882
rect 131 4886 135 4887
rect 131 4881 135 4882
rect 267 4886 271 4887
rect 267 4881 271 4882
rect 403 4886 407 4887
rect 403 4881 407 4882
rect 539 4886 543 4887
rect 539 4881 543 4882
rect 675 4886 679 4887
rect 675 4881 679 4882
rect 1935 4886 1939 4887
rect 1935 4881 1939 4882
rect 112 4821 114 4881
rect 110 4820 116 4821
rect 132 4820 134 4881
rect 268 4820 270 4881
rect 404 4820 406 4881
rect 540 4820 542 4881
rect 676 4820 678 4881
rect 1936 4821 1938 4881
rect 1934 4820 1940 4821
rect 110 4816 111 4820
rect 115 4816 116 4820
rect 110 4815 116 4816
rect 130 4819 136 4820
rect 130 4815 131 4819
rect 135 4815 136 4819
rect 130 4814 136 4815
rect 266 4819 272 4820
rect 266 4815 267 4819
rect 271 4815 272 4819
rect 266 4814 272 4815
rect 402 4819 408 4820
rect 402 4815 403 4819
rect 407 4815 408 4819
rect 402 4814 408 4815
rect 538 4819 544 4820
rect 538 4815 539 4819
rect 543 4815 544 4819
rect 538 4814 544 4815
rect 674 4819 680 4820
rect 674 4815 675 4819
rect 679 4815 680 4819
rect 1934 4816 1935 4820
rect 1939 4816 1940 4820
rect 1934 4815 1940 4816
rect 674 4814 680 4815
rect 158 4804 164 4805
rect 110 4803 116 4804
rect 110 4799 111 4803
rect 115 4799 116 4803
rect 158 4800 159 4804
rect 163 4800 164 4804
rect 158 4799 164 4800
rect 294 4804 300 4805
rect 294 4800 295 4804
rect 299 4800 300 4804
rect 294 4799 300 4800
rect 430 4804 436 4805
rect 430 4800 431 4804
rect 435 4800 436 4804
rect 430 4799 436 4800
rect 566 4804 572 4805
rect 566 4800 567 4804
rect 571 4800 572 4804
rect 566 4799 572 4800
rect 702 4804 708 4805
rect 702 4800 703 4804
rect 707 4800 708 4804
rect 702 4799 708 4800
rect 1934 4803 1940 4804
rect 1976 4803 1978 4891
rect 3108 4803 3110 4892
rect 3244 4803 3246 4892
rect 3380 4803 3382 4892
rect 3516 4803 3518 4892
rect 3652 4803 3654 4892
rect 3798 4891 3804 4892
rect 3800 4803 3802 4891
rect 3840 4883 3842 4955
rect 4836 4883 4838 4956
rect 4972 4883 4974 4956
rect 5108 4883 5110 4956
rect 5244 4883 5246 4956
rect 5380 4883 5382 4956
rect 5516 4883 5518 4956
rect 5662 4955 5668 4956
rect 5664 4883 5666 4955
rect 3839 4882 3843 4883
rect 3839 4877 3843 4878
rect 4483 4882 4487 4883
rect 4483 4877 4487 4878
rect 4675 4882 4679 4883
rect 4675 4877 4679 4878
rect 4835 4882 4839 4883
rect 4835 4877 4839 4878
rect 4875 4882 4879 4883
rect 4875 4877 4879 4878
rect 4971 4882 4975 4883
rect 4971 4877 4975 4878
rect 5091 4882 5095 4883
rect 5091 4877 5095 4878
rect 5107 4882 5111 4883
rect 5107 4877 5111 4878
rect 5243 4882 5247 4883
rect 5243 4877 5247 4878
rect 5315 4882 5319 4883
rect 5315 4877 5319 4878
rect 5379 4882 5383 4883
rect 5379 4877 5383 4878
rect 5515 4882 5519 4883
rect 5515 4877 5519 4878
rect 5663 4882 5667 4883
rect 5663 4877 5667 4878
rect 3840 4817 3842 4877
rect 3838 4816 3844 4817
rect 4484 4816 4486 4877
rect 4676 4816 4678 4877
rect 4876 4816 4878 4877
rect 5092 4816 5094 4877
rect 5316 4816 5318 4877
rect 5516 4816 5518 4877
rect 5664 4817 5666 4877
rect 5662 4816 5668 4817
rect 3838 4812 3839 4816
rect 3843 4812 3844 4816
rect 3838 4811 3844 4812
rect 4482 4815 4488 4816
rect 4482 4811 4483 4815
rect 4487 4811 4488 4815
rect 4482 4810 4488 4811
rect 4674 4815 4680 4816
rect 4674 4811 4675 4815
rect 4679 4811 4680 4815
rect 4674 4810 4680 4811
rect 4874 4815 4880 4816
rect 4874 4811 4875 4815
rect 4879 4811 4880 4815
rect 4874 4810 4880 4811
rect 5090 4815 5096 4816
rect 5090 4811 5091 4815
rect 5095 4811 5096 4815
rect 5090 4810 5096 4811
rect 5314 4815 5320 4816
rect 5314 4811 5315 4815
rect 5319 4811 5320 4815
rect 5314 4810 5320 4811
rect 5514 4815 5520 4816
rect 5514 4811 5515 4815
rect 5519 4811 5520 4815
rect 5662 4812 5663 4816
rect 5667 4812 5668 4816
rect 5662 4811 5668 4812
rect 5514 4810 5520 4811
rect 1934 4799 1935 4803
rect 1939 4799 1940 4803
rect 110 4798 116 4799
rect 112 4771 114 4798
rect 160 4771 162 4799
rect 296 4771 298 4799
rect 432 4771 434 4799
rect 568 4771 570 4799
rect 704 4771 706 4799
rect 1934 4798 1940 4799
rect 1975 4802 1979 4803
rect 1936 4771 1938 4798
rect 1975 4797 1979 4798
rect 3107 4802 3111 4803
rect 3107 4797 3111 4798
rect 3243 4802 3247 4803
rect 3243 4797 3247 4798
rect 3379 4802 3383 4803
rect 3379 4797 3383 4798
rect 3515 4802 3519 4803
rect 3515 4797 3519 4798
rect 3651 4802 3655 4803
rect 3651 4797 3655 4798
rect 3799 4802 3803 4803
rect 4510 4800 4516 4801
rect 3799 4797 3803 4798
rect 3838 4799 3844 4800
rect 111 4770 115 4771
rect 111 4765 115 4766
rect 159 4770 163 4771
rect 159 4765 163 4766
rect 295 4770 299 4771
rect 295 4765 299 4766
rect 431 4770 435 4771
rect 431 4765 435 4766
rect 567 4770 571 4771
rect 567 4765 571 4766
rect 703 4770 707 4771
rect 703 4765 707 4766
rect 1935 4770 1939 4771
rect 1935 4765 1939 4766
rect 112 4742 114 4765
rect 110 4741 116 4742
rect 160 4741 162 4765
rect 296 4741 298 4765
rect 432 4741 434 4765
rect 568 4741 570 4765
rect 704 4741 706 4765
rect 1936 4742 1938 4765
rect 1934 4741 1940 4742
rect 110 4737 111 4741
rect 115 4737 116 4741
rect 110 4736 116 4737
rect 158 4740 164 4741
rect 158 4736 159 4740
rect 163 4736 164 4740
rect 158 4735 164 4736
rect 294 4740 300 4741
rect 294 4736 295 4740
rect 299 4736 300 4740
rect 294 4735 300 4736
rect 430 4740 436 4741
rect 430 4736 431 4740
rect 435 4736 436 4740
rect 430 4735 436 4736
rect 566 4740 572 4741
rect 566 4736 567 4740
rect 571 4736 572 4740
rect 566 4735 572 4736
rect 702 4740 708 4741
rect 702 4736 703 4740
rect 707 4736 708 4740
rect 1934 4737 1935 4741
rect 1939 4737 1940 4741
rect 1976 4737 1978 4797
rect 1934 4736 1940 4737
rect 1974 4736 1980 4737
rect 3108 4736 3110 4797
rect 3244 4736 3246 4797
rect 3380 4736 3382 4797
rect 3516 4736 3518 4797
rect 3652 4736 3654 4797
rect 3800 4737 3802 4797
rect 3838 4795 3839 4799
rect 3843 4795 3844 4799
rect 4510 4796 4511 4800
rect 4515 4796 4516 4800
rect 4510 4795 4516 4796
rect 4702 4800 4708 4801
rect 4702 4796 4703 4800
rect 4707 4796 4708 4800
rect 4702 4795 4708 4796
rect 4902 4800 4908 4801
rect 4902 4796 4903 4800
rect 4907 4796 4908 4800
rect 4902 4795 4908 4796
rect 5118 4800 5124 4801
rect 5118 4796 5119 4800
rect 5123 4796 5124 4800
rect 5118 4795 5124 4796
rect 5342 4800 5348 4801
rect 5342 4796 5343 4800
rect 5347 4796 5348 4800
rect 5342 4795 5348 4796
rect 5542 4800 5548 4801
rect 5542 4796 5543 4800
rect 5547 4796 5548 4800
rect 5542 4795 5548 4796
rect 5662 4799 5668 4800
rect 5662 4795 5663 4799
rect 5667 4795 5668 4799
rect 3838 4794 3844 4795
rect 3840 4751 3842 4794
rect 4512 4751 4514 4795
rect 4704 4751 4706 4795
rect 4904 4751 4906 4795
rect 5120 4751 5122 4795
rect 5344 4751 5346 4795
rect 5544 4751 5546 4795
rect 5662 4794 5668 4795
rect 5664 4751 5666 4794
rect 3839 4750 3843 4751
rect 3839 4745 3843 4746
rect 4119 4750 4123 4751
rect 4119 4745 4123 4746
rect 4375 4750 4379 4751
rect 4375 4745 4379 4746
rect 4511 4750 4515 4751
rect 4511 4745 4515 4746
rect 4647 4750 4651 4751
rect 4647 4745 4651 4746
rect 4703 4750 4707 4751
rect 4703 4745 4707 4746
rect 4903 4750 4907 4751
rect 4903 4745 4907 4746
rect 4943 4750 4947 4751
rect 4943 4745 4947 4746
rect 5119 4750 5123 4751
rect 5119 4745 5123 4746
rect 5255 4750 5259 4751
rect 5255 4745 5259 4746
rect 5343 4750 5347 4751
rect 5343 4745 5347 4746
rect 5543 4750 5547 4751
rect 5543 4745 5547 4746
rect 5663 4750 5667 4751
rect 5663 4745 5667 4746
rect 3798 4736 3804 4737
rect 702 4735 708 4736
rect 1974 4732 1975 4736
rect 1979 4732 1980 4736
rect 1974 4731 1980 4732
rect 3106 4735 3112 4736
rect 3106 4731 3107 4735
rect 3111 4731 3112 4735
rect 3106 4730 3112 4731
rect 3242 4735 3248 4736
rect 3242 4731 3243 4735
rect 3247 4731 3248 4735
rect 3242 4730 3248 4731
rect 3378 4735 3384 4736
rect 3378 4731 3379 4735
rect 3383 4731 3384 4735
rect 3378 4730 3384 4731
rect 3514 4735 3520 4736
rect 3514 4731 3515 4735
rect 3519 4731 3520 4735
rect 3514 4730 3520 4731
rect 3650 4735 3656 4736
rect 3650 4731 3651 4735
rect 3655 4731 3656 4735
rect 3798 4732 3799 4736
rect 3803 4732 3804 4736
rect 3798 4731 3804 4732
rect 3650 4730 3656 4731
rect 130 4725 136 4726
rect 110 4724 116 4725
rect 110 4720 111 4724
rect 115 4720 116 4724
rect 130 4721 131 4725
rect 135 4721 136 4725
rect 130 4720 136 4721
rect 266 4725 272 4726
rect 266 4721 267 4725
rect 271 4721 272 4725
rect 266 4720 272 4721
rect 402 4725 408 4726
rect 402 4721 403 4725
rect 407 4721 408 4725
rect 402 4720 408 4721
rect 538 4725 544 4726
rect 538 4721 539 4725
rect 543 4721 544 4725
rect 538 4720 544 4721
rect 674 4725 680 4726
rect 674 4721 675 4725
rect 679 4721 680 4725
rect 674 4720 680 4721
rect 1934 4724 1940 4725
rect 1934 4720 1935 4724
rect 1939 4720 1940 4724
rect 3840 4722 3842 4745
rect 3838 4721 3844 4722
rect 4120 4721 4122 4745
rect 4376 4721 4378 4745
rect 4648 4721 4650 4745
rect 4944 4721 4946 4745
rect 5256 4721 5258 4745
rect 5544 4721 5546 4745
rect 5664 4722 5666 4745
rect 5662 4721 5668 4722
rect 3134 4720 3140 4721
rect 110 4719 116 4720
rect 112 4651 114 4719
rect 132 4651 134 4720
rect 268 4651 270 4720
rect 404 4651 406 4720
rect 540 4651 542 4720
rect 676 4651 678 4720
rect 1934 4719 1940 4720
rect 1974 4719 1980 4720
rect 1936 4651 1938 4719
rect 1974 4715 1975 4719
rect 1979 4715 1980 4719
rect 3134 4716 3135 4720
rect 3139 4716 3140 4720
rect 3134 4715 3140 4716
rect 3270 4720 3276 4721
rect 3270 4716 3271 4720
rect 3275 4716 3276 4720
rect 3270 4715 3276 4716
rect 3406 4720 3412 4721
rect 3406 4716 3407 4720
rect 3411 4716 3412 4720
rect 3406 4715 3412 4716
rect 3542 4720 3548 4721
rect 3542 4716 3543 4720
rect 3547 4716 3548 4720
rect 3542 4715 3548 4716
rect 3678 4720 3684 4721
rect 3678 4716 3679 4720
rect 3683 4716 3684 4720
rect 3678 4715 3684 4716
rect 3798 4719 3804 4720
rect 3798 4715 3799 4719
rect 3803 4715 3804 4719
rect 3838 4717 3839 4721
rect 3843 4717 3844 4721
rect 3838 4716 3844 4717
rect 4118 4720 4124 4721
rect 4118 4716 4119 4720
rect 4123 4716 4124 4720
rect 4118 4715 4124 4716
rect 4374 4720 4380 4721
rect 4374 4716 4375 4720
rect 4379 4716 4380 4720
rect 4374 4715 4380 4716
rect 4646 4720 4652 4721
rect 4646 4716 4647 4720
rect 4651 4716 4652 4720
rect 4646 4715 4652 4716
rect 4942 4720 4948 4721
rect 4942 4716 4943 4720
rect 4947 4716 4948 4720
rect 4942 4715 4948 4716
rect 5254 4720 5260 4721
rect 5254 4716 5255 4720
rect 5259 4716 5260 4720
rect 5254 4715 5260 4716
rect 5542 4720 5548 4721
rect 5542 4716 5543 4720
rect 5547 4716 5548 4720
rect 5662 4717 5663 4721
rect 5667 4717 5668 4721
rect 5662 4716 5668 4717
rect 5542 4715 5548 4716
rect 1974 4714 1980 4715
rect 1976 4651 1978 4714
rect 3136 4651 3138 4715
rect 3272 4651 3274 4715
rect 3408 4651 3410 4715
rect 3544 4651 3546 4715
rect 3680 4651 3682 4715
rect 3798 4714 3804 4715
rect 3800 4651 3802 4714
rect 4090 4705 4096 4706
rect 3838 4704 3844 4705
rect 3838 4700 3839 4704
rect 3843 4700 3844 4704
rect 4090 4701 4091 4705
rect 4095 4701 4096 4705
rect 4090 4700 4096 4701
rect 4346 4705 4352 4706
rect 4346 4701 4347 4705
rect 4351 4701 4352 4705
rect 4346 4700 4352 4701
rect 4618 4705 4624 4706
rect 4618 4701 4619 4705
rect 4623 4701 4624 4705
rect 4618 4700 4624 4701
rect 4914 4705 4920 4706
rect 4914 4701 4915 4705
rect 4919 4701 4920 4705
rect 4914 4700 4920 4701
rect 5226 4705 5232 4706
rect 5226 4701 5227 4705
rect 5231 4701 5232 4705
rect 5226 4700 5232 4701
rect 5514 4705 5520 4706
rect 5514 4701 5515 4705
rect 5519 4701 5520 4705
rect 5514 4700 5520 4701
rect 5662 4704 5668 4705
rect 5662 4700 5663 4704
rect 5667 4700 5668 4704
rect 3838 4699 3844 4700
rect 111 4650 115 4651
rect 111 4645 115 4646
rect 131 4650 135 4651
rect 131 4645 135 4646
rect 211 4650 215 4651
rect 211 4645 215 4646
rect 267 4650 271 4651
rect 267 4645 271 4646
rect 403 4650 407 4651
rect 403 4645 407 4646
rect 427 4650 431 4651
rect 427 4645 431 4646
rect 539 4650 543 4651
rect 539 4645 543 4646
rect 667 4650 671 4651
rect 667 4645 671 4646
rect 675 4650 679 4651
rect 675 4645 679 4646
rect 931 4650 935 4651
rect 931 4645 935 4646
rect 1219 4650 1223 4651
rect 1219 4645 1223 4646
rect 1515 4650 1519 4651
rect 1515 4645 1519 4646
rect 1787 4650 1791 4651
rect 1787 4645 1791 4646
rect 1935 4650 1939 4651
rect 1935 4645 1939 4646
rect 1975 4650 1979 4651
rect 1975 4645 1979 4646
rect 2023 4650 2027 4651
rect 2023 4645 2027 4646
rect 2159 4650 2163 4651
rect 2159 4645 2163 4646
rect 2311 4650 2315 4651
rect 2311 4645 2315 4646
rect 2479 4650 2483 4651
rect 2479 4645 2483 4646
rect 2655 4650 2659 4651
rect 2655 4645 2659 4646
rect 2831 4650 2835 4651
rect 2831 4645 2835 4646
rect 3007 4650 3011 4651
rect 3007 4645 3011 4646
rect 3135 4650 3139 4651
rect 3135 4645 3139 4646
rect 3183 4650 3187 4651
rect 3183 4645 3187 4646
rect 3271 4650 3275 4651
rect 3271 4645 3275 4646
rect 3351 4650 3355 4651
rect 3351 4645 3355 4646
rect 3407 4650 3411 4651
rect 3407 4645 3411 4646
rect 3527 4650 3531 4651
rect 3527 4645 3531 4646
rect 3543 4650 3547 4651
rect 3543 4645 3547 4646
rect 3679 4650 3683 4651
rect 3679 4645 3683 4646
rect 3799 4650 3803 4651
rect 3799 4645 3803 4646
rect 112 4585 114 4645
rect 110 4584 116 4585
rect 212 4584 214 4645
rect 428 4584 430 4645
rect 668 4584 670 4645
rect 932 4584 934 4645
rect 1220 4584 1222 4645
rect 1516 4584 1518 4645
rect 1788 4584 1790 4645
rect 1936 4585 1938 4645
rect 1976 4622 1978 4645
rect 1974 4621 1980 4622
rect 2024 4621 2026 4645
rect 2160 4621 2162 4645
rect 2312 4621 2314 4645
rect 2480 4621 2482 4645
rect 2656 4621 2658 4645
rect 2832 4621 2834 4645
rect 3008 4621 3010 4645
rect 3184 4621 3186 4645
rect 3352 4621 3354 4645
rect 3528 4621 3530 4645
rect 3680 4621 3682 4645
rect 3800 4622 3802 4645
rect 3798 4621 3804 4622
rect 1974 4617 1975 4621
rect 1979 4617 1980 4621
rect 1974 4616 1980 4617
rect 2022 4620 2028 4621
rect 2022 4616 2023 4620
rect 2027 4616 2028 4620
rect 2022 4615 2028 4616
rect 2158 4620 2164 4621
rect 2158 4616 2159 4620
rect 2163 4616 2164 4620
rect 2158 4615 2164 4616
rect 2310 4620 2316 4621
rect 2310 4616 2311 4620
rect 2315 4616 2316 4620
rect 2310 4615 2316 4616
rect 2478 4620 2484 4621
rect 2478 4616 2479 4620
rect 2483 4616 2484 4620
rect 2478 4615 2484 4616
rect 2654 4620 2660 4621
rect 2654 4616 2655 4620
rect 2659 4616 2660 4620
rect 2654 4615 2660 4616
rect 2830 4620 2836 4621
rect 2830 4616 2831 4620
rect 2835 4616 2836 4620
rect 2830 4615 2836 4616
rect 3006 4620 3012 4621
rect 3006 4616 3007 4620
rect 3011 4616 3012 4620
rect 3006 4615 3012 4616
rect 3182 4620 3188 4621
rect 3182 4616 3183 4620
rect 3187 4616 3188 4620
rect 3182 4615 3188 4616
rect 3350 4620 3356 4621
rect 3350 4616 3351 4620
rect 3355 4616 3356 4620
rect 3350 4615 3356 4616
rect 3526 4620 3532 4621
rect 3526 4616 3527 4620
rect 3531 4616 3532 4620
rect 3526 4615 3532 4616
rect 3678 4620 3684 4621
rect 3678 4616 3679 4620
rect 3683 4616 3684 4620
rect 3798 4617 3799 4621
rect 3803 4617 3804 4621
rect 3840 4619 3842 4699
rect 4092 4619 4094 4700
rect 4348 4619 4350 4700
rect 4620 4619 4622 4700
rect 4916 4619 4918 4700
rect 5228 4619 5230 4700
rect 5516 4619 5518 4700
rect 5662 4699 5668 4700
rect 5664 4619 5666 4699
rect 3798 4616 3804 4617
rect 3839 4618 3843 4619
rect 3678 4615 3684 4616
rect 3839 4613 3843 4614
rect 4035 4618 4039 4619
rect 4035 4613 4039 4614
rect 4091 4618 4095 4619
rect 4091 4613 4095 4614
rect 4331 4618 4335 4619
rect 4331 4613 4335 4614
rect 4347 4618 4351 4619
rect 4347 4613 4351 4614
rect 4619 4618 4623 4619
rect 4619 4613 4623 4614
rect 4627 4618 4631 4619
rect 4627 4613 4631 4614
rect 4915 4618 4919 4619
rect 4915 4613 4919 4614
rect 4931 4618 4935 4619
rect 4931 4613 4935 4614
rect 5227 4618 5231 4619
rect 5227 4613 5231 4614
rect 5235 4618 5239 4619
rect 5235 4613 5239 4614
rect 5515 4618 5519 4619
rect 5515 4613 5519 4614
rect 5663 4618 5667 4619
rect 5663 4613 5667 4614
rect 1994 4605 2000 4606
rect 1974 4604 1980 4605
rect 1974 4600 1975 4604
rect 1979 4600 1980 4604
rect 1994 4601 1995 4605
rect 1999 4601 2000 4605
rect 1994 4600 2000 4601
rect 2130 4605 2136 4606
rect 2130 4601 2131 4605
rect 2135 4601 2136 4605
rect 2130 4600 2136 4601
rect 2282 4605 2288 4606
rect 2282 4601 2283 4605
rect 2287 4601 2288 4605
rect 2282 4600 2288 4601
rect 2450 4605 2456 4606
rect 2450 4601 2451 4605
rect 2455 4601 2456 4605
rect 2450 4600 2456 4601
rect 2626 4605 2632 4606
rect 2626 4601 2627 4605
rect 2631 4601 2632 4605
rect 2626 4600 2632 4601
rect 2802 4605 2808 4606
rect 2802 4601 2803 4605
rect 2807 4601 2808 4605
rect 2802 4600 2808 4601
rect 2978 4605 2984 4606
rect 2978 4601 2979 4605
rect 2983 4601 2984 4605
rect 2978 4600 2984 4601
rect 3154 4605 3160 4606
rect 3154 4601 3155 4605
rect 3159 4601 3160 4605
rect 3154 4600 3160 4601
rect 3322 4605 3328 4606
rect 3322 4601 3323 4605
rect 3327 4601 3328 4605
rect 3322 4600 3328 4601
rect 3498 4605 3504 4606
rect 3498 4601 3499 4605
rect 3503 4601 3504 4605
rect 3498 4600 3504 4601
rect 3650 4605 3656 4606
rect 3650 4601 3651 4605
rect 3655 4601 3656 4605
rect 3650 4600 3656 4601
rect 3798 4604 3804 4605
rect 3798 4600 3799 4604
rect 3803 4600 3804 4604
rect 1974 4599 1980 4600
rect 1934 4584 1940 4585
rect 110 4580 111 4584
rect 115 4580 116 4584
rect 110 4579 116 4580
rect 210 4583 216 4584
rect 210 4579 211 4583
rect 215 4579 216 4583
rect 210 4578 216 4579
rect 426 4583 432 4584
rect 426 4579 427 4583
rect 431 4579 432 4583
rect 426 4578 432 4579
rect 666 4583 672 4584
rect 666 4579 667 4583
rect 671 4579 672 4583
rect 666 4578 672 4579
rect 930 4583 936 4584
rect 930 4579 931 4583
rect 935 4579 936 4583
rect 930 4578 936 4579
rect 1218 4583 1224 4584
rect 1218 4579 1219 4583
rect 1223 4579 1224 4583
rect 1218 4578 1224 4579
rect 1514 4583 1520 4584
rect 1514 4579 1515 4583
rect 1519 4579 1520 4583
rect 1514 4578 1520 4579
rect 1786 4583 1792 4584
rect 1786 4579 1787 4583
rect 1791 4579 1792 4583
rect 1934 4580 1935 4584
rect 1939 4580 1940 4584
rect 1934 4579 1940 4580
rect 1786 4578 1792 4579
rect 238 4568 244 4569
rect 110 4567 116 4568
rect 110 4563 111 4567
rect 115 4563 116 4567
rect 238 4564 239 4568
rect 243 4564 244 4568
rect 238 4563 244 4564
rect 454 4568 460 4569
rect 454 4564 455 4568
rect 459 4564 460 4568
rect 454 4563 460 4564
rect 694 4568 700 4569
rect 694 4564 695 4568
rect 699 4564 700 4568
rect 694 4563 700 4564
rect 958 4568 964 4569
rect 958 4564 959 4568
rect 963 4564 964 4568
rect 958 4563 964 4564
rect 1246 4568 1252 4569
rect 1246 4564 1247 4568
rect 1251 4564 1252 4568
rect 1246 4563 1252 4564
rect 1542 4568 1548 4569
rect 1542 4564 1543 4568
rect 1547 4564 1548 4568
rect 1542 4563 1548 4564
rect 1814 4568 1820 4569
rect 1814 4564 1815 4568
rect 1819 4564 1820 4568
rect 1814 4563 1820 4564
rect 1934 4567 1940 4568
rect 1934 4563 1935 4567
rect 1939 4563 1940 4567
rect 110 4562 116 4563
rect 112 4539 114 4562
rect 240 4539 242 4563
rect 456 4539 458 4563
rect 696 4539 698 4563
rect 960 4539 962 4563
rect 1248 4539 1250 4563
rect 1544 4539 1546 4563
rect 1816 4539 1818 4563
rect 1934 4562 1940 4563
rect 1936 4539 1938 4562
rect 1976 4539 1978 4599
rect 1996 4539 1998 4600
rect 2132 4539 2134 4600
rect 2284 4539 2286 4600
rect 2452 4539 2454 4600
rect 2628 4539 2630 4600
rect 2804 4539 2806 4600
rect 2980 4539 2982 4600
rect 3156 4539 3158 4600
rect 3324 4539 3326 4600
rect 3500 4539 3502 4600
rect 3652 4539 3654 4600
rect 3798 4599 3804 4600
rect 3800 4539 3802 4599
rect 3840 4553 3842 4613
rect 3838 4552 3844 4553
rect 4036 4552 4038 4613
rect 4332 4552 4334 4613
rect 4628 4552 4630 4613
rect 4932 4552 4934 4613
rect 5236 4552 5238 4613
rect 5516 4552 5518 4613
rect 5664 4553 5666 4613
rect 5662 4552 5668 4553
rect 3838 4548 3839 4552
rect 3843 4548 3844 4552
rect 3838 4547 3844 4548
rect 4034 4551 4040 4552
rect 4034 4547 4035 4551
rect 4039 4547 4040 4551
rect 4034 4546 4040 4547
rect 4330 4551 4336 4552
rect 4330 4547 4331 4551
rect 4335 4547 4336 4551
rect 4330 4546 4336 4547
rect 4626 4551 4632 4552
rect 4626 4547 4627 4551
rect 4631 4547 4632 4551
rect 4626 4546 4632 4547
rect 4930 4551 4936 4552
rect 4930 4547 4931 4551
rect 4935 4547 4936 4551
rect 4930 4546 4936 4547
rect 5234 4551 5240 4552
rect 5234 4547 5235 4551
rect 5239 4547 5240 4551
rect 5234 4546 5240 4547
rect 5514 4551 5520 4552
rect 5514 4547 5515 4551
rect 5519 4547 5520 4551
rect 5662 4548 5663 4552
rect 5667 4548 5668 4552
rect 5662 4547 5668 4548
rect 5514 4546 5520 4547
rect 111 4538 115 4539
rect 111 4533 115 4534
rect 239 4538 243 4539
rect 239 4533 243 4534
rect 447 4538 451 4539
rect 447 4533 451 4534
rect 455 4538 459 4539
rect 455 4533 459 4534
rect 623 4538 627 4539
rect 623 4533 627 4534
rect 695 4538 699 4539
rect 695 4533 699 4534
rect 807 4538 811 4539
rect 807 4533 811 4534
rect 959 4538 963 4539
rect 959 4533 963 4534
rect 999 4538 1003 4539
rect 999 4533 1003 4534
rect 1199 4538 1203 4539
rect 1199 4533 1203 4534
rect 1247 4538 1251 4539
rect 1247 4533 1251 4534
rect 1407 4538 1411 4539
rect 1407 4533 1411 4534
rect 1543 4538 1547 4539
rect 1543 4533 1547 4534
rect 1623 4538 1627 4539
rect 1623 4533 1627 4534
rect 1815 4538 1819 4539
rect 1815 4533 1819 4534
rect 1935 4538 1939 4539
rect 1935 4533 1939 4534
rect 1975 4538 1979 4539
rect 1975 4533 1979 4534
rect 1995 4538 1999 4539
rect 1995 4533 1999 4534
rect 2131 4538 2135 4539
rect 2131 4533 2135 4534
rect 2227 4538 2231 4539
rect 2227 4533 2231 4534
rect 2283 4538 2287 4539
rect 2283 4533 2287 4534
rect 2451 4538 2455 4539
rect 2451 4533 2455 4534
rect 2459 4538 2463 4539
rect 2459 4533 2463 4534
rect 2627 4538 2631 4539
rect 2627 4533 2631 4534
rect 2691 4538 2695 4539
rect 2691 4533 2695 4534
rect 2803 4538 2807 4539
rect 2803 4533 2807 4534
rect 2915 4538 2919 4539
rect 2915 4533 2919 4534
rect 2979 4538 2983 4539
rect 2979 4533 2983 4534
rect 3131 4538 3135 4539
rect 3131 4533 3135 4534
rect 3155 4538 3159 4539
rect 3155 4533 3159 4534
rect 3323 4538 3327 4539
rect 3323 4533 3327 4534
rect 3355 4538 3359 4539
rect 3355 4533 3359 4534
rect 3499 4538 3503 4539
rect 3499 4533 3503 4534
rect 3579 4538 3583 4539
rect 3579 4533 3583 4534
rect 3651 4538 3655 4539
rect 3651 4533 3655 4534
rect 3799 4538 3803 4539
rect 4062 4536 4068 4537
rect 3799 4533 3803 4534
rect 3838 4535 3844 4536
rect 112 4510 114 4533
rect 110 4509 116 4510
rect 448 4509 450 4533
rect 624 4509 626 4533
rect 808 4509 810 4533
rect 1000 4509 1002 4533
rect 1200 4509 1202 4533
rect 1408 4509 1410 4533
rect 1624 4509 1626 4533
rect 1816 4509 1818 4533
rect 1936 4510 1938 4533
rect 1934 4509 1940 4510
rect 110 4505 111 4509
rect 115 4505 116 4509
rect 110 4504 116 4505
rect 446 4508 452 4509
rect 446 4504 447 4508
rect 451 4504 452 4508
rect 446 4503 452 4504
rect 622 4508 628 4509
rect 622 4504 623 4508
rect 627 4504 628 4508
rect 622 4503 628 4504
rect 806 4508 812 4509
rect 806 4504 807 4508
rect 811 4504 812 4508
rect 806 4503 812 4504
rect 998 4508 1004 4509
rect 998 4504 999 4508
rect 1003 4504 1004 4508
rect 998 4503 1004 4504
rect 1198 4508 1204 4509
rect 1198 4504 1199 4508
rect 1203 4504 1204 4508
rect 1198 4503 1204 4504
rect 1406 4508 1412 4509
rect 1406 4504 1407 4508
rect 1411 4504 1412 4508
rect 1406 4503 1412 4504
rect 1622 4508 1628 4509
rect 1622 4504 1623 4508
rect 1627 4504 1628 4508
rect 1622 4503 1628 4504
rect 1814 4508 1820 4509
rect 1814 4504 1815 4508
rect 1819 4504 1820 4508
rect 1934 4505 1935 4509
rect 1939 4505 1940 4509
rect 1934 4504 1940 4505
rect 1814 4503 1820 4504
rect 418 4493 424 4494
rect 110 4492 116 4493
rect 110 4488 111 4492
rect 115 4488 116 4492
rect 418 4489 419 4493
rect 423 4489 424 4493
rect 418 4488 424 4489
rect 594 4493 600 4494
rect 594 4489 595 4493
rect 599 4489 600 4493
rect 594 4488 600 4489
rect 778 4493 784 4494
rect 778 4489 779 4493
rect 783 4489 784 4493
rect 778 4488 784 4489
rect 970 4493 976 4494
rect 970 4489 971 4493
rect 975 4489 976 4493
rect 970 4488 976 4489
rect 1170 4493 1176 4494
rect 1170 4489 1171 4493
rect 1175 4489 1176 4493
rect 1170 4488 1176 4489
rect 1378 4493 1384 4494
rect 1378 4489 1379 4493
rect 1383 4489 1384 4493
rect 1378 4488 1384 4489
rect 1594 4493 1600 4494
rect 1594 4489 1595 4493
rect 1599 4489 1600 4493
rect 1594 4488 1600 4489
rect 1786 4493 1792 4494
rect 1786 4489 1787 4493
rect 1791 4489 1792 4493
rect 1786 4488 1792 4489
rect 1934 4492 1940 4493
rect 1934 4488 1935 4492
rect 1939 4488 1940 4492
rect 110 4487 116 4488
rect 112 4423 114 4487
rect 420 4423 422 4488
rect 596 4423 598 4488
rect 780 4423 782 4488
rect 972 4423 974 4488
rect 1172 4423 1174 4488
rect 1380 4423 1382 4488
rect 1596 4423 1598 4488
rect 1788 4423 1790 4488
rect 1934 4487 1940 4488
rect 1936 4423 1938 4487
rect 1976 4473 1978 4533
rect 1974 4472 1980 4473
rect 1996 4472 1998 4533
rect 2228 4472 2230 4533
rect 2460 4472 2462 4533
rect 2692 4472 2694 4533
rect 2916 4472 2918 4533
rect 3132 4472 3134 4533
rect 3356 4472 3358 4533
rect 3580 4472 3582 4533
rect 3800 4473 3802 4533
rect 3838 4531 3839 4535
rect 3843 4531 3844 4535
rect 4062 4532 4063 4536
rect 4067 4532 4068 4536
rect 4062 4531 4068 4532
rect 4358 4536 4364 4537
rect 4358 4532 4359 4536
rect 4363 4532 4364 4536
rect 4358 4531 4364 4532
rect 4654 4536 4660 4537
rect 4654 4532 4655 4536
rect 4659 4532 4660 4536
rect 4654 4531 4660 4532
rect 4958 4536 4964 4537
rect 4958 4532 4959 4536
rect 4963 4532 4964 4536
rect 4958 4531 4964 4532
rect 5262 4536 5268 4537
rect 5262 4532 5263 4536
rect 5267 4532 5268 4536
rect 5262 4531 5268 4532
rect 5542 4536 5548 4537
rect 5542 4532 5543 4536
rect 5547 4532 5548 4536
rect 5542 4531 5548 4532
rect 5662 4535 5668 4536
rect 5662 4531 5663 4535
rect 5667 4531 5668 4535
rect 3838 4530 3844 4531
rect 3840 4491 3842 4530
rect 4064 4491 4066 4531
rect 4360 4491 4362 4531
rect 4656 4491 4658 4531
rect 4960 4491 4962 4531
rect 5264 4491 5266 4531
rect 5544 4491 5546 4531
rect 5662 4530 5668 4531
rect 5664 4491 5666 4530
rect 3839 4490 3843 4491
rect 3839 4485 3843 4486
rect 4063 4490 4067 4491
rect 4063 4485 4067 4486
rect 4311 4490 4315 4491
rect 4311 4485 4315 4486
rect 4359 4490 4363 4491
rect 4359 4485 4363 4486
rect 4535 4490 4539 4491
rect 4535 4485 4539 4486
rect 4655 4490 4659 4491
rect 4655 4485 4659 4486
rect 4775 4490 4779 4491
rect 4775 4485 4779 4486
rect 4959 4490 4963 4491
rect 4959 4485 4963 4486
rect 5023 4490 5027 4491
rect 5023 4485 5027 4486
rect 5263 4490 5267 4491
rect 5263 4485 5267 4486
rect 5279 4490 5283 4491
rect 5279 4485 5283 4486
rect 5543 4490 5547 4491
rect 5543 4485 5547 4486
rect 5663 4490 5667 4491
rect 5663 4485 5667 4486
rect 3798 4472 3804 4473
rect 1974 4468 1975 4472
rect 1979 4468 1980 4472
rect 1974 4467 1980 4468
rect 1994 4471 2000 4472
rect 1994 4467 1995 4471
rect 1999 4467 2000 4471
rect 1994 4466 2000 4467
rect 2226 4471 2232 4472
rect 2226 4467 2227 4471
rect 2231 4467 2232 4471
rect 2226 4466 2232 4467
rect 2458 4471 2464 4472
rect 2458 4467 2459 4471
rect 2463 4467 2464 4471
rect 2458 4466 2464 4467
rect 2690 4471 2696 4472
rect 2690 4467 2691 4471
rect 2695 4467 2696 4471
rect 2690 4466 2696 4467
rect 2914 4471 2920 4472
rect 2914 4467 2915 4471
rect 2919 4467 2920 4471
rect 2914 4466 2920 4467
rect 3130 4471 3136 4472
rect 3130 4467 3131 4471
rect 3135 4467 3136 4471
rect 3130 4466 3136 4467
rect 3354 4471 3360 4472
rect 3354 4467 3355 4471
rect 3359 4467 3360 4471
rect 3354 4466 3360 4467
rect 3578 4471 3584 4472
rect 3578 4467 3579 4471
rect 3583 4467 3584 4471
rect 3798 4468 3799 4472
rect 3803 4468 3804 4472
rect 3798 4467 3804 4468
rect 3578 4466 3584 4467
rect 3840 4462 3842 4485
rect 3838 4461 3844 4462
rect 4312 4461 4314 4485
rect 4536 4461 4538 4485
rect 4776 4461 4778 4485
rect 5024 4461 5026 4485
rect 5280 4461 5282 4485
rect 5544 4461 5546 4485
rect 5664 4462 5666 4485
rect 5662 4461 5668 4462
rect 3838 4457 3839 4461
rect 3843 4457 3844 4461
rect 2022 4456 2028 4457
rect 1974 4455 1980 4456
rect 1974 4451 1975 4455
rect 1979 4451 1980 4455
rect 2022 4452 2023 4456
rect 2027 4452 2028 4456
rect 2022 4451 2028 4452
rect 2254 4456 2260 4457
rect 2254 4452 2255 4456
rect 2259 4452 2260 4456
rect 2254 4451 2260 4452
rect 2486 4456 2492 4457
rect 2486 4452 2487 4456
rect 2491 4452 2492 4456
rect 2486 4451 2492 4452
rect 2718 4456 2724 4457
rect 2718 4452 2719 4456
rect 2723 4452 2724 4456
rect 2718 4451 2724 4452
rect 2942 4456 2948 4457
rect 2942 4452 2943 4456
rect 2947 4452 2948 4456
rect 2942 4451 2948 4452
rect 3158 4456 3164 4457
rect 3158 4452 3159 4456
rect 3163 4452 3164 4456
rect 3158 4451 3164 4452
rect 3382 4456 3388 4457
rect 3382 4452 3383 4456
rect 3387 4452 3388 4456
rect 3382 4451 3388 4452
rect 3606 4456 3612 4457
rect 3838 4456 3844 4457
rect 4310 4460 4316 4461
rect 4310 4456 4311 4460
rect 4315 4456 4316 4460
rect 3606 4452 3607 4456
rect 3611 4452 3612 4456
rect 3606 4451 3612 4452
rect 3798 4455 3804 4456
rect 4310 4455 4316 4456
rect 4534 4460 4540 4461
rect 4534 4456 4535 4460
rect 4539 4456 4540 4460
rect 4534 4455 4540 4456
rect 4774 4460 4780 4461
rect 4774 4456 4775 4460
rect 4779 4456 4780 4460
rect 4774 4455 4780 4456
rect 5022 4460 5028 4461
rect 5022 4456 5023 4460
rect 5027 4456 5028 4460
rect 5022 4455 5028 4456
rect 5278 4460 5284 4461
rect 5278 4456 5279 4460
rect 5283 4456 5284 4460
rect 5278 4455 5284 4456
rect 5542 4460 5548 4461
rect 5542 4456 5543 4460
rect 5547 4456 5548 4460
rect 5662 4457 5663 4461
rect 5667 4457 5668 4461
rect 5662 4456 5668 4457
rect 5542 4455 5548 4456
rect 3798 4451 3799 4455
rect 3803 4451 3804 4455
rect 1974 4450 1980 4451
rect 1976 4423 1978 4450
rect 2024 4423 2026 4451
rect 2256 4423 2258 4451
rect 2488 4423 2490 4451
rect 2720 4423 2722 4451
rect 2944 4423 2946 4451
rect 3160 4423 3162 4451
rect 3384 4423 3386 4451
rect 3608 4423 3610 4451
rect 3798 4450 3804 4451
rect 3800 4423 3802 4450
rect 4282 4445 4288 4446
rect 3838 4444 3844 4445
rect 3838 4440 3839 4444
rect 3843 4440 3844 4444
rect 4282 4441 4283 4445
rect 4287 4441 4288 4445
rect 4282 4440 4288 4441
rect 4506 4445 4512 4446
rect 4506 4441 4507 4445
rect 4511 4441 4512 4445
rect 4506 4440 4512 4441
rect 4746 4445 4752 4446
rect 4746 4441 4747 4445
rect 4751 4441 4752 4445
rect 4746 4440 4752 4441
rect 4994 4445 5000 4446
rect 4994 4441 4995 4445
rect 4999 4441 5000 4445
rect 4994 4440 5000 4441
rect 5250 4445 5256 4446
rect 5250 4441 5251 4445
rect 5255 4441 5256 4445
rect 5250 4440 5256 4441
rect 5514 4445 5520 4446
rect 5514 4441 5515 4445
rect 5519 4441 5520 4445
rect 5514 4440 5520 4441
rect 5662 4444 5668 4445
rect 5662 4440 5663 4444
rect 5667 4440 5668 4444
rect 3838 4439 3844 4440
rect 111 4422 115 4423
rect 111 4417 115 4418
rect 419 4422 423 4423
rect 419 4417 423 4418
rect 571 4422 575 4423
rect 571 4417 575 4418
rect 595 4422 599 4423
rect 595 4417 599 4418
rect 739 4422 743 4423
rect 739 4417 743 4418
rect 779 4422 783 4423
rect 779 4417 783 4418
rect 915 4422 919 4423
rect 915 4417 919 4418
rect 971 4422 975 4423
rect 971 4417 975 4418
rect 1107 4422 1111 4423
rect 1107 4417 1111 4418
rect 1171 4422 1175 4423
rect 1171 4417 1175 4418
rect 1299 4422 1303 4423
rect 1299 4417 1303 4418
rect 1379 4422 1383 4423
rect 1379 4417 1383 4418
rect 1499 4422 1503 4423
rect 1499 4417 1503 4418
rect 1595 4422 1599 4423
rect 1595 4417 1599 4418
rect 1707 4422 1711 4423
rect 1707 4417 1711 4418
rect 1787 4422 1791 4423
rect 1787 4417 1791 4418
rect 1935 4422 1939 4423
rect 1935 4417 1939 4418
rect 1975 4422 1979 4423
rect 1975 4417 1979 4418
rect 2023 4422 2027 4423
rect 2023 4417 2027 4418
rect 2119 4422 2123 4423
rect 2119 4417 2123 4418
rect 2255 4422 2259 4423
rect 2255 4417 2259 4418
rect 2343 4422 2347 4423
rect 2343 4417 2347 4418
rect 2487 4422 2491 4423
rect 2487 4417 2491 4418
rect 2567 4422 2571 4423
rect 2567 4417 2571 4418
rect 2719 4422 2723 4423
rect 2719 4417 2723 4418
rect 2783 4422 2787 4423
rect 2783 4417 2787 4418
rect 2943 4422 2947 4423
rect 2943 4417 2947 4418
rect 2991 4422 2995 4423
rect 2991 4417 2995 4418
rect 3159 4422 3163 4423
rect 3159 4417 3163 4418
rect 3199 4422 3203 4423
rect 3199 4417 3203 4418
rect 3383 4422 3387 4423
rect 3383 4417 3387 4418
rect 3407 4422 3411 4423
rect 3407 4417 3411 4418
rect 3607 4422 3611 4423
rect 3607 4417 3611 4418
rect 3799 4422 3803 4423
rect 3799 4417 3803 4418
rect 112 4357 114 4417
rect 110 4356 116 4357
rect 572 4356 574 4417
rect 740 4356 742 4417
rect 916 4356 918 4417
rect 1108 4356 1110 4417
rect 1300 4356 1302 4417
rect 1500 4356 1502 4417
rect 1708 4356 1710 4417
rect 1936 4357 1938 4417
rect 1976 4394 1978 4417
rect 1974 4393 1980 4394
rect 2120 4393 2122 4417
rect 2344 4393 2346 4417
rect 2568 4393 2570 4417
rect 2784 4393 2786 4417
rect 2992 4393 2994 4417
rect 3200 4393 3202 4417
rect 3408 4393 3410 4417
rect 3800 4394 3802 4417
rect 3798 4393 3804 4394
rect 1974 4389 1975 4393
rect 1979 4389 1980 4393
rect 1974 4388 1980 4389
rect 2118 4392 2124 4393
rect 2118 4388 2119 4392
rect 2123 4388 2124 4392
rect 2118 4387 2124 4388
rect 2342 4392 2348 4393
rect 2342 4388 2343 4392
rect 2347 4388 2348 4392
rect 2342 4387 2348 4388
rect 2566 4392 2572 4393
rect 2566 4388 2567 4392
rect 2571 4388 2572 4392
rect 2566 4387 2572 4388
rect 2782 4392 2788 4393
rect 2782 4388 2783 4392
rect 2787 4388 2788 4392
rect 2782 4387 2788 4388
rect 2990 4392 2996 4393
rect 2990 4388 2991 4392
rect 2995 4388 2996 4392
rect 2990 4387 2996 4388
rect 3198 4392 3204 4393
rect 3198 4388 3199 4392
rect 3203 4388 3204 4392
rect 3198 4387 3204 4388
rect 3406 4392 3412 4393
rect 3406 4388 3407 4392
rect 3411 4388 3412 4392
rect 3798 4389 3799 4393
rect 3803 4389 3804 4393
rect 3798 4388 3804 4389
rect 3406 4387 3412 4388
rect 2090 4377 2096 4378
rect 1974 4376 1980 4377
rect 1974 4372 1975 4376
rect 1979 4372 1980 4376
rect 2090 4373 2091 4377
rect 2095 4373 2096 4377
rect 2090 4372 2096 4373
rect 2314 4377 2320 4378
rect 2314 4373 2315 4377
rect 2319 4373 2320 4377
rect 2314 4372 2320 4373
rect 2538 4377 2544 4378
rect 2538 4373 2539 4377
rect 2543 4373 2544 4377
rect 2538 4372 2544 4373
rect 2754 4377 2760 4378
rect 2754 4373 2755 4377
rect 2759 4373 2760 4377
rect 2754 4372 2760 4373
rect 2962 4377 2968 4378
rect 2962 4373 2963 4377
rect 2967 4373 2968 4377
rect 2962 4372 2968 4373
rect 3170 4377 3176 4378
rect 3170 4373 3171 4377
rect 3175 4373 3176 4377
rect 3170 4372 3176 4373
rect 3378 4377 3384 4378
rect 3378 4373 3379 4377
rect 3383 4373 3384 4377
rect 3378 4372 3384 4373
rect 3798 4376 3804 4377
rect 3798 4372 3799 4376
rect 3803 4372 3804 4376
rect 1974 4371 1980 4372
rect 1934 4356 1940 4357
rect 110 4352 111 4356
rect 115 4352 116 4356
rect 110 4351 116 4352
rect 570 4355 576 4356
rect 570 4351 571 4355
rect 575 4351 576 4355
rect 570 4350 576 4351
rect 738 4355 744 4356
rect 738 4351 739 4355
rect 743 4351 744 4355
rect 738 4350 744 4351
rect 914 4355 920 4356
rect 914 4351 915 4355
rect 919 4351 920 4355
rect 914 4350 920 4351
rect 1106 4355 1112 4356
rect 1106 4351 1107 4355
rect 1111 4351 1112 4355
rect 1106 4350 1112 4351
rect 1298 4355 1304 4356
rect 1298 4351 1299 4355
rect 1303 4351 1304 4355
rect 1298 4350 1304 4351
rect 1498 4355 1504 4356
rect 1498 4351 1499 4355
rect 1503 4351 1504 4355
rect 1498 4350 1504 4351
rect 1706 4355 1712 4356
rect 1706 4351 1707 4355
rect 1711 4351 1712 4355
rect 1934 4352 1935 4356
rect 1939 4352 1940 4356
rect 1934 4351 1940 4352
rect 1706 4350 1712 4351
rect 598 4340 604 4341
rect 110 4339 116 4340
rect 110 4335 111 4339
rect 115 4335 116 4339
rect 598 4336 599 4340
rect 603 4336 604 4340
rect 598 4335 604 4336
rect 766 4340 772 4341
rect 766 4336 767 4340
rect 771 4336 772 4340
rect 766 4335 772 4336
rect 942 4340 948 4341
rect 942 4336 943 4340
rect 947 4336 948 4340
rect 942 4335 948 4336
rect 1134 4340 1140 4341
rect 1134 4336 1135 4340
rect 1139 4336 1140 4340
rect 1134 4335 1140 4336
rect 1326 4340 1332 4341
rect 1326 4336 1327 4340
rect 1331 4336 1332 4340
rect 1326 4335 1332 4336
rect 1526 4340 1532 4341
rect 1526 4336 1527 4340
rect 1531 4336 1532 4340
rect 1526 4335 1532 4336
rect 1734 4340 1740 4341
rect 1734 4336 1735 4340
rect 1739 4336 1740 4340
rect 1734 4335 1740 4336
rect 1934 4339 1940 4340
rect 1934 4335 1935 4339
rect 1939 4335 1940 4339
rect 110 4334 116 4335
rect 112 4311 114 4334
rect 600 4311 602 4335
rect 768 4311 770 4335
rect 944 4311 946 4335
rect 1136 4311 1138 4335
rect 1328 4311 1330 4335
rect 1528 4311 1530 4335
rect 1736 4311 1738 4335
rect 1934 4334 1940 4335
rect 1936 4311 1938 4334
rect 111 4310 115 4311
rect 111 4305 115 4306
rect 599 4310 603 4311
rect 599 4305 603 4306
rect 655 4310 659 4311
rect 655 4305 659 4306
rect 767 4310 771 4311
rect 767 4305 771 4306
rect 823 4310 827 4311
rect 823 4305 827 4306
rect 943 4310 947 4311
rect 943 4305 947 4306
rect 991 4310 995 4311
rect 991 4305 995 4306
rect 1135 4310 1139 4311
rect 1135 4305 1139 4306
rect 1167 4310 1171 4311
rect 1167 4305 1171 4306
rect 1327 4310 1331 4311
rect 1327 4305 1331 4306
rect 1343 4310 1347 4311
rect 1343 4305 1347 4306
rect 1519 4310 1523 4311
rect 1519 4305 1523 4306
rect 1527 4310 1531 4311
rect 1527 4305 1531 4306
rect 1703 4310 1707 4311
rect 1703 4305 1707 4306
rect 1735 4310 1739 4311
rect 1735 4305 1739 4306
rect 1935 4310 1939 4311
rect 1935 4305 1939 4306
rect 112 4282 114 4305
rect 110 4281 116 4282
rect 656 4281 658 4305
rect 824 4281 826 4305
rect 992 4281 994 4305
rect 1168 4281 1170 4305
rect 1344 4281 1346 4305
rect 1520 4281 1522 4305
rect 1704 4281 1706 4305
rect 1936 4282 1938 4305
rect 1976 4303 1978 4371
rect 2092 4303 2094 4372
rect 2316 4303 2318 4372
rect 2540 4303 2542 4372
rect 2756 4303 2758 4372
rect 2964 4303 2966 4372
rect 3172 4303 3174 4372
rect 3380 4303 3382 4372
rect 3798 4371 3804 4372
rect 3800 4303 3802 4371
rect 3840 4359 3842 4439
rect 4284 4359 4286 4440
rect 4508 4359 4510 4440
rect 4748 4359 4750 4440
rect 4996 4359 4998 4440
rect 5252 4359 5254 4440
rect 5516 4359 5518 4440
rect 5662 4439 5668 4440
rect 5664 4359 5666 4439
rect 3839 4358 3843 4359
rect 3839 4353 3843 4354
rect 4283 4358 4287 4359
rect 4283 4353 4287 4354
rect 4507 4358 4511 4359
rect 4507 4353 4511 4354
rect 4515 4358 4519 4359
rect 4515 4353 4519 4354
rect 4691 4358 4695 4359
rect 4691 4353 4695 4354
rect 4747 4358 4751 4359
rect 4747 4353 4751 4354
rect 4875 4358 4879 4359
rect 4875 4353 4879 4354
rect 4995 4358 4999 4359
rect 4995 4353 4999 4354
rect 5067 4358 5071 4359
rect 5067 4353 5071 4354
rect 5251 4358 5255 4359
rect 5251 4353 5255 4354
rect 5267 4358 5271 4359
rect 5267 4353 5271 4354
rect 5467 4358 5471 4359
rect 5467 4353 5471 4354
rect 5515 4358 5519 4359
rect 5515 4353 5519 4354
rect 5663 4358 5667 4359
rect 5663 4353 5667 4354
rect 1975 4302 1979 4303
rect 1975 4297 1979 4298
rect 2019 4302 2023 4303
rect 2019 4297 2023 4298
rect 2091 4302 2095 4303
rect 2091 4297 2095 4298
rect 2243 4302 2247 4303
rect 2243 4297 2247 4298
rect 2315 4302 2319 4303
rect 2315 4297 2319 4298
rect 2459 4302 2463 4303
rect 2459 4297 2463 4298
rect 2539 4302 2543 4303
rect 2539 4297 2543 4298
rect 2667 4302 2671 4303
rect 2667 4297 2671 4298
rect 2755 4302 2759 4303
rect 2755 4297 2759 4298
rect 2875 4302 2879 4303
rect 2875 4297 2879 4298
rect 2963 4302 2967 4303
rect 2963 4297 2967 4298
rect 3083 4302 3087 4303
rect 3083 4297 3087 4298
rect 3171 4302 3175 4303
rect 3171 4297 3175 4298
rect 3291 4302 3295 4303
rect 3291 4297 3295 4298
rect 3379 4302 3383 4303
rect 3379 4297 3383 4298
rect 3799 4302 3803 4303
rect 3799 4297 3803 4298
rect 1934 4281 1940 4282
rect 110 4277 111 4281
rect 115 4277 116 4281
rect 110 4276 116 4277
rect 654 4280 660 4281
rect 654 4276 655 4280
rect 659 4276 660 4280
rect 654 4275 660 4276
rect 822 4280 828 4281
rect 822 4276 823 4280
rect 827 4276 828 4280
rect 822 4275 828 4276
rect 990 4280 996 4281
rect 990 4276 991 4280
rect 995 4276 996 4280
rect 990 4275 996 4276
rect 1166 4280 1172 4281
rect 1166 4276 1167 4280
rect 1171 4276 1172 4280
rect 1166 4275 1172 4276
rect 1342 4280 1348 4281
rect 1342 4276 1343 4280
rect 1347 4276 1348 4280
rect 1342 4275 1348 4276
rect 1518 4280 1524 4281
rect 1518 4276 1519 4280
rect 1523 4276 1524 4280
rect 1518 4275 1524 4276
rect 1702 4280 1708 4281
rect 1702 4276 1703 4280
rect 1707 4276 1708 4280
rect 1934 4277 1935 4281
rect 1939 4277 1940 4281
rect 1934 4276 1940 4277
rect 1702 4275 1708 4276
rect 626 4265 632 4266
rect 110 4264 116 4265
rect 110 4260 111 4264
rect 115 4260 116 4264
rect 626 4261 627 4265
rect 631 4261 632 4265
rect 626 4260 632 4261
rect 794 4265 800 4266
rect 794 4261 795 4265
rect 799 4261 800 4265
rect 794 4260 800 4261
rect 962 4265 968 4266
rect 962 4261 963 4265
rect 967 4261 968 4265
rect 962 4260 968 4261
rect 1138 4265 1144 4266
rect 1138 4261 1139 4265
rect 1143 4261 1144 4265
rect 1138 4260 1144 4261
rect 1314 4265 1320 4266
rect 1314 4261 1315 4265
rect 1319 4261 1320 4265
rect 1314 4260 1320 4261
rect 1490 4265 1496 4266
rect 1490 4261 1491 4265
rect 1495 4261 1496 4265
rect 1490 4260 1496 4261
rect 1674 4265 1680 4266
rect 1674 4261 1675 4265
rect 1679 4261 1680 4265
rect 1674 4260 1680 4261
rect 1934 4264 1940 4265
rect 1934 4260 1935 4264
rect 1939 4260 1940 4264
rect 110 4259 116 4260
rect 112 4187 114 4259
rect 628 4187 630 4260
rect 796 4187 798 4260
rect 964 4187 966 4260
rect 1140 4187 1142 4260
rect 1316 4187 1318 4260
rect 1492 4187 1494 4260
rect 1676 4187 1678 4260
rect 1934 4259 1940 4260
rect 1936 4187 1938 4259
rect 1976 4237 1978 4297
rect 1974 4236 1980 4237
rect 2020 4236 2022 4297
rect 2244 4236 2246 4297
rect 2460 4236 2462 4297
rect 2668 4236 2670 4297
rect 2876 4236 2878 4297
rect 3084 4236 3086 4297
rect 3292 4236 3294 4297
rect 3800 4237 3802 4297
rect 3840 4293 3842 4353
rect 3838 4292 3844 4293
rect 4516 4292 4518 4353
rect 4692 4292 4694 4353
rect 4876 4292 4878 4353
rect 5068 4292 5070 4353
rect 5268 4292 5270 4353
rect 5468 4292 5470 4353
rect 5664 4293 5666 4353
rect 5662 4292 5668 4293
rect 3838 4288 3839 4292
rect 3843 4288 3844 4292
rect 3838 4287 3844 4288
rect 4514 4291 4520 4292
rect 4514 4287 4515 4291
rect 4519 4287 4520 4291
rect 4514 4286 4520 4287
rect 4690 4291 4696 4292
rect 4690 4287 4691 4291
rect 4695 4287 4696 4291
rect 4690 4286 4696 4287
rect 4874 4291 4880 4292
rect 4874 4287 4875 4291
rect 4879 4287 4880 4291
rect 4874 4286 4880 4287
rect 5066 4291 5072 4292
rect 5066 4287 5067 4291
rect 5071 4287 5072 4291
rect 5066 4286 5072 4287
rect 5266 4291 5272 4292
rect 5266 4287 5267 4291
rect 5271 4287 5272 4291
rect 5266 4286 5272 4287
rect 5466 4291 5472 4292
rect 5466 4287 5467 4291
rect 5471 4287 5472 4291
rect 5662 4288 5663 4292
rect 5667 4288 5668 4292
rect 5662 4287 5668 4288
rect 5466 4286 5472 4287
rect 4542 4276 4548 4277
rect 3838 4275 3844 4276
rect 3838 4271 3839 4275
rect 3843 4271 3844 4275
rect 4542 4272 4543 4276
rect 4547 4272 4548 4276
rect 4542 4271 4548 4272
rect 4718 4276 4724 4277
rect 4718 4272 4719 4276
rect 4723 4272 4724 4276
rect 4718 4271 4724 4272
rect 4902 4276 4908 4277
rect 4902 4272 4903 4276
rect 4907 4272 4908 4276
rect 4902 4271 4908 4272
rect 5094 4276 5100 4277
rect 5094 4272 5095 4276
rect 5099 4272 5100 4276
rect 5094 4271 5100 4272
rect 5294 4276 5300 4277
rect 5294 4272 5295 4276
rect 5299 4272 5300 4276
rect 5294 4271 5300 4272
rect 5494 4276 5500 4277
rect 5494 4272 5495 4276
rect 5499 4272 5500 4276
rect 5494 4271 5500 4272
rect 5662 4275 5668 4276
rect 5662 4271 5663 4275
rect 5667 4271 5668 4275
rect 3838 4270 3844 4271
rect 3798 4236 3804 4237
rect 1974 4232 1975 4236
rect 1979 4232 1980 4236
rect 1974 4231 1980 4232
rect 2018 4235 2024 4236
rect 2018 4231 2019 4235
rect 2023 4231 2024 4235
rect 2018 4230 2024 4231
rect 2242 4235 2248 4236
rect 2242 4231 2243 4235
rect 2247 4231 2248 4235
rect 2242 4230 2248 4231
rect 2458 4235 2464 4236
rect 2458 4231 2459 4235
rect 2463 4231 2464 4235
rect 2458 4230 2464 4231
rect 2666 4235 2672 4236
rect 2666 4231 2667 4235
rect 2671 4231 2672 4235
rect 2666 4230 2672 4231
rect 2874 4235 2880 4236
rect 2874 4231 2875 4235
rect 2879 4231 2880 4235
rect 2874 4230 2880 4231
rect 3082 4235 3088 4236
rect 3082 4231 3083 4235
rect 3087 4231 3088 4235
rect 3082 4230 3088 4231
rect 3290 4235 3296 4236
rect 3290 4231 3291 4235
rect 3295 4231 3296 4235
rect 3798 4232 3799 4236
rect 3803 4232 3804 4236
rect 3798 4231 3804 4232
rect 3290 4230 3296 4231
rect 3840 4227 3842 4270
rect 4544 4227 4546 4271
rect 4720 4227 4722 4271
rect 4904 4227 4906 4271
rect 5096 4227 5098 4271
rect 5296 4227 5298 4271
rect 5496 4227 5498 4271
rect 5662 4270 5668 4271
rect 5664 4227 5666 4270
rect 3839 4226 3843 4227
rect 3839 4221 3843 4222
rect 4543 4226 4547 4227
rect 4543 4221 4547 4222
rect 4719 4226 4723 4227
rect 4719 4221 4723 4222
rect 4815 4226 4819 4227
rect 4815 4221 4819 4222
rect 4903 4226 4907 4227
rect 4903 4221 4907 4222
rect 4951 4226 4955 4227
rect 4951 4221 4955 4222
rect 5087 4226 5091 4227
rect 5087 4221 5091 4222
rect 5095 4226 5099 4227
rect 5095 4221 5099 4222
rect 5223 4226 5227 4227
rect 5223 4221 5227 4222
rect 5295 4226 5299 4227
rect 5295 4221 5299 4222
rect 5359 4226 5363 4227
rect 5359 4221 5363 4222
rect 5495 4226 5499 4227
rect 5495 4221 5499 4222
rect 5663 4226 5667 4227
rect 5663 4221 5667 4222
rect 2046 4220 2052 4221
rect 1974 4219 1980 4220
rect 1974 4215 1975 4219
rect 1979 4215 1980 4219
rect 2046 4216 2047 4220
rect 2051 4216 2052 4220
rect 2046 4215 2052 4216
rect 2270 4220 2276 4221
rect 2270 4216 2271 4220
rect 2275 4216 2276 4220
rect 2270 4215 2276 4216
rect 2486 4220 2492 4221
rect 2486 4216 2487 4220
rect 2491 4216 2492 4220
rect 2486 4215 2492 4216
rect 2694 4220 2700 4221
rect 2694 4216 2695 4220
rect 2699 4216 2700 4220
rect 2694 4215 2700 4216
rect 2902 4220 2908 4221
rect 2902 4216 2903 4220
rect 2907 4216 2908 4220
rect 2902 4215 2908 4216
rect 3110 4220 3116 4221
rect 3110 4216 3111 4220
rect 3115 4216 3116 4220
rect 3110 4215 3116 4216
rect 3318 4220 3324 4221
rect 3318 4216 3319 4220
rect 3323 4216 3324 4220
rect 3318 4215 3324 4216
rect 3798 4219 3804 4220
rect 3798 4215 3799 4219
rect 3803 4215 3804 4219
rect 1974 4214 1980 4215
rect 1976 4187 1978 4214
rect 2048 4187 2050 4215
rect 2272 4187 2274 4215
rect 2488 4187 2490 4215
rect 2696 4187 2698 4215
rect 2904 4187 2906 4215
rect 3112 4187 3114 4215
rect 3320 4187 3322 4215
rect 3798 4214 3804 4215
rect 3800 4187 3802 4214
rect 3840 4198 3842 4221
rect 3838 4197 3844 4198
rect 4816 4197 4818 4221
rect 4952 4197 4954 4221
rect 5088 4197 5090 4221
rect 5224 4197 5226 4221
rect 5360 4197 5362 4221
rect 5496 4197 5498 4221
rect 5664 4198 5666 4221
rect 5662 4197 5668 4198
rect 3838 4193 3839 4197
rect 3843 4193 3844 4197
rect 3838 4192 3844 4193
rect 4814 4196 4820 4197
rect 4814 4192 4815 4196
rect 4819 4192 4820 4196
rect 4814 4191 4820 4192
rect 4950 4196 4956 4197
rect 4950 4192 4951 4196
rect 4955 4192 4956 4196
rect 4950 4191 4956 4192
rect 5086 4196 5092 4197
rect 5086 4192 5087 4196
rect 5091 4192 5092 4196
rect 5086 4191 5092 4192
rect 5222 4196 5228 4197
rect 5222 4192 5223 4196
rect 5227 4192 5228 4196
rect 5222 4191 5228 4192
rect 5358 4196 5364 4197
rect 5358 4192 5359 4196
rect 5363 4192 5364 4196
rect 5358 4191 5364 4192
rect 5494 4196 5500 4197
rect 5494 4192 5495 4196
rect 5499 4192 5500 4196
rect 5662 4193 5663 4197
rect 5667 4193 5668 4197
rect 5662 4192 5668 4193
rect 5494 4191 5500 4192
rect 111 4186 115 4187
rect 111 4181 115 4182
rect 347 4186 351 4187
rect 347 4181 351 4182
rect 515 4186 519 4187
rect 515 4181 519 4182
rect 627 4186 631 4187
rect 627 4181 631 4182
rect 699 4186 703 4187
rect 699 4181 703 4182
rect 795 4186 799 4187
rect 795 4181 799 4182
rect 891 4186 895 4187
rect 891 4181 895 4182
rect 963 4186 967 4187
rect 963 4181 967 4182
rect 1099 4186 1103 4187
rect 1099 4181 1103 4182
rect 1139 4186 1143 4187
rect 1139 4181 1143 4182
rect 1315 4186 1319 4187
rect 1315 4181 1319 4182
rect 1491 4186 1495 4187
rect 1491 4181 1495 4182
rect 1531 4186 1535 4187
rect 1531 4181 1535 4182
rect 1675 4186 1679 4187
rect 1675 4181 1679 4182
rect 1935 4186 1939 4187
rect 1935 4181 1939 4182
rect 1975 4186 1979 4187
rect 1975 4181 1979 4182
rect 2023 4186 2027 4187
rect 2023 4181 2027 4182
rect 2047 4186 2051 4187
rect 2047 4181 2051 4182
rect 2271 4186 2275 4187
rect 2271 4181 2275 4182
rect 2287 4186 2291 4187
rect 2287 4181 2291 4182
rect 2487 4186 2491 4187
rect 2487 4181 2491 4182
rect 2551 4186 2555 4187
rect 2551 4181 2555 4182
rect 2695 4186 2699 4187
rect 2695 4181 2699 4182
rect 2799 4186 2803 4187
rect 2799 4181 2803 4182
rect 2903 4186 2907 4187
rect 2903 4181 2907 4182
rect 3039 4186 3043 4187
rect 3039 4181 3043 4182
rect 3111 4186 3115 4187
rect 3111 4181 3115 4182
rect 3279 4186 3283 4187
rect 3279 4181 3283 4182
rect 3319 4186 3323 4187
rect 3319 4181 3323 4182
rect 3519 4186 3523 4187
rect 3519 4181 3523 4182
rect 3799 4186 3803 4187
rect 3799 4181 3803 4182
rect 4786 4181 4792 4182
rect 112 4121 114 4181
rect 110 4120 116 4121
rect 348 4120 350 4181
rect 516 4120 518 4181
rect 700 4120 702 4181
rect 892 4120 894 4181
rect 1100 4120 1102 4181
rect 1316 4120 1318 4181
rect 1532 4120 1534 4181
rect 1936 4121 1938 4181
rect 1976 4158 1978 4181
rect 1974 4157 1980 4158
rect 2024 4157 2026 4181
rect 2288 4157 2290 4181
rect 2552 4157 2554 4181
rect 2800 4157 2802 4181
rect 3040 4157 3042 4181
rect 3280 4157 3282 4181
rect 3520 4157 3522 4181
rect 3800 4158 3802 4181
rect 3838 4180 3844 4181
rect 3838 4176 3839 4180
rect 3843 4176 3844 4180
rect 4786 4177 4787 4181
rect 4791 4177 4792 4181
rect 4786 4176 4792 4177
rect 4922 4181 4928 4182
rect 4922 4177 4923 4181
rect 4927 4177 4928 4181
rect 4922 4176 4928 4177
rect 5058 4181 5064 4182
rect 5058 4177 5059 4181
rect 5063 4177 5064 4181
rect 5058 4176 5064 4177
rect 5194 4181 5200 4182
rect 5194 4177 5195 4181
rect 5199 4177 5200 4181
rect 5194 4176 5200 4177
rect 5330 4181 5336 4182
rect 5330 4177 5331 4181
rect 5335 4177 5336 4181
rect 5330 4176 5336 4177
rect 5466 4181 5472 4182
rect 5466 4177 5467 4181
rect 5471 4177 5472 4181
rect 5466 4176 5472 4177
rect 5662 4180 5668 4181
rect 5662 4176 5663 4180
rect 5667 4176 5668 4180
rect 3838 4175 3844 4176
rect 3798 4157 3804 4158
rect 1974 4153 1975 4157
rect 1979 4153 1980 4157
rect 1974 4152 1980 4153
rect 2022 4156 2028 4157
rect 2022 4152 2023 4156
rect 2027 4152 2028 4156
rect 2022 4151 2028 4152
rect 2286 4156 2292 4157
rect 2286 4152 2287 4156
rect 2291 4152 2292 4156
rect 2286 4151 2292 4152
rect 2550 4156 2556 4157
rect 2550 4152 2551 4156
rect 2555 4152 2556 4156
rect 2550 4151 2556 4152
rect 2798 4156 2804 4157
rect 2798 4152 2799 4156
rect 2803 4152 2804 4156
rect 2798 4151 2804 4152
rect 3038 4156 3044 4157
rect 3038 4152 3039 4156
rect 3043 4152 3044 4156
rect 3038 4151 3044 4152
rect 3278 4156 3284 4157
rect 3278 4152 3279 4156
rect 3283 4152 3284 4156
rect 3278 4151 3284 4152
rect 3518 4156 3524 4157
rect 3518 4152 3519 4156
rect 3523 4152 3524 4156
rect 3798 4153 3799 4157
rect 3803 4153 3804 4157
rect 3798 4152 3804 4153
rect 3518 4151 3524 4152
rect 1994 4141 2000 4142
rect 1974 4140 1980 4141
rect 1974 4136 1975 4140
rect 1979 4136 1980 4140
rect 1994 4137 1995 4141
rect 1999 4137 2000 4141
rect 1994 4136 2000 4137
rect 2258 4141 2264 4142
rect 2258 4137 2259 4141
rect 2263 4137 2264 4141
rect 2258 4136 2264 4137
rect 2522 4141 2528 4142
rect 2522 4137 2523 4141
rect 2527 4137 2528 4141
rect 2522 4136 2528 4137
rect 2770 4141 2776 4142
rect 2770 4137 2771 4141
rect 2775 4137 2776 4141
rect 2770 4136 2776 4137
rect 3010 4141 3016 4142
rect 3010 4137 3011 4141
rect 3015 4137 3016 4141
rect 3010 4136 3016 4137
rect 3250 4141 3256 4142
rect 3250 4137 3251 4141
rect 3255 4137 3256 4141
rect 3250 4136 3256 4137
rect 3490 4141 3496 4142
rect 3490 4137 3491 4141
rect 3495 4137 3496 4141
rect 3490 4136 3496 4137
rect 3798 4140 3804 4141
rect 3798 4136 3799 4140
rect 3803 4136 3804 4140
rect 1974 4135 1980 4136
rect 1934 4120 1940 4121
rect 110 4116 111 4120
rect 115 4116 116 4120
rect 110 4115 116 4116
rect 346 4119 352 4120
rect 346 4115 347 4119
rect 351 4115 352 4119
rect 346 4114 352 4115
rect 514 4119 520 4120
rect 514 4115 515 4119
rect 519 4115 520 4119
rect 514 4114 520 4115
rect 698 4119 704 4120
rect 698 4115 699 4119
rect 703 4115 704 4119
rect 698 4114 704 4115
rect 890 4119 896 4120
rect 890 4115 891 4119
rect 895 4115 896 4119
rect 890 4114 896 4115
rect 1098 4119 1104 4120
rect 1098 4115 1099 4119
rect 1103 4115 1104 4119
rect 1098 4114 1104 4115
rect 1314 4119 1320 4120
rect 1314 4115 1315 4119
rect 1319 4115 1320 4119
rect 1314 4114 1320 4115
rect 1530 4119 1536 4120
rect 1530 4115 1531 4119
rect 1535 4115 1536 4119
rect 1934 4116 1935 4120
rect 1939 4116 1940 4120
rect 1934 4115 1940 4116
rect 1530 4114 1536 4115
rect 374 4104 380 4105
rect 110 4103 116 4104
rect 110 4099 111 4103
rect 115 4099 116 4103
rect 374 4100 375 4104
rect 379 4100 380 4104
rect 374 4099 380 4100
rect 542 4104 548 4105
rect 542 4100 543 4104
rect 547 4100 548 4104
rect 542 4099 548 4100
rect 726 4104 732 4105
rect 726 4100 727 4104
rect 731 4100 732 4104
rect 726 4099 732 4100
rect 918 4104 924 4105
rect 918 4100 919 4104
rect 923 4100 924 4104
rect 918 4099 924 4100
rect 1126 4104 1132 4105
rect 1126 4100 1127 4104
rect 1131 4100 1132 4104
rect 1126 4099 1132 4100
rect 1342 4104 1348 4105
rect 1342 4100 1343 4104
rect 1347 4100 1348 4104
rect 1342 4099 1348 4100
rect 1558 4104 1564 4105
rect 1558 4100 1559 4104
rect 1563 4100 1564 4104
rect 1558 4099 1564 4100
rect 1934 4103 1940 4104
rect 1934 4099 1935 4103
rect 1939 4099 1940 4103
rect 110 4098 116 4099
rect 112 4059 114 4098
rect 376 4059 378 4099
rect 544 4059 546 4099
rect 728 4059 730 4099
rect 920 4059 922 4099
rect 1128 4059 1130 4099
rect 1344 4059 1346 4099
rect 1560 4059 1562 4099
rect 1934 4098 1940 4099
rect 1936 4059 1938 4098
rect 1976 4075 1978 4135
rect 1996 4075 1998 4136
rect 2260 4075 2262 4136
rect 2524 4075 2526 4136
rect 2772 4075 2774 4136
rect 3012 4075 3014 4136
rect 3252 4075 3254 4136
rect 3492 4075 3494 4136
rect 3798 4135 3804 4136
rect 3800 4075 3802 4135
rect 3840 4111 3842 4175
rect 4788 4111 4790 4176
rect 4924 4111 4926 4176
rect 5060 4111 5062 4176
rect 5196 4111 5198 4176
rect 5332 4111 5334 4176
rect 5468 4111 5470 4176
rect 5662 4175 5668 4176
rect 5664 4111 5666 4175
rect 3839 4110 3843 4111
rect 3839 4105 3843 4106
rect 4787 4110 4791 4111
rect 4787 4105 4791 4106
rect 4923 4110 4927 4111
rect 4923 4105 4927 4106
rect 4939 4110 4943 4111
rect 4939 4105 4943 4106
rect 5059 4110 5063 4111
rect 5059 4105 5063 4106
rect 5075 4110 5079 4111
rect 5075 4105 5079 4106
rect 5195 4110 5199 4111
rect 5195 4105 5199 4106
rect 5211 4110 5215 4111
rect 5211 4105 5215 4106
rect 5331 4110 5335 4111
rect 5331 4105 5335 4106
rect 5347 4110 5351 4111
rect 5347 4105 5351 4106
rect 5467 4110 5471 4111
rect 5467 4105 5471 4106
rect 5483 4110 5487 4111
rect 5483 4105 5487 4106
rect 5663 4110 5667 4111
rect 5663 4105 5667 4106
rect 1975 4074 1979 4075
rect 1975 4069 1979 4070
rect 1995 4074 1999 4075
rect 1995 4069 1999 4070
rect 2259 4074 2263 4075
rect 2259 4069 2263 4070
rect 2283 4074 2287 4075
rect 2283 4069 2287 4070
rect 2523 4074 2527 4075
rect 2523 4069 2527 4070
rect 2587 4074 2591 4075
rect 2587 4069 2591 4070
rect 2771 4074 2775 4075
rect 2771 4069 2775 4070
rect 2875 4074 2879 4075
rect 2875 4069 2879 4070
rect 3011 4074 3015 4075
rect 3011 4069 3015 4070
rect 3163 4074 3167 4075
rect 3163 4069 3167 4070
rect 3251 4074 3255 4075
rect 3251 4069 3255 4070
rect 3451 4074 3455 4075
rect 3451 4069 3455 4070
rect 3491 4074 3495 4075
rect 3491 4069 3495 4070
rect 3799 4074 3803 4075
rect 3799 4069 3803 4070
rect 111 4058 115 4059
rect 111 4053 115 4054
rect 231 4058 235 4059
rect 231 4053 235 4054
rect 375 4058 379 4059
rect 375 4053 379 4054
rect 423 4058 427 4059
rect 423 4053 427 4054
rect 543 4058 547 4059
rect 543 4053 547 4054
rect 615 4058 619 4059
rect 615 4053 619 4054
rect 727 4058 731 4059
rect 727 4053 731 4054
rect 807 4058 811 4059
rect 807 4053 811 4054
rect 919 4058 923 4059
rect 919 4053 923 4054
rect 991 4058 995 4059
rect 991 4053 995 4054
rect 1127 4058 1131 4059
rect 1127 4053 1131 4054
rect 1167 4058 1171 4059
rect 1167 4053 1171 4054
rect 1335 4058 1339 4059
rect 1335 4053 1339 4054
rect 1343 4058 1347 4059
rect 1343 4053 1347 4054
rect 1503 4058 1507 4059
rect 1503 4053 1507 4054
rect 1559 4058 1563 4059
rect 1559 4053 1563 4054
rect 1671 4058 1675 4059
rect 1671 4053 1675 4054
rect 1815 4058 1819 4059
rect 1815 4053 1819 4054
rect 1935 4058 1939 4059
rect 1935 4053 1939 4054
rect 112 4030 114 4053
rect 110 4029 116 4030
rect 232 4029 234 4053
rect 424 4029 426 4053
rect 616 4029 618 4053
rect 808 4029 810 4053
rect 992 4029 994 4053
rect 1168 4029 1170 4053
rect 1336 4029 1338 4053
rect 1504 4029 1506 4053
rect 1672 4029 1674 4053
rect 1816 4029 1818 4053
rect 1936 4030 1938 4053
rect 1934 4029 1940 4030
rect 110 4025 111 4029
rect 115 4025 116 4029
rect 110 4024 116 4025
rect 230 4028 236 4029
rect 230 4024 231 4028
rect 235 4024 236 4028
rect 230 4023 236 4024
rect 422 4028 428 4029
rect 422 4024 423 4028
rect 427 4024 428 4028
rect 422 4023 428 4024
rect 614 4028 620 4029
rect 614 4024 615 4028
rect 619 4024 620 4028
rect 614 4023 620 4024
rect 806 4028 812 4029
rect 806 4024 807 4028
rect 811 4024 812 4028
rect 806 4023 812 4024
rect 990 4028 996 4029
rect 990 4024 991 4028
rect 995 4024 996 4028
rect 990 4023 996 4024
rect 1166 4028 1172 4029
rect 1166 4024 1167 4028
rect 1171 4024 1172 4028
rect 1166 4023 1172 4024
rect 1334 4028 1340 4029
rect 1334 4024 1335 4028
rect 1339 4024 1340 4028
rect 1334 4023 1340 4024
rect 1502 4028 1508 4029
rect 1502 4024 1503 4028
rect 1507 4024 1508 4028
rect 1502 4023 1508 4024
rect 1670 4028 1676 4029
rect 1670 4024 1671 4028
rect 1675 4024 1676 4028
rect 1670 4023 1676 4024
rect 1814 4028 1820 4029
rect 1814 4024 1815 4028
rect 1819 4024 1820 4028
rect 1934 4025 1935 4029
rect 1939 4025 1940 4029
rect 1934 4024 1940 4025
rect 1814 4023 1820 4024
rect 202 4013 208 4014
rect 110 4012 116 4013
rect 110 4008 111 4012
rect 115 4008 116 4012
rect 202 4009 203 4013
rect 207 4009 208 4013
rect 202 4008 208 4009
rect 394 4013 400 4014
rect 394 4009 395 4013
rect 399 4009 400 4013
rect 394 4008 400 4009
rect 586 4013 592 4014
rect 586 4009 587 4013
rect 591 4009 592 4013
rect 586 4008 592 4009
rect 778 4013 784 4014
rect 778 4009 779 4013
rect 783 4009 784 4013
rect 778 4008 784 4009
rect 962 4013 968 4014
rect 962 4009 963 4013
rect 967 4009 968 4013
rect 962 4008 968 4009
rect 1138 4013 1144 4014
rect 1138 4009 1139 4013
rect 1143 4009 1144 4013
rect 1138 4008 1144 4009
rect 1306 4013 1312 4014
rect 1306 4009 1307 4013
rect 1311 4009 1312 4013
rect 1306 4008 1312 4009
rect 1474 4013 1480 4014
rect 1474 4009 1475 4013
rect 1479 4009 1480 4013
rect 1474 4008 1480 4009
rect 1642 4013 1648 4014
rect 1642 4009 1643 4013
rect 1647 4009 1648 4013
rect 1642 4008 1648 4009
rect 1786 4013 1792 4014
rect 1786 4009 1787 4013
rect 1791 4009 1792 4013
rect 1786 4008 1792 4009
rect 1934 4012 1940 4013
rect 1934 4008 1935 4012
rect 1939 4008 1940 4012
rect 1976 4009 1978 4069
rect 110 4007 116 4008
rect 112 3947 114 4007
rect 204 3947 206 4008
rect 396 3947 398 4008
rect 588 3947 590 4008
rect 780 3947 782 4008
rect 964 3947 966 4008
rect 1140 3947 1142 4008
rect 1308 3947 1310 4008
rect 1476 3947 1478 4008
rect 1644 3947 1646 4008
rect 1788 3947 1790 4008
rect 1934 4007 1940 4008
rect 1974 4008 1980 4009
rect 1996 4008 1998 4069
rect 2284 4008 2286 4069
rect 2588 4008 2590 4069
rect 2876 4008 2878 4069
rect 3164 4008 3166 4069
rect 3452 4008 3454 4069
rect 3800 4009 3802 4069
rect 3840 4045 3842 4105
rect 3838 4044 3844 4045
rect 4940 4044 4942 4105
rect 5076 4044 5078 4105
rect 5212 4044 5214 4105
rect 5348 4044 5350 4105
rect 5484 4044 5486 4105
rect 5664 4045 5666 4105
rect 5662 4044 5668 4045
rect 3838 4040 3839 4044
rect 3843 4040 3844 4044
rect 3838 4039 3844 4040
rect 4938 4043 4944 4044
rect 4938 4039 4939 4043
rect 4943 4039 4944 4043
rect 4938 4038 4944 4039
rect 5074 4043 5080 4044
rect 5074 4039 5075 4043
rect 5079 4039 5080 4043
rect 5074 4038 5080 4039
rect 5210 4043 5216 4044
rect 5210 4039 5211 4043
rect 5215 4039 5216 4043
rect 5210 4038 5216 4039
rect 5346 4043 5352 4044
rect 5346 4039 5347 4043
rect 5351 4039 5352 4043
rect 5346 4038 5352 4039
rect 5482 4043 5488 4044
rect 5482 4039 5483 4043
rect 5487 4039 5488 4043
rect 5662 4040 5663 4044
rect 5667 4040 5668 4044
rect 5662 4039 5668 4040
rect 5482 4038 5488 4039
rect 4966 4028 4972 4029
rect 3838 4027 3844 4028
rect 3838 4023 3839 4027
rect 3843 4023 3844 4027
rect 4966 4024 4967 4028
rect 4971 4024 4972 4028
rect 4966 4023 4972 4024
rect 5102 4028 5108 4029
rect 5102 4024 5103 4028
rect 5107 4024 5108 4028
rect 5102 4023 5108 4024
rect 5238 4028 5244 4029
rect 5238 4024 5239 4028
rect 5243 4024 5244 4028
rect 5238 4023 5244 4024
rect 5374 4028 5380 4029
rect 5374 4024 5375 4028
rect 5379 4024 5380 4028
rect 5374 4023 5380 4024
rect 5510 4028 5516 4029
rect 5510 4024 5511 4028
rect 5515 4024 5516 4028
rect 5510 4023 5516 4024
rect 5662 4027 5668 4028
rect 5662 4023 5663 4027
rect 5667 4023 5668 4027
rect 3838 4022 3844 4023
rect 3798 4008 3804 4009
rect 1936 3947 1938 4007
rect 1974 4004 1975 4008
rect 1979 4004 1980 4008
rect 1974 4003 1980 4004
rect 1994 4007 2000 4008
rect 1994 4003 1995 4007
rect 1999 4003 2000 4007
rect 1994 4002 2000 4003
rect 2282 4007 2288 4008
rect 2282 4003 2283 4007
rect 2287 4003 2288 4007
rect 2282 4002 2288 4003
rect 2586 4007 2592 4008
rect 2586 4003 2587 4007
rect 2591 4003 2592 4007
rect 2586 4002 2592 4003
rect 2874 4007 2880 4008
rect 2874 4003 2875 4007
rect 2879 4003 2880 4007
rect 2874 4002 2880 4003
rect 3162 4007 3168 4008
rect 3162 4003 3163 4007
rect 3167 4003 3168 4007
rect 3162 4002 3168 4003
rect 3450 4007 3456 4008
rect 3450 4003 3451 4007
rect 3455 4003 3456 4007
rect 3798 4004 3799 4008
rect 3803 4004 3804 4008
rect 3798 4003 3804 4004
rect 3450 4002 3456 4003
rect 2022 3992 2028 3993
rect 1974 3991 1980 3992
rect 1974 3987 1975 3991
rect 1979 3987 1980 3991
rect 2022 3988 2023 3992
rect 2027 3988 2028 3992
rect 2022 3987 2028 3988
rect 2310 3992 2316 3993
rect 2310 3988 2311 3992
rect 2315 3988 2316 3992
rect 2310 3987 2316 3988
rect 2614 3992 2620 3993
rect 2614 3988 2615 3992
rect 2619 3988 2620 3992
rect 2614 3987 2620 3988
rect 2902 3992 2908 3993
rect 2902 3988 2903 3992
rect 2907 3988 2908 3992
rect 2902 3987 2908 3988
rect 3190 3992 3196 3993
rect 3190 3988 3191 3992
rect 3195 3988 3196 3992
rect 3190 3987 3196 3988
rect 3478 3992 3484 3993
rect 3478 3988 3479 3992
rect 3483 3988 3484 3992
rect 3478 3987 3484 3988
rect 3798 3991 3804 3992
rect 3840 3991 3842 4022
rect 4968 3991 4970 4023
rect 5104 3991 5106 4023
rect 5240 3991 5242 4023
rect 5376 3991 5378 4023
rect 5512 3991 5514 4023
rect 5662 4022 5668 4023
rect 5664 3991 5666 4022
rect 3798 3987 3799 3991
rect 3803 3987 3804 3991
rect 1974 3986 1980 3987
rect 111 3946 115 3947
rect 111 3941 115 3942
rect 203 3946 207 3947
rect 203 3941 207 3942
rect 251 3946 255 3947
rect 251 3941 255 3942
rect 395 3946 399 3947
rect 395 3941 399 3942
rect 451 3946 455 3947
rect 451 3941 455 3942
rect 587 3946 591 3947
rect 587 3941 591 3942
rect 643 3946 647 3947
rect 643 3941 647 3942
rect 779 3946 783 3947
rect 779 3941 783 3942
rect 827 3946 831 3947
rect 827 3941 831 3942
rect 963 3946 967 3947
rect 963 3941 967 3942
rect 1003 3946 1007 3947
rect 1003 3941 1007 3942
rect 1139 3946 1143 3947
rect 1139 3941 1143 3942
rect 1171 3946 1175 3947
rect 1171 3941 1175 3942
rect 1307 3946 1311 3947
rect 1307 3941 1311 3942
rect 1331 3946 1335 3947
rect 1331 3941 1335 3942
rect 1475 3946 1479 3947
rect 1475 3941 1479 3942
rect 1491 3946 1495 3947
rect 1491 3941 1495 3942
rect 1643 3946 1647 3947
rect 1643 3941 1647 3942
rect 1651 3946 1655 3947
rect 1651 3941 1655 3942
rect 1787 3946 1791 3947
rect 1787 3941 1791 3942
rect 1935 3946 1939 3947
rect 1976 3943 1978 3986
rect 2024 3943 2026 3987
rect 2312 3943 2314 3987
rect 2616 3943 2618 3987
rect 2904 3943 2906 3987
rect 3192 3943 3194 3987
rect 3480 3943 3482 3987
rect 3798 3986 3804 3987
rect 3839 3990 3843 3991
rect 3800 3943 3802 3986
rect 3839 3985 3843 3986
rect 4831 3990 4835 3991
rect 4831 3985 4835 3986
rect 4967 3990 4971 3991
rect 4967 3985 4971 3986
rect 5103 3990 5107 3991
rect 5103 3985 5107 3986
rect 5111 3990 5115 3991
rect 5111 3985 5115 3986
rect 5239 3990 5243 3991
rect 5239 3985 5243 3986
rect 5255 3990 5259 3991
rect 5255 3985 5259 3986
rect 5375 3990 5379 3991
rect 5375 3985 5379 3986
rect 5407 3990 5411 3991
rect 5407 3985 5411 3986
rect 5511 3990 5515 3991
rect 5511 3985 5515 3986
rect 5543 3990 5547 3991
rect 5543 3985 5547 3986
rect 5663 3990 5667 3991
rect 5663 3985 5667 3986
rect 3840 3962 3842 3985
rect 3838 3961 3844 3962
rect 4832 3961 4834 3985
rect 4968 3961 4970 3985
rect 5112 3961 5114 3985
rect 5256 3961 5258 3985
rect 5408 3961 5410 3985
rect 5544 3961 5546 3985
rect 5664 3962 5666 3985
rect 5662 3961 5668 3962
rect 3838 3957 3839 3961
rect 3843 3957 3844 3961
rect 3838 3956 3844 3957
rect 4830 3960 4836 3961
rect 4830 3956 4831 3960
rect 4835 3956 4836 3960
rect 4830 3955 4836 3956
rect 4966 3960 4972 3961
rect 4966 3956 4967 3960
rect 4971 3956 4972 3960
rect 4966 3955 4972 3956
rect 5110 3960 5116 3961
rect 5110 3956 5111 3960
rect 5115 3956 5116 3960
rect 5110 3955 5116 3956
rect 5254 3960 5260 3961
rect 5254 3956 5255 3960
rect 5259 3956 5260 3960
rect 5254 3955 5260 3956
rect 5406 3960 5412 3961
rect 5406 3956 5407 3960
rect 5411 3956 5412 3960
rect 5406 3955 5412 3956
rect 5542 3960 5548 3961
rect 5542 3956 5543 3960
rect 5547 3956 5548 3960
rect 5662 3957 5663 3961
rect 5667 3957 5668 3961
rect 5662 3956 5668 3957
rect 5542 3955 5548 3956
rect 4802 3945 4808 3946
rect 3838 3944 3844 3945
rect 1935 3941 1939 3942
rect 1975 3942 1979 3943
rect 112 3881 114 3941
rect 110 3880 116 3881
rect 252 3880 254 3941
rect 452 3880 454 3941
rect 644 3880 646 3941
rect 828 3880 830 3941
rect 1004 3880 1006 3941
rect 1172 3880 1174 3941
rect 1332 3880 1334 3941
rect 1492 3880 1494 3941
rect 1652 3880 1654 3941
rect 1788 3880 1790 3941
rect 1936 3881 1938 3941
rect 1975 3937 1979 3938
rect 2023 3942 2027 3943
rect 2023 3937 2027 3938
rect 2311 3942 2315 3943
rect 2311 3937 2315 3938
rect 2615 3942 2619 3943
rect 2615 3937 2619 3938
rect 2671 3942 2675 3943
rect 2671 3937 2675 3938
rect 2807 3942 2811 3943
rect 2807 3937 2811 3938
rect 2903 3942 2907 3943
rect 2903 3937 2907 3938
rect 2943 3942 2947 3943
rect 2943 3937 2947 3938
rect 3079 3942 3083 3943
rect 3079 3937 3083 3938
rect 3191 3942 3195 3943
rect 3191 3937 3195 3938
rect 3215 3942 3219 3943
rect 3215 3937 3219 3938
rect 3479 3942 3483 3943
rect 3479 3937 3483 3938
rect 3799 3942 3803 3943
rect 3838 3940 3839 3944
rect 3843 3940 3844 3944
rect 4802 3941 4803 3945
rect 4807 3941 4808 3945
rect 4802 3940 4808 3941
rect 4938 3945 4944 3946
rect 4938 3941 4939 3945
rect 4943 3941 4944 3945
rect 4938 3940 4944 3941
rect 5082 3945 5088 3946
rect 5082 3941 5083 3945
rect 5087 3941 5088 3945
rect 5082 3940 5088 3941
rect 5226 3945 5232 3946
rect 5226 3941 5227 3945
rect 5231 3941 5232 3945
rect 5226 3940 5232 3941
rect 5378 3945 5384 3946
rect 5378 3941 5379 3945
rect 5383 3941 5384 3945
rect 5378 3940 5384 3941
rect 5514 3945 5520 3946
rect 5514 3941 5515 3945
rect 5519 3941 5520 3945
rect 5514 3940 5520 3941
rect 5662 3944 5668 3945
rect 5662 3940 5663 3944
rect 5667 3940 5668 3944
rect 3838 3939 3844 3940
rect 3799 3937 3803 3938
rect 1976 3914 1978 3937
rect 1974 3913 1980 3914
rect 2672 3913 2674 3937
rect 2808 3913 2810 3937
rect 2944 3913 2946 3937
rect 3080 3913 3082 3937
rect 3216 3913 3218 3937
rect 3800 3914 3802 3937
rect 3798 3913 3804 3914
rect 1974 3909 1975 3913
rect 1979 3909 1980 3913
rect 1974 3908 1980 3909
rect 2670 3912 2676 3913
rect 2670 3908 2671 3912
rect 2675 3908 2676 3912
rect 2670 3907 2676 3908
rect 2806 3912 2812 3913
rect 2806 3908 2807 3912
rect 2811 3908 2812 3912
rect 2806 3907 2812 3908
rect 2942 3912 2948 3913
rect 2942 3908 2943 3912
rect 2947 3908 2948 3912
rect 2942 3907 2948 3908
rect 3078 3912 3084 3913
rect 3078 3908 3079 3912
rect 3083 3908 3084 3912
rect 3078 3907 3084 3908
rect 3214 3912 3220 3913
rect 3214 3908 3215 3912
rect 3219 3908 3220 3912
rect 3798 3909 3799 3913
rect 3803 3909 3804 3913
rect 3798 3908 3804 3909
rect 3214 3907 3220 3908
rect 2642 3897 2648 3898
rect 1974 3896 1980 3897
rect 1974 3892 1975 3896
rect 1979 3892 1980 3896
rect 2642 3893 2643 3897
rect 2647 3893 2648 3897
rect 2642 3892 2648 3893
rect 2778 3897 2784 3898
rect 2778 3893 2779 3897
rect 2783 3893 2784 3897
rect 2778 3892 2784 3893
rect 2914 3897 2920 3898
rect 2914 3893 2915 3897
rect 2919 3893 2920 3897
rect 2914 3892 2920 3893
rect 3050 3897 3056 3898
rect 3050 3893 3051 3897
rect 3055 3893 3056 3897
rect 3050 3892 3056 3893
rect 3186 3897 3192 3898
rect 3186 3893 3187 3897
rect 3191 3893 3192 3897
rect 3186 3892 3192 3893
rect 3798 3896 3804 3897
rect 3798 3892 3799 3896
rect 3803 3892 3804 3896
rect 1974 3891 1980 3892
rect 1934 3880 1940 3881
rect 110 3876 111 3880
rect 115 3876 116 3880
rect 110 3875 116 3876
rect 250 3879 256 3880
rect 250 3875 251 3879
rect 255 3875 256 3879
rect 250 3874 256 3875
rect 450 3879 456 3880
rect 450 3875 451 3879
rect 455 3875 456 3879
rect 450 3874 456 3875
rect 642 3879 648 3880
rect 642 3875 643 3879
rect 647 3875 648 3879
rect 642 3874 648 3875
rect 826 3879 832 3880
rect 826 3875 827 3879
rect 831 3875 832 3879
rect 826 3874 832 3875
rect 1002 3879 1008 3880
rect 1002 3875 1003 3879
rect 1007 3875 1008 3879
rect 1002 3874 1008 3875
rect 1170 3879 1176 3880
rect 1170 3875 1171 3879
rect 1175 3875 1176 3879
rect 1170 3874 1176 3875
rect 1330 3879 1336 3880
rect 1330 3875 1331 3879
rect 1335 3875 1336 3879
rect 1330 3874 1336 3875
rect 1490 3879 1496 3880
rect 1490 3875 1491 3879
rect 1495 3875 1496 3879
rect 1490 3874 1496 3875
rect 1650 3879 1656 3880
rect 1650 3875 1651 3879
rect 1655 3875 1656 3879
rect 1650 3874 1656 3875
rect 1786 3879 1792 3880
rect 1786 3875 1787 3879
rect 1791 3875 1792 3879
rect 1934 3876 1935 3880
rect 1939 3876 1940 3880
rect 1934 3875 1940 3876
rect 1786 3874 1792 3875
rect 278 3864 284 3865
rect 110 3863 116 3864
rect 110 3859 111 3863
rect 115 3859 116 3863
rect 278 3860 279 3864
rect 283 3860 284 3864
rect 278 3859 284 3860
rect 478 3864 484 3865
rect 478 3860 479 3864
rect 483 3860 484 3864
rect 478 3859 484 3860
rect 670 3864 676 3865
rect 670 3860 671 3864
rect 675 3860 676 3864
rect 670 3859 676 3860
rect 854 3864 860 3865
rect 854 3860 855 3864
rect 859 3860 860 3864
rect 854 3859 860 3860
rect 1030 3864 1036 3865
rect 1030 3860 1031 3864
rect 1035 3860 1036 3864
rect 1030 3859 1036 3860
rect 1198 3864 1204 3865
rect 1198 3860 1199 3864
rect 1203 3860 1204 3864
rect 1198 3859 1204 3860
rect 1358 3864 1364 3865
rect 1358 3860 1359 3864
rect 1363 3860 1364 3864
rect 1358 3859 1364 3860
rect 1518 3864 1524 3865
rect 1518 3860 1519 3864
rect 1523 3860 1524 3864
rect 1518 3859 1524 3860
rect 1678 3864 1684 3865
rect 1678 3860 1679 3864
rect 1683 3860 1684 3864
rect 1678 3859 1684 3860
rect 1814 3864 1820 3865
rect 1814 3860 1815 3864
rect 1819 3860 1820 3864
rect 1814 3859 1820 3860
rect 1934 3863 1940 3864
rect 1934 3859 1935 3863
rect 1939 3859 1940 3863
rect 110 3858 116 3859
rect 112 3835 114 3858
rect 280 3835 282 3859
rect 480 3835 482 3859
rect 672 3835 674 3859
rect 856 3835 858 3859
rect 1032 3835 1034 3859
rect 1200 3835 1202 3859
rect 1360 3835 1362 3859
rect 1520 3835 1522 3859
rect 1680 3835 1682 3859
rect 1816 3835 1818 3859
rect 1934 3858 1940 3859
rect 1936 3835 1938 3858
rect 111 3834 115 3835
rect 111 3829 115 3830
rect 279 3834 283 3835
rect 279 3829 283 3830
rect 311 3834 315 3835
rect 311 3829 315 3830
rect 479 3834 483 3835
rect 479 3829 483 3830
rect 511 3834 515 3835
rect 511 3829 515 3830
rect 671 3834 675 3835
rect 671 3829 675 3830
rect 735 3834 739 3835
rect 735 3829 739 3830
rect 855 3834 859 3835
rect 855 3829 859 3830
rect 991 3834 995 3835
rect 991 3829 995 3830
rect 1031 3834 1035 3835
rect 1031 3829 1035 3830
rect 1199 3834 1203 3835
rect 1199 3829 1203 3830
rect 1263 3834 1267 3835
rect 1263 3829 1267 3830
rect 1359 3834 1363 3835
rect 1359 3829 1363 3830
rect 1519 3834 1523 3835
rect 1519 3829 1523 3830
rect 1551 3834 1555 3835
rect 1551 3829 1555 3830
rect 1679 3834 1683 3835
rect 1679 3829 1683 3830
rect 1815 3834 1819 3835
rect 1815 3829 1819 3830
rect 1935 3834 1939 3835
rect 1935 3829 1939 3830
rect 112 3806 114 3829
rect 110 3805 116 3806
rect 312 3805 314 3829
rect 512 3805 514 3829
rect 736 3805 738 3829
rect 992 3805 994 3829
rect 1264 3805 1266 3829
rect 1552 3805 1554 3829
rect 1816 3805 1818 3829
rect 1936 3806 1938 3829
rect 1976 3819 1978 3891
rect 2644 3819 2646 3892
rect 2780 3819 2782 3892
rect 2916 3819 2918 3892
rect 3052 3819 3054 3892
rect 3188 3819 3190 3892
rect 3798 3891 3804 3892
rect 3800 3819 3802 3891
rect 3840 3859 3842 3939
rect 4804 3859 4806 3940
rect 4940 3859 4942 3940
rect 5084 3859 5086 3940
rect 5228 3859 5230 3940
rect 5380 3859 5382 3940
rect 5516 3859 5518 3940
rect 5662 3939 5668 3940
rect 5664 3859 5666 3939
rect 3839 3858 3843 3859
rect 3839 3853 3843 3854
rect 4499 3858 4503 3859
rect 4499 3853 4503 3854
rect 4675 3858 4679 3859
rect 4675 3853 4679 3854
rect 4803 3858 4807 3859
rect 4803 3853 4807 3854
rect 4875 3858 4879 3859
rect 4875 3853 4879 3854
rect 4939 3858 4943 3859
rect 4939 3853 4943 3854
rect 5083 3858 5087 3859
rect 5083 3853 5087 3854
rect 5091 3858 5095 3859
rect 5091 3853 5095 3854
rect 5227 3858 5231 3859
rect 5227 3853 5231 3854
rect 5315 3858 5319 3859
rect 5315 3853 5319 3854
rect 5379 3858 5383 3859
rect 5379 3853 5383 3854
rect 5515 3858 5519 3859
rect 5515 3853 5519 3854
rect 5663 3858 5667 3859
rect 5663 3853 5667 3854
rect 1975 3818 1979 3819
rect 1975 3813 1979 3814
rect 1995 3818 1999 3819
rect 1995 3813 1999 3814
rect 2131 3818 2135 3819
rect 2131 3813 2135 3814
rect 2283 3818 2287 3819
rect 2283 3813 2287 3814
rect 2443 3818 2447 3819
rect 2443 3813 2447 3814
rect 2603 3818 2607 3819
rect 2603 3813 2607 3814
rect 2643 3818 2647 3819
rect 2643 3813 2647 3814
rect 2763 3818 2767 3819
rect 2763 3813 2767 3814
rect 2779 3818 2783 3819
rect 2779 3813 2783 3814
rect 2915 3818 2919 3819
rect 2915 3813 2919 3814
rect 2923 3818 2927 3819
rect 2923 3813 2927 3814
rect 3051 3818 3055 3819
rect 3051 3813 3055 3814
rect 3083 3818 3087 3819
rect 3083 3813 3087 3814
rect 3187 3818 3191 3819
rect 3187 3813 3191 3814
rect 3243 3818 3247 3819
rect 3243 3813 3247 3814
rect 3411 3818 3415 3819
rect 3411 3813 3415 3814
rect 3799 3818 3803 3819
rect 3799 3813 3803 3814
rect 1934 3805 1940 3806
rect 110 3801 111 3805
rect 115 3801 116 3805
rect 110 3800 116 3801
rect 310 3804 316 3805
rect 310 3800 311 3804
rect 315 3800 316 3804
rect 310 3799 316 3800
rect 510 3804 516 3805
rect 510 3800 511 3804
rect 515 3800 516 3804
rect 510 3799 516 3800
rect 734 3804 740 3805
rect 734 3800 735 3804
rect 739 3800 740 3804
rect 734 3799 740 3800
rect 990 3804 996 3805
rect 990 3800 991 3804
rect 995 3800 996 3804
rect 990 3799 996 3800
rect 1262 3804 1268 3805
rect 1262 3800 1263 3804
rect 1267 3800 1268 3804
rect 1262 3799 1268 3800
rect 1550 3804 1556 3805
rect 1550 3800 1551 3804
rect 1555 3800 1556 3804
rect 1550 3799 1556 3800
rect 1814 3804 1820 3805
rect 1814 3800 1815 3804
rect 1819 3800 1820 3804
rect 1934 3801 1935 3805
rect 1939 3801 1940 3805
rect 1934 3800 1940 3801
rect 1814 3799 1820 3800
rect 282 3789 288 3790
rect 110 3788 116 3789
rect 110 3784 111 3788
rect 115 3784 116 3788
rect 282 3785 283 3789
rect 287 3785 288 3789
rect 282 3784 288 3785
rect 482 3789 488 3790
rect 482 3785 483 3789
rect 487 3785 488 3789
rect 482 3784 488 3785
rect 706 3789 712 3790
rect 706 3785 707 3789
rect 711 3785 712 3789
rect 706 3784 712 3785
rect 962 3789 968 3790
rect 962 3785 963 3789
rect 967 3785 968 3789
rect 962 3784 968 3785
rect 1234 3789 1240 3790
rect 1234 3785 1235 3789
rect 1239 3785 1240 3789
rect 1234 3784 1240 3785
rect 1522 3789 1528 3790
rect 1522 3785 1523 3789
rect 1527 3785 1528 3789
rect 1522 3784 1528 3785
rect 1786 3789 1792 3790
rect 1786 3785 1787 3789
rect 1791 3785 1792 3789
rect 1786 3784 1792 3785
rect 1934 3788 1940 3789
rect 1934 3784 1935 3788
rect 1939 3784 1940 3788
rect 110 3783 116 3784
rect 112 3699 114 3783
rect 284 3699 286 3784
rect 484 3699 486 3784
rect 708 3699 710 3784
rect 964 3699 966 3784
rect 1236 3699 1238 3784
rect 1524 3699 1526 3784
rect 1788 3699 1790 3784
rect 1934 3783 1940 3784
rect 1936 3699 1938 3783
rect 1976 3753 1978 3813
rect 1974 3752 1980 3753
rect 1996 3752 1998 3813
rect 2132 3752 2134 3813
rect 2284 3752 2286 3813
rect 2444 3752 2446 3813
rect 2604 3752 2606 3813
rect 2764 3752 2766 3813
rect 2924 3752 2926 3813
rect 3084 3752 3086 3813
rect 3244 3752 3246 3813
rect 3412 3752 3414 3813
rect 3800 3753 3802 3813
rect 3840 3793 3842 3853
rect 3838 3792 3844 3793
rect 4500 3792 4502 3853
rect 4676 3792 4678 3853
rect 4876 3792 4878 3853
rect 5092 3792 5094 3853
rect 5316 3792 5318 3853
rect 5516 3792 5518 3853
rect 5664 3793 5666 3853
rect 5662 3792 5668 3793
rect 3838 3788 3839 3792
rect 3843 3788 3844 3792
rect 3838 3787 3844 3788
rect 4498 3791 4504 3792
rect 4498 3787 4499 3791
rect 4503 3787 4504 3791
rect 4498 3786 4504 3787
rect 4674 3791 4680 3792
rect 4674 3787 4675 3791
rect 4679 3787 4680 3791
rect 4674 3786 4680 3787
rect 4874 3791 4880 3792
rect 4874 3787 4875 3791
rect 4879 3787 4880 3791
rect 4874 3786 4880 3787
rect 5090 3791 5096 3792
rect 5090 3787 5091 3791
rect 5095 3787 5096 3791
rect 5090 3786 5096 3787
rect 5314 3791 5320 3792
rect 5314 3787 5315 3791
rect 5319 3787 5320 3791
rect 5314 3786 5320 3787
rect 5514 3791 5520 3792
rect 5514 3787 5515 3791
rect 5519 3787 5520 3791
rect 5662 3788 5663 3792
rect 5667 3788 5668 3792
rect 5662 3787 5668 3788
rect 5514 3786 5520 3787
rect 4526 3776 4532 3777
rect 3838 3775 3844 3776
rect 3838 3771 3839 3775
rect 3843 3771 3844 3775
rect 4526 3772 4527 3776
rect 4531 3772 4532 3776
rect 4526 3771 4532 3772
rect 4702 3776 4708 3777
rect 4702 3772 4703 3776
rect 4707 3772 4708 3776
rect 4702 3771 4708 3772
rect 4902 3776 4908 3777
rect 4902 3772 4903 3776
rect 4907 3772 4908 3776
rect 4902 3771 4908 3772
rect 5118 3776 5124 3777
rect 5118 3772 5119 3776
rect 5123 3772 5124 3776
rect 5118 3771 5124 3772
rect 5342 3776 5348 3777
rect 5342 3772 5343 3776
rect 5347 3772 5348 3776
rect 5342 3771 5348 3772
rect 5542 3776 5548 3777
rect 5542 3772 5543 3776
rect 5547 3772 5548 3776
rect 5542 3771 5548 3772
rect 5662 3775 5668 3776
rect 5662 3771 5663 3775
rect 5667 3771 5668 3775
rect 3838 3770 3844 3771
rect 3798 3752 3804 3753
rect 1974 3748 1975 3752
rect 1979 3748 1980 3752
rect 1974 3747 1980 3748
rect 1994 3751 2000 3752
rect 1994 3747 1995 3751
rect 1999 3747 2000 3751
rect 1994 3746 2000 3747
rect 2130 3751 2136 3752
rect 2130 3747 2131 3751
rect 2135 3747 2136 3751
rect 2130 3746 2136 3747
rect 2282 3751 2288 3752
rect 2282 3747 2283 3751
rect 2287 3747 2288 3751
rect 2282 3746 2288 3747
rect 2442 3751 2448 3752
rect 2442 3747 2443 3751
rect 2447 3747 2448 3751
rect 2442 3746 2448 3747
rect 2602 3751 2608 3752
rect 2602 3747 2603 3751
rect 2607 3747 2608 3751
rect 2602 3746 2608 3747
rect 2762 3751 2768 3752
rect 2762 3747 2763 3751
rect 2767 3747 2768 3751
rect 2762 3746 2768 3747
rect 2922 3751 2928 3752
rect 2922 3747 2923 3751
rect 2927 3747 2928 3751
rect 2922 3746 2928 3747
rect 3082 3751 3088 3752
rect 3082 3747 3083 3751
rect 3087 3747 3088 3751
rect 3082 3746 3088 3747
rect 3242 3751 3248 3752
rect 3242 3747 3243 3751
rect 3247 3747 3248 3751
rect 3242 3746 3248 3747
rect 3410 3751 3416 3752
rect 3410 3747 3411 3751
rect 3415 3747 3416 3751
rect 3798 3748 3799 3752
rect 3803 3748 3804 3752
rect 3798 3747 3804 3748
rect 3410 3746 3416 3747
rect 2022 3736 2028 3737
rect 1974 3735 1980 3736
rect 1974 3731 1975 3735
rect 1979 3731 1980 3735
rect 2022 3732 2023 3736
rect 2027 3732 2028 3736
rect 2022 3731 2028 3732
rect 2158 3736 2164 3737
rect 2158 3732 2159 3736
rect 2163 3732 2164 3736
rect 2158 3731 2164 3732
rect 2310 3736 2316 3737
rect 2310 3732 2311 3736
rect 2315 3732 2316 3736
rect 2310 3731 2316 3732
rect 2470 3736 2476 3737
rect 2470 3732 2471 3736
rect 2475 3732 2476 3736
rect 2470 3731 2476 3732
rect 2630 3736 2636 3737
rect 2630 3732 2631 3736
rect 2635 3732 2636 3736
rect 2630 3731 2636 3732
rect 2790 3736 2796 3737
rect 2790 3732 2791 3736
rect 2795 3732 2796 3736
rect 2790 3731 2796 3732
rect 2950 3736 2956 3737
rect 2950 3732 2951 3736
rect 2955 3732 2956 3736
rect 2950 3731 2956 3732
rect 3110 3736 3116 3737
rect 3110 3732 3111 3736
rect 3115 3732 3116 3736
rect 3110 3731 3116 3732
rect 3270 3736 3276 3737
rect 3270 3732 3271 3736
rect 3275 3732 3276 3736
rect 3270 3731 3276 3732
rect 3438 3736 3444 3737
rect 3438 3732 3439 3736
rect 3443 3732 3444 3736
rect 3438 3731 3444 3732
rect 3798 3735 3804 3736
rect 3798 3731 3799 3735
rect 3803 3731 3804 3735
rect 1974 3730 1980 3731
rect 1976 3699 1978 3730
rect 2024 3699 2026 3731
rect 2160 3699 2162 3731
rect 2312 3699 2314 3731
rect 2472 3699 2474 3731
rect 2632 3699 2634 3731
rect 2792 3699 2794 3731
rect 2952 3699 2954 3731
rect 3112 3699 3114 3731
rect 3272 3699 3274 3731
rect 3440 3699 3442 3731
rect 3798 3730 3804 3731
rect 3800 3699 3802 3730
rect 3840 3723 3842 3770
rect 4528 3723 4530 3771
rect 4704 3723 4706 3771
rect 4904 3723 4906 3771
rect 5120 3723 5122 3771
rect 5344 3723 5346 3771
rect 5544 3723 5546 3771
rect 5662 3770 5668 3771
rect 5664 3723 5666 3770
rect 3839 3722 3843 3723
rect 3839 3717 3843 3718
rect 4271 3722 4275 3723
rect 4271 3717 4275 3718
rect 4471 3722 4475 3723
rect 4471 3717 4475 3718
rect 4527 3722 4531 3723
rect 4527 3717 4531 3718
rect 4695 3722 4699 3723
rect 4695 3717 4699 3718
rect 4703 3722 4707 3723
rect 4703 3717 4707 3718
rect 4903 3722 4907 3723
rect 4903 3717 4907 3718
rect 4935 3722 4939 3723
rect 4935 3717 4939 3718
rect 5119 3722 5123 3723
rect 5119 3717 5123 3718
rect 5191 3722 5195 3723
rect 5191 3717 5195 3718
rect 5343 3722 5347 3723
rect 5343 3717 5347 3718
rect 5447 3722 5451 3723
rect 5447 3717 5451 3718
rect 5543 3722 5547 3723
rect 5543 3717 5547 3718
rect 5663 3722 5667 3723
rect 5663 3717 5667 3718
rect 111 3698 115 3699
rect 111 3693 115 3694
rect 155 3698 159 3699
rect 155 3693 159 3694
rect 283 3698 287 3699
rect 283 3693 287 3694
rect 291 3698 295 3699
rect 291 3693 295 3694
rect 427 3698 431 3699
rect 427 3693 431 3694
rect 483 3698 487 3699
rect 483 3693 487 3694
rect 563 3698 567 3699
rect 563 3693 567 3694
rect 699 3698 703 3699
rect 699 3693 703 3694
rect 707 3698 711 3699
rect 707 3693 711 3694
rect 835 3698 839 3699
rect 835 3693 839 3694
rect 963 3698 967 3699
rect 963 3693 967 3694
rect 971 3698 975 3699
rect 971 3693 975 3694
rect 1107 3698 1111 3699
rect 1107 3693 1111 3694
rect 1235 3698 1239 3699
rect 1235 3693 1239 3694
rect 1243 3698 1247 3699
rect 1243 3693 1247 3694
rect 1379 3698 1383 3699
rect 1379 3693 1383 3694
rect 1515 3698 1519 3699
rect 1515 3693 1519 3694
rect 1523 3698 1527 3699
rect 1523 3693 1527 3694
rect 1787 3698 1791 3699
rect 1787 3693 1791 3694
rect 1935 3698 1939 3699
rect 1935 3693 1939 3694
rect 1975 3698 1979 3699
rect 1975 3693 1979 3694
rect 2023 3698 2027 3699
rect 2023 3693 2027 3694
rect 2047 3698 2051 3699
rect 2047 3693 2051 3694
rect 2159 3698 2163 3699
rect 2159 3693 2163 3694
rect 2223 3698 2227 3699
rect 2223 3693 2227 3694
rect 2311 3698 2315 3699
rect 2311 3693 2315 3694
rect 2407 3698 2411 3699
rect 2407 3693 2411 3694
rect 2471 3698 2475 3699
rect 2471 3693 2475 3694
rect 2591 3698 2595 3699
rect 2591 3693 2595 3694
rect 2631 3698 2635 3699
rect 2631 3693 2635 3694
rect 2783 3698 2787 3699
rect 2783 3693 2787 3694
rect 2791 3698 2795 3699
rect 2791 3693 2795 3694
rect 2951 3698 2955 3699
rect 2951 3693 2955 3694
rect 2967 3698 2971 3699
rect 2967 3693 2971 3694
rect 3111 3698 3115 3699
rect 3111 3693 3115 3694
rect 3151 3698 3155 3699
rect 3151 3693 3155 3694
rect 3271 3698 3275 3699
rect 3271 3693 3275 3694
rect 3335 3698 3339 3699
rect 3335 3693 3339 3694
rect 3439 3698 3443 3699
rect 3439 3693 3443 3694
rect 3519 3698 3523 3699
rect 3519 3693 3523 3694
rect 3679 3698 3683 3699
rect 3679 3693 3683 3694
rect 3799 3698 3803 3699
rect 3840 3694 3842 3717
rect 3799 3693 3803 3694
rect 3838 3693 3844 3694
rect 4272 3693 4274 3717
rect 4472 3693 4474 3717
rect 4696 3693 4698 3717
rect 4936 3693 4938 3717
rect 5192 3693 5194 3717
rect 5448 3693 5450 3717
rect 5664 3694 5666 3717
rect 5662 3693 5668 3694
rect 112 3633 114 3693
rect 110 3632 116 3633
rect 156 3632 158 3693
rect 292 3632 294 3693
rect 428 3632 430 3693
rect 564 3632 566 3693
rect 700 3632 702 3693
rect 836 3632 838 3693
rect 972 3632 974 3693
rect 1108 3632 1110 3693
rect 1244 3632 1246 3693
rect 1380 3632 1382 3693
rect 1516 3632 1518 3693
rect 1936 3633 1938 3693
rect 1976 3670 1978 3693
rect 1974 3669 1980 3670
rect 2048 3669 2050 3693
rect 2224 3669 2226 3693
rect 2408 3669 2410 3693
rect 2592 3669 2594 3693
rect 2784 3669 2786 3693
rect 2968 3669 2970 3693
rect 3152 3669 3154 3693
rect 3336 3669 3338 3693
rect 3520 3669 3522 3693
rect 3680 3669 3682 3693
rect 3800 3670 3802 3693
rect 3838 3689 3839 3693
rect 3843 3689 3844 3693
rect 3838 3688 3844 3689
rect 4270 3692 4276 3693
rect 4270 3688 4271 3692
rect 4275 3688 4276 3692
rect 4270 3687 4276 3688
rect 4470 3692 4476 3693
rect 4470 3688 4471 3692
rect 4475 3688 4476 3692
rect 4470 3687 4476 3688
rect 4694 3692 4700 3693
rect 4694 3688 4695 3692
rect 4699 3688 4700 3692
rect 4694 3687 4700 3688
rect 4934 3692 4940 3693
rect 4934 3688 4935 3692
rect 4939 3688 4940 3692
rect 4934 3687 4940 3688
rect 5190 3692 5196 3693
rect 5190 3688 5191 3692
rect 5195 3688 5196 3692
rect 5190 3687 5196 3688
rect 5446 3692 5452 3693
rect 5446 3688 5447 3692
rect 5451 3688 5452 3692
rect 5662 3689 5663 3693
rect 5667 3689 5668 3693
rect 5662 3688 5668 3689
rect 5446 3687 5452 3688
rect 4242 3677 4248 3678
rect 3838 3676 3844 3677
rect 3838 3672 3839 3676
rect 3843 3672 3844 3676
rect 4242 3673 4243 3677
rect 4247 3673 4248 3677
rect 4242 3672 4248 3673
rect 4442 3677 4448 3678
rect 4442 3673 4443 3677
rect 4447 3673 4448 3677
rect 4442 3672 4448 3673
rect 4666 3677 4672 3678
rect 4666 3673 4667 3677
rect 4671 3673 4672 3677
rect 4666 3672 4672 3673
rect 4906 3677 4912 3678
rect 4906 3673 4907 3677
rect 4911 3673 4912 3677
rect 4906 3672 4912 3673
rect 5162 3677 5168 3678
rect 5162 3673 5163 3677
rect 5167 3673 5168 3677
rect 5162 3672 5168 3673
rect 5418 3677 5424 3678
rect 5418 3673 5419 3677
rect 5423 3673 5424 3677
rect 5418 3672 5424 3673
rect 5662 3676 5668 3677
rect 5662 3672 5663 3676
rect 5667 3672 5668 3676
rect 3838 3671 3844 3672
rect 3798 3669 3804 3670
rect 1974 3665 1975 3669
rect 1979 3665 1980 3669
rect 1974 3664 1980 3665
rect 2046 3668 2052 3669
rect 2046 3664 2047 3668
rect 2051 3664 2052 3668
rect 2046 3663 2052 3664
rect 2222 3668 2228 3669
rect 2222 3664 2223 3668
rect 2227 3664 2228 3668
rect 2222 3663 2228 3664
rect 2406 3668 2412 3669
rect 2406 3664 2407 3668
rect 2411 3664 2412 3668
rect 2406 3663 2412 3664
rect 2590 3668 2596 3669
rect 2590 3664 2591 3668
rect 2595 3664 2596 3668
rect 2590 3663 2596 3664
rect 2782 3668 2788 3669
rect 2782 3664 2783 3668
rect 2787 3664 2788 3668
rect 2782 3663 2788 3664
rect 2966 3668 2972 3669
rect 2966 3664 2967 3668
rect 2971 3664 2972 3668
rect 2966 3663 2972 3664
rect 3150 3668 3156 3669
rect 3150 3664 3151 3668
rect 3155 3664 3156 3668
rect 3150 3663 3156 3664
rect 3334 3668 3340 3669
rect 3334 3664 3335 3668
rect 3339 3664 3340 3668
rect 3334 3663 3340 3664
rect 3518 3668 3524 3669
rect 3518 3664 3519 3668
rect 3523 3664 3524 3668
rect 3518 3663 3524 3664
rect 3678 3668 3684 3669
rect 3678 3664 3679 3668
rect 3683 3664 3684 3668
rect 3798 3665 3799 3669
rect 3803 3665 3804 3669
rect 3798 3664 3804 3665
rect 3678 3663 3684 3664
rect 2018 3653 2024 3654
rect 1974 3652 1980 3653
rect 1974 3648 1975 3652
rect 1979 3648 1980 3652
rect 2018 3649 2019 3653
rect 2023 3649 2024 3653
rect 2018 3648 2024 3649
rect 2194 3653 2200 3654
rect 2194 3649 2195 3653
rect 2199 3649 2200 3653
rect 2194 3648 2200 3649
rect 2378 3653 2384 3654
rect 2378 3649 2379 3653
rect 2383 3649 2384 3653
rect 2378 3648 2384 3649
rect 2562 3653 2568 3654
rect 2562 3649 2563 3653
rect 2567 3649 2568 3653
rect 2562 3648 2568 3649
rect 2754 3653 2760 3654
rect 2754 3649 2755 3653
rect 2759 3649 2760 3653
rect 2754 3648 2760 3649
rect 2938 3653 2944 3654
rect 2938 3649 2939 3653
rect 2943 3649 2944 3653
rect 2938 3648 2944 3649
rect 3122 3653 3128 3654
rect 3122 3649 3123 3653
rect 3127 3649 3128 3653
rect 3122 3648 3128 3649
rect 3306 3653 3312 3654
rect 3306 3649 3307 3653
rect 3311 3649 3312 3653
rect 3306 3648 3312 3649
rect 3490 3653 3496 3654
rect 3490 3649 3491 3653
rect 3495 3649 3496 3653
rect 3490 3648 3496 3649
rect 3650 3653 3656 3654
rect 3650 3649 3651 3653
rect 3655 3649 3656 3653
rect 3650 3648 3656 3649
rect 3798 3652 3804 3653
rect 3798 3648 3799 3652
rect 3803 3648 3804 3652
rect 1974 3647 1980 3648
rect 1934 3632 1940 3633
rect 110 3628 111 3632
rect 115 3628 116 3632
rect 110 3627 116 3628
rect 154 3631 160 3632
rect 154 3627 155 3631
rect 159 3627 160 3631
rect 154 3626 160 3627
rect 290 3631 296 3632
rect 290 3627 291 3631
rect 295 3627 296 3631
rect 290 3626 296 3627
rect 426 3631 432 3632
rect 426 3627 427 3631
rect 431 3627 432 3631
rect 426 3626 432 3627
rect 562 3631 568 3632
rect 562 3627 563 3631
rect 567 3627 568 3631
rect 562 3626 568 3627
rect 698 3631 704 3632
rect 698 3627 699 3631
rect 703 3627 704 3631
rect 698 3626 704 3627
rect 834 3631 840 3632
rect 834 3627 835 3631
rect 839 3627 840 3631
rect 834 3626 840 3627
rect 970 3631 976 3632
rect 970 3627 971 3631
rect 975 3627 976 3631
rect 970 3626 976 3627
rect 1106 3631 1112 3632
rect 1106 3627 1107 3631
rect 1111 3627 1112 3631
rect 1106 3626 1112 3627
rect 1242 3631 1248 3632
rect 1242 3627 1243 3631
rect 1247 3627 1248 3631
rect 1242 3626 1248 3627
rect 1378 3631 1384 3632
rect 1378 3627 1379 3631
rect 1383 3627 1384 3631
rect 1378 3626 1384 3627
rect 1514 3631 1520 3632
rect 1514 3627 1515 3631
rect 1519 3627 1520 3631
rect 1934 3628 1935 3632
rect 1939 3628 1940 3632
rect 1934 3627 1940 3628
rect 1514 3626 1520 3627
rect 182 3616 188 3617
rect 110 3615 116 3616
rect 110 3611 111 3615
rect 115 3611 116 3615
rect 182 3612 183 3616
rect 187 3612 188 3616
rect 182 3611 188 3612
rect 318 3616 324 3617
rect 318 3612 319 3616
rect 323 3612 324 3616
rect 318 3611 324 3612
rect 454 3616 460 3617
rect 454 3612 455 3616
rect 459 3612 460 3616
rect 454 3611 460 3612
rect 590 3616 596 3617
rect 590 3612 591 3616
rect 595 3612 596 3616
rect 590 3611 596 3612
rect 726 3616 732 3617
rect 726 3612 727 3616
rect 731 3612 732 3616
rect 726 3611 732 3612
rect 862 3616 868 3617
rect 862 3612 863 3616
rect 867 3612 868 3616
rect 862 3611 868 3612
rect 998 3616 1004 3617
rect 998 3612 999 3616
rect 1003 3612 1004 3616
rect 998 3611 1004 3612
rect 1134 3616 1140 3617
rect 1134 3612 1135 3616
rect 1139 3612 1140 3616
rect 1134 3611 1140 3612
rect 1270 3616 1276 3617
rect 1270 3612 1271 3616
rect 1275 3612 1276 3616
rect 1270 3611 1276 3612
rect 1406 3616 1412 3617
rect 1406 3612 1407 3616
rect 1411 3612 1412 3616
rect 1406 3611 1412 3612
rect 1542 3616 1548 3617
rect 1542 3612 1543 3616
rect 1547 3612 1548 3616
rect 1542 3611 1548 3612
rect 1934 3615 1940 3616
rect 1934 3611 1935 3615
rect 1939 3611 1940 3615
rect 110 3610 116 3611
rect 112 3299 114 3610
rect 184 3299 186 3611
rect 320 3299 322 3611
rect 456 3299 458 3611
rect 592 3299 594 3611
rect 728 3299 730 3611
rect 864 3299 866 3611
rect 1000 3299 1002 3611
rect 1136 3299 1138 3611
rect 1272 3299 1274 3611
rect 1408 3299 1410 3611
rect 1544 3299 1546 3611
rect 1934 3610 1940 3611
rect 1936 3299 1938 3610
rect 1976 3575 1978 3647
rect 2020 3575 2022 3648
rect 2196 3575 2198 3648
rect 2380 3575 2382 3648
rect 2564 3575 2566 3648
rect 2756 3575 2758 3648
rect 2940 3575 2942 3648
rect 3124 3575 3126 3648
rect 3308 3575 3310 3648
rect 3492 3575 3494 3648
rect 3652 3575 3654 3648
rect 3798 3647 3804 3648
rect 3800 3575 3802 3647
rect 3840 3607 3842 3671
rect 4244 3607 4246 3672
rect 4444 3607 4446 3672
rect 4668 3607 4670 3672
rect 4908 3607 4910 3672
rect 5164 3607 5166 3672
rect 5420 3607 5422 3672
rect 5662 3671 5668 3672
rect 5664 3607 5666 3671
rect 3839 3606 3843 3607
rect 3839 3601 3843 3602
rect 3859 3606 3863 3607
rect 3859 3601 3863 3602
rect 3995 3606 3999 3607
rect 3995 3601 3999 3602
rect 4131 3606 4135 3607
rect 4131 3601 4135 3602
rect 4243 3606 4247 3607
rect 4243 3601 4247 3602
rect 4267 3606 4271 3607
rect 4267 3601 4271 3602
rect 4403 3606 4407 3607
rect 4403 3601 4407 3602
rect 4443 3606 4447 3607
rect 4443 3601 4447 3602
rect 4539 3606 4543 3607
rect 4539 3601 4543 3602
rect 4667 3606 4671 3607
rect 4667 3601 4671 3602
rect 4675 3606 4679 3607
rect 4675 3601 4679 3602
rect 4811 3606 4815 3607
rect 4811 3601 4815 3602
rect 4907 3606 4911 3607
rect 4907 3601 4911 3602
rect 4947 3606 4951 3607
rect 4947 3601 4951 3602
rect 5163 3606 5167 3607
rect 5163 3601 5167 3602
rect 5419 3606 5423 3607
rect 5419 3601 5423 3602
rect 5663 3606 5667 3607
rect 5663 3601 5667 3602
rect 1975 3574 1979 3575
rect 1975 3569 1979 3570
rect 2019 3574 2023 3575
rect 2019 3569 2023 3570
rect 2195 3574 2199 3575
rect 2195 3569 2199 3570
rect 2307 3574 2311 3575
rect 2307 3569 2311 3570
rect 2379 3574 2383 3575
rect 2379 3569 2383 3570
rect 2443 3574 2447 3575
rect 2443 3569 2447 3570
rect 2563 3574 2567 3575
rect 2563 3569 2567 3570
rect 2579 3574 2583 3575
rect 2579 3569 2583 3570
rect 2715 3574 2719 3575
rect 2715 3569 2719 3570
rect 2755 3574 2759 3575
rect 2755 3569 2759 3570
rect 2939 3574 2943 3575
rect 2939 3569 2943 3570
rect 3123 3574 3127 3575
rect 3123 3569 3127 3570
rect 3307 3574 3311 3575
rect 3307 3569 3311 3570
rect 3491 3574 3495 3575
rect 3491 3569 3495 3570
rect 3651 3574 3655 3575
rect 3651 3569 3655 3570
rect 3799 3574 3803 3575
rect 3799 3569 3803 3570
rect 1976 3509 1978 3569
rect 1974 3508 1980 3509
rect 2308 3508 2310 3569
rect 2444 3508 2446 3569
rect 2580 3508 2582 3569
rect 2716 3508 2718 3569
rect 3800 3509 3802 3569
rect 3840 3541 3842 3601
rect 3838 3540 3844 3541
rect 3860 3540 3862 3601
rect 3996 3540 3998 3601
rect 4132 3540 4134 3601
rect 4268 3540 4270 3601
rect 4404 3540 4406 3601
rect 4540 3540 4542 3601
rect 4676 3540 4678 3601
rect 4812 3540 4814 3601
rect 4948 3540 4950 3601
rect 5664 3541 5666 3601
rect 5662 3540 5668 3541
rect 3838 3536 3839 3540
rect 3843 3536 3844 3540
rect 3838 3535 3844 3536
rect 3858 3539 3864 3540
rect 3858 3535 3859 3539
rect 3863 3535 3864 3539
rect 3858 3534 3864 3535
rect 3994 3539 4000 3540
rect 3994 3535 3995 3539
rect 3999 3535 4000 3539
rect 3994 3534 4000 3535
rect 4130 3539 4136 3540
rect 4130 3535 4131 3539
rect 4135 3535 4136 3539
rect 4130 3534 4136 3535
rect 4266 3539 4272 3540
rect 4266 3535 4267 3539
rect 4271 3535 4272 3539
rect 4266 3534 4272 3535
rect 4402 3539 4408 3540
rect 4402 3535 4403 3539
rect 4407 3535 4408 3539
rect 4402 3534 4408 3535
rect 4538 3539 4544 3540
rect 4538 3535 4539 3539
rect 4543 3535 4544 3539
rect 4538 3534 4544 3535
rect 4674 3539 4680 3540
rect 4674 3535 4675 3539
rect 4679 3535 4680 3539
rect 4674 3534 4680 3535
rect 4810 3539 4816 3540
rect 4810 3535 4811 3539
rect 4815 3535 4816 3539
rect 4810 3534 4816 3535
rect 4946 3539 4952 3540
rect 4946 3535 4947 3539
rect 4951 3535 4952 3539
rect 5662 3536 5663 3540
rect 5667 3536 5668 3540
rect 5662 3535 5668 3536
rect 4946 3534 4952 3535
rect 3886 3524 3892 3525
rect 3838 3523 3844 3524
rect 3838 3519 3839 3523
rect 3843 3519 3844 3523
rect 3886 3520 3887 3524
rect 3891 3520 3892 3524
rect 3886 3519 3892 3520
rect 4022 3524 4028 3525
rect 4022 3520 4023 3524
rect 4027 3520 4028 3524
rect 4022 3519 4028 3520
rect 4158 3524 4164 3525
rect 4158 3520 4159 3524
rect 4163 3520 4164 3524
rect 4158 3519 4164 3520
rect 4294 3524 4300 3525
rect 4294 3520 4295 3524
rect 4299 3520 4300 3524
rect 4294 3519 4300 3520
rect 4430 3524 4436 3525
rect 4430 3520 4431 3524
rect 4435 3520 4436 3524
rect 4430 3519 4436 3520
rect 4566 3524 4572 3525
rect 4566 3520 4567 3524
rect 4571 3520 4572 3524
rect 4566 3519 4572 3520
rect 4702 3524 4708 3525
rect 4702 3520 4703 3524
rect 4707 3520 4708 3524
rect 4702 3519 4708 3520
rect 4838 3524 4844 3525
rect 4838 3520 4839 3524
rect 4843 3520 4844 3524
rect 4838 3519 4844 3520
rect 4974 3524 4980 3525
rect 4974 3520 4975 3524
rect 4979 3520 4980 3524
rect 4974 3519 4980 3520
rect 5662 3523 5668 3524
rect 5662 3519 5663 3523
rect 5667 3519 5668 3523
rect 3838 3518 3844 3519
rect 3798 3508 3804 3509
rect 1974 3504 1975 3508
rect 1979 3504 1980 3508
rect 1974 3503 1980 3504
rect 2306 3507 2312 3508
rect 2306 3503 2307 3507
rect 2311 3503 2312 3507
rect 2306 3502 2312 3503
rect 2442 3507 2448 3508
rect 2442 3503 2443 3507
rect 2447 3503 2448 3507
rect 2442 3502 2448 3503
rect 2578 3507 2584 3508
rect 2578 3503 2579 3507
rect 2583 3503 2584 3507
rect 2578 3502 2584 3503
rect 2714 3507 2720 3508
rect 2714 3503 2715 3507
rect 2719 3503 2720 3507
rect 3798 3504 3799 3508
rect 3803 3504 3804 3508
rect 3798 3503 3804 3504
rect 2714 3502 2720 3503
rect 3840 3495 3842 3518
rect 3888 3495 3890 3519
rect 4024 3495 4026 3519
rect 4160 3495 4162 3519
rect 4296 3495 4298 3519
rect 4432 3495 4434 3519
rect 4568 3495 4570 3519
rect 4704 3495 4706 3519
rect 4840 3495 4842 3519
rect 4976 3495 4978 3519
rect 5662 3518 5668 3519
rect 5664 3495 5666 3518
rect 3839 3494 3843 3495
rect 2334 3492 2340 3493
rect 1974 3491 1980 3492
rect 1974 3487 1975 3491
rect 1979 3487 1980 3491
rect 2334 3488 2335 3492
rect 2339 3488 2340 3492
rect 2334 3487 2340 3488
rect 2470 3492 2476 3493
rect 2470 3488 2471 3492
rect 2475 3488 2476 3492
rect 2470 3487 2476 3488
rect 2606 3492 2612 3493
rect 2606 3488 2607 3492
rect 2611 3488 2612 3492
rect 2606 3487 2612 3488
rect 2742 3492 2748 3493
rect 2742 3488 2743 3492
rect 2747 3488 2748 3492
rect 2742 3487 2748 3488
rect 3798 3491 3804 3492
rect 3798 3487 3799 3491
rect 3803 3487 3804 3491
rect 3839 3489 3843 3490
rect 3887 3494 3891 3495
rect 3887 3489 3891 3490
rect 4023 3494 4027 3495
rect 4023 3489 4027 3490
rect 4159 3494 4163 3495
rect 4159 3489 4163 3490
rect 4295 3494 4299 3495
rect 4295 3489 4299 3490
rect 4431 3494 4435 3495
rect 4431 3489 4435 3490
rect 4567 3494 4571 3495
rect 4567 3489 4571 3490
rect 4703 3494 4707 3495
rect 4703 3489 4707 3490
rect 4839 3494 4843 3495
rect 4839 3489 4843 3490
rect 4975 3494 4979 3495
rect 4975 3489 4979 3490
rect 5111 3494 5115 3495
rect 5111 3489 5115 3490
rect 5247 3494 5251 3495
rect 5247 3489 5251 3490
rect 5383 3494 5387 3495
rect 5383 3489 5387 3490
rect 5519 3494 5523 3495
rect 5519 3489 5523 3490
rect 5663 3494 5667 3495
rect 5663 3489 5667 3490
rect 1974 3486 1980 3487
rect 1976 3427 1978 3486
rect 2336 3427 2338 3487
rect 2472 3427 2474 3487
rect 2608 3427 2610 3487
rect 2744 3427 2746 3487
rect 3798 3486 3804 3487
rect 3800 3427 3802 3486
rect 3840 3466 3842 3489
rect 3838 3465 3844 3466
rect 3888 3465 3890 3489
rect 4024 3465 4026 3489
rect 4160 3465 4162 3489
rect 4296 3465 4298 3489
rect 4432 3465 4434 3489
rect 4568 3465 4570 3489
rect 4704 3465 4706 3489
rect 4840 3465 4842 3489
rect 4976 3465 4978 3489
rect 5112 3465 5114 3489
rect 5248 3465 5250 3489
rect 5384 3465 5386 3489
rect 5520 3465 5522 3489
rect 5664 3466 5666 3489
rect 5662 3465 5668 3466
rect 3838 3461 3839 3465
rect 3843 3461 3844 3465
rect 3838 3460 3844 3461
rect 3886 3464 3892 3465
rect 3886 3460 3887 3464
rect 3891 3460 3892 3464
rect 3886 3459 3892 3460
rect 4022 3464 4028 3465
rect 4022 3460 4023 3464
rect 4027 3460 4028 3464
rect 4022 3459 4028 3460
rect 4158 3464 4164 3465
rect 4158 3460 4159 3464
rect 4163 3460 4164 3464
rect 4158 3459 4164 3460
rect 4294 3464 4300 3465
rect 4294 3460 4295 3464
rect 4299 3460 4300 3464
rect 4294 3459 4300 3460
rect 4430 3464 4436 3465
rect 4430 3460 4431 3464
rect 4435 3460 4436 3464
rect 4430 3459 4436 3460
rect 4566 3464 4572 3465
rect 4566 3460 4567 3464
rect 4571 3460 4572 3464
rect 4566 3459 4572 3460
rect 4702 3464 4708 3465
rect 4702 3460 4703 3464
rect 4707 3460 4708 3464
rect 4702 3459 4708 3460
rect 4838 3464 4844 3465
rect 4838 3460 4839 3464
rect 4843 3460 4844 3464
rect 4838 3459 4844 3460
rect 4974 3464 4980 3465
rect 4974 3460 4975 3464
rect 4979 3460 4980 3464
rect 4974 3459 4980 3460
rect 5110 3464 5116 3465
rect 5110 3460 5111 3464
rect 5115 3460 5116 3464
rect 5110 3459 5116 3460
rect 5246 3464 5252 3465
rect 5246 3460 5247 3464
rect 5251 3460 5252 3464
rect 5246 3459 5252 3460
rect 5382 3464 5388 3465
rect 5382 3460 5383 3464
rect 5387 3460 5388 3464
rect 5382 3459 5388 3460
rect 5518 3464 5524 3465
rect 5518 3460 5519 3464
rect 5523 3460 5524 3464
rect 5662 3461 5663 3465
rect 5667 3461 5668 3465
rect 5662 3460 5668 3461
rect 5518 3459 5524 3460
rect 3858 3449 3864 3450
rect 3838 3448 3844 3449
rect 3838 3444 3839 3448
rect 3843 3444 3844 3448
rect 3858 3445 3859 3449
rect 3863 3445 3864 3449
rect 3858 3444 3864 3445
rect 3994 3449 4000 3450
rect 3994 3445 3995 3449
rect 3999 3445 4000 3449
rect 3994 3444 4000 3445
rect 4130 3449 4136 3450
rect 4130 3445 4131 3449
rect 4135 3445 4136 3449
rect 4130 3444 4136 3445
rect 4266 3449 4272 3450
rect 4266 3445 4267 3449
rect 4271 3445 4272 3449
rect 4266 3444 4272 3445
rect 4402 3449 4408 3450
rect 4402 3445 4403 3449
rect 4407 3445 4408 3449
rect 4402 3444 4408 3445
rect 4538 3449 4544 3450
rect 4538 3445 4539 3449
rect 4543 3445 4544 3449
rect 4538 3444 4544 3445
rect 4674 3449 4680 3450
rect 4674 3445 4675 3449
rect 4679 3445 4680 3449
rect 4674 3444 4680 3445
rect 4810 3449 4816 3450
rect 4810 3445 4811 3449
rect 4815 3445 4816 3449
rect 4810 3444 4816 3445
rect 4946 3449 4952 3450
rect 4946 3445 4947 3449
rect 4951 3445 4952 3449
rect 4946 3444 4952 3445
rect 5082 3449 5088 3450
rect 5082 3445 5083 3449
rect 5087 3445 5088 3449
rect 5082 3444 5088 3445
rect 5218 3449 5224 3450
rect 5218 3445 5219 3449
rect 5223 3445 5224 3449
rect 5218 3444 5224 3445
rect 5354 3449 5360 3450
rect 5354 3445 5355 3449
rect 5359 3445 5360 3449
rect 5354 3444 5360 3445
rect 5490 3449 5496 3450
rect 5490 3445 5491 3449
rect 5495 3445 5496 3449
rect 5490 3444 5496 3445
rect 5662 3448 5668 3449
rect 5662 3444 5663 3448
rect 5667 3444 5668 3448
rect 3838 3443 3844 3444
rect 1975 3426 1979 3427
rect 1975 3421 1979 3422
rect 2167 3426 2171 3427
rect 2167 3421 2171 3422
rect 2303 3426 2307 3427
rect 2303 3421 2307 3422
rect 2335 3426 2339 3427
rect 2335 3421 2339 3422
rect 2439 3426 2443 3427
rect 2439 3421 2443 3422
rect 2471 3426 2475 3427
rect 2471 3421 2475 3422
rect 2575 3426 2579 3427
rect 2575 3421 2579 3422
rect 2607 3426 2611 3427
rect 2607 3421 2611 3422
rect 2711 3426 2715 3427
rect 2711 3421 2715 3422
rect 2743 3426 2747 3427
rect 2743 3421 2747 3422
rect 2847 3426 2851 3427
rect 2847 3421 2851 3422
rect 2983 3426 2987 3427
rect 2983 3421 2987 3422
rect 3799 3426 3803 3427
rect 3799 3421 3803 3422
rect 1976 3398 1978 3421
rect 1974 3397 1980 3398
rect 2168 3397 2170 3421
rect 2304 3397 2306 3421
rect 2440 3397 2442 3421
rect 2576 3397 2578 3421
rect 2712 3397 2714 3421
rect 2848 3397 2850 3421
rect 2984 3397 2986 3421
rect 3800 3398 3802 3421
rect 3798 3397 3804 3398
rect 1974 3393 1975 3397
rect 1979 3393 1980 3397
rect 1974 3392 1980 3393
rect 2166 3396 2172 3397
rect 2166 3392 2167 3396
rect 2171 3392 2172 3396
rect 2166 3391 2172 3392
rect 2302 3396 2308 3397
rect 2302 3392 2303 3396
rect 2307 3392 2308 3396
rect 2302 3391 2308 3392
rect 2438 3396 2444 3397
rect 2438 3392 2439 3396
rect 2443 3392 2444 3396
rect 2438 3391 2444 3392
rect 2574 3396 2580 3397
rect 2574 3392 2575 3396
rect 2579 3392 2580 3396
rect 2574 3391 2580 3392
rect 2710 3396 2716 3397
rect 2710 3392 2711 3396
rect 2715 3392 2716 3396
rect 2710 3391 2716 3392
rect 2846 3396 2852 3397
rect 2846 3392 2847 3396
rect 2851 3392 2852 3396
rect 2846 3391 2852 3392
rect 2982 3396 2988 3397
rect 2982 3392 2983 3396
rect 2987 3392 2988 3396
rect 3798 3393 3799 3397
rect 3803 3393 3804 3397
rect 3798 3392 3804 3393
rect 2982 3391 2988 3392
rect 2138 3381 2144 3382
rect 1974 3380 1980 3381
rect 1974 3376 1975 3380
rect 1979 3376 1980 3380
rect 2138 3377 2139 3381
rect 2143 3377 2144 3381
rect 2138 3376 2144 3377
rect 2274 3381 2280 3382
rect 2274 3377 2275 3381
rect 2279 3377 2280 3381
rect 2274 3376 2280 3377
rect 2410 3381 2416 3382
rect 2410 3377 2411 3381
rect 2415 3377 2416 3381
rect 2410 3376 2416 3377
rect 2546 3381 2552 3382
rect 2546 3377 2547 3381
rect 2551 3377 2552 3381
rect 2546 3376 2552 3377
rect 2682 3381 2688 3382
rect 2682 3377 2683 3381
rect 2687 3377 2688 3381
rect 2682 3376 2688 3377
rect 2818 3381 2824 3382
rect 2818 3377 2819 3381
rect 2823 3377 2824 3381
rect 2818 3376 2824 3377
rect 2954 3381 2960 3382
rect 2954 3377 2955 3381
rect 2959 3377 2960 3381
rect 2954 3376 2960 3377
rect 3798 3380 3804 3381
rect 3798 3376 3799 3380
rect 3803 3376 3804 3380
rect 1974 3375 1980 3376
rect 1976 3315 1978 3375
rect 2140 3315 2142 3376
rect 2276 3315 2278 3376
rect 2412 3315 2414 3376
rect 2548 3315 2550 3376
rect 2684 3315 2686 3376
rect 2820 3315 2822 3376
rect 2956 3315 2958 3376
rect 3798 3375 3804 3376
rect 3840 3375 3842 3443
rect 3860 3375 3862 3444
rect 3996 3375 3998 3444
rect 4132 3375 4134 3444
rect 4268 3375 4270 3444
rect 4404 3375 4406 3444
rect 4540 3375 4542 3444
rect 4676 3375 4678 3444
rect 4812 3375 4814 3444
rect 4948 3375 4950 3444
rect 5084 3375 5086 3444
rect 5220 3375 5222 3444
rect 5356 3375 5358 3444
rect 5492 3375 5494 3444
rect 5662 3443 5668 3444
rect 5664 3375 5666 3443
rect 3800 3315 3802 3375
rect 3839 3374 3843 3375
rect 3839 3369 3843 3370
rect 3859 3374 3863 3375
rect 3859 3369 3863 3370
rect 3995 3374 3999 3375
rect 3995 3369 3999 3370
rect 4131 3374 4135 3375
rect 4131 3369 4135 3370
rect 4155 3374 4159 3375
rect 4155 3369 4159 3370
rect 4267 3374 4271 3375
rect 4267 3369 4271 3370
rect 4315 3374 4319 3375
rect 4315 3369 4319 3370
rect 4403 3374 4407 3375
rect 4403 3369 4407 3370
rect 4467 3374 4471 3375
rect 4467 3369 4471 3370
rect 4539 3374 4543 3375
rect 4539 3369 4543 3370
rect 4627 3374 4631 3375
rect 4627 3369 4631 3370
rect 4675 3374 4679 3375
rect 4675 3369 4679 3370
rect 4787 3374 4791 3375
rect 4787 3369 4791 3370
rect 4811 3374 4815 3375
rect 4811 3369 4815 3370
rect 4947 3374 4951 3375
rect 4947 3369 4951 3370
rect 5083 3374 5087 3375
rect 5083 3369 5087 3370
rect 5219 3374 5223 3375
rect 5219 3369 5223 3370
rect 5355 3374 5359 3375
rect 5355 3369 5359 3370
rect 5491 3374 5495 3375
rect 5491 3369 5495 3370
rect 5663 3374 5667 3375
rect 5663 3369 5667 3370
rect 1975 3314 1979 3315
rect 1975 3309 1979 3310
rect 2059 3314 2063 3315
rect 2059 3309 2063 3310
rect 2139 3314 2143 3315
rect 2139 3309 2143 3310
rect 2203 3314 2207 3315
rect 2203 3309 2207 3310
rect 2275 3314 2279 3315
rect 2275 3309 2279 3310
rect 2363 3314 2367 3315
rect 2363 3309 2367 3310
rect 2411 3314 2415 3315
rect 2411 3309 2415 3310
rect 2539 3314 2543 3315
rect 2539 3309 2543 3310
rect 2547 3314 2551 3315
rect 2547 3309 2551 3310
rect 2683 3314 2687 3315
rect 2683 3309 2687 3310
rect 2739 3314 2743 3315
rect 2739 3309 2743 3310
rect 2819 3314 2823 3315
rect 2819 3309 2823 3310
rect 2955 3314 2959 3315
rect 2955 3309 2959 3310
rect 3187 3314 3191 3315
rect 3187 3309 3191 3310
rect 3427 3314 3431 3315
rect 3427 3309 3431 3310
rect 3651 3314 3655 3315
rect 3651 3309 3655 3310
rect 3799 3314 3803 3315
rect 3799 3309 3803 3310
rect 3840 3309 3842 3369
rect 111 3298 115 3299
rect 111 3293 115 3294
rect 159 3298 163 3299
rect 159 3293 163 3294
rect 183 3298 187 3299
rect 183 3293 187 3294
rect 295 3298 299 3299
rect 295 3293 299 3294
rect 319 3298 323 3299
rect 319 3293 323 3294
rect 431 3298 435 3299
rect 431 3293 435 3294
rect 455 3298 459 3299
rect 455 3293 459 3294
rect 567 3298 571 3299
rect 567 3293 571 3294
rect 591 3298 595 3299
rect 591 3293 595 3294
rect 703 3298 707 3299
rect 703 3293 707 3294
rect 727 3298 731 3299
rect 727 3293 731 3294
rect 839 3298 843 3299
rect 839 3293 843 3294
rect 863 3298 867 3299
rect 863 3293 867 3294
rect 975 3298 979 3299
rect 975 3293 979 3294
rect 999 3298 1003 3299
rect 999 3293 1003 3294
rect 1111 3298 1115 3299
rect 1111 3293 1115 3294
rect 1135 3298 1139 3299
rect 1135 3293 1139 3294
rect 1247 3298 1251 3299
rect 1247 3293 1251 3294
rect 1271 3298 1275 3299
rect 1271 3293 1275 3294
rect 1383 3298 1387 3299
rect 1383 3293 1387 3294
rect 1407 3298 1411 3299
rect 1407 3293 1411 3294
rect 1519 3298 1523 3299
rect 1519 3293 1523 3294
rect 1543 3298 1547 3299
rect 1543 3293 1547 3294
rect 1935 3298 1939 3299
rect 1935 3293 1939 3294
rect 112 3270 114 3293
rect 110 3269 116 3270
rect 160 3269 162 3293
rect 296 3269 298 3293
rect 432 3269 434 3293
rect 568 3269 570 3293
rect 704 3269 706 3293
rect 840 3269 842 3293
rect 976 3269 978 3293
rect 1112 3269 1114 3293
rect 1248 3269 1250 3293
rect 1384 3269 1386 3293
rect 1520 3269 1522 3293
rect 1936 3270 1938 3293
rect 1934 3269 1940 3270
rect 110 3265 111 3269
rect 115 3265 116 3269
rect 110 3264 116 3265
rect 158 3268 164 3269
rect 158 3264 159 3268
rect 163 3264 164 3268
rect 158 3263 164 3264
rect 294 3268 300 3269
rect 294 3264 295 3268
rect 299 3264 300 3268
rect 294 3263 300 3264
rect 430 3268 436 3269
rect 430 3264 431 3268
rect 435 3264 436 3268
rect 430 3263 436 3264
rect 566 3268 572 3269
rect 566 3264 567 3268
rect 571 3264 572 3268
rect 566 3263 572 3264
rect 702 3268 708 3269
rect 702 3264 703 3268
rect 707 3264 708 3268
rect 702 3263 708 3264
rect 838 3268 844 3269
rect 838 3264 839 3268
rect 843 3264 844 3268
rect 838 3263 844 3264
rect 974 3268 980 3269
rect 974 3264 975 3268
rect 979 3264 980 3268
rect 974 3263 980 3264
rect 1110 3268 1116 3269
rect 1110 3264 1111 3268
rect 1115 3264 1116 3268
rect 1110 3263 1116 3264
rect 1246 3268 1252 3269
rect 1246 3264 1247 3268
rect 1251 3264 1252 3268
rect 1246 3263 1252 3264
rect 1382 3268 1388 3269
rect 1382 3264 1383 3268
rect 1387 3264 1388 3268
rect 1382 3263 1388 3264
rect 1518 3268 1524 3269
rect 1518 3264 1519 3268
rect 1523 3264 1524 3268
rect 1934 3265 1935 3269
rect 1939 3265 1940 3269
rect 1934 3264 1940 3265
rect 1518 3263 1524 3264
rect 130 3253 136 3254
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 130 3249 131 3253
rect 135 3249 136 3253
rect 130 3248 136 3249
rect 266 3253 272 3254
rect 266 3249 267 3253
rect 271 3249 272 3253
rect 266 3248 272 3249
rect 402 3253 408 3254
rect 402 3249 403 3253
rect 407 3249 408 3253
rect 402 3248 408 3249
rect 538 3253 544 3254
rect 538 3249 539 3253
rect 543 3249 544 3253
rect 538 3248 544 3249
rect 674 3253 680 3254
rect 674 3249 675 3253
rect 679 3249 680 3253
rect 674 3248 680 3249
rect 810 3253 816 3254
rect 810 3249 811 3253
rect 815 3249 816 3253
rect 810 3248 816 3249
rect 946 3253 952 3254
rect 946 3249 947 3253
rect 951 3249 952 3253
rect 946 3248 952 3249
rect 1082 3253 1088 3254
rect 1082 3249 1083 3253
rect 1087 3249 1088 3253
rect 1082 3248 1088 3249
rect 1218 3253 1224 3254
rect 1218 3249 1219 3253
rect 1223 3249 1224 3253
rect 1218 3248 1224 3249
rect 1354 3253 1360 3254
rect 1354 3249 1355 3253
rect 1359 3249 1360 3253
rect 1354 3248 1360 3249
rect 1490 3253 1496 3254
rect 1490 3249 1491 3253
rect 1495 3249 1496 3253
rect 1490 3248 1496 3249
rect 1934 3252 1940 3253
rect 1934 3248 1935 3252
rect 1939 3248 1940 3252
rect 1976 3249 1978 3309
rect 110 3247 116 3248
rect 112 3159 114 3247
rect 132 3159 134 3248
rect 268 3159 270 3248
rect 404 3159 406 3248
rect 540 3159 542 3248
rect 676 3159 678 3248
rect 812 3159 814 3248
rect 948 3159 950 3248
rect 1084 3159 1086 3248
rect 1220 3159 1222 3248
rect 1356 3159 1358 3248
rect 1492 3159 1494 3248
rect 1934 3247 1940 3248
rect 1974 3248 1980 3249
rect 2060 3248 2062 3309
rect 2204 3248 2206 3309
rect 2364 3248 2366 3309
rect 2540 3248 2542 3309
rect 2740 3248 2742 3309
rect 2956 3248 2958 3309
rect 3188 3248 3190 3309
rect 3428 3248 3430 3309
rect 3652 3248 3654 3309
rect 3800 3249 3802 3309
rect 3838 3308 3844 3309
rect 3860 3308 3862 3369
rect 3996 3308 3998 3369
rect 4156 3308 4158 3369
rect 4316 3308 4318 3369
rect 4468 3308 4470 3369
rect 4628 3308 4630 3369
rect 4788 3308 4790 3369
rect 4948 3308 4950 3369
rect 5664 3309 5666 3369
rect 5662 3308 5668 3309
rect 3838 3304 3839 3308
rect 3843 3304 3844 3308
rect 3838 3303 3844 3304
rect 3858 3307 3864 3308
rect 3858 3303 3859 3307
rect 3863 3303 3864 3307
rect 3858 3302 3864 3303
rect 3994 3307 4000 3308
rect 3994 3303 3995 3307
rect 3999 3303 4000 3307
rect 3994 3302 4000 3303
rect 4154 3307 4160 3308
rect 4154 3303 4155 3307
rect 4159 3303 4160 3307
rect 4154 3302 4160 3303
rect 4314 3307 4320 3308
rect 4314 3303 4315 3307
rect 4319 3303 4320 3307
rect 4314 3302 4320 3303
rect 4466 3307 4472 3308
rect 4466 3303 4467 3307
rect 4471 3303 4472 3307
rect 4466 3302 4472 3303
rect 4626 3307 4632 3308
rect 4626 3303 4627 3307
rect 4631 3303 4632 3307
rect 4626 3302 4632 3303
rect 4786 3307 4792 3308
rect 4786 3303 4787 3307
rect 4791 3303 4792 3307
rect 4786 3302 4792 3303
rect 4946 3307 4952 3308
rect 4946 3303 4947 3307
rect 4951 3303 4952 3307
rect 5662 3304 5663 3308
rect 5667 3304 5668 3308
rect 5662 3303 5668 3304
rect 4946 3302 4952 3303
rect 3886 3292 3892 3293
rect 3838 3291 3844 3292
rect 3838 3287 3839 3291
rect 3843 3287 3844 3291
rect 3886 3288 3887 3292
rect 3891 3288 3892 3292
rect 3886 3287 3892 3288
rect 4022 3292 4028 3293
rect 4022 3288 4023 3292
rect 4027 3288 4028 3292
rect 4022 3287 4028 3288
rect 4182 3292 4188 3293
rect 4182 3288 4183 3292
rect 4187 3288 4188 3292
rect 4182 3287 4188 3288
rect 4342 3292 4348 3293
rect 4342 3288 4343 3292
rect 4347 3288 4348 3292
rect 4342 3287 4348 3288
rect 4494 3292 4500 3293
rect 4494 3288 4495 3292
rect 4499 3288 4500 3292
rect 4494 3287 4500 3288
rect 4654 3292 4660 3293
rect 4654 3288 4655 3292
rect 4659 3288 4660 3292
rect 4654 3287 4660 3288
rect 4814 3292 4820 3293
rect 4814 3288 4815 3292
rect 4819 3288 4820 3292
rect 4814 3287 4820 3288
rect 4974 3292 4980 3293
rect 4974 3288 4975 3292
rect 4979 3288 4980 3292
rect 4974 3287 4980 3288
rect 5662 3291 5668 3292
rect 5662 3287 5663 3291
rect 5667 3287 5668 3291
rect 3838 3286 3844 3287
rect 3840 3251 3842 3286
rect 3888 3251 3890 3287
rect 4024 3251 4026 3287
rect 4184 3251 4186 3287
rect 4344 3251 4346 3287
rect 4496 3251 4498 3287
rect 4656 3251 4658 3287
rect 4816 3251 4818 3287
rect 4976 3251 4978 3287
rect 5662 3286 5668 3287
rect 5664 3251 5666 3286
rect 3839 3250 3843 3251
rect 3798 3248 3804 3249
rect 1936 3159 1938 3247
rect 1974 3244 1975 3248
rect 1979 3244 1980 3248
rect 1974 3243 1980 3244
rect 2058 3247 2064 3248
rect 2058 3243 2059 3247
rect 2063 3243 2064 3247
rect 2058 3242 2064 3243
rect 2202 3247 2208 3248
rect 2202 3243 2203 3247
rect 2207 3243 2208 3247
rect 2202 3242 2208 3243
rect 2362 3247 2368 3248
rect 2362 3243 2363 3247
rect 2367 3243 2368 3247
rect 2362 3242 2368 3243
rect 2538 3247 2544 3248
rect 2538 3243 2539 3247
rect 2543 3243 2544 3247
rect 2538 3242 2544 3243
rect 2738 3247 2744 3248
rect 2738 3243 2739 3247
rect 2743 3243 2744 3247
rect 2738 3242 2744 3243
rect 2954 3247 2960 3248
rect 2954 3243 2955 3247
rect 2959 3243 2960 3247
rect 2954 3242 2960 3243
rect 3186 3247 3192 3248
rect 3186 3243 3187 3247
rect 3191 3243 3192 3247
rect 3186 3242 3192 3243
rect 3426 3247 3432 3248
rect 3426 3243 3427 3247
rect 3431 3243 3432 3247
rect 3426 3242 3432 3243
rect 3650 3247 3656 3248
rect 3650 3243 3651 3247
rect 3655 3243 3656 3247
rect 3798 3244 3799 3248
rect 3803 3244 3804 3248
rect 3839 3245 3843 3246
rect 3887 3250 3891 3251
rect 3887 3245 3891 3246
rect 4023 3250 4027 3251
rect 4023 3245 4027 3246
rect 4183 3250 4187 3251
rect 4183 3245 4187 3246
rect 4343 3250 4347 3251
rect 4343 3245 4347 3246
rect 4495 3250 4499 3251
rect 4495 3245 4499 3246
rect 4655 3250 4659 3251
rect 4655 3245 4659 3246
rect 4807 3250 4811 3251
rect 4807 3245 4811 3246
rect 4815 3250 4819 3251
rect 4815 3245 4819 3246
rect 4943 3250 4947 3251
rect 4943 3245 4947 3246
rect 4975 3250 4979 3251
rect 4975 3245 4979 3246
rect 5079 3250 5083 3251
rect 5079 3245 5083 3246
rect 5215 3250 5219 3251
rect 5215 3245 5219 3246
rect 5351 3250 5355 3251
rect 5351 3245 5355 3246
rect 5663 3250 5667 3251
rect 5663 3245 5667 3246
rect 3798 3243 3804 3244
rect 3650 3242 3656 3243
rect 2086 3232 2092 3233
rect 1974 3231 1980 3232
rect 1974 3227 1975 3231
rect 1979 3227 1980 3231
rect 2086 3228 2087 3232
rect 2091 3228 2092 3232
rect 2086 3227 2092 3228
rect 2230 3232 2236 3233
rect 2230 3228 2231 3232
rect 2235 3228 2236 3232
rect 2230 3227 2236 3228
rect 2390 3232 2396 3233
rect 2390 3228 2391 3232
rect 2395 3228 2396 3232
rect 2390 3227 2396 3228
rect 2566 3232 2572 3233
rect 2566 3228 2567 3232
rect 2571 3228 2572 3232
rect 2566 3227 2572 3228
rect 2766 3232 2772 3233
rect 2766 3228 2767 3232
rect 2771 3228 2772 3232
rect 2766 3227 2772 3228
rect 2982 3232 2988 3233
rect 2982 3228 2983 3232
rect 2987 3228 2988 3232
rect 2982 3227 2988 3228
rect 3214 3232 3220 3233
rect 3214 3228 3215 3232
rect 3219 3228 3220 3232
rect 3214 3227 3220 3228
rect 3454 3232 3460 3233
rect 3454 3228 3455 3232
rect 3459 3228 3460 3232
rect 3454 3227 3460 3228
rect 3678 3232 3684 3233
rect 3678 3228 3679 3232
rect 3683 3228 3684 3232
rect 3678 3227 3684 3228
rect 3798 3231 3804 3232
rect 3798 3227 3799 3231
rect 3803 3227 3804 3231
rect 1974 3226 1980 3227
rect 1976 3199 1978 3226
rect 2088 3199 2090 3227
rect 2232 3199 2234 3227
rect 2392 3199 2394 3227
rect 2568 3199 2570 3227
rect 2768 3199 2770 3227
rect 2984 3199 2986 3227
rect 3216 3199 3218 3227
rect 3456 3199 3458 3227
rect 3680 3199 3682 3227
rect 3798 3226 3804 3227
rect 3800 3199 3802 3226
rect 3840 3222 3842 3245
rect 3838 3221 3844 3222
rect 4808 3221 4810 3245
rect 4944 3221 4946 3245
rect 5080 3221 5082 3245
rect 5216 3221 5218 3245
rect 5352 3221 5354 3245
rect 5664 3222 5666 3245
rect 5662 3221 5668 3222
rect 3838 3217 3839 3221
rect 3843 3217 3844 3221
rect 3838 3216 3844 3217
rect 4806 3220 4812 3221
rect 4806 3216 4807 3220
rect 4811 3216 4812 3220
rect 4806 3215 4812 3216
rect 4942 3220 4948 3221
rect 4942 3216 4943 3220
rect 4947 3216 4948 3220
rect 4942 3215 4948 3216
rect 5078 3220 5084 3221
rect 5078 3216 5079 3220
rect 5083 3216 5084 3220
rect 5078 3215 5084 3216
rect 5214 3220 5220 3221
rect 5214 3216 5215 3220
rect 5219 3216 5220 3220
rect 5214 3215 5220 3216
rect 5350 3220 5356 3221
rect 5350 3216 5351 3220
rect 5355 3216 5356 3220
rect 5662 3217 5663 3221
rect 5667 3217 5668 3221
rect 5662 3216 5668 3217
rect 5350 3215 5356 3216
rect 4778 3205 4784 3206
rect 3838 3204 3844 3205
rect 3838 3200 3839 3204
rect 3843 3200 3844 3204
rect 4778 3201 4779 3205
rect 4783 3201 4784 3205
rect 4778 3200 4784 3201
rect 4914 3205 4920 3206
rect 4914 3201 4915 3205
rect 4919 3201 4920 3205
rect 4914 3200 4920 3201
rect 5050 3205 5056 3206
rect 5050 3201 5051 3205
rect 5055 3201 5056 3205
rect 5050 3200 5056 3201
rect 5186 3205 5192 3206
rect 5186 3201 5187 3205
rect 5191 3201 5192 3205
rect 5186 3200 5192 3201
rect 5322 3205 5328 3206
rect 5322 3201 5323 3205
rect 5327 3201 5328 3205
rect 5322 3200 5328 3201
rect 5662 3204 5668 3205
rect 5662 3200 5663 3204
rect 5667 3200 5668 3204
rect 3838 3199 3844 3200
rect 1975 3198 1979 3199
rect 1975 3193 1979 3194
rect 2023 3198 2027 3199
rect 2023 3193 2027 3194
rect 2087 3198 2091 3199
rect 2087 3193 2091 3194
rect 2159 3198 2163 3199
rect 2159 3193 2163 3194
rect 2231 3198 2235 3199
rect 2231 3193 2235 3194
rect 2303 3198 2307 3199
rect 2303 3193 2307 3194
rect 2391 3198 2395 3199
rect 2391 3193 2395 3194
rect 2455 3198 2459 3199
rect 2455 3193 2459 3194
rect 2567 3198 2571 3199
rect 2567 3193 2571 3194
rect 2615 3198 2619 3199
rect 2615 3193 2619 3194
rect 2767 3198 2771 3199
rect 2767 3193 2771 3194
rect 2783 3198 2787 3199
rect 2783 3193 2787 3194
rect 2951 3198 2955 3199
rect 2951 3193 2955 3194
rect 2983 3198 2987 3199
rect 2983 3193 2987 3194
rect 3127 3198 3131 3199
rect 3127 3193 3131 3194
rect 3215 3198 3219 3199
rect 3215 3193 3219 3194
rect 3311 3198 3315 3199
rect 3311 3193 3315 3194
rect 3455 3198 3459 3199
rect 3455 3193 3459 3194
rect 3503 3198 3507 3199
rect 3503 3193 3507 3194
rect 3679 3198 3683 3199
rect 3679 3193 3683 3194
rect 3799 3198 3803 3199
rect 3799 3193 3803 3194
rect 1976 3170 1978 3193
rect 1974 3169 1980 3170
rect 2024 3169 2026 3193
rect 2160 3169 2162 3193
rect 2304 3169 2306 3193
rect 2456 3169 2458 3193
rect 2616 3169 2618 3193
rect 2784 3169 2786 3193
rect 2952 3169 2954 3193
rect 3128 3169 3130 3193
rect 3312 3169 3314 3193
rect 3504 3169 3506 3193
rect 3680 3169 3682 3193
rect 3800 3170 3802 3193
rect 3798 3169 3804 3170
rect 1974 3165 1975 3169
rect 1979 3165 1980 3169
rect 1974 3164 1980 3165
rect 2022 3168 2028 3169
rect 2022 3164 2023 3168
rect 2027 3164 2028 3168
rect 2022 3163 2028 3164
rect 2158 3168 2164 3169
rect 2158 3164 2159 3168
rect 2163 3164 2164 3168
rect 2158 3163 2164 3164
rect 2302 3168 2308 3169
rect 2302 3164 2303 3168
rect 2307 3164 2308 3168
rect 2302 3163 2308 3164
rect 2454 3168 2460 3169
rect 2454 3164 2455 3168
rect 2459 3164 2460 3168
rect 2454 3163 2460 3164
rect 2614 3168 2620 3169
rect 2614 3164 2615 3168
rect 2619 3164 2620 3168
rect 2614 3163 2620 3164
rect 2782 3168 2788 3169
rect 2782 3164 2783 3168
rect 2787 3164 2788 3168
rect 2782 3163 2788 3164
rect 2950 3168 2956 3169
rect 2950 3164 2951 3168
rect 2955 3164 2956 3168
rect 2950 3163 2956 3164
rect 3126 3168 3132 3169
rect 3126 3164 3127 3168
rect 3131 3164 3132 3168
rect 3126 3163 3132 3164
rect 3310 3168 3316 3169
rect 3310 3164 3311 3168
rect 3315 3164 3316 3168
rect 3310 3163 3316 3164
rect 3502 3168 3508 3169
rect 3502 3164 3503 3168
rect 3507 3164 3508 3168
rect 3502 3163 3508 3164
rect 3678 3168 3684 3169
rect 3678 3164 3679 3168
rect 3683 3164 3684 3168
rect 3798 3165 3799 3169
rect 3803 3165 3804 3169
rect 3798 3164 3804 3165
rect 3678 3163 3684 3164
rect 111 3158 115 3159
rect 111 3153 115 3154
rect 131 3158 135 3159
rect 131 3153 135 3154
rect 267 3158 271 3159
rect 267 3153 271 3154
rect 291 3158 295 3159
rect 291 3153 295 3154
rect 403 3158 407 3159
rect 403 3153 407 3154
rect 459 3158 463 3159
rect 459 3153 463 3154
rect 539 3158 543 3159
rect 539 3153 543 3154
rect 627 3158 631 3159
rect 627 3153 631 3154
rect 675 3158 679 3159
rect 675 3153 679 3154
rect 811 3158 815 3159
rect 811 3153 815 3154
rect 947 3158 951 3159
rect 947 3153 951 3154
rect 995 3158 999 3159
rect 995 3153 999 3154
rect 1083 3158 1087 3159
rect 1083 3153 1087 3154
rect 1187 3158 1191 3159
rect 1187 3153 1191 3154
rect 1219 3158 1223 3159
rect 1219 3153 1223 3154
rect 1355 3158 1359 3159
rect 1355 3153 1359 3154
rect 1387 3158 1391 3159
rect 1387 3153 1391 3154
rect 1491 3158 1495 3159
rect 1491 3153 1495 3154
rect 1595 3158 1599 3159
rect 1595 3153 1599 3154
rect 1787 3158 1791 3159
rect 1787 3153 1791 3154
rect 1935 3158 1939 3159
rect 1935 3153 1939 3154
rect 1994 3153 2000 3154
rect 112 3093 114 3153
rect 110 3092 116 3093
rect 292 3092 294 3153
rect 460 3092 462 3153
rect 628 3092 630 3153
rect 812 3092 814 3153
rect 996 3092 998 3153
rect 1188 3092 1190 3153
rect 1388 3092 1390 3153
rect 1596 3092 1598 3153
rect 1788 3092 1790 3153
rect 1936 3093 1938 3153
rect 1974 3152 1980 3153
rect 1974 3148 1975 3152
rect 1979 3148 1980 3152
rect 1994 3149 1995 3153
rect 1999 3149 2000 3153
rect 1994 3148 2000 3149
rect 2130 3153 2136 3154
rect 2130 3149 2131 3153
rect 2135 3149 2136 3153
rect 2130 3148 2136 3149
rect 2274 3153 2280 3154
rect 2274 3149 2275 3153
rect 2279 3149 2280 3153
rect 2274 3148 2280 3149
rect 2426 3153 2432 3154
rect 2426 3149 2427 3153
rect 2431 3149 2432 3153
rect 2426 3148 2432 3149
rect 2586 3153 2592 3154
rect 2586 3149 2587 3153
rect 2591 3149 2592 3153
rect 2586 3148 2592 3149
rect 2754 3153 2760 3154
rect 2754 3149 2755 3153
rect 2759 3149 2760 3153
rect 2754 3148 2760 3149
rect 2922 3153 2928 3154
rect 2922 3149 2923 3153
rect 2927 3149 2928 3153
rect 2922 3148 2928 3149
rect 3098 3153 3104 3154
rect 3098 3149 3099 3153
rect 3103 3149 3104 3153
rect 3098 3148 3104 3149
rect 3282 3153 3288 3154
rect 3282 3149 3283 3153
rect 3287 3149 3288 3153
rect 3282 3148 3288 3149
rect 3474 3153 3480 3154
rect 3474 3149 3475 3153
rect 3479 3149 3480 3153
rect 3474 3148 3480 3149
rect 3650 3153 3656 3154
rect 3650 3149 3651 3153
rect 3655 3149 3656 3153
rect 3650 3148 3656 3149
rect 3798 3152 3804 3153
rect 3798 3148 3799 3152
rect 3803 3148 3804 3152
rect 1974 3147 1980 3148
rect 1934 3092 1940 3093
rect 110 3088 111 3092
rect 115 3088 116 3092
rect 110 3087 116 3088
rect 290 3091 296 3092
rect 290 3087 291 3091
rect 295 3087 296 3091
rect 290 3086 296 3087
rect 458 3091 464 3092
rect 458 3087 459 3091
rect 463 3087 464 3091
rect 458 3086 464 3087
rect 626 3091 632 3092
rect 626 3087 627 3091
rect 631 3087 632 3091
rect 626 3086 632 3087
rect 810 3091 816 3092
rect 810 3087 811 3091
rect 815 3087 816 3091
rect 810 3086 816 3087
rect 994 3091 1000 3092
rect 994 3087 995 3091
rect 999 3087 1000 3091
rect 994 3086 1000 3087
rect 1186 3091 1192 3092
rect 1186 3087 1187 3091
rect 1191 3087 1192 3091
rect 1186 3086 1192 3087
rect 1386 3091 1392 3092
rect 1386 3087 1387 3091
rect 1391 3087 1392 3091
rect 1386 3086 1392 3087
rect 1594 3091 1600 3092
rect 1594 3087 1595 3091
rect 1599 3087 1600 3091
rect 1594 3086 1600 3087
rect 1786 3091 1792 3092
rect 1786 3087 1787 3091
rect 1791 3087 1792 3091
rect 1934 3088 1935 3092
rect 1939 3088 1940 3092
rect 1934 3087 1940 3088
rect 1786 3086 1792 3087
rect 318 3076 324 3077
rect 110 3075 116 3076
rect 110 3071 111 3075
rect 115 3071 116 3075
rect 318 3072 319 3076
rect 323 3072 324 3076
rect 318 3071 324 3072
rect 486 3076 492 3077
rect 486 3072 487 3076
rect 491 3072 492 3076
rect 486 3071 492 3072
rect 654 3076 660 3077
rect 654 3072 655 3076
rect 659 3072 660 3076
rect 654 3071 660 3072
rect 838 3076 844 3077
rect 838 3072 839 3076
rect 843 3072 844 3076
rect 838 3071 844 3072
rect 1022 3076 1028 3077
rect 1022 3072 1023 3076
rect 1027 3072 1028 3076
rect 1022 3071 1028 3072
rect 1214 3076 1220 3077
rect 1214 3072 1215 3076
rect 1219 3072 1220 3076
rect 1214 3071 1220 3072
rect 1414 3076 1420 3077
rect 1414 3072 1415 3076
rect 1419 3072 1420 3076
rect 1414 3071 1420 3072
rect 1622 3076 1628 3077
rect 1622 3072 1623 3076
rect 1627 3072 1628 3076
rect 1622 3071 1628 3072
rect 1814 3076 1820 3077
rect 1814 3072 1815 3076
rect 1819 3072 1820 3076
rect 1814 3071 1820 3072
rect 1934 3075 1940 3076
rect 1934 3071 1935 3075
rect 1939 3071 1940 3075
rect 110 3070 116 3071
rect 112 3047 114 3070
rect 320 3047 322 3071
rect 488 3047 490 3071
rect 656 3047 658 3071
rect 840 3047 842 3071
rect 1024 3047 1026 3071
rect 1216 3047 1218 3071
rect 1416 3047 1418 3071
rect 1624 3047 1626 3071
rect 1816 3047 1818 3071
rect 1934 3070 1940 3071
rect 1936 3047 1938 3070
rect 1976 3067 1978 3147
rect 1996 3067 1998 3148
rect 2132 3067 2134 3148
rect 2276 3067 2278 3148
rect 2428 3067 2430 3148
rect 2588 3067 2590 3148
rect 2756 3067 2758 3148
rect 2924 3067 2926 3148
rect 3100 3067 3102 3148
rect 3284 3067 3286 3148
rect 3476 3067 3478 3148
rect 3652 3067 3654 3148
rect 3798 3147 3804 3148
rect 3800 3067 3802 3147
rect 3840 3135 3842 3199
rect 4780 3135 4782 3200
rect 4916 3135 4918 3200
rect 5052 3135 5054 3200
rect 5188 3135 5190 3200
rect 5324 3135 5326 3200
rect 5662 3199 5668 3200
rect 5664 3135 5666 3199
rect 3839 3134 3843 3135
rect 3839 3129 3843 3130
rect 4699 3134 4703 3135
rect 4699 3129 4703 3130
rect 4779 3134 4783 3135
rect 4779 3129 4783 3130
rect 4835 3134 4839 3135
rect 4835 3129 4839 3130
rect 4915 3134 4919 3135
rect 4915 3129 4919 3130
rect 4971 3134 4975 3135
rect 4971 3129 4975 3130
rect 5051 3134 5055 3135
rect 5051 3129 5055 3130
rect 5107 3134 5111 3135
rect 5107 3129 5111 3130
rect 5187 3134 5191 3135
rect 5187 3129 5191 3130
rect 5243 3134 5247 3135
rect 5243 3129 5247 3130
rect 5323 3134 5327 3135
rect 5323 3129 5327 3130
rect 5379 3134 5383 3135
rect 5379 3129 5383 3130
rect 5515 3134 5519 3135
rect 5515 3129 5519 3130
rect 5663 3134 5667 3135
rect 5663 3129 5667 3130
rect 3840 3069 3842 3129
rect 3838 3068 3844 3069
rect 4700 3068 4702 3129
rect 4836 3068 4838 3129
rect 4972 3068 4974 3129
rect 5108 3068 5110 3129
rect 5244 3068 5246 3129
rect 5380 3068 5382 3129
rect 5516 3068 5518 3129
rect 5664 3069 5666 3129
rect 5662 3068 5668 3069
rect 1975 3066 1979 3067
rect 1975 3061 1979 3062
rect 1995 3066 1999 3067
rect 1995 3061 1999 3062
rect 2131 3066 2135 3067
rect 2131 3061 2135 3062
rect 2275 3066 2279 3067
rect 2275 3061 2279 3062
rect 2427 3066 2431 3067
rect 2427 3061 2431 3062
rect 2587 3066 2591 3067
rect 2587 3061 2591 3062
rect 2755 3066 2759 3067
rect 2755 3061 2759 3062
rect 2811 3066 2815 3067
rect 2811 3061 2815 3062
rect 2923 3066 2927 3067
rect 2923 3061 2927 3062
rect 3003 3066 3007 3067
rect 3003 3061 3007 3062
rect 3099 3066 3103 3067
rect 3099 3061 3103 3062
rect 3203 3066 3207 3067
rect 3203 3061 3207 3062
rect 3283 3066 3287 3067
rect 3283 3061 3287 3062
rect 3403 3066 3407 3067
rect 3403 3061 3407 3062
rect 3475 3066 3479 3067
rect 3475 3061 3479 3062
rect 3603 3066 3607 3067
rect 3603 3061 3607 3062
rect 3651 3066 3655 3067
rect 3651 3061 3655 3062
rect 3799 3066 3803 3067
rect 3838 3064 3839 3068
rect 3843 3064 3844 3068
rect 3838 3063 3844 3064
rect 4698 3067 4704 3068
rect 4698 3063 4699 3067
rect 4703 3063 4704 3067
rect 4698 3062 4704 3063
rect 4834 3067 4840 3068
rect 4834 3063 4835 3067
rect 4839 3063 4840 3067
rect 4834 3062 4840 3063
rect 4970 3067 4976 3068
rect 4970 3063 4971 3067
rect 4975 3063 4976 3067
rect 4970 3062 4976 3063
rect 5106 3067 5112 3068
rect 5106 3063 5107 3067
rect 5111 3063 5112 3067
rect 5106 3062 5112 3063
rect 5242 3067 5248 3068
rect 5242 3063 5243 3067
rect 5247 3063 5248 3067
rect 5242 3062 5248 3063
rect 5378 3067 5384 3068
rect 5378 3063 5379 3067
rect 5383 3063 5384 3067
rect 5378 3062 5384 3063
rect 5514 3067 5520 3068
rect 5514 3063 5515 3067
rect 5519 3063 5520 3067
rect 5662 3064 5663 3068
rect 5667 3064 5668 3068
rect 5662 3063 5668 3064
rect 5514 3062 5520 3063
rect 3799 3061 3803 3062
rect 111 3046 115 3047
rect 111 3041 115 3042
rect 319 3046 323 3047
rect 319 3041 323 3042
rect 327 3046 331 3047
rect 327 3041 331 3042
rect 487 3046 491 3047
rect 487 3041 491 3042
rect 647 3046 651 3047
rect 647 3041 651 3042
rect 655 3046 659 3047
rect 655 3041 659 3042
rect 807 3046 811 3047
rect 807 3041 811 3042
rect 839 3046 843 3047
rect 839 3041 843 3042
rect 959 3046 963 3047
rect 959 3041 963 3042
rect 1023 3046 1027 3047
rect 1023 3041 1027 3042
rect 1103 3046 1107 3047
rect 1103 3041 1107 3042
rect 1215 3046 1219 3047
rect 1215 3041 1219 3042
rect 1247 3046 1251 3047
rect 1247 3041 1251 3042
rect 1391 3046 1395 3047
rect 1391 3041 1395 3042
rect 1415 3046 1419 3047
rect 1415 3041 1419 3042
rect 1535 3046 1539 3047
rect 1535 3041 1539 3042
rect 1623 3046 1627 3047
rect 1623 3041 1627 3042
rect 1679 3046 1683 3047
rect 1679 3041 1683 3042
rect 1815 3046 1819 3047
rect 1815 3041 1819 3042
rect 1935 3046 1939 3047
rect 1935 3041 1939 3042
rect 112 3018 114 3041
rect 110 3017 116 3018
rect 328 3017 330 3041
rect 488 3017 490 3041
rect 648 3017 650 3041
rect 808 3017 810 3041
rect 960 3017 962 3041
rect 1104 3017 1106 3041
rect 1248 3017 1250 3041
rect 1392 3017 1394 3041
rect 1536 3017 1538 3041
rect 1680 3017 1682 3041
rect 1816 3017 1818 3041
rect 1936 3018 1938 3041
rect 1934 3017 1940 3018
rect 110 3013 111 3017
rect 115 3013 116 3017
rect 110 3012 116 3013
rect 326 3016 332 3017
rect 326 3012 327 3016
rect 331 3012 332 3016
rect 326 3011 332 3012
rect 486 3016 492 3017
rect 486 3012 487 3016
rect 491 3012 492 3016
rect 486 3011 492 3012
rect 646 3016 652 3017
rect 646 3012 647 3016
rect 651 3012 652 3016
rect 646 3011 652 3012
rect 806 3016 812 3017
rect 806 3012 807 3016
rect 811 3012 812 3016
rect 806 3011 812 3012
rect 958 3016 964 3017
rect 958 3012 959 3016
rect 963 3012 964 3016
rect 958 3011 964 3012
rect 1102 3016 1108 3017
rect 1102 3012 1103 3016
rect 1107 3012 1108 3016
rect 1102 3011 1108 3012
rect 1246 3016 1252 3017
rect 1246 3012 1247 3016
rect 1251 3012 1252 3016
rect 1246 3011 1252 3012
rect 1390 3016 1396 3017
rect 1390 3012 1391 3016
rect 1395 3012 1396 3016
rect 1390 3011 1396 3012
rect 1534 3016 1540 3017
rect 1534 3012 1535 3016
rect 1539 3012 1540 3016
rect 1534 3011 1540 3012
rect 1678 3016 1684 3017
rect 1678 3012 1679 3016
rect 1683 3012 1684 3016
rect 1678 3011 1684 3012
rect 1814 3016 1820 3017
rect 1814 3012 1815 3016
rect 1819 3012 1820 3016
rect 1934 3013 1935 3017
rect 1939 3013 1940 3017
rect 1934 3012 1940 3013
rect 1814 3011 1820 3012
rect 298 3001 304 3002
rect 110 3000 116 3001
rect 110 2996 111 3000
rect 115 2996 116 3000
rect 298 2997 299 3001
rect 303 2997 304 3001
rect 298 2996 304 2997
rect 458 3001 464 3002
rect 458 2997 459 3001
rect 463 2997 464 3001
rect 458 2996 464 2997
rect 618 3001 624 3002
rect 618 2997 619 3001
rect 623 2997 624 3001
rect 618 2996 624 2997
rect 778 3001 784 3002
rect 778 2997 779 3001
rect 783 2997 784 3001
rect 778 2996 784 2997
rect 930 3001 936 3002
rect 930 2997 931 3001
rect 935 2997 936 3001
rect 930 2996 936 2997
rect 1074 3001 1080 3002
rect 1074 2997 1075 3001
rect 1079 2997 1080 3001
rect 1074 2996 1080 2997
rect 1218 3001 1224 3002
rect 1218 2997 1219 3001
rect 1223 2997 1224 3001
rect 1218 2996 1224 2997
rect 1362 3001 1368 3002
rect 1362 2997 1363 3001
rect 1367 2997 1368 3001
rect 1362 2996 1368 2997
rect 1506 3001 1512 3002
rect 1506 2997 1507 3001
rect 1511 2997 1512 3001
rect 1506 2996 1512 2997
rect 1650 3001 1656 3002
rect 1650 2997 1651 3001
rect 1655 2997 1656 3001
rect 1650 2996 1656 2997
rect 1786 3001 1792 3002
rect 1976 3001 1978 3061
rect 1786 2997 1787 3001
rect 1791 2997 1792 3001
rect 1786 2996 1792 2997
rect 1934 3000 1940 3001
rect 1934 2996 1935 3000
rect 1939 2996 1940 3000
rect 110 2995 116 2996
rect 112 2935 114 2995
rect 300 2935 302 2996
rect 460 2935 462 2996
rect 620 2935 622 2996
rect 780 2935 782 2996
rect 932 2935 934 2996
rect 1076 2935 1078 2996
rect 1220 2935 1222 2996
rect 1364 2935 1366 2996
rect 1508 2935 1510 2996
rect 1652 2935 1654 2996
rect 1788 2935 1790 2996
rect 1934 2995 1940 2996
rect 1974 3000 1980 3001
rect 2812 3000 2814 3061
rect 3004 3000 3006 3061
rect 3204 3000 3206 3061
rect 3404 3000 3406 3061
rect 3604 3000 3606 3061
rect 3800 3001 3802 3061
rect 4726 3052 4732 3053
rect 3838 3051 3844 3052
rect 3838 3047 3839 3051
rect 3843 3047 3844 3051
rect 4726 3048 4727 3052
rect 4731 3048 4732 3052
rect 4726 3047 4732 3048
rect 4862 3052 4868 3053
rect 4862 3048 4863 3052
rect 4867 3048 4868 3052
rect 4862 3047 4868 3048
rect 4998 3052 5004 3053
rect 4998 3048 4999 3052
rect 5003 3048 5004 3052
rect 4998 3047 5004 3048
rect 5134 3052 5140 3053
rect 5134 3048 5135 3052
rect 5139 3048 5140 3052
rect 5134 3047 5140 3048
rect 5270 3052 5276 3053
rect 5270 3048 5271 3052
rect 5275 3048 5276 3052
rect 5270 3047 5276 3048
rect 5406 3052 5412 3053
rect 5406 3048 5407 3052
rect 5411 3048 5412 3052
rect 5406 3047 5412 3048
rect 5542 3052 5548 3053
rect 5542 3048 5543 3052
rect 5547 3048 5548 3052
rect 5542 3047 5548 3048
rect 5662 3051 5668 3052
rect 5662 3047 5663 3051
rect 5667 3047 5668 3051
rect 3838 3046 3844 3047
rect 3840 3023 3842 3046
rect 4728 3023 4730 3047
rect 4864 3023 4866 3047
rect 5000 3023 5002 3047
rect 5136 3023 5138 3047
rect 5272 3023 5274 3047
rect 5408 3023 5410 3047
rect 5544 3023 5546 3047
rect 5662 3046 5668 3047
rect 5664 3023 5666 3046
rect 3839 3022 3843 3023
rect 3839 3017 3843 3018
rect 4367 3022 4371 3023
rect 4367 3017 4371 3018
rect 4567 3022 4571 3023
rect 4567 3017 4571 3018
rect 4727 3022 4731 3023
rect 4727 3017 4731 3018
rect 4783 3022 4787 3023
rect 4783 3017 4787 3018
rect 4863 3022 4867 3023
rect 4863 3017 4867 3018
rect 4999 3022 5003 3023
rect 4999 3017 5003 3018
rect 5023 3022 5027 3023
rect 5023 3017 5027 3018
rect 5135 3022 5139 3023
rect 5135 3017 5139 3018
rect 5271 3022 5275 3023
rect 5271 3017 5275 3018
rect 5279 3022 5283 3023
rect 5279 3017 5283 3018
rect 5407 3022 5411 3023
rect 5407 3017 5411 3018
rect 5535 3022 5539 3023
rect 5535 3017 5539 3018
rect 5543 3022 5547 3023
rect 5543 3017 5547 3018
rect 5663 3022 5667 3023
rect 5663 3017 5667 3018
rect 3798 3000 3804 3001
rect 1974 2996 1975 3000
rect 1979 2996 1980 3000
rect 1974 2995 1980 2996
rect 2810 2999 2816 3000
rect 2810 2995 2811 2999
rect 2815 2995 2816 2999
rect 1936 2935 1938 2995
rect 2810 2994 2816 2995
rect 3002 2999 3008 3000
rect 3002 2995 3003 2999
rect 3007 2995 3008 2999
rect 3002 2994 3008 2995
rect 3202 2999 3208 3000
rect 3202 2995 3203 2999
rect 3207 2995 3208 2999
rect 3202 2994 3208 2995
rect 3402 2999 3408 3000
rect 3402 2995 3403 2999
rect 3407 2995 3408 2999
rect 3402 2994 3408 2995
rect 3602 2999 3608 3000
rect 3602 2995 3603 2999
rect 3607 2995 3608 2999
rect 3798 2996 3799 3000
rect 3803 2996 3804 3000
rect 3798 2995 3804 2996
rect 3602 2994 3608 2995
rect 3840 2994 3842 3017
rect 3838 2993 3844 2994
rect 4368 2993 4370 3017
rect 4568 2993 4570 3017
rect 4784 2993 4786 3017
rect 5024 2993 5026 3017
rect 5280 2993 5282 3017
rect 5536 2993 5538 3017
rect 5664 2994 5666 3017
rect 5662 2993 5668 2994
rect 3838 2989 3839 2993
rect 3843 2989 3844 2993
rect 3838 2988 3844 2989
rect 4366 2992 4372 2993
rect 4366 2988 4367 2992
rect 4371 2988 4372 2992
rect 4366 2987 4372 2988
rect 4566 2992 4572 2993
rect 4566 2988 4567 2992
rect 4571 2988 4572 2992
rect 4566 2987 4572 2988
rect 4782 2992 4788 2993
rect 4782 2988 4783 2992
rect 4787 2988 4788 2992
rect 4782 2987 4788 2988
rect 5022 2992 5028 2993
rect 5022 2988 5023 2992
rect 5027 2988 5028 2992
rect 5022 2987 5028 2988
rect 5278 2992 5284 2993
rect 5278 2988 5279 2992
rect 5283 2988 5284 2992
rect 5278 2987 5284 2988
rect 5534 2992 5540 2993
rect 5534 2988 5535 2992
rect 5539 2988 5540 2992
rect 5662 2989 5663 2993
rect 5667 2989 5668 2993
rect 5662 2988 5668 2989
rect 5534 2987 5540 2988
rect 2838 2984 2844 2985
rect 1974 2983 1980 2984
rect 1974 2979 1975 2983
rect 1979 2979 1980 2983
rect 2838 2980 2839 2984
rect 2843 2980 2844 2984
rect 2838 2979 2844 2980
rect 3030 2984 3036 2985
rect 3030 2980 3031 2984
rect 3035 2980 3036 2984
rect 3030 2979 3036 2980
rect 3230 2984 3236 2985
rect 3230 2980 3231 2984
rect 3235 2980 3236 2984
rect 3230 2979 3236 2980
rect 3430 2984 3436 2985
rect 3430 2980 3431 2984
rect 3435 2980 3436 2984
rect 3430 2979 3436 2980
rect 3630 2984 3636 2985
rect 3630 2980 3631 2984
rect 3635 2980 3636 2984
rect 3630 2979 3636 2980
rect 3798 2983 3804 2984
rect 3798 2979 3799 2983
rect 3803 2979 3804 2983
rect 1974 2978 1980 2979
rect 1976 2947 1978 2978
rect 2840 2947 2842 2979
rect 3032 2947 3034 2979
rect 3232 2947 3234 2979
rect 3432 2947 3434 2979
rect 3632 2947 3634 2979
rect 3798 2978 3804 2979
rect 3800 2947 3802 2978
rect 4338 2977 4344 2978
rect 3838 2976 3844 2977
rect 3838 2972 3839 2976
rect 3843 2972 3844 2976
rect 4338 2973 4339 2977
rect 4343 2973 4344 2977
rect 4338 2972 4344 2973
rect 4538 2977 4544 2978
rect 4538 2973 4539 2977
rect 4543 2973 4544 2977
rect 4538 2972 4544 2973
rect 4754 2977 4760 2978
rect 4754 2973 4755 2977
rect 4759 2973 4760 2977
rect 4754 2972 4760 2973
rect 4994 2977 5000 2978
rect 4994 2973 4995 2977
rect 4999 2973 5000 2977
rect 4994 2972 5000 2973
rect 5250 2977 5256 2978
rect 5250 2973 5251 2977
rect 5255 2973 5256 2977
rect 5250 2972 5256 2973
rect 5506 2977 5512 2978
rect 5506 2973 5507 2977
rect 5511 2973 5512 2977
rect 5506 2972 5512 2973
rect 5662 2976 5668 2977
rect 5662 2972 5663 2976
rect 5667 2972 5668 2976
rect 3838 2971 3844 2972
rect 1975 2946 1979 2947
rect 1975 2941 1979 2942
rect 2839 2946 2843 2947
rect 2839 2941 2843 2942
rect 2847 2946 2851 2947
rect 2847 2941 2851 2942
rect 2983 2946 2987 2947
rect 2983 2941 2987 2942
rect 3031 2946 3035 2947
rect 3031 2941 3035 2942
rect 3119 2946 3123 2947
rect 3119 2941 3123 2942
rect 3231 2946 3235 2947
rect 3231 2941 3235 2942
rect 3255 2946 3259 2947
rect 3255 2941 3259 2942
rect 3391 2946 3395 2947
rect 3391 2941 3395 2942
rect 3431 2946 3435 2947
rect 3431 2941 3435 2942
rect 3527 2946 3531 2947
rect 3527 2941 3531 2942
rect 3631 2946 3635 2947
rect 3631 2941 3635 2942
rect 3671 2946 3675 2947
rect 3671 2941 3675 2942
rect 3799 2946 3803 2947
rect 3799 2941 3803 2942
rect 111 2934 115 2935
rect 111 2929 115 2930
rect 155 2934 159 2935
rect 155 2929 159 2930
rect 299 2934 303 2935
rect 299 2929 303 2930
rect 379 2934 383 2935
rect 379 2929 383 2930
rect 459 2934 463 2935
rect 459 2929 463 2930
rect 595 2934 599 2935
rect 595 2929 599 2930
rect 619 2934 623 2935
rect 619 2929 623 2930
rect 779 2934 783 2935
rect 779 2929 783 2930
rect 811 2934 815 2935
rect 811 2929 815 2930
rect 931 2934 935 2935
rect 931 2929 935 2930
rect 1019 2934 1023 2935
rect 1019 2929 1023 2930
rect 1075 2934 1079 2935
rect 1075 2929 1079 2930
rect 1219 2934 1223 2935
rect 1219 2929 1223 2930
rect 1363 2934 1367 2935
rect 1363 2929 1367 2930
rect 1411 2934 1415 2935
rect 1411 2929 1415 2930
rect 1507 2934 1511 2935
rect 1507 2929 1511 2930
rect 1611 2934 1615 2935
rect 1611 2929 1615 2930
rect 1651 2934 1655 2935
rect 1651 2929 1655 2930
rect 1787 2934 1791 2935
rect 1787 2929 1791 2930
rect 1935 2934 1939 2935
rect 1935 2929 1939 2930
rect 112 2869 114 2929
rect 110 2868 116 2869
rect 156 2868 158 2929
rect 380 2868 382 2929
rect 596 2868 598 2929
rect 812 2868 814 2929
rect 1020 2868 1022 2929
rect 1220 2868 1222 2929
rect 1412 2868 1414 2929
rect 1612 2868 1614 2929
rect 1788 2868 1790 2929
rect 1936 2869 1938 2929
rect 1976 2918 1978 2941
rect 1974 2917 1980 2918
rect 2848 2917 2850 2941
rect 2984 2917 2986 2941
rect 3120 2917 3122 2941
rect 3256 2917 3258 2941
rect 3392 2917 3394 2941
rect 3528 2917 3530 2941
rect 3672 2917 3674 2941
rect 3800 2918 3802 2941
rect 3798 2917 3804 2918
rect 1974 2913 1975 2917
rect 1979 2913 1980 2917
rect 1974 2912 1980 2913
rect 2846 2916 2852 2917
rect 2846 2912 2847 2916
rect 2851 2912 2852 2916
rect 2846 2911 2852 2912
rect 2982 2916 2988 2917
rect 2982 2912 2983 2916
rect 2987 2912 2988 2916
rect 2982 2911 2988 2912
rect 3118 2916 3124 2917
rect 3118 2912 3119 2916
rect 3123 2912 3124 2916
rect 3118 2911 3124 2912
rect 3254 2916 3260 2917
rect 3254 2912 3255 2916
rect 3259 2912 3260 2916
rect 3254 2911 3260 2912
rect 3390 2916 3396 2917
rect 3390 2912 3391 2916
rect 3395 2912 3396 2916
rect 3390 2911 3396 2912
rect 3526 2916 3532 2917
rect 3526 2912 3527 2916
rect 3531 2912 3532 2916
rect 3526 2911 3532 2912
rect 3670 2916 3676 2917
rect 3670 2912 3671 2916
rect 3675 2912 3676 2916
rect 3798 2913 3799 2917
rect 3803 2913 3804 2917
rect 3798 2912 3804 2913
rect 3670 2911 3676 2912
rect 3840 2911 3842 2971
rect 4340 2911 4342 2972
rect 4540 2911 4542 2972
rect 4756 2911 4758 2972
rect 4996 2911 4998 2972
rect 5252 2911 5254 2972
rect 5508 2911 5510 2972
rect 5662 2971 5668 2972
rect 5664 2911 5666 2971
rect 3839 2910 3843 2911
rect 3839 2905 3843 2906
rect 4035 2910 4039 2911
rect 4035 2905 4039 2906
rect 4315 2910 4319 2911
rect 4315 2905 4319 2906
rect 4339 2910 4343 2911
rect 4339 2905 4343 2906
rect 4539 2910 4543 2911
rect 4539 2905 4543 2906
rect 4603 2910 4607 2911
rect 4603 2905 4607 2906
rect 4755 2910 4759 2911
rect 4755 2905 4759 2906
rect 4907 2910 4911 2911
rect 4907 2905 4911 2906
rect 4995 2910 4999 2911
rect 4995 2905 4999 2906
rect 5219 2910 5223 2911
rect 5219 2905 5223 2906
rect 5251 2910 5255 2911
rect 5251 2905 5255 2906
rect 5507 2910 5511 2911
rect 5507 2905 5511 2906
rect 5515 2910 5519 2911
rect 5515 2905 5519 2906
rect 5663 2910 5667 2911
rect 5663 2905 5667 2906
rect 2818 2901 2824 2902
rect 1974 2900 1980 2901
rect 1974 2896 1975 2900
rect 1979 2896 1980 2900
rect 2818 2897 2819 2901
rect 2823 2897 2824 2901
rect 2818 2896 2824 2897
rect 2954 2901 2960 2902
rect 2954 2897 2955 2901
rect 2959 2897 2960 2901
rect 2954 2896 2960 2897
rect 3090 2901 3096 2902
rect 3090 2897 3091 2901
rect 3095 2897 3096 2901
rect 3090 2896 3096 2897
rect 3226 2901 3232 2902
rect 3226 2897 3227 2901
rect 3231 2897 3232 2901
rect 3226 2896 3232 2897
rect 3362 2901 3368 2902
rect 3362 2897 3363 2901
rect 3367 2897 3368 2901
rect 3362 2896 3368 2897
rect 3498 2901 3504 2902
rect 3498 2897 3499 2901
rect 3503 2897 3504 2901
rect 3498 2896 3504 2897
rect 3642 2901 3648 2902
rect 3642 2897 3643 2901
rect 3647 2897 3648 2901
rect 3642 2896 3648 2897
rect 3798 2900 3804 2901
rect 3798 2896 3799 2900
rect 3803 2896 3804 2900
rect 1974 2895 1980 2896
rect 1934 2868 1940 2869
rect 110 2864 111 2868
rect 115 2864 116 2868
rect 110 2863 116 2864
rect 154 2867 160 2868
rect 154 2863 155 2867
rect 159 2863 160 2867
rect 154 2862 160 2863
rect 378 2867 384 2868
rect 378 2863 379 2867
rect 383 2863 384 2867
rect 378 2862 384 2863
rect 594 2867 600 2868
rect 594 2863 595 2867
rect 599 2863 600 2867
rect 594 2862 600 2863
rect 810 2867 816 2868
rect 810 2863 811 2867
rect 815 2863 816 2867
rect 810 2862 816 2863
rect 1018 2867 1024 2868
rect 1018 2863 1019 2867
rect 1023 2863 1024 2867
rect 1018 2862 1024 2863
rect 1218 2867 1224 2868
rect 1218 2863 1219 2867
rect 1223 2863 1224 2867
rect 1218 2862 1224 2863
rect 1410 2867 1416 2868
rect 1410 2863 1411 2867
rect 1415 2863 1416 2867
rect 1410 2862 1416 2863
rect 1610 2867 1616 2868
rect 1610 2863 1611 2867
rect 1615 2863 1616 2867
rect 1610 2862 1616 2863
rect 1786 2867 1792 2868
rect 1786 2863 1787 2867
rect 1791 2863 1792 2867
rect 1934 2864 1935 2868
rect 1939 2864 1940 2868
rect 1934 2863 1940 2864
rect 1786 2862 1792 2863
rect 182 2852 188 2853
rect 110 2851 116 2852
rect 110 2847 111 2851
rect 115 2847 116 2851
rect 182 2848 183 2852
rect 187 2848 188 2852
rect 182 2847 188 2848
rect 406 2852 412 2853
rect 406 2848 407 2852
rect 411 2848 412 2852
rect 406 2847 412 2848
rect 622 2852 628 2853
rect 622 2848 623 2852
rect 627 2848 628 2852
rect 622 2847 628 2848
rect 838 2852 844 2853
rect 838 2848 839 2852
rect 843 2848 844 2852
rect 838 2847 844 2848
rect 1046 2852 1052 2853
rect 1046 2848 1047 2852
rect 1051 2848 1052 2852
rect 1046 2847 1052 2848
rect 1246 2852 1252 2853
rect 1246 2848 1247 2852
rect 1251 2848 1252 2852
rect 1246 2847 1252 2848
rect 1438 2852 1444 2853
rect 1438 2848 1439 2852
rect 1443 2848 1444 2852
rect 1438 2847 1444 2848
rect 1638 2852 1644 2853
rect 1638 2848 1639 2852
rect 1643 2848 1644 2852
rect 1638 2847 1644 2848
rect 1814 2852 1820 2853
rect 1814 2848 1815 2852
rect 1819 2848 1820 2852
rect 1814 2847 1820 2848
rect 1934 2851 1940 2852
rect 1934 2847 1935 2851
rect 1939 2847 1940 2851
rect 110 2846 116 2847
rect 112 2791 114 2846
rect 184 2791 186 2847
rect 408 2791 410 2847
rect 624 2791 626 2847
rect 840 2791 842 2847
rect 1048 2791 1050 2847
rect 1248 2791 1250 2847
rect 1440 2791 1442 2847
rect 1640 2791 1642 2847
rect 1816 2791 1818 2847
rect 1934 2846 1940 2847
rect 1936 2791 1938 2846
rect 1976 2835 1978 2895
rect 2820 2835 2822 2896
rect 2956 2835 2958 2896
rect 3092 2835 3094 2896
rect 3228 2835 3230 2896
rect 3364 2835 3366 2896
rect 3500 2835 3502 2896
rect 3644 2835 3646 2896
rect 3798 2895 3804 2896
rect 3800 2835 3802 2895
rect 3840 2845 3842 2905
rect 3838 2844 3844 2845
rect 4036 2844 4038 2905
rect 4316 2844 4318 2905
rect 4604 2844 4606 2905
rect 4908 2844 4910 2905
rect 5220 2844 5222 2905
rect 5516 2844 5518 2905
rect 5664 2845 5666 2905
rect 5662 2844 5668 2845
rect 3838 2840 3839 2844
rect 3843 2840 3844 2844
rect 3838 2839 3844 2840
rect 4034 2843 4040 2844
rect 4034 2839 4035 2843
rect 4039 2839 4040 2843
rect 4034 2838 4040 2839
rect 4314 2843 4320 2844
rect 4314 2839 4315 2843
rect 4319 2839 4320 2843
rect 4314 2838 4320 2839
rect 4602 2843 4608 2844
rect 4602 2839 4603 2843
rect 4607 2839 4608 2843
rect 4602 2838 4608 2839
rect 4906 2843 4912 2844
rect 4906 2839 4907 2843
rect 4911 2839 4912 2843
rect 4906 2838 4912 2839
rect 5218 2843 5224 2844
rect 5218 2839 5219 2843
rect 5223 2839 5224 2843
rect 5218 2838 5224 2839
rect 5514 2843 5520 2844
rect 5514 2839 5515 2843
rect 5519 2839 5520 2843
rect 5662 2840 5663 2844
rect 5667 2840 5668 2844
rect 5662 2839 5668 2840
rect 5514 2838 5520 2839
rect 1975 2834 1979 2835
rect 1975 2829 1979 2830
rect 2011 2834 2015 2835
rect 2011 2829 2015 2830
rect 2251 2834 2255 2835
rect 2251 2829 2255 2830
rect 2491 2834 2495 2835
rect 2491 2829 2495 2830
rect 2731 2834 2735 2835
rect 2731 2829 2735 2830
rect 2819 2834 2823 2835
rect 2819 2829 2823 2830
rect 2955 2834 2959 2835
rect 2955 2829 2959 2830
rect 2971 2834 2975 2835
rect 2971 2829 2975 2830
rect 3091 2834 3095 2835
rect 3091 2829 3095 2830
rect 3227 2834 3231 2835
rect 3227 2829 3231 2830
rect 3363 2834 3367 2835
rect 3363 2829 3367 2830
rect 3499 2834 3503 2835
rect 3499 2829 3503 2830
rect 3643 2834 3647 2835
rect 3643 2829 3647 2830
rect 3799 2834 3803 2835
rect 3799 2829 3803 2830
rect 111 2790 115 2791
rect 111 2785 115 2786
rect 183 2790 187 2791
rect 183 2785 187 2786
rect 287 2790 291 2791
rect 287 2785 291 2786
rect 407 2790 411 2791
rect 407 2785 411 2786
rect 423 2790 427 2791
rect 423 2785 427 2786
rect 559 2790 563 2791
rect 559 2785 563 2786
rect 623 2790 627 2791
rect 623 2785 627 2786
rect 695 2790 699 2791
rect 695 2785 699 2786
rect 831 2790 835 2791
rect 831 2785 835 2786
rect 839 2790 843 2791
rect 839 2785 843 2786
rect 1047 2790 1051 2791
rect 1047 2785 1051 2786
rect 1247 2790 1251 2791
rect 1247 2785 1251 2786
rect 1439 2790 1443 2791
rect 1439 2785 1443 2786
rect 1639 2790 1643 2791
rect 1639 2785 1643 2786
rect 1815 2790 1819 2791
rect 1815 2785 1819 2786
rect 1935 2790 1939 2791
rect 1935 2785 1939 2786
rect 112 2762 114 2785
rect 110 2761 116 2762
rect 288 2761 290 2785
rect 424 2761 426 2785
rect 560 2761 562 2785
rect 696 2761 698 2785
rect 832 2761 834 2785
rect 1936 2762 1938 2785
rect 1976 2769 1978 2829
rect 1974 2768 1980 2769
rect 2012 2768 2014 2829
rect 2252 2768 2254 2829
rect 2492 2768 2494 2829
rect 2732 2768 2734 2829
rect 2972 2768 2974 2829
rect 3800 2769 3802 2829
rect 4062 2828 4068 2829
rect 3838 2827 3844 2828
rect 3838 2823 3839 2827
rect 3843 2823 3844 2827
rect 4062 2824 4063 2828
rect 4067 2824 4068 2828
rect 4062 2823 4068 2824
rect 4342 2828 4348 2829
rect 4342 2824 4343 2828
rect 4347 2824 4348 2828
rect 4342 2823 4348 2824
rect 4630 2828 4636 2829
rect 4630 2824 4631 2828
rect 4635 2824 4636 2828
rect 4630 2823 4636 2824
rect 4934 2828 4940 2829
rect 4934 2824 4935 2828
rect 4939 2824 4940 2828
rect 4934 2823 4940 2824
rect 5246 2828 5252 2829
rect 5246 2824 5247 2828
rect 5251 2824 5252 2828
rect 5246 2823 5252 2824
rect 5542 2828 5548 2829
rect 5542 2824 5543 2828
rect 5547 2824 5548 2828
rect 5542 2823 5548 2824
rect 5662 2827 5668 2828
rect 5662 2823 5663 2827
rect 5667 2823 5668 2827
rect 3838 2822 3844 2823
rect 3840 2791 3842 2822
rect 4064 2791 4066 2823
rect 4344 2791 4346 2823
rect 4632 2791 4634 2823
rect 4936 2791 4938 2823
rect 5248 2791 5250 2823
rect 5544 2791 5546 2823
rect 5662 2822 5668 2823
rect 5664 2791 5666 2822
rect 3839 2790 3843 2791
rect 3839 2785 3843 2786
rect 3967 2790 3971 2791
rect 3967 2785 3971 2786
rect 4063 2790 4067 2791
rect 4063 2785 4067 2786
rect 4255 2790 4259 2791
rect 4255 2785 4259 2786
rect 4343 2790 4347 2791
rect 4343 2785 4347 2786
rect 4567 2790 4571 2791
rect 4567 2785 4571 2786
rect 4631 2790 4635 2791
rect 4631 2785 4635 2786
rect 4895 2790 4899 2791
rect 4895 2785 4899 2786
rect 4935 2790 4939 2791
rect 4935 2785 4939 2786
rect 5231 2790 5235 2791
rect 5231 2785 5235 2786
rect 5247 2790 5251 2791
rect 5247 2785 5251 2786
rect 5543 2790 5547 2791
rect 5543 2785 5547 2786
rect 5663 2790 5667 2791
rect 5663 2785 5667 2786
rect 3798 2768 3804 2769
rect 1974 2764 1975 2768
rect 1979 2764 1980 2768
rect 1974 2763 1980 2764
rect 2010 2767 2016 2768
rect 2010 2763 2011 2767
rect 2015 2763 2016 2767
rect 2010 2762 2016 2763
rect 2250 2767 2256 2768
rect 2250 2763 2251 2767
rect 2255 2763 2256 2767
rect 2250 2762 2256 2763
rect 2490 2767 2496 2768
rect 2490 2763 2491 2767
rect 2495 2763 2496 2767
rect 2490 2762 2496 2763
rect 2730 2767 2736 2768
rect 2730 2763 2731 2767
rect 2735 2763 2736 2767
rect 2730 2762 2736 2763
rect 2970 2767 2976 2768
rect 2970 2763 2971 2767
rect 2975 2763 2976 2767
rect 3798 2764 3799 2768
rect 3803 2764 3804 2768
rect 3798 2763 3804 2764
rect 2970 2762 2976 2763
rect 3840 2762 3842 2785
rect 1934 2761 1940 2762
rect 110 2757 111 2761
rect 115 2757 116 2761
rect 110 2756 116 2757
rect 286 2760 292 2761
rect 286 2756 287 2760
rect 291 2756 292 2760
rect 286 2755 292 2756
rect 422 2760 428 2761
rect 422 2756 423 2760
rect 427 2756 428 2760
rect 422 2755 428 2756
rect 558 2760 564 2761
rect 558 2756 559 2760
rect 563 2756 564 2760
rect 558 2755 564 2756
rect 694 2760 700 2761
rect 694 2756 695 2760
rect 699 2756 700 2760
rect 694 2755 700 2756
rect 830 2760 836 2761
rect 830 2756 831 2760
rect 835 2756 836 2760
rect 1934 2757 1935 2761
rect 1939 2757 1940 2761
rect 1934 2756 1940 2757
rect 3838 2761 3844 2762
rect 3968 2761 3970 2785
rect 4256 2761 4258 2785
rect 4568 2761 4570 2785
rect 4896 2761 4898 2785
rect 5232 2761 5234 2785
rect 5544 2761 5546 2785
rect 5664 2762 5666 2785
rect 5662 2761 5668 2762
rect 3838 2757 3839 2761
rect 3843 2757 3844 2761
rect 3838 2756 3844 2757
rect 3966 2760 3972 2761
rect 3966 2756 3967 2760
rect 3971 2756 3972 2760
rect 830 2755 836 2756
rect 3966 2755 3972 2756
rect 4254 2760 4260 2761
rect 4254 2756 4255 2760
rect 4259 2756 4260 2760
rect 4254 2755 4260 2756
rect 4566 2760 4572 2761
rect 4566 2756 4567 2760
rect 4571 2756 4572 2760
rect 4566 2755 4572 2756
rect 4894 2760 4900 2761
rect 4894 2756 4895 2760
rect 4899 2756 4900 2760
rect 4894 2755 4900 2756
rect 5230 2760 5236 2761
rect 5230 2756 5231 2760
rect 5235 2756 5236 2760
rect 5230 2755 5236 2756
rect 5542 2760 5548 2761
rect 5542 2756 5543 2760
rect 5547 2756 5548 2760
rect 5662 2757 5663 2761
rect 5667 2757 5668 2761
rect 5662 2756 5668 2757
rect 5542 2755 5548 2756
rect 2038 2752 2044 2753
rect 1974 2751 1980 2752
rect 1974 2747 1975 2751
rect 1979 2747 1980 2751
rect 2038 2748 2039 2752
rect 2043 2748 2044 2752
rect 2038 2747 2044 2748
rect 2278 2752 2284 2753
rect 2278 2748 2279 2752
rect 2283 2748 2284 2752
rect 2278 2747 2284 2748
rect 2518 2752 2524 2753
rect 2518 2748 2519 2752
rect 2523 2748 2524 2752
rect 2518 2747 2524 2748
rect 2758 2752 2764 2753
rect 2758 2748 2759 2752
rect 2763 2748 2764 2752
rect 2758 2747 2764 2748
rect 2998 2752 3004 2753
rect 2998 2748 2999 2752
rect 3003 2748 3004 2752
rect 2998 2747 3004 2748
rect 3798 2751 3804 2752
rect 3798 2747 3799 2751
rect 3803 2747 3804 2751
rect 1974 2746 1980 2747
rect 258 2745 264 2746
rect 110 2744 116 2745
rect 110 2740 111 2744
rect 115 2740 116 2744
rect 258 2741 259 2745
rect 263 2741 264 2745
rect 258 2740 264 2741
rect 394 2745 400 2746
rect 394 2741 395 2745
rect 399 2741 400 2745
rect 394 2740 400 2741
rect 530 2745 536 2746
rect 530 2741 531 2745
rect 535 2741 536 2745
rect 530 2740 536 2741
rect 666 2745 672 2746
rect 666 2741 667 2745
rect 671 2741 672 2745
rect 666 2740 672 2741
rect 802 2745 808 2746
rect 802 2741 803 2745
rect 807 2741 808 2745
rect 802 2740 808 2741
rect 1934 2744 1940 2745
rect 1934 2740 1935 2744
rect 1939 2740 1940 2744
rect 110 2739 116 2740
rect 112 2659 114 2739
rect 260 2659 262 2740
rect 396 2659 398 2740
rect 532 2659 534 2740
rect 668 2659 670 2740
rect 804 2659 806 2740
rect 1934 2739 1940 2740
rect 1936 2659 1938 2739
rect 1976 2723 1978 2746
rect 2040 2723 2042 2747
rect 2280 2723 2282 2747
rect 2520 2723 2522 2747
rect 2760 2723 2762 2747
rect 3000 2723 3002 2747
rect 3798 2746 3804 2747
rect 3800 2723 3802 2746
rect 3938 2745 3944 2746
rect 3838 2744 3844 2745
rect 3838 2740 3839 2744
rect 3843 2740 3844 2744
rect 3938 2741 3939 2745
rect 3943 2741 3944 2745
rect 3938 2740 3944 2741
rect 4226 2745 4232 2746
rect 4226 2741 4227 2745
rect 4231 2741 4232 2745
rect 4226 2740 4232 2741
rect 4538 2745 4544 2746
rect 4538 2741 4539 2745
rect 4543 2741 4544 2745
rect 4538 2740 4544 2741
rect 4866 2745 4872 2746
rect 4866 2741 4867 2745
rect 4871 2741 4872 2745
rect 4866 2740 4872 2741
rect 5202 2745 5208 2746
rect 5202 2741 5203 2745
rect 5207 2741 5208 2745
rect 5202 2740 5208 2741
rect 5514 2745 5520 2746
rect 5514 2741 5515 2745
rect 5519 2741 5520 2745
rect 5514 2740 5520 2741
rect 5662 2744 5668 2745
rect 5662 2740 5663 2744
rect 5667 2740 5668 2744
rect 3838 2739 3844 2740
rect 1975 2722 1979 2723
rect 1975 2717 1979 2718
rect 2023 2722 2027 2723
rect 2023 2717 2027 2718
rect 2039 2722 2043 2723
rect 2039 2717 2043 2718
rect 2159 2722 2163 2723
rect 2159 2717 2163 2718
rect 2279 2722 2283 2723
rect 2279 2717 2283 2718
rect 2295 2722 2299 2723
rect 2295 2717 2299 2718
rect 2431 2722 2435 2723
rect 2431 2717 2435 2718
rect 2519 2722 2523 2723
rect 2519 2717 2523 2718
rect 2567 2722 2571 2723
rect 2567 2717 2571 2718
rect 2703 2722 2707 2723
rect 2703 2717 2707 2718
rect 2759 2722 2763 2723
rect 2759 2717 2763 2718
rect 2839 2722 2843 2723
rect 2839 2717 2843 2718
rect 2975 2722 2979 2723
rect 2975 2717 2979 2718
rect 2999 2722 3003 2723
rect 2999 2717 3003 2718
rect 3111 2722 3115 2723
rect 3111 2717 3115 2718
rect 3247 2722 3251 2723
rect 3247 2717 3251 2718
rect 3383 2722 3387 2723
rect 3383 2717 3387 2718
rect 3799 2722 3803 2723
rect 3799 2717 3803 2718
rect 1976 2694 1978 2717
rect 1974 2693 1980 2694
rect 2024 2693 2026 2717
rect 2160 2693 2162 2717
rect 2296 2693 2298 2717
rect 2432 2693 2434 2717
rect 2568 2693 2570 2717
rect 2704 2693 2706 2717
rect 2840 2693 2842 2717
rect 2976 2693 2978 2717
rect 3112 2693 3114 2717
rect 3248 2693 3250 2717
rect 3384 2693 3386 2717
rect 3800 2694 3802 2717
rect 3798 2693 3804 2694
rect 1974 2689 1975 2693
rect 1979 2689 1980 2693
rect 1974 2688 1980 2689
rect 2022 2692 2028 2693
rect 2022 2688 2023 2692
rect 2027 2688 2028 2692
rect 2022 2687 2028 2688
rect 2158 2692 2164 2693
rect 2158 2688 2159 2692
rect 2163 2688 2164 2692
rect 2158 2687 2164 2688
rect 2294 2692 2300 2693
rect 2294 2688 2295 2692
rect 2299 2688 2300 2692
rect 2294 2687 2300 2688
rect 2430 2692 2436 2693
rect 2430 2688 2431 2692
rect 2435 2688 2436 2692
rect 2430 2687 2436 2688
rect 2566 2692 2572 2693
rect 2566 2688 2567 2692
rect 2571 2688 2572 2692
rect 2566 2687 2572 2688
rect 2702 2692 2708 2693
rect 2702 2688 2703 2692
rect 2707 2688 2708 2692
rect 2702 2687 2708 2688
rect 2838 2692 2844 2693
rect 2838 2688 2839 2692
rect 2843 2688 2844 2692
rect 2838 2687 2844 2688
rect 2974 2692 2980 2693
rect 2974 2688 2975 2692
rect 2979 2688 2980 2692
rect 2974 2687 2980 2688
rect 3110 2692 3116 2693
rect 3110 2688 3111 2692
rect 3115 2688 3116 2692
rect 3110 2687 3116 2688
rect 3246 2692 3252 2693
rect 3246 2688 3247 2692
rect 3251 2688 3252 2692
rect 3246 2687 3252 2688
rect 3382 2692 3388 2693
rect 3382 2688 3383 2692
rect 3387 2688 3388 2692
rect 3798 2689 3799 2693
rect 3803 2689 3804 2693
rect 3798 2688 3804 2689
rect 3382 2687 3388 2688
rect 1994 2677 2000 2678
rect 1974 2676 1980 2677
rect 1974 2672 1975 2676
rect 1979 2672 1980 2676
rect 1994 2673 1995 2677
rect 1999 2673 2000 2677
rect 1994 2672 2000 2673
rect 2130 2677 2136 2678
rect 2130 2673 2131 2677
rect 2135 2673 2136 2677
rect 2130 2672 2136 2673
rect 2266 2677 2272 2678
rect 2266 2673 2267 2677
rect 2271 2673 2272 2677
rect 2266 2672 2272 2673
rect 2402 2677 2408 2678
rect 2402 2673 2403 2677
rect 2407 2673 2408 2677
rect 2402 2672 2408 2673
rect 2538 2677 2544 2678
rect 2538 2673 2539 2677
rect 2543 2673 2544 2677
rect 2538 2672 2544 2673
rect 2674 2677 2680 2678
rect 2674 2673 2675 2677
rect 2679 2673 2680 2677
rect 2674 2672 2680 2673
rect 2810 2677 2816 2678
rect 2810 2673 2811 2677
rect 2815 2673 2816 2677
rect 2810 2672 2816 2673
rect 2946 2677 2952 2678
rect 2946 2673 2947 2677
rect 2951 2673 2952 2677
rect 2946 2672 2952 2673
rect 3082 2677 3088 2678
rect 3082 2673 3083 2677
rect 3087 2673 3088 2677
rect 3082 2672 3088 2673
rect 3218 2677 3224 2678
rect 3218 2673 3219 2677
rect 3223 2673 3224 2677
rect 3218 2672 3224 2673
rect 3354 2677 3360 2678
rect 3354 2673 3355 2677
rect 3359 2673 3360 2677
rect 3354 2672 3360 2673
rect 3798 2676 3804 2677
rect 3798 2672 3799 2676
rect 3803 2672 3804 2676
rect 3840 2675 3842 2739
rect 3940 2675 3942 2740
rect 4228 2675 4230 2740
rect 4540 2675 4542 2740
rect 4868 2675 4870 2740
rect 5204 2675 5206 2740
rect 5516 2675 5518 2740
rect 5662 2739 5668 2740
rect 5664 2675 5666 2739
rect 1974 2671 1980 2672
rect 111 2658 115 2659
rect 111 2653 115 2654
rect 259 2658 263 2659
rect 259 2653 263 2654
rect 395 2658 399 2659
rect 395 2653 399 2654
rect 531 2658 535 2659
rect 531 2653 535 2654
rect 539 2658 543 2659
rect 539 2653 543 2654
rect 667 2658 671 2659
rect 667 2653 671 2654
rect 699 2658 703 2659
rect 699 2653 703 2654
rect 803 2658 807 2659
rect 803 2653 807 2654
rect 883 2658 887 2659
rect 883 2653 887 2654
rect 1091 2658 1095 2659
rect 1091 2653 1095 2654
rect 1323 2658 1327 2659
rect 1323 2653 1327 2654
rect 1563 2658 1567 2659
rect 1563 2653 1567 2654
rect 1787 2658 1791 2659
rect 1787 2653 1791 2654
rect 1935 2658 1939 2659
rect 1935 2653 1939 2654
rect 112 2593 114 2653
rect 110 2592 116 2593
rect 540 2592 542 2653
rect 700 2592 702 2653
rect 884 2592 886 2653
rect 1092 2592 1094 2653
rect 1324 2592 1326 2653
rect 1564 2592 1566 2653
rect 1788 2592 1790 2653
rect 1936 2593 1938 2653
rect 1976 2611 1978 2671
rect 1996 2611 1998 2672
rect 2132 2611 2134 2672
rect 2268 2611 2270 2672
rect 2404 2611 2406 2672
rect 2540 2611 2542 2672
rect 2676 2611 2678 2672
rect 2812 2611 2814 2672
rect 2948 2611 2950 2672
rect 3084 2611 3086 2672
rect 3220 2611 3222 2672
rect 3356 2611 3358 2672
rect 3798 2671 3804 2672
rect 3839 2674 3843 2675
rect 3800 2611 3802 2671
rect 3839 2669 3843 2670
rect 3939 2674 3943 2675
rect 3939 2669 3943 2670
rect 4027 2674 4031 2675
rect 4027 2669 4031 2670
rect 4227 2674 4231 2675
rect 4227 2669 4231 2670
rect 4275 2674 4279 2675
rect 4275 2669 4279 2670
rect 4539 2674 4543 2675
rect 4539 2669 4543 2670
rect 4555 2674 4559 2675
rect 4555 2669 4559 2670
rect 4867 2674 4871 2675
rect 4867 2669 4871 2670
rect 5203 2674 5207 2675
rect 5203 2669 5207 2670
rect 5515 2674 5519 2675
rect 5515 2669 5519 2670
rect 5663 2674 5667 2675
rect 5663 2669 5667 2670
rect 1975 2610 1979 2611
rect 1975 2605 1979 2606
rect 1995 2610 1999 2611
rect 1995 2605 1999 2606
rect 2131 2610 2135 2611
rect 2131 2605 2135 2606
rect 2203 2610 2207 2611
rect 2203 2605 2207 2606
rect 2267 2610 2271 2611
rect 2267 2605 2271 2606
rect 2403 2610 2407 2611
rect 2403 2605 2407 2606
rect 2419 2610 2423 2611
rect 2419 2605 2423 2606
rect 2539 2610 2543 2611
rect 2539 2605 2543 2606
rect 2627 2610 2631 2611
rect 2627 2605 2631 2606
rect 2675 2610 2679 2611
rect 2675 2605 2679 2606
rect 2811 2610 2815 2611
rect 2811 2605 2815 2606
rect 2827 2610 2831 2611
rect 2827 2605 2831 2606
rect 2947 2610 2951 2611
rect 2947 2605 2951 2606
rect 3019 2610 3023 2611
rect 3019 2605 3023 2606
rect 3083 2610 3087 2611
rect 3083 2605 3087 2606
rect 3211 2610 3215 2611
rect 3211 2605 3215 2606
rect 3219 2610 3223 2611
rect 3219 2605 3223 2606
rect 3355 2610 3359 2611
rect 3355 2605 3359 2606
rect 3403 2610 3407 2611
rect 3403 2605 3407 2606
rect 3799 2610 3803 2611
rect 3840 2609 3842 2669
rect 3799 2605 3803 2606
rect 3838 2608 3844 2609
rect 4028 2608 4030 2669
rect 4276 2608 4278 2669
rect 4556 2608 4558 2669
rect 4868 2608 4870 2669
rect 5204 2608 5206 2669
rect 5516 2608 5518 2669
rect 5664 2609 5666 2669
rect 5662 2608 5668 2609
rect 1934 2592 1940 2593
rect 110 2588 111 2592
rect 115 2588 116 2592
rect 110 2587 116 2588
rect 538 2591 544 2592
rect 538 2587 539 2591
rect 543 2587 544 2591
rect 538 2586 544 2587
rect 698 2591 704 2592
rect 698 2587 699 2591
rect 703 2587 704 2591
rect 698 2586 704 2587
rect 882 2591 888 2592
rect 882 2587 883 2591
rect 887 2587 888 2591
rect 882 2586 888 2587
rect 1090 2591 1096 2592
rect 1090 2587 1091 2591
rect 1095 2587 1096 2591
rect 1090 2586 1096 2587
rect 1322 2591 1328 2592
rect 1322 2587 1323 2591
rect 1327 2587 1328 2591
rect 1322 2586 1328 2587
rect 1562 2591 1568 2592
rect 1562 2587 1563 2591
rect 1567 2587 1568 2591
rect 1562 2586 1568 2587
rect 1786 2591 1792 2592
rect 1786 2587 1787 2591
rect 1791 2587 1792 2591
rect 1934 2588 1935 2592
rect 1939 2588 1940 2592
rect 1934 2587 1940 2588
rect 1786 2586 1792 2587
rect 566 2576 572 2577
rect 110 2575 116 2576
rect 110 2571 111 2575
rect 115 2571 116 2575
rect 566 2572 567 2576
rect 571 2572 572 2576
rect 566 2571 572 2572
rect 726 2576 732 2577
rect 726 2572 727 2576
rect 731 2572 732 2576
rect 726 2571 732 2572
rect 910 2576 916 2577
rect 910 2572 911 2576
rect 915 2572 916 2576
rect 910 2571 916 2572
rect 1118 2576 1124 2577
rect 1118 2572 1119 2576
rect 1123 2572 1124 2576
rect 1118 2571 1124 2572
rect 1350 2576 1356 2577
rect 1350 2572 1351 2576
rect 1355 2572 1356 2576
rect 1350 2571 1356 2572
rect 1590 2576 1596 2577
rect 1590 2572 1591 2576
rect 1595 2572 1596 2576
rect 1590 2571 1596 2572
rect 1814 2576 1820 2577
rect 1814 2572 1815 2576
rect 1819 2572 1820 2576
rect 1814 2571 1820 2572
rect 1934 2575 1940 2576
rect 1934 2571 1935 2575
rect 1939 2571 1940 2575
rect 110 2570 116 2571
rect 112 2535 114 2570
rect 568 2535 570 2571
rect 728 2535 730 2571
rect 912 2535 914 2571
rect 1120 2535 1122 2571
rect 1352 2535 1354 2571
rect 1592 2535 1594 2571
rect 1816 2535 1818 2571
rect 1934 2570 1940 2571
rect 1936 2535 1938 2570
rect 1976 2545 1978 2605
rect 1974 2544 1980 2545
rect 1996 2544 1998 2605
rect 2204 2544 2206 2605
rect 2420 2544 2422 2605
rect 2628 2544 2630 2605
rect 2828 2544 2830 2605
rect 3020 2544 3022 2605
rect 3212 2544 3214 2605
rect 3404 2544 3406 2605
rect 3800 2545 3802 2605
rect 3838 2604 3839 2608
rect 3843 2604 3844 2608
rect 3838 2603 3844 2604
rect 4026 2607 4032 2608
rect 4026 2603 4027 2607
rect 4031 2603 4032 2607
rect 4026 2602 4032 2603
rect 4274 2607 4280 2608
rect 4274 2603 4275 2607
rect 4279 2603 4280 2607
rect 4274 2602 4280 2603
rect 4554 2607 4560 2608
rect 4554 2603 4555 2607
rect 4559 2603 4560 2607
rect 4554 2602 4560 2603
rect 4866 2607 4872 2608
rect 4866 2603 4867 2607
rect 4871 2603 4872 2607
rect 4866 2602 4872 2603
rect 5202 2607 5208 2608
rect 5202 2603 5203 2607
rect 5207 2603 5208 2607
rect 5202 2602 5208 2603
rect 5514 2607 5520 2608
rect 5514 2603 5515 2607
rect 5519 2603 5520 2607
rect 5662 2604 5663 2608
rect 5667 2604 5668 2608
rect 5662 2603 5668 2604
rect 5514 2602 5520 2603
rect 4054 2592 4060 2593
rect 3838 2591 3844 2592
rect 3838 2587 3839 2591
rect 3843 2587 3844 2591
rect 4054 2588 4055 2592
rect 4059 2588 4060 2592
rect 4054 2587 4060 2588
rect 4302 2592 4308 2593
rect 4302 2588 4303 2592
rect 4307 2588 4308 2592
rect 4302 2587 4308 2588
rect 4582 2592 4588 2593
rect 4582 2588 4583 2592
rect 4587 2588 4588 2592
rect 4582 2587 4588 2588
rect 4894 2592 4900 2593
rect 4894 2588 4895 2592
rect 4899 2588 4900 2592
rect 4894 2587 4900 2588
rect 5230 2592 5236 2593
rect 5230 2588 5231 2592
rect 5235 2588 5236 2592
rect 5230 2587 5236 2588
rect 5542 2592 5548 2593
rect 5542 2588 5543 2592
rect 5547 2588 5548 2592
rect 5542 2587 5548 2588
rect 5662 2591 5668 2592
rect 5662 2587 5663 2591
rect 5667 2587 5668 2591
rect 3838 2586 3844 2587
rect 3840 2559 3842 2586
rect 4056 2559 4058 2587
rect 4304 2559 4306 2587
rect 4584 2559 4586 2587
rect 4896 2559 4898 2587
rect 5232 2559 5234 2587
rect 5544 2559 5546 2587
rect 5662 2586 5668 2587
rect 5664 2559 5666 2586
rect 3839 2558 3843 2559
rect 3839 2553 3843 2554
rect 4055 2558 4059 2559
rect 4055 2553 4059 2554
rect 4303 2558 4307 2559
rect 4303 2553 4307 2554
rect 4335 2558 4339 2559
rect 4335 2553 4339 2554
rect 4559 2558 4563 2559
rect 4559 2553 4563 2554
rect 4583 2558 4587 2559
rect 4583 2553 4587 2554
rect 4799 2558 4803 2559
rect 4799 2553 4803 2554
rect 4895 2558 4899 2559
rect 4895 2553 4899 2554
rect 5047 2558 5051 2559
rect 5047 2553 5051 2554
rect 5231 2558 5235 2559
rect 5231 2553 5235 2554
rect 5303 2558 5307 2559
rect 5303 2553 5307 2554
rect 5543 2558 5547 2559
rect 5543 2553 5547 2554
rect 5663 2558 5667 2559
rect 5663 2553 5667 2554
rect 3798 2544 3804 2545
rect 1974 2540 1975 2544
rect 1979 2540 1980 2544
rect 1974 2539 1980 2540
rect 1994 2543 2000 2544
rect 1994 2539 1995 2543
rect 1999 2539 2000 2543
rect 1994 2538 2000 2539
rect 2202 2543 2208 2544
rect 2202 2539 2203 2543
rect 2207 2539 2208 2543
rect 2202 2538 2208 2539
rect 2418 2543 2424 2544
rect 2418 2539 2419 2543
rect 2423 2539 2424 2543
rect 2418 2538 2424 2539
rect 2626 2543 2632 2544
rect 2626 2539 2627 2543
rect 2631 2539 2632 2543
rect 2626 2538 2632 2539
rect 2826 2543 2832 2544
rect 2826 2539 2827 2543
rect 2831 2539 2832 2543
rect 2826 2538 2832 2539
rect 3018 2543 3024 2544
rect 3018 2539 3019 2543
rect 3023 2539 3024 2543
rect 3018 2538 3024 2539
rect 3210 2543 3216 2544
rect 3210 2539 3211 2543
rect 3215 2539 3216 2543
rect 3210 2538 3216 2539
rect 3402 2543 3408 2544
rect 3402 2539 3403 2543
rect 3407 2539 3408 2543
rect 3798 2540 3799 2544
rect 3803 2540 3804 2544
rect 3798 2539 3804 2540
rect 3402 2538 3408 2539
rect 111 2534 115 2535
rect 111 2529 115 2530
rect 567 2534 571 2535
rect 567 2529 571 2530
rect 695 2534 699 2535
rect 695 2529 699 2530
rect 727 2534 731 2535
rect 727 2529 731 2530
rect 847 2534 851 2535
rect 847 2529 851 2530
rect 911 2534 915 2535
rect 911 2529 915 2530
rect 999 2534 1003 2535
rect 999 2529 1003 2530
rect 1119 2534 1123 2535
rect 1119 2529 1123 2530
rect 1159 2534 1163 2535
rect 1159 2529 1163 2530
rect 1327 2534 1331 2535
rect 1327 2529 1331 2530
rect 1351 2534 1355 2535
rect 1351 2529 1355 2530
rect 1495 2534 1499 2535
rect 1495 2529 1499 2530
rect 1591 2534 1595 2535
rect 1591 2529 1595 2530
rect 1663 2534 1667 2535
rect 1663 2529 1667 2530
rect 1815 2534 1819 2535
rect 1815 2529 1819 2530
rect 1935 2534 1939 2535
rect 3840 2530 3842 2553
rect 1935 2529 1939 2530
rect 3838 2529 3844 2530
rect 4336 2529 4338 2553
rect 4560 2529 4562 2553
rect 4800 2529 4802 2553
rect 5048 2529 5050 2553
rect 5304 2529 5306 2553
rect 5544 2529 5546 2553
rect 5664 2530 5666 2553
rect 5662 2529 5668 2530
rect 112 2506 114 2529
rect 110 2505 116 2506
rect 696 2505 698 2529
rect 848 2505 850 2529
rect 1000 2505 1002 2529
rect 1160 2505 1162 2529
rect 1328 2505 1330 2529
rect 1496 2505 1498 2529
rect 1664 2505 1666 2529
rect 1816 2505 1818 2529
rect 1936 2506 1938 2529
rect 2022 2528 2028 2529
rect 1974 2527 1980 2528
rect 1974 2523 1975 2527
rect 1979 2523 1980 2527
rect 2022 2524 2023 2528
rect 2027 2524 2028 2528
rect 2022 2523 2028 2524
rect 2230 2528 2236 2529
rect 2230 2524 2231 2528
rect 2235 2524 2236 2528
rect 2230 2523 2236 2524
rect 2446 2528 2452 2529
rect 2446 2524 2447 2528
rect 2451 2524 2452 2528
rect 2446 2523 2452 2524
rect 2654 2528 2660 2529
rect 2654 2524 2655 2528
rect 2659 2524 2660 2528
rect 2654 2523 2660 2524
rect 2854 2528 2860 2529
rect 2854 2524 2855 2528
rect 2859 2524 2860 2528
rect 2854 2523 2860 2524
rect 3046 2528 3052 2529
rect 3046 2524 3047 2528
rect 3051 2524 3052 2528
rect 3046 2523 3052 2524
rect 3238 2528 3244 2529
rect 3238 2524 3239 2528
rect 3243 2524 3244 2528
rect 3238 2523 3244 2524
rect 3430 2528 3436 2529
rect 3430 2524 3431 2528
rect 3435 2524 3436 2528
rect 3430 2523 3436 2524
rect 3798 2527 3804 2528
rect 3798 2523 3799 2527
rect 3803 2523 3804 2527
rect 3838 2525 3839 2529
rect 3843 2525 3844 2529
rect 3838 2524 3844 2525
rect 4334 2528 4340 2529
rect 4334 2524 4335 2528
rect 4339 2524 4340 2528
rect 4334 2523 4340 2524
rect 4558 2528 4564 2529
rect 4558 2524 4559 2528
rect 4563 2524 4564 2528
rect 4558 2523 4564 2524
rect 4798 2528 4804 2529
rect 4798 2524 4799 2528
rect 4803 2524 4804 2528
rect 4798 2523 4804 2524
rect 5046 2528 5052 2529
rect 5046 2524 5047 2528
rect 5051 2524 5052 2528
rect 5046 2523 5052 2524
rect 5302 2528 5308 2529
rect 5302 2524 5303 2528
rect 5307 2524 5308 2528
rect 5302 2523 5308 2524
rect 5542 2528 5548 2529
rect 5542 2524 5543 2528
rect 5547 2524 5548 2528
rect 5662 2525 5663 2529
rect 5667 2525 5668 2529
rect 5662 2524 5668 2525
rect 5542 2523 5548 2524
rect 1974 2522 1980 2523
rect 1934 2505 1940 2506
rect 110 2501 111 2505
rect 115 2501 116 2505
rect 110 2500 116 2501
rect 694 2504 700 2505
rect 694 2500 695 2504
rect 699 2500 700 2504
rect 694 2499 700 2500
rect 846 2504 852 2505
rect 846 2500 847 2504
rect 851 2500 852 2504
rect 846 2499 852 2500
rect 998 2504 1004 2505
rect 998 2500 999 2504
rect 1003 2500 1004 2504
rect 998 2499 1004 2500
rect 1158 2504 1164 2505
rect 1158 2500 1159 2504
rect 1163 2500 1164 2504
rect 1158 2499 1164 2500
rect 1326 2504 1332 2505
rect 1326 2500 1327 2504
rect 1331 2500 1332 2504
rect 1326 2499 1332 2500
rect 1494 2504 1500 2505
rect 1494 2500 1495 2504
rect 1499 2500 1500 2504
rect 1494 2499 1500 2500
rect 1662 2504 1668 2505
rect 1662 2500 1663 2504
rect 1667 2500 1668 2504
rect 1662 2499 1668 2500
rect 1814 2504 1820 2505
rect 1814 2500 1815 2504
rect 1819 2500 1820 2504
rect 1934 2501 1935 2505
rect 1939 2501 1940 2505
rect 1934 2500 1940 2501
rect 1814 2499 1820 2500
rect 1976 2491 1978 2522
rect 2024 2491 2026 2523
rect 2232 2491 2234 2523
rect 2448 2491 2450 2523
rect 2656 2491 2658 2523
rect 2856 2491 2858 2523
rect 3048 2491 3050 2523
rect 3240 2491 3242 2523
rect 3432 2491 3434 2523
rect 3798 2522 3804 2523
rect 3800 2491 3802 2522
rect 4306 2513 4312 2514
rect 3838 2512 3844 2513
rect 3838 2508 3839 2512
rect 3843 2508 3844 2512
rect 4306 2509 4307 2513
rect 4311 2509 4312 2513
rect 4306 2508 4312 2509
rect 4530 2513 4536 2514
rect 4530 2509 4531 2513
rect 4535 2509 4536 2513
rect 4530 2508 4536 2509
rect 4770 2513 4776 2514
rect 4770 2509 4771 2513
rect 4775 2509 4776 2513
rect 4770 2508 4776 2509
rect 5018 2513 5024 2514
rect 5018 2509 5019 2513
rect 5023 2509 5024 2513
rect 5018 2508 5024 2509
rect 5274 2513 5280 2514
rect 5274 2509 5275 2513
rect 5279 2509 5280 2513
rect 5274 2508 5280 2509
rect 5514 2513 5520 2514
rect 5514 2509 5515 2513
rect 5519 2509 5520 2513
rect 5514 2508 5520 2509
rect 5662 2512 5668 2513
rect 5662 2508 5663 2512
rect 5667 2508 5668 2512
rect 3838 2507 3844 2508
rect 1975 2490 1979 2491
rect 666 2489 672 2490
rect 110 2488 116 2489
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 666 2485 667 2489
rect 671 2485 672 2489
rect 666 2484 672 2485
rect 818 2489 824 2490
rect 818 2485 819 2489
rect 823 2485 824 2489
rect 818 2484 824 2485
rect 970 2489 976 2490
rect 970 2485 971 2489
rect 975 2485 976 2489
rect 970 2484 976 2485
rect 1130 2489 1136 2490
rect 1130 2485 1131 2489
rect 1135 2485 1136 2489
rect 1130 2484 1136 2485
rect 1298 2489 1304 2490
rect 1298 2485 1299 2489
rect 1303 2485 1304 2489
rect 1298 2484 1304 2485
rect 1466 2489 1472 2490
rect 1466 2485 1467 2489
rect 1471 2485 1472 2489
rect 1466 2484 1472 2485
rect 1634 2489 1640 2490
rect 1634 2485 1635 2489
rect 1639 2485 1640 2489
rect 1634 2484 1640 2485
rect 1786 2489 1792 2490
rect 1786 2485 1787 2489
rect 1791 2485 1792 2489
rect 1786 2484 1792 2485
rect 1934 2488 1940 2489
rect 1934 2484 1935 2488
rect 1939 2484 1940 2488
rect 1975 2485 1979 2486
rect 2023 2490 2027 2491
rect 2023 2485 2027 2486
rect 2231 2490 2235 2491
rect 2231 2485 2235 2486
rect 2319 2490 2323 2491
rect 2319 2485 2323 2486
rect 2447 2490 2451 2491
rect 2447 2485 2451 2486
rect 2567 2490 2571 2491
rect 2567 2485 2571 2486
rect 2655 2490 2659 2491
rect 2655 2485 2659 2486
rect 2799 2490 2803 2491
rect 2799 2485 2803 2486
rect 2855 2490 2859 2491
rect 2855 2485 2859 2486
rect 3023 2490 3027 2491
rect 3023 2485 3027 2486
rect 3047 2490 3051 2491
rect 3047 2485 3051 2486
rect 3239 2490 3243 2491
rect 3239 2485 3243 2486
rect 3431 2490 3435 2491
rect 3431 2485 3435 2486
rect 3455 2490 3459 2491
rect 3455 2485 3459 2486
rect 3671 2490 3675 2491
rect 3671 2485 3675 2486
rect 3799 2490 3803 2491
rect 3799 2485 3803 2486
rect 110 2483 116 2484
rect 112 2415 114 2483
rect 668 2415 670 2484
rect 820 2415 822 2484
rect 972 2415 974 2484
rect 1132 2415 1134 2484
rect 1300 2415 1302 2484
rect 1468 2415 1470 2484
rect 1636 2415 1638 2484
rect 1788 2415 1790 2484
rect 1934 2483 1940 2484
rect 1936 2415 1938 2483
rect 1976 2462 1978 2485
rect 1974 2461 1980 2462
rect 2320 2461 2322 2485
rect 2568 2461 2570 2485
rect 2800 2461 2802 2485
rect 3024 2461 3026 2485
rect 3240 2461 3242 2485
rect 3456 2461 3458 2485
rect 3672 2461 3674 2485
rect 3800 2462 3802 2485
rect 3798 2461 3804 2462
rect 1974 2457 1975 2461
rect 1979 2457 1980 2461
rect 1974 2456 1980 2457
rect 2318 2460 2324 2461
rect 2318 2456 2319 2460
rect 2323 2456 2324 2460
rect 2318 2455 2324 2456
rect 2566 2460 2572 2461
rect 2566 2456 2567 2460
rect 2571 2456 2572 2460
rect 2566 2455 2572 2456
rect 2798 2460 2804 2461
rect 2798 2456 2799 2460
rect 2803 2456 2804 2460
rect 2798 2455 2804 2456
rect 3022 2460 3028 2461
rect 3022 2456 3023 2460
rect 3027 2456 3028 2460
rect 3022 2455 3028 2456
rect 3238 2460 3244 2461
rect 3238 2456 3239 2460
rect 3243 2456 3244 2460
rect 3238 2455 3244 2456
rect 3454 2460 3460 2461
rect 3454 2456 3455 2460
rect 3459 2456 3460 2460
rect 3454 2455 3460 2456
rect 3670 2460 3676 2461
rect 3670 2456 3671 2460
rect 3675 2456 3676 2460
rect 3798 2457 3799 2461
rect 3803 2457 3804 2461
rect 3798 2456 3804 2457
rect 3670 2455 3676 2456
rect 2290 2445 2296 2446
rect 1974 2444 1980 2445
rect 1974 2440 1975 2444
rect 1979 2440 1980 2444
rect 2290 2441 2291 2445
rect 2295 2441 2296 2445
rect 2290 2440 2296 2441
rect 2538 2445 2544 2446
rect 2538 2441 2539 2445
rect 2543 2441 2544 2445
rect 2538 2440 2544 2441
rect 2770 2445 2776 2446
rect 2770 2441 2771 2445
rect 2775 2441 2776 2445
rect 2770 2440 2776 2441
rect 2994 2445 3000 2446
rect 2994 2441 2995 2445
rect 2999 2441 3000 2445
rect 2994 2440 3000 2441
rect 3210 2445 3216 2446
rect 3210 2441 3211 2445
rect 3215 2441 3216 2445
rect 3210 2440 3216 2441
rect 3426 2445 3432 2446
rect 3426 2441 3427 2445
rect 3431 2441 3432 2445
rect 3426 2440 3432 2441
rect 3642 2445 3648 2446
rect 3642 2441 3643 2445
rect 3647 2441 3648 2445
rect 3642 2440 3648 2441
rect 3798 2444 3804 2445
rect 3798 2440 3799 2444
rect 3803 2440 3804 2444
rect 1974 2439 1980 2440
rect 111 2414 115 2415
rect 111 2409 115 2410
rect 355 2414 359 2415
rect 355 2409 359 2410
rect 507 2414 511 2415
rect 507 2409 511 2410
rect 667 2414 671 2415
rect 667 2409 671 2410
rect 675 2414 679 2415
rect 675 2409 679 2410
rect 819 2414 823 2415
rect 819 2409 823 2410
rect 859 2414 863 2415
rect 859 2409 863 2410
rect 971 2414 975 2415
rect 971 2409 975 2410
rect 1059 2414 1063 2415
rect 1059 2409 1063 2410
rect 1131 2414 1135 2415
rect 1131 2409 1135 2410
rect 1267 2414 1271 2415
rect 1267 2409 1271 2410
rect 1299 2414 1303 2415
rect 1299 2409 1303 2410
rect 1467 2414 1471 2415
rect 1467 2409 1471 2410
rect 1483 2414 1487 2415
rect 1483 2409 1487 2410
rect 1635 2414 1639 2415
rect 1635 2409 1639 2410
rect 1699 2414 1703 2415
rect 1699 2409 1703 2410
rect 1787 2414 1791 2415
rect 1787 2409 1791 2410
rect 1935 2414 1939 2415
rect 1935 2409 1939 2410
rect 112 2349 114 2409
rect 110 2348 116 2349
rect 356 2348 358 2409
rect 508 2348 510 2409
rect 676 2348 678 2409
rect 860 2348 862 2409
rect 1060 2348 1062 2409
rect 1268 2348 1270 2409
rect 1484 2348 1486 2409
rect 1700 2348 1702 2409
rect 1936 2349 1938 2409
rect 1976 2371 1978 2439
rect 2292 2371 2294 2440
rect 2540 2371 2542 2440
rect 2772 2371 2774 2440
rect 2996 2371 2998 2440
rect 3212 2371 3214 2440
rect 3428 2371 3430 2440
rect 3644 2371 3646 2440
rect 3798 2439 3804 2440
rect 3800 2371 3802 2439
rect 3840 2431 3842 2507
rect 4308 2431 4310 2508
rect 4532 2431 4534 2508
rect 4772 2431 4774 2508
rect 5020 2431 5022 2508
rect 5276 2431 5278 2508
rect 5516 2431 5518 2508
rect 5662 2507 5668 2508
rect 5664 2431 5666 2507
rect 3839 2430 3843 2431
rect 3839 2425 3843 2426
rect 4307 2430 4311 2431
rect 4307 2425 4311 2426
rect 4491 2430 4495 2431
rect 4491 2425 4495 2426
rect 4531 2430 4535 2431
rect 4531 2425 4535 2426
rect 4635 2430 4639 2431
rect 4635 2425 4639 2426
rect 4771 2430 4775 2431
rect 4771 2425 4775 2426
rect 4795 2430 4799 2431
rect 4795 2425 4799 2426
rect 4963 2430 4967 2431
rect 4963 2425 4967 2426
rect 5019 2430 5023 2431
rect 5019 2425 5023 2426
rect 5139 2430 5143 2431
rect 5139 2425 5143 2426
rect 5275 2430 5279 2431
rect 5275 2425 5279 2426
rect 5323 2430 5327 2431
rect 5323 2425 5327 2426
rect 5515 2430 5519 2431
rect 5515 2425 5519 2426
rect 5663 2430 5667 2431
rect 5663 2425 5667 2426
rect 1975 2370 1979 2371
rect 1975 2365 1979 2366
rect 2291 2370 2295 2371
rect 2291 2365 2295 2366
rect 2331 2370 2335 2371
rect 2331 2365 2335 2366
rect 2539 2370 2543 2371
rect 2539 2365 2543 2366
rect 2739 2370 2743 2371
rect 2739 2365 2743 2366
rect 2771 2370 2775 2371
rect 2771 2365 2775 2366
rect 2931 2370 2935 2371
rect 2931 2365 2935 2366
rect 2995 2370 2999 2371
rect 2995 2365 2999 2366
rect 3123 2370 3127 2371
rect 3123 2365 3127 2366
rect 3211 2370 3215 2371
rect 3211 2365 3215 2366
rect 3307 2370 3311 2371
rect 3307 2365 3311 2366
rect 3427 2370 3431 2371
rect 3427 2365 3431 2366
rect 3491 2370 3495 2371
rect 3491 2365 3495 2366
rect 3643 2370 3647 2371
rect 3643 2365 3647 2366
rect 3651 2370 3655 2371
rect 3651 2365 3655 2366
rect 3799 2370 3803 2371
rect 3799 2365 3803 2366
rect 3840 2365 3842 2425
rect 1934 2348 1940 2349
rect 110 2344 111 2348
rect 115 2344 116 2348
rect 110 2343 116 2344
rect 354 2347 360 2348
rect 354 2343 355 2347
rect 359 2343 360 2347
rect 354 2342 360 2343
rect 506 2347 512 2348
rect 506 2343 507 2347
rect 511 2343 512 2347
rect 506 2342 512 2343
rect 674 2347 680 2348
rect 674 2343 675 2347
rect 679 2343 680 2347
rect 674 2342 680 2343
rect 858 2347 864 2348
rect 858 2343 859 2347
rect 863 2343 864 2347
rect 858 2342 864 2343
rect 1058 2347 1064 2348
rect 1058 2343 1059 2347
rect 1063 2343 1064 2347
rect 1058 2342 1064 2343
rect 1266 2347 1272 2348
rect 1266 2343 1267 2347
rect 1271 2343 1272 2347
rect 1266 2342 1272 2343
rect 1482 2347 1488 2348
rect 1482 2343 1483 2347
rect 1487 2343 1488 2347
rect 1482 2342 1488 2343
rect 1698 2347 1704 2348
rect 1698 2343 1699 2347
rect 1703 2343 1704 2347
rect 1934 2344 1935 2348
rect 1939 2344 1940 2348
rect 1934 2343 1940 2344
rect 1698 2342 1704 2343
rect 382 2332 388 2333
rect 110 2331 116 2332
rect 110 2327 111 2331
rect 115 2327 116 2331
rect 382 2328 383 2332
rect 387 2328 388 2332
rect 382 2327 388 2328
rect 534 2332 540 2333
rect 534 2328 535 2332
rect 539 2328 540 2332
rect 534 2327 540 2328
rect 702 2332 708 2333
rect 702 2328 703 2332
rect 707 2328 708 2332
rect 702 2327 708 2328
rect 886 2332 892 2333
rect 886 2328 887 2332
rect 891 2328 892 2332
rect 886 2327 892 2328
rect 1086 2332 1092 2333
rect 1086 2328 1087 2332
rect 1091 2328 1092 2332
rect 1086 2327 1092 2328
rect 1294 2332 1300 2333
rect 1294 2328 1295 2332
rect 1299 2328 1300 2332
rect 1294 2327 1300 2328
rect 1510 2332 1516 2333
rect 1510 2328 1511 2332
rect 1515 2328 1516 2332
rect 1510 2327 1516 2328
rect 1726 2332 1732 2333
rect 1726 2328 1727 2332
rect 1731 2328 1732 2332
rect 1726 2327 1732 2328
rect 1934 2331 1940 2332
rect 1934 2327 1935 2331
rect 1939 2327 1940 2331
rect 110 2326 116 2327
rect 112 2295 114 2326
rect 384 2295 386 2327
rect 536 2295 538 2327
rect 704 2295 706 2327
rect 888 2295 890 2327
rect 1088 2295 1090 2327
rect 1296 2295 1298 2327
rect 1512 2295 1514 2327
rect 1728 2295 1730 2327
rect 1934 2326 1940 2327
rect 1936 2295 1938 2326
rect 1976 2305 1978 2365
rect 1974 2304 1980 2305
rect 2332 2304 2334 2365
rect 2540 2304 2542 2365
rect 2740 2304 2742 2365
rect 2932 2304 2934 2365
rect 3124 2304 3126 2365
rect 3308 2304 3310 2365
rect 3492 2304 3494 2365
rect 3652 2304 3654 2365
rect 3800 2305 3802 2365
rect 3838 2364 3844 2365
rect 4492 2364 4494 2425
rect 4636 2364 4638 2425
rect 4796 2364 4798 2425
rect 4964 2364 4966 2425
rect 5140 2364 5142 2425
rect 5324 2364 5326 2425
rect 5516 2364 5518 2425
rect 5664 2365 5666 2425
rect 5662 2364 5668 2365
rect 3838 2360 3839 2364
rect 3843 2360 3844 2364
rect 3838 2359 3844 2360
rect 4490 2363 4496 2364
rect 4490 2359 4491 2363
rect 4495 2359 4496 2363
rect 4490 2358 4496 2359
rect 4634 2363 4640 2364
rect 4634 2359 4635 2363
rect 4639 2359 4640 2363
rect 4634 2358 4640 2359
rect 4794 2363 4800 2364
rect 4794 2359 4795 2363
rect 4799 2359 4800 2363
rect 4794 2358 4800 2359
rect 4962 2363 4968 2364
rect 4962 2359 4963 2363
rect 4967 2359 4968 2363
rect 4962 2358 4968 2359
rect 5138 2363 5144 2364
rect 5138 2359 5139 2363
rect 5143 2359 5144 2363
rect 5138 2358 5144 2359
rect 5322 2363 5328 2364
rect 5322 2359 5323 2363
rect 5327 2359 5328 2363
rect 5322 2358 5328 2359
rect 5514 2363 5520 2364
rect 5514 2359 5515 2363
rect 5519 2359 5520 2363
rect 5662 2360 5663 2364
rect 5667 2360 5668 2364
rect 5662 2359 5668 2360
rect 5514 2358 5520 2359
rect 4518 2348 4524 2349
rect 3838 2347 3844 2348
rect 3838 2343 3839 2347
rect 3843 2343 3844 2347
rect 4518 2344 4519 2348
rect 4523 2344 4524 2348
rect 4518 2343 4524 2344
rect 4662 2348 4668 2349
rect 4662 2344 4663 2348
rect 4667 2344 4668 2348
rect 4662 2343 4668 2344
rect 4822 2348 4828 2349
rect 4822 2344 4823 2348
rect 4827 2344 4828 2348
rect 4822 2343 4828 2344
rect 4990 2348 4996 2349
rect 4990 2344 4991 2348
rect 4995 2344 4996 2348
rect 4990 2343 4996 2344
rect 5166 2348 5172 2349
rect 5166 2344 5167 2348
rect 5171 2344 5172 2348
rect 5166 2343 5172 2344
rect 5350 2348 5356 2349
rect 5350 2344 5351 2348
rect 5355 2344 5356 2348
rect 5350 2343 5356 2344
rect 5542 2348 5548 2349
rect 5542 2344 5543 2348
rect 5547 2344 5548 2348
rect 5542 2343 5548 2344
rect 5662 2347 5668 2348
rect 5662 2343 5663 2347
rect 5667 2343 5668 2347
rect 3838 2342 3844 2343
rect 3798 2304 3804 2305
rect 1974 2300 1975 2304
rect 1979 2300 1980 2304
rect 1974 2299 1980 2300
rect 2330 2303 2336 2304
rect 2330 2299 2331 2303
rect 2335 2299 2336 2303
rect 2330 2298 2336 2299
rect 2538 2303 2544 2304
rect 2538 2299 2539 2303
rect 2543 2299 2544 2303
rect 2538 2298 2544 2299
rect 2738 2303 2744 2304
rect 2738 2299 2739 2303
rect 2743 2299 2744 2303
rect 2738 2298 2744 2299
rect 2930 2303 2936 2304
rect 2930 2299 2931 2303
rect 2935 2299 2936 2303
rect 2930 2298 2936 2299
rect 3122 2303 3128 2304
rect 3122 2299 3123 2303
rect 3127 2299 3128 2303
rect 3122 2298 3128 2299
rect 3306 2303 3312 2304
rect 3306 2299 3307 2303
rect 3311 2299 3312 2303
rect 3306 2298 3312 2299
rect 3490 2303 3496 2304
rect 3490 2299 3491 2303
rect 3495 2299 3496 2303
rect 3490 2298 3496 2299
rect 3650 2303 3656 2304
rect 3650 2299 3651 2303
rect 3655 2299 3656 2303
rect 3798 2300 3799 2304
rect 3803 2300 3804 2304
rect 3798 2299 3804 2300
rect 3840 2299 3842 2342
rect 4520 2299 4522 2343
rect 4664 2299 4666 2343
rect 4824 2299 4826 2343
rect 4992 2299 4994 2343
rect 5168 2299 5170 2343
rect 5352 2299 5354 2343
rect 5544 2299 5546 2343
rect 5662 2342 5668 2343
rect 5664 2299 5666 2342
rect 3650 2298 3656 2299
rect 3839 2298 3843 2299
rect 111 2294 115 2295
rect 111 2289 115 2290
rect 159 2294 163 2295
rect 159 2289 163 2290
rect 335 2294 339 2295
rect 335 2289 339 2290
rect 383 2294 387 2295
rect 383 2289 387 2290
rect 535 2294 539 2295
rect 535 2289 539 2290
rect 543 2294 547 2295
rect 543 2289 547 2290
rect 703 2294 707 2295
rect 703 2289 707 2290
rect 759 2294 763 2295
rect 759 2289 763 2290
rect 887 2294 891 2295
rect 887 2289 891 2290
rect 975 2294 979 2295
rect 975 2289 979 2290
rect 1087 2294 1091 2295
rect 1087 2289 1091 2290
rect 1199 2294 1203 2295
rect 1199 2289 1203 2290
rect 1295 2294 1299 2295
rect 1295 2289 1299 2290
rect 1431 2294 1435 2295
rect 1431 2289 1435 2290
rect 1511 2294 1515 2295
rect 1511 2289 1515 2290
rect 1671 2294 1675 2295
rect 1671 2289 1675 2290
rect 1727 2294 1731 2295
rect 1727 2289 1731 2290
rect 1935 2294 1939 2295
rect 3839 2293 3843 2294
rect 3887 2298 3891 2299
rect 3887 2293 3891 2294
rect 4071 2298 4075 2299
rect 4071 2293 4075 2294
rect 4271 2298 4275 2299
rect 4271 2293 4275 2294
rect 4463 2298 4467 2299
rect 4463 2293 4467 2294
rect 4519 2298 4523 2299
rect 4519 2293 4523 2294
rect 4655 2298 4659 2299
rect 4655 2293 4659 2294
rect 4663 2298 4667 2299
rect 4663 2293 4667 2294
rect 4823 2298 4827 2299
rect 4823 2293 4827 2294
rect 4839 2298 4843 2299
rect 4839 2293 4843 2294
rect 4991 2298 4995 2299
rect 4991 2293 4995 2294
rect 5015 2298 5019 2299
rect 5015 2293 5019 2294
rect 5167 2298 5171 2299
rect 5167 2293 5171 2294
rect 5183 2298 5187 2299
rect 5183 2293 5187 2294
rect 5351 2298 5355 2299
rect 5351 2293 5355 2294
rect 5359 2298 5363 2299
rect 5359 2293 5363 2294
rect 5535 2298 5539 2299
rect 5535 2293 5539 2294
rect 5543 2298 5547 2299
rect 5543 2293 5547 2294
rect 5663 2298 5667 2299
rect 5663 2293 5667 2294
rect 1935 2289 1939 2290
rect 112 2266 114 2289
rect 110 2265 116 2266
rect 160 2265 162 2289
rect 336 2265 338 2289
rect 544 2265 546 2289
rect 760 2265 762 2289
rect 976 2265 978 2289
rect 1200 2265 1202 2289
rect 1432 2265 1434 2289
rect 1672 2265 1674 2289
rect 1936 2266 1938 2289
rect 2358 2288 2364 2289
rect 1974 2287 1980 2288
rect 1974 2283 1975 2287
rect 1979 2283 1980 2287
rect 2358 2284 2359 2288
rect 2363 2284 2364 2288
rect 2358 2283 2364 2284
rect 2566 2288 2572 2289
rect 2566 2284 2567 2288
rect 2571 2284 2572 2288
rect 2566 2283 2572 2284
rect 2766 2288 2772 2289
rect 2766 2284 2767 2288
rect 2771 2284 2772 2288
rect 2766 2283 2772 2284
rect 2958 2288 2964 2289
rect 2958 2284 2959 2288
rect 2963 2284 2964 2288
rect 2958 2283 2964 2284
rect 3150 2288 3156 2289
rect 3150 2284 3151 2288
rect 3155 2284 3156 2288
rect 3150 2283 3156 2284
rect 3334 2288 3340 2289
rect 3334 2284 3335 2288
rect 3339 2284 3340 2288
rect 3334 2283 3340 2284
rect 3518 2288 3524 2289
rect 3518 2284 3519 2288
rect 3523 2284 3524 2288
rect 3518 2283 3524 2284
rect 3678 2288 3684 2289
rect 3678 2284 3679 2288
rect 3683 2284 3684 2288
rect 3678 2283 3684 2284
rect 3798 2287 3804 2288
rect 3798 2283 3799 2287
rect 3803 2283 3804 2287
rect 1974 2282 1980 2283
rect 1934 2265 1940 2266
rect 110 2261 111 2265
rect 115 2261 116 2265
rect 110 2260 116 2261
rect 158 2264 164 2265
rect 158 2260 159 2264
rect 163 2260 164 2264
rect 158 2259 164 2260
rect 334 2264 340 2265
rect 334 2260 335 2264
rect 339 2260 340 2264
rect 334 2259 340 2260
rect 542 2264 548 2265
rect 542 2260 543 2264
rect 547 2260 548 2264
rect 542 2259 548 2260
rect 758 2264 764 2265
rect 758 2260 759 2264
rect 763 2260 764 2264
rect 758 2259 764 2260
rect 974 2264 980 2265
rect 974 2260 975 2264
rect 979 2260 980 2264
rect 974 2259 980 2260
rect 1198 2264 1204 2265
rect 1198 2260 1199 2264
rect 1203 2260 1204 2264
rect 1198 2259 1204 2260
rect 1430 2264 1436 2265
rect 1430 2260 1431 2264
rect 1435 2260 1436 2264
rect 1430 2259 1436 2260
rect 1670 2264 1676 2265
rect 1670 2260 1671 2264
rect 1675 2260 1676 2264
rect 1934 2261 1935 2265
rect 1939 2261 1940 2265
rect 1934 2260 1940 2261
rect 1670 2259 1676 2260
rect 130 2249 136 2250
rect 110 2248 116 2249
rect 110 2244 111 2248
rect 115 2244 116 2248
rect 130 2245 131 2249
rect 135 2245 136 2249
rect 130 2244 136 2245
rect 306 2249 312 2250
rect 306 2245 307 2249
rect 311 2245 312 2249
rect 306 2244 312 2245
rect 514 2249 520 2250
rect 514 2245 515 2249
rect 519 2245 520 2249
rect 514 2244 520 2245
rect 730 2249 736 2250
rect 730 2245 731 2249
rect 735 2245 736 2249
rect 730 2244 736 2245
rect 946 2249 952 2250
rect 946 2245 947 2249
rect 951 2245 952 2249
rect 946 2244 952 2245
rect 1170 2249 1176 2250
rect 1170 2245 1171 2249
rect 1175 2245 1176 2249
rect 1170 2244 1176 2245
rect 1402 2249 1408 2250
rect 1402 2245 1403 2249
rect 1407 2245 1408 2249
rect 1402 2244 1408 2245
rect 1642 2249 1648 2250
rect 1642 2245 1643 2249
rect 1647 2245 1648 2249
rect 1642 2244 1648 2245
rect 1934 2248 1940 2249
rect 1934 2244 1935 2248
rect 1939 2244 1940 2248
rect 110 2243 116 2244
rect 112 2163 114 2243
rect 132 2163 134 2244
rect 308 2163 310 2244
rect 516 2163 518 2244
rect 732 2163 734 2244
rect 948 2163 950 2244
rect 1172 2163 1174 2244
rect 1404 2163 1406 2244
rect 1644 2163 1646 2244
rect 1934 2243 1940 2244
rect 1936 2163 1938 2243
rect 1976 2231 1978 2282
rect 2360 2231 2362 2283
rect 2568 2231 2570 2283
rect 2768 2231 2770 2283
rect 2960 2231 2962 2283
rect 3152 2231 3154 2283
rect 3336 2231 3338 2283
rect 3520 2231 3522 2283
rect 3680 2231 3682 2283
rect 3798 2282 3804 2283
rect 3800 2231 3802 2282
rect 3840 2270 3842 2293
rect 3838 2269 3844 2270
rect 3888 2269 3890 2293
rect 4072 2269 4074 2293
rect 4272 2269 4274 2293
rect 4464 2269 4466 2293
rect 4656 2269 4658 2293
rect 4840 2269 4842 2293
rect 5016 2269 5018 2293
rect 5184 2269 5186 2293
rect 5360 2269 5362 2293
rect 5536 2269 5538 2293
rect 5664 2270 5666 2293
rect 5662 2269 5668 2270
rect 3838 2265 3839 2269
rect 3843 2265 3844 2269
rect 3838 2264 3844 2265
rect 3886 2268 3892 2269
rect 3886 2264 3887 2268
rect 3891 2264 3892 2268
rect 3886 2263 3892 2264
rect 4070 2268 4076 2269
rect 4070 2264 4071 2268
rect 4075 2264 4076 2268
rect 4070 2263 4076 2264
rect 4270 2268 4276 2269
rect 4270 2264 4271 2268
rect 4275 2264 4276 2268
rect 4270 2263 4276 2264
rect 4462 2268 4468 2269
rect 4462 2264 4463 2268
rect 4467 2264 4468 2268
rect 4462 2263 4468 2264
rect 4654 2268 4660 2269
rect 4654 2264 4655 2268
rect 4659 2264 4660 2268
rect 4654 2263 4660 2264
rect 4838 2268 4844 2269
rect 4838 2264 4839 2268
rect 4843 2264 4844 2268
rect 4838 2263 4844 2264
rect 5014 2268 5020 2269
rect 5014 2264 5015 2268
rect 5019 2264 5020 2268
rect 5014 2263 5020 2264
rect 5182 2268 5188 2269
rect 5182 2264 5183 2268
rect 5187 2264 5188 2268
rect 5182 2263 5188 2264
rect 5358 2268 5364 2269
rect 5358 2264 5359 2268
rect 5363 2264 5364 2268
rect 5358 2263 5364 2264
rect 5534 2268 5540 2269
rect 5534 2264 5535 2268
rect 5539 2264 5540 2268
rect 5662 2265 5663 2269
rect 5667 2265 5668 2269
rect 5662 2264 5668 2265
rect 5534 2263 5540 2264
rect 3858 2253 3864 2254
rect 3838 2252 3844 2253
rect 3838 2248 3839 2252
rect 3843 2248 3844 2252
rect 3858 2249 3859 2253
rect 3863 2249 3864 2253
rect 3858 2248 3864 2249
rect 4042 2253 4048 2254
rect 4042 2249 4043 2253
rect 4047 2249 4048 2253
rect 4042 2248 4048 2249
rect 4242 2253 4248 2254
rect 4242 2249 4243 2253
rect 4247 2249 4248 2253
rect 4242 2248 4248 2249
rect 4434 2253 4440 2254
rect 4434 2249 4435 2253
rect 4439 2249 4440 2253
rect 4434 2248 4440 2249
rect 4626 2253 4632 2254
rect 4626 2249 4627 2253
rect 4631 2249 4632 2253
rect 4626 2248 4632 2249
rect 4810 2253 4816 2254
rect 4810 2249 4811 2253
rect 4815 2249 4816 2253
rect 4810 2248 4816 2249
rect 4986 2253 4992 2254
rect 4986 2249 4987 2253
rect 4991 2249 4992 2253
rect 4986 2248 4992 2249
rect 5154 2253 5160 2254
rect 5154 2249 5155 2253
rect 5159 2249 5160 2253
rect 5154 2248 5160 2249
rect 5330 2253 5336 2254
rect 5330 2249 5331 2253
rect 5335 2249 5336 2253
rect 5330 2248 5336 2249
rect 5506 2253 5512 2254
rect 5506 2249 5507 2253
rect 5511 2249 5512 2253
rect 5506 2248 5512 2249
rect 5662 2252 5668 2253
rect 5662 2248 5663 2252
rect 5667 2248 5668 2252
rect 3838 2247 3844 2248
rect 1975 2230 1979 2231
rect 1975 2225 1979 2226
rect 2359 2230 2363 2231
rect 2359 2225 2363 2226
rect 2463 2230 2467 2231
rect 2463 2225 2467 2226
rect 2567 2230 2571 2231
rect 2567 2225 2571 2226
rect 2599 2230 2603 2231
rect 2599 2225 2603 2226
rect 2735 2230 2739 2231
rect 2735 2225 2739 2226
rect 2767 2230 2771 2231
rect 2767 2225 2771 2226
rect 2959 2230 2963 2231
rect 2959 2225 2963 2226
rect 3151 2230 3155 2231
rect 3151 2225 3155 2226
rect 3335 2230 3339 2231
rect 3335 2225 3339 2226
rect 3519 2230 3523 2231
rect 3519 2225 3523 2226
rect 3679 2230 3683 2231
rect 3679 2225 3683 2226
rect 3799 2230 3803 2231
rect 3799 2225 3803 2226
rect 1976 2202 1978 2225
rect 1974 2201 1980 2202
rect 2464 2201 2466 2225
rect 2600 2201 2602 2225
rect 2736 2201 2738 2225
rect 3800 2202 3802 2225
rect 3798 2201 3804 2202
rect 1974 2197 1975 2201
rect 1979 2197 1980 2201
rect 1974 2196 1980 2197
rect 2462 2200 2468 2201
rect 2462 2196 2463 2200
rect 2467 2196 2468 2200
rect 2462 2195 2468 2196
rect 2598 2200 2604 2201
rect 2598 2196 2599 2200
rect 2603 2196 2604 2200
rect 2598 2195 2604 2196
rect 2734 2200 2740 2201
rect 2734 2196 2735 2200
rect 2739 2196 2740 2200
rect 3798 2197 3799 2201
rect 3803 2197 3804 2201
rect 3798 2196 3804 2197
rect 2734 2195 2740 2196
rect 3840 2187 3842 2247
rect 3860 2187 3862 2248
rect 4044 2187 4046 2248
rect 4244 2187 4246 2248
rect 4436 2187 4438 2248
rect 4628 2187 4630 2248
rect 4812 2187 4814 2248
rect 4988 2187 4990 2248
rect 5156 2187 5158 2248
rect 5332 2187 5334 2248
rect 5508 2187 5510 2248
rect 5662 2247 5668 2248
rect 5664 2187 5666 2247
rect 3839 2186 3843 2187
rect 2434 2185 2440 2186
rect 1974 2184 1980 2185
rect 1974 2180 1975 2184
rect 1979 2180 1980 2184
rect 2434 2181 2435 2185
rect 2439 2181 2440 2185
rect 2434 2180 2440 2181
rect 2570 2185 2576 2186
rect 2570 2181 2571 2185
rect 2575 2181 2576 2185
rect 2570 2180 2576 2181
rect 2706 2185 2712 2186
rect 2706 2181 2707 2185
rect 2711 2181 2712 2185
rect 2706 2180 2712 2181
rect 3798 2184 3804 2185
rect 3798 2180 3799 2184
rect 3803 2180 3804 2184
rect 3839 2181 3843 2182
rect 3859 2186 3863 2187
rect 3859 2181 3863 2182
rect 4043 2186 4047 2187
rect 4043 2181 4047 2182
rect 4243 2186 4247 2187
rect 4243 2181 4247 2182
rect 4251 2186 4255 2187
rect 4251 2181 4255 2182
rect 4435 2186 4439 2187
rect 4435 2181 4439 2182
rect 4459 2186 4463 2187
rect 4459 2181 4463 2182
rect 4627 2186 4631 2187
rect 4627 2181 4631 2182
rect 4659 2186 4663 2187
rect 4659 2181 4663 2182
rect 4811 2186 4815 2187
rect 4811 2181 4815 2182
rect 4851 2186 4855 2187
rect 4851 2181 4855 2182
rect 4987 2186 4991 2187
rect 4987 2181 4991 2182
rect 5035 2186 5039 2187
rect 5035 2181 5039 2182
rect 5155 2186 5159 2187
rect 5155 2181 5159 2182
rect 5219 2186 5223 2187
rect 5219 2181 5223 2182
rect 5331 2186 5335 2187
rect 5331 2181 5335 2182
rect 5411 2186 5415 2187
rect 5411 2181 5415 2182
rect 5507 2186 5511 2187
rect 5507 2181 5511 2182
rect 5663 2186 5667 2187
rect 5663 2181 5667 2182
rect 1974 2179 1980 2180
rect 111 2162 115 2163
rect 111 2157 115 2158
rect 131 2162 135 2163
rect 131 2157 135 2158
rect 299 2162 303 2163
rect 299 2157 303 2158
rect 307 2162 311 2163
rect 307 2157 311 2158
rect 499 2162 503 2163
rect 499 2157 503 2158
rect 515 2162 519 2163
rect 515 2157 519 2158
rect 715 2162 719 2163
rect 715 2157 719 2158
rect 731 2162 735 2163
rect 731 2157 735 2158
rect 931 2162 935 2163
rect 931 2157 935 2158
rect 947 2162 951 2163
rect 947 2157 951 2158
rect 1155 2162 1159 2163
rect 1155 2157 1159 2158
rect 1171 2162 1175 2163
rect 1171 2157 1175 2158
rect 1387 2162 1391 2163
rect 1387 2157 1391 2158
rect 1403 2162 1407 2163
rect 1403 2157 1407 2158
rect 1627 2162 1631 2163
rect 1627 2157 1631 2158
rect 1643 2162 1647 2163
rect 1643 2157 1647 2158
rect 1935 2162 1939 2163
rect 1935 2157 1939 2158
rect 112 2097 114 2157
rect 110 2096 116 2097
rect 132 2096 134 2157
rect 300 2096 302 2157
rect 500 2096 502 2157
rect 716 2096 718 2157
rect 932 2096 934 2157
rect 1156 2096 1158 2157
rect 1388 2096 1390 2157
rect 1628 2096 1630 2157
rect 1936 2097 1938 2157
rect 1934 2096 1940 2097
rect 110 2092 111 2096
rect 115 2092 116 2096
rect 110 2091 116 2092
rect 130 2095 136 2096
rect 130 2091 131 2095
rect 135 2091 136 2095
rect 130 2090 136 2091
rect 298 2095 304 2096
rect 298 2091 299 2095
rect 303 2091 304 2095
rect 298 2090 304 2091
rect 498 2095 504 2096
rect 498 2091 499 2095
rect 503 2091 504 2095
rect 498 2090 504 2091
rect 714 2095 720 2096
rect 714 2091 715 2095
rect 719 2091 720 2095
rect 714 2090 720 2091
rect 930 2095 936 2096
rect 930 2091 931 2095
rect 935 2091 936 2095
rect 930 2090 936 2091
rect 1154 2095 1160 2096
rect 1154 2091 1155 2095
rect 1159 2091 1160 2095
rect 1154 2090 1160 2091
rect 1386 2095 1392 2096
rect 1386 2091 1387 2095
rect 1391 2091 1392 2095
rect 1386 2090 1392 2091
rect 1626 2095 1632 2096
rect 1626 2091 1627 2095
rect 1631 2091 1632 2095
rect 1934 2092 1935 2096
rect 1939 2092 1940 2096
rect 1934 2091 1940 2092
rect 1626 2090 1632 2091
rect 1976 2087 1978 2179
rect 2436 2087 2438 2180
rect 2572 2087 2574 2180
rect 2708 2087 2710 2180
rect 3798 2179 3804 2180
rect 3800 2087 3802 2179
rect 3840 2121 3842 2181
rect 3838 2120 3844 2121
rect 3860 2120 3862 2181
rect 4044 2120 4046 2181
rect 4252 2120 4254 2181
rect 4460 2120 4462 2181
rect 4660 2120 4662 2181
rect 4852 2120 4854 2181
rect 5036 2120 5038 2181
rect 5220 2120 5222 2181
rect 5412 2120 5414 2181
rect 5664 2121 5666 2181
rect 5662 2120 5668 2121
rect 3838 2116 3839 2120
rect 3843 2116 3844 2120
rect 3838 2115 3844 2116
rect 3858 2119 3864 2120
rect 3858 2115 3859 2119
rect 3863 2115 3864 2119
rect 3858 2114 3864 2115
rect 4042 2119 4048 2120
rect 4042 2115 4043 2119
rect 4047 2115 4048 2119
rect 4042 2114 4048 2115
rect 4250 2119 4256 2120
rect 4250 2115 4251 2119
rect 4255 2115 4256 2119
rect 4250 2114 4256 2115
rect 4458 2119 4464 2120
rect 4458 2115 4459 2119
rect 4463 2115 4464 2119
rect 4458 2114 4464 2115
rect 4658 2119 4664 2120
rect 4658 2115 4659 2119
rect 4663 2115 4664 2119
rect 4658 2114 4664 2115
rect 4850 2119 4856 2120
rect 4850 2115 4851 2119
rect 4855 2115 4856 2119
rect 4850 2114 4856 2115
rect 5034 2119 5040 2120
rect 5034 2115 5035 2119
rect 5039 2115 5040 2119
rect 5034 2114 5040 2115
rect 5218 2119 5224 2120
rect 5218 2115 5219 2119
rect 5223 2115 5224 2119
rect 5218 2114 5224 2115
rect 5410 2119 5416 2120
rect 5410 2115 5411 2119
rect 5415 2115 5416 2119
rect 5662 2116 5663 2120
rect 5667 2116 5668 2120
rect 5662 2115 5668 2116
rect 5410 2114 5416 2115
rect 3886 2104 3892 2105
rect 3838 2103 3844 2104
rect 3838 2099 3839 2103
rect 3843 2099 3844 2103
rect 3886 2100 3887 2104
rect 3891 2100 3892 2104
rect 3886 2099 3892 2100
rect 4070 2104 4076 2105
rect 4070 2100 4071 2104
rect 4075 2100 4076 2104
rect 4070 2099 4076 2100
rect 4278 2104 4284 2105
rect 4278 2100 4279 2104
rect 4283 2100 4284 2104
rect 4278 2099 4284 2100
rect 4486 2104 4492 2105
rect 4486 2100 4487 2104
rect 4491 2100 4492 2104
rect 4486 2099 4492 2100
rect 4686 2104 4692 2105
rect 4686 2100 4687 2104
rect 4691 2100 4692 2104
rect 4686 2099 4692 2100
rect 4878 2104 4884 2105
rect 4878 2100 4879 2104
rect 4883 2100 4884 2104
rect 4878 2099 4884 2100
rect 5062 2104 5068 2105
rect 5062 2100 5063 2104
rect 5067 2100 5068 2104
rect 5062 2099 5068 2100
rect 5246 2104 5252 2105
rect 5246 2100 5247 2104
rect 5251 2100 5252 2104
rect 5246 2099 5252 2100
rect 5438 2104 5444 2105
rect 5438 2100 5439 2104
rect 5443 2100 5444 2104
rect 5438 2099 5444 2100
rect 5662 2103 5668 2104
rect 5662 2099 5663 2103
rect 5667 2099 5668 2103
rect 3838 2098 3844 2099
rect 1975 2086 1979 2087
rect 1975 2081 1979 2082
rect 2419 2086 2423 2087
rect 2419 2081 2423 2082
rect 2435 2086 2439 2087
rect 2435 2081 2439 2082
rect 2571 2086 2575 2087
rect 2571 2081 2575 2082
rect 2611 2086 2615 2087
rect 2611 2081 2615 2082
rect 2707 2086 2711 2087
rect 2707 2081 2711 2082
rect 2795 2086 2799 2087
rect 2795 2081 2799 2082
rect 2979 2086 2983 2087
rect 2979 2081 2983 2082
rect 3155 2086 3159 2087
rect 3155 2081 3159 2082
rect 3323 2086 3327 2087
rect 3323 2081 3327 2082
rect 3499 2086 3503 2087
rect 3499 2081 3503 2082
rect 3651 2086 3655 2087
rect 3651 2081 3655 2082
rect 3799 2086 3803 2087
rect 3799 2081 3803 2082
rect 158 2080 164 2081
rect 110 2079 116 2080
rect 110 2075 111 2079
rect 115 2075 116 2079
rect 158 2076 159 2080
rect 163 2076 164 2080
rect 158 2075 164 2076
rect 326 2080 332 2081
rect 326 2076 327 2080
rect 331 2076 332 2080
rect 326 2075 332 2076
rect 526 2080 532 2081
rect 526 2076 527 2080
rect 531 2076 532 2080
rect 526 2075 532 2076
rect 742 2080 748 2081
rect 742 2076 743 2080
rect 747 2076 748 2080
rect 742 2075 748 2076
rect 958 2080 964 2081
rect 958 2076 959 2080
rect 963 2076 964 2080
rect 958 2075 964 2076
rect 1182 2080 1188 2081
rect 1182 2076 1183 2080
rect 1187 2076 1188 2080
rect 1182 2075 1188 2076
rect 1414 2080 1420 2081
rect 1414 2076 1415 2080
rect 1419 2076 1420 2080
rect 1414 2075 1420 2076
rect 1654 2080 1660 2081
rect 1654 2076 1655 2080
rect 1659 2076 1660 2080
rect 1654 2075 1660 2076
rect 1934 2079 1940 2080
rect 1934 2075 1935 2079
rect 1939 2075 1940 2079
rect 110 2074 116 2075
rect 112 2043 114 2074
rect 160 2043 162 2075
rect 328 2043 330 2075
rect 528 2043 530 2075
rect 744 2043 746 2075
rect 960 2043 962 2075
rect 1184 2043 1186 2075
rect 1416 2043 1418 2075
rect 1656 2043 1658 2075
rect 1934 2074 1940 2075
rect 1936 2043 1938 2074
rect 111 2042 115 2043
rect 111 2037 115 2038
rect 159 2042 163 2043
rect 159 2037 163 2038
rect 327 2042 331 2043
rect 327 2037 331 2038
rect 343 2042 347 2043
rect 343 2037 347 2038
rect 527 2042 531 2043
rect 527 2037 531 2038
rect 567 2042 571 2043
rect 567 2037 571 2038
rect 743 2042 747 2043
rect 743 2037 747 2038
rect 807 2042 811 2043
rect 807 2037 811 2038
rect 959 2042 963 2043
rect 959 2037 963 2038
rect 1063 2042 1067 2043
rect 1063 2037 1067 2038
rect 1183 2042 1187 2043
rect 1183 2037 1187 2038
rect 1335 2042 1339 2043
rect 1335 2037 1339 2038
rect 1415 2042 1419 2043
rect 1415 2037 1419 2038
rect 1607 2042 1611 2043
rect 1607 2037 1611 2038
rect 1655 2042 1659 2043
rect 1655 2037 1659 2038
rect 1935 2042 1939 2043
rect 1935 2037 1939 2038
rect 112 2014 114 2037
rect 110 2013 116 2014
rect 160 2013 162 2037
rect 344 2013 346 2037
rect 568 2013 570 2037
rect 808 2013 810 2037
rect 1064 2013 1066 2037
rect 1336 2013 1338 2037
rect 1608 2013 1610 2037
rect 1936 2014 1938 2037
rect 1976 2021 1978 2081
rect 1974 2020 1980 2021
rect 2420 2020 2422 2081
rect 2612 2020 2614 2081
rect 2796 2020 2798 2081
rect 2980 2020 2982 2081
rect 3156 2020 3158 2081
rect 3324 2020 3326 2081
rect 3500 2020 3502 2081
rect 3652 2020 3654 2081
rect 3800 2021 3802 2081
rect 3840 2055 3842 2098
rect 3888 2055 3890 2099
rect 4072 2055 4074 2099
rect 4280 2055 4282 2099
rect 4488 2055 4490 2099
rect 4688 2055 4690 2099
rect 4880 2055 4882 2099
rect 5064 2055 5066 2099
rect 5248 2055 5250 2099
rect 5440 2055 5442 2099
rect 5662 2098 5668 2099
rect 5664 2055 5666 2098
rect 3839 2054 3843 2055
rect 3839 2049 3843 2050
rect 3887 2054 3891 2055
rect 3887 2049 3891 2050
rect 4071 2054 4075 2055
rect 4071 2049 4075 2050
rect 4279 2054 4283 2055
rect 4279 2049 4283 2050
rect 4287 2054 4291 2055
rect 4287 2049 4291 2050
rect 4423 2054 4427 2055
rect 4423 2049 4427 2050
rect 4487 2054 4491 2055
rect 4487 2049 4491 2050
rect 4559 2054 4563 2055
rect 4559 2049 4563 2050
rect 4687 2054 4691 2055
rect 4687 2049 4691 2050
rect 4695 2054 4699 2055
rect 4695 2049 4699 2050
rect 4839 2054 4843 2055
rect 4839 2049 4843 2050
rect 4879 2054 4883 2055
rect 4879 2049 4883 2050
rect 5063 2054 5067 2055
rect 5063 2049 5067 2050
rect 5247 2054 5251 2055
rect 5247 2049 5251 2050
rect 5439 2054 5443 2055
rect 5439 2049 5443 2050
rect 5663 2054 5667 2055
rect 5663 2049 5667 2050
rect 3840 2026 3842 2049
rect 3838 2025 3844 2026
rect 4288 2025 4290 2049
rect 4424 2025 4426 2049
rect 4560 2025 4562 2049
rect 4696 2025 4698 2049
rect 4840 2025 4842 2049
rect 5664 2026 5666 2049
rect 5662 2025 5668 2026
rect 3838 2021 3839 2025
rect 3843 2021 3844 2025
rect 3798 2020 3804 2021
rect 3838 2020 3844 2021
rect 4286 2024 4292 2025
rect 4286 2020 4287 2024
rect 4291 2020 4292 2024
rect 1974 2016 1975 2020
rect 1979 2016 1980 2020
rect 1974 2015 1980 2016
rect 2418 2019 2424 2020
rect 2418 2015 2419 2019
rect 2423 2015 2424 2019
rect 2418 2014 2424 2015
rect 2610 2019 2616 2020
rect 2610 2015 2611 2019
rect 2615 2015 2616 2019
rect 2610 2014 2616 2015
rect 2794 2019 2800 2020
rect 2794 2015 2795 2019
rect 2799 2015 2800 2019
rect 2794 2014 2800 2015
rect 2978 2019 2984 2020
rect 2978 2015 2979 2019
rect 2983 2015 2984 2019
rect 2978 2014 2984 2015
rect 3154 2019 3160 2020
rect 3154 2015 3155 2019
rect 3159 2015 3160 2019
rect 3154 2014 3160 2015
rect 3322 2019 3328 2020
rect 3322 2015 3323 2019
rect 3327 2015 3328 2019
rect 3322 2014 3328 2015
rect 3498 2019 3504 2020
rect 3498 2015 3499 2019
rect 3503 2015 3504 2019
rect 3498 2014 3504 2015
rect 3650 2019 3656 2020
rect 3650 2015 3651 2019
rect 3655 2015 3656 2019
rect 3798 2016 3799 2020
rect 3803 2016 3804 2020
rect 4286 2019 4292 2020
rect 4422 2024 4428 2025
rect 4422 2020 4423 2024
rect 4427 2020 4428 2024
rect 4422 2019 4428 2020
rect 4558 2024 4564 2025
rect 4558 2020 4559 2024
rect 4563 2020 4564 2024
rect 4558 2019 4564 2020
rect 4694 2024 4700 2025
rect 4694 2020 4695 2024
rect 4699 2020 4700 2024
rect 4694 2019 4700 2020
rect 4838 2024 4844 2025
rect 4838 2020 4839 2024
rect 4843 2020 4844 2024
rect 5662 2021 5663 2025
rect 5667 2021 5668 2025
rect 5662 2020 5668 2021
rect 4838 2019 4844 2020
rect 3798 2015 3804 2016
rect 3650 2014 3656 2015
rect 1934 2013 1940 2014
rect 110 2009 111 2013
rect 115 2009 116 2013
rect 110 2008 116 2009
rect 158 2012 164 2013
rect 158 2008 159 2012
rect 163 2008 164 2012
rect 158 2007 164 2008
rect 342 2012 348 2013
rect 342 2008 343 2012
rect 347 2008 348 2012
rect 342 2007 348 2008
rect 566 2012 572 2013
rect 566 2008 567 2012
rect 571 2008 572 2012
rect 566 2007 572 2008
rect 806 2012 812 2013
rect 806 2008 807 2012
rect 811 2008 812 2012
rect 806 2007 812 2008
rect 1062 2012 1068 2013
rect 1062 2008 1063 2012
rect 1067 2008 1068 2012
rect 1062 2007 1068 2008
rect 1334 2012 1340 2013
rect 1334 2008 1335 2012
rect 1339 2008 1340 2012
rect 1334 2007 1340 2008
rect 1606 2012 1612 2013
rect 1606 2008 1607 2012
rect 1611 2008 1612 2012
rect 1934 2009 1935 2013
rect 1939 2009 1940 2013
rect 4258 2009 4264 2010
rect 1934 2008 1940 2009
rect 3838 2008 3844 2009
rect 1606 2007 1612 2008
rect 2446 2004 2452 2005
rect 1974 2003 1980 2004
rect 1974 1999 1975 2003
rect 1979 1999 1980 2003
rect 2446 2000 2447 2004
rect 2451 2000 2452 2004
rect 2446 1999 2452 2000
rect 2638 2004 2644 2005
rect 2638 2000 2639 2004
rect 2643 2000 2644 2004
rect 2638 1999 2644 2000
rect 2822 2004 2828 2005
rect 2822 2000 2823 2004
rect 2827 2000 2828 2004
rect 2822 1999 2828 2000
rect 3006 2004 3012 2005
rect 3006 2000 3007 2004
rect 3011 2000 3012 2004
rect 3006 1999 3012 2000
rect 3182 2004 3188 2005
rect 3182 2000 3183 2004
rect 3187 2000 3188 2004
rect 3182 1999 3188 2000
rect 3350 2004 3356 2005
rect 3350 2000 3351 2004
rect 3355 2000 3356 2004
rect 3350 1999 3356 2000
rect 3526 2004 3532 2005
rect 3526 2000 3527 2004
rect 3531 2000 3532 2004
rect 3526 1999 3532 2000
rect 3678 2004 3684 2005
rect 3838 2004 3839 2008
rect 3843 2004 3844 2008
rect 4258 2005 4259 2009
rect 4263 2005 4264 2009
rect 4258 2004 4264 2005
rect 4394 2009 4400 2010
rect 4394 2005 4395 2009
rect 4399 2005 4400 2009
rect 4394 2004 4400 2005
rect 4530 2009 4536 2010
rect 4530 2005 4531 2009
rect 4535 2005 4536 2009
rect 4530 2004 4536 2005
rect 4666 2009 4672 2010
rect 4666 2005 4667 2009
rect 4671 2005 4672 2009
rect 4666 2004 4672 2005
rect 4810 2009 4816 2010
rect 4810 2005 4811 2009
rect 4815 2005 4816 2009
rect 4810 2004 4816 2005
rect 5662 2008 5668 2009
rect 5662 2004 5663 2008
rect 5667 2004 5668 2008
rect 3678 2000 3679 2004
rect 3683 2000 3684 2004
rect 3678 1999 3684 2000
rect 3798 2003 3804 2004
rect 3838 2003 3844 2004
rect 3798 1999 3799 2003
rect 3803 1999 3804 2003
rect 1974 1998 1980 1999
rect 130 1997 136 1998
rect 110 1996 116 1997
rect 110 1992 111 1996
rect 115 1992 116 1996
rect 130 1993 131 1997
rect 135 1993 136 1997
rect 130 1992 136 1993
rect 314 1997 320 1998
rect 314 1993 315 1997
rect 319 1993 320 1997
rect 314 1992 320 1993
rect 538 1997 544 1998
rect 538 1993 539 1997
rect 543 1993 544 1997
rect 538 1992 544 1993
rect 778 1997 784 1998
rect 778 1993 779 1997
rect 783 1993 784 1997
rect 778 1992 784 1993
rect 1034 1997 1040 1998
rect 1034 1993 1035 1997
rect 1039 1993 1040 1997
rect 1034 1992 1040 1993
rect 1306 1997 1312 1998
rect 1306 1993 1307 1997
rect 1311 1993 1312 1997
rect 1306 1992 1312 1993
rect 1578 1997 1584 1998
rect 1578 1993 1579 1997
rect 1583 1993 1584 1997
rect 1578 1992 1584 1993
rect 1934 1996 1940 1997
rect 1934 1992 1935 1996
rect 1939 1992 1940 1996
rect 110 1991 116 1992
rect 112 1927 114 1991
rect 132 1927 134 1992
rect 316 1927 318 1992
rect 540 1927 542 1992
rect 780 1927 782 1992
rect 1036 1927 1038 1992
rect 1308 1927 1310 1992
rect 1580 1927 1582 1992
rect 1934 1991 1940 1992
rect 1936 1927 1938 1991
rect 1976 1963 1978 1998
rect 2448 1963 2450 1999
rect 2640 1963 2642 1999
rect 2824 1963 2826 1999
rect 3008 1963 3010 1999
rect 3184 1963 3186 1999
rect 3352 1963 3354 1999
rect 3528 1963 3530 1999
rect 3680 1963 3682 1999
rect 3798 1998 3804 1999
rect 3800 1963 3802 1998
rect 1975 1962 1979 1963
rect 1975 1957 1979 1958
rect 2359 1962 2363 1963
rect 2359 1957 2363 1958
rect 2447 1962 2451 1963
rect 2447 1957 2451 1958
rect 2495 1962 2499 1963
rect 2495 1957 2499 1958
rect 2631 1962 2635 1963
rect 2631 1957 2635 1958
rect 2639 1962 2643 1963
rect 2639 1957 2643 1958
rect 2767 1962 2771 1963
rect 2767 1957 2771 1958
rect 2823 1962 2827 1963
rect 2823 1957 2827 1958
rect 2903 1962 2907 1963
rect 2903 1957 2907 1958
rect 3007 1962 3011 1963
rect 3007 1957 3011 1958
rect 3039 1962 3043 1963
rect 3039 1957 3043 1958
rect 3175 1962 3179 1963
rect 3175 1957 3179 1958
rect 3183 1962 3187 1963
rect 3183 1957 3187 1958
rect 3319 1962 3323 1963
rect 3319 1957 3323 1958
rect 3351 1962 3355 1963
rect 3351 1957 3355 1958
rect 3527 1962 3531 1963
rect 3527 1957 3531 1958
rect 3679 1962 3683 1963
rect 3679 1957 3683 1958
rect 3799 1962 3803 1963
rect 3799 1957 3803 1958
rect 1976 1934 1978 1957
rect 1974 1933 1980 1934
rect 2360 1933 2362 1957
rect 2496 1933 2498 1957
rect 2632 1933 2634 1957
rect 2768 1933 2770 1957
rect 2904 1933 2906 1957
rect 3040 1933 3042 1957
rect 3176 1933 3178 1957
rect 3320 1933 3322 1957
rect 3800 1934 3802 1957
rect 3798 1933 3804 1934
rect 1974 1929 1975 1933
rect 1979 1929 1980 1933
rect 1974 1928 1980 1929
rect 2358 1932 2364 1933
rect 2358 1928 2359 1932
rect 2363 1928 2364 1932
rect 2358 1927 2364 1928
rect 2494 1932 2500 1933
rect 2494 1928 2495 1932
rect 2499 1928 2500 1932
rect 2494 1927 2500 1928
rect 2630 1932 2636 1933
rect 2630 1928 2631 1932
rect 2635 1928 2636 1932
rect 2630 1927 2636 1928
rect 2766 1932 2772 1933
rect 2766 1928 2767 1932
rect 2771 1928 2772 1932
rect 2766 1927 2772 1928
rect 2902 1932 2908 1933
rect 2902 1928 2903 1932
rect 2907 1928 2908 1932
rect 2902 1927 2908 1928
rect 3038 1932 3044 1933
rect 3038 1928 3039 1932
rect 3043 1928 3044 1932
rect 3038 1927 3044 1928
rect 3174 1932 3180 1933
rect 3174 1928 3175 1932
rect 3179 1928 3180 1932
rect 3174 1927 3180 1928
rect 3318 1932 3324 1933
rect 3318 1928 3319 1932
rect 3323 1928 3324 1932
rect 3798 1929 3799 1933
rect 3803 1929 3804 1933
rect 3798 1928 3804 1929
rect 3318 1927 3324 1928
rect 111 1926 115 1927
rect 111 1921 115 1922
rect 131 1926 135 1927
rect 131 1921 135 1922
rect 315 1926 319 1927
rect 315 1921 319 1922
rect 331 1926 335 1927
rect 331 1921 335 1922
rect 499 1926 503 1927
rect 499 1921 503 1922
rect 539 1926 543 1927
rect 539 1921 543 1922
rect 667 1926 671 1927
rect 667 1921 671 1922
rect 779 1926 783 1927
rect 779 1921 783 1922
rect 843 1926 847 1927
rect 843 1921 847 1922
rect 1027 1926 1031 1927
rect 1027 1921 1031 1922
rect 1035 1926 1039 1927
rect 1035 1921 1039 1922
rect 1219 1926 1223 1927
rect 1219 1921 1223 1922
rect 1307 1926 1311 1927
rect 1307 1921 1311 1922
rect 1411 1926 1415 1927
rect 1411 1921 1415 1922
rect 1579 1926 1583 1927
rect 1579 1921 1583 1922
rect 1603 1926 1607 1927
rect 1603 1921 1607 1922
rect 1935 1926 1939 1927
rect 3840 1923 3842 2003
rect 4260 1923 4262 2004
rect 4396 1923 4398 2004
rect 4532 1923 4534 2004
rect 4668 1923 4670 2004
rect 4812 1923 4814 2004
rect 5662 2003 5668 2004
rect 5664 1923 5666 2003
rect 1935 1921 1939 1922
rect 3839 1922 3843 1923
rect 112 1861 114 1921
rect 110 1860 116 1861
rect 332 1860 334 1921
rect 500 1860 502 1921
rect 668 1860 670 1921
rect 844 1860 846 1921
rect 1028 1860 1030 1921
rect 1220 1860 1222 1921
rect 1412 1860 1414 1921
rect 1604 1860 1606 1921
rect 1936 1861 1938 1921
rect 2330 1917 2336 1918
rect 1974 1916 1980 1917
rect 1974 1912 1975 1916
rect 1979 1912 1980 1916
rect 2330 1913 2331 1917
rect 2335 1913 2336 1917
rect 2330 1912 2336 1913
rect 2466 1917 2472 1918
rect 2466 1913 2467 1917
rect 2471 1913 2472 1917
rect 2466 1912 2472 1913
rect 2602 1917 2608 1918
rect 2602 1913 2603 1917
rect 2607 1913 2608 1917
rect 2602 1912 2608 1913
rect 2738 1917 2744 1918
rect 2738 1913 2739 1917
rect 2743 1913 2744 1917
rect 2738 1912 2744 1913
rect 2874 1917 2880 1918
rect 2874 1913 2875 1917
rect 2879 1913 2880 1917
rect 2874 1912 2880 1913
rect 3010 1917 3016 1918
rect 3010 1913 3011 1917
rect 3015 1913 3016 1917
rect 3010 1912 3016 1913
rect 3146 1917 3152 1918
rect 3146 1913 3147 1917
rect 3151 1913 3152 1917
rect 3146 1912 3152 1913
rect 3290 1917 3296 1918
rect 3839 1917 3843 1918
rect 3955 1922 3959 1923
rect 3955 1917 3959 1918
rect 4195 1922 4199 1923
rect 4195 1917 4199 1918
rect 4259 1922 4263 1923
rect 4259 1917 4263 1918
rect 4395 1922 4399 1923
rect 4395 1917 4399 1918
rect 4467 1922 4471 1923
rect 4467 1917 4471 1918
rect 4531 1922 4535 1923
rect 4531 1917 4535 1918
rect 4667 1922 4671 1923
rect 4667 1917 4671 1918
rect 4771 1922 4775 1923
rect 4771 1917 4775 1918
rect 4811 1922 4815 1923
rect 4811 1917 4815 1918
rect 5091 1922 5095 1923
rect 5091 1917 5095 1918
rect 5411 1922 5415 1923
rect 5411 1917 5415 1918
rect 5663 1922 5667 1923
rect 5663 1917 5667 1918
rect 3290 1913 3291 1917
rect 3295 1913 3296 1917
rect 3290 1912 3296 1913
rect 3798 1916 3804 1917
rect 3798 1912 3799 1916
rect 3803 1912 3804 1916
rect 1974 1911 1980 1912
rect 1934 1860 1940 1861
rect 110 1856 111 1860
rect 115 1856 116 1860
rect 110 1855 116 1856
rect 330 1859 336 1860
rect 330 1855 331 1859
rect 335 1855 336 1859
rect 330 1854 336 1855
rect 498 1859 504 1860
rect 498 1855 499 1859
rect 503 1855 504 1859
rect 498 1854 504 1855
rect 666 1859 672 1860
rect 666 1855 667 1859
rect 671 1855 672 1859
rect 666 1854 672 1855
rect 842 1859 848 1860
rect 842 1855 843 1859
rect 847 1855 848 1859
rect 842 1854 848 1855
rect 1026 1859 1032 1860
rect 1026 1855 1027 1859
rect 1031 1855 1032 1859
rect 1026 1854 1032 1855
rect 1218 1859 1224 1860
rect 1218 1855 1219 1859
rect 1223 1855 1224 1859
rect 1218 1854 1224 1855
rect 1410 1859 1416 1860
rect 1410 1855 1411 1859
rect 1415 1855 1416 1859
rect 1410 1854 1416 1855
rect 1602 1859 1608 1860
rect 1602 1855 1603 1859
rect 1607 1855 1608 1859
rect 1934 1856 1935 1860
rect 1939 1856 1940 1860
rect 1934 1855 1940 1856
rect 1602 1854 1608 1855
rect 1976 1851 1978 1911
rect 2332 1851 2334 1912
rect 2468 1851 2470 1912
rect 2604 1851 2606 1912
rect 2740 1851 2742 1912
rect 2876 1851 2878 1912
rect 3012 1851 3014 1912
rect 3148 1851 3150 1912
rect 3292 1851 3294 1912
rect 3798 1911 3804 1912
rect 3800 1851 3802 1911
rect 3840 1857 3842 1917
rect 3838 1856 3844 1857
rect 3956 1856 3958 1917
rect 4196 1856 4198 1917
rect 4468 1856 4470 1917
rect 4772 1856 4774 1917
rect 5092 1856 5094 1917
rect 5412 1856 5414 1917
rect 5664 1857 5666 1917
rect 5662 1856 5668 1857
rect 3838 1852 3839 1856
rect 3843 1852 3844 1856
rect 3838 1851 3844 1852
rect 3954 1855 3960 1856
rect 3954 1851 3955 1855
rect 3959 1851 3960 1855
rect 1975 1850 1979 1851
rect 1975 1845 1979 1846
rect 2211 1850 2215 1851
rect 2211 1845 2215 1846
rect 2331 1850 2335 1851
rect 2331 1845 2335 1846
rect 2355 1850 2359 1851
rect 2355 1845 2359 1846
rect 2467 1850 2471 1851
rect 2467 1845 2471 1846
rect 2499 1850 2503 1851
rect 2499 1845 2503 1846
rect 2603 1850 2607 1851
rect 2603 1845 2607 1846
rect 2643 1850 2647 1851
rect 2643 1845 2647 1846
rect 2739 1850 2743 1851
rect 2739 1845 2743 1846
rect 2787 1850 2791 1851
rect 2787 1845 2791 1846
rect 2875 1850 2879 1851
rect 2875 1845 2879 1846
rect 2931 1850 2935 1851
rect 2931 1845 2935 1846
rect 3011 1850 3015 1851
rect 3011 1845 3015 1846
rect 3083 1850 3087 1851
rect 3083 1845 3087 1846
rect 3147 1850 3151 1851
rect 3147 1845 3151 1846
rect 3291 1850 3295 1851
rect 3291 1845 3295 1846
rect 3799 1850 3803 1851
rect 3954 1850 3960 1851
rect 4194 1855 4200 1856
rect 4194 1851 4195 1855
rect 4199 1851 4200 1855
rect 4194 1850 4200 1851
rect 4466 1855 4472 1856
rect 4466 1851 4467 1855
rect 4471 1851 4472 1855
rect 4466 1850 4472 1851
rect 4770 1855 4776 1856
rect 4770 1851 4771 1855
rect 4775 1851 4776 1855
rect 4770 1850 4776 1851
rect 5090 1855 5096 1856
rect 5090 1851 5091 1855
rect 5095 1851 5096 1855
rect 5090 1850 5096 1851
rect 5410 1855 5416 1856
rect 5410 1851 5411 1855
rect 5415 1851 5416 1855
rect 5662 1852 5663 1856
rect 5667 1852 5668 1856
rect 5662 1851 5668 1852
rect 5410 1850 5416 1851
rect 3799 1845 3803 1846
rect 358 1844 364 1845
rect 110 1843 116 1844
rect 110 1839 111 1843
rect 115 1839 116 1843
rect 358 1840 359 1844
rect 363 1840 364 1844
rect 358 1839 364 1840
rect 526 1844 532 1845
rect 526 1840 527 1844
rect 531 1840 532 1844
rect 526 1839 532 1840
rect 694 1844 700 1845
rect 694 1840 695 1844
rect 699 1840 700 1844
rect 694 1839 700 1840
rect 870 1844 876 1845
rect 870 1840 871 1844
rect 875 1840 876 1844
rect 870 1839 876 1840
rect 1054 1844 1060 1845
rect 1054 1840 1055 1844
rect 1059 1840 1060 1844
rect 1054 1839 1060 1840
rect 1246 1844 1252 1845
rect 1246 1840 1247 1844
rect 1251 1840 1252 1844
rect 1246 1839 1252 1840
rect 1438 1844 1444 1845
rect 1438 1840 1439 1844
rect 1443 1840 1444 1844
rect 1438 1839 1444 1840
rect 1630 1844 1636 1845
rect 1630 1840 1631 1844
rect 1635 1840 1636 1844
rect 1630 1839 1636 1840
rect 1934 1843 1940 1844
rect 1934 1839 1935 1843
rect 1939 1839 1940 1843
rect 110 1838 116 1839
rect 112 1803 114 1838
rect 360 1803 362 1839
rect 528 1803 530 1839
rect 696 1803 698 1839
rect 872 1803 874 1839
rect 1056 1803 1058 1839
rect 1248 1803 1250 1839
rect 1440 1803 1442 1839
rect 1632 1803 1634 1839
rect 1934 1838 1940 1839
rect 1936 1803 1938 1838
rect 111 1802 115 1803
rect 111 1797 115 1798
rect 359 1802 363 1803
rect 359 1797 363 1798
rect 527 1802 531 1803
rect 527 1797 531 1798
rect 535 1802 539 1803
rect 535 1797 539 1798
rect 695 1802 699 1803
rect 695 1797 699 1798
rect 855 1802 859 1803
rect 855 1797 859 1798
rect 871 1802 875 1803
rect 871 1797 875 1798
rect 1015 1802 1019 1803
rect 1015 1797 1019 1798
rect 1055 1802 1059 1803
rect 1055 1797 1059 1798
rect 1183 1802 1187 1803
rect 1183 1797 1187 1798
rect 1247 1802 1251 1803
rect 1247 1797 1251 1798
rect 1351 1802 1355 1803
rect 1351 1797 1355 1798
rect 1439 1802 1443 1803
rect 1439 1797 1443 1798
rect 1519 1802 1523 1803
rect 1519 1797 1523 1798
rect 1631 1802 1635 1803
rect 1631 1797 1635 1798
rect 1935 1802 1939 1803
rect 1935 1797 1939 1798
rect 112 1774 114 1797
rect 110 1773 116 1774
rect 536 1773 538 1797
rect 696 1773 698 1797
rect 856 1773 858 1797
rect 1016 1773 1018 1797
rect 1184 1773 1186 1797
rect 1352 1773 1354 1797
rect 1520 1773 1522 1797
rect 1936 1774 1938 1797
rect 1976 1785 1978 1845
rect 1974 1784 1980 1785
rect 2212 1784 2214 1845
rect 2356 1784 2358 1845
rect 2500 1784 2502 1845
rect 2644 1784 2646 1845
rect 2788 1784 2790 1845
rect 2932 1784 2934 1845
rect 3084 1784 3086 1845
rect 3800 1785 3802 1845
rect 3982 1840 3988 1841
rect 3838 1839 3844 1840
rect 3838 1835 3839 1839
rect 3843 1835 3844 1839
rect 3982 1836 3983 1840
rect 3987 1836 3988 1840
rect 3982 1835 3988 1836
rect 4222 1840 4228 1841
rect 4222 1836 4223 1840
rect 4227 1836 4228 1840
rect 4222 1835 4228 1836
rect 4494 1840 4500 1841
rect 4494 1836 4495 1840
rect 4499 1836 4500 1840
rect 4494 1835 4500 1836
rect 4798 1840 4804 1841
rect 4798 1836 4799 1840
rect 4803 1836 4804 1840
rect 4798 1835 4804 1836
rect 5118 1840 5124 1841
rect 5118 1836 5119 1840
rect 5123 1836 5124 1840
rect 5118 1835 5124 1836
rect 5438 1840 5444 1841
rect 5438 1836 5439 1840
rect 5443 1836 5444 1840
rect 5438 1835 5444 1836
rect 5662 1839 5668 1840
rect 5662 1835 5663 1839
rect 5667 1835 5668 1839
rect 3838 1834 3844 1835
rect 3840 1811 3842 1834
rect 3984 1811 3986 1835
rect 4224 1811 4226 1835
rect 4496 1811 4498 1835
rect 4800 1811 4802 1835
rect 5120 1811 5122 1835
rect 5440 1811 5442 1835
rect 5662 1834 5668 1835
rect 5664 1811 5666 1834
rect 3839 1810 3843 1811
rect 3839 1805 3843 1806
rect 3983 1810 3987 1811
rect 3983 1805 3987 1806
rect 4223 1810 4227 1811
rect 4223 1805 4227 1806
rect 4367 1810 4371 1811
rect 4367 1805 4371 1806
rect 4495 1810 4499 1811
rect 4495 1805 4499 1806
rect 4575 1810 4579 1811
rect 4575 1805 4579 1806
rect 4783 1810 4787 1811
rect 4783 1805 4787 1806
rect 4799 1810 4803 1811
rect 4799 1805 4803 1806
rect 4983 1810 4987 1811
rect 4983 1805 4987 1806
rect 5119 1810 5123 1811
rect 5119 1805 5123 1806
rect 5175 1810 5179 1811
rect 5175 1805 5179 1806
rect 5367 1810 5371 1811
rect 5367 1805 5371 1806
rect 5439 1810 5443 1811
rect 5439 1805 5443 1806
rect 5543 1810 5547 1811
rect 5543 1805 5547 1806
rect 5663 1810 5667 1811
rect 5663 1805 5667 1806
rect 3798 1784 3804 1785
rect 1974 1780 1975 1784
rect 1979 1780 1980 1784
rect 1974 1779 1980 1780
rect 2210 1783 2216 1784
rect 2210 1779 2211 1783
rect 2215 1779 2216 1783
rect 2210 1778 2216 1779
rect 2354 1783 2360 1784
rect 2354 1779 2355 1783
rect 2359 1779 2360 1783
rect 2354 1778 2360 1779
rect 2498 1783 2504 1784
rect 2498 1779 2499 1783
rect 2503 1779 2504 1783
rect 2498 1778 2504 1779
rect 2642 1783 2648 1784
rect 2642 1779 2643 1783
rect 2647 1779 2648 1783
rect 2642 1778 2648 1779
rect 2786 1783 2792 1784
rect 2786 1779 2787 1783
rect 2791 1779 2792 1783
rect 2786 1778 2792 1779
rect 2930 1783 2936 1784
rect 2930 1779 2931 1783
rect 2935 1779 2936 1783
rect 2930 1778 2936 1779
rect 3082 1783 3088 1784
rect 3082 1779 3083 1783
rect 3087 1779 3088 1783
rect 3798 1780 3799 1784
rect 3803 1780 3804 1784
rect 3840 1782 3842 1805
rect 3798 1779 3804 1780
rect 3838 1781 3844 1782
rect 4368 1781 4370 1805
rect 4576 1781 4578 1805
rect 4784 1781 4786 1805
rect 4984 1781 4986 1805
rect 5176 1781 5178 1805
rect 5368 1781 5370 1805
rect 5544 1781 5546 1805
rect 5664 1782 5666 1805
rect 5662 1781 5668 1782
rect 3082 1778 3088 1779
rect 3838 1777 3839 1781
rect 3843 1777 3844 1781
rect 3838 1776 3844 1777
rect 4366 1780 4372 1781
rect 4366 1776 4367 1780
rect 4371 1776 4372 1780
rect 4366 1775 4372 1776
rect 4574 1780 4580 1781
rect 4574 1776 4575 1780
rect 4579 1776 4580 1780
rect 4574 1775 4580 1776
rect 4782 1780 4788 1781
rect 4782 1776 4783 1780
rect 4787 1776 4788 1780
rect 4782 1775 4788 1776
rect 4982 1780 4988 1781
rect 4982 1776 4983 1780
rect 4987 1776 4988 1780
rect 4982 1775 4988 1776
rect 5174 1780 5180 1781
rect 5174 1776 5175 1780
rect 5179 1776 5180 1780
rect 5174 1775 5180 1776
rect 5366 1780 5372 1781
rect 5366 1776 5367 1780
rect 5371 1776 5372 1780
rect 5366 1775 5372 1776
rect 5542 1780 5548 1781
rect 5542 1776 5543 1780
rect 5547 1776 5548 1780
rect 5662 1777 5663 1781
rect 5667 1777 5668 1781
rect 5662 1776 5668 1777
rect 5542 1775 5548 1776
rect 1934 1773 1940 1774
rect 110 1769 111 1773
rect 115 1769 116 1773
rect 110 1768 116 1769
rect 534 1772 540 1773
rect 534 1768 535 1772
rect 539 1768 540 1772
rect 534 1767 540 1768
rect 694 1772 700 1773
rect 694 1768 695 1772
rect 699 1768 700 1772
rect 694 1767 700 1768
rect 854 1772 860 1773
rect 854 1768 855 1772
rect 859 1768 860 1772
rect 854 1767 860 1768
rect 1014 1772 1020 1773
rect 1014 1768 1015 1772
rect 1019 1768 1020 1772
rect 1014 1767 1020 1768
rect 1182 1772 1188 1773
rect 1182 1768 1183 1772
rect 1187 1768 1188 1772
rect 1182 1767 1188 1768
rect 1350 1772 1356 1773
rect 1350 1768 1351 1772
rect 1355 1768 1356 1772
rect 1350 1767 1356 1768
rect 1518 1772 1524 1773
rect 1518 1768 1519 1772
rect 1523 1768 1524 1772
rect 1934 1769 1935 1773
rect 1939 1769 1940 1773
rect 1934 1768 1940 1769
rect 2238 1768 2244 1769
rect 1518 1767 1524 1768
rect 1974 1767 1980 1768
rect 1974 1763 1975 1767
rect 1979 1763 1980 1767
rect 2238 1764 2239 1768
rect 2243 1764 2244 1768
rect 2238 1763 2244 1764
rect 2382 1768 2388 1769
rect 2382 1764 2383 1768
rect 2387 1764 2388 1768
rect 2382 1763 2388 1764
rect 2526 1768 2532 1769
rect 2526 1764 2527 1768
rect 2531 1764 2532 1768
rect 2526 1763 2532 1764
rect 2670 1768 2676 1769
rect 2670 1764 2671 1768
rect 2675 1764 2676 1768
rect 2670 1763 2676 1764
rect 2814 1768 2820 1769
rect 2814 1764 2815 1768
rect 2819 1764 2820 1768
rect 2814 1763 2820 1764
rect 2958 1768 2964 1769
rect 2958 1764 2959 1768
rect 2963 1764 2964 1768
rect 2958 1763 2964 1764
rect 3110 1768 3116 1769
rect 3110 1764 3111 1768
rect 3115 1764 3116 1768
rect 3110 1763 3116 1764
rect 3798 1767 3804 1768
rect 3798 1763 3799 1767
rect 3803 1763 3804 1767
rect 4338 1765 4344 1766
rect 1974 1762 1980 1763
rect 506 1757 512 1758
rect 110 1756 116 1757
rect 110 1752 111 1756
rect 115 1752 116 1756
rect 506 1753 507 1757
rect 511 1753 512 1757
rect 506 1752 512 1753
rect 666 1757 672 1758
rect 666 1753 667 1757
rect 671 1753 672 1757
rect 666 1752 672 1753
rect 826 1757 832 1758
rect 826 1753 827 1757
rect 831 1753 832 1757
rect 826 1752 832 1753
rect 986 1757 992 1758
rect 986 1753 987 1757
rect 991 1753 992 1757
rect 986 1752 992 1753
rect 1154 1757 1160 1758
rect 1154 1753 1155 1757
rect 1159 1753 1160 1757
rect 1154 1752 1160 1753
rect 1322 1757 1328 1758
rect 1322 1753 1323 1757
rect 1327 1753 1328 1757
rect 1322 1752 1328 1753
rect 1490 1757 1496 1758
rect 1490 1753 1491 1757
rect 1495 1753 1496 1757
rect 1490 1752 1496 1753
rect 1934 1756 1940 1757
rect 1934 1752 1935 1756
rect 1939 1752 1940 1756
rect 110 1751 116 1752
rect 112 1675 114 1751
rect 508 1675 510 1752
rect 668 1675 670 1752
rect 828 1675 830 1752
rect 988 1675 990 1752
rect 1156 1675 1158 1752
rect 1324 1675 1326 1752
rect 1492 1675 1494 1752
rect 1934 1751 1940 1752
rect 1936 1675 1938 1751
rect 1976 1739 1978 1762
rect 2240 1739 2242 1763
rect 2384 1739 2386 1763
rect 2528 1739 2530 1763
rect 2672 1739 2674 1763
rect 2816 1739 2818 1763
rect 2960 1739 2962 1763
rect 3112 1739 3114 1763
rect 3798 1762 3804 1763
rect 3838 1764 3844 1765
rect 3800 1739 3802 1762
rect 3838 1760 3839 1764
rect 3843 1760 3844 1764
rect 4338 1761 4339 1765
rect 4343 1761 4344 1765
rect 4338 1760 4344 1761
rect 4546 1765 4552 1766
rect 4546 1761 4547 1765
rect 4551 1761 4552 1765
rect 4546 1760 4552 1761
rect 4754 1765 4760 1766
rect 4754 1761 4755 1765
rect 4759 1761 4760 1765
rect 4754 1760 4760 1761
rect 4954 1765 4960 1766
rect 4954 1761 4955 1765
rect 4959 1761 4960 1765
rect 4954 1760 4960 1761
rect 5146 1765 5152 1766
rect 5146 1761 5147 1765
rect 5151 1761 5152 1765
rect 5146 1760 5152 1761
rect 5338 1765 5344 1766
rect 5338 1761 5339 1765
rect 5343 1761 5344 1765
rect 5338 1760 5344 1761
rect 5514 1765 5520 1766
rect 5514 1761 5515 1765
rect 5519 1761 5520 1765
rect 5514 1760 5520 1761
rect 5662 1764 5668 1765
rect 5662 1760 5663 1764
rect 5667 1760 5668 1764
rect 3838 1759 3844 1760
rect 1975 1738 1979 1739
rect 1975 1733 1979 1734
rect 2023 1738 2027 1739
rect 2023 1733 2027 1734
rect 2215 1738 2219 1739
rect 2215 1733 2219 1734
rect 2239 1738 2243 1739
rect 2239 1733 2243 1734
rect 2383 1738 2387 1739
rect 2383 1733 2387 1734
rect 2407 1738 2411 1739
rect 2407 1733 2411 1734
rect 2527 1738 2531 1739
rect 2527 1733 2531 1734
rect 2599 1738 2603 1739
rect 2599 1733 2603 1734
rect 2671 1738 2675 1739
rect 2671 1733 2675 1734
rect 2791 1738 2795 1739
rect 2791 1733 2795 1734
rect 2815 1738 2819 1739
rect 2815 1733 2819 1734
rect 2959 1738 2963 1739
rect 2959 1733 2963 1734
rect 2975 1738 2979 1739
rect 2975 1733 2979 1734
rect 3111 1738 3115 1739
rect 3111 1733 3115 1734
rect 3151 1738 3155 1739
rect 3151 1733 3155 1734
rect 3335 1738 3339 1739
rect 3335 1733 3339 1734
rect 3519 1738 3523 1739
rect 3519 1733 3523 1734
rect 3799 1738 3803 1739
rect 3799 1733 3803 1734
rect 1976 1710 1978 1733
rect 1974 1709 1980 1710
rect 2024 1709 2026 1733
rect 2216 1709 2218 1733
rect 2408 1709 2410 1733
rect 2600 1709 2602 1733
rect 2792 1709 2794 1733
rect 2976 1709 2978 1733
rect 3152 1709 3154 1733
rect 3336 1709 3338 1733
rect 3520 1709 3522 1733
rect 3800 1710 3802 1733
rect 3798 1709 3804 1710
rect 1974 1705 1975 1709
rect 1979 1705 1980 1709
rect 1974 1704 1980 1705
rect 2022 1708 2028 1709
rect 2022 1704 2023 1708
rect 2027 1704 2028 1708
rect 2022 1703 2028 1704
rect 2214 1708 2220 1709
rect 2214 1704 2215 1708
rect 2219 1704 2220 1708
rect 2214 1703 2220 1704
rect 2406 1708 2412 1709
rect 2406 1704 2407 1708
rect 2411 1704 2412 1708
rect 2406 1703 2412 1704
rect 2598 1708 2604 1709
rect 2598 1704 2599 1708
rect 2603 1704 2604 1708
rect 2598 1703 2604 1704
rect 2790 1708 2796 1709
rect 2790 1704 2791 1708
rect 2795 1704 2796 1708
rect 2790 1703 2796 1704
rect 2974 1708 2980 1709
rect 2974 1704 2975 1708
rect 2979 1704 2980 1708
rect 2974 1703 2980 1704
rect 3150 1708 3156 1709
rect 3150 1704 3151 1708
rect 3155 1704 3156 1708
rect 3150 1703 3156 1704
rect 3334 1708 3340 1709
rect 3334 1704 3335 1708
rect 3339 1704 3340 1708
rect 3334 1703 3340 1704
rect 3518 1708 3524 1709
rect 3518 1704 3519 1708
rect 3523 1704 3524 1708
rect 3798 1705 3799 1709
rect 3803 1705 3804 1709
rect 3798 1704 3804 1705
rect 3518 1703 3524 1704
rect 1994 1693 2000 1694
rect 1974 1692 1980 1693
rect 1974 1688 1975 1692
rect 1979 1688 1980 1692
rect 1994 1689 1995 1693
rect 1999 1689 2000 1693
rect 1994 1688 2000 1689
rect 2186 1693 2192 1694
rect 2186 1689 2187 1693
rect 2191 1689 2192 1693
rect 2186 1688 2192 1689
rect 2378 1693 2384 1694
rect 2378 1689 2379 1693
rect 2383 1689 2384 1693
rect 2378 1688 2384 1689
rect 2570 1693 2576 1694
rect 2570 1689 2571 1693
rect 2575 1689 2576 1693
rect 2570 1688 2576 1689
rect 2762 1693 2768 1694
rect 2762 1689 2763 1693
rect 2767 1689 2768 1693
rect 2762 1688 2768 1689
rect 2946 1693 2952 1694
rect 2946 1689 2947 1693
rect 2951 1689 2952 1693
rect 2946 1688 2952 1689
rect 3122 1693 3128 1694
rect 3122 1689 3123 1693
rect 3127 1689 3128 1693
rect 3122 1688 3128 1689
rect 3306 1693 3312 1694
rect 3306 1689 3307 1693
rect 3311 1689 3312 1693
rect 3306 1688 3312 1689
rect 3490 1693 3496 1694
rect 3490 1689 3491 1693
rect 3495 1689 3496 1693
rect 3490 1688 3496 1689
rect 3798 1692 3804 1693
rect 3798 1688 3799 1692
rect 3803 1688 3804 1692
rect 1974 1687 1980 1688
rect 111 1674 115 1675
rect 111 1669 115 1670
rect 427 1674 431 1675
rect 427 1669 431 1670
rect 507 1674 511 1675
rect 507 1669 511 1670
rect 611 1674 615 1675
rect 611 1669 615 1670
rect 667 1674 671 1675
rect 667 1669 671 1670
rect 803 1674 807 1675
rect 803 1669 807 1670
rect 827 1674 831 1675
rect 827 1669 831 1670
rect 987 1674 991 1675
rect 987 1669 991 1670
rect 995 1674 999 1675
rect 995 1669 999 1670
rect 1155 1674 1159 1675
rect 1155 1669 1159 1670
rect 1187 1674 1191 1675
rect 1187 1669 1191 1670
rect 1323 1674 1327 1675
rect 1323 1669 1327 1670
rect 1379 1674 1383 1675
rect 1379 1669 1383 1670
rect 1491 1674 1495 1675
rect 1491 1669 1495 1670
rect 1935 1674 1939 1675
rect 1935 1669 1939 1670
rect 112 1609 114 1669
rect 110 1608 116 1609
rect 428 1608 430 1669
rect 612 1608 614 1669
rect 804 1608 806 1669
rect 996 1608 998 1669
rect 1188 1608 1190 1669
rect 1380 1608 1382 1669
rect 1936 1609 1938 1669
rect 1976 1627 1978 1687
rect 1996 1627 1998 1688
rect 2188 1627 2190 1688
rect 2380 1627 2382 1688
rect 2572 1627 2574 1688
rect 2764 1627 2766 1688
rect 2948 1627 2950 1688
rect 3124 1627 3126 1688
rect 3308 1627 3310 1688
rect 3492 1627 3494 1688
rect 3798 1687 3804 1688
rect 3800 1627 3802 1687
rect 3840 1683 3842 1759
rect 4340 1683 4342 1760
rect 4548 1683 4550 1760
rect 4756 1683 4758 1760
rect 4956 1683 4958 1760
rect 5148 1683 5150 1760
rect 5340 1683 5342 1760
rect 5516 1683 5518 1760
rect 5662 1759 5668 1760
rect 5664 1683 5666 1759
rect 3839 1682 3843 1683
rect 3839 1677 3843 1678
rect 4339 1682 4343 1683
rect 4339 1677 4343 1678
rect 4547 1682 4551 1683
rect 4547 1677 4551 1678
rect 4603 1682 4607 1683
rect 4603 1677 4607 1678
rect 4755 1682 4759 1683
rect 4755 1677 4759 1678
rect 4787 1682 4791 1683
rect 4787 1677 4791 1678
rect 4955 1682 4959 1683
rect 4955 1677 4959 1678
rect 4971 1682 4975 1683
rect 4971 1677 4975 1678
rect 5147 1682 5151 1683
rect 5147 1677 5151 1678
rect 5155 1682 5159 1683
rect 5155 1677 5159 1678
rect 5339 1682 5343 1683
rect 5339 1677 5343 1678
rect 5515 1682 5519 1683
rect 5515 1677 5519 1678
rect 5663 1682 5667 1683
rect 5663 1677 5667 1678
rect 1975 1626 1979 1627
rect 1975 1621 1979 1622
rect 1995 1626 1999 1627
rect 1995 1621 1999 1622
rect 2163 1626 2167 1627
rect 2163 1621 2167 1622
rect 2187 1626 2191 1627
rect 2187 1621 2191 1622
rect 2371 1626 2375 1627
rect 2371 1621 2375 1622
rect 2379 1626 2383 1627
rect 2379 1621 2383 1622
rect 2571 1626 2575 1627
rect 2571 1621 2575 1622
rect 2587 1626 2591 1627
rect 2587 1621 2591 1622
rect 2763 1626 2767 1627
rect 2763 1621 2767 1622
rect 2803 1626 2807 1627
rect 2803 1621 2807 1622
rect 2947 1626 2951 1627
rect 2947 1621 2951 1622
rect 3019 1626 3023 1627
rect 3019 1621 3023 1622
rect 3123 1626 3127 1627
rect 3123 1621 3127 1622
rect 3235 1626 3239 1627
rect 3235 1621 3239 1622
rect 3307 1626 3311 1627
rect 3307 1621 3311 1622
rect 3451 1626 3455 1627
rect 3451 1621 3455 1622
rect 3491 1626 3495 1627
rect 3491 1621 3495 1622
rect 3651 1626 3655 1627
rect 3651 1621 3655 1622
rect 3799 1626 3803 1627
rect 3799 1621 3803 1622
rect 1934 1608 1940 1609
rect 110 1604 111 1608
rect 115 1604 116 1608
rect 110 1603 116 1604
rect 426 1607 432 1608
rect 426 1603 427 1607
rect 431 1603 432 1607
rect 426 1602 432 1603
rect 610 1607 616 1608
rect 610 1603 611 1607
rect 615 1603 616 1607
rect 610 1602 616 1603
rect 802 1607 808 1608
rect 802 1603 803 1607
rect 807 1603 808 1607
rect 802 1602 808 1603
rect 994 1607 1000 1608
rect 994 1603 995 1607
rect 999 1603 1000 1607
rect 994 1602 1000 1603
rect 1186 1607 1192 1608
rect 1186 1603 1187 1607
rect 1191 1603 1192 1607
rect 1186 1602 1192 1603
rect 1378 1607 1384 1608
rect 1378 1603 1379 1607
rect 1383 1603 1384 1607
rect 1934 1604 1935 1608
rect 1939 1604 1940 1608
rect 1934 1603 1940 1604
rect 1378 1602 1384 1603
rect 454 1592 460 1593
rect 110 1591 116 1592
rect 110 1587 111 1591
rect 115 1587 116 1591
rect 454 1588 455 1592
rect 459 1588 460 1592
rect 454 1587 460 1588
rect 638 1592 644 1593
rect 638 1588 639 1592
rect 643 1588 644 1592
rect 638 1587 644 1588
rect 830 1592 836 1593
rect 830 1588 831 1592
rect 835 1588 836 1592
rect 830 1587 836 1588
rect 1022 1592 1028 1593
rect 1022 1588 1023 1592
rect 1027 1588 1028 1592
rect 1022 1587 1028 1588
rect 1214 1592 1220 1593
rect 1214 1588 1215 1592
rect 1219 1588 1220 1592
rect 1214 1587 1220 1588
rect 1406 1592 1412 1593
rect 1406 1588 1407 1592
rect 1411 1588 1412 1592
rect 1406 1587 1412 1588
rect 1934 1591 1940 1592
rect 1934 1587 1935 1591
rect 1939 1587 1940 1591
rect 110 1586 116 1587
rect 112 1555 114 1586
rect 456 1555 458 1587
rect 640 1555 642 1587
rect 832 1555 834 1587
rect 1024 1555 1026 1587
rect 1216 1555 1218 1587
rect 1408 1555 1410 1587
rect 1934 1586 1940 1587
rect 1936 1555 1938 1586
rect 1976 1561 1978 1621
rect 1974 1560 1980 1561
rect 1996 1560 1998 1621
rect 2164 1560 2166 1621
rect 2372 1560 2374 1621
rect 2588 1560 2590 1621
rect 2804 1560 2806 1621
rect 3020 1560 3022 1621
rect 3236 1560 3238 1621
rect 3452 1560 3454 1621
rect 3652 1560 3654 1621
rect 3800 1561 3802 1621
rect 3840 1617 3842 1677
rect 3838 1616 3844 1617
rect 4604 1616 4606 1677
rect 4788 1616 4790 1677
rect 4972 1616 4974 1677
rect 5156 1616 5158 1677
rect 5340 1616 5342 1677
rect 5516 1616 5518 1677
rect 5664 1617 5666 1677
rect 5662 1616 5668 1617
rect 3838 1612 3839 1616
rect 3843 1612 3844 1616
rect 3838 1611 3844 1612
rect 4602 1615 4608 1616
rect 4602 1611 4603 1615
rect 4607 1611 4608 1615
rect 4602 1610 4608 1611
rect 4786 1615 4792 1616
rect 4786 1611 4787 1615
rect 4791 1611 4792 1615
rect 4786 1610 4792 1611
rect 4970 1615 4976 1616
rect 4970 1611 4971 1615
rect 4975 1611 4976 1615
rect 4970 1610 4976 1611
rect 5154 1615 5160 1616
rect 5154 1611 5155 1615
rect 5159 1611 5160 1615
rect 5154 1610 5160 1611
rect 5338 1615 5344 1616
rect 5338 1611 5339 1615
rect 5343 1611 5344 1615
rect 5338 1610 5344 1611
rect 5514 1615 5520 1616
rect 5514 1611 5515 1615
rect 5519 1611 5520 1615
rect 5662 1612 5663 1616
rect 5667 1612 5668 1616
rect 5662 1611 5668 1612
rect 5514 1610 5520 1611
rect 4630 1600 4636 1601
rect 3838 1599 3844 1600
rect 3838 1595 3839 1599
rect 3843 1595 3844 1599
rect 4630 1596 4631 1600
rect 4635 1596 4636 1600
rect 4630 1595 4636 1596
rect 4814 1600 4820 1601
rect 4814 1596 4815 1600
rect 4819 1596 4820 1600
rect 4814 1595 4820 1596
rect 4998 1600 5004 1601
rect 4998 1596 4999 1600
rect 5003 1596 5004 1600
rect 4998 1595 5004 1596
rect 5182 1600 5188 1601
rect 5182 1596 5183 1600
rect 5187 1596 5188 1600
rect 5182 1595 5188 1596
rect 5366 1600 5372 1601
rect 5366 1596 5367 1600
rect 5371 1596 5372 1600
rect 5366 1595 5372 1596
rect 5542 1600 5548 1601
rect 5542 1596 5543 1600
rect 5547 1596 5548 1600
rect 5542 1595 5548 1596
rect 5662 1599 5668 1600
rect 5662 1595 5663 1599
rect 5667 1595 5668 1599
rect 3838 1594 3844 1595
rect 3798 1560 3804 1561
rect 1974 1556 1975 1560
rect 1979 1556 1980 1560
rect 1974 1555 1980 1556
rect 1994 1559 2000 1560
rect 1994 1555 1995 1559
rect 1999 1555 2000 1559
rect 111 1554 115 1555
rect 111 1549 115 1550
rect 359 1554 363 1555
rect 359 1549 363 1550
rect 455 1554 459 1555
rect 455 1549 459 1550
rect 631 1554 635 1555
rect 631 1549 635 1550
rect 639 1554 643 1555
rect 639 1549 643 1550
rect 831 1554 835 1555
rect 831 1549 835 1550
rect 887 1554 891 1555
rect 887 1549 891 1550
rect 1023 1554 1027 1555
rect 1023 1549 1027 1550
rect 1135 1554 1139 1555
rect 1135 1549 1139 1550
rect 1215 1554 1219 1555
rect 1215 1549 1219 1550
rect 1367 1554 1371 1555
rect 1367 1549 1371 1550
rect 1407 1554 1411 1555
rect 1407 1549 1411 1550
rect 1599 1554 1603 1555
rect 1599 1549 1603 1550
rect 1815 1554 1819 1555
rect 1815 1549 1819 1550
rect 1935 1554 1939 1555
rect 1994 1554 2000 1555
rect 2162 1559 2168 1560
rect 2162 1555 2163 1559
rect 2167 1555 2168 1559
rect 2162 1554 2168 1555
rect 2370 1559 2376 1560
rect 2370 1555 2371 1559
rect 2375 1555 2376 1559
rect 2370 1554 2376 1555
rect 2586 1559 2592 1560
rect 2586 1555 2587 1559
rect 2591 1555 2592 1559
rect 2586 1554 2592 1555
rect 2802 1559 2808 1560
rect 2802 1555 2803 1559
rect 2807 1555 2808 1559
rect 2802 1554 2808 1555
rect 3018 1559 3024 1560
rect 3018 1555 3019 1559
rect 3023 1555 3024 1559
rect 3018 1554 3024 1555
rect 3234 1559 3240 1560
rect 3234 1555 3235 1559
rect 3239 1555 3240 1559
rect 3234 1554 3240 1555
rect 3450 1559 3456 1560
rect 3450 1555 3451 1559
rect 3455 1555 3456 1559
rect 3450 1554 3456 1555
rect 3650 1559 3656 1560
rect 3650 1555 3651 1559
rect 3655 1555 3656 1559
rect 3798 1556 3799 1560
rect 3803 1556 3804 1560
rect 3798 1555 3804 1556
rect 3840 1555 3842 1594
rect 4632 1555 4634 1595
rect 4816 1555 4818 1595
rect 5000 1555 5002 1595
rect 5184 1555 5186 1595
rect 5368 1555 5370 1595
rect 5544 1555 5546 1595
rect 5662 1594 5668 1595
rect 5664 1555 5666 1594
rect 3650 1554 3656 1555
rect 3839 1554 3843 1555
rect 1935 1549 1939 1550
rect 3839 1549 3843 1550
rect 3887 1554 3891 1555
rect 3887 1549 3891 1550
rect 4031 1554 4035 1555
rect 4031 1549 4035 1550
rect 4199 1554 4203 1555
rect 4199 1549 4203 1550
rect 4367 1554 4371 1555
rect 4367 1549 4371 1550
rect 4527 1554 4531 1555
rect 4527 1549 4531 1550
rect 4631 1554 4635 1555
rect 4631 1549 4635 1550
rect 4695 1554 4699 1555
rect 4695 1549 4699 1550
rect 4815 1554 4819 1555
rect 4815 1549 4819 1550
rect 4863 1554 4867 1555
rect 4863 1549 4867 1550
rect 4999 1554 5003 1555
rect 4999 1549 5003 1550
rect 5031 1554 5035 1555
rect 5031 1549 5035 1550
rect 5183 1554 5187 1555
rect 5183 1549 5187 1550
rect 5207 1554 5211 1555
rect 5207 1549 5211 1550
rect 5367 1554 5371 1555
rect 5367 1549 5371 1550
rect 5383 1554 5387 1555
rect 5383 1549 5387 1550
rect 5543 1554 5547 1555
rect 5543 1549 5547 1550
rect 5663 1554 5667 1555
rect 5663 1549 5667 1550
rect 112 1526 114 1549
rect 110 1525 116 1526
rect 360 1525 362 1549
rect 632 1525 634 1549
rect 888 1525 890 1549
rect 1136 1525 1138 1549
rect 1368 1525 1370 1549
rect 1600 1525 1602 1549
rect 1816 1525 1818 1549
rect 1936 1526 1938 1549
rect 2022 1544 2028 1545
rect 1974 1543 1980 1544
rect 1974 1539 1975 1543
rect 1979 1539 1980 1543
rect 2022 1540 2023 1544
rect 2027 1540 2028 1544
rect 2022 1539 2028 1540
rect 2190 1544 2196 1545
rect 2190 1540 2191 1544
rect 2195 1540 2196 1544
rect 2190 1539 2196 1540
rect 2398 1544 2404 1545
rect 2398 1540 2399 1544
rect 2403 1540 2404 1544
rect 2398 1539 2404 1540
rect 2614 1544 2620 1545
rect 2614 1540 2615 1544
rect 2619 1540 2620 1544
rect 2614 1539 2620 1540
rect 2830 1544 2836 1545
rect 2830 1540 2831 1544
rect 2835 1540 2836 1544
rect 2830 1539 2836 1540
rect 3046 1544 3052 1545
rect 3046 1540 3047 1544
rect 3051 1540 3052 1544
rect 3046 1539 3052 1540
rect 3262 1544 3268 1545
rect 3262 1540 3263 1544
rect 3267 1540 3268 1544
rect 3262 1539 3268 1540
rect 3478 1544 3484 1545
rect 3478 1540 3479 1544
rect 3483 1540 3484 1544
rect 3478 1539 3484 1540
rect 3678 1544 3684 1545
rect 3678 1540 3679 1544
rect 3683 1540 3684 1544
rect 3678 1539 3684 1540
rect 3798 1543 3804 1544
rect 3798 1539 3799 1543
rect 3803 1539 3804 1543
rect 1974 1538 1980 1539
rect 1934 1525 1940 1526
rect 110 1521 111 1525
rect 115 1521 116 1525
rect 110 1520 116 1521
rect 358 1524 364 1525
rect 358 1520 359 1524
rect 363 1520 364 1524
rect 358 1519 364 1520
rect 630 1524 636 1525
rect 630 1520 631 1524
rect 635 1520 636 1524
rect 630 1519 636 1520
rect 886 1524 892 1525
rect 886 1520 887 1524
rect 891 1520 892 1524
rect 886 1519 892 1520
rect 1134 1524 1140 1525
rect 1134 1520 1135 1524
rect 1139 1520 1140 1524
rect 1134 1519 1140 1520
rect 1366 1524 1372 1525
rect 1366 1520 1367 1524
rect 1371 1520 1372 1524
rect 1366 1519 1372 1520
rect 1598 1524 1604 1525
rect 1598 1520 1599 1524
rect 1603 1520 1604 1524
rect 1598 1519 1604 1520
rect 1814 1524 1820 1525
rect 1814 1520 1815 1524
rect 1819 1520 1820 1524
rect 1934 1521 1935 1525
rect 1939 1521 1940 1525
rect 1934 1520 1940 1521
rect 1814 1519 1820 1520
rect 330 1509 336 1510
rect 110 1508 116 1509
rect 110 1504 111 1508
rect 115 1504 116 1508
rect 330 1505 331 1509
rect 335 1505 336 1509
rect 330 1504 336 1505
rect 602 1509 608 1510
rect 602 1505 603 1509
rect 607 1505 608 1509
rect 602 1504 608 1505
rect 858 1509 864 1510
rect 858 1505 859 1509
rect 863 1505 864 1509
rect 858 1504 864 1505
rect 1106 1509 1112 1510
rect 1106 1505 1107 1509
rect 1111 1505 1112 1509
rect 1106 1504 1112 1505
rect 1338 1509 1344 1510
rect 1338 1505 1339 1509
rect 1343 1505 1344 1509
rect 1338 1504 1344 1505
rect 1570 1509 1576 1510
rect 1570 1505 1571 1509
rect 1575 1505 1576 1509
rect 1570 1504 1576 1505
rect 1786 1509 1792 1510
rect 1786 1505 1787 1509
rect 1791 1505 1792 1509
rect 1786 1504 1792 1505
rect 1934 1508 1940 1509
rect 1934 1504 1935 1508
rect 1939 1504 1940 1508
rect 110 1503 116 1504
rect 112 1443 114 1503
rect 332 1443 334 1504
rect 604 1443 606 1504
rect 860 1443 862 1504
rect 1108 1443 1110 1504
rect 1340 1443 1342 1504
rect 1572 1443 1574 1504
rect 1788 1443 1790 1504
rect 1934 1503 1940 1504
rect 1936 1443 1938 1503
rect 111 1442 115 1443
rect 111 1437 115 1438
rect 131 1442 135 1443
rect 131 1437 135 1438
rect 307 1442 311 1443
rect 307 1437 311 1438
rect 331 1442 335 1443
rect 331 1437 335 1438
rect 499 1442 503 1443
rect 499 1437 503 1438
rect 603 1442 607 1443
rect 603 1437 607 1438
rect 683 1442 687 1443
rect 683 1437 687 1438
rect 859 1442 863 1443
rect 859 1437 863 1438
rect 1027 1442 1031 1443
rect 1027 1437 1031 1438
rect 1107 1442 1111 1443
rect 1107 1437 1111 1438
rect 1187 1442 1191 1443
rect 1187 1437 1191 1438
rect 1339 1442 1343 1443
rect 1339 1437 1343 1438
rect 1491 1442 1495 1443
rect 1491 1437 1495 1438
rect 1571 1442 1575 1443
rect 1571 1437 1575 1438
rect 1651 1442 1655 1443
rect 1651 1437 1655 1438
rect 1787 1442 1791 1443
rect 1787 1437 1791 1438
rect 1935 1442 1939 1443
rect 1935 1437 1939 1438
rect 112 1377 114 1437
rect 110 1376 116 1377
rect 132 1376 134 1437
rect 308 1376 310 1437
rect 500 1376 502 1437
rect 684 1376 686 1437
rect 860 1376 862 1437
rect 1028 1376 1030 1437
rect 1188 1376 1190 1437
rect 1340 1376 1342 1437
rect 1492 1376 1494 1437
rect 1652 1376 1654 1437
rect 1788 1376 1790 1437
rect 1936 1377 1938 1437
rect 1934 1376 1940 1377
rect 110 1372 111 1376
rect 115 1372 116 1376
rect 110 1371 116 1372
rect 130 1375 136 1376
rect 130 1371 131 1375
rect 135 1371 136 1375
rect 130 1370 136 1371
rect 306 1375 312 1376
rect 306 1371 307 1375
rect 311 1371 312 1375
rect 306 1370 312 1371
rect 498 1375 504 1376
rect 498 1371 499 1375
rect 503 1371 504 1375
rect 498 1370 504 1371
rect 682 1375 688 1376
rect 682 1371 683 1375
rect 687 1371 688 1375
rect 682 1370 688 1371
rect 858 1375 864 1376
rect 858 1371 859 1375
rect 863 1371 864 1375
rect 858 1370 864 1371
rect 1026 1375 1032 1376
rect 1026 1371 1027 1375
rect 1031 1371 1032 1375
rect 1026 1370 1032 1371
rect 1186 1375 1192 1376
rect 1186 1371 1187 1375
rect 1191 1371 1192 1375
rect 1186 1370 1192 1371
rect 1338 1375 1344 1376
rect 1338 1371 1339 1375
rect 1343 1371 1344 1375
rect 1338 1370 1344 1371
rect 1490 1375 1496 1376
rect 1490 1371 1491 1375
rect 1495 1371 1496 1375
rect 1490 1370 1496 1371
rect 1650 1375 1656 1376
rect 1650 1371 1651 1375
rect 1655 1371 1656 1375
rect 1650 1370 1656 1371
rect 1786 1375 1792 1376
rect 1786 1371 1787 1375
rect 1791 1371 1792 1375
rect 1934 1372 1935 1376
rect 1939 1372 1940 1376
rect 1934 1371 1940 1372
rect 1786 1370 1792 1371
rect 158 1360 164 1361
rect 110 1359 116 1360
rect 110 1355 111 1359
rect 115 1355 116 1359
rect 158 1356 159 1360
rect 163 1356 164 1360
rect 158 1355 164 1356
rect 334 1360 340 1361
rect 334 1356 335 1360
rect 339 1356 340 1360
rect 334 1355 340 1356
rect 526 1360 532 1361
rect 526 1356 527 1360
rect 531 1356 532 1360
rect 526 1355 532 1356
rect 710 1360 716 1361
rect 710 1356 711 1360
rect 715 1356 716 1360
rect 710 1355 716 1356
rect 886 1360 892 1361
rect 886 1356 887 1360
rect 891 1356 892 1360
rect 886 1355 892 1356
rect 1054 1360 1060 1361
rect 1054 1356 1055 1360
rect 1059 1356 1060 1360
rect 1054 1355 1060 1356
rect 1214 1360 1220 1361
rect 1214 1356 1215 1360
rect 1219 1356 1220 1360
rect 1214 1355 1220 1356
rect 1366 1360 1372 1361
rect 1366 1356 1367 1360
rect 1371 1356 1372 1360
rect 1366 1355 1372 1356
rect 1518 1360 1524 1361
rect 1518 1356 1519 1360
rect 1523 1356 1524 1360
rect 1518 1355 1524 1356
rect 1678 1360 1684 1361
rect 1678 1356 1679 1360
rect 1683 1356 1684 1360
rect 1678 1355 1684 1356
rect 1814 1360 1820 1361
rect 1814 1356 1815 1360
rect 1819 1356 1820 1360
rect 1814 1355 1820 1356
rect 1934 1359 1940 1360
rect 1934 1355 1935 1359
rect 1939 1355 1940 1359
rect 110 1354 116 1355
rect 112 1323 114 1354
rect 160 1323 162 1355
rect 336 1323 338 1355
rect 528 1323 530 1355
rect 712 1323 714 1355
rect 888 1323 890 1355
rect 1056 1323 1058 1355
rect 1216 1323 1218 1355
rect 1368 1323 1370 1355
rect 1520 1323 1522 1355
rect 1680 1323 1682 1355
rect 1816 1323 1818 1355
rect 1934 1354 1940 1355
rect 1936 1323 1938 1354
rect 111 1322 115 1323
rect 111 1317 115 1318
rect 159 1322 163 1323
rect 159 1317 163 1318
rect 335 1322 339 1323
rect 335 1317 339 1318
rect 375 1322 379 1323
rect 375 1317 379 1318
rect 527 1322 531 1323
rect 527 1317 531 1318
rect 599 1322 603 1323
rect 599 1317 603 1318
rect 711 1322 715 1323
rect 711 1317 715 1318
rect 807 1322 811 1323
rect 807 1317 811 1318
rect 887 1322 891 1323
rect 887 1317 891 1318
rect 999 1322 1003 1323
rect 999 1317 1003 1318
rect 1055 1322 1059 1323
rect 1055 1317 1059 1318
rect 1175 1322 1179 1323
rect 1175 1317 1179 1318
rect 1215 1322 1219 1323
rect 1215 1317 1219 1318
rect 1343 1322 1347 1323
rect 1343 1317 1347 1318
rect 1367 1322 1371 1323
rect 1367 1317 1371 1318
rect 1511 1322 1515 1323
rect 1511 1317 1515 1318
rect 1519 1322 1523 1323
rect 1519 1317 1523 1318
rect 1671 1322 1675 1323
rect 1671 1317 1675 1318
rect 1679 1322 1683 1323
rect 1679 1317 1683 1318
rect 1815 1322 1819 1323
rect 1815 1317 1819 1318
rect 1935 1322 1939 1323
rect 1935 1317 1939 1318
rect 112 1294 114 1317
rect 110 1293 116 1294
rect 160 1293 162 1317
rect 376 1293 378 1317
rect 600 1293 602 1317
rect 808 1293 810 1317
rect 1000 1293 1002 1317
rect 1176 1293 1178 1317
rect 1344 1293 1346 1317
rect 1512 1293 1514 1317
rect 1672 1293 1674 1317
rect 1816 1293 1818 1317
rect 1936 1294 1938 1317
rect 1976 1311 1978 1538
rect 2024 1311 2026 1539
rect 2192 1311 2194 1539
rect 2400 1311 2402 1539
rect 2616 1311 2618 1539
rect 2832 1311 2834 1539
rect 3048 1311 3050 1539
rect 3264 1311 3266 1539
rect 3480 1311 3482 1539
rect 3680 1311 3682 1539
rect 3798 1538 3804 1539
rect 3800 1311 3802 1538
rect 3840 1526 3842 1549
rect 3838 1525 3844 1526
rect 3888 1525 3890 1549
rect 4032 1525 4034 1549
rect 4200 1525 4202 1549
rect 4368 1525 4370 1549
rect 4528 1525 4530 1549
rect 4696 1525 4698 1549
rect 4864 1525 4866 1549
rect 5032 1525 5034 1549
rect 5208 1525 5210 1549
rect 5384 1525 5386 1549
rect 5544 1525 5546 1549
rect 5664 1526 5666 1549
rect 5662 1525 5668 1526
rect 3838 1521 3839 1525
rect 3843 1521 3844 1525
rect 3838 1520 3844 1521
rect 3886 1524 3892 1525
rect 3886 1520 3887 1524
rect 3891 1520 3892 1524
rect 3886 1519 3892 1520
rect 4030 1524 4036 1525
rect 4030 1520 4031 1524
rect 4035 1520 4036 1524
rect 4030 1519 4036 1520
rect 4198 1524 4204 1525
rect 4198 1520 4199 1524
rect 4203 1520 4204 1524
rect 4198 1519 4204 1520
rect 4366 1524 4372 1525
rect 4366 1520 4367 1524
rect 4371 1520 4372 1524
rect 4366 1519 4372 1520
rect 4526 1524 4532 1525
rect 4526 1520 4527 1524
rect 4531 1520 4532 1524
rect 4526 1519 4532 1520
rect 4694 1524 4700 1525
rect 4694 1520 4695 1524
rect 4699 1520 4700 1524
rect 4694 1519 4700 1520
rect 4862 1524 4868 1525
rect 4862 1520 4863 1524
rect 4867 1520 4868 1524
rect 4862 1519 4868 1520
rect 5030 1524 5036 1525
rect 5030 1520 5031 1524
rect 5035 1520 5036 1524
rect 5030 1519 5036 1520
rect 5206 1524 5212 1525
rect 5206 1520 5207 1524
rect 5211 1520 5212 1524
rect 5206 1519 5212 1520
rect 5382 1524 5388 1525
rect 5382 1520 5383 1524
rect 5387 1520 5388 1524
rect 5382 1519 5388 1520
rect 5542 1524 5548 1525
rect 5542 1520 5543 1524
rect 5547 1520 5548 1524
rect 5662 1521 5663 1525
rect 5667 1521 5668 1525
rect 5662 1520 5668 1521
rect 5542 1519 5548 1520
rect 3858 1509 3864 1510
rect 3838 1508 3844 1509
rect 3838 1504 3839 1508
rect 3843 1504 3844 1508
rect 3858 1505 3859 1509
rect 3863 1505 3864 1509
rect 3858 1504 3864 1505
rect 4002 1509 4008 1510
rect 4002 1505 4003 1509
rect 4007 1505 4008 1509
rect 4002 1504 4008 1505
rect 4170 1509 4176 1510
rect 4170 1505 4171 1509
rect 4175 1505 4176 1509
rect 4170 1504 4176 1505
rect 4338 1509 4344 1510
rect 4338 1505 4339 1509
rect 4343 1505 4344 1509
rect 4338 1504 4344 1505
rect 4498 1509 4504 1510
rect 4498 1505 4499 1509
rect 4503 1505 4504 1509
rect 4498 1504 4504 1505
rect 4666 1509 4672 1510
rect 4666 1505 4667 1509
rect 4671 1505 4672 1509
rect 4666 1504 4672 1505
rect 4834 1509 4840 1510
rect 4834 1505 4835 1509
rect 4839 1505 4840 1509
rect 4834 1504 4840 1505
rect 5002 1509 5008 1510
rect 5002 1505 5003 1509
rect 5007 1505 5008 1509
rect 5002 1504 5008 1505
rect 5178 1509 5184 1510
rect 5178 1505 5179 1509
rect 5183 1505 5184 1509
rect 5178 1504 5184 1505
rect 5354 1509 5360 1510
rect 5354 1505 5355 1509
rect 5359 1505 5360 1509
rect 5354 1504 5360 1505
rect 5514 1509 5520 1510
rect 5514 1505 5515 1509
rect 5519 1505 5520 1509
rect 5514 1504 5520 1505
rect 5662 1508 5668 1509
rect 5662 1504 5663 1508
rect 5667 1504 5668 1508
rect 3838 1503 3844 1504
rect 3840 1439 3842 1503
rect 3860 1439 3862 1504
rect 4004 1439 4006 1504
rect 4172 1439 4174 1504
rect 4340 1439 4342 1504
rect 4500 1439 4502 1504
rect 4668 1439 4670 1504
rect 4836 1439 4838 1504
rect 5004 1439 5006 1504
rect 5180 1439 5182 1504
rect 5356 1439 5358 1504
rect 5516 1439 5518 1504
rect 5662 1503 5668 1504
rect 5664 1439 5666 1503
rect 3839 1438 3843 1439
rect 3839 1433 3843 1434
rect 3859 1438 3863 1439
rect 3859 1433 3863 1434
rect 4003 1438 4007 1439
rect 4003 1433 4007 1434
rect 4171 1438 4175 1439
rect 4171 1433 4175 1434
rect 4179 1438 4183 1439
rect 4179 1433 4183 1434
rect 4339 1438 4343 1439
rect 4339 1433 4343 1434
rect 4355 1438 4359 1439
rect 4355 1433 4359 1434
rect 4499 1438 4503 1439
rect 4499 1433 4503 1434
rect 4531 1438 4535 1439
rect 4531 1433 4535 1434
rect 4667 1438 4671 1439
rect 4667 1433 4671 1434
rect 4707 1438 4711 1439
rect 4707 1433 4711 1434
rect 4835 1438 4839 1439
rect 4835 1433 4839 1434
rect 4875 1438 4879 1439
rect 4875 1433 4879 1434
rect 5003 1438 5007 1439
rect 5003 1433 5007 1434
rect 5043 1438 5047 1439
rect 5043 1433 5047 1434
rect 5179 1438 5183 1439
rect 5179 1433 5183 1434
rect 5203 1438 5207 1439
rect 5203 1433 5207 1434
rect 5355 1438 5359 1439
rect 5355 1433 5359 1434
rect 5371 1438 5375 1439
rect 5371 1433 5375 1434
rect 5515 1438 5519 1439
rect 5515 1433 5519 1434
rect 5663 1438 5667 1439
rect 5663 1433 5667 1434
rect 3840 1373 3842 1433
rect 3838 1372 3844 1373
rect 3860 1372 3862 1433
rect 4004 1372 4006 1433
rect 4180 1372 4182 1433
rect 4356 1372 4358 1433
rect 4532 1372 4534 1433
rect 4708 1372 4710 1433
rect 4876 1372 4878 1433
rect 5044 1372 5046 1433
rect 5204 1372 5206 1433
rect 5372 1372 5374 1433
rect 5516 1372 5518 1433
rect 5664 1373 5666 1433
rect 5662 1372 5668 1373
rect 3838 1368 3839 1372
rect 3843 1368 3844 1372
rect 3838 1367 3844 1368
rect 3858 1371 3864 1372
rect 3858 1367 3859 1371
rect 3863 1367 3864 1371
rect 3858 1366 3864 1367
rect 4002 1371 4008 1372
rect 4002 1367 4003 1371
rect 4007 1367 4008 1371
rect 4002 1366 4008 1367
rect 4178 1371 4184 1372
rect 4178 1367 4179 1371
rect 4183 1367 4184 1371
rect 4178 1366 4184 1367
rect 4354 1371 4360 1372
rect 4354 1367 4355 1371
rect 4359 1367 4360 1371
rect 4354 1366 4360 1367
rect 4530 1371 4536 1372
rect 4530 1367 4531 1371
rect 4535 1367 4536 1371
rect 4530 1366 4536 1367
rect 4706 1371 4712 1372
rect 4706 1367 4707 1371
rect 4711 1367 4712 1371
rect 4706 1366 4712 1367
rect 4874 1371 4880 1372
rect 4874 1367 4875 1371
rect 4879 1367 4880 1371
rect 4874 1366 4880 1367
rect 5042 1371 5048 1372
rect 5042 1367 5043 1371
rect 5047 1367 5048 1371
rect 5042 1366 5048 1367
rect 5202 1371 5208 1372
rect 5202 1367 5203 1371
rect 5207 1367 5208 1371
rect 5202 1366 5208 1367
rect 5370 1371 5376 1372
rect 5370 1367 5371 1371
rect 5375 1367 5376 1371
rect 5370 1366 5376 1367
rect 5514 1371 5520 1372
rect 5514 1367 5515 1371
rect 5519 1367 5520 1371
rect 5662 1368 5663 1372
rect 5667 1368 5668 1372
rect 5662 1367 5668 1368
rect 5514 1366 5520 1367
rect 3886 1356 3892 1357
rect 3838 1355 3844 1356
rect 3838 1351 3839 1355
rect 3843 1351 3844 1355
rect 3886 1352 3887 1356
rect 3891 1352 3892 1356
rect 3886 1351 3892 1352
rect 4030 1356 4036 1357
rect 4030 1352 4031 1356
rect 4035 1352 4036 1356
rect 4030 1351 4036 1352
rect 4206 1356 4212 1357
rect 4206 1352 4207 1356
rect 4211 1352 4212 1356
rect 4206 1351 4212 1352
rect 4382 1356 4388 1357
rect 4382 1352 4383 1356
rect 4387 1352 4388 1356
rect 4382 1351 4388 1352
rect 4558 1356 4564 1357
rect 4558 1352 4559 1356
rect 4563 1352 4564 1356
rect 4558 1351 4564 1352
rect 4734 1356 4740 1357
rect 4734 1352 4735 1356
rect 4739 1352 4740 1356
rect 4734 1351 4740 1352
rect 4902 1356 4908 1357
rect 4902 1352 4903 1356
rect 4907 1352 4908 1356
rect 4902 1351 4908 1352
rect 5070 1356 5076 1357
rect 5070 1352 5071 1356
rect 5075 1352 5076 1356
rect 5070 1351 5076 1352
rect 5230 1356 5236 1357
rect 5230 1352 5231 1356
rect 5235 1352 5236 1356
rect 5230 1351 5236 1352
rect 5398 1356 5404 1357
rect 5398 1352 5399 1356
rect 5403 1352 5404 1356
rect 5398 1351 5404 1352
rect 5542 1356 5548 1357
rect 5542 1352 5543 1356
rect 5547 1352 5548 1356
rect 5542 1351 5548 1352
rect 5662 1355 5668 1356
rect 5662 1351 5663 1355
rect 5667 1351 5668 1355
rect 3838 1350 3844 1351
rect 3840 1327 3842 1350
rect 3888 1327 3890 1351
rect 4032 1327 4034 1351
rect 4208 1327 4210 1351
rect 4384 1327 4386 1351
rect 4560 1327 4562 1351
rect 4736 1327 4738 1351
rect 4904 1327 4906 1351
rect 5072 1327 5074 1351
rect 5232 1327 5234 1351
rect 5400 1327 5402 1351
rect 5544 1327 5546 1351
rect 5662 1350 5668 1351
rect 5664 1327 5666 1350
rect 3839 1326 3843 1327
rect 3839 1321 3843 1322
rect 3887 1326 3891 1327
rect 3887 1321 3891 1322
rect 4031 1326 4035 1327
rect 4031 1321 4035 1322
rect 4175 1326 4179 1327
rect 4175 1321 4179 1322
rect 4207 1326 4211 1327
rect 4207 1321 4211 1322
rect 4383 1326 4387 1327
rect 4383 1321 4387 1322
rect 4471 1326 4475 1327
rect 4471 1321 4475 1322
rect 4559 1326 4563 1327
rect 4559 1321 4563 1322
rect 4735 1326 4739 1327
rect 4735 1321 4739 1322
rect 4751 1326 4755 1327
rect 4751 1321 4755 1322
rect 4903 1326 4907 1327
rect 4903 1321 4907 1322
rect 5023 1326 5027 1327
rect 5023 1321 5027 1322
rect 5071 1326 5075 1327
rect 5071 1321 5075 1322
rect 5231 1326 5235 1327
rect 5231 1321 5235 1322
rect 5287 1326 5291 1327
rect 5287 1321 5291 1322
rect 5399 1326 5403 1327
rect 5399 1321 5403 1322
rect 5543 1326 5547 1327
rect 5543 1321 5547 1322
rect 5663 1326 5667 1327
rect 5663 1321 5667 1322
rect 1975 1310 1979 1311
rect 1975 1305 1979 1306
rect 2023 1310 2027 1311
rect 2023 1305 2027 1306
rect 2191 1310 2195 1311
rect 2191 1305 2195 1306
rect 2399 1310 2403 1311
rect 2399 1305 2403 1306
rect 2615 1310 2619 1311
rect 2615 1305 2619 1306
rect 2831 1310 2835 1311
rect 2831 1305 2835 1306
rect 3047 1310 3051 1311
rect 3047 1305 3051 1306
rect 3263 1310 3267 1311
rect 3263 1305 3267 1306
rect 3271 1310 3275 1311
rect 3271 1305 3275 1306
rect 3407 1310 3411 1311
rect 3407 1305 3411 1306
rect 3479 1310 3483 1311
rect 3479 1305 3483 1306
rect 3543 1310 3547 1311
rect 3543 1305 3547 1306
rect 3679 1310 3683 1311
rect 3679 1305 3683 1306
rect 3799 1310 3803 1311
rect 3799 1305 3803 1306
rect 1934 1293 1940 1294
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 158 1292 164 1293
rect 158 1288 159 1292
rect 163 1288 164 1292
rect 158 1287 164 1288
rect 374 1292 380 1293
rect 374 1288 375 1292
rect 379 1288 380 1292
rect 374 1287 380 1288
rect 598 1292 604 1293
rect 598 1288 599 1292
rect 603 1288 604 1292
rect 598 1287 604 1288
rect 806 1292 812 1293
rect 806 1288 807 1292
rect 811 1288 812 1292
rect 806 1287 812 1288
rect 998 1292 1004 1293
rect 998 1288 999 1292
rect 1003 1288 1004 1292
rect 998 1287 1004 1288
rect 1174 1292 1180 1293
rect 1174 1288 1175 1292
rect 1179 1288 1180 1292
rect 1174 1287 1180 1288
rect 1342 1292 1348 1293
rect 1342 1288 1343 1292
rect 1347 1288 1348 1292
rect 1342 1287 1348 1288
rect 1510 1292 1516 1293
rect 1510 1288 1511 1292
rect 1515 1288 1516 1292
rect 1510 1287 1516 1288
rect 1670 1292 1676 1293
rect 1670 1288 1671 1292
rect 1675 1288 1676 1292
rect 1670 1287 1676 1288
rect 1814 1292 1820 1293
rect 1814 1288 1815 1292
rect 1819 1288 1820 1292
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 1934 1288 1940 1289
rect 1814 1287 1820 1288
rect 1976 1282 1978 1305
rect 1974 1281 1980 1282
rect 3272 1281 3274 1305
rect 3408 1281 3410 1305
rect 3544 1281 3546 1305
rect 3680 1281 3682 1305
rect 3800 1282 3802 1305
rect 3840 1298 3842 1321
rect 3838 1297 3844 1298
rect 3888 1297 3890 1321
rect 4176 1297 4178 1321
rect 4472 1297 4474 1321
rect 4752 1297 4754 1321
rect 5024 1297 5026 1321
rect 5288 1297 5290 1321
rect 5544 1297 5546 1321
rect 5664 1298 5666 1321
rect 5662 1297 5668 1298
rect 3838 1293 3839 1297
rect 3843 1293 3844 1297
rect 3838 1292 3844 1293
rect 3886 1296 3892 1297
rect 3886 1292 3887 1296
rect 3891 1292 3892 1296
rect 3886 1291 3892 1292
rect 4174 1296 4180 1297
rect 4174 1292 4175 1296
rect 4179 1292 4180 1296
rect 4174 1291 4180 1292
rect 4470 1296 4476 1297
rect 4470 1292 4471 1296
rect 4475 1292 4476 1296
rect 4470 1291 4476 1292
rect 4750 1296 4756 1297
rect 4750 1292 4751 1296
rect 4755 1292 4756 1296
rect 4750 1291 4756 1292
rect 5022 1296 5028 1297
rect 5022 1292 5023 1296
rect 5027 1292 5028 1296
rect 5022 1291 5028 1292
rect 5286 1296 5292 1297
rect 5286 1292 5287 1296
rect 5291 1292 5292 1296
rect 5286 1291 5292 1292
rect 5542 1296 5548 1297
rect 5542 1292 5543 1296
rect 5547 1292 5548 1296
rect 5662 1293 5663 1297
rect 5667 1293 5668 1297
rect 5662 1292 5668 1293
rect 5542 1291 5548 1292
rect 3798 1281 3804 1282
rect 3858 1281 3864 1282
rect 130 1277 136 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 130 1273 131 1277
rect 135 1273 136 1277
rect 130 1272 136 1273
rect 346 1277 352 1278
rect 346 1273 347 1277
rect 351 1273 352 1277
rect 346 1272 352 1273
rect 570 1277 576 1278
rect 570 1273 571 1277
rect 575 1273 576 1277
rect 570 1272 576 1273
rect 778 1277 784 1278
rect 778 1273 779 1277
rect 783 1273 784 1277
rect 778 1272 784 1273
rect 970 1277 976 1278
rect 970 1273 971 1277
rect 975 1273 976 1277
rect 970 1272 976 1273
rect 1146 1277 1152 1278
rect 1146 1273 1147 1277
rect 1151 1273 1152 1277
rect 1146 1272 1152 1273
rect 1314 1277 1320 1278
rect 1314 1273 1315 1277
rect 1319 1273 1320 1277
rect 1314 1272 1320 1273
rect 1482 1277 1488 1278
rect 1482 1273 1483 1277
rect 1487 1273 1488 1277
rect 1482 1272 1488 1273
rect 1642 1277 1648 1278
rect 1642 1273 1643 1277
rect 1647 1273 1648 1277
rect 1642 1272 1648 1273
rect 1786 1277 1792 1278
rect 1974 1277 1975 1281
rect 1979 1277 1980 1281
rect 1786 1273 1787 1277
rect 1791 1273 1792 1277
rect 1786 1272 1792 1273
rect 1934 1276 1940 1277
rect 1974 1276 1980 1277
rect 3270 1280 3276 1281
rect 3270 1276 3271 1280
rect 3275 1276 3276 1280
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 3270 1275 3276 1276
rect 3406 1280 3412 1281
rect 3406 1276 3407 1280
rect 3411 1276 3412 1280
rect 3406 1275 3412 1276
rect 3542 1280 3548 1281
rect 3542 1276 3543 1280
rect 3547 1276 3548 1280
rect 3542 1275 3548 1276
rect 3678 1280 3684 1281
rect 3678 1276 3679 1280
rect 3683 1276 3684 1280
rect 3798 1277 3799 1281
rect 3803 1277 3804 1281
rect 3798 1276 3804 1277
rect 3838 1280 3844 1281
rect 3838 1276 3839 1280
rect 3843 1276 3844 1280
rect 3858 1277 3859 1281
rect 3863 1277 3864 1281
rect 3858 1276 3864 1277
rect 4146 1281 4152 1282
rect 4146 1277 4147 1281
rect 4151 1277 4152 1281
rect 4146 1276 4152 1277
rect 4442 1281 4448 1282
rect 4442 1277 4443 1281
rect 4447 1277 4448 1281
rect 4442 1276 4448 1277
rect 4722 1281 4728 1282
rect 4722 1277 4723 1281
rect 4727 1277 4728 1281
rect 4722 1276 4728 1277
rect 4994 1281 5000 1282
rect 4994 1277 4995 1281
rect 4999 1277 5000 1281
rect 4994 1276 5000 1277
rect 5258 1281 5264 1282
rect 5258 1277 5259 1281
rect 5263 1277 5264 1281
rect 5258 1276 5264 1277
rect 5514 1281 5520 1282
rect 5514 1277 5515 1281
rect 5519 1277 5520 1281
rect 5514 1276 5520 1277
rect 5662 1280 5668 1281
rect 5662 1276 5663 1280
rect 5667 1276 5668 1280
rect 3678 1275 3684 1276
rect 3838 1275 3844 1276
rect 110 1271 116 1272
rect 112 1211 114 1271
rect 132 1211 134 1272
rect 348 1211 350 1272
rect 572 1211 574 1272
rect 780 1211 782 1272
rect 972 1211 974 1272
rect 1148 1211 1150 1272
rect 1316 1211 1318 1272
rect 1484 1211 1486 1272
rect 1644 1211 1646 1272
rect 1788 1211 1790 1272
rect 1934 1271 1940 1272
rect 1936 1211 1938 1271
rect 3242 1265 3248 1266
rect 1974 1264 1980 1265
rect 1974 1260 1975 1264
rect 1979 1260 1980 1264
rect 3242 1261 3243 1265
rect 3247 1261 3248 1265
rect 3242 1260 3248 1261
rect 3378 1265 3384 1266
rect 3378 1261 3379 1265
rect 3383 1261 3384 1265
rect 3378 1260 3384 1261
rect 3514 1265 3520 1266
rect 3514 1261 3515 1265
rect 3519 1261 3520 1265
rect 3514 1260 3520 1261
rect 3650 1265 3656 1266
rect 3650 1261 3651 1265
rect 3655 1261 3656 1265
rect 3650 1260 3656 1261
rect 3798 1264 3804 1265
rect 3798 1260 3799 1264
rect 3803 1260 3804 1264
rect 1974 1259 1980 1260
rect 111 1210 115 1211
rect 111 1205 115 1206
rect 131 1210 135 1211
rect 131 1205 135 1206
rect 347 1210 351 1211
rect 347 1205 351 1206
rect 563 1210 567 1211
rect 563 1205 567 1206
rect 571 1210 575 1211
rect 571 1205 575 1206
rect 779 1210 783 1211
rect 779 1205 783 1206
rect 971 1210 975 1211
rect 971 1205 975 1206
rect 987 1210 991 1211
rect 987 1205 991 1206
rect 1147 1210 1151 1211
rect 1147 1205 1151 1206
rect 1195 1210 1199 1211
rect 1195 1205 1199 1206
rect 1315 1210 1319 1211
rect 1315 1205 1319 1206
rect 1395 1210 1399 1211
rect 1395 1205 1399 1206
rect 1483 1210 1487 1211
rect 1483 1205 1487 1206
rect 1603 1210 1607 1211
rect 1603 1205 1607 1206
rect 1643 1210 1647 1211
rect 1643 1205 1647 1206
rect 1787 1210 1791 1211
rect 1787 1205 1791 1206
rect 1935 1210 1939 1211
rect 1935 1205 1939 1206
rect 112 1145 114 1205
rect 110 1144 116 1145
rect 132 1144 134 1205
rect 348 1144 350 1205
rect 564 1144 566 1205
rect 780 1144 782 1205
rect 988 1144 990 1205
rect 1196 1144 1198 1205
rect 1396 1144 1398 1205
rect 1604 1144 1606 1205
rect 1788 1144 1790 1205
rect 1936 1145 1938 1205
rect 1976 1187 1978 1259
rect 3244 1187 3246 1260
rect 3380 1187 3382 1260
rect 3516 1187 3518 1260
rect 3652 1187 3654 1260
rect 3798 1259 3804 1260
rect 3800 1187 3802 1259
rect 3840 1203 3842 1275
rect 3860 1203 3862 1276
rect 4148 1203 4150 1276
rect 4444 1203 4446 1276
rect 4724 1203 4726 1276
rect 4996 1203 4998 1276
rect 5260 1203 5262 1276
rect 5516 1203 5518 1276
rect 5662 1275 5668 1276
rect 5664 1203 5666 1275
rect 3839 1202 3843 1203
rect 3839 1197 3843 1198
rect 3859 1202 3863 1203
rect 3859 1197 3863 1198
rect 4147 1202 4151 1203
rect 4147 1197 4151 1198
rect 4427 1202 4431 1203
rect 4427 1197 4431 1198
rect 4443 1202 4447 1203
rect 4443 1197 4447 1198
rect 4563 1202 4567 1203
rect 4563 1197 4567 1198
rect 4699 1202 4703 1203
rect 4699 1197 4703 1198
rect 4723 1202 4727 1203
rect 4723 1197 4727 1198
rect 4835 1202 4839 1203
rect 4835 1197 4839 1198
rect 4971 1202 4975 1203
rect 4971 1197 4975 1198
rect 4995 1202 4999 1203
rect 4995 1197 4999 1198
rect 5107 1202 5111 1203
rect 5107 1197 5111 1198
rect 5243 1202 5247 1203
rect 5243 1197 5247 1198
rect 5259 1202 5263 1203
rect 5259 1197 5263 1198
rect 5379 1202 5383 1203
rect 5379 1197 5383 1198
rect 5515 1202 5519 1203
rect 5515 1197 5519 1198
rect 5663 1202 5667 1203
rect 5663 1197 5667 1198
rect 1975 1186 1979 1187
rect 1975 1181 1979 1182
rect 1995 1186 1999 1187
rect 1995 1181 1999 1182
rect 2227 1186 2231 1187
rect 2227 1181 2231 1182
rect 2467 1186 2471 1187
rect 2467 1181 2471 1182
rect 2691 1186 2695 1187
rect 2691 1181 2695 1182
rect 2907 1186 2911 1187
rect 2907 1181 2911 1182
rect 3107 1186 3111 1187
rect 3107 1181 3111 1182
rect 3243 1186 3247 1187
rect 3243 1181 3247 1182
rect 3299 1186 3303 1187
rect 3299 1181 3303 1182
rect 3379 1186 3383 1187
rect 3379 1181 3383 1182
rect 3483 1186 3487 1187
rect 3483 1181 3487 1182
rect 3515 1186 3519 1187
rect 3515 1181 3519 1182
rect 3651 1186 3655 1187
rect 3651 1181 3655 1182
rect 3799 1186 3803 1187
rect 3799 1181 3803 1182
rect 1934 1144 1940 1145
rect 110 1140 111 1144
rect 115 1140 116 1144
rect 110 1139 116 1140
rect 130 1143 136 1144
rect 130 1139 131 1143
rect 135 1139 136 1143
rect 130 1138 136 1139
rect 346 1143 352 1144
rect 346 1139 347 1143
rect 351 1139 352 1143
rect 346 1138 352 1139
rect 562 1143 568 1144
rect 562 1139 563 1143
rect 567 1139 568 1143
rect 562 1138 568 1139
rect 778 1143 784 1144
rect 778 1139 779 1143
rect 783 1139 784 1143
rect 778 1138 784 1139
rect 986 1143 992 1144
rect 986 1139 987 1143
rect 991 1139 992 1143
rect 986 1138 992 1139
rect 1194 1143 1200 1144
rect 1194 1139 1195 1143
rect 1199 1139 1200 1143
rect 1194 1138 1200 1139
rect 1394 1143 1400 1144
rect 1394 1139 1395 1143
rect 1399 1139 1400 1143
rect 1394 1138 1400 1139
rect 1602 1143 1608 1144
rect 1602 1139 1603 1143
rect 1607 1139 1608 1143
rect 1602 1138 1608 1139
rect 1786 1143 1792 1144
rect 1786 1139 1787 1143
rect 1791 1139 1792 1143
rect 1934 1140 1935 1144
rect 1939 1140 1940 1144
rect 1934 1139 1940 1140
rect 1786 1138 1792 1139
rect 158 1128 164 1129
rect 110 1127 116 1128
rect 110 1123 111 1127
rect 115 1123 116 1127
rect 158 1124 159 1128
rect 163 1124 164 1128
rect 158 1123 164 1124
rect 374 1128 380 1129
rect 374 1124 375 1128
rect 379 1124 380 1128
rect 374 1123 380 1124
rect 590 1128 596 1129
rect 590 1124 591 1128
rect 595 1124 596 1128
rect 590 1123 596 1124
rect 806 1128 812 1129
rect 806 1124 807 1128
rect 811 1124 812 1128
rect 806 1123 812 1124
rect 1014 1128 1020 1129
rect 1014 1124 1015 1128
rect 1019 1124 1020 1128
rect 1014 1123 1020 1124
rect 1222 1128 1228 1129
rect 1222 1124 1223 1128
rect 1227 1124 1228 1128
rect 1222 1123 1228 1124
rect 1422 1128 1428 1129
rect 1422 1124 1423 1128
rect 1427 1124 1428 1128
rect 1422 1123 1428 1124
rect 1630 1128 1636 1129
rect 1630 1124 1631 1128
rect 1635 1124 1636 1128
rect 1630 1123 1636 1124
rect 1814 1128 1820 1129
rect 1814 1124 1815 1128
rect 1819 1124 1820 1128
rect 1814 1123 1820 1124
rect 1934 1127 1940 1128
rect 1934 1123 1935 1127
rect 1939 1123 1940 1127
rect 110 1122 116 1123
rect 112 1075 114 1122
rect 160 1075 162 1123
rect 376 1075 378 1123
rect 592 1075 594 1123
rect 808 1075 810 1123
rect 1016 1075 1018 1123
rect 1224 1075 1226 1123
rect 1424 1075 1426 1123
rect 1632 1075 1634 1123
rect 1816 1075 1818 1123
rect 1934 1122 1940 1123
rect 1936 1075 1938 1122
rect 1976 1121 1978 1181
rect 1974 1120 1980 1121
rect 1996 1120 1998 1181
rect 2228 1120 2230 1181
rect 2468 1120 2470 1181
rect 2692 1120 2694 1181
rect 2908 1120 2910 1181
rect 3108 1120 3110 1181
rect 3300 1120 3302 1181
rect 3484 1120 3486 1181
rect 3652 1120 3654 1181
rect 3800 1121 3802 1181
rect 3840 1137 3842 1197
rect 3838 1136 3844 1137
rect 4428 1136 4430 1197
rect 4564 1136 4566 1197
rect 4700 1136 4702 1197
rect 4836 1136 4838 1197
rect 4972 1136 4974 1197
rect 5108 1136 5110 1197
rect 5244 1136 5246 1197
rect 5380 1136 5382 1197
rect 5516 1136 5518 1197
rect 5664 1137 5666 1197
rect 5662 1136 5668 1137
rect 3838 1132 3839 1136
rect 3843 1132 3844 1136
rect 3838 1131 3844 1132
rect 4426 1135 4432 1136
rect 4426 1131 4427 1135
rect 4431 1131 4432 1135
rect 4426 1130 4432 1131
rect 4562 1135 4568 1136
rect 4562 1131 4563 1135
rect 4567 1131 4568 1135
rect 4562 1130 4568 1131
rect 4698 1135 4704 1136
rect 4698 1131 4699 1135
rect 4703 1131 4704 1135
rect 4698 1130 4704 1131
rect 4834 1135 4840 1136
rect 4834 1131 4835 1135
rect 4839 1131 4840 1135
rect 4834 1130 4840 1131
rect 4970 1135 4976 1136
rect 4970 1131 4971 1135
rect 4975 1131 4976 1135
rect 4970 1130 4976 1131
rect 5106 1135 5112 1136
rect 5106 1131 5107 1135
rect 5111 1131 5112 1135
rect 5106 1130 5112 1131
rect 5242 1135 5248 1136
rect 5242 1131 5243 1135
rect 5247 1131 5248 1135
rect 5242 1130 5248 1131
rect 5378 1135 5384 1136
rect 5378 1131 5379 1135
rect 5383 1131 5384 1135
rect 5378 1130 5384 1131
rect 5514 1135 5520 1136
rect 5514 1131 5515 1135
rect 5519 1131 5520 1135
rect 5662 1132 5663 1136
rect 5667 1132 5668 1136
rect 5662 1131 5668 1132
rect 5514 1130 5520 1131
rect 3798 1120 3804 1121
rect 4454 1120 4460 1121
rect 1974 1116 1975 1120
rect 1979 1116 1980 1120
rect 1974 1115 1980 1116
rect 1994 1119 2000 1120
rect 1994 1115 1995 1119
rect 1999 1115 2000 1119
rect 1994 1114 2000 1115
rect 2226 1119 2232 1120
rect 2226 1115 2227 1119
rect 2231 1115 2232 1119
rect 2226 1114 2232 1115
rect 2466 1119 2472 1120
rect 2466 1115 2467 1119
rect 2471 1115 2472 1119
rect 2466 1114 2472 1115
rect 2690 1119 2696 1120
rect 2690 1115 2691 1119
rect 2695 1115 2696 1119
rect 2690 1114 2696 1115
rect 2906 1119 2912 1120
rect 2906 1115 2907 1119
rect 2911 1115 2912 1119
rect 2906 1114 2912 1115
rect 3106 1119 3112 1120
rect 3106 1115 3107 1119
rect 3111 1115 3112 1119
rect 3106 1114 3112 1115
rect 3298 1119 3304 1120
rect 3298 1115 3299 1119
rect 3303 1115 3304 1119
rect 3298 1114 3304 1115
rect 3482 1119 3488 1120
rect 3482 1115 3483 1119
rect 3487 1115 3488 1119
rect 3482 1114 3488 1115
rect 3650 1119 3656 1120
rect 3650 1115 3651 1119
rect 3655 1115 3656 1119
rect 3798 1116 3799 1120
rect 3803 1116 3804 1120
rect 3798 1115 3804 1116
rect 3838 1119 3844 1120
rect 3838 1115 3839 1119
rect 3843 1115 3844 1119
rect 4454 1116 4455 1120
rect 4459 1116 4460 1120
rect 4454 1115 4460 1116
rect 4590 1120 4596 1121
rect 4590 1116 4591 1120
rect 4595 1116 4596 1120
rect 4590 1115 4596 1116
rect 4726 1120 4732 1121
rect 4726 1116 4727 1120
rect 4731 1116 4732 1120
rect 4726 1115 4732 1116
rect 4862 1120 4868 1121
rect 4862 1116 4863 1120
rect 4867 1116 4868 1120
rect 4862 1115 4868 1116
rect 4998 1120 5004 1121
rect 4998 1116 4999 1120
rect 5003 1116 5004 1120
rect 4998 1115 5004 1116
rect 5134 1120 5140 1121
rect 5134 1116 5135 1120
rect 5139 1116 5140 1120
rect 5134 1115 5140 1116
rect 5270 1120 5276 1121
rect 5270 1116 5271 1120
rect 5275 1116 5276 1120
rect 5270 1115 5276 1116
rect 5406 1120 5412 1121
rect 5406 1116 5407 1120
rect 5411 1116 5412 1120
rect 5406 1115 5412 1116
rect 5542 1120 5548 1121
rect 5542 1116 5543 1120
rect 5547 1116 5548 1120
rect 5542 1115 5548 1116
rect 5662 1119 5668 1120
rect 5662 1115 5663 1119
rect 5667 1115 5668 1119
rect 3650 1114 3656 1115
rect 3838 1114 3844 1115
rect 2022 1104 2028 1105
rect 1974 1103 1980 1104
rect 1974 1099 1975 1103
rect 1979 1099 1980 1103
rect 2022 1100 2023 1104
rect 2027 1100 2028 1104
rect 2022 1099 2028 1100
rect 2254 1104 2260 1105
rect 2254 1100 2255 1104
rect 2259 1100 2260 1104
rect 2254 1099 2260 1100
rect 2494 1104 2500 1105
rect 2494 1100 2495 1104
rect 2499 1100 2500 1104
rect 2494 1099 2500 1100
rect 2718 1104 2724 1105
rect 2718 1100 2719 1104
rect 2723 1100 2724 1104
rect 2718 1099 2724 1100
rect 2934 1104 2940 1105
rect 2934 1100 2935 1104
rect 2939 1100 2940 1104
rect 2934 1099 2940 1100
rect 3134 1104 3140 1105
rect 3134 1100 3135 1104
rect 3139 1100 3140 1104
rect 3134 1099 3140 1100
rect 3326 1104 3332 1105
rect 3326 1100 3327 1104
rect 3331 1100 3332 1104
rect 3326 1099 3332 1100
rect 3510 1104 3516 1105
rect 3510 1100 3511 1104
rect 3515 1100 3516 1104
rect 3510 1099 3516 1100
rect 3678 1104 3684 1105
rect 3678 1100 3679 1104
rect 3683 1100 3684 1104
rect 3678 1099 3684 1100
rect 3798 1103 3804 1104
rect 3798 1099 3799 1103
rect 3803 1099 3804 1103
rect 1974 1098 1980 1099
rect 1976 1075 1978 1098
rect 2024 1075 2026 1099
rect 2256 1075 2258 1099
rect 2496 1075 2498 1099
rect 2720 1075 2722 1099
rect 2936 1075 2938 1099
rect 3136 1075 3138 1099
rect 3328 1075 3330 1099
rect 3512 1075 3514 1099
rect 3680 1075 3682 1099
rect 3798 1098 3804 1099
rect 3800 1075 3802 1098
rect 3840 1075 3842 1114
rect 4456 1075 4458 1115
rect 4592 1075 4594 1115
rect 4728 1075 4730 1115
rect 4864 1075 4866 1115
rect 5000 1075 5002 1115
rect 5136 1075 5138 1115
rect 5272 1075 5274 1115
rect 5408 1075 5410 1115
rect 5544 1075 5546 1115
rect 5662 1114 5668 1115
rect 5664 1075 5666 1114
rect 111 1074 115 1075
rect 111 1069 115 1070
rect 159 1074 163 1075
rect 159 1069 163 1070
rect 375 1074 379 1075
rect 375 1069 379 1070
rect 471 1074 475 1075
rect 471 1069 475 1070
rect 591 1074 595 1075
rect 591 1069 595 1070
rect 607 1074 611 1075
rect 607 1069 611 1070
rect 743 1074 747 1075
rect 743 1069 747 1070
rect 807 1074 811 1075
rect 807 1069 811 1070
rect 887 1074 891 1075
rect 887 1069 891 1070
rect 1015 1074 1019 1075
rect 1015 1069 1019 1070
rect 1031 1074 1035 1075
rect 1031 1069 1035 1070
rect 1223 1074 1227 1075
rect 1223 1069 1227 1070
rect 1423 1074 1427 1075
rect 1423 1069 1427 1070
rect 1631 1074 1635 1075
rect 1631 1069 1635 1070
rect 1815 1074 1819 1075
rect 1815 1069 1819 1070
rect 1935 1074 1939 1075
rect 1935 1069 1939 1070
rect 1975 1074 1979 1075
rect 1975 1069 1979 1070
rect 2023 1074 2027 1075
rect 2023 1069 2027 1070
rect 2183 1074 2187 1075
rect 2183 1069 2187 1070
rect 2255 1074 2259 1075
rect 2255 1069 2259 1070
rect 2319 1074 2323 1075
rect 2319 1069 2323 1070
rect 2455 1074 2459 1075
rect 2455 1069 2459 1070
rect 2495 1074 2499 1075
rect 2495 1069 2499 1070
rect 2599 1074 2603 1075
rect 2599 1069 2603 1070
rect 2719 1074 2723 1075
rect 2719 1069 2723 1070
rect 2743 1074 2747 1075
rect 2743 1069 2747 1070
rect 2887 1074 2891 1075
rect 2887 1069 2891 1070
rect 2935 1074 2939 1075
rect 2935 1069 2939 1070
rect 3031 1074 3035 1075
rect 3031 1069 3035 1070
rect 3135 1074 3139 1075
rect 3135 1069 3139 1070
rect 3175 1074 3179 1075
rect 3175 1069 3179 1070
rect 3319 1074 3323 1075
rect 3319 1069 3323 1070
rect 3327 1074 3331 1075
rect 3327 1069 3331 1070
rect 3463 1074 3467 1075
rect 3463 1069 3467 1070
rect 3511 1074 3515 1075
rect 3511 1069 3515 1070
rect 3679 1074 3683 1075
rect 3679 1069 3683 1070
rect 3799 1074 3803 1075
rect 3799 1069 3803 1070
rect 3839 1074 3843 1075
rect 3839 1069 3843 1070
rect 4367 1074 4371 1075
rect 4367 1069 4371 1070
rect 4455 1074 4459 1075
rect 4455 1069 4459 1070
rect 4503 1074 4507 1075
rect 4503 1069 4507 1070
rect 4591 1074 4595 1075
rect 4591 1069 4595 1070
rect 4639 1074 4643 1075
rect 4639 1069 4643 1070
rect 4727 1074 4731 1075
rect 4727 1069 4731 1070
rect 4775 1074 4779 1075
rect 4775 1069 4779 1070
rect 4863 1074 4867 1075
rect 4863 1069 4867 1070
rect 4911 1074 4915 1075
rect 4911 1069 4915 1070
rect 4999 1074 5003 1075
rect 4999 1069 5003 1070
rect 5135 1074 5139 1075
rect 5135 1069 5139 1070
rect 5271 1074 5275 1075
rect 5271 1069 5275 1070
rect 5407 1074 5411 1075
rect 5407 1069 5411 1070
rect 5543 1074 5547 1075
rect 5543 1069 5547 1070
rect 5663 1074 5667 1075
rect 5663 1069 5667 1070
rect 112 1046 114 1069
rect 110 1045 116 1046
rect 472 1045 474 1069
rect 608 1045 610 1069
rect 744 1045 746 1069
rect 888 1045 890 1069
rect 1032 1045 1034 1069
rect 1936 1046 1938 1069
rect 1976 1046 1978 1069
rect 1934 1045 1940 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 470 1044 476 1045
rect 470 1040 471 1044
rect 475 1040 476 1044
rect 470 1039 476 1040
rect 606 1044 612 1045
rect 606 1040 607 1044
rect 611 1040 612 1044
rect 606 1039 612 1040
rect 742 1044 748 1045
rect 742 1040 743 1044
rect 747 1040 748 1044
rect 742 1039 748 1040
rect 886 1044 892 1045
rect 886 1040 887 1044
rect 891 1040 892 1044
rect 886 1039 892 1040
rect 1030 1044 1036 1045
rect 1030 1040 1031 1044
rect 1035 1040 1036 1044
rect 1934 1041 1935 1045
rect 1939 1041 1940 1045
rect 1934 1040 1940 1041
rect 1974 1045 1980 1046
rect 2184 1045 2186 1069
rect 2320 1045 2322 1069
rect 2456 1045 2458 1069
rect 2600 1045 2602 1069
rect 2744 1045 2746 1069
rect 2888 1045 2890 1069
rect 3032 1045 3034 1069
rect 3176 1045 3178 1069
rect 3320 1045 3322 1069
rect 3464 1045 3466 1069
rect 3800 1046 3802 1069
rect 3840 1046 3842 1069
rect 3798 1045 3804 1046
rect 1974 1041 1975 1045
rect 1979 1041 1980 1045
rect 1974 1040 1980 1041
rect 2182 1044 2188 1045
rect 2182 1040 2183 1044
rect 2187 1040 2188 1044
rect 1030 1039 1036 1040
rect 2182 1039 2188 1040
rect 2318 1044 2324 1045
rect 2318 1040 2319 1044
rect 2323 1040 2324 1044
rect 2318 1039 2324 1040
rect 2454 1044 2460 1045
rect 2454 1040 2455 1044
rect 2459 1040 2460 1044
rect 2454 1039 2460 1040
rect 2598 1044 2604 1045
rect 2598 1040 2599 1044
rect 2603 1040 2604 1044
rect 2598 1039 2604 1040
rect 2742 1044 2748 1045
rect 2742 1040 2743 1044
rect 2747 1040 2748 1044
rect 2742 1039 2748 1040
rect 2886 1044 2892 1045
rect 2886 1040 2887 1044
rect 2891 1040 2892 1044
rect 2886 1039 2892 1040
rect 3030 1044 3036 1045
rect 3030 1040 3031 1044
rect 3035 1040 3036 1044
rect 3030 1039 3036 1040
rect 3174 1044 3180 1045
rect 3174 1040 3175 1044
rect 3179 1040 3180 1044
rect 3174 1039 3180 1040
rect 3318 1044 3324 1045
rect 3318 1040 3319 1044
rect 3323 1040 3324 1044
rect 3318 1039 3324 1040
rect 3462 1044 3468 1045
rect 3462 1040 3463 1044
rect 3467 1040 3468 1044
rect 3798 1041 3799 1045
rect 3803 1041 3804 1045
rect 3798 1040 3804 1041
rect 3838 1045 3844 1046
rect 4368 1045 4370 1069
rect 4504 1045 4506 1069
rect 4640 1045 4642 1069
rect 4776 1045 4778 1069
rect 4912 1045 4914 1069
rect 5664 1046 5666 1069
rect 5662 1045 5668 1046
rect 3838 1041 3839 1045
rect 3843 1041 3844 1045
rect 3838 1040 3844 1041
rect 4366 1044 4372 1045
rect 4366 1040 4367 1044
rect 4371 1040 4372 1044
rect 3462 1039 3468 1040
rect 4366 1039 4372 1040
rect 4502 1044 4508 1045
rect 4502 1040 4503 1044
rect 4507 1040 4508 1044
rect 4502 1039 4508 1040
rect 4638 1044 4644 1045
rect 4638 1040 4639 1044
rect 4643 1040 4644 1044
rect 4638 1039 4644 1040
rect 4774 1044 4780 1045
rect 4774 1040 4775 1044
rect 4779 1040 4780 1044
rect 4774 1039 4780 1040
rect 4910 1044 4916 1045
rect 4910 1040 4911 1044
rect 4915 1040 4916 1044
rect 5662 1041 5663 1045
rect 5667 1041 5668 1045
rect 5662 1040 5668 1041
rect 4910 1039 4916 1040
rect 442 1029 448 1030
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 442 1025 443 1029
rect 447 1025 448 1029
rect 442 1024 448 1025
rect 578 1029 584 1030
rect 578 1025 579 1029
rect 583 1025 584 1029
rect 578 1024 584 1025
rect 714 1029 720 1030
rect 714 1025 715 1029
rect 719 1025 720 1029
rect 714 1024 720 1025
rect 858 1029 864 1030
rect 858 1025 859 1029
rect 863 1025 864 1029
rect 858 1024 864 1025
rect 1002 1029 1008 1030
rect 2154 1029 2160 1030
rect 1002 1025 1003 1029
rect 1007 1025 1008 1029
rect 1002 1024 1008 1025
rect 1934 1028 1940 1029
rect 1934 1024 1935 1028
rect 1939 1024 1940 1028
rect 110 1023 116 1024
rect 112 951 114 1023
rect 444 951 446 1024
rect 580 951 582 1024
rect 716 951 718 1024
rect 860 951 862 1024
rect 1004 951 1006 1024
rect 1934 1023 1940 1024
rect 1974 1028 1980 1029
rect 1974 1024 1975 1028
rect 1979 1024 1980 1028
rect 2154 1025 2155 1029
rect 2159 1025 2160 1029
rect 2154 1024 2160 1025
rect 2290 1029 2296 1030
rect 2290 1025 2291 1029
rect 2295 1025 2296 1029
rect 2290 1024 2296 1025
rect 2426 1029 2432 1030
rect 2426 1025 2427 1029
rect 2431 1025 2432 1029
rect 2426 1024 2432 1025
rect 2570 1029 2576 1030
rect 2570 1025 2571 1029
rect 2575 1025 2576 1029
rect 2570 1024 2576 1025
rect 2714 1029 2720 1030
rect 2714 1025 2715 1029
rect 2719 1025 2720 1029
rect 2714 1024 2720 1025
rect 2858 1029 2864 1030
rect 2858 1025 2859 1029
rect 2863 1025 2864 1029
rect 2858 1024 2864 1025
rect 3002 1029 3008 1030
rect 3002 1025 3003 1029
rect 3007 1025 3008 1029
rect 3002 1024 3008 1025
rect 3146 1029 3152 1030
rect 3146 1025 3147 1029
rect 3151 1025 3152 1029
rect 3146 1024 3152 1025
rect 3290 1029 3296 1030
rect 3290 1025 3291 1029
rect 3295 1025 3296 1029
rect 3290 1024 3296 1025
rect 3434 1029 3440 1030
rect 4338 1029 4344 1030
rect 3434 1025 3435 1029
rect 3439 1025 3440 1029
rect 3434 1024 3440 1025
rect 3798 1028 3804 1029
rect 3798 1024 3799 1028
rect 3803 1024 3804 1028
rect 1974 1023 1980 1024
rect 1936 951 1938 1023
rect 1976 951 1978 1023
rect 2156 951 2158 1024
rect 2292 951 2294 1024
rect 2428 951 2430 1024
rect 2572 951 2574 1024
rect 2716 951 2718 1024
rect 2860 951 2862 1024
rect 3004 951 3006 1024
rect 3148 951 3150 1024
rect 3292 951 3294 1024
rect 3436 951 3438 1024
rect 3798 1023 3804 1024
rect 3838 1028 3844 1029
rect 3838 1024 3839 1028
rect 3843 1024 3844 1028
rect 4338 1025 4339 1029
rect 4343 1025 4344 1029
rect 4338 1024 4344 1025
rect 4474 1029 4480 1030
rect 4474 1025 4475 1029
rect 4479 1025 4480 1029
rect 4474 1024 4480 1025
rect 4610 1029 4616 1030
rect 4610 1025 4611 1029
rect 4615 1025 4616 1029
rect 4610 1024 4616 1025
rect 4746 1029 4752 1030
rect 4746 1025 4747 1029
rect 4751 1025 4752 1029
rect 4746 1024 4752 1025
rect 4882 1029 4888 1030
rect 4882 1025 4883 1029
rect 4887 1025 4888 1029
rect 4882 1024 4888 1025
rect 5662 1028 5668 1029
rect 5662 1024 5663 1028
rect 5667 1024 5668 1028
rect 3838 1023 3844 1024
rect 3800 951 3802 1023
rect 3840 951 3842 1023
rect 4340 951 4342 1024
rect 4476 951 4478 1024
rect 4612 951 4614 1024
rect 4748 951 4750 1024
rect 4884 951 4886 1024
rect 5662 1023 5668 1024
rect 5664 951 5666 1023
rect 111 950 115 951
rect 111 945 115 946
rect 259 950 263 951
rect 259 945 263 946
rect 395 950 399 951
rect 395 945 399 946
rect 443 950 447 951
rect 443 945 447 946
rect 531 950 535 951
rect 531 945 535 946
rect 579 950 583 951
rect 579 945 583 946
rect 667 950 671 951
rect 667 945 671 946
rect 715 950 719 951
rect 715 945 719 946
rect 803 950 807 951
rect 803 945 807 946
rect 859 950 863 951
rect 859 945 863 946
rect 939 950 943 951
rect 939 945 943 946
rect 1003 950 1007 951
rect 1003 945 1007 946
rect 1935 950 1939 951
rect 1935 945 1939 946
rect 1975 950 1979 951
rect 1975 945 1979 946
rect 1995 950 1999 951
rect 1995 945 1999 946
rect 2131 950 2135 951
rect 2131 945 2135 946
rect 2155 950 2159 951
rect 2155 945 2159 946
rect 2267 950 2271 951
rect 2267 945 2271 946
rect 2291 950 2295 951
rect 2291 945 2295 946
rect 2403 950 2407 951
rect 2403 945 2407 946
rect 2427 950 2431 951
rect 2427 945 2431 946
rect 2539 950 2543 951
rect 2539 945 2543 946
rect 2571 950 2575 951
rect 2571 945 2575 946
rect 2675 950 2679 951
rect 2675 945 2679 946
rect 2715 950 2719 951
rect 2715 945 2719 946
rect 2811 950 2815 951
rect 2811 945 2815 946
rect 2859 950 2863 951
rect 2859 945 2863 946
rect 2947 950 2951 951
rect 2947 945 2951 946
rect 3003 950 3007 951
rect 3003 945 3007 946
rect 3083 950 3087 951
rect 3083 945 3087 946
rect 3147 950 3151 951
rect 3147 945 3151 946
rect 3219 950 3223 951
rect 3219 945 3223 946
rect 3291 950 3295 951
rect 3291 945 3295 946
rect 3355 950 3359 951
rect 3355 945 3359 946
rect 3435 950 3439 951
rect 3435 945 3439 946
rect 3491 950 3495 951
rect 3491 945 3495 946
rect 3799 950 3803 951
rect 3799 945 3803 946
rect 3839 950 3843 951
rect 3839 945 3843 946
rect 4019 950 4023 951
rect 4019 945 4023 946
rect 4155 950 4159 951
rect 4155 945 4159 946
rect 4291 950 4295 951
rect 4291 945 4295 946
rect 4339 950 4343 951
rect 4339 945 4343 946
rect 4427 950 4431 951
rect 4427 945 4431 946
rect 4475 950 4479 951
rect 4475 945 4479 946
rect 4563 950 4567 951
rect 4563 945 4567 946
rect 4611 950 4615 951
rect 4611 945 4615 946
rect 4699 950 4703 951
rect 4699 945 4703 946
rect 4747 950 4751 951
rect 4747 945 4751 946
rect 4883 950 4887 951
rect 4883 945 4887 946
rect 5663 950 5667 951
rect 5663 945 5667 946
rect 112 885 114 945
rect 110 884 116 885
rect 260 884 262 945
rect 396 884 398 945
rect 532 884 534 945
rect 668 884 670 945
rect 804 884 806 945
rect 940 884 942 945
rect 1936 885 1938 945
rect 1976 885 1978 945
rect 1934 884 1940 885
rect 110 880 111 884
rect 115 880 116 884
rect 110 879 116 880
rect 258 883 264 884
rect 258 879 259 883
rect 263 879 264 883
rect 258 878 264 879
rect 394 883 400 884
rect 394 879 395 883
rect 399 879 400 883
rect 394 878 400 879
rect 530 883 536 884
rect 530 879 531 883
rect 535 879 536 883
rect 530 878 536 879
rect 666 883 672 884
rect 666 879 667 883
rect 671 879 672 883
rect 666 878 672 879
rect 802 883 808 884
rect 802 879 803 883
rect 807 879 808 883
rect 802 878 808 879
rect 938 883 944 884
rect 938 879 939 883
rect 943 879 944 883
rect 1934 880 1935 884
rect 1939 880 1940 884
rect 1934 879 1940 880
rect 1974 884 1980 885
rect 1996 884 1998 945
rect 2132 884 2134 945
rect 2268 884 2270 945
rect 2404 884 2406 945
rect 2540 884 2542 945
rect 2676 884 2678 945
rect 2812 884 2814 945
rect 2948 884 2950 945
rect 3084 884 3086 945
rect 3220 884 3222 945
rect 3356 884 3358 945
rect 3492 884 3494 945
rect 3800 885 3802 945
rect 3840 885 3842 945
rect 3798 884 3804 885
rect 1974 880 1975 884
rect 1979 880 1980 884
rect 1974 879 1980 880
rect 1994 883 2000 884
rect 1994 879 1995 883
rect 1999 879 2000 883
rect 938 878 944 879
rect 1994 878 2000 879
rect 2130 883 2136 884
rect 2130 879 2131 883
rect 2135 879 2136 883
rect 2130 878 2136 879
rect 2266 883 2272 884
rect 2266 879 2267 883
rect 2271 879 2272 883
rect 2266 878 2272 879
rect 2402 883 2408 884
rect 2402 879 2403 883
rect 2407 879 2408 883
rect 2402 878 2408 879
rect 2538 883 2544 884
rect 2538 879 2539 883
rect 2543 879 2544 883
rect 2538 878 2544 879
rect 2674 883 2680 884
rect 2674 879 2675 883
rect 2679 879 2680 883
rect 2674 878 2680 879
rect 2810 883 2816 884
rect 2810 879 2811 883
rect 2815 879 2816 883
rect 2810 878 2816 879
rect 2946 883 2952 884
rect 2946 879 2947 883
rect 2951 879 2952 883
rect 2946 878 2952 879
rect 3082 883 3088 884
rect 3082 879 3083 883
rect 3087 879 3088 883
rect 3082 878 3088 879
rect 3218 883 3224 884
rect 3218 879 3219 883
rect 3223 879 3224 883
rect 3218 878 3224 879
rect 3354 883 3360 884
rect 3354 879 3355 883
rect 3359 879 3360 883
rect 3354 878 3360 879
rect 3490 883 3496 884
rect 3490 879 3491 883
rect 3495 879 3496 883
rect 3798 880 3799 884
rect 3803 880 3804 884
rect 3798 879 3804 880
rect 3838 884 3844 885
rect 4020 884 4022 945
rect 4156 884 4158 945
rect 4292 884 4294 945
rect 4428 884 4430 945
rect 4564 884 4566 945
rect 4700 884 4702 945
rect 5664 885 5666 945
rect 5662 884 5668 885
rect 3838 880 3839 884
rect 3843 880 3844 884
rect 3838 879 3844 880
rect 4018 883 4024 884
rect 4018 879 4019 883
rect 4023 879 4024 883
rect 3490 878 3496 879
rect 4018 878 4024 879
rect 4154 883 4160 884
rect 4154 879 4155 883
rect 4159 879 4160 883
rect 4154 878 4160 879
rect 4290 883 4296 884
rect 4290 879 4291 883
rect 4295 879 4296 883
rect 4290 878 4296 879
rect 4426 883 4432 884
rect 4426 879 4427 883
rect 4431 879 4432 883
rect 4426 878 4432 879
rect 4562 883 4568 884
rect 4562 879 4563 883
rect 4567 879 4568 883
rect 4562 878 4568 879
rect 4698 883 4704 884
rect 4698 879 4699 883
rect 4703 879 4704 883
rect 5662 880 5663 884
rect 5667 880 5668 884
rect 5662 879 5668 880
rect 4698 878 4704 879
rect 286 868 292 869
rect 110 867 116 868
rect 110 863 111 867
rect 115 863 116 867
rect 286 864 287 868
rect 291 864 292 868
rect 286 863 292 864
rect 422 868 428 869
rect 422 864 423 868
rect 427 864 428 868
rect 422 863 428 864
rect 558 868 564 869
rect 558 864 559 868
rect 563 864 564 868
rect 558 863 564 864
rect 694 868 700 869
rect 694 864 695 868
rect 699 864 700 868
rect 694 863 700 864
rect 830 868 836 869
rect 830 864 831 868
rect 835 864 836 868
rect 830 863 836 864
rect 966 868 972 869
rect 2022 868 2028 869
rect 966 864 967 868
rect 971 864 972 868
rect 966 863 972 864
rect 1934 867 1940 868
rect 1934 863 1935 867
rect 1939 863 1940 867
rect 110 862 116 863
rect 112 827 114 862
rect 288 827 290 863
rect 424 827 426 863
rect 560 827 562 863
rect 696 827 698 863
rect 832 827 834 863
rect 968 827 970 863
rect 1934 862 1940 863
rect 1974 867 1980 868
rect 1974 863 1975 867
rect 1979 863 1980 867
rect 2022 864 2023 868
rect 2027 864 2028 868
rect 2022 863 2028 864
rect 2158 868 2164 869
rect 2158 864 2159 868
rect 2163 864 2164 868
rect 2158 863 2164 864
rect 2294 868 2300 869
rect 2294 864 2295 868
rect 2299 864 2300 868
rect 2294 863 2300 864
rect 2430 868 2436 869
rect 2430 864 2431 868
rect 2435 864 2436 868
rect 2430 863 2436 864
rect 2566 868 2572 869
rect 2566 864 2567 868
rect 2571 864 2572 868
rect 2566 863 2572 864
rect 2702 868 2708 869
rect 2702 864 2703 868
rect 2707 864 2708 868
rect 2702 863 2708 864
rect 2838 868 2844 869
rect 2838 864 2839 868
rect 2843 864 2844 868
rect 2838 863 2844 864
rect 2974 868 2980 869
rect 2974 864 2975 868
rect 2979 864 2980 868
rect 2974 863 2980 864
rect 3110 868 3116 869
rect 3110 864 3111 868
rect 3115 864 3116 868
rect 3110 863 3116 864
rect 3246 868 3252 869
rect 3246 864 3247 868
rect 3251 864 3252 868
rect 3246 863 3252 864
rect 3382 868 3388 869
rect 3382 864 3383 868
rect 3387 864 3388 868
rect 3382 863 3388 864
rect 3518 868 3524 869
rect 4046 868 4052 869
rect 3518 864 3519 868
rect 3523 864 3524 868
rect 3518 863 3524 864
rect 3798 867 3804 868
rect 3798 863 3799 867
rect 3803 863 3804 867
rect 1974 862 1980 863
rect 1936 827 1938 862
rect 1976 839 1978 862
rect 2024 839 2026 863
rect 2160 839 2162 863
rect 2296 839 2298 863
rect 2432 839 2434 863
rect 2568 839 2570 863
rect 2704 839 2706 863
rect 2840 839 2842 863
rect 2976 839 2978 863
rect 3112 839 3114 863
rect 3248 839 3250 863
rect 3384 839 3386 863
rect 3520 839 3522 863
rect 3798 862 3804 863
rect 3838 867 3844 868
rect 3838 863 3839 867
rect 3843 863 3844 867
rect 4046 864 4047 868
rect 4051 864 4052 868
rect 4046 863 4052 864
rect 4182 868 4188 869
rect 4182 864 4183 868
rect 4187 864 4188 868
rect 4182 863 4188 864
rect 4318 868 4324 869
rect 4318 864 4319 868
rect 4323 864 4324 868
rect 4318 863 4324 864
rect 4454 868 4460 869
rect 4454 864 4455 868
rect 4459 864 4460 868
rect 4454 863 4460 864
rect 4590 868 4596 869
rect 4590 864 4591 868
rect 4595 864 4596 868
rect 4590 863 4596 864
rect 4726 868 4732 869
rect 4726 864 4727 868
rect 4731 864 4732 868
rect 4726 863 4732 864
rect 5662 867 5668 868
rect 5662 863 5663 867
rect 5667 863 5668 867
rect 3838 862 3844 863
rect 3800 839 3802 862
rect 1975 838 1979 839
rect 1975 833 1979 834
rect 2023 838 2027 839
rect 2023 833 2027 834
rect 2159 838 2163 839
rect 2159 833 2163 834
rect 2167 838 2171 839
rect 2167 833 2171 834
rect 2295 838 2299 839
rect 2295 833 2299 834
rect 2335 838 2339 839
rect 2335 833 2339 834
rect 2431 838 2435 839
rect 2431 833 2435 834
rect 2495 838 2499 839
rect 2495 833 2499 834
rect 2567 838 2571 839
rect 2567 833 2571 834
rect 2655 838 2659 839
rect 2655 833 2659 834
rect 2703 838 2707 839
rect 2703 833 2707 834
rect 2823 838 2827 839
rect 2823 833 2827 834
rect 2839 838 2843 839
rect 2839 833 2843 834
rect 2975 838 2979 839
rect 2975 833 2979 834
rect 2991 838 2995 839
rect 2991 833 2995 834
rect 3111 838 3115 839
rect 3111 833 3115 834
rect 3247 838 3251 839
rect 3247 833 3251 834
rect 3383 838 3387 839
rect 3383 833 3387 834
rect 3519 838 3523 839
rect 3519 833 3523 834
rect 3799 838 3803 839
rect 3799 833 3803 834
rect 111 826 115 827
rect 111 821 115 822
rect 239 826 243 827
rect 239 821 243 822
rect 287 826 291 827
rect 287 821 291 822
rect 423 826 427 827
rect 423 821 427 822
rect 439 826 443 827
rect 439 821 443 822
rect 559 826 563 827
rect 559 821 563 822
rect 647 826 651 827
rect 647 821 651 822
rect 695 826 699 827
rect 695 821 699 822
rect 831 826 835 827
rect 831 821 835 822
rect 855 826 859 827
rect 855 821 859 822
rect 967 826 971 827
rect 967 821 971 822
rect 1063 826 1067 827
rect 1063 821 1067 822
rect 1935 826 1939 827
rect 1935 821 1939 822
rect 112 798 114 821
rect 110 797 116 798
rect 240 797 242 821
rect 440 797 442 821
rect 648 797 650 821
rect 856 797 858 821
rect 1064 797 1066 821
rect 1936 798 1938 821
rect 1976 810 1978 833
rect 1974 809 1980 810
rect 2024 809 2026 833
rect 2168 809 2170 833
rect 2336 809 2338 833
rect 2496 809 2498 833
rect 2656 809 2658 833
rect 2824 809 2826 833
rect 2992 809 2994 833
rect 3800 810 3802 833
rect 3840 823 3842 862
rect 4048 823 4050 863
rect 4184 823 4186 863
rect 4320 823 4322 863
rect 4456 823 4458 863
rect 4592 823 4594 863
rect 4728 823 4730 863
rect 5662 862 5668 863
rect 5664 823 5666 862
rect 3839 822 3843 823
rect 3839 817 3843 818
rect 3887 822 3891 823
rect 3887 817 3891 818
rect 4023 822 4027 823
rect 4023 817 4027 818
rect 4047 822 4051 823
rect 4047 817 4051 818
rect 4159 822 4163 823
rect 4159 817 4163 818
rect 4183 822 4187 823
rect 4183 817 4187 818
rect 4295 822 4299 823
rect 4295 817 4299 818
rect 4319 822 4323 823
rect 4319 817 4323 818
rect 4431 822 4435 823
rect 4431 817 4435 818
rect 4455 822 4459 823
rect 4455 817 4459 818
rect 4567 822 4571 823
rect 4567 817 4571 818
rect 4591 822 4595 823
rect 4591 817 4595 818
rect 4703 822 4707 823
rect 4703 817 4707 818
rect 4727 822 4731 823
rect 4727 817 4731 818
rect 4839 822 4843 823
rect 4839 817 4843 818
rect 5663 822 5667 823
rect 5663 817 5667 818
rect 3798 809 3804 810
rect 1974 805 1975 809
rect 1979 805 1980 809
rect 1974 804 1980 805
rect 2022 808 2028 809
rect 2022 804 2023 808
rect 2027 804 2028 808
rect 2022 803 2028 804
rect 2166 808 2172 809
rect 2166 804 2167 808
rect 2171 804 2172 808
rect 2166 803 2172 804
rect 2334 808 2340 809
rect 2334 804 2335 808
rect 2339 804 2340 808
rect 2334 803 2340 804
rect 2494 808 2500 809
rect 2494 804 2495 808
rect 2499 804 2500 808
rect 2494 803 2500 804
rect 2654 808 2660 809
rect 2654 804 2655 808
rect 2659 804 2660 808
rect 2654 803 2660 804
rect 2822 808 2828 809
rect 2822 804 2823 808
rect 2827 804 2828 808
rect 2822 803 2828 804
rect 2990 808 2996 809
rect 2990 804 2991 808
rect 2995 804 2996 808
rect 3798 805 3799 809
rect 3803 805 3804 809
rect 3798 804 3804 805
rect 2990 803 2996 804
rect 1934 797 1940 798
rect 110 793 111 797
rect 115 793 116 797
rect 110 792 116 793
rect 238 796 244 797
rect 238 792 239 796
rect 243 792 244 796
rect 238 791 244 792
rect 438 796 444 797
rect 438 792 439 796
rect 443 792 444 796
rect 438 791 444 792
rect 646 796 652 797
rect 646 792 647 796
rect 651 792 652 796
rect 646 791 652 792
rect 854 796 860 797
rect 854 792 855 796
rect 859 792 860 796
rect 854 791 860 792
rect 1062 796 1068 797
rect 1062 792 1063 796
rect 1067 792 1068 796
rect 1934 793 1935 797
rect 1939 793 1940 797
rect 3840 794 3842 817
rect 1994 793 2000 794
rect 1934 792 1940 793
rect 1974 792 1980 793
rect 1062 791 1068 792
rect 1974 788 1975 792
rect 1979 788 1980 792
rect 1994 789 1995 793
rect 1999 789 2000 793
rect 1994 788 2000 789
rect 2138 793 2144 794
rect 2138 789 2139 793
rect 2143 789 2144 793
rect 2138 788 2144 789
rect 2306 793 2312 794
rect 2306 789 2307 793
rect 2311 789 2312 793
rect 2306 788 2312 789
rect 2466 793 2472 794
rect 2466 789 2467 793
rect 2471 789 2472 793
rect 2466 788 2472 789
rect 2626 793 2632 794
rect 2626 789 2627 793
rect 2631 789 2632 793
rect 2626 788 2632 789
rect 2794 793 2800 794
rect 2794 789 2795 793
rect 2799 789 2800 793
rect 2794 788 2800 789
rect 2962 793 2968 794
rect 3838 793 3844 794
rect 3888 793 3890 817
rect 4024 793 4026 817
rect 4160 793 4162 817
rect 4296 793 4298 817
rect 4432 793 4434 817
rect 4568 793 4570 817
rect 4704 793 4706 817
rect 4840 793 4842 817
rect 5664 794 5666 817
rect 5662 793 5668 794
rect 2962 789 2963 793
rect 2967 789 2968 793
rect 2962 788 2968 789
rect 3798 792 3804 793
rect 3798 788 3799 792
rect 3803 788 3804 792
rect 3838 789 3839 793
rect 3843 789 3844 793
rect 3838 788 3844 789
rect 3886 792 3892 793
rect 3886 788 3887 792
rect 3891 788 3892 792
rect 1974 787 1980 788
rect 210 781 216 782
rect 110 780 116 781
rect 110 776 111 780
rect 115 776 116 780
rect 210 777 211 781
rect 215 777 216 781
rect 210 776 216 777
rect 410 781 416 782
rect 410 777 411 781
rect 415 777 416 781
rect 410 776 416 777
rect 618 781 624 782
rect 618 777 619 781
rect 623 777 624 781
rect 618 776 624 777
rect 826 781 832 782
rect 826 777 827 781
rect 831 777 832 781
rect 826 776 832 777
rect 1034 781 1040 782
rect 1034 777 1035 781
rect 1039 777 1040 781
rect 1034 776 1040 777
rect 1934 780 1940 781
rect 1934 776 1935 780
rect 1939 776 1940 780
rect 110 775 116 776
rect 112 695 114 775
rect 212 695 214 776
rect 412 695 414 776
rect 620 695 622 776
rect 828 695 830 776
rect 1036 695 1038 776
rect 1934 775 1940 776
rect 1936 695 1938 775
rect 1976 699 1978 787
rect 1996 699 1998 788
rect 2140 699 2142 788
rect 2308 699 2310 788
rect 2468 699 2470 788
rect 2628 699 2630 788
rect 2796 699 2798 788
rect 2964 699 2966 788
rect 3798 787 3804 788
rect 3886 787 3892 788
rect 4022 792 4028 793
rect 4022 788 4023 792
rect 4027 788 4028 792
rect 4022 787 4028 788
rect 4158 792 4164 793
rect 4158 788 4159 792
rect 4163 788 4164 792
rect 4158 787 4164 788
rect 4294 792 4300 793
rect 4294 788 4295 792
rect 4299 788 4300 792
rect 4294 787 4300 788
rect 4430 792 4436 793
rect 4430 788 4431 792
rect 4435 788 4436 792
rect 4430 787 4436 788
rect 4566 792 4572 793
rect 4566 788 4567 792
rect 4571 788 4572 792
rect 4566 787 4572 788
rect 4702 792 4708 793
rect 4702 788 4703 792
rect 4707 788 4708 792
rect 4702 787 4708 788
rect 4838 792 4844 793
rect 4838 788 4839 792
rect 4843 788 4844 792
rect 5662 789 5663 793
rect 5667 789 5668 793
rect 5662 788 5668 789
rect 4838 787 4844 788
rect 3800 699 3802 787
rect 3858 777 3864 778
rect 3838 776 3844 777
rect 3838 772 3839 776
rect 3843 772 3844 776
rect 3858 773 3859 777
rect 3863 773 3864 777
rect 3858 772 3864 773
rect 3994 777 4000 778
rect 3994 773 3995 777
rect 3999 773 4000 777
rect 3994 772 4000 773
rect 4130 777 4136 778
rect 4130 773 4131 777
rect 4135 773 4136 777
rect 4130 772 4136 773
rect 4266 777 4272 778
rect 4266 773 4267 777
rect 4271 773 4272 777
rect 4266 772 4272 773
rect 4402 777 4408 778
rect 4402 773 4403 777
rect 4407 773 4408 777
rect 4402 772 4408 773
rect 4538 777 4544 778
rect 4538 773 4539 777
rect 4543 773 4544 777
rect 4538 772 4544 773
rect 4674 777 4680 778
rect 4674 773 4675 777
rect 4679 773 4680 777
rect 4674 772 4680 773
rect 4810 777 4816 778
rect 4810 773 4811 777
rect 4815 773 4816 777
rect 4810 772 4816 773
rect 5662 776 5668 777
rect 5662 772 5663 776
rect 5667 772 5668 776
rect 3838 771 3844 772
rect 3840 711 3842 771
rect 3860 711 3862 772
rect 3996 711 3998 772
rect 4132 711 4134 772
rect 4268 711 4270 772
rect 4404 711 4406 772
rect 4540 711 4542 772
rect 4676 711 4678 772
rect 4812 711 4814 772
rect 5662 771 5668 772
rect 5664 711 5666 771
rect 3839 710 3843 711
rect 3839 705 3843 706
rect 3859 710 3863 711
rect 3859 705 3863 706
rect 3995 710 3999 711
rect 3995 705 3999 706
rect 4131 710 4135 711
rect 4131 705 4135 706
rect 4267 710 4271 711
rect 4267 705 4271 706
rect 4403 710 4407 711
rect 4403 705 4407 706
rect 4539 710 4543 711
rect 4539 705 4543 706
rect 4675 710 4679 711
rect 4675 705 4679 706
rect 4811 710 4815 711
rect 4811 705 4815 706
rect 4947 710 4951 711
rect 4947 705 4951 706
rect 5083 710 5087 711
rect 5083 705 5087 706
rect 5663 710 5667 711
rect 5663 705 5667 706
rect 1975 698 1979 699
rect 111 694 115 695
rect 111 689 115 690
rect 131 694 135 695
rect 131 689 135 690
rect 211 694 215 695
rect 211 689 215 690
rect 347 694 351 695
rect 347 689 351 690
rect 411 694 415 695
rect 411 689 415 690
rect 587 694 591 695
rect 587 689 591 690
rect 619 694 623 695
rect 619 689 623 690
rect 827 694 831 695
rect 827 689 831 690
rect 1035 694 1039 695
rect 1035 689 1039 690
rect 1067 694 1071 695
rect 1067 689 1071 690
rect 1315 694 1319 695
rect 1315 689 1319 690
rect 1563 694 1567 695
rect 1563 689 1567 690
rect 1787 694 1791 695
rect 1787 689 1791 690
rect 1935 694 1939 695
rect 1975 693 1979 694
rect 1995 698 1999 699
rect 1995 693 1999 694
rect 2139 698 2143 699
rect 2139 693 2143 694
rect 2299 698 2303 699
rect 2299 693 2303 694
rect 2307 698 2311 699
rect 2307 693 2311 694
rect 2467 698 2471 699
rect 2467 693 2471 694
rect 2627 698 2631 699
rect 2627 693 2631 694
rect 2635 698 2639 699
rect 2635 693 2639 694
rect 2795 698 2799 699
rect 2795 693 2799 694
rect 2963 698 2967 699
rect 2963 693 2967 694
rect 2979 698 2983 699
rect 2979 693 2983 694
rect 3323 698 3327 699
rect 3323 693 3327 694
rect 3651 698 3655 699
rect 3651 693 3655 694
rect 3799 698 3803 699
rect 3799 693 3803 694
rect 1935 689 1939 690
rect 112 629 114 689
rect 110 628 116 629
rect 132 628 134 689
rect 348 628 350 689
rect 588 628 590 689
rect 828 628 830 689
rect 1068 628 1070 689
rect 1316 628 1318 689
rect 1564 628 1566 689
rect 1788 628 1790 689
rect 1936 629 1938 689
rect 1976 633 1978 693
rect 1974 632 1980 633
rect 1996 632 1998 693
rect 2300 632 2302 693
rect 2636 632 2638 693
rect 2980 632 2982 693
rect 3324 632 3326 693
rect 3652 632 3654 693
rect 3800 633 3802 693
rect 3840 645 3842 705
rect 3838 644 3844 645
rect 3860 644 3862 705
rect 3996 644 3998 705
rect 4132 644 4134 705
rect 4268 644 4270 705
rect 4404 644 4406 705
rect 4540 644 4542 705
rect 4676 644 4678 705
rect 4812 644 4814 705
rect 4948 644 4950 705
rect 5084 644 5086 705
rect 5664 645 5666 705
rect 5662 644 5668 645
rect 3838 640 3839 644
rect 3843 640 3844 644
rect 3838 639 3844 640
rect 3858 643 3864 644
rect 3858 639 3859 643
rect 3863 639 3864 643
rect 3858 638 3864 639
rect 3994 643 4000 644
rect 3994 639 3995 643
rect 3999 639 4000 643
rect 3994 638 4000 639
rect 4130 643 4136 644
rect 4130 639 4131 643
rect 4135 639 4136 643
rect 4130 638 4136 639
rect 4266 643 4272 644
rect 4266 639 4267 643
rect 4271 639 4272 643
rect 4266 638 4272 639
rect 4402 643 4408 644
rect 4402 639 4403 643
rect 4407 639 4408 643
rect 4402 638 4408 639
rect 4538 643 4544 644
rect 4538 639 4539 643
rect 4543 639 4544 643
rect 4538 638 4544 639
rect 4674 643 4680 644
rect 4674 639 4675 643
rect 4679 639 4680 643
rect 4674 638 4680 639
rect 4810 643 4816 644
rect 4810 639 4811 643
rect 4815 639 4816 643
rect 4810 638 4816 639
rect 4946 643 4952 644
rect 4946 639 4947 643
rect 4951 639 4952 643
rect 4946 638 4952 639
rect 5082 643 5088 644
rect 5082 639 5083 643
rect 5087 639 5088 643
rect 5662 640 5663 644
rect 5667 640 5668 644
rect 5662 639 5668 640
rect 5082 638 5088 639
rect 3798 632 3804 633
rect 1934 628 1940 629
rect 110 624 111 628
rect 115 624 116 628
rect 110 623 116 624
rect 130 627 136 628
rect 130 623 131 627
rect 135 623 136 627
rect 130 622 136 623
rect 346 627 352 628
rect 346 623 347 627
rect 351 623 352 627
rect 346 622 352 623
rect 586 627 592 628
rect 586 623 587 627
rect 591 623 592 627
rect 586 622 592 623
rect 826 627 832 628
rect 826 623 827 627
rect 831 623 832 627
rect 826 622 832 623
rect 1066 627 1072 628
rect 1066 623 1067 627
rect 1071 623 1072 627
rect 1066 622 1072 623
rect 1314 627 1320 628
rect 1314 623 1315 627
rect 1319 623 1320 627
rect 1314 622 1320 623
rect 1562 627 1568 628
rect 1562 623 1563 627
rect 1567 623 1568 627
rect 1562 622 1568 623
rect 1786 627 1792 628
rect 1786 623 1787 627
rect 1791 623 1792 627
rect 1934 624 1935 628
rect 1939 624 1940 628
rect 1974 628 1975 632
rect 1979 628 1980 632
rect 1974 627 1980 628
rect 1994 631 2000 632
rect 1994 627 1995 631
rect 1999 627 2000 631
rect 1994 626 2000 627
rect 2298 631 2304 632
rect 2298 627 2299 631
rect 2303 627 2304 631
rect 2298 626 2304 627
rect 2634 631 2640 632
rect 2634 627 2635 631
rect 2639 627 2640 631
rect 2634 626 2640 627
rect 2978 631 2984 632
rect 2978 627 2979 631
rect 2983 627 2984 631
rect 2978 626 2984 627
rect 3322 631 3328 632
rect 3322 627 3323 631
rect 3327 627 3328 631
rect 3322 626 3328 627
rect 3650 631 3656 632
rect 3650 627 3651 631
rect 3655 627 3656 631
rect 3798 628 3799 632
rect 3803 628 3804 632
rect 3886 628 3892 629
rect 3798 627 3804 628
rect 3838 627 3844 628
rect 3650 626 3656 627
rect 1934 623 1940 624
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3886 624 3887 628
rect 3891 624 3892 628
rect 3886 623 3892 624
rect 4022 628 4028 629
rect 4022 624 4023 628
rect 4027 624 4028 628
rect 4022 623 4028 624
rect 4158 628 4164 629
rect 4158 624 4159 628
rect 4163 624 4164 628
rect 4158 623 4164 624
rect 4294 628 4300 629
rect 4294 624 4295 628
rect 4299 624 4300 628
rect 4294 623 4300 624
rect 4430 628 4436 629
rect 4430 624 4431 628
rect 4435 624 4436 628
rect 4430 623 4436 624
rect 4566 628 4572 629
rect 4566 624 4567 628
rect 4571 624 4572 628
rect 4566 623 4572 624
rect 4702 628 4708 629
rect 4702 624 4703 628
rect 4707 624 4708 628
rect 4702 623 4708 624
rect 4838 628 4844 629
rect 4838 624 4839 628
rect 4843 624 4844 628
rect 4838 623 4844 624
rect 4974 628 4980 629
rect 4974 624 4975 628
rect 4979 624 4980 628
rect 4974 623 4980 624
rect 5110 628 5116 629
rect 5110 624 5111 628
rect 5115 624 5116 628
rect 5110 623 5116 624
rect 5662 627 5668 628
rect 5662 623 5663 627
rect 5667 623 5668 627
rect 1786 622 1792 623
rect 3838 622 3844 623
rect 2022 616 2028 617
rect 1974 615 1980 616
rect 158 612 164 613
rect 110 611 116 612
rect 110 607 111 611
rect 115 607 116 611
rect 158 608 159 612
rect 163 608 164 612
rect 158 607 164 608
rect 374 612 380 613
rect 374 608 375 612
rect 379 608 380 612
rect 374 607 380 608
rect 614 612 620 613
rect 614 608 615 612
rect 619 608 620 612
rect 614 607 620 608
rect 854 612 860 613
rect 854 608 855 612
rect 859 608 860 612
rect 854 607 860 608
rect 1094 612 1100 613
rect 1094 608 1095 612
rect 1099 608 1100 612
rect 1094 607 1100 608
rect 1342 612 1348 613
rect 1342 608 1343 612
rect 1347 608 1348 612
rect 1342 607 1348 608
rect 1590 612 1596 613
rect 1590 608 1591 612
rect 1595 608 1596 612
rect 1590 607 1596 608
rect 1814 612 1820 613
rect 1814 608 1815 612
rect 1819 608 1820 612
rect 1814 607 1820 608
rect 1934 611 1940 612
rect 1934 607 1935 611
rect 1939 607 1940 611
rect 1974 611 1975 615
rect 1979 611 1980 615
rect 2022 612 2023 616
rect 2027 612 2028 616
rect 2022 611 2028 612
rect 2326 616 2332 617
rect 2326 612 2327 616
rect 2331 612 2332 616
rect 2326 611 2332 612
rect 2662 616 2668 617
rect 2662 612 2663 616
rect 2667 612 2668 616
rect 2662 611 2668 612
rect 3006 616 3012 617
rect 3006 612 3007 616
rect 3011 612 3012 616
rect 3006 611 3012 612
rect 3350 616 3356 617
rect 3350 612 3351 616
rect 3355 612 3356 616
rect 3350 611 3356 612
rect 3678 616 3684 617
rect 3678 612 3679 616
rect 3683 612 3684 616
rect 3678 611 3684 612
rect 3798 615 3804 616
rect 3798 611 3799 615
rect 3803 611 3804 615
rect 1974 610 1980 611
rect 110 606 116 607
rect 112 579 114 606
rect 160 579 162 607
rect 376 579 378 607
rect 616 579 618 607
rect 856 579 858 607
rect 1096 579 1098 607
rect 1344 579 1346 607
rect 1592 579 1594 607
rect 1816 579 1818 607
rect 1934 606 1940 607
rect 1936 579 1938 606
rect 1976 587 1978 610
rect 2024 587 2026 611
rect 2328 587 2330 611
rect 2664 587 2666 611
rect 3008 587 3010 611
rect 3352 587 3354 611
rect 3680 587 3682 611
rect 3798 610 3804 611
rect 3800 587 3802 610
rect 1975 586 1979 587
rect 1975 581 1979 582
rect 2023 586 2027 587
rect 2023 581 2027 582
rect 2327 586 2331 587
rect 2327 581 2331 582
rect 2335 586 2339 587
rect 2335 581 2339 582
rect 2527 586 2531 587
rect 2527 581 2531 582
rect 2663 586 2667 587
rect 2663 581 2667 582
rect 2711 586 2715 587
rect 2711 581 2715 582
rect 2887 586 2891 587
rect 2887 581 2891 582
rect 3007 586 3011 587
rect 3007 581 3011 582
rect 3063 586 3067 587
rect 3063 581 3067 582
rect 3231 586 3235 587
rect 3231 581 3235 582
rect 3351 586 3355 587
rect 3351 581 3355 582
rect 3407 586 3411 587
rect 3407 581 3411 582
rect 3583 586 3587 587
rect 3583 581 3587 582
rect 3679 586 3683 587
rect 3679 581 3683 582
rect 3799 586 3803 587
rect 3799 581 3803 582
rect 111 578 115 579
rect 111 573 115 574
rect 159 578 163 579
rect 159 573 163 574
rect 375 578 379 579
rect 375 573 379 574
rect 407 578 411 579
rect 407 573 411 574
rect 615 578 619 579
rect 615 573 619 574
rect 671 578 675 579
rect 671 573 675 574
rect 855 578 859 579
rect 855 573 859 574
rect 935 578 939 579
rect 935 573 939 574
rect 1095 578 1099 579
rect 1095 573 1099 574
rect 1191 578 1195 579
rect 1191 573 1195 574
rect 1343 578 1347 579
rect 1343 573 1347 574
rect 1447 578 1451 579
rect 1447 573 1451 574
rect 1591 578 1595 579
rect 1591 573 1595 574
rect 1711 578 1715 579
rect 1711 573 1715 574
rect 1815 578 1819 579
rect 1815 573 1819 574
rect 1935 578 1939 579
rect 1935 573 1939 574
rect 112 550 114 573
rect 110 549 116 550
rect 160 549 162 573
rect 408 549 410 573
rect 672 549 674 573
rect 936 549 938 573
rect 1192 549 1194 573
rect 1448 549 1450 573
rect 1712 549 1714 573
rect 1936 550 1938 573
rect 1976 558 1978 581
rect 1974 557 1980 558
rect 2336 557 2338 581
rect 2528 557 2530 581
rect 2712 557 2714 581
rect 2888 557 2890 581
rect 3064 557 3066 581
rect 3232 557 3234 581
rect 3408 557 3410 581
rect 3584 557 3586 581
rect 3800 558 3802 581
rect 3840 579 3842 622
rect 3888 579 3890 623
rect 4024 579 4026 623
rect 4160 579 4162 623
rect 4296 579 4298 623
rect 4432 579 4434 623
rect 4568 579 4570 623
rect 4704 579 4706 623
rect 4840 579 4842 623
rect 4976 579 4978 623
rect 5112 579 5114 623
rect 5662 622 5668 623
rect 5664 579 5666 622
rect 3839 578 3843 579
rect 3839 573 3843 574
rect 3887 578 3891 579
rect 3887 573 3891 574
rect 4023 578 4027 579
rect 4023 573 4027 574
rect 4047 578 4051 579
rect 4047 573 4051 574
rect 4159 578 4163 579
rect 4159 573 4163 574
rect 4207 578 4211 579
rect 4207 573 4211 574
rect 4295 578 4299 579
rect 4295 573 4299 574
rect 4367 578 4371 579
rect 4367 573 4371 574
rect 4431 578 4435 579
rect 4431 573 4435 574
rect 4527 578 4531 579
rect 4527 573 4531 574
rect 4567 578 4571 579
rect 4567 573 4571 574
rect 4687 578 4691 579
rect 4687 573 4691 574
rect 4703 578 4707 579
rect 4703 573 4707 574
rect 4839 578 4843 579
rect 4839 573 4843 574
rect 4975 578 4979 579
rect 4975 573 4979 574
rect 5111 578 5115 579
rect 5111 573 5115 574
rect 5663 578 5667 579
rect 5663 573 5667 574
rect 3798 557 3804 558
rect 1974 553 1975 557
rect 1979 553 1980 557
rect 1974 552 1980 553
rect 2334 556 2340 557
rect 2334 552 2335 556
rect 2339 552 2340 556
rect 2334 551 2340 552
rect 2526 556 2532 557
rect 2526 552 2527 556
rect 2531 552 2532 556
rect 2526 551 2532 552
rect 2710 556 2716 557
rect 2710 552 2711 556
rect 2715 552 2716 556
rect 2710 551 2716 552
rect 2886 556 2892 557
rect 2886 552 2887 556
rect 2891 552 2892 556
rect 2886 551 2892 552
rect 3062 556 3068 557
rect 3062 552 3063 556
rect 3067 552 3068 556
rect 3062 551 3068 552
rect 3230 556 3236 557
rect 3230 552 3231 556
rect 3235 552 3236 556
rect 3230 551 3236 552
rect 3406 556 3412 557
rect 3406 552 3407 556
rect 3411 552 3412 556
rect 3406 551 3412 552
rect 3582 556 3588 557
rect 3582 552 3583 556
rect 3587 552 3588 556
rect 3798 553 3799 557
rect 3803 553 3804 557
rect 3798 552 3804 553
rect 3582 551 3588 552
rect 3840 550 3842 573
rect 1934 549 1940 550
rect 110 545 111 549
rect 115 545 116 549
rect 110 544 116 545
rect 158 548 164 549
rect 158 544 159 548
rect 163 544 164 548
rect 158 543 164 544
rect 406 548 412 549
rect 406 544 407 548
rect 411 544 412 548
rect 406 543 412 544
rect 670 548 676 549
rect 670 544 671 548
rect 675 544 676 548
rect 670 543 676 544
rect 934 548 940 549
rect 934 544 935 548
rect 939 544 940 548
rect 934 543 940 544
rect 1190 548 1196 549
rect 1190 544 1191 548
rect 1195 544 1196 548
rect 1190 543 1196 544
rect 1446 548 1452 549
rect 1446 544 1447 548
rect 1451 544 1452 548
rect 1446 543 1452 544
rect 1710 548 1716 549
rect 1710 544 1711 548
rect 1715 544 1716 548
rect 1934 545 1935 549
rect 1939 545 1940 549
rect 1934 544 1940 545
rect 3838 549 3844 550
rect 4048 549 4050 573
rect 4208 549 4210 573
rect 4368 549 4370 573
rect 4528 549 4530 573
rect 4688 549 4690 573
rect 5664 550 5666 573
rect 5662 549 5668 550
rect 3838 545 3839 549
rect 3843 545 3844 549
rect 3838 544 3844 545
rect 4046 548 4052 549
rect 4046 544 4047 548
rect 4051 544 4052 548
rect 1710 543 1716 544
rect 4046 543 4052 544
rect 4206 548 4212 549
rect 4206 544 4207 548
rect 4211 544 4212 548
rect 4206 543 4212 544
rect 4366 548 4372 549
rect 4366 544 4367 548
rect 4371 544 4372 548
rect 4366 543 4372 544
rect 4526 548 4532 549
rect 4526 544 4527 548
rect 4531 544 4532 548
rect 4526 543 4532 544
rect 4686 548 4692 549
rect 4686 544 4687 548
rect 4691 544 4692 548
rect 5662 545 5663 549
rect 5667 545 5668 549
rect 5662 544 5668 545
rect 4686 543 4692 544
rect 2306 541 2312 542
rect 1974 540 1980 541
rect 1974 536 1975 540
rect 1979 536 1980 540
rect 2306 537 2307 541
rect 2311 537 2312 541
rect 2306 536 2312 537
rect 2498 541 2504 542
rect 2498 537 2499 541
rect 2503 537 2504 541
rect 2498 536 2504 537
rect 2682 541 2688 542
rect 2682 537 2683 541
rect 2687 537 2688 541
rect 2682 536 2688 537
rect 2858 541 2864 542
rect 2858 537 2859 541
rect 2863 537 2864 541
rect 2858 536 2864 537
rect 3034 541 3040 542
rect 3034 537 3035 541
rect 3039 537 3040 541
rect 3034 536 3040 537
rect 3202 541 3208 542
rect 3202 537 3203 541
rect 3207 537 3208 541
rect 3202 536 3208 537
rect 3378 541 3384 542
rect 3378 537 3379 541
rect 3383 537 3384 541
rect 3378 536 3384 537
rect 3554 541 3560 542
rect 3554 537 3555 541
rect 3559 537 3560 541
rect 3554 536 3560 537
rect 3798 540 3804 541
rect 3798 536 3799 540
rect 3803 536 3804 540
rect 1974 535 1980 536
rect 130 533 136 534
rect 110 532 116 533
rect 110 528 111 532
rect 115 528 116 532
rect 130 529 131 533
rect 135 529 136 533
rect 130 528 136 529
rect 378 533 384 534
rect 378 529 379 533
rect 383 529 384 533
rect 378 528 384 529
rect 642 533 648 534
rect 642 529 643 533
rect 647 529 648 533
rect 642 528 648 529
rect 906 533 912 534
rect 906 529 907 533
rect 911 529 912 533
rect 906 528 912 529
rect 1162 533 1168 534
rect 1162 529 1163 533
rect 1167 529 1168 533
rect 1162 528 1168 529
rect 1418 533 1424 534
rect 1418 529 1419 533
rect 1423 529 1424 533
rect 1418 528 1424 529
rect 1682 533 1688 534
rect 1682 529 1683 533
rect 1687 529 1688 533
rect 1682 528 1688 529
rect 1934 532 1940 533
rect 1934 528 1935 532
rect 1939 528 1940 532
rect 110 527 116 528
rect 112 467 114 527
rect 132 467 134 528
rect 380 467 382 528
rect 644 467 646 528
rect 908 467 910 528
rect 1164 467 1166 528
rect 1420 467 1422 528
rect 1684 467 1686 528
rect 1934 527 1940 528
rect 1936 467 1938 527
rect 1976 475 1978 535
rect 2308 475 2310 536
rect 2500 475 2502 536
rect 2684 475 2686 536
rect 2860 475 2862 536
rect 3036 475 3038 536
rect 3204 475 3206 536
rect 3380 475 3382 536
rect 3556 475 3558 536
rect 3798 535 3804 536
rect 3800 475 3802 535
rect 4018 533 4024 534
rect 3838 532 3844 533
rect 3838 528 3839 532
rect 3843 528 3844 532
rect 4018 529 4019 533
rect 4023 529 4024 533
rect 4018 528 4024 529
rect 4178 533 4184 534
rect 4178 529 4179 533
rect 4183 529 4184 533
rect 4178 528 4184 529
rect 4338 533 4344 534
rect 4338 529 4339 533
rect 4343 529 4344 533
rect 4338 528 4344 529
rect 4498 533 4504 534
rect 4498 529 4499 533
rect 4503 529 4504 533
rect 4498 528 4504 529
rect 4658 533 4664 534
rect 4658 529 4659 533
rect 4663 529 4664 533
rect 4658 528 4664 529
rect 5662 532 5668 533
rect 5662 528 5663 532
rect 5667 528 5668 532
rect 3838 527 3844 528
rect 1975 474 1979 475
rect 1975 469 1979 470
rect 2171 474 2175 475
rect 2171 469 2175 470
rect 2307 474 2311 475
rect 2307 469 2311 470
rect 2315 474 2319 475
rect 2315 469 2319 470
rect 2459 474 2463 475
rect 2459 469 2463 470
rect 2499 474 2503 475
rect 2499 469 2503 470
rect 2603 474 2607 475
rect 2603 469 2607 470
rect 2683 474 2687 475
rect 2683 469 2687 470
rect 2747 474 2751 475
rect 2747 469 2751 470
rect 2859 474 2863 475
rect 2859 469 2863 470
rect 2891 474 2895 475
rect 2891 469 2895 470
rect 3035 474 3039 475
rect 3035 469 3039 470
rect 3203 474 3207 475
rect 3203 469 3207 470
rect 3379 474 3383 475
rect 3379 469 3383 470
rect 3555 474 3559 475
rect 3555 469 3559 470
rect 3799 474 3803 475
rect 3799 469 3803 470
rect 111 466 115 467
rect 111 461 115 462
rect 131 466 135 467
rect 131 461 135 462
rect 195 466 199 467
rect 195 461 199 462
rect 379 466 383 467
rect 379 461 383 462
rect 427 466 431 467
rect 427 461 431 462
rect 643 466 647 467
rect 643 461 647 462
rect 659 466 663 467
rect 659 461 663 462
rect 883 466 887 467
rect 883 461 887 462
rect 907 466 911 467
rect 907 461 911 462
rect 1099 466 1103 467
rect 1099 461 1103 462
rect 1163 466 1167 467
rect 1163 461 1167 462
rect 1323 466 1327 467
rect 1323 461 1327 462
rect 1419 466 1423 467
rect 1419 461 1423 462
rect 1547 466 1551 467
rect 1547 461 1551 462
rect 1683 466 1687 467
rect 1683 461 1687 462
rect 1935 466 1939 467
rect 1935 461 1939 462
rect 112 401 114 461
rect 110 400 116 401
rect 196 400 198 461
rect 428 400 430 461
rect 660 400 662 461
rect 884 400 886 461
rect 1100 400 1102 461
rect 1324 400 1326 461
rect 1548 400 1550 461
rect 1936 401 1938 461
rect 1976 409 1978 469
rect 1974 408 1980 409
rect 2172 408 2174 469
rect 2316 408 2318 469
rect 2460 408 2462 469
rect 2604 408 2606 469
rect 2748 408 2750 469
rect 2892 408 2894 469
rect 3036 408 3038 469
rect 3800 409 3802 469
rect 3840 459 3842 527
rect 4020 459 4022 528
rect 4180 459 4182 528
rect 4340 459 4342 528
rect 4500 459 4502 528
rect 4660 459 4662 528
rect 5662 527 5668 528
rect 5664 459 5666 527
rect 3839 458 3843 459
rect 3839 453 3843 454
rect 3931 458 3935 459
rect 3931 453 3935 454
rect 4019 458 4023 459
rect 4019 453 4023 454
rect 4131 458 4135 459
rect 4131 453 4135 454
rect 4179 458 4183 459
rect 4179 453 4183 454
rect 4331 458 4335 459
rect 4331 453 4335 454
rect 4339 458 4343 459
rect 4339 453 4343 454
rect 4499 458 4503 459
rect 4499 453 4503 454
rect 4523 458 4527 459
rect 4523 453 4527 454
rect 4659 458 4663 459
rect 4659 453 4663 454
rect 4723 458 4727 459
rect 4723 453 4727 454
rect 4923 458 4927 459
rect 4923 453 4927 454
rect 5663 458 5667 459
rect 5663 453 5667 454
rect 3798 408 3804 409
rect 1974 404 1975 408
rect 1979 404 1980 408
rect 1974 403 1980 404
rect 2170 407 2176 408
rect 2170 403 2171 407
rect 2175 403 2176 407
rect 2170 402 2176 403
rect 2314 407 2320 408
rect 2314 403 2315 407
rect 2319 403 2320 407
rect 2314 402 2320 403
rect 2458 407 2464 408
rect 2458 403 2459 407
rect 2463 403 2464 407
rect 2458 402 2464 403
rect 2602 407 2608 408
rect 2602 403 2603 407
rect 2607 403 2608 407
rect 2602 402 2608 403
rect 2746 407 2752 408
rect 2746 403 2747 407
rect 2751 403 2752 407
rect 2746 402 2752 403
rect 2890 407 2896 408
rect 2890 403 2891 407
rect 2895 403 2896 407
rect 2890 402 2896 403
rect 3034 407 3040 408
rect 3034 403 3035 407
rect 3039 403 3040 407
rect 3798 404 3799 408
rect 3803 404 3804 408
rect 3798 403 3804 404
rect 3034 402 3040 403
rect 1934 400 1940 401
rect 110 396 111 400
rect 115 396 116 400
rect 110 395 116 396
rect 194 399 200 400
rect 194 395 195 399
rect 199 395 200 399
rect 194 394 200 395
rect 426 399 432 400
rect 426 395 427 399
rect 431 395 432 399
rect 426 394 432 395
rect 658 399 664 400
rect 658 395 659 399
rect 663 395 664 399
rect 658 394 664 395
rect 882 399 888 400
rect 882 395 883 399
rect 887 395 888 399
rect 882 394 888 395
rect 1098 399 1104 400
rect 1098 395 1099 399
rect 1103 395 1104 399
rect 1098 394 1104 395
rect 1322 399 1328 400
rect 1322 395 1323 399
rect 1327 395 1328 399
rect 1322 394 1328 395
rect 1546 399 1552 400
rect 1546 395 1547 399
rect 1551 395 1552 399
rect 1934 396 1935 400
rect 1939 396 1940 400
rect 1934 395 1940 396
rect 1546 394 1552 395
rect 3840 393 3842 453
rect 2198 392 2204 393
rect 1974 391 1980 392
rect 1974 387 1975 391
rect 1979 387 1980 391
rect 2198 388 2199 392
rect 2203 388 2204 392
rect 2198 387 2204 388
rect 2342 392 2348 393
rect 2342 388 2343 392
rect 2347 388 2348 392
rect 2342 387 2348 388
rect 2486 392 2492 393
rect 2486 388 2487 392
rect 2491 388 2492 392
rect 2486 387 2492 388
rect 2630 392 2636 393
rect 2630 388 2631 392
rect 2635 388 2636 392
rect 2630 387 2636 388
rect 2774 392 2780 393
rect 2774 388 2775 392
rect 2779 388 2780 392
rect 2774 387 2780 388
rect 2918 392 2924 393
rect 2918 388 2919 392
rect 2923 388 2924 392
rect 2918 387 2924 388
rect 3062 392 3068 393
rect 3838 392 3844 393
rect 3932 392 3934 453
rect 4132 392 4134 453
rect 4332 392 4334 453
rect 4524 392 4526 453
rect 4724 392 4726 453
rect 4924 392 4926 453
rect 5664 393 5666 453
rect 5662 392 5668 393
rect 3062 388 3063 392
rect 3067 388 3068 392
rect 3062 387 3068 388
rect 3798 391 3804 392
rect 3798 387 3799 391
rect 3803 387 3804 391
rect 3838 388 3839 392
rect 3843 388 3844 392
rect 3838 387 3844 388
rect 3930 391 3936 392
rect 3930 387 3931 391
rect 3935 387 3936 391
rect 1974 386 1980 387
rect 222 384 228 385
rect 110 383 116 384
rect 110 379 111 383
rect 115 379 116 383
rect 222 380 223 384
rect 227 380 228 384
rect 222 379 228 380
rect 454 384 460 385
rect 454 380 455 384
rect 459 380 460 384
rect 454 379 460 380
rect 686 384 692 385
rect 686 380 687 384
rect 691 380 692 384
rect 686 379 692 380
rect 910 384 916 385
rect 910 380 911 384
rect 915 380 916 384
rect 910 379 916 380
rect 1126 384 1132 385
rect 1126 380 1127 384
rect 1131 380 1132 384
rect 1126 379 1132 380
rect 1350 384 1356 385
rect 1350 380 1351 384
rect 1355 380 1356 384
rect 1350 379 1356 380
rect 1574 384 1580 385
rect 1574 380 1575 384
rect 1579 380 1580 384
rect 1574 379 1580 380
rect 1934 383 1940 384
rect 1934 379 1935 383
rect 1939 379 1940 383
rect 110 378 116 379
rect 112 347 114 378
rect 224 347 226 379
rect 456 347 458 379
rect 688 347 690 379
rect 912 347 914 379
rect 1128 347 1130 379
rect 1352 347 1354 379
rect 1576 347 1578 379
rect 1934 378 1940 379
rect 1936 347 1938 378
rect 1976 359 1978 386
rect 2200 359 2202 387
rect 2344 359 2346 387
rect 2488 359 2490 387
rect 2632 359 2634 387
rect 2776 359 2778 387
rect 2920 359 2922 387
rect 3064 359 3066 387
rect 3798 386 3804 387
rect 3930 386 3936 387
rect 4130 391 4136 392
rect 4130 387 4131 391
rect 4135 387 4136 391
rect 4130 386 4136 387
rect 4330 391 4336 392
rect 4330 387 4331 391
rect 4335 387 4336 391
rect 4330 386 4336 387
rect 4522 391 4528 392
rect 4522 387 4523 391
rect 4527 387 4528 391
rect 4522 386 4528 387
rect 4722 391 4728 392
rect 4722 387 4723 391
rect 4727 387 4728 391
rect 4722 386 4728 387
rect 4922 391 4928 392
rect 4922 387 4923 391
rect 4927 387 4928 391
rect 5662 388 5663 392
rect 5667 388 5668 392
rect 5662 387 5668 388
rect 4922 386 4928 387
rect 3800 359 3802 386
rect 3958 376 3964 377
rect 3838 375 3844 376
rect 3838 371 3839 375
rect 3843 371 3844 375
rect 3958 372 3959 376
rect 3963 372 3964 376
rect 3958 371 3964 372
rect 4158 376 4164 377
rect 4158 372 4159 376
rect 4163 372 4164 376
rect 4158 371 4164 372
rect 4358 376 4364 377
rect 4358 372 4359 376
rect 4363 372 4364 376
rect 4358 371 4364 372
rect 4550 376 4556 377
rect 4550 372 4551 376
rect 4555 372 4556 376
rect 4550 371 4556 372
rect 4750 376 4756 377
rect 4750 372 4751 376
rect 4755 372 4756 376
rect 4750 371 4756 372
rect 4950 376 4956 377
rect 4950 372 4951 376
rect 4955 372 4956 376
rect 4950 371 4956 372
rect 5662 375 5668 376
rect 5662 371 5663 375
rect 5667 371 5668 375
rect 3838 370 3844 371
rect 1975 358 1979 359
rect 1975 353 1979 354
rect 2023 358 2027 359
rect 2023 353 2027 354
rect 2175 358 2179 359
rect 2175 353 2179 354
rect 2199 358 2203 359
rect 2199 353 2203 354
rect 2343 358 2347 359
rect 2343 353 2347 354
rect 2367 358 2371 359
rect 2367 353 2371 354
rect 2487 358 2491 359
rect 2487 353 2491 354
rect 2591 358 2595 359
rect 2591 353 2595 354
rect 2631 358 2635 359
rect 2631 353 2635 354
rect 2775 358 2779 359
rect 2775 353 2779 354
rect 2847 358 2851 359
rect 2847 353 2851 354
rect 2919 358 2923 359
rect 2919 353 2923 354
rect 3063 358 3067 359
rect 3063 353 3067 354
rect 3119 358 3123 359
rect 3119 353 3123 354
rect 3407 358 3411 359
rect 3407 353 3411 354
rect 3679 358 3683 359
rect 3679 353 3683 354
rect 3799 358 3803 359
rect 3799 353 3803 354
rect 111 346 115 347
rect 111 341 115 342
rect 223 346 227 347
rect 223 341 227 342
rect 351 346 355 347
rect 351 341 355 342
rect 455 346 459 347
rect 455 341 459 342
rect 575 346 579 347
rect 575 341 579 342
rect 687 346 691 347
rect 687 341 691 342
rect 799 346 803 347
rect 799 341 803 342
rect 911 346 915 347
rect 911 341 915 342
rect 1015 346 1019 347
rect 1015 341 1019 342
rect 1127 346 1131 347
rect 1127 341 1131 342
rect 1231 346 1235 347
rect 1231 341 1235 342
rect 1351 346 1355 347
rect 1351 341 1355 342
rect 1455 346 1459 347
rect 1455 341 1459 342
rect 1575 346 1579 347
rect 1575 341 1579 342
rect 1935 346 1939 347
rect 1935 341 1939 342
rect 112 318 114 341
rect 110 317 116 318
rect 352 317 354 341
rect 576 317 578 341
rect 800 317 802 341
rect 1016 317 1018 341
rect 1232 317 1234 341
rect 1456 317 1458 341
rect 1936 318 1938 341
rect 1976 330 1978 353
rect 1974 329 1980 330
rect 2024 329 2026 353
rect 2176 329 2178 353
rect 2368 329 2370 353
rect 2592 329 2594 353
rect 2848 329 2850 353
rect 3120 329 3122 353
rect 3408 329 3410 353
rect 3680 329 3682 353
rect 3800 330 3802 353
rect 3840 347 3842 370
rect 3960 347 3962 371
rect 4160 347 4162 371
rect 4360 347 4362 371
rect 4552 347 4554 371
rect 4752 347 4754 371
rect 4952 347 4954 371
rect 5662 370 5668 371
rect 5664 347 5666 370
rect 3839 346 3843 347
rect 3839 341 3843 342
rect 3887 346 3891 347
rect 3887 341 3891 342
rect 3959 346 3963 347
rect 3959 341 3963 342
rect 4135 346 4139 347
rect 4135 341 4139 342
rect 4159 346 4163 347
rect 4159 341 4163 342
rect 4359 346 4363 347
rect 4359 341 4363 342
rect 4383 346 4387 347
rect 4383 341 4387 342
rect 4551 346 4555 347
rect 4551 341 4555 342
rect 4615 346 4619 347
rect 4615 341 4619 342
rect 4751 346 4755 347
rect 4751 341 4755 342
rect 4823 346 4827 347
rect 4823 341 4827 342
rect 4951 346 4955 347
rect 4951 341 4955 342
rect 5015 346 5019 347
rect 5015 341 5019 342
rect 5199 346 5203 347
rect 5199 341 5203 342
rect 5383 346 5387 347
rect 5383 341 5387 342
rect 5543 346 5547 347
rect 5543 341 5547 342
rect 5663 346 5667 347
rect 5663 341 5667 342
rect 3798 329 3804 330
rect 1974 325 1975 329
rect 1979 325 1980 329
rect 1974 324 1980 325
rect 2022 328 2028 329
rect 2022 324 2023 328
rect 2027 324 2028 328
rect 2022 323 2028 324
rect 2174 328 2180 329
rect 2174 324 2175 328
rect 2179 324 2180 328
rect 2174 323 2180 324
rect 2366 328 2372 329
rect 2366 324 2367 328
rect 2371 324 2372 328
rect 2366 323 2372 324
rect 2590 328 2596 329
rect 2590 324 2591 328
rect 2595 324 2596 328
rect 2590 323 2596 324
rect 2846 328 2852 329
rect 2846 324 2847 328
rect 2851 324 2852 328
rect 2846 323 2852 324
rect 3118 328 3124 329
rect 3118 324 3119 328
rect 3123 324 3124 328
rect 3118 323 3124 324
rect 3406 328 3412 329
rect 3406 324 3407 328
rect 3411 324 3412 328
rect 3406 323 3412 324
rect 3678 328 3684 329
rect 3678 324 3679 328
rect 3683 324 3684 328
rect 3798 325 3799 329
rect 3803 325 3804 329
rect 3798 324 3804 325
rect 3678 323 3684 324
rect 3840 318 3842 341
rect 1934 317 1940 318
rect 110 313 111 317
rect 115 313 116 317
rect 110 312 116 313
rect 350 316 356 317
rect 350 312 351 316
rect 355 312 356 316
rect 350 311 356 312
rect 574 316 580 317
rect 574 312 575 316
rect 579 312 580 316
rect 574 311 580 312
rect 798 316 804 317
rect 798 312 799 316
rect 803 312 804 316
rect 798 311 804 312
rect 1014 316 1020 317
rect 1014 312 1015 316
rect 1019 312 1020 316
rect 1014 311 1020 312
rect 1230 316 1236 317
rect 1230 312 1231 316
rect 1235 312 1236 316
rect 1230 311 1236 312
rect 1454 316 1460 317
rect 1454 312 1455 316
rect 1459 312 1460 316
rect 1934 313 1935 317
rect 1939 313 1940 317
rect 3838 317 3844 318
rect 3888 317 3890 341
rect 4136 317 4138 341
rect 4384 317 4386 341
rect 4616 317 4618 341
rect 4824 317 4826 341
rect 5016 317 5018 341
rect 5200 317 5202 341
rect 5384 317 5386 341
rect 5544 317 5546 341
rect 5664 318 5666 341
rect 5662 317 5668 318
rect 1994 313 2000 314
rect 1934 312 1940 313
rect 1974 312 1980 313
rect 1454 311 1460 312
rect 1974 308 1975 312
rect 1979 308 1980 312
rect 1994 309 1995 313
rect 1999 309 2000 313
rect 1994 308 2000 309
rect 2146 313 2152 314
rect 2146 309 2147 313
rect 2151 309 2152 313
rect 2146 308 2152 309
rect 2338 313 2344 314
rect 2338 309 2339 313
rect 2343 309 2344 313
rect 2338 308 2344 309
rect 2562 313 2568 314
rect 2562 309 2563 313
rect 2567 309 2568 313
rect 2562 308 2568 309
rect 2818 313 2824 314
rect 2818 309 2819 313
rect 2823 309 2824 313
rect 2818 308 2824 309
rect 3090 313 3096 314
rect 3090 309 3091 313
rect 3095 309 3096 313
rect 3090 308 3096 309
rect 3378 313 3384 314
rect 3378 309 3379 313
rect 3383 309 3384 313
rect 3378 308 3384 309
rect 3650 313 3656 314
rect 3838 313 3839 317
rect 3843 313 3844 317
rect 3650 309 3651 313
rect 3655 309 3656 313
rect 3650 308 3656 309
rect 3798 312 3804 313
rect 3838 312 3844 313
rect 3886 316 3892 317
rect 3886 312 3887 316
rect 3891 312 3892 316
rect 3798 308 3799 312
rect 3803 308 3804 312
rect 3886 311 3892 312
rect 4134 316 4140 317
rect 4134 312 4135 316
rect 4139 312 4140 316
rect 4134 311 4140 312
rect 4382 316 4388 317
rect 4382 312 4383 316
rect 4387 312 4388 316
rect 4382 311 4388 312
rect 4614 316 4620 317
rect 4614 312 4615 316
rect 4619 312 4620 316
rect 4614 311 4620 312
rect 4822 316 4828 317
rect 4822 312 4823 316
rect 4827 312 4828 316
rect 4822 311 4828 312
rect 5014 316 5020 317
rect 5014 312 5015 316
rect 5019 312 5020 316
rect 5014 311 5020 312
rect 5198 316 5204 317
rect 5198 312 5199 316
rect 5203 312 5204 316
rect 5198 311 5204 312
rect 5382 316 5388 317
rect 5382 312 5383 316
rect 5387 312 5388 316
rect 5382 311 5388 312
rect 5542 316 5548 317
rect 5542 312 5543 316
rect 5547 312 5548 316
rect 5662 313 5663 317
rect 5667 313 5668 317
rect 5662 312 5668 313
rect 5542 311 5548 312
rect 1974 307 1980 308
rect 322 301 328 302
rect 110 300 116 301
rect 110 296 111 300
rect 115 296 116 300
rect 322 297 323 301
rect 327 297 328 301
rect 322 296 328 297
rect 546 301 552 302
rect 546 297 547 301
rect 551 297 552 301
rect 546 296 552 297
rect 770 301 776 302
rect 770 297 771 301
rect 775 297 776 301
rect 770 296 776 297
rect 986 301 992 302
rect 986 297 987 301
rect 991 297 992 301
rect 986 296 992 297
rect 1202 301 1208 302
rect 1202 297 1203 301
rect 1207 297 1208 301
rect 1202 296 1208 297
rect 1426 301 1432 302
rect 1426 297 1427 301
rect 1431 297 1432 301
rect 1426 296 1432 297
rect 1934 300 1940 301
rect 1934 296 1935 300
rect 1939 296 1940 300
rect 110 295 116 296
rect 112 199 114 295
rect 324 199 326 296
rect 548 199 550 296
rect 772 199 774 296
rect 988 199 990 296
rect 1204 199 1206 296
rect 1428 199 1430 296
rect 1934 295 1940 296
rect 1936 199 1938 295
rect 1976 219 1978 307
rect 1996 219 1998 308
rect 2148 219 2150 308
rect 2340 219 2342 308
rect 2564 219 2566 308
rect 2820 219 2822 308
rect 3092 219 3094 308
rect 3380 219 3382 308
rect 3652 219 3654 308
rect 3798 307 3804 308
rect 3800 219 3802 307
rect 3858 301 3864 302
rect 3838 300 3844 301
rect 3838 296 3839 300
rect 3843 296 3844 300
rect 3858 297 3859 301
rect 3863 297 3864 301
rect 3858 296 3864 297
rect 4106 301 4112 302
rect 4106 297 4107 301
rect 4111 297 4112 301
rect 4106 296 4112 297
rect 4354 301 4360 302
rect 4354 297 4355 301
rect 4359 297 4360 301
rect 4354 296 4360 297
rect 4586 301 4592 302
rect 4586 297 4587 301
rect 4591 297 4592 301
rect 4586 296 4592 297
rect 4794 301 4800 302
rect 4794 297 4795 301
rect 4799 297 4800 301
rect 4794 296 4800 297
rect 4986 301 4992 302
rect 4986 297 4987 301
rect 4991 297 4992 301
rect 4986 296 4992 297
rect 5170 301 5176 302
rect 5170 297 5171 301
rect 5175 297 5176 301
rect 5170 296 5176 297
rect 5354 301 5360 302
rect 5354 297 5355 301
rect 5359 297 5360 301
rect 5354 296 5360 297
rect 5514 301 5520 302
rect 5514 297 5515 301
rect 5519 297 5520 301
rect 5514 296 5520 297
rect 5662 300 5668 301
rect 5662 296 5663 300
rect 5667 296 5668 300
rect 3838 295 3844 296
rect 3840 223 3842 295
rect 3860 223 3862 296
rect 4108 223 4110 296
rect 4356 223 4358 296
rect 4588 223 4590 296
rect 4796 223 4798 296
rect 4988 223 4990 296
rect 5172 223 5174 296
rect 5356 223 5358 296
rect 5516 223 5518 296
rect 5662 295 5668 296
rect 5664 223 5666 295
rect 3839 222 3843 223
rect 1975 218 1979 219
rect 1975 213 1979 214
rect 1995 218 1999 219
rect 1995 213 1999 214
rect 2147 218 2151 219
rect 2147 213 2151 214
rect 2171 218 2175 219
rect 2171 213 2175 214
rect 2339 218 2343 219
rect 2339 213 2343 214
rect 2363 218 2367 219
rect 2363 213 2367 214
rect 2547 218 2551 219
rect 2547 213 2551 214
rect 2563 218 2567 219
rect 2563 213 2567 214
rect 2723 218 2727 219
rect 2723 213 2727 214
rect 2819 218 2823 219
rect 2819 213 2823 214
rect 2891 218 2895 219
rect 2891 213 2895 214
rect 3051 218 3055 219
rect 3051 213 3055 214
rect 3091 218 3095 219
rect 3091 213 3095 214
rect 3203 218 3207 219
rect 3203 213 3207 214
rect 3355 218 3359 219
rect 3355 213 3359 214
rect 3379 218 3383 219
rect 3379 213 3383 214
rect 3515 218 3519 219
rect 3515 213 3519 214
rect 3651 218 3655 219
rect 3651 213 3655 214
rect 3799 218 3803 219
rect 3839 217 3843 218
rect 3859 222 3863 223
rect 3859 217 3863 218
rect 4107 222 4111 223
rect 4107 217 4111 218
rect 4291 222 4295 223
rect 4291 217 4295 218
rect 4355 222 4359 223
rect 4355 217 4359 218
rect 4427 222 4431 223
rect 4427 217 4431 218
rect 4563 222 4567 223
rect 4563 217 4567 218
rect 4587 222 4591 223
rect 4587 217 4591 218
rect 4699 222 4703 223
rect 4699 217 4703 218
rect 4795 222 4799 223
rect 4795 217 4799 218
rect 4835 222 4839 223
rect 4835 217 4839 218
rect 4971 222 4975 223
rect 4971 217 4975 218
rect 4987 222 4991 223
rect 4987 217 4991 218
rect 5107 222 5111 223
rect 5107 217 5111 218
rect 5171 222 5175 223
rect 5171 217 5175 218
rect 5243 222 5247 223
rect 5243 217 5247 218
rect 5355 222 5359 223
rect 5355 217 5359 218
rect 5379 222 5383 223
rect 5379 217 5383 218
rect 5515 222 5519 223
rect 5515 217 5519 218
rect 5663 222 5667 223
rect 5663 217 5667 218
rect 3799 213 3803 214
rect 111 198 115 199
rect 111 193 115 194
rect 131 198 135 199
rect 131 193 135 194
rect 267 198 271 199
rect 267 193 271 194
rect 323 198 327 199
rect 323 193 327 194
rect 403 198 407 199
rect 403 193 407 194
rect 539 198 543 199
rect 539 193 543 194
rect 547 198 551 199
rect 547 193 551 194
rect 675 198 679 199
rect 675 193 679 194
rect 771 198 775 199
rect 771 193 775 194
rect 811 198 815 199
rect 811 193 815 194
rect 947 198 951 199
rect 947 193 951 194
rect 987 198 991 199
rect 987 193 991 194
rect 1083 198 1087 199
rect 1083 193 1087 194
rect 1203 198 1207 199
rect 1203 193 1207 194
rect 1227 198 1231 199
rect 1227 193 1231 194
rect 1371 198 1375 199
rect 1371 193 1375 194
rect 1427 198 1431 199
rect 1427 193 1431 194
rect 1515 198 1519 199
rect 1515 193 1519 194
rect 1651 198 1655 199
rect 1651 193 1655 194
rect 1787 198 1791 199
rect 1787 193 1791 194
rect 1935 198 1939 199
rect 1935 193 1939 194
rect 112 133 114 193
rect 110 132 116 133
rect 132 132 134 193
rect 268 132 270 193
rect 404 132 406 193
rect 540 132 542 193
rect 676 132 678 193
rect 812 132 814 193
rect 948 132 950 193
rect 1084 132 1086 193
rect 1228 132 1230 193
rect 1372 132 1374 193
rect 1516 132 1518 193
rect 1652 132 1654 193
rect 1788 132 1790 193
rect 1936 133 1938 193
rect 1976 153 1978 213
rect 1974 152 1980 153
rect 1996 152 1998 213
rect 2172 152 2174 213
rect 2364 152 2366 213
rect 2548 152 2550 213
rect 2724 152 2726 213
rect 2892 152 2894 213
rect 3052 152 3054 213
rect 3204 152 3206 213
rect 3356 152 3358 213
rect 3516 152 3518 213
rect 3652 152 3654 213
rect 3800 153 3802 213
rect 3840 157 3842 217
rect 3838 156 3844 157
rect 4292 156 4294 217
rect 4428 156 4430 217
rect 4564 156 4566 217
rect 4700 156 4702 217
rect 4836 156 4838 217
rect 4972 156 4974 217
rect 5108 156 5110 217
rect 5244 156 5246 217
rect 5380 156 5382 217
rect 5516 156 5518 217
rect 5664 157 5666 217
rect 5662 156 5668 157
rect 3798 152 3804 153
rect 1974 148 1975 152
rect 1979 148 1980 152
rect 1974 147 1980 148
rect 1994 151 2000 152
rect 1994 147 1995 151
rect 1999 147 2000 151
rect 1994 146 2000 147
rect 2170 151 2176 152
rect 2170 147 2171 151
rect 2175 147 2176 151
rect 2170 146 2176 147
rect 2362 151 2368 152
rect 2362 147 2363 151
rect 2367 147 2368 151
rect 2362 146 2368 147
rect 2546 151 2552 152
rect 2546 147 2547 151
rect 2551 147 2552 151
rect 2546 146 2552 147
rect 2722 151 2728 152
rect 2722 147 2723 151
rect 2727 147 2728 151
rect 2722 146 2728 147
rect 2890 151 2896 152
rect 2890 147 2891 151
rect 2895 147 2896 151
rect 2890 146 2896 147
rect 3050 151 3056 152
rect 3050 147 3051 151
rect 3055 147 3056 151
rect 3050 146 3056 147
rect 3202 151 3208 152
rect 3202 147 3203 151
rect 3207 147 3208 151
rect 3202 146 3208 147
rect 3354 151 3360 152
rect 3354 147 3355 151
rect 3359 147 3360 151
rect 3354 146 3360 147
rect 3514 151 3520 152
rect 3514 147 3515 151
rect 3519 147 3520 151
rect 3514 146 3520 147
rect 3650 151 3656 152
rect 3650 147 3651 151
rect 3655 147 3656 151
rect 3798 148 3799 152
rect 3803 148 3804 152
rect 3838 152 3839 156
rect 3843 152 3844 156
rect 3838 151 3844 152
rect 4290 155 4296 156
rect 4290 151 4291 155
rect 4295 151 4296 155
rect 4290 150 4296 151
rect 4426 155 4432 156
rect 4426 151 4427 155
rect 4431 151 4432 155
rect 4426 150 4432 151
rect 4562 155 4568 156
rect 4562 151 4563 155
rect 4567 151 4568 155
rect 4562 150 4568 151
rect 4698 155 4704 156
rect 4698 151 4699 155
rect 4703 151 4704 155
rect 4698 150 4704 151
rect 4834 155 4840 156
rect 4834 151 4835 155
rect 4839 151 4840 155
rect 4834 150 4840 151
rect 4970 155 4976 156
rect 4970 151 4971 155
rect 4975 151 4976 155
rect 4970 150 4976 151
rect 5106 155 5112 156
rect 5106 151 5107 155
rect 5111 151 5112 155
rect 5106 150 5112 151
rect 5242 155 5248 156
rect 5242 151 5243 155
rect 5247 151 5248 155
rect 5242 150 5248 151
rect 5378 155 5384 156
rect 5378 151 5379 155
rect 5383 151 5384 155
rect 5378 150 5384 151
rect 5514 155 5520 156
rect 5514 151 5515 155
rect 5519 151 5520 155
rect 5662 152 5663 156
rect 5667 152 5668 156
rect 5662 151 5668 152
rect 5514 150 5520 151
rect 3798 147 3804 148
rect 3650 146 3656 147
rect 4318 140 4324 141
rect 3838 139 3844 140
rect 2022 136 2028 137
rect 1974 135 1980 136
rect 1934 132 1940 133
rect 110 128 111 132
rect 115 128 116 132
rect 110 127 116 128
rect 130 131 136 132
rect 130 127 131 131
rect 135 127 136 131
rect 130 126 136 127
rect 266 131 272 132
rect 266 127 267 131
rect 271 127 272 131
rect 266 126 272 127
rect 402 131 408 132
rect 402 127 403 131
rect 407 127 408 131
rect 402 126 408 127
rect 538 131 544 132
rect 538 127 539 131
rect 543 127 544 131
rect 538 126 544 127
rect 674 131 680 132
rect 674 127 675 131
rect 679 127 680 131
rect 674 126 680 127
rect 810 131 816 132
rect 810 127 811 131
rect 815 127 816 131
rect 810 126 816 127
rect 946 131 952 132
rect 946 127 947 131
rect 951 127 952 131
rect 946 126 952 127
rect 1082 131 1088 132
rect 1082 127 1083 131
rect 1087 127 1088 131
rect 1082 126 1088 127
rect 1226 131 1232 132
rect 1226 127 1227 131
rect 1231 127 1232 131
rect 1226 126 1232 127
rect 1370 131 1376 132
rect 1370 127 1371 131
rect 1375 127 1376 131
rect 1370 126 1376 127
rect 1514 131 1520 132
rect 1514 127 1515 131
rect 1519 127 1520 131
rect 1514 126 1520 127
rect 1650 131 1656 132
rect 1650 127 1651 131
rect 1655 127 1656 131
rect 1650 126 1656 127
rect 1786 131 1792 132
rect 1786 127 1787 131
rect 1791 127 1792 131
rect 1934 128 1935 132
rect 1939 128 1940 132
rect 1974 131 1975 135
rect 1979 131 1980 135
rect 2022 132 2023 136
rect 2027 132 2028 136
rect 2022 131 2028 132
rect 2198 136 2204 137
rect 2198 132 2199 136
rect 2203 132 2204 136
rect 2198 131 2204 132
rect 2390 136 2396 137
rect 2390 132 2391 136
rect 2395 132 2396 136
rect 2390 131 2396 132
rect 2574 136 2580 137
rect 2574 132 2575 136
rect 2579 132 2580 136
rect 2574 131 2580 132
rect 2750 136 2756 137
rect 2750 132 2751 136
rect 2755 132 2756 136
rect 2750 131 2756 132
rect 2918 136 2924 137
rect 2918 132 2919 136
rect 2923 132 2924 136
rect 2918 131 2924 132
rect 3078 136 3084 137
rect 3078 132 3079 136
rect 3083 132 3084 136
rect 3078 131 3084 132
rect 3230 136 3236 137
rect 3230 132 3231 136
rect 3235 132 3236 136
rect 3230 131 3236 132
rect 3382 136 3388 137
rect 3382 132 3383 136
rect 3387 132 3388 136
rect 3382 131 3388 132
rect 3542 136 3548 137
rect 3542 132 3543 136
rect 3547 132 3548 136
rect 3542 131 3548 132
rect 3678 136 3684 137
rect 3678 132 3679 136
rect 3683 132 3684 136
rect 3678 131 3684 132
rect 3798 135 3804 136
rect 3798 131 3799 135
rect 3803 131 3804 135
rect 3838 135 3839 139
rect 3843 135 3844 139
rect 4318 136 4319 140
rect 4323 136 4324 140
rect 4318 135 4324 136
rect 4454 140 4460 141
rect 4454 136 4455 140
rect 4459 136 4460 140
rect 4454 135 4460 136
rect 4590 140 4596 141
rect 4590 136 4591 140
rect 4595 136 4596 140
rect 4590 135 4596 136
rect 4726 140 4732 141
rect 4726 136 4727 140
rect 4731 136 4732 140
rect 4726 135 4732 136
rect 4862 140 4868 141
rect 4862 136 4863 140
rect 4867 136 4868 140
rect 4862 135 4868 136
rect 4998 140 5004 141
rect 4998 136 4999 140
rect 5003 136 5004 140
rect 4998 135 5004 136
rect 5134 140 5140 141
rect 5134 136 5135 140
rect 5139 136 5140 140
rect 5134 135 5140 136
rect 5270 140 5276 141
rect 5270 136 5271 140
rect 5275 136 5276 140
rect 5270 135 5276 136
rect 5406 140 5412 141
rect 5406 136 5407 140
rect 5411 136 5412 140
rect 5406 135 5412 136
rect 5542 140 5548 141
rect 5542 136 5543 140
rect 5547 136 5548 140
rect 5542 135 5548 136
rect 5662 139 5668 140
rect 5662 135 5663 139
rect 5667 135 5668 139
rect 3838 134 3844 135
rect 1974 130 1980 131
rect 1934 127 1940 128
rect 1786 126 1792 127
rect 158 116 164 117
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 158 112 159 116
rect 163 112 164 116
rect 158 111 164 112
rect 294 116 300 117
rect 294 112 295 116
rect 299 112 300 116
rect 294 111 300 112
rect 430 116 436 117
rect 430 112 431 116
rect 435 112 436 116
rect 430 111 436 112
rect 566 116 572 117
rect 566 112 567 116
rect 571 112 572 116
rect 566 111 572 112
rect 702 116 708 117
rect 702 112 703 116
rect 707 112 708 116
rect 702 111 708 112
rect 838 116 844 117
rect 838 112 839 116
rect 843 112 844 116
rect 838 111 844 112
rect 974 116 980 117
rect 974 112 975 116
rect 979 112 980 116
rect 974 111 980 112
rect 1110 116 1116 117
rect 1110 112 1111 116
rect 1115 112 1116 116
rect 1110 111 1116 112
rect 1254 116 1260 117
rect 1254 112 1255 116
rect 1259 112 1260 116
rect 1254 111 1260 112
rect 1398 116 1404 117
rect 1398 112 1399 116
rect 1403 112 1404 116
rect 1398 111 1404 112
rect 1542 116 1548 117
rect 1542 112 1543 116
rect 1547 112 1548 116
rect 1542 111 1548 112
rect 1678 116 1684 117
rect 1678 112 1679 116
rect 1683 112 1684 116
rect 1678 111 1684 112
rect 1814 116 1820 117
rect 1814 112 1815 116
rect 1819 112 1820 116
rect 1814 111 1820 112
rect 1934 115 1940 116
rect 1934 111 1935 115
rect 1939 111 1940 115
rect 110 110 116 111
rect 112 87 114 110
rect 160 87 162 111
rect 296 87 298 111
rect 432 87 434 111
rect 568 87 570 111
rect 704 87 706 111
rect 840 87 842 111
rect 976 87 978 111
rect 1112 87 1114 111
rect 1256 87 1258 111
rect 1400 87 1402 111
rect 1544 87 1546 111
rect 1680 87 1682 111
rect 1816 87 1818 111
rect 1934 110 1940 111
rect 1936 87 1938 110
rect 1976 107 1978 130
rect 2024 107 2026 131
rect 2200 107 2202 131
rect 2392 107 2394 131
rect 2576 107 2578 131
rect 2752 107 2754 131
rect 2920 107 2922 131
rect 3080 107 3082 131
rect 3232 107 3234 131
rect 3384 107 3386 131
rect 3544 107 3546 131
rect 3680 107 3682 131
rect 3798 130 3804 131
rect 3800 107 3802 130
rect 3840 111 3842 134
rect 4320 111 4322 135
rect 4456 111 4458 135
rect 4592 111 4594 135
rect 4728 111 4730 135
rect 4864 111 4866 135
rect 5000 111 5002 135
rect 5136 111 5138 135
rect 5272 111 5274 135
rect 5408 111 5410 135
rect 5544 111 5546 135
rect 5662 134 5668 135
rect 5664 111 5666 134
rect 3839 110 3843 111
rect 1975 106 1979 107
rect 1975 101 1979 102
rect 2023 106 2027 107
rect 2023 101 2027 102
rect 2199 106 2203 107
rect 2199 101 2203 102
rect 2391 106 2395 107
rect 2391 101 2395 102
rect 2575 106 2579 107
rect 2575 101 2579 102
rect 2751 106 2755 107
rect 2751 101 2755 102
rect 2919 106 2923 107
rect 2919 101 2923 102
rect 3079 106 3083 107
rect 3079 101 3083 102
rect 3231 106 3235 107
rect 3231 101 3235 102
rect 3383 106 3387 107
rect 3383 101 3387 102
rect 3543 106 3547 107
rect 3543 101 3547 102
rect 3679 106 3683 107
rect 3679 101 3683 102
rect 3799 106 3803 107
rect 3839 105 3843 106
rect 4319 110 4323 111
rect 4319 105 4323 106
rect 4455 110 4459 111
rect 4455 105 4459 106
rect 4591 110 4595 111
rect 4591 105 4595 106
rect 4727 110 4731 111
rect 4727 105 4731 106
rect 4863 110 4867 111
rect 4863 105 4867 106
rect 4999 110 5003 111
rect 4999 105 5003 106
rect 5135 110 5139 111
rect 5135 105 5139 106
rect 5271 110 5275 111
rect 5271 105 5275 106
rect 5407 110 5411 111
rect 5407 105 5411 106
rect 5543 110 5547 111
rect 5543 105 5547 106
rect 5663 110 5667 111
rect 5663 105 5667 106
rect 3799 101 3803 102
rect 111 86 115 87
rect 111 81 115 82
rect 159 86 163 87
rect 159 81 163 82
rect 295 86 299 87
rect 295 81 299 82
rect 431 86 435 87
rect 431 81 435 82
rect 567 86 571 87
rect 567 81 571 82
rect 703 86 707 87
rect 703 81 707 82
rect 839 86 843 87
rect 839 81 843 82
rect 975 86 979 87
rect 975 81 979 82
rect 1111 86 1115 87
rect 1111 81 1115 82
rect 1255 86 1259 87
rect 1255 81 1259 82
rect 1399 86 1403 87
rect 1399 81 1403 82
rect 1543 86 1547 87
rect 1543 81 1547 82
rect 1679 86 1683 87
rect 1679 81 1683 82
rect 1815 86 1819 87
rect 1815 81 1819 82
rect 1935 86 1939 87
rect 1935 81 1939 82
<< m4c >>
rect 111 5730 115 5734
rect 159 5730 163 5734
rect 295 5730 299 5734
rect 431 5730 435 5734
rect 567 5730 571 5734
rect 703 5730 707 5734
rect 839 5730 843 5734
rect 975 5730 979 5734
rect 1935 5730 1939 5734
rect 1975 5670 1979 5674
rect 2103 5670 2107 5674
rect 2239 5670 2243 5674
rect 2375 5670 2379 5674
rect 2511 5670 2515 5674
rect 2647 5670 2651 5674
rect 2783 5670 2787 5674
rect 2919 5670 2923 5674
rect 3055 5670 3059 5674
rect 3191 5670 3195 5674
rect 3327 5670 3331 5674
rect 3463 5670 3467 5674
rect 3599 5670 3603 5674
rect 3799 5670 3803 5674
rect 111 5602 115 5606
rect 131 5602 135 5606
rect 267 5602 271 5606
rect 403 5602 407 5606
rect 539 5602 543 5606
rect 675 5602 679 5606
rect 755 5602 759 5606
rect 811 5602 815 5606
rect 891 5602 895 5606
rect 947 5602 951 5606
rect 1027 5602 1031 5606
rect 1163 5602 1167 5606
rect 1935 5602 1939 5606
rect 3839 5606 3843 5610
rect 4243 5606 4247 5610
rect 4379 5606 4383 5610
rect 4515 5606 4519 5610
rect 4651 5606 4655 5610
rect 4787 5606 4791 5610
rect 4923 5606 4927 5610
rect 5059 5606 5063 5610
rect 5663 5606 5667 5610
rect 1975 5558 1979 5562
rect 1995 5558 1999 5562
rect 2075 5558 2079 5562
rect 2131 5558 2135 5562
rect 2211 5558 2215 5562
rect 2267 5558 2271 5562
rect 2347 5558 2351 5562
rect 2403 5558 2407 5562
rect 2483 5558 2487 5562
rect 2555 5558 2559 5562
rect 2619 5558 2623 5562
rect 2707 5558 2711 5562
rect 2755 5558 2759 5562
rect 2859 5558 2863 5562
rect 2891 5558 2895 5562
rect 3011 5558 3015 5562
rect 3027 5558 3031 5562
rect 3163 5558 3167 5562
rect 3299 5558 3303 5562
rect 3323 5558 3327 5562
rect 3435 5558 3439 5562
rect 3483 5558 3487 5562
rect 3571 5558 3575 5562
rect 3799 5558 3803 5562
rect 3839 5494 3843 5498
rect 4271 5494 4275 5498
rect 4407 5494 4411 5498
rect 4455 5494 4459 5498
rect 4543 5494 4547 5498
rect 4591 5494 4595 5498
rect 4679 5494 4683 5498
rect 4727 5494 4731 5498
rect 4815 5494 4819 5498
rect 4863 5494 4867 5498
rect 4951 5494 4955 5498
rect 5087 5494 5091 5498
rect 5663 5494 5667 5498
rect 111 5478 115 5482
rect 783 5478 787 5482
rect 863 5478 867 5482
rect 919 5478 923 5482
rect 999 5478 1003 5482
rect 1055 5478 1059 5482
rect 1135 5478 1139 5482
rect 1191 5478 1195 5482
rect 1271 5478 1275 5482
rect 1407 5478 1411 5482
rect 1543 5478 1547 5482
rect 1679 5478 1683 5482
rect 1815 5478 1819 5482
rect 1935 5478 1939 5482
rect 1975 5434 1979 5438
rect 2023 5434 2027 5438
rect 2159 5434 2163 5438
rect 2295 5434 2299 5438
rect 2431 5434 2435 5438
rect 2583 5434 2587 5438
rect 2735 5434 2739 5438
rect 2831 5434 2835 5438
rect 2887 5434 2891 5438
rect 2967 5434 2971 5438
rect 3039 5434 3043 5438
rect 3103 5434 3107 5438
rect 3191 5434 3195 5438
rect 3239 5434 3243 5438
rect 3351 5434 3355 5438
rect 3511 5434 3515 5438
rect 3799 5434 3803 5438
rect 111 5366 115 5370
rect 427 5366 431 5370
rect 563 5366 567 5370
rect 699 5366 703 5370
rect 835 5366 839 5370
rect 971 5366 975 5370
rect 1107 5366 1111 5370
rect 1243 5366 1247 5370
rect 1379 5366 1383 5370
rect 1515 5366 1519 5370
rect 1651 5366 1655 5370
rect 1787 5366 1791 5370
rect 1935 5366 1939 5370
rect 3839 5382 3843 5386
rect 4283 5382 4287 5386
rect 4427 5382 4431 5386
rect 4483 5382 4487 5386
rect 4563 5382 4567 5386
rect 4699 5382 4703 5386
rect 4835 5382 4839 5386
rect 4931 5382 4935 5386
rect 5171 5382 5175 5386
rect 5419 5382 5423 5386
rect 5663 5382 5667 5386
rect 1975 5286 1979 5290
rect 1995 5286 1999 5290
rect 2219 5286 2223 5290
rect 2467 5286 2471 5290
rect 2715 5286 2719 5290
rect 2803 5286 2807 5290
rect 2939 5286 2943 5290
rect 2971 5286 2975 5290
rect 3075 5286 3079 5290
rect 3211 5286 3215 5290
rect 3799 5286 3803 5290
rect 111 5254 115 5258
rect 455 5254 459 5258
rect 591 5254 595 5258
rect 727 5254 731 5258
rect 863 5254 867 5258
rect 999 5254 1003 5258
rect 1135 5254 1139 5258
rect 1271 5254 1275 5258
rect 1407 5254 1411 5258
rect 1543 5254 1547 5258
rect 1679 5254 1683 5258
rect 1815 5254 1819 5258
rect 1935 5254 1939 5258
rect 3839 5242 3843 5246
rect 3887 5242 3891 5246
rect 4023 5242 4027 5246
rect 4159 5242 4163 5246
rect 4295 5242 4299 5246
rect 4311 5242 4315 5246
rect 4431 5242 4435 5246
rect 4511 5242 4515 5246
rect 4567 5242 4571 5246
rect 4703 5242 4707 5246
rect 4727 5242 4731 5246
rect 4839 5242 4843 5246
rect 4959 5242 4963 5246
rect 4991 5242 4995 5246
rect 5151 5242 5155 5246
rect 5199 5242 5203 5246
rect 5319 5242 5323 5246
rect 5447 5242 5451 5246
rect 5495 5242 5499 5246
rect 5663 5242 5667 5246
rect 1975 5170 1979 5174
rect 2023 5170 2027 5174
rect 2159 5170 2163 5174
rect 2247 5170 2251 5174
rect 2295 5170 2299 5174
rect 2431 5170 2435 5174
rect 2495 5170 2499 5174
rect 2567 5170 2571 5174
rect 2703 5170 2707 5174
rect 2743 5170 2747 5174
rect 2839 5170 2843 5174
rect 2975 5170 2979 5174
rect 2999 5170 3003 5174
rect 3111 5170 3115 5174
rect 3247 5170 3251 5174
rect 3391 5170 3395 5174
rect 3543 5170 3547 5174
rect 3679 5170 3683 5174
rect 3799 5170 3803 5174
rect 111 5126 115 5130
rect 267 5126 271 5130
rect 403 5126 407 5130
rect 427 5126 431 5130
rect 539 5126 543 5130
rect 563 5126 567 5130
rect 675 5126 679 5130
rect 699 5126 703 5130
rect 811 5126 815 5130
rect 835 5126 839 5130
rect 947 5126 951 5130
rect 971 5126 975 5130
rect 1107 5126 1111 5130
rect 1243 5126 1247 5130
rect 1379 5126 1383 5130
rect 1515 5126 1519 5130
rect 1651 5126 1655 5130
rect 1787 5126 1791 5130
rect 3839 5130 3843 5134
rect 1935 5126 1939 5130
rect 3859 5130 3863 5134
rect 3979 5130 3983 5134
rect 3995 5130 3999 5134
rect 4131 5130 4135 5134
rect 4267 5130 4271 5134
rect 4275 5130 4279 5134
rect 4403 5130 4407 5134
rect 4539 5130 4543 5134
rect 4579 5130 4583 5134
rect 4675 5130 4679 5134
rect 4811 5130 4815 5134
rect 4883 5130 4887 5134
rect 4963 5130 4967 5134
rect 5123 5130 5127 5134
rect 5195 5130 5199 5134
rect 5291 5130 5295 5134
rect 5467 5130 5471 5134
rect 5515 5130 5519 5134
rect 5663 5130 5667 5134
rect 1975 5058 1979 5062
rect 1995 5058 1999 5062
rect 2131 5058 2135 5062
rect 2267 5058 2271 5062
rect 2403 5058 2407 5062
rect 2539 5058 2543 5062
rect 2675 5058 2679 5062
rect 2811 5058 2815 5062
rect 2947 5058 2951 5062
rect 3083 5058 3087 5062
rect 3107 5058 3111 5062
rect 3219 5058 3223 5062
rect 3243 5058 3247 5062
rect 3363 5058 3367 5062
rect 3379 5058 3383 5062
rect 3515 5058 3519 5062
rect 3651 5058 3655 5062
rect 3799 5058 3803 5062
rect 111 5002 115 5006
rect 159 5002 163 5006
rect 295 5002 299 5006
rect 431 5002 435 5006
rect 567 5002 571 5006
rect 703 5002 707 5006
rect 839 5002 843 5006
rect 975 5002 979 5006
rect 1935 5002 1939 5006
rect 3839 5002 3843 5006
rect 4007 5002 4011 5006
rect 4303 5002 4307 5006
rect 4607 5002 4611 5006
rect 4863 5002 4867 5006
rect 4911 5002 4915 5006
rect 4999 5002 5003 5006
rect 5135 5002 5139 5006
rect 5223 5002 5227 5006
rect 5271 5002 5275 5006
rect 5407 5002 5411 5006
rect 5543 5002 5547 5006
rect 5663 5002 5667 5006
rect 1975 4938 1979 4942
rect 3135 4938 3139 4942
rect 3271 4938 3275 4942
rect 3407 4938 3411 4942
rect 3543 4938 3547 4942
rect 3679 4938 3683 4942
rect 3799 4938 3803 4942
rect 111 4882 115 4886
rect 131 4882 135 4886
rect 267 4882 271 4886
rect 403 4882 407 4886
rect 539 4882 543 4886
rect 675 4882 679 4886
rect 1935 4882 1939 4886
rect 3839 4878 3843 4882
rect 4483 4878 4487 4882
rect 4675 4878 4679 4882
rect 4835 4878 4839 4882
rect 4875 4878 4879 4882
rect 4971 4878 4975 4882
rect 5091 4878 5095 4882
rect 5107 4878 5111 4882
rect 5243 4878 5247 4882
rect 5315 4878 5319 4882
rect 5379 4878 5383 4882
rect 5515 4878 5519 4882
rect 5663 4878 5667 4882
rect 1975 4798 1979 4802
rect 3107 4798 3111 4802
rect 3243 4798 3247 4802
rect 3379 4798 3383 4802
rect 3515 4798 3519 4802
rect 3651 4798 3655 4802
rect 3799 4798 3803 4802
rect 111 4766 115 4770
rect 159 4766 163 4770
rect 295 4766 299 4770
rect 431 4766 435 4770
rect 567 4766 571 4770
rect 703 4766 707 4770
rect 1935 4766 1939 4770
rect 3839 4746 3843 4750
rect 4119 4746 4123 4750
rect 4375 4746 4379 4750
rect 4511 4746 4515 4750
rect 4647 4746 4651 4750
rect 4703 4746 4707 4750
rect 4903 4746 4907 4750
rect 4943 4746 4947 4750
rect 5119 4746 5123 4750
rect 5255 4746 5259 4750
rect 5343 4746 5347 4750
rect 5543 4746 5547 4750
rect 5663 4746 5667 4750
rect 111 4646 115 4650
rect 131 4646 135 4650
rect 211 4646 215 4650
rect 267 4646 271 4650
rect 403 4646 407 4650
rect 427 4646 431 4650
rect 539 4646 543 4650
rect 667 4646 671 4650
rect 675 4646 679 4650
rect 931 4646 935 4650
rect 1219 4646 1223 4650
rect 1515 4646 1519 4650
rect 1787 4646 1791 4650
rect 1935 4646 1939 4650
rect 1975 4646 1979 4650
rect 2023 4646 2027 4650
rect 2159 4646 2163 4650
rect 2311 4646 2315 4650
rect 2479 4646 2483 4650
rect 2655 4646 2659 4650
rect 2831 4646 2835 4650
rect 3007 4646 3011 4650
rect 3135 4646 3139 4650
rect 3183 4646 3187 4650
rect 3271 4646 3275 4650
rect 3351 4646 3355 4650
rect 3407 4646 3411 4650
rect 3527 4646 3531 4650
rect 3543 4646 3547 4650
rect 3679 4646 3683 4650
rect 3799 4646 3803 4650
rect 3839 4614 3843 4618
rect 4035 4614 4039 4618
rect 4091 4614 4095 4618
rect 4331 4614 4335 4618
rect 4347 4614 4351 4618
rect 4619 4614 4623 4618
rect 4627 4614 4631 4618
rect 4915 4614 4919 4618
rect 4931 4614 4935 4618
rect 5227 4614 5231 4618
rect 5235 4614 5239 4618
rect 5515 4614 5519 4618
rect 5663 4614 5667 4618
rect 111 4534 115 4538
rect 239 4534 243 4538
rect 447 4534 451 4538
rect 455 4534 459 4538
rect 623 4534 627 4538
rect 695 4534 699 4538
rect 807 4534 811 4538
rect 959 4534 963 4538
rect 999 4534 1003 4538
rect 1199 4534 1203 4538
rect 1247 4534 1251 4538
rect 1407 4534 1411 4538
rect 1543 4534 1547 4538
rect 1623 4534 1627 4538
rect 1815 4534 1819 4538
rect 1935 4534 1939 4538
rect 1975 4534 1979 4538
rect 1995 4534 1999 4538
rect 2131 4534 2135 4538
rect 2227 4534 2231 4538
rect 2283 4534 2287 4538
rect 2451 4534 2455 4538
rect 2459 4534 2463 4538
rect 2627 4534 2631 4538
rect 2691 4534 2695 4538
rect 2803 4534 2807 4538
rect 2915 4534 2919 4538
rect 2979 4534 2983 4538
rect 3131 4534 3135 4538
rect 3155 4534 3159 4538
rect 3323 4534 3327 4538
rect 3355 4534 3359 4538
rect 3499 4534 3503 4538
rect 3579 4534 3583 4538
rect 3651 4534 3655 4538
rect 3799 4534 3803 4538
rect 3839 4486 3843 4490
rect 4063 4486 4067 4490
rect 4311 4486 4315 4490
rect 4359 4486 4363 4490
rect 4535 4486 4539 4490
rect 4655 4486 4659 4490
rect 4775 4486 4779 4490
rect 4959 4486 4963 4490
rect 5023 4486 5027 4490
rect 5263 4486 5267 4490
rect 5279 4486 5283 4490
rect 5543 4486 5547 4490
rect 5663 4486 5667 4490
rect 111 4418 115 4422
rect 419 4418 423 4422
rect 571 4418 575 4422
rect 595 4418 599 4422
rect 739 4418 743 4422
rect 779 4418 783 4422
rect 915 4418 919 4422
rect 971 4418 975 4422
rect 1107 4418 1111 4422
rect 1171 4418 1175 4422
rect 1299 4418 1303 4422
rect 1379 4418 1383 4422
rect 1499 4418 1503 4422
rect 1595 4418 1599 4422
rect 1707 4418 1711 4422
rect 1787 4418 1791 4422
rect 1935 4418 1939 4422
rect 1975 4418 1979 4422
rect 2023 4418 2027 4422
rect 2119 4418 2123 4422
rect 2255 4418 2259 4422
rect 2343 4418 2347 4422
rect 2487 4418 2491 4422
rect 2567 4418 2571 4422
rect 2719 4418 2723 4422
rect 2783 4418 2787 4422
rect 2943 4418 2947 4422
rect 2991 4418 2995 4422
rect 3159 4418 3163 4422
rect 3199 4418 3203 4422
rect 3383 4418 3387 4422
rect 3407 4418 3411 4422
rect 3607 4418 3611 4422
rect 3799 4418 3803 4422
rect 111 4306 115 4310
rect 599 4306 603 4310
rect 655 4306 659 4310
rect 767 4306 771 4310
rect 823 4306 827 4310
rect 943 4306 947 4310
rect 991 4306 995 4310
rect 1135 4306 1139 4310
rect 1167 4306 1171 4310
rect 1327 4306 1331 4310
rect 1343 4306 1347 4310
rect 1519 4306 1523 4310
rect 1527 4306 1531 4310
rect 1703 4306 1707 4310
rect 1735 4306 1739 4310
rect 1935 4306 1939 4310
rect 3839 4354 3843 4358
rect 4283 4354 4287 4358
rect 4507 4354 4511 4358
rect 4515 4354 4519 4358
rect 4691 4354 4695 4358
rect 4747 4354 4751 4358
rect 4875 4354 4879 4358
rect 4995 4354 4999 4358
rect 5067 4354 5071 4358
rect 5251 4354 5255 4358
rect 5267 4354 5271 4358
rect 5467 4354 5471 4358
rect 5515 4354 5519 4358
rect 5663 4354 5667 4358
rect 1975 4298 1979 4302
rect 2019 4298 2023 4302
rect 2091 4298 2095 4302
rect 2243 4298 2247 4302
rect 2315 4298 2319 4302
rect 2459 4298 2463 4302
rect 2539 4298 2543 4302
rect 2667 4298 2671 4302
rect 2755 4298 2759 4302
rect 2875 4298 2879 4302
rect 2963 4298 2967 4302
rect 3083 4298 3087 4302
rect 3171 4298 3175 4302
rect 3291 4298 3295 4302
rect 3379 4298 3383 4302
rect 3799 4298 3803 4302
rect 3839 4222 3843 4226
rect 4543 4222 4547 4226
rect 4719 4222 4723 4226
rect 4815 4222 4819 4226
rect 4903 4222 4907 4226
rect 4951 4222 4955 4226
rect 5087 4222 5091 4226
rect 5095 4222 5099 4226
rect 5223 4222 5227 4226
rect 5295 4222 5299 4226
rect 5359 4222 5363 4226
rect 5495 4222 5499 4226
rect 5663 4222 5667 4226
rect 111 4182 115 4186
rect 347 4182 351 4186
rect 515 4182 519 4186
rect 627 4182 631 4186
rect 699 4182 703 4186
rect 795 4182 799 4186
rect 891 4182 895 4186
rect 963 4182 967 4186
rect 1099 4182 1103 4186
rect 1139 4182 1143 4186
rect 1315 4182 1319 4186
rect 1491 4182 1495 4186
rect 1531 4182 1535 4186
rect 1675 4182 1679 4186
rect 1935 4182 1939 4186
rect 1975 4182 1979 4186
rect 2023 4182 2027 4186
rect 2047 4182 2051 4186
rect 2271 4182 2275 4186
rect 2287 4182 2291 4186
rect 2487 4182 2491 4186
rect 2551 4182 2555 4186
rect 2695 4182 2699 4186
rect 2799 4182 2803 4186
rect 2903 4182 2907 4186
rect 3039 4182 3043 4186
rect 3111 4182 3115 4186
rect 3279 4182 3283 4186
rect 3319 4182 3323 4186
rect 3519 4182 3523 4186
rect 3799 4182 3803 4186
rect 3839 4106 3843 4110
rect 4787 4106 4791 4110
rect 4923 4106 4927 4110
rect 4939 4106 4943 4110
rect 5059 4106 5063 4110
rect 5075 4106 5079 4110
rect 5195 4106 5199 4110
rect 5211 4106 5215 4110
rect 5331 4106 5335 4110
rect 5347 4106 5351 4110
rect 5467 4106 5471 4110
rect 5483 4106 5487 4110
rect 5663 4106 5667 4110
rect 1975 4070 1979 4074
rect 1995 4070 1999 4074
rect 2259 4070 2263 4074
rect 2283 4070 2287 4074
rect 2523 4070 2527 4074
rect 2587 4070 2591 4074
rect 2771 4070 2775 4074
rect 2875 4070 2879 4074
rect 3011 4070 3015 4074
rect 3163 4070 3167 4074
rect 3251 4070 3255 4074
rect 3451 4070 3455 4074
rect 3491 4070 3495 4074
rect 3799 4070 3803 4074
rect 111 4054 115 4058
rect 231 4054 235 4058
rect 375 4054 379 4058
rect 423 4054 427 4058
rect 543 4054 547 4058
rect 615 4054 619 4058
rect 727 4054 731 4058
rect 807 4054 811 4058
rect 919 4054 923 4058
rect 991 4054 995 4058
rect 1127 4054 1131 4058
rect 1167 4054 1171 4058
rect 1335 4054 1339 4058
rect 1343 4054 1347 4058
rect 1503 4054 1507 4058
rect 1559 4054 1563 4058
rect 1671 4054 1675 4058
rect 1815 4054 1819 4058
rect 1935 4054 1939 4058
rect 111 3942 115 3946
rect 203 3942 207 3946
rect 251 3942 255 3946
rect 395 3942 399 3946
rect 451 3942 455 3946
rect 587 3942 591 3946
rect 643 3942 647 3946
rect 779 3942 783 3946
rect 827 3942 831 3946
rect 963 3942 967 3946
rect 1003 3942 1007 3946
rect 1139 3942 1143 3946
rect 1171 3942 1175 3946
rect 1307 3942 1311 3946
rect 1331 3942 1335 3946
rect 1475 3942 1479 3946
rect 1491 3942 1495 3946
rect 1643 3942 1647 3946
rect 1651 3942 1655 3946
rect 1787 3942 1791 3946
rect 1935 3942 1939 3946
rect 3839 3986 3843 3990
rect 4831 3986 4835 3990
rect 4967 3986 4971 3990
rect 5103 3986 5107 3990
rect 5111 3986 5115 3990
rect 5239 3986 5243 3990
rect 5255 3986 5259 3990
rect 5375 3986 5379 3990
rect 5407 3986 5411 3990
rect 5511 3986 5515 3990
rect 5543 3986 5547 3990
rect 5663 3986 5667 3990
rect 1975 3938 1979 3942
rect 2023 3938 2027 3942
rect 2311 3938 2315 3942
rect 2615 3938 2619 3942
rect 2671 3938 2675 3942
rect 2807 3938 2811 3942
rect 2903 3938 2907 3942
rect 2943 3938 2947 3942
rect 3079 3938 3083 3942
rect 3191 3938 3195 3942
rect 3215 3938 3219 3942
rect 3479 3938 3483 3942
rect 3799 3938 3803 3942
rect 111 3830 115 3834
rect 279 3830 283 3834
rect 311 3830 315 3834
rect 479 3830 483 3834
rect 511 3830 515 3834
rect 671 3830 675 3834
rect 735 3830 739 3834
rect 855 3830 859 3834
rect 991 3830 995 3834
rect 1031 3830 1035 3834
rect 1199 3830 1203 3834
rect 1263 3830 1267 3834
rect 1359 3830 1363 3834
rect 1519 3830 1523 3834
rect 1551 3830 1555 3834
rect 1679 3830 1683 3834
rect 1815 3830 1819 3834
rect 1935 3830 1939 3834
rect 3839 3854 3843 3858
rect 4499 3854 4503 3858
rect 4675 3854 4679 3858
rect 4803 3854 4807 3858
rect 4875 3854 4879 3858
rect 4939 3854 4943 3858
rect 5083 3854 5087 3858
rect 5091 3854 5095 3858
rect 5227 3854 5231 3858
rect 5315 3854 5319 3858
rect 5379 3854 5383 3858
rect 5515 3854 5519 3858
rect 5663 3854 5667 3858
rect 1975 3814 1979 3818
rect 1995 3814 1999 3818
rect 2131 3814 2135 3818
rect 2283 3814 2287 3818
rect 2443 3814 2447 3818
rect 2603 3814 2607 3818
rect 2643 3814 2647 3818
rect 2763 3814 2767 3818
rect 2779 3814 2783 3818
rect 2915 3814 2919 3818
rect 2923 3814 2927 3818
rect 3051 3814 3055 3818
rect 3083 3814 3087 3818
rect 3187 3814 3191 3818
rect 3243 3814 3247 3818
rect 3411 3814 3415 3818
rect 3799 3814 3803 3818
rect 3839 3718 3843 3722
rect 4271 3718 4275 3722
rect 4471 3718 4475 3722
rect 4527 3718 4531 3722
rect 4695 3718 4699 3722
rect 4703 3718 4707 3722
rect 4903 3718 4907 3722
rect 4935 3718 4939 3722
rect 5119 3718 5123 3722
rect 5191 3718 5195 3722
rect 5343 3718 5347 3722
rect 5447 3718 5451 3722
rect 5543 3718 5547 3722
rect 5663 3718 5667 3722
rect 111 3694 115 3698
rect 155 3694 159 3698
rect 283 3694 287 3698
rect 291 3694 295 3698
rect 427 3694 431 3698
rect 483 3694 487 3698
rect 563 3694 567 3698
rect 699 3694 703 3698
rect 707 3694 711 3698
rect 835 3694 839 3698
rect 963 3694 967 3698
rect 971 3694 975 3698
rect 1107 3694 1111 3698
rect 1235 3694 1239 3698
rect 1243 3694 1247 3698
rect 1379 3694 1383 3698
rect 1515 3694 1519 3698
rect 1523 3694 1527 3698
rect 1787 3694 1791 3698
rect 1935 3694 1939 3698
rect 1975 3694 1979 3698
rect 2023 3694 2027 3698
rect 2047 3694 2051 3698
rect 2159 3694 2163 3698
rect 2223 3694 2227 3698
rect 2311 3694 2315 3698
rect 2407 3694 2411 3698
rect 2471 3694 2475 3698
rect 2591 3694 2595 3698
rect 2631 3694 2635 3698
rect 2783 3694 2787 3698
rect 2791 3694 2795 3698
rect 2951 3694 2955 3698
rect 2967 3694 2971 3698
rect 3111 3694 3115 3698
rect 3151 3694 3155 3698
rect 3271 3694 3275 3698
rect 3335 3694 3339 3698
rect 3439 3694 3443 3698
rect 3519 3694 3523 3698
rect 3679 3694 3683 3698
rect 3799 3694 3803 3698
rect 3839 3602 3843 3606
rect 3859 3602 3863 3606
rect 3995 3602 3999 3606
rect 4131 3602 4135 3606
rect 4243 3602 4247 3606
rect 4267 3602 4271 3606
rect 4403 3602 4407 3606
rect 4443 3602 4447 3606
rect 4539 3602 4543 3606
rect 4667 3602 4671 3606
rect 4675 3602 4679 3606
rect 4811 3602 4815 3606
rect 4907 3602 4911 3606
rect 4947 3602 4951 3606
rect 5163 3602 5167 3606
rect 5419 3602 5423 3606
rect 5663 3602 5667 3606
rect 1975 3570 1979 3574
rect 2019 3570 2023 3574
rect 2195 3570 2199 3574
rect 2307 3570 2311 3574
rect 2379 3570 2383 3574
rect 2443 3570 2447 3574
rect 2563 3570 2567 3574
rect 2579 3570 2583 3574
rect 2715 3570 2719 3574
rect 2755 3570 2759 3574
rect 2939 3570 2943 3574
rect 3123 3570 3127 3574
rect 3307 3570 3311 3574
rect 3491 3570 3495 3574
rect 3651 3570 3655 3574
rect 3799 3570 3803 3574
rect 3839 3490 3843 3494
rect 3887 3490 3891 3494
rect 4023 3490 4027 3494
rect 4159 3490 4163 3494
rect 4295 3490 4299 3494
rect 4431 3490 4435 3494
rect 4567 3490 4571 3494
rect 4703 3490 4707 3494
rect 4839 3490 4843 3494
rect 4975 3490 4979 3494
rect 5111 3490 5115 3494
rect 5247 3490 5251 3494
rect 5383 3490 5387 3494
rect 5519 3490 5523 3494
rect 5663 3490 5667 3494
rect 1975 3422 1979 3426
rect 2167 3422 2171 3426
rect 2303 3422 2307 3426
rect 2335 3422 2339 3426
rect 2439 3422 2443 3426
rect 2471 3422 2475 3426
rect 2575 3422 2579 3426
rect 2607 3422 2611 3426
rect 2711 3422 2715 3426
rect 2743 3422 2747 3426
rect 2847 3422 2851 3426
rect 2983 3422 2987 3426
rect 3799 3422 3803 3426
rect 3839 3370 3843 3374
rect 3859 3370 3863 3374
rect 3995 3370 3999 3374
rect 4131 3370 4135 3374
rect 4155 3370 4159 3374
rect 4267 3370 4271 3374
rect 4315 3370 4319 3374
rect 4403 3370 4407 3374
rect 4467 3370 4471 3374
rect 4539 3370 4543 3374
rect 4627 3370 4631 3374
rect 4675 3370 4679 3374
rect 4787 3370 4791 3374
rect 4811 3370 4815 3374
rect 4947 3370 4951 3374
rect 5083 3370 5087 3374
rect 5219 3370 5223 3374
rect 5355 3370 5359 3374
rect 5491 3370 5495 3374
rect 5663 3370 5667 3374
rect 1975 3310 1979 3314
rect 2059 3310 2063 3314
rect 2139 3310 2143 3314
rect 2203 3310 2207 3314
rect 2275 3310 2279 3314
rect 2363 3310 2367 3314
rect 2411 3310 2415 3314
rect 2539 3310 2543 3314
rect 2547 3310 2551 3314
rect 2683 3310 2687 3314
rect 2739 3310 2743 3314
rect 2819 3310 2823 3314
rect 2955 3310 2959 3314
rect 3187 3310 3191 3314
rect 3427 3310 3431 3314
rect 3651 3310 3655 3314
rect 3799 3310 3803 3314
rect 111 3294 115 3298
rect 159 3294 163 3298
rect 183 3294 187 3298
rect 295 3294 299 3298
rect 319 3294 323 3298
rect 431 3294 435 3298
rect 455 3294 459 3298
rect 567 3294 571 3298
rect 591 3294 595 3298
rect 703 3294 707 3298
rect 727 3294 731 3298
rect 839 3294 843 3298
rect 863 3294 867 3298
rect 975 3294 979 3298
rect 999 3294 1003 3298
rect 1111 3294 1115 3298
rect 1135 3294 1139 3298
rect 1247 3294 1251 3298
rect 1271 3294 1275 3298
rect 1383 3294 1387 3298
rect 1407 3294 1411 3298
rect 1519 3294 1523 3298
rect 1543 3294 1547 3298
rect 1935 3294 1939 3298
rect 3839 3246 3843 3250
rect 3887 3246 3891 3250
rect 4023 3246 4027 3250
rect 4183 3246 4187 3250
rect 4343 3246 4347 3250
rect 4495 3246 4499 3250
rect 4655 3246 4659 3250
rect 4807 3246 4811 3250
rect 4815 3246 4819 3250
rect 4943 3246 4947 3250
rect 4975 3246 4979 3250
rect 5079 3246 5083 3250
rect 5215 3246 5219 3250
rect 5351 3246 5355 3250
rect 5663 3246 5667 3250
rect 1975 3194 1979 3198
rect 2023 3194 2027 3198
rect 2087 3194 2091 3198
rect 2159 3194 2163 3198
rect 2231 3194 2235 3198
rect 2303 3194 2307 3198
rect 2391 3194 2395 3198
rect 2455 3194 2459 3198
rect 2567 3194 2571 3198
rect 2615 3194 2619 3198
rect 2767 3194 2771 3198
rect 2783 3194 2787 3198
rect 2951 3194 2955 3198
rect 2983 3194 2987 3198
rect 3127 3194 3131 3198
rect 3215 3194 3219 3198
rect 3311 3194 3315 3198
rect 3455 3194 3459 3198
rect 3503 3194 3507 3198
rect 3679 3194 3683 3198
rect 3799 3194 3803 3198
rect 111 3154 115 3158
rect 131 3154 135 3158
rect 267 3154 271 3158
rect 291 3154 295 3158
rect 403 3154 407 3158
rect 459 3154 463 3158
rect 539 3154 543 3158
rect 627 3154 631 3158
rect 675 3154 679 3158
rect 811 3154 815 3158
rect 947 3154 951 3158
rect 995 3154 999 3158
rect 1083 3154 1087 3158
rect 1187 3154 1191 3158
rect 1219 3154 1223 3158
rect 1355 3154 1359 3158
rect 1387 3154 1391 3158
rect 1491 3154 1495 3158
rect 1595 3154 1599 3158
rect 1787 3154 1791 3158
rect 1935 3154 1939 3158
rect 3839 3130 3843 3134
rect 4699 3130 4703 3134
rect 4779 3130 4783 3134
rect 4835 3130 4839 3134
rect 4915 3130 4919 3134
rect 4971 3130 4975 3134
rect 5051 3130 5055 3134
rect 5107 3130 5111 3134
rect 5187 3130 5191 3134
rect 5243 3130 5247 3134
rect 5323 3130 5327 3134
rect 5379 3130 5383 3134
rect 5515 3130 5519 3134
rect 5663 3130 5667 3134
rect 1975 3062 1979 3066
rect 1995 3062 1999 3066
rect 2131 3062 2135 3066
rect 2275 3062 2279 3066
rect 2427 3062 2431 3066
rect 2587 3062 2591 3066
rect 2755 3062 2759 3066
rect 2811 3062 2815 3066
rect 2923 3062 2927 3066
rect 3003 3062 3007 3066
rect 3099 3062 3103 3066
rect 3203 3062 3207 3066
rect 3283 3062 3287 3066
rect 3403 3062 3407 3066
rect 3475 3062 3479 3066
rect 3603 3062 3607 3066
rect 3651 3062 3655 3066
rect 3799 3062 3803 3066
rect 111 3042 115 3046
rect 319 3042 323 3046
rect 327 3042 331 3046
rect 487 3042 491 3046
rect 647 3042 651 3046
rect 655 3042 659 3046
rect 807 3042 811 3046
rect 839 3042 843 3046
rect 959 3042 963 3046
rect 1023 3042 1027 3046
rect 1103 3042 1107 3046
rect 1215 3042 1219 3046
rect 1247 3042 1251 3046
rect 1391 3042 1395 3046
rect 1415 3042 1419 3046
rect 1535 3042 1539 3046
rect 1623 3042 1627 3046
rect 1679 3042 1683 3046
rect 1815 3042 1819 3046
rect 1935 3042 1939 3046
rect 3839 3018 3843 3022
rect 4367 3018 4371 3022
rect 4567 3018 4571 3022
rect 4727 3018 4731 3022
rect 4783 3018 4787 3022
rect 4863 3018 4867 3022
rect 4999 3018 5003 3022
rect 5023 3018 5027 3022
rect 5135 3018 5139 3022
rect 5271 3018 5275 3022
rect 5279 3018 5283 3022
rect 5407 3018 5411 3022
rect 5535 3018 5539 3022
rect 5543 3018 5547 3022
rect 5663 3018 5667 3022
rect 1975 2942 1979 2946
rect 2839 2942 2843 2946
rect 2847 2942 2851 2946
rect 2983 2942 2987 2946
rect 3031 2942 3035 2946
rect 3119 2942 3123 2946
rect 3231 2942 3235 2946
rect 3255 2942 3259 2946
rect 3391 2942 3395 2946
rect 3431 2942 3435 2946
rect 3527 2942 3531 2946
rect 3631 2942 3635 2946
rect 3671 2942 3675 2946
rect 3799 2942 3803 2946
rect 111 2930 115 2934
rect 155 2930 159 2934
rect 299 2930 303 2934
rect 379 2930 383 2934
rect 459 2930 463 2934
rect 595 2930 599 2934
rect 619 2930 623 2934
rect 779 2930 783 2934
rect 811 2930 815 2934
rect 931 2930 935 2934
rect 1019 2930 1023 2934
rect 1075 2930 1079 2934
rect 1219 2930 1223 2934
rect 1363 2930 1367 2934
rect 1411 2930 1415 2934
rect 1507 2930 1511 2934
rect 1611 2930 1615 2934
rect 1651 2930 1655 2934
rect 1787 2930 1791 2934
rect 1935 2930 1939 2934
rect 3839 2906 3843 2910
rect 4035 2906 4039 2910
rect 4315 2906 4319 2910
rect 4339 2906 4343 2910
rect 4539 2906 4543 2910
rect 4603 2906 4607 2910
rect 4755 2906 4759 2910
rect 4907 2906 4911 2910
rect 4995 2906 4999 2910
rect 5219 2906 5223 2910
rect 5251 2906 5255 2910
rect 5507 2906 5511 2910
rect 5515 2906 5519 2910
rect 5663 2906 5667 2910
rect 1975 2830 1979 2834
rect 2011 2830 2015 2834
rect 2251 2830 2255 2834
rect 2491 2830 2495 2834
rect 2731 2830 2735 2834
rect 2819 2830 2823 2834
rect 2955 2830 2959 2834
rect 2971 2830 2975 2834
rect 3091 2830 3095 2834
rect 3227 2830 3231 2834
rect 3363 2830 3367 2834
rect 3499 2830 3503 2834
rect 3643 2830 3647 2834
rect 3799 2830 3803 2834
rect 111 2786 115 2790
rect 183 2786 187 2790
rect 287 2786 291 2790
rect 407 2786 411 2790
rect 423 2786 427 2790
rect 559 2786 563 2790
rect 623 2786 627 2790
rect 695 2786 699 2790
rect 831 2786 835 2790
rect 839 2786 843 2790
rect 1047 2786 1051 2790
rect 1247 2786 1251 2790
rect 1439 2786 1443 2790
rect 1639 2786 1643 2790
rect 1815 2786 1819 2790
rect 1935 2786 1939 2790
rect 3839 2786 3843 2790
rect 3967 2786 3971 2790
rect 4063 2786 4067 2790
rect 4255 2786 4259 2790
rect 4343 2786 4347 2790
rect 4567 2786 4571 2790
rect 4631 2786 4635 2790
rect 4895 2786 4899 2790
rect 4935 2786 4939 2790
rect 5231 2786 5235 2790
rect 5247 2786 5251 2790
rect 5543 2786 5547 2790
rect 5663 2786 5667 2790
rect 1975 2718 1979 2722
rect 2023 2718 2027 2722
rect 2039 2718 2043 2722
rect 2159 2718 2163 2722
rect 2279 2718 2283 2722
rect 2295 2718 2299 2722
rect 2431 2718 2435 2722
rect 2519 2718 2523 2722
rect 2567 2718 2571 2722
rect 2703 2718 2707 2722
rect 2759 2718 2763 2722
rect 2839 2718 2843 2722
rect 2975 2718 2979 2722
rect 2999 2718 3003 2722
rect 3111 2718 3115 2722
rect 3247 2718 3251 2722
rect 3383 2718 3387 2722
rect 3799 2718 3803 2722
rect 111 2654 115 2658
rect 259 2654 263 2658
rect 395 2654 399 2658
rect 531 2654 535 2658
rect 539 2654 543 2658
rect 667 2654 671 2658
rect 699 2654 703 2658
rect 803 2654 807 2658
rect 883 2654 887 2658
rect 1091 2654 1095 2658
rect 1323 2654 1327 2658
rect 1563 2654 1567 2658
rect 1787 2654 1791 2658
rect 1935 2654 1939 2658
rect 3839 2670 3843 2674
rect 3939 2670 3943 2674
rect 4027 2670 4031 2674
rect 4227 2670 4231 2674
rect 4275 2670 4279 2674
rect 4539 2670 4543 2674
rect 4555 2670 4559 2674
rect 4867 2670 4871 2674
rect 5203 2670 5207 2674
rect 5515 2670 5519 2674
rect 5663 2670 5667 2674
rect 1975 2606 1979 2610
rect 1995 2606 1999 2610
rect 2131 2606 2135 2610
rect 2203 2606 2207 2610
rect 2267 2606 2271 2610
rect 2403 2606 2407 2610
rect 2419 2606 2423 2610
rect 2539 2606 2543 2610
rect 2627 2606 2631 2610
rect 2675 2606 2679 2610
rect 2811 2606 2815 2610
rect 2827 2606 2831 2610
rect 2947 2606 2951 2610
rect 3019 2606 3023 2610
rect 3083 2606 3087 2610
rect 3211 2606 3215 2610
rect 3219 2606 3223 2610
rect 3355 2606 3359 2610
rect 3403 2606 3407 2610
rect 3799 2606 3803 2610
rect 3839 2554 3843 2558
rect 4055 2554 4059 2558
rect 4303 2554 4307 2558
rect 4335 2554 4339 2558
rect 4559 2554 4563 2558
rect 4583 2554 4587 2558
rect 4799 2554 4803 2558
rect 4895 2554 4899 2558
rect 5047 2554 5051 2558
rect 5231 2554 5235 2558
rect 5303 2554 5307 2558
rect 5543 2554 5547 2558
rect 5663 2554 5667 2558
rect 111 2530 115 2534
rect 567 2530 571 2534
rect 695 2530 699 2534
rect 727 2530 731 2534
rect 847 2530 851 2534
rect 911 2530 915 2534
rect 999 2530 1003 2534
rect 1119 2530 1123 2534
rect 1159 2530 1163 2534
rect 1327 2530 1331 2534
rect 1351 2530 1355 2534
rect 1495 2530 1499 2534
rect 1591 2530 1595 2534
rect 1663 2530 1667 2534
rect 1815 2530 1819 2534
rect 1935 2530 1939 2534
rect 1975 2486 1979 2490
rect 2023 2486 2027 2490
rect 2231 2486 2235 2490
rect 2319 2486 2323 2490
rect 2447 2486 2451 2490
rect 2567 2486 2571 2490
rect 2655 2486 2659 2490
rect 2799 2486 2803 2490
rect 2855 2486 2859 2490
rect 3023 2486 3027 2490
rect 3047 2486 3051 2490
rect 3239 2486 3243 2490
rect 3431 2486 3435 2490
rect 3455 2486 3459 2490
rect 3671 2486 3675 2490
rect 3799 2486 3803 2490
rect 111 2410 115 2414
rect 355 2410 359 2414
rect 507 2410 511 2414
rect 667 2410 671 2414
rect 675 2410 679 2414
rect 819 2410 823 2414
rect 859 2410 863 2414
rect 971 2410 975 2414
rect 1059 2410 1063 2414
rect 1131 2410 1135 2414
rect 1267 2410 1271 2414
rect 1299 2410 1303 2414
rect 1467 2410 1471 2414
rect 1483 2410 1487 2414
rect 1635 2410 1639 2414
rect 1699 2410 1703 2414
rect 1787 2410 1791 2414
rect 1935 2410 1939 2414
rect 3839 2426 3843 2430
rect 4307 2426 4311 2430
rect 4491 2426 4495 2430
rect 4531 2426 4535 2430
rect 4635 2426 4639 2430
rect 4771 2426 4775 2430
rect 4795 2426 4799 2430
rect 4963 2426 4967 2430
rect 5019 2426 5023 2430
rect 5139 2426 5143 2430
rect 5275 2426 5279 2430
rect 5323 2426 5327 2430
rect 5515 2426 5519 2430
rect 5663 2426 5667 2430
rect 1975 2366 1979 2370
rect 2291 2366 2295 2370
rect 2331 2366 2335 2370
rect 2539 2366 2543 2370
rect 2739 2366 2743 2370
rect 2771 2366 2775 2370
rect 2931 2366 2935 2370
rect 2995 2366 2999 2370
rect 3123 2366 3127 2370
rect 3211 2366 3215 2370
rect 3307 2366 3311 2370
rect 3427 2366 3431 2370
rect 3491 2366 3495 2370
rect 3643 2366 3647 2370
rect 3651 2366 3655 2370
rect 3799 2366 3803 2370
rect 111 2290 115 2294
rect 159 2290 163 2294
rect 335 2290 339 2294
rect 383 2290 387 2294
rect 535 2290 539 2294
rect 543 2290 547 2294
rect 703 2290 707 2294
rect 759 2290 763 2294
rect 887 2290 891 2294
rect 975 2290 979 2294
rect 1087 2290 1091 2294
rect 1199 2290 1203 2294
rect 1295 2290 1299 2294
rect 1431 2290 1435 2294
rect 1511 2290 1515 2294
rect 1671 2290 1675 2294
rect 1727 2290 1731 2294
rect 1935 2290 1939 2294
rect 3839 2294 3843 2298
rect 3887 2294 3891 2298
rect 4071 2294 4075 2298
rect 4271 2294 4275 2298
rect 4463 2294 4467 2298
rect 4519 2294 4523 2298
rect 4655 2294 4659 2298
rect 4663 2294 4667 2298
rect 4823 2294 4827 2298
rect 4839 2294 4843 2298
rect 4991 2294 4995 2298
rect 5015 2294 5019 2298
rect 5167 2294 5171 2298
rect 5183 2294 5187 2298
rect 5351 2294 5355 2298
rect 5359 2294 5363 2298
rect 5535 2294 5539 2298
rect 5543 2294 5547 2298
rect 5663 2294 5667 2298
rect 1975 2226 1979 2230
rect 2359 2226 2363 2230
rect 2463 2226 2467 2230
rect 2567 2226 2571 2230
rect 2599 2226 2603 2230
rect 2735 2226 2739 2230
rect 2767 2226 2771 2230
rect 2959 2226 2963 2230
rect 3151 2226 3155 2230
rect 3335 2226 3339 2230
rect 3519 2226 3523 2230
rect 3679 2226 3683 2230
rect 3799 2226 3803 2230
rect 3839 2182 3843 2186
rect 3859 2182 3863 2186
rect 4043 2182 4047 2186
rect 4243 2182 4247 2186
rect 4251 2182 4255 2186
rect 4435 2182 4439 2186
rect 4459 2182 4463 2186
rect 4627 2182 4631 2186
rect 4659 2182 4663 2186
rect 4811 2182 4815 2186
rect 4851 2182 4855 2186
rect 4987 2182 4991 2186
rect 5035 2182 5039 2186
rect 5155 2182 5159 2186
rect 5219 2182 5223 2186
rect 5331 2182 5335 2186
rect 5411 2182 5415 2186
rect 5507 2182 5511 2186
rect 5663 2182 5667 2186
rect 111 2158 115 2162
rect 131 2158 135 2162
rect 299 2158 303 2162
rect 307 2158 311 2162
rect 499 2158 503 2162
rect 515 2158 519 2162
rect 715 2158 719 2162
rect 731 2158 735 2162
rect 931 2158 935 2162
rect 947 2158 951 2162
rect 1155 2158 1159 2162
rect 1171 2158 1175 2162
rect 1387 2158 1391 2162
rect 1403 2158 1407 2162
rect 1627 2158 1631 2162
rect 1643 2158 1647 2162
rect 1935 2158 1939 2162
rect 1975 2082 1979 2086
rect 2419 2082 2423 2086
rect 2435 2082 2439 2086
rect 2571 2082 2575 2086
rect 2611 2082 2615 2086
rect 2707 2082 2711 2086
rect 2795 2082 2799 2086
rect 2979 2082 2983 2086
rect 3155 2082 3159 2086
rect 3323 2082 3327 2086
rect 3499 2082 3503 2086
rect 3651 2082 3655 2086
rect 3799 2082 3803 2086
rect 111 2038 115 2042
rect 159 2038 163 2042
rect 327 2038 331 2042
rect 343 2038 347 2042
rect 527 2038 531 2042
rect 567 2038 571 2042
rect 743 2038 747 2042
rect 807 2038 811 2042
rect 959 2038 963 2042
rect 1063 2038 1067 2042
rect 1183 2038 1187 2042
rect 1335 2038 1339 2042
rect 1415 2038 1419 2042
rect 1607 2038 1611 2042
rect 1655 2038 1659 2042
rect 1935 2038 1939 2042
rect 3839 2050 3843 2054
rect 3887 2050 3891 2054
rect 4071 2050 4075 2054
rect 4279 2050 4283 2054
rect 4287 2050 4291 2054
rect 4423 2050 4427 2054
rect 4487 2050 4491 2054
rect 4559 2050 4563 2054
rect 4687 2050 4691 2054
rect 4695 2050 4699 2054
rect 4839 2050 4843 2054
rect 4879 2050 4883 2054
rect 5063 2050 5067 2054
rect 5247 2050 5251 2054
rect 5439 2050 5443 2054
rect 5663 2050 5667 2054
rect 1975 1958 1979 1962
rect 2359 1958 2363 1962
rect 2447 1958 2451 1962
rect 2495 1958 2499 1962
rect 2631 1958 2635 1962
rect 2639 1958 2643 1962
rect 2767 1958 2771 1962
rect 2823 1958 2827 1962
rect 2903 1958 2907 1962
rect 3007 1958 3011 1962
rect 3039 1958 3043 1962
rect 3175 1958 3179 1962
rect 3183 1958 3187 1962
rect 3319 1958 3323 1962
rect 3351 1958 3355 1962
rect 3527 1958 3531 1962
rect 3679 1958 3683 1962
rect 3799 1958 3803 1962
rect 111 1922 115 1926
rect 131 1922 135 1926
rect 315 1922 319 1926
rect 331 1922 335 1926
rect 499 1922 503 1926
rect 539 1922 543 1926
rect 667 1922 671 1926
rect 779 1922 783 1926
rect 843 1922 847 1926
rect 1027 1922 1031 1926
rect 1035 1922 1039 1926
rect 1219 1922 1223 1926
rect 1307 1922 1311 1926
rect 1411 1922 1415 1926
rect 1579 1922 1583 1926
rect 1603 1922 1607 1926
rect 1935 1922 1939 1926
rect 3839 1918 3843 1922
rect 3955 1918 3959 1922
rect 4195 1918 4199 1922
rect 4259 1918 4263 1922
rect 4395 1918 4399 1922
rect 4467 1918 4471 1922
rect 4531 1918 4535 1922
rect 4667 1918 4671 1922
rect 4771 1918 4775 1922
rect 4811 1918 4815 1922
rect 5091 1918 5095 1922
rect 5411 1918 5415 1922
rect 5663 1918 5667 1922
rect 1975 1846 1979 1850
rect 2211 1846 2215 1850
rect 2331 1846 2335 1850
rect 2355 1846 2359 1850
rect 2467 1846 2471 1850
rect 2499 1846 2503 1850
rect 2603 1846 2607 1850
rect 2643 1846 2647 1850
rect 2739 1846 2743 1850
rect 2787 1846 2791 1850
rect 2875 1846 2879 1850
rect 2931 1846 2935 1850
rect 3011 1846 3015 1850
rect 3083 1846 3087 1850
rect 3147 1846 3151 1850
rect 3291 1846 3295 1850
rect 3799 1846 3803 1850
rect 111 1798 115 1802
rect 359 1798 363 1802
rect 527 1798 531 1802
rect 535 1798 539 1802
rect 695 1798 699 1802
rect 855 1798 859 1802
rect 871 1798 875 1802
rect 1015 1798 1019 1802
rect 1055 1798 1059 1802
rect 1183 1798 1187 1802
rect 1247 1798 1251 1802
rect 1351 1798 1355 1802
rect 1439 1798 1443 1802
rect 1519 1798 1523 1802
rect 1631 1798 1635 1802
rect 1935 1798 1939 1802
rect 3839 1806 3843 1810
rect 3983 1806 3987 1810
rect 4223 1806 4227 1810
rect 4367 1806 4371 1810
rect 4495 1806 4499 1810
rect 4575 1806 4579 1810
rect 4783 1806 4787 1810
rect 4799 1806 4803 1810
rect 4983 1806 4987 1810
rect 5119 1806 5123 1810
rect 5175 1806 5179 1810
rect 5367 1806 5371 1810
rect 5439 1806 5443 1810
rect 5543 1806 5547 1810
rect 5663 1806 5667 1810
rect 1975 1734 1979 1738
rect 2023 1734 2027 1738
rect 2215 1734 2219 1738
rect 2239 1734 2243 1738
rect 2383 1734 2387 1738
rect 2407 1734 2411 1738
rect 2527 1734 2531 1738
rect 2599 1734 2603 1738
rect 2671 1734 2675 1738
rect 2791 1734 2795 1738
rect 2815 1734 2819 1738
rect 2959 1734 2963 1738
rect 2975 1734 2979 1738
rect 3111 1734 3115 1738
rect 3151 1734 3155 1738
rect 3335 1734 3339 1738
rect 3519 1734 3523 1738
rect 3799 1734 3803 1738
rect 111 1670 115 1674
rect 427 1670 431 1674
rect 507 1670 511 1674
rect 611 1670 615 1674
rect 667 1670 671 1674
rect 803 1670 807 1674
rect 827 1670 831 1674
rect 987 1670 991 1674
rect 995 1670 999 1674
rect 1155 1670 1159 1674
rect 1187 1670 1191 1674
rect 1323 1670 1327 1674
rect 1379 1670 1383 1674
rect 1491 1670 1495 1674
rect 1935 1670 1939 1674
rect 3839 1678 3843 1682
rect 4339 1678 4343 1682
rect 4547 1678 4551 1682
rect 4603 1678 4607 1682
rect 4755 1678 4759 1682
rect 4787 1678 4791 1682
rect 4955 1678 4959 1682
rect 4971 1678 4975 1682
rect 5147 1678 5151 1682
rect 5155 1678 5159 1682
rect 5339 1678 5343 1682
rect 5515 1678 5519 1682
rect 5663 1678 5667 1682
rect 1975 1622 1979 1626
rect 1995 1622 1999 1626
rect 2163 1622 2167 1626
rect 2187 1622 2191 1626
rect 2371 1622 2375 1626
rect 2379 1622 2383 1626
rect 2571 1622 2575 1626
rect 2587 1622 2591 1626
rect 2763 1622 2767 1626
rect 2803 1622 2807 1626
rect 2947 1622 2951 1626
rect 3019 1622 3023 1626
rect 3123 1622 3127 1626
rect 3235 1622 3239 1626
rect 3307 1622 3311 1626
rect 3451 1622 3455 1626
rect 3491 1622 3495 1626
rect 3651 1622 3655 1626
rect 3799 1622 3803 1626
rect 111 1550 115 1554
rect 359 1550 363 1554
rect 455 1550 459 1554
rect 631 1550 635 1554
rect 639 1550 643 1554
rect 831 1550 835 1554
rect 887 1550 891 1554
rect 1023 1550 1027 1554
rect 1135 1550 1139 1554
rect 1215 1550 1219 1554
rect 1367 1550 1371 1554
rect 1407 1550 1411 1554
rect 1599 1550 1603 1554
rect 1815 1550 1819 1554
rect 1935 1550 1939 1554
rect 3839 1550 3843 1554
rect 3887 1550 3891 1554
rect 4031 1550 4035 1554
rect 4199 1550 4203 1554
rect 4367 1550 4371 1554
rect 4527 1550 4531 1554
rect 4631 1550 4635 1554
rect 4695 1550 4699 1554
rect 4815 1550 4819 1554
rect 4863 1550 4867 1554
rect 4999 1550 5003 1554
rect 5031 1550 5035 1554
rect 5183 1550 5187 1554
rect 5207 1550 5211 1554
rect 5367 1550 5371 1554
rect 5383 1550 5387 1554
rect 5543 1550 5547 1554
rect 5663 1550 5667 1554
rect 111 1438 115 1442
rect 131 1438 135 1442
rect 307 1438 311 1442
rect 331 1438 335 1442
rect 499 1438 503 1442
rect 603 1438 607 1442
rect 683 1438 687 1442
rect 859 1438 863 1442
rect 1027 1438 1031 1442
rect 1107 1438 1111 1442
rect 1187 1438 1191 1442
rect 1339 1438 1343 1442
rect 1491 1438 1495 1442
rect 1571 1438 1575 1442
rect 1651 1438 1655 1442
rect 1787 1438 1791 1442
rect 1935 1438 1939 1442
rect 111 1318 115 1322
rect 159 1318 163 1322
rect 335 1318 339 1322
rect 375 1318 379 1322
rect 527 1318 531 1322
rect 599 1318 603 1322
rect 711 1318 715 1322
rect 807 1318 811 1322
rect 887 1318 891 1322
rect 999 1318 1003 1322
rect 1055 1318 1059 1322
rect 1175 1318 1179 1322
rect 1215 1318 1219 1322
rect 1343 1318 1347 1322
rect 1367 1318 1371 1322
rect 1511 1318 1515 1322
rect 1519 1318 1523 1322
rect 1671 1318 1675 1322
rect 1679 1318 1683 1322
rect 1815 1318 1819 1322
rect 1935 1318 1939 1322
rect 3839 1434 3843 1438
rect 3859 1434 3863 1438
rect 4003 1434 4007 1438
rect 4171 1434 4175 1438
rect 4179 1434 4183 1438
rect 4339 1434 4343 1438
rect 4355 1434 4359 1438
rect 4499 1434 4503 1438
rect 4531 1434 4535 1438
rect 4667 1434 4671 1438
rect 4707 1434 4711 1438
rect 4835 1434 4839 1438
rect 4875 1434 4879 1438
rect 5003 1434 5007 1438
rect 5043 1434 5047 1438
rect 5179 1434 5183 1438
rect 5203 1434 5207 1438
rect 5355 1434 5359 1438
rect 5371 1434 5375 1438
rect 5515 1434 5519 1438
rect 5663 1434 5667 1438
rect 3839 1322 3843 1326
rect 3887 1322 3891 1326
rect 4031 1322 4035 1326
rect 4175 1322 4179 1326
rect 4207 1322 4211 1326
rect 4383 1322 4387 1326
rect 4471 1322 4475 1326
rect 4559 1322 4563 1326
rect 4735 1322 4739 1326
rect 4751 1322 4755 1326
rect 4903 1322 4907 1326
rect 5023 1322 5027 1326
rect 5071 1322 5075 1326
rect 5231 1322 5235 1326
rect 5287 1322 5291 1326
rect 5399 1322 5403 1326
rect 5543 1322 5547 1326
rect 5663 1322 5667 1326
rect 1975 1306 1979 1310
rect 2023 1306 2027 1310
rect 2191 1306 2195 1310
rect 2399 1306 2403 1310
rect 2615 1306 2619 1310
rect 2831 1306 2835 1310
rect 3047 1306 3051 1310
rect 3263 1306 3267 1310
rect 3271 1306 3275 1310
rect 3407 1306 3411 1310
rect 3479 1306 3483 1310
rect 3543 1306 3547 1310
rect 3679 1306 3683 1310
rect 3799 1306 3803 1310
rect 111 1206 115 1210
rect 131 1206 135 1210
rect 347 1206 351 1210
rect 563 1206 567 1210
rect 571 1206 575 1210
rect 779 1206 783 1210
rect 971 1206 975 1210
rect 987 1206 991 1210
rect 1147 1206 1151 1210
rect 1195 1206 1199 1210
rect 1315 1206 1319 1210
rect 1395 1206 1399 1210
rect 1483 1206 1487 1210
rect 1603 1206 1607 1210
rect 1643 1206 1647 1210
rect 1787 1206 1791 1210
rect 1935 1206 1939 1210
rect 3839 1198 3843 1202
rect 3859 1198 3863 1202
rect 4147 1198 4151 1202
rect 4427 1198 4431 1202
rect 4443 1198 4447 1202
rect 4563 1198 4567 1202
rect 4699 1198 4703 1202
rect 4723 1198 4727 1202
rect 4835 1198 4839 1202
rect 4971 1198 4975 1202
rect 4995 1198 4999 1202
rect 5107 1198 5111 1202
rect 5243 1198 5247 1202
rect 5259 1198 5263 1202
rect 5379 1198 5383 1202
rect 5515 1198 5519 1202
rect 5663 1198 5667 1202
rect 1975 1182 1979 1186
rect 1995 1182 1999 1186
rect 2227 1182 2231 1186
rect 2467 1182 2471 1186
rect 2691 1182 2695 1186
rect 2907 1182 2911 1186
rect 3107 1182 3111 1186
rect 3243 1182 3247 1186
rect 3299 1182 3303 1186
rect 3379 1182 3383 1186
rect 3483 1182 3487 1186
rect 3515 1182 3519 1186
rect 3651 1182 3655 1186
rect 3799 1182 3803 1186
rect 111 1070 115 1074
rect 159 1070 163 1074
rect 375 1070 379 1074
rect 471 1070 475 1074
rect 591 1070 595 1074
rect 607 1070 611 1074
rect 743 1070 747 1074
rect 807 1070 811 1074
rect 887 1070 891 1074
rect 1015 1070 1019 1074
rect 1031 1070 1035 1074
rect 1223 1070 1227 1074
rect 1423 1070 1427 1074
rect 1631 1070 1635 1074
rect 1815 1070 1819 1074
rect 1935 1070 1939 1074
rect 1975 1070 1979 1074
rect 2023 1070 2027 1074
rect 2183 1070 2187 1074
rect 2255 1070 2259 1074
rect 2319 1070 2323 1074
rect 2455 1070 2459 1074
rect 2495 1070 2499 1074
rect 2599 1070 2603 1074
rect 2719 1070 2723 1074
rect 2743 1070 2747 1074
rect 2887 1070 2891 1074
rect 2935 1070 2939 1074
rect 3031 1070 3035 1074
rect 3135 1070 3139 1074
rect 3175 1070 3179 1074
rect 3319 1070 3323 1074
rect 3327 1070 3331 1074
rect 3463 1070 3467 1074
rect 3511 1070 3515 1074
rect 3679 1070 3683 1074
rect 3799 1070 3803 1074
rect 3839 1070 3843 1074
rect 4367 1070 4371 1074
rect 4455 1070 4459 1074
rect 4503 1070 4507 1074
rect 4591 1070 4595 1074
rect 4639 1070 4643 1074
rect 4727 1070 4731 1074
rect 4775 1070 4779 1074
rect 4863 1070 4867 1074
rect 4911 1070 4915 1074
rect 4999 1070 5003 1074
rect 5135 1070 5139 1074
rect 5271 1070 5275 1074
rect 5407 1070 5411 1074
rect 5543 1070 5547 1074
rect 5663 1070 5667 1074
rect 111 946 115 950
rect 259 946 263 950
rect 395 946 399 950
rect 443 946 447 950
rect 531 946 535 950
rect 579 946 583 950
rect 667 946 671 950
rect 715 946 719 950
rect 803 946 807 950
rect 859 946 863 950
rect 939 946 943 950
rect 1003 946 1007 950
rect 1935 946 1939 950
rect 1975 946 1979 950
rect 1995 946 1999 950
rect 2131 946 2135 950
rect 2155 946 2159 950
rect 2267 946 2271 950
rect 2291 946 2295 950
rect 2403 946 2407 950
rect 2427 946 2431 950
rect 2539 946 2543 950
rect 2571 946 2575 950
rect 2675 946 2679 950
rect 2715 946 2719 950
rect 2811 946 2815 950
rect 2859 946 2863 950
rect 2947 946 2951 950
rect 3003 946 3007 950
rect 3083 946 3087 950
rect 3147 946 3151 950
rect 3219 946 3223 950
rect 3291 946 3295 950
rect 3355 946 3359 950
rect 3435 946 3439 950
rect 3491 946 3495 950
rect 3799 946 3803 950
rect 3839 946 3843 950
rect 4019 946 4023 950
rect 4155 946 4159 950
rect 4291 946 4295 950
rect 4339 946 4343 950
rect 4427 946 4431 950
rect 4475 946 4479 950
rect 4563 946 4567 950
rect 4611 946 4615 950
rect 4699 946 4703 950
rect 4747 946 4751 950
rect 4883 946 4887 950
rect 5663 946 5667 950
rect 1975 834 1979 838
rect 2023 834 2027 838
rect 2159 834 2163 838
rect 2167 834 2171 838
rect 2295 834 2299 838
rect 2335 834 2339 838
rect 2431 834 2435 838
rect 2495 834 2499 838
rect 2567 834 2571 838
rect 2655 834 2659 838
rect 2703 834 2707 838
rect 2823 834 2827 838
rect 2839 834 2843 838
rect 2975 834 2979 838
rect 2991 834 2995 838
rect 3111 834 3115 838
rect 3247 834 3251 838
rect 3383 834 3387 838
rect 3519 834 3523 838
rect 3799 834 3803 838
rect 111 822 115 826
rect 239 822 243 826
rect 287 822 291 826
rect 423 822 427 826
rect 439 822 443 826
rect 559 822 563 826
rect 647 822 651 826
rect 695 822 699 826
rect 831 822 835 826
rect 855 822 859 826
rect 967 822 971 826
rect 1063 822 1067 826
rect 1935 822 1939 826
rect 3839 818 3843 822
rect 3887 818 3891 822
rect 4023 818 4027 822
rect 4047 818 4051 822
rect 4159 818 4163 822
rect 4183 818 4187 822
rect 4295 818 4299 822
rect 4319 818 4323 822
rect 4431 818 4435 822
rect 4455 818 4459 822
rect 4567 818 4571 822
rect 4591 818 4595 822
rect 4703 818 4707 822
rect 4727 818 4731 822
rect 4839 818 4843 822
rect 5663 818 5667 822
rect 3839 706 3843 710
rect 3859 706 3863 710
rect 3995 706 3999 710
rect 4131 706 4135 710
rect 4267 706 4271 710
rect 4403 706 4407 710
rect 4539 706 4543 710
rect 4675 706 4679 710
rect 4811 706 4815 710
rect 4947 706 4951 710
rect 5083 706 5087 710
rect 5663 706 5667 710
rect 111 690 115 694
rect 131 690 135 694
rect 211 690 215 694
rect 347 690 351 694
rect 411 690 415 694
rect 587 690 591 694
rect 619 690 623 694
rect 827 690 831 694
rect 1035 690 1039 694
rect 1067 690 1071 694
rect 1315 690 1319 694
rect 1563 690 1567 694
rect 1787 690 1791 694
rect 1935 690 1939 694
rect 1975 694 1979 698
rect 1995 694 1999 698
rect 2139 694 2143 698
rect 2299 694 2303 698
rect 2307 694 2311 698
rect 2467 694 2471 698
rect 2627 694 2631 698
rect 2635 694 2639 698
rect 2795 694 2799 698
rect 2963 694 2967 698
rect 2979 694 2983 698
rect 3323 694 3327 698
rect 3651 694 3655 698
rect 3799 694 3803 698
rect 1975 582 1979 586
rect 2023 582 2027 586
rect 2327 582 2331 586
rect 2335 582 2339 586
rect 2527 582 2531 586
rect 2663 582 2667 586
rect 2711 582 2715 586
rect 2887 582 2891 586
rect 3007 582 3011 586
rect 3063 582 3067 586
rect 3231 582 3235 586
rect 3351 582 3355 586
rect 3407 582 3411 586
rect 3583 582 3587 586
rect 3679 582 3683 586
rect 3799 582 3803 586
rect 111 574 115 578
rect 159 574 163 578
rect 375 574 379 578
rect 407 574 411 578
rect 615 574 619 578
rect 671 574 675 578
rect 855 574 859 578
rect 935 574 939 578
rect 1095 574 1099 578
rect 1191 574 1195 578
rect 1343 574 1347 578
rect 1447 574 1451 578
rect 1591 574 1595 578
rect 1711 574 1715 578
rect 1815 574 1819 578
rect 1935 574 1939 578
rect 3839 574 3843 578
rect 3887 574 3891 578
rect 4023 574 4027 578
rect 4047 574 4051 578
rect 4159 574 4163 578
rect 4207 574 4211 578
rect 4295 574 4299 578
rect 4367 574 4371 578
rect 4431 574 4435 578
rect 4527 574 4531 578
rect 4567 574 4571 578
rect 4687 574 4691 578
rect 4703 574 4707 578
rect 4839 574 4843 578
rect 4975 574 4979 578
rect 5111 574 5115 578
rect 5663 574 5667 578
rect 1975 470 1979 474
rect 2171 470 2175 474
rect 2307 470 2311 474
rect 2315 470 2319 474
rect 2459 470 2463 474
rect 2499 470 2503 474
rect 2603 470 2607 474
rect 2683 470 2687 474
rect 2747 470 2751 474
rect 2859 470 2863 474
rect 2891 470 2895 474
rect 3035 470 3039 474
rect 3203 470 3207 474
rect 3379 470 3383 474
rect 3555 470 3559 474
rect 3799 470 3803 474
rect 111 462 115 466
rect 131 462 135 466
rect 195 462 199 466
rect 379 462 383 466
rect 427 462 431 466
rect 643 462 647 466
rect 659 462 663 466
rect 883 462 887 466
rect 907 462 911 466
rect 1099 462 1103 466
rect 1163 462 1167 466
rect 1323 462 1327 466
rect 1419 462 1423 466
rect 1547 462 1551 466
rect 1683 462 1687 466
rect 1935 462 1939 466
rect 3839 454 3843 458
rect 3931 454 3935 458
rect 4019 454 4023 458
rect 4131 454 4135 458
rect 4179 454 4183 458
rect 4331 454 4335 458
rect 4339 454 4343 458
rect 4499 454 4503 458
rect 4523 454 4527 458
rect 4659 454 4663 458
rect 4723 454 4727 458
rect 4923 454 4927 458
rect 5663 454 5667 458
rect 1975 354 1979 358
rect 2023 354 2027 358
rect 2175 354 2179 358
rect 2199 354 2203 358
rect 2343 354 2347 358
rect 2367 354 2371 358
rect 2487 354 2491 358
rect 2591 354 2595 358
rect 2631 354 2635 358
rect 2775 354 2779 358
rect 2847 354 2851 358
rect 2919 354 2923 358
rect 3063 354 3067 358
rect 3119 354 3123 358
rect 3407 354 3411 358
rect 3679 354 3683 358
rect 3799 354 3803 358
rect 111 342 115 346
rect 223 342 227 346
rect 351 342 355 346
rect 455 342 459 346
rect 575 342 579 346
rect 687 342 691 346
rect 799 342 803 346
rect 911 342 915 346
rect 1015 342 1019 346
rect 1127 342 1131 346
rect 1231 342 1235 346
rect 1351 342 1355 346
rect 1455 342 1459 346
rect 1575 342 1579 346
rect 1935 342 1939 346
rect 3839 342 3843 346
rect 3887 342 3891 346
rect 3959 342 3963 346
rect 4135 342 4139 346
rect 4159 342 4163 346
rect 4359 342 4363 346
rect 4383 342 4387 346
rect 4551 342 4555 346
rect 4615 342 4619 346
rect 4751 342 4755 346
rect 4823 342 4827 346
rect 4951 342 4955 346
rect 5015 342 5019 346
rect 5199 342 5203 346
rect 5383 342 5387 346
rect 5543 342 5547 346
rect 5663 342 5667 346
rect 1975 214 1979 218
rect 1995 214 1999 218
rect 2147 214 2151 218
rect 2171 214 2175 218
rect 2339 214 2343 218
rect 2363 214 2367 218
rect 2547 214 2551 218
rect 2563 214 2567 218
rect 2723 214 2727 218
rect 2819 214 2823 218
rect 2891 214 2895 218
rect 3051 214 3055 218
rect 3091 214 3095 218
rect 3203 214 3207 218
rect 3355 214 3359 218
rect 3379 214 3383 218
rect 3515 214 3519 218
rect 3651 214 3655 218
rect 3799 214 3803 218
rect 3839 218 3843 222
rect 3859 218 3863 222
rect 4107 218 4111 222
rect 4291 218 4295 222
rect 4355 218 4359 222
rect 4427 218 4431 222
rect 4563 218 4567 222
rect 4587 218 4591 222
rect 4699 218 4703 222
rect 4795 218 4799 222
rect 4835 218 4839 222
rect 4971 218 4975 222
rect 4987 218 4991 222
rect 5107 218 5111 222
rect 5171 218 5175 222
rect 5243 218 5247 222
rect 5355 218 5359 222
rect 5379 218 5383 222
rect 5515 218 5519 222
rect 5663 218 5667 222
rect 111 194 115 198
rect 131 194 135 198
rect 267 194 271 198
rect 323 194 327 198
rect 403 194 407 198
rect 539 194 543 198
rect 547 194 551 198
rect 675 194 679 198
rect 771 194 775 198
rect 811 194 815 198
rect 947 194 951 198
rect 987 194 991 198
rect 1083 194 1087 198
rect 1203 194 1207 198
rect 1227 194 1231 198
rect 1371 194 1375 198
rect 1427 194 1431 198
rect 1515 194 1519 198
rect 1651 194 1655 198
rect 1787 194 1791 198
rect 1935 194 1939 198
rect 1975 102 1979 106
rect 2023 102 2027 106
rect 2199 102 2203 106
rect 2391 102 2395 106
rect 2575 102 2579 106
rect 2751 102 2755 106
rect 2919 102 2923 106
rect 3079 102 3083 106
rect 3231 102 3235 106
rect 3383 102 3387 106
rect 3543 102 3547 106
rect 3679 102 3683 106
rect 3799 102 3803 106
rect 3839 106 3843 110
rect 4319 106 4323 110
rect 4455 106 4459 110
rect 4591 106 4595 110
rect 4727 106 4731 110
rect 4863 106 4867 110
rect 4999 106 5003 110
rect 5135 106 5139 110
rect 5271 106 5275 110
rect 5407 106 5411 110
rect 5543 106 5547 110
rect 5663 106 5667 110
rect 111 82 115 86
rect 159 82 163 86
rect 295 82 299 86
rect 431 82 435 86
rect 567 82 571 86
rect 703 82 707 86
rect 839 82 843 86
rect 975 82 979 86
rect 1111 82 1115 86
rect 1255 82 1259 86
rect 1399 82 1403 86
rect 1543 82 1547 86
rect 1679 82 1683 86
rect 1815 82 1819 86
rect 1935 82 1939 86
<< m4 >>
rect 84 5729 85 5735
rect 91 5734 1947 5735
rect 91 5730 111 5734
rect 115 5730 159 5734
rect 163 5730 295 5734
rect 299 5730 431 5734
rect 435 5730 567 5734
rect 571 5730 703 5734
rect 707 5730 839 5734
rect 843 5730 975 5734
rect 979 5730 1935 5734
rect 1939 5730 1947 5734
rect 91 5729 1947 5730
rect 1953 5729 1954 5735
rect 1946 5669 1947 5675
rect 1953 5674 3811 5675
rect 1953 5670 1975 5674
rect 1979 5670 2103 5674
rect 2107 5670 2239 5674
rect 2243 5670 2375 5674
rect 2379 5670 2511 5674
rect 2515 5670 2647 5674
rect 2651 5670 2783 5674
rect 2787 5670 2919 5674
rect 2923 5670 3055 5674
rect 3059 5670 3191 5674
rect 3195 5670 3327 5674
rect 3331 5670 3463 5674
rect 3467 5670 3599 5674
rect 3603 5670 3799 5674
rect 3803 5670 3811 5674
rect 1953 5669 3811 5670
rect 3817 5669 3818 5675
rect 96 5601 97 5607
rect 103 5606 1959 5607
rect 103 5602 111 5606
rect 115 5602 131 5606
rect 135 5602 267 5606
rect 271 5602 403 5606
rect 407 5602 539 5606
rect 543 5602 675 5606
rect 679 5602 755 5606
rect 759 5602 811 5606
rect 815 5602 891 5606
rect 895 5602 947 5606
rect 951 5602 1027 5606
rect 1031 5602 1163 5606
rect 1167 5602 1935 5606
rect 1939 5602 1959 5606
rect 103 5601 1959 5602
rect 1965 5601 1966 5607
rect 3822 5605 3823 5611
rect 3829 5610 5707 5611
rect 3829 5606 3839 5610
rect 3843 5606 4243 5610
rect 4247 5606 4379 5610
rect 4383 5606 4515 5610
rect 4519 5606 4651 5610
rect 4655 5606 4787 5610
rect 4791 5606 4923 5610
rect 4927 5606 5059 5610
rect 5063 5606 5663 5610
rect 5667 5606 5707 5610
rect 3829 5605 5707 5606
rect 5713 5605 5714 5611
rect 1958 5557 1959 5563
rect 1965 5562 3823 5563
rect 1965 5558 1975 5562
rect 1979 5558 1995 5562
rect 1999 5558 2075 5562
rect 2079 5558 2131 5562
rect 2135 5558 2211 5562
rect 2215 5558 2267 5562
rect 2271 5558 2347 5562
rect 2351 5558 2403 5562
rect 2407 5558 2483 5562
rect 2487 5558 2555 5562
rect 2559 5558 2619 5562
rect 2623 5558 2707 5562
rect 2711 5558 2755 5562
rect 2759 5558 2859 5562
rect 2863 5558 2891 5562
rect 2895 5558 3011 5562
rect 3015 5558 3027 5562
rect 3031 5558 3163 5562
rect 3167 5558 3299 5562
rect 3303 5558 3323 5562
rect 3327 5558 3435 5562
rect 3439 5558 3483 5562
rect 3487 5558 3571 5562
rect 3575 5558 3799 5562
rect 3803 5558 3823 5562
rect 1965 5557 3823 5558
rect 3829 5557 3830 5563
rect 3810 5493 3811 5499
rect 3817 5498 5695 5499
rect 3817 5494 3839 5498
rect 3843 5494 4271 5498
rect 4275 5494 4407 5498
rect 4411 5494 4455 5498
rect 4459 5494 4543 5498
rect 4547 5494 4591 5498
rect 4595 5494 4679 5498
rect 4683 5494 4727 5498
rect 4731 5494 4815 5498
rect 4819 5494 4863 5498
rect 4867 5494 4951 5498
rect 4955 5494 5087 5498
rect 5091 5494 5663 5498
rect 5667 5494 5695 5498
rect 3817 5493 5695 5494
rect 5701 5493 5702 5499
rect 84 5477 85 5483
rect 91 5482 1947 5483
rect 91 5478 111 5482
rect 115 5478 783 5482
rect 787 5478 863 5482
rect 867 5478 919 5482
rect 923 5478 999 5482
rect 1003 5478 1055 5482
rect 1059 5478 1135 5482
rect 1139 5478 1191 5482
rect 1195 5478 1271 5482
rect 1275 5478 1407 5482
rect 1411 5478 1543 5482
rect 1547 5478 1679 5482
rect 1683 5478 1815 5482
rect 1819 5478 1935 5482
rect 1939 5478 1947 5482
rect 91 5477 1947 5478
rect 1953 5477 1954 5483
rect 1946 5433 1947 5439
rect 1953 5438 3811 5439
rect 1953 5434 1975 5438
rect 1979 5434 2023 5438
rect 2027 5434 2159 5438
rect 2163 5434 2295 5438
rect 2299 5434 2431 5438
rect 2435 5434 2583 5438
rect 2587 5434 2735 5438
rect 2739 5434 2831 5438
rect 2835 5434 2887 5438
rect 2891 5434 2967 5438
rect 2971 5434 3039 5438
rect 3043 5434 3103 5438
rect 3107 5434 3191 5438
rect 3195 5434 3239 5438
rect 3243 5434 3351 5438
rect 3355 5434 3511 5438
rect 3515 5434 3799 5438
rect 3803 5434 3811 5438
rect 1953 5433 3811 5434
rect 3817 5433 3818 5439
rect 3822 5381 3823 5387
rect 3829 5386 5707 5387
rect 3829 5382 3839 5386
rect 3843 5382 4283 5386
rect 4287 5382 4427 5386
rect 4431 5382 4483 5386
rect 4487 5382 4563 5386
rect 4567 5382 4699 5386
rect 4703 5382 4835 5386
rect 4839 5382 4931 5386
rect 4935 5382 5171 5386
rect 5175 5382 5419 5386
rect 5423 5382 5663 5386
rect 5667 5382 5707 5386
rect 3829 5381 5707 5382
rect 5713 5381 5714 5387
rect 96 5365 97 5371
rect 103 5370 1959 5371
rect 103 5366 111 5370
rect 115 5366 427 5370
rect 431 5366 563 5370
rect 567 5366 699 5370
rect 703 5366 835 5370
rect 839 5366 971 5370
rect 975 5366 1107 5370
rect 1111 5366 1243 5370
rect 1247 5366 1379 5370
rect 1383 5366 1515 5370
rect 1519 5366 1651 5370
rect 1655 5366 1787 5370
rect 1791 5366 1935 5370
rect 1939 5366 1959 5370
rect 103 5365 1959 5366
rect 1965 5365 1966 5371
rect 1958 5285 1959 5291
rect 1965 5290 3823 5291
rect 1965 5286 1975 5290
rect 1979 5286 1995 5290
rect 1999 5286 2219 5290
rect 2223 5286 2467 5290
rect 2471 5286 2715 5290
rect 2719 5286 2803 5290
rect 2807 5286 2939 5290
rect 2943 5286 2971 5290
rect 2975 5286 3075 5290
rect 3079 5286 3211 5290
rect 3215 5286 3799 5290
rect 3803 5286 3823 5290
rect 1965 5285 3823 5286
rect 3829 5285 3830 5291
rect 84 5253 85 5259
rect 91 5258 1947 5259
rect 91 5254 111 5258
rect 115 5254 455 5258
rect 459 5254 591 5258
rect 595 5254 727 5258
rect 731 5254 863 5258
rect 867 5254 999 5258
rect 1003 5254 1135 5258
rect 1139 5254 1271 5258
rect 1275 5254 1407 5258
rect 1411 5254 1543 5258
rect 1547 5254 1679 5258
rect 1683 5254 1815 5258
rect 1819 5254 1935 5258
rect 1939 5254 1947 5258
rect 91 5253 1947 5254
rect 1953 5253 1954 5259
rect 3810 5241 3811 5247
rect 3817 5246 5695 5247
rect 3817 5242 3839 5246
rect 3843 5242 3887 5246
rect 3891 5242 4023 5246
rect 4027 5242 4159 5246
rect 4163 5242 4295 5246
rect 4299 5242 4311 5246
rect 4315 5242 4431 5246
rect 4435 5242 4511 5246
rect 4515 5242 4567 5246
rect 4571 5242 4703 5246
rect 4707 5242 4727 5246
rect 4731 5242 4839 5246
rect 4843 5242 4959 5246
rect 4963 5242 4991 5246
rect 4995 5242 5151 5246
rect 5155 5242 5199 5246
rect 5203 5242 5319 5246
rect 5323 5242 5447 5246
rect 5451 5242 5495 5246
rect 5499 5242 5663 5246
rect 5667 5242 5695 5246
rect 3817 5241 5695 5242
rect 5701 5241 5702 5247
rect 1946 5169 1947 5175
rect 1953 5174 3811 5175
rect 1953 5170 1975 5174
rect 1979 5170 2023 5174
rect 2027 5170 2159 5174
rect 2163 5170 2247 5174
rect 2251 5170 2295 5174
rect 2299 5170 2431 5174
rect 2435 5170 2495 5174
rect 2499 5170 2567 5174
rect 2571 5170 2703 5174
rect 2707 5170 2743 5174
rect 2747 5170 2839 5174
rect 2843 5170 2975 5174
rect 2979 5170 2999 5174
rect 3003 5170 3111 5174
rect 3115 5170 3247 5174
rect 3251 5170 3391 5174
rect 3395 5170 3543 5174
rect 3547 5170 3679 5174
rect 3683 5170 3799 5174
rect 3803 5170 3811 5174
rect 1953 5169 3811 5170
rect 3817 5169 3818 5175
rect 96 5125 97 5131
rect 103 5130 1959 5131
rect 103 5126 111 5130
rect 115 5126 267 5130
rect 271 5126 403 5130
rect 407 5126 427 5130
rect 431 5126 539 5130
rect 543 5126 563 5130
rect 567 5126 675 5130
rect 679 5126 699 5130
rect 703 5126 811 5130
rect 815 5126 835 5130
rect 839 5126 947 5130
rect 951 5126 971 5130
rect 975 5126 1107 5130
rect 1111 5126 1243 5130
rect 1247 5126 1379 5130
rect 1383 5126 1515 5130
rect 1519 5126 1651 5130
rect 1655 5126 1787 5130
rect 1791 5126 1935 5130
rect 1939 5126 1959 5130
rect 103 5125 1959 5126
rect 1965 5125 1966 5131
rect 3822 5129 3823 5135
rect 3829 5134 5707 5135
rect 3829 5130 3839 5134
rect 3843 5130 3859 5134
rect 3863 5130 3979 5134
rect 3983 5130 3995 5134
rect 3999 5130 4131 5134
rect 4135 5130 4267 5134
rect 4271 5130 4275 5134
rect 4279 5130 4403 5134
rect 4407 5130 4539 5134
rect 4543 5130 4579 5134
rect 4583 5130 4675 5134
rect 4679 5130 4811 5134
rect 4815 5130 4883 5134
rect 4887 5130 4963 5134
rect 4967 5130 5123 5134
rect 5127 5130 5195 5134
rect 5199 5130 5291 5134
rect 5295 5130 5467 5134
rect 5471 5130 5515 5134
rect 5519 5130 5663 5134
rect 5667 5130 5707 5134
rect 3829 5129 5707 5130
rect 5713 5129 5714 5135
rect 1958 5057 1959 5063
rect 1965 5062 3823 5063
rect 1965 5058 1975 5062
rect 1979 5058 1995 5062
rect 1999 5058 2131 5062
rect 2135 5058 2267 5062
rect 2271 5058 2403 5062
rect 2407 5058 2539 5062
rect 2543 5058 2675 5062
rect 2679 5058 2811 5062
rect 2815 5058 2947 5062
rect 2951 5058 3083 5062
rect 3087 5058 3107 5062
rect 3111 5058 3219 5062
rect 3223 5058 3243 5062
rect 3247 5058 3363 5062
rect 3367 5058 3379 5062
rect 3383 5058 3515 5062
rect 3519 5058 3651 5062
rect 3655 5058 3799 5062
rect 3803 5058 3823 5062
rect 1965 5057 3823 5058
rect 3829 5057 3830 5063
rect 84 5001 85 5007
rect 91 5006 1947 5007
rect 91 5002 111 5006
rect 115 5002 159 5006
rect 163 5002 295 5006
rect 299 5002 431 5006
rect 435 5002 567 5006
rect 571 5002 703 5006
rect 707 5002 839 5006
rect 843 5002 975 5006
rect 979 5002 1935 5006
rect 1939 5002 1947 5006
rect 91 5001 1947 5002
rect 1953 5001 1954 5007
rect 3810 5001 3811 5007
rect 3817 5006 5695 5007
rect 3817 5002 3839 5006
rect 3843 5002 4007 5006
rect 4011 5002 4303 5006
rect 4307 5002 4607 5006
rect 4611 5002 4863 5006
rect 4867 5002 4911 5006
rect 4915 5002 4999 5006
rect 5003 5002 5135 5006
rect 5139 5002 5223 5006
rect 5227 5002 5271 5006
rect 5275 5002 5407 5006
rect 5411 5002 5543 5006
rect 5547 5002 5663 5006
rect 5667 5002 5695 5006
rect 3817 5001 5695 5002
rect 5701 5001 5702 5007
rect 1946 4937 1947 4943
rect 1953 4942 3811 4943
rect 1953 4938 1975 4942
rect 1979 4938 3135 4942
rect 3139 4938 3271 4942
rect 3275 4938 3407 4942
rect 3411 4938 3543 4942
rect 3547 4938 3679 4942
rect 3683 4938 3799 4942
rect 3803 4938 3811 4942
rect 1953 4937 3811 4938
rect 3817 4937 3818 4943
rect 96 4881 97 4887
rect 103 4886 1959 4887
rect 103 4882 111 4886
rect 115 4882 131 4886
rect 135 4882 267 4886
rect 271 4882 403 4886
rect 407 4882 539 4886
rect 543 4882 675 4886
rect 679 4882 1935 4886
rect 1939 4882 1959 4886
rect 103 4881 1959 4882
rect 1965 4881 1966 4887
rect 3822 4877 3823 4883
rect 3829 4882 5707 4883
rect 3829 4878 3839 4882
rect 3843 4878 4483 4882
rect 4487 4878 4675 4882
rect 4679 4878 4835 4882
rect 4839 4878 4875 4882
rect 4879 4878 4971 4882
rect 4975 4878 5091 4882
rect 5095 4878 5107 4882
rect 5111 4878 5243 4882
rect 5247 4878 5315 4882
rect 5319 4878 5379 4882
rect 5383 4878 5515 4882
rect 5519 4878 5663 4882
rect 5667 4878 5707 4882
rect 3829 4877 5707 4878
rect 5713 4877 5714 4883
rect 1958 4797 1959 4803
rect 1965 4802 3823 4803
rect 1965 4798 1975 4802
rect 1979 4798 3107 4802
rect 3111 4798 3243 4802
rect 3247 4798 3379 4802
rect 3383 4798 3515 4802
rect 3519 4798 3651 4802
rect 3655 4798 3799 4802
rect 3803 4798 3823 4802
rect 1965 4797 3823 4798
rect 3829 4797 3830 4803
rect 84 4765 85 4771
rect 91 4770 1947 4771
rect 91 4766 111 4770
rect 115 4766 159 4770
rect 163 4766 295 4770
rect 299 4766 431 4770
rect 435 4766 567 4770
rect 571 4766 703 4770
rect 707 4766 1935 4770
rect 1939 4766 1947 4770
rect 91 4765 1947 4766
rect 1953 4765 1954 4771
rect 3810 4745 3811 4751
rect 3817 4750 5695 4751
rect 3817 4746 3839 4750
rect 3843 4746 4119 4750
rect 4123 4746 4375 4750
rect 4379 4746 4511 4750
rect 4515 4746 4647 4750
rect 4651 4746 4703 4750
rect 4707 4746 4903 4750
rect 4907 4746 4943 4750
rect 4947 4746 5119 4750
rect 5123 4746 5255 4750
rect 5259 4746 5343 4750
rect 5347 4746 5543 4750
rect 5547 4746 5663 4750
rect 5667 4746 5695 4750
rect 3817 4745 5695 4746
rect 5701 4745 5702 4751
rect 1946 4655 1947 4661
rect 1953 4655 1978 4661
rect 1972 4651 1978 4655
rect 96 4645 97 4651
rect 103 4650 1959 4651
rect 103 4646 111 4650
rect 115 4646 131 4650
rect 135 4646 211 4650
rect 215 4646 267 4650
rect 271 4646 403 4650
rect 407 4646 427 4650
rect 431 4646 539 4650
rect 543 4646 667 4650
rect 671 4646 675 4650
rect 679 4646 931 4650
rect 935 4646 1219 4650
rect 1223 4646 1515 4650
rect 1519 4646 1787 4650
rect 1791 4646 1935 4650
rect 1939 4646 1959 4650
rect 103 4645 1959 4646
rect 1965 4645 1966 4651
rect 1972 4650 3811 4651
rect 1972 4646 1975 4650
rect 1979 4646 2023 4650
rect 2027 4646 2159 4650
rect 2163 4646 2311 4650
rect 2315 4646 2479 4650
rect 2483 4646 2655 4650
rect 2659 4646 2831 4650
rect 2835 4646 3007 4650
rect 3011 4646 3135 4650
rect 3139 4646 3183 4650
rect 3187 4646 3271 4650
rect 3275 4646 3351 4650
rect 3355 4646 3407 4650
rect 3411 4646 3527 4650
rect 3531 4646 3543 4650
rect 3547 4646 3679 4650
rect 3683 4646 3799 4650
rect 3803 4646 3811 4650
rect 1972 4645 3811 4646
rect 3817 4645 3818 4651
rect 3822 4613 3823 4619
rect 3829 4618 5707 4619
rect 3829 4614 3839 4618
rect 3843 4614 4035 4618
rect 4039 4614 4091 4618
rect 4095 4614 4331 4618
rect 4335 4614 4347 4618
rect 4351 4614 4619 4618
rect 4623 4614 4627 4618
rect 4631 4614 4915 4618
rect 4919 4614 4931 4618
rect 4935 4614 5227 4618
rect 5231 4614 5235 4618
rect 5239 4614 5515 4618
rect 5519 4614 5663 4618
rect 5667 4614 5707 4618
rect 3829 4613 5707 4614
rect 5713 4613 5714 4619
rect 84 4533 85 4539
rect 91 4538 1947 4539
rect 91 4534 111 4538
rect 115 4534 239 4538
rect 243 4534 447 4538
rect 451 4534 455 4538
rect 459 4534 623 4538
rect 627 4534 695 4538
rect 699 4534 807 4538
rect 811 4534 959 4538
rect 963 4534 999 4538
rect 1003 4534 1199 4538
rect 1203 4534 1247 4538
rect 1251 4534 1407 4538
rect 1411 4534 1543 4538
rect 1547 4534 1623 4538
rect 1627 4534 1815 4538
rect 1819 4534 1935 4538
rect 1939 4534 1947 4538
rect 91 4533 1947 4534
rect 1953 4533 1954 4539
rect 1958 4533 1959 4539
rect 1965 4538 3823 4539
rect 1965 4534 1975 4538
rect 1979 4534 1995 4538
rect 1999 4534 2131 4538
rect 2135 4534 2227 4538
rect 2231 4534 2283 4538
rect 2287 4534 2451 4538
rect 2455 4534 2459 4538
rect 2463 4534 2627 4538
rect 2631 4534 2691 4538
rect 2695 4534 2803 4538
rect 2807 4534 2915 4538
rect 2919 4534 2979 4538
rect 2983 4534 3131 4538
rect 3135 4534 3155 4538
rect 3159 4534 3323 4538
rect 3327 4534 3355 4538
rect 3359 4534 3499 4538
rect 3503 4534 3579 4538
rect 3583 4534 3651 4538
rect 3655 4534 3799 4538
rect 3803 4534 3823 4538
rect 1965 4533 3823 4534
rect 3829 4533 3830 4539
rect 3810 4485 3811 4491
rect 3817 4490 5695 4491
rect 3817 4486 3839 4490
rect 3843 4486 4063 4490
rect 4067 4486 4311 4490
rect 4315 4486 4359 4490
rect 4363 4486 4535 4490
rect 4539 4486 4655 4490
rect 4659 4486 4775 4490
rect 4779 4486 4959 4490
rect 4963 4486 5023 4490
rect 5027 4486 5263 4490
rect 5267 4486 5279 4490
rect 5283 4486 5543 4490
rect 5547 4486 5663 4490
rect 5667 4486 5695 4490
rect 3817 4485 5695 4486
rect 5701 4485 5702 4491
rect 1946 4427 1947 4433
rect 1953 4427 1978 4433
rect 1972 4423 1978 4427
rect 96 4417 97 4423
rect 103 4422 1959 4423
rect 103 4418 111 4422
rect 115 4418 419 4422
rect 423 4418 571 4422
rect 575 4418 595 4422
rect 599 4418 739 4422
rect 743 4418 779 4422
rect 783 4418 915 4422
rect 919 4418 971 4422
rect 975 4418 1107 4422
rect 1111 4418 1171 4422
rect 1175 4418 1299 4422
rect 1303 4418 1379 4422
rect 1383 4418 1499 4422
rect 1503 4418 1595 4422
rect 1599 4418 1707 4422
rect 1711 4418 1787 4422
rect 1791 4418 1935 4422
rect 1939 4418 1959 4422
rect 103 4417 1959 4418
rect 1965 4417 1966 4423
rect 1972 4422 3811 4423
rect 1972 4418 1975 4422
rect 1979 4418 2023 4422
rect 2027 4418 2119 4422
rect 2123 4418 2255 4422
rect 2259 4418 2343 4422
rect 2347 4418 2487 4422
rect 2491 4418 2567 4422
rect 2571 4418 2719 4422
rect 2723 4418 2783 4422
rect 2787 4418 2943 4422
rect 2947 4418 2991 4422
rect 2995 4418 3159 4422
rect 3163 4418 3199 4422
rect 3203 4418 3383 4422
rect 3387 4418 3407 4422
rect 3411 4418 3607 4422
rect 3611 4418 3799 4422
rect 3803 4418 3811 4422
rect 1972 4417 3811 4418
rect 3817 4417 3818 4423
rect 3822 4353 3823 4359
rect 3829 4358 5707 4359
rect 3829 4354 3839 4358
rect 3843 4354 4283 4358
rect 4287 4354 4507 4358
rect 4511 4354 4515 4358
rect 4519 4354 4691 4358
rect 4695 4354 4747 4358
rect 4751 4354 4875 4358
rect 4879 4354 4995 4358
rect 4999 4354 5067 4358
rect 5071 4354 5251 4358
rect 5255 4354 5267 4358
rect 5271 4354 5467 4358
rect 5471 4354 5515 4358
rect 5519 4354 5663 4358
rect 5667 4354 5707 4358
rect 3829 4353 5707 4354
rect 5713 4353 5714 4359
rect 84 4305 85 4311
rect 91 4310 1947 4311
rect 91 4306 111 4310
rect 115 4306 599 4310
rect 603 4306 655 4310
rect 659 4306 767 4310
rect 771 4306 823 4310
rect 827 4306 943 4310
rect 947 4306 991 4310
rect 995 4306 1135 4310
rect 1139 4306 1167 4310
rect 1171 4306 1327 4310
rect 1331 4306 1343 4310
rect 1347 4306 1519 4310
rect 1523 4306 1527 4310
rect 1531 4306 1703 4310
rect 1707 4306 1735 4310
rect 1739 4306 1935 4310
rect 1939 4306 1947 4310
rect 91 4305 1947 4306
rect 1953 4305 1954 4311
rect 1958 4297 1959 4303
rect 1965 4302 3823 4303
rect 1965 4298 1975 4302
rect 1979 4298 2019 4302
rect 2023 4298 2091 4302
rect 2095 4298 2243 4302
rect 2247 4298 2315 4302
rect 2319 4298 2459 4302
rect 2463 4298 2539 4302
rect 2543 4298 2667 4302
rect 2671 4298 2755 4302
rect 2759 4298 2875 4302
rect 2879 4298 2963 4302
rect 2967 4298 3083 4302
rect 3087 4298 3171 4302
rect 3175 4298 3291 4302
rect 3295 4298 3379 4302
rect 3383 4298 3799 4302
rect 3803 4298 3823 4302
rect 1965 4297 3823 4298
rect 3829 4297 3830 4303
rect 3810 4221 3811 4227
rect 3817 4226 5695 4227
rect 3817 4222 3839 4226
rect 3843 4222 4543 4226
rect 4547 4222 4719 4226
rect 4723 4222 4815 4226
rect 4819 4222 4903 4226
rect 4907 4222 4951 4226
rect 4955 4222 5087 4226
rect 5091 4222 5095 4226
rect 5099 4222 5223 4226
rect 5227 4222 5295 4226
rect 5299 4222 5359 4226
rect 5363 4222 5495 4226
rect 5499 4222 5663 4226
rect 5667 4222 5695 4226
rect 3817 4221 5695 4222
rect 5701 4221 5702 4227
rect 1946 4191 1947 4197
rect 1953 4191 1978 4197
rect 1972 4187 1978 4191
rect 96 4181 97 4187
rect 103 4186 1959 4187
rect 103 4182 111 4186
rect 115 4182 347 4186
rect 351 4182 515 4186
rect 519 4182 627 4186
rect 631 4182 699 4186
rect 703 4182 795 4186
rect 799 4182 891 4186
rect 895 4182 963 4186
rect 967 4182 1099 4186
rect 1103 4182 1139 4186
rect 1143 4182 1315 4186
rect 1319 4182 1491 4186
rect 1495 4182 1531 4186
rect 1535 4182 1675 4186
rect 1679 4182 1935 4186
rect 1939 4182 1959 4186
rect 103 4181 1959 4182
rect 1965 4181 1966 4187
rect 1972 4186 3811 4187
rect 1972 4182 1975 4186
rect 1979 4182 2023 4186
rect 2027 4182 2047 4186
rect 2051 4182 2271 4186
rect 2275 4182 2287 4186
rect 2291 4182 2487 4186
rect 2491 4182 2551 4186
rect 2555 4182 2695 4186
rect 2699 4182 2799 4186
rect 2803 4182 2903 4186
rect 2907 4182 3039 4186
rect 3043 4182 3111 4186
rect 3115 4182 3279 4186
rect 3283 4182 3319 4186
rect 3323 4182 3519 4186
rect 3523 4182 3799 4186
rect 3803 4182 3811 4186
rect 1972 4181 3811 4182
rect 3817 4181 3818 4187
rect 3822 4105 3823 4111
rect 3829 4110 5707 4111
rect 3829 4106 3839 4110
rect 3843 4106 4787 4110
rect 4791 4106 4923 4110
rect 4927 4106 4939 4110
rect 4943 4106 5059 4110
rect 5063 4106 5075 4110
rect 5079 4106 5195 4110
rect 5199 4106 5211 4110
rect 5215 4106 5331 4110
rect 5335 4106 5347 4110
rect 5351 4106 5467 4110
rect 5471 4106 5483 4110
rect 5487 4106 5663 4110
rect 5667 4106 5707 4110
rect 3829 4105 5707 4106
rect 5713 4105 5714 4111
rect 1958 4069 1959 4075
rect 1965 4074 3823 4075
rect 1965 4070 1975 4074
rect 1979 4070 1995 4074
rect 1999 4070 2259 4074
rect 2263 4070 2283 4074
rect 2287 4070 2523 4074
rect 2527 4070 2587 4074
rect 2591 4070 2771 4074
rect 2775 4070 2875 4074
rect 2879 4070 3011 4074
rect 3015 4070 3163 4074
rect 3167 4070 3251 4074
rect 3255 4070 3451 4074
rect 3455 4070 3491 4074
rect 3495 4070 3799 4074
rect 3803 4070 3823 4074
rect 1965 4069 3823 4070
rect 3829 4069 3830 4075
rect 84 4053 85 4059
rect 91 4058 1947 4059
rect 91 4054 111 4058
rect 115 4054 231 4058
rect 235 4054 375 4058
rect 379 4054 423 4058
rect 427 4054 543 4058
rect 547 4054 615 4058
rect 619 4054 727 4058
rect 731 4054 807 4058
rect 811 4054 919 4058
rect 923 4054 991 4058
rect 995 4054 1127 4058
rect 1131 4054 1167 4058
rect 1171 4054 1335 4058
rect 1339 4054 1343 4058
rect 1347 4054 1503 4058
rect 1507 4054 1559 4058
rect 1563 4054 1671 4058
rect 1675 4054 1815 4058
rect 1819 4054 1935 4058
rect 1939 4054 1947 4058
rect 91 4053 1947 4054
rect 1953 4053 1954 4059
rect 3810 3985 3811 3991
rect 3817 3990 5695 3991
rect 3817 3986 3839 3990
rect 3843 3986 4831 3990
rect 4835 3986 4967 3990
rect 4971 3986 5103 3990
rect 5107 3986 5111 3990
rect 5115 3986 5239 3990
rect 5243 3986 5255 3990
rect 5259 3986 5375 3990
rect 5379 3986 5407 3990
rect 5411 3986 5511 3990
rect 5515 3986 5543 3990
rect 5547 3986 5663 3990
rect 5667 3986 5695 3990
rect 3817 3985 5695 3986
rect 5701 3985 5702 3991
rect 1946 3951 1947 3957
rect 1953 3951 1978 3957
rect 96 3941 97 3947
rect 103 3946 1959 3947
rect 103 3942 111 3946
rect 115 3942 203 3946
rect 207 3942 251 3946
rect 255 3942 395 3946
rect 399 3942 451 3946
rect 455 3942 587 3946
rect 591 3942 643 3946
rect 647 3942 779 3946
rect 783 3942 827 3946
rect 831 3942 963 3946
rect 967 3942 1003 3946
rect 1007 3942 1139 3946
rect 1143 3942 1171 3946
rect 1175 3942 1307 3946
rect 1311 3942 1331 3946
rect 1335 3942 1475 3946
rect 1479 3942 1491 3946
rect 1495 3942 1643 3946
rect 1647 3942 1651 3946
rect 1655 3942 1787 3946
rect 1791 3942 1935 3946
rect 1939 3942 1959 3946
rect 103 3941 1959 3942
rect 1965 3941 1966 3947
rect 1972 3943 1978 3951
rect 1972 3942 3811 3943
rect 1972 3938 1975 3942
rect 1979 3938 2023 3942
rect 2027 3938 2311 3942
rect 2315 3938 2615 3942
rect 2619 3938 2671 3942
rect 2675 3938 2807 3942
rect 2811 3938 2903 3942
rect 2907 3938 2943 3942
rect 2947 3938 3079 3942
rect 3083 3938 3191 3942
rect 3195 3938 3215 3942
rect 3219 3938 3479 3942
rect 3483 3938 3799 3942
rect 3803 3938 3811 3942
rect 1972 3937 3811 3938
rect 3817 3937 3818 3943
rect 3822 3853 3823 3859
rect 3829 3858 5707 3859
rect 3829 3854 3839 3858
rect 3843 3854 4499 3858
rect 4503 3854 4675 3858
rect 4679 3854 4803 3858
rect 4807 3854 4875 3858
rect 4879 3854 4939 3858
rect 4943 3854 5083 3858
rect 5087 3854 5091 3858
rect 5095 3854 5227 3858
rect 5231 3854 5315 3858
rect 5319 3854 5379 3858
rect 5383 3854 5515 3858
rect 5519 3854 5663 3858
rect 5667 3854 5707 3858
rect 3829 3853 5707 3854
rect 5713 3853 5714 3859
rect 84 3829 85 3835
rect 91 3834 1947 3835
rect 91 3830 111 3834
rect 115 3830 279 3834
rect 283 3830 311 3834
rect 315 3830 479 3834
rect 483 3830 511 3834
rect 515 3830 671 3834
rect 675 3830 735 3834
rect 739 3830 855 3834
rect 859 3830 991 3834
rect 995 3830 1031 3834
rect 1035 3830 1199 3834
rect 1203 3830 1263 3834
rect 1267 3830 1359 3834
rect 1363 3830 1519 3834
rect 1523 3830 1551 3834
rect 1555 3830 1679 3834
rect 1683 3830 1815 3834
rect 1819 3830 1935 3834
rect 1939 3830 1947 3834
rect 91 3829 1947 3830
rect 1953 3829 1954 3835
rect 1958 3813 1959 3819
rect 1965 3818 3823 3819
rect 1965 3814 1975 3818
rect 1979 3814 1995 3818
rect 1999 3814 2131 3818
rect 2135 3814 2283 3818
rect 2287 3814 2443 3818
rect 2447 3814 2603 3818
rect 2607 3814 2643 3818
rect 2647 3814 2763 3818
rect 2767 3814 2779 3818
rect 2783 3814 2915 3818
rect 2919 3814 2923 3818
rect 2927 3814 3051 3818
rect 3055 3814 3083 3818
rect 3087 3814 3187 3818
rect 3191 3814 3243 3818
rect 3247 3814 3411 3818
rect 3415 3814 3799 3818
rect 3803 3814 3823 3818
rect 1965 3813 3823 3814
rect 3829 3813 3830 3819
rect 3810 3717 3811 3723
rect 3817 3722 5695 3723
rect 3817 3718 3839 3722
rect 3843 3718 4271 3722
rect 4275 3718 4471 3722
rect 4475 3718 4527 3722
rect 4531 3718 4695 3722
rect 4699 3718 4703 3722
rect 4707 3718 4903 3722
rect 4907 3718 4935 3722
rect 4939 3718 5119 3722
rect 5123 3718 5191 3722
rect 5195 3718 5343 3722
rect 5347 3718 5447 3722
rect 5451 3718 5543 3722
rect 5547 3718 5663 3722
rect 5667 3718 5695 3722
rect 3817 3717 5695 3718
rect 5701 3717 5702 3723
rect 1946 3703 1947 3709
rect 1953 3703 1978 3709
rect 1972 3699 1978 3703
rect 96 3693 97 3699
rect 103 3698 1959 3699
rect 103 3694 111 3698
rect 115 3694 155 3698
rect 159 3694 283 3698
rect 287 3694 291 3698
rect 295 3694 427 3698
rect 431 3694 483 3698
rect 487 3694 563 3698
rect 567 3694 699 3698
rect 703 3694 707 3698
rect 711 3694 835 3698
rect 839 3694 963 3698
rect 967 3694 971 3698
rect 975 3694 1107 3698
rect 1111 3694 1235 3698
rect 1239 3694 1243 3698
rect 1247 3694 1379 3698
rect 1383 3694 1515 3698
rect 1519 3694 1523 3698
rect 1527 3694 1787 3698
rect 1791 3694 1935 3698
rect 1939 3694 1959 3698
rect 103 3693 1959 3694
rect 1965 3693 1966 3699
rect 1972 3698 3811 3699
rect 1972 3694 1975 3698
rect 1979 3694 2023 3698
rect 2027 3694 2047 3698
rect 2051 3694 2159 3698
rect 2163 3694 2223 3698
rect 2227 3694 2311 3698
rect 2315 3694 2407 3698
rect 2411 3694 2471 3698
rect 2475 3694 2591 3698
rect 2595 3694 2631 3698
rect 2635 3694 2783 3698
rect 2787 3694 2791 3698
rect 2795 3694 2951 3698
rect 2955 3694 2967 3698
rect 2971 3694 3111 3698
rect 3115 3694 3151 3698
rect 3155 3694 3271 3698
rect 3275 3694 3335 3698
rect 3339 3694 3439 3698
rect 3443 3694 3519 3698
rect 3523 3694 3679 3698
rect 3683 3694 3799 3698
rect 3803 3694 3811 3698
rect 1972 3693 3811 3694
rect 3817 3693 3818 3699
rect 3822 3601 3823 3607
rect 3829 3606 5707 3607
rect 3829 3602 3839 3606
rect 3843 3602 3859 3606
rect 3863 3602 3995 3606
rect 3999 3602 4131 3606
rect 4135 3602 4243 3606
rect 4247 3602 4267 3606
rect 4271 3602 4403 3606
rect 4407 3602 4443 3606
rect 4447 3602 4539 3606
rect 4543 3602 4667 3606
rect 4671 3602 4675 3606
rect 4679 3602 4811 3606
rect 4815 3602 4907 3606
rect 4911 3602 4947 3606
rect 4951 3602 5163 3606
rect 5167 3602 5419 3606
rect 5423 3602 5663 3606
rect 5667 3602 5707 3606
rect 3829 3601 5707 3602
rect 5713 3601 5714 3607
rect 1958 3569 1959 3575
rect 1965 3574 3823 3575
rect 1965 3570 1975 3574
rect 1979 3570 2019 3574
rect 2023 3570 2195 3574
rect 2199 3570 2307 3574
rect 2311 3570 2379 3574
rect 2383 3570 2443 3574
rect 2447 3570 2563 3574
rect 2567 3570 2579 3574
rect 2583 3570 2715 3574
rect 2719 3570 2755 3574
rect 2759 3570 2939 3574
rect 2943 3570 3123 3574
rect 3127 3570 3307 3574
rect 3311 3570 3491 3574
rect 3495 3570 3651 3574
rect 3655 3570 3799 3574
rect 3803 3570 3823 3574
rect 1965 3569 3823 3570
rect 3829 3569 3830 3575
rect 3810 3489 3811 3495
rect 3817 3494 5695 3495
rect 3817 3490 3839 3494
rect 3843 3490 3887 3494
rect 3891 3490 4023 3494
rect 4027 3490 4159 3494
rect 4163 3490 4295 3494
rect 4299 3490 4431 3494
rect 4435 3490 4567 3494
rect 4571 3490 4703 3494
rect 4707 3490 4839 3494
rect 4843 3490 4975 3494
rect 4979 3490 5111 3494
rect 5115 3490 5247 3494
rect 5251 3490 5383 3494
rect 5387 3490 5519 3494
rect 5523 3490 5663 3494
rect 5667 3490 5695 3494
rect 3817 3489 5695 3490
rect 5701 3489 5702 3495
rect 1946 3421 1947 3427
rect 1953 3426 3811 3427
rect 1953 3422 1975 3426
rect 1979 3422 2167 3426
rect 2171 3422 2303 3426
rect 2307 3422 2335 3426
rect 2339 3422 2439 3426
rect 2443 3422 2471 3426
rect 2475 3422 2575 3426
rect 2579 3422 2607 3426
rect 2611 3422 2711 3426
rect 2715 3422 2743 3426
rect 2747 3422 2847 3426
rect 2851 3422 2983 3426
rect 2987 3422 3799 3426
rect 3803 3422 3811 3426
rect 1953 3421 3811 3422
rect 3817 3421 3818 3427
rect 3822 3369 3823 3375
rect 3829 3374 5707 3375
rect 3829 3370 3839 3374
rect 3843 3370 3859 3374
rect 3863 3370 3995 3374
rect 3999 3370 4131 3374
rect 4135 3370 4155 3374
rect 4159 3370 4267 3374
rect 4271 3370 4315 3374
rect 4319 3370 4403 3374
rect 4407 3370 4467 3374
rect 4471 3370 4539 3374
rect 4543 3370 4627 3374
rect 4631 3370 4675 3374
rect 4679 3370 4787 3374
rect 4791 3370 4811 3374
rect 4815 3370 4947 3374
rect 4951 3370 5083 3374
rect 5087 3370 5219 3374
rect 5223 3370 5355 3374
rect 5359 3370 5491 3374
rect 5495 3370 5663 3374
rect 5667 3370 5707 3374
rect 3829 3369 5707 3370
rect 5713 3369 5714 3375
rect 1958 3309 1959 3315
rect 1965 3314 3823 3315
rect 1965 3310 1975 3314
rect 1979 3310 2059 3314
rect 2063 3310 2139 3314
rect 2143 3310 2203 3314
rect 2207 3310 2275 3314
rect 2279 3310 2363 3314
rect 2367 3310 2411 3314
rect 2415 3310 2539 3314
rect 2543 3310 2547 3314
rect 2551 3310 2683 3314
rect 2687 3310 2739 3314
rect 2743 3310 2819 3314
rect 2823 3310 2955 3314
rect 2959 3310 3187 3314
rect 3191 3310 3427 3314
rect 3431 3310 3651 3314
rect 3655 3310 3799 3314
rect 3803 3310 3823 3314
rect 1965 3309 3823 3310
rect 3829 3309 3830 3315
rect 84 3293 85 3299
rect 91 3298 1947 3299
rect 91 3294 111 3298
rect 115 3294 159 3298
rect 163 3294 183 3298
rect 187 3294 295 3298
rect 299 3294 319 3298
rect 323 3294 431 3298
rect 435 3294 455 3298
rect 459 3294 567 3298
rect 571 3294 591 3298
rect 595 3294 703 3298
rect 707 3294 727 3298
rect 731 3294 839 3298
rect 843 3294 863 3298
rect 867 3294 975 3298
rect 979 3294 999 3298
rect 1003 3294 1111 3298
rect 1115 3294 1135 3298
rect 1139 3294 1247 3298
rect 1251 3294 1271 3298
rect 1275 3294 1383 3298
rect 1387 3294 1407 3298
rect 1411 3294 1519 3298
rect 1523 3294 1543 3298
rect 1547 3294 1935 3298
rect 1939 3294 1947 3298
rect 91 3293 1947 3294
rect 1953 3293 1954 3299
rect 3810 3245 3811 3251
rect 3817 3250 5695 3251
rect 3817 3246 3839 3250
rect 3843 3246 3887 3250
rect 3891 3246 4023 3250
rect 4027 3246 4183 3250
rect 4187 3246 4343 3250
rect 4347 3246 4495 3250
rect 4499 3246 4655 3250
rect 4659 3246 4807 3250
rect 4811 3246 4815 3250
rect 4819 3246 4943 3250
rect 4947 3246 4975 3250
rect 4979 3246 5079 3250
rect 5083 3246 5215 3250
rect 5219 3246 5351 3250
rect 5355 3246 5663 3250
rect 5667 3246 5695 3250
rect 3817 3245 5695 3246
rect 5701 3245 5702 3251
rect 1946 3193 1947 3199
rect 1953 3198 3811 3199
rect 1953 3194 1975 3198
rect 1979 3194 2023 3198
rect 2027 3194 2087 3198
rect 2091 3194 2159 3198
rect 2163 3194 2231 3198
rect 2235 3194 2303 3198
rect 2307 3194 2391 3198
rect 2395 3194 2455 3198
rect 2459 3194 2567 3198
rect 2571 3194 2615 3198
rect 2619 3194 2767 3198
rect 2771 3194 2783 3198
rect 2787 3194 2951 3198
rect 2955 3194 2983 3198
rect 2987 3194 3127 3198
rect 3131 3194 3215 3198
rect 3219 3194 3311 3198
rect 3315 3194 3455 3198
rect 3459 3194 3503 3198
rect 3507 3194 3679 3198
rect 3683 3194 3799 3198
rect 3803 3194 3811 3198
rect 1953 3193 3811 3194
rect 3817 3193 3818 3199
rect 96 3153 97 3159
rect 103 3158 1959 3159
rect 103 3154 111 3158
rect 115 3154 131 3158
rect 135 3154 267 3158
rect 271 3154 291 3158
rect 295 3154 403 3158
rect 407 3154 459 3158
rect 463 3154 539 3158
rect 543 3154 627 3158
rect 631 3154 675 3158
rect 679 3154 811 3158
rect 815 3154 947 3158
rect 951 3154 995 3158
rect 999 3154 1083 3158
rect 1087 3154 1187 3158
rect 1191 3154 1219 3158
rect 1223 3154 1355 3158
rect 1359 3154 1387 3158
rect 1391 3154 1491 3158
rect 1495 3154 1595 3158
rect 1599 3154 1787 3158
rect 1791 3154 1935 3158
rect 1939 3154 1959 3158
rect 103 3153 1959 3154
rect 1965 3153 1966 3159
rect 3822 3129 3823 3135
rect 3829 3134 5707 3135
rect 3829 3130 3839 3134
rect 3843 3130 4699 3134
rect 4703 3130 4779 3134
rect 4783 3130 4835 3134
rect 4839 3130 4915 3134
rect 4919 3130 4971 3134
rect 4975 3130 5051 3134
rect 5055 3130 5107 3134
rect 5111 3130 5187 3134
rect 5191 3130 5243 3134
rect 5247 3130 5323 3134
rect 5327 3130 5379 3134
rect 5383 3130 5515 3134
rect 5519 3130 5663 3134
rect 5667 3130 5707 3134
rect 3829 3129 5707 3130
rect 5713 3129 5714 3135
rect 1958 3061 1959 3067
rect 1965 3066 3823 3067
rect 1965 3062 1975 3066
rect 1979 3062 1995 3066
rect 1999 3062 2131 3066
rect 2135 3062 2275 3066
rect 2279 3062 2427 3066
rect 2431 3062 2587 3066
rect 2591 3062 2755 3066
rect 2759 3062 2811 3066
rect 2815 3062 2923 3066
rect 2927 3062 3003 3066
rect 3007 3062 3099 3066
rect 3103 3062 3203 3066
rect 3207 3062 3283 3066
rect 3287 3062 3403 3066
rect 3407 3062 3475 3066
rect 3479 3062 3603 3066
rect 3607 3062 3651 3066
rect 3655 3062 3799 3066
rect 3803 3062 3823 3066
rect 1965 3061 3823 3062
rect 3829 3061 3830 3067
rect 84 3041 85 3047
rect 91 3046 1947 3047
rect 91 3042 111 3046
rect 115 3042 319 3046
rect 323 3042 327 3046
rect 331 3042 487 3046
rect 491 3042 647 3046
rect 651 3042 655 3046
rect 659 3042 807 3046
rect 811 3042 839 3046
rect 843 3042 959 3046
rect 963 3042 1023 3046
rect 1027 3042 1103 3046
rect 1107 3042 1215 3046
rect 1219 3042 1247 3046
rect 1251 3042 1391 3046
rect 1395 3042 1415 3046
rect 1419 3042 1535 3046
rect 1539 3042 1623 3046
rect 1627 3042 1679 3046
rect 1683 3042 1815 3046
rect 1819 3042 1935 3046
rect 1939 3042 1947 3046
rect 91 3041 1947 3042
rect 1953 3041 1954 3047
rect 3810 3017 3811 3023
rect 3817 3022 5695 3023
rect 3817 3018 3839 3022
rect 3843 3018 4367 3022
rect 4371 3018 4567 3022
rect 4571 3018 4727 3022
rect 4731 3018 4783 3022
rect 4787 3018 4863 3022
rect 4867 3018 4999 3022
rect 5003 3018 5023 3022
rect 5027 3018 5135 3022
rect 5139 3018 5271 3022
rect 5275 3018 5279 3022
rect 5283 3018 5407 3022
rect 5411 3018 5535 3022
rect 5539 3018 5543 3022
rect 5547 3018 5663 3022
rect 5667 3018 5695 3022
rect 3817 3017 5695 3018
rect 5701 3017 5702 3023
rect 1946 2941 1947 2947
rect 1953 2946 3811 2947
rect 1953 2942 1975 2946
rect 1979 2942 2839 2946
rect 2843 2942 2847 2946
rect 2851 2942 2983 2946
rect 2987 2942 3031 2946
rect 3035 2942 3119 2946
rect 3123 2942 3231 2946
rect 3235 2942 3255 2946
rect 3259 2942 3391 2946
rect 3395 2942 3431 2946
rect 3435 2942 3527 2946
rect 3531 2942 3631 2946
rect 3635 2942 3671 2946
rect 3675 2942 3799 2946
rect 3803 2942 3811 2946
rect 1953 2941 3811 2942
rect 3817 2941 3818 2947
rect 96 2929 97 2935
rect 103 2934 1959 2935
rect 103 2930 111 2934
rect 115 2930 155 2934
rect 159 2930 299 2934
rect 303 2930 379 2934
rect 383 2930 459 2934
rect 463 2930 595 2934
rect 599 2930 619 2934
rect 623 2930 779 2934
rect 783 2930 811 2934
rect 815 2930 931 2934
rect 935 2930 1019 2934
rect 1023 2930 1075 2934
rect 1079 2930 1219 2934
rect 1223 2930 1363 2934
rect 1367 2930 1411 2934
rect 1415 2930 1507 2934
rect 1511 2930 1611 2934
rect 1615 2930 1651 2934
rect 1655 2930 1787 2934
rect 1791 2930 1935 2934
rect 1939 2930 1959 2934
rect 103 2929 1959 2930
rect 1965 2929 1966 2935
rect 3822 2905 3823 2911
rect 3829 2910 5707 2911
rect 3829 2906 3839 2910
rect 3843 2906 4035 2910
rect 4039 2906 4315 2910
rect 4319 2906 4339 2910
rect 4343 2906 4539 2910
rect 4543 2906 4603 2910
rect 4607 2906 4755 2910
rect 4759 2906 4907 2910
rect 4911 2906 4995 2910
rect 4999 2906 5219 2910
rect 5223 2906 5251 2910
rect 5255 2906 5507 2910
rect 5511 2906 5515 2910
rect 5519 2906 5663 2910
rect 5667 2906 5707 2910
rect 3829 2905 5707 2906
rect 5713 2905 5714 2911
rect 1958 2829 1959 2835
rect 1965 2834 3823 2835
rect 1965 2830 1975 2834
rect 1979 2830 2011 2834
rect 2015 2830 2251 2834
rect 2255 2830 2491 2834
rect 2495 2830 2731 2834
rect 2735 2830 2819 2834
rect 2823 2830 2955 2834
rect 2959 2830 2971 2834
rect 2975 2830 3091 2834
rect 3095 2830 3227 2834
rect 3231 2830 3363 2834
rect 3367 2830 3499 2834
rect 3503 2830 3643 2834
rect 3647 2830 3799 2834
rect 3803 2830 3823 2834
rect 1965 2829 3823 2830
rect 3829 2829 3830 2835
rect 84 2785 85 2791
rect 91 2790 1947 2791
rect 91 2786 111 2790
rect 115 2786 183 2790
rect 187 2786 287 2790
rect 291 2786 407 2790
rect 411 2786 423 2790
rect 427 2786 559 2790
rect 563 2786 623 2790
rect 627 2786 695 2790
rect 699 2786 831 2790
rect 835 2786 839 2790
rect 843 2786 1047 2790
rect 1051 2786 1247 2790
rect 1251 2786 1439 2790
rect 1443 2786 1639 2790
rect 1643 2786 1815 2790
rect 1819 2786 1935 2790
rect 1939 2786 1947 2790
rect 91 2785 1947 2786
rect 1953 2785 1954 2791
rect 3810 2785 3811 2791
rect 3817 2790 5695 2791
rect 3817 2786 3839 2790
rect 3843 2786 3967 2790
rect 3971 2786 4063 2790
rect 4067 2786 4255 2790
rect 4259 2786 4343 2790
rect 4347 2786 4567 2790
rect 4571 2786 4631 2790
rect 4635 2786 4895 2790
rect 4899 2786 4935 2790
rect 4939 2786 5231 2790
rect 5235 2786 5247 2790
rect 5251 2786 5543 2790
rect 5547 2786 5663 2790
rect 5667 2786 5695 2790
rect 3817 2785 5695 2786
rect 5701 2785 5702 2791
rect 1946 2717 1947 2723
rect 1953 2722 3811 2723
rect 1953 2718 1975 2722
rect 1979 2718 2023 2722
rect 2027 2718 2039 2722
rect 2043 2718 2159 2722
rect 2163 2718 2279 2722
rect 2283 2718 2295 2722
rect 2299 2718 2431 2722
rect 2435 2718 2519 2722
rect 2523 2718 2567 2722
rect 2571 2718 2703 2722
rect 2707 2718 2759 2722
rect 2763 2718 2839 2722
rect 2843 2718 2975 2722
rect 2979 2718 2999 2722
rect 3003 2718 3111 2722
rect 3115 2718 3247 2722
rect 3251 2718 3383 2722
rect 3387 2718 3799 2722
rect 3803 2718 3811 2722
rect 1953 2717 3811 2718
rect 3817 2717 3818 2723
rect 3822 2669 3823 2675
rect 3829 2674 5707 2675
rect 3829 2670 3839 2674
rect 3843 2670 3939 2674
rect 3943 2670 4027 2674
rect 4031 2670 4227 2674
rect 4231 2670 4275 2674
rect 4279 2670 4539 2674
rect 4543 2670 4555 2674
rect 4559 2670 4867 2674
rect 4871 2670 5203 2674
rect 5207 2670 5515 2674
rect 5519 2670 5663 2674
rect 5667 2670 5707 2674
rect 3829 2669 5707 2670
rect 5713 2669 5714 2675
rect 96 2653 97 2659
rect 103 2658 1959 2659
rect 103 2654 111 2658
rect 115 2654 259 2658
rect 263 2654 395 2658
rect 399 2654 531 2658
rect 535 2654 539 2658
rect 543 2654 667 2658
rect 671 2654 699 2658
rect 703 2654 803 2658
rect 807 2654 883 2658
rect 887 2654 1091 2658
rect 1095 2654 1323 2658
rect 1327 2654 1563 2658
rect 1567 2654 1787 2658
rect 1791 2654 1935 2658
rect 1939 2654 1959 2658
rect 103 2653 1959 2654
rect 1965 2653 1966 2659
rect 1958 2605 1959 2611
rect 1965 2610 3823 2611
rect 1965 2606 1975 2610
rect 1979 2606 1995 2610
rect 1999 2606 2131 2610
rect 2135 2606 2203 2610
rect 2207 2606 2267 2610
rect 2271 2606 2403 2610
rect 2407 2606 2419 2610
rect 2423 2606 2539 2610
rect 2543 2606 2627 2610
rect 2631 2606 2675 2610
rect 2679 2606 2811 2610
rect 2815 2606 2827 2610
rect 2831 2606 2947 2610
rect 2951 2606 3019 2610
rect 3023 2606 3083 2610
rect 3087 2606 3211 2610
rect 3215 2606 3219 2610
rect 3223 2606 3355 2610
rect 3359 2606 3403 2610
rect 3407 2606 3799 2610
rect 3803 2606 3823 2610
rect 1965 2605 3823 2606
rect 3829 2605 3830 2611
rect 3810 2553 3811 2559
rect 3817 2558 5695 2559
rect 3817 2554 3839 2558
rect 3843 2554 4055 2558
rect 4059 2554 4303 2558
rect 4307 2554 4335 2558
rect 4339 2554 4559 2558
rect 4563 2554 4583 2558
rect 4587 2554 4799 2558
rect 4803 2554 4895 2558
rect 4899 2554 5047 2558
rect 5051 2554 5231 2558
rect 5235 2554 5303 2558
rect 5307 2554 5543 2558
rect 5547 2554 5663 2558
rect 5667 2554 5695 2558
rect 3817 2553 5695 2554
rect 5701 2553 5702 2559
rect 84 2529 85 2535
rect 91 2534 1947 2535
rect 91 2530 111 2534
rect 115 2530 567 2534
rect 571 2530 695 2534
rect 699 2530 727 2534
rect 731 2530 847 2534
rect 851 2530 911 2534
rect 915 2530 999 2534
rect 1003 2530 1119 2534
rect 1123 2530 1159 2534
rect 1163 2530 1327 2534
rect 1331 2530 1351 2534
rect 1355 2530 1495 2534
rect 1499 2530 1591 2534
rect 1595 2530 1663 2534
rect 1667 2530 1815 2534
rect 1819 2530 1935 2534
rect 1939 2530 1947 2534
rect 91 2529 1947 2530
rect 1953 2529 1954 2535
rect 1946 2485 1947 2491
rect 1953 2490 3811 2491
rect 1953 2486 1975 2490
rect 1979 2486 2023 2490
rect 2027 2486 2231 2490
rect 2235 2486 2319 2490
rect 2323 2486 2447 2490
rect 2451 2486 2567 2490
rect 2571 2486 2655 2490
rect 2659 2486 2799 2490
rect 2803 2486 2855 2490
rect 2859 2486 3023 2490
rect 3027 2486 3047 2490
rect 3051 2486 3239 2490
rect 3243 2486 3431 2490
rect 3435 2486 3455 2490
rect 3459 2486 3671 2490
rect 3675 2486 3799 2490
rect 3803 2486 3811 2490
rect 1953 2485 3811 2486
rect 3817 2485 3818 2491
rect 3822 2425 3823 2431
rect 3829 2430 5707 2431
rect 3829 2426 3839 2430
rect 3843 2426 4307 2430
rect 4311 2426 4491 2430
rect 4495 2426 4531 2430
rect 4535 2426 4635 2430
rect 4639 2426 4771 2430
rect 4775 2426 4795 2430
rect 4799 2426 4963 2430
rect 4967 2426 5019 2430
rect 5023 2426 5139 2430
rect 5143 2426 5275 2430
rect 5279 2426 5323 2430
rect 5327 2426 5515 2430
rect 5519 2426 5663 2430
rect 5667 2426 5707 2430
rect 3829 2425 5707 2426
rect 5713 2425 5714 2431
rect 96 2409 97 2415
rect 103 2414 1959 2415
rect 103 2410 111 2414
rect 115 2410 355 2414
rect 359 2410 507 2414
rect 511 2410 667 2414
rect 671 2410 675 2414
rect 679 2410 819 2414
rect 823 2410 859 2414
rect 863 2410 971 2414
rect 975 2410 1059 2414
rect 1063 2410 1131 2414
rect 1135 2410 1267 2414
rect 1271 2410 1299 2414
rect 1303 2410 1467 2414
rect 1471 2410 1483 2414
rect 1487 2410 1635 2414
rect 1639 2410 1699 2414
rect 1703 2410 1787 2414
rect 1791 2410 1935 2414
rect 1939 2410 1959 2414
rect 103 2409 1959 2410
rect 1965 2409 1966 2415
rect 1958 2365 1959 2371
rect 1965 2370 3823 2371
rect 1965 2366 1975 2370
rect 1979 2366 2291 2370
rect 2295 2366 2331 2370
rect 2335 2366 2539 2370
rect 2543 2366 2739 2370
rect 2743 2366 2771 2370
rect 2775 2366 2931 2370
rect 2935 2366 2995 2370
rect 2999 2366 3123 2370
rect 3127 2366 3211 2370
rect 3215 2366 3307 2370
rect 3311 2366 3427 2370
rect 3431 2366 3491 2370
rect 3495 2366 3643 2370
rect 3647 2366 3651 2370
rect 3655 2366 3799 2370
rect 3803 2366 3823 2370
rect 1965 2365 3823 2366
rect 3829 2365 3830 2371
rect 84 2289 85 2295
rect 91 2294 1947 2295
rect 91 2290 111 2294
rect 115 2290 159 2294
rect 163 2290 335 2294
rect 339 2290 383 2294
rect 387 2290 535 2294
rect 539 2290 543 2294
rect 547 2290 703 2294
rect 707 2290 759 2294
rect 763 2290 887 2294
rect 891 2290 975 2294
rect 979 2290 1087 2294
rect 1091 2290 1199 2294
rect 1203 2290 1295 2294
rect 1299 2290 1431 2294
rect 1435 2290 1511 2294
rect 1515 2290 1671 2294
rect 1675 2290 1727 2294
rect 1731 2290 1935 2294
rect 1939 2290 1947 2294
rect 91 2289 1947 2290
rect 1953 2289 1954 2295
rect 3810 2293 3811 2299
rect 3817 2298 5695 2299
rect 3817 2294 3839 2298
rect 3843 2294 3887 2298
rect 3891 2294 4071 2298
rect 4075 2294 4271 2298
rect 4275 2294 4463 2298
rect 4467 2294 4519 2298
rect 4523 2294 4655 2298
rect 4659 2294 4663 2298
rect 4667 2294 4823 2298
rect 4827 2294 4839 2298
rect 4843 2294 4991 2298
rect 4995 2294 5015 2298
rect 5019 2294 5167 2298
rect 5171 2294 5183 2298
rect 5187 2294 5351 2298
rect 5355 2294 5359 2298
rect 5363 2294 5535 2298
rect 5539 2294 5543 2298
rect 5547 2294 5663 2298
rect 5667 2294 5695 2298
rect 3817 2293 5695 2294
rect 5701 2293 5702 2299
rect 1946 2225 1947 2231
rect 1953 2230 3811 2231
rect 1953 2226 1975 2230
rect 1979 2226 2359 2230
rect 2363 2226 2463 2230
rect 2467 2226 2567 2230
rect 2571 2226 2599 2230
rect 2603 2226 2735 2230
rect 2739 2226 2767 2230
rect 2771 2226 2959 2230
rect 2963 2226 3151 2230
rect 3155 2226 3335 2230
rect 3339 2226 3519 2230
rect 3523 2226 3679 2230
rect 3683 2226 3799 2230
rect 3803 2226 3811 2230
rect 1953 2225 3811 2226
rect 3817 2225 3818 2231
rect 3822 2181 3823 2187
rect 3829 2186 5707 2187
rect 3829 2182 3839 2186
rect 3843 2182 3859 2186
rect 3863 2182 4043 2186
rect 4047 2182 4243 2186
rect 4247 2182 4251 2186
rect 4255 2182 4435 2186
rect 4439 2182 4459 2186
rect 4463 2182 4627 2186
rect 4631 2182 4659 2186
rect 4663 2182 4811 2186
rect 4815 2182 4851 2186
rect 4855 2182 4987 2186
rect 4991 2182 5035 2186
rect 5039 2182 5155 2186
rect 5159 2182 5219 2186
rect 5223 2182 5331 2186
rect 5335 2182 5411 2186
rect 5415 2182 5507 2186
rect 5511 2182 5663 2186
rect 5667 2182 5707 2186
rect 3829 2181 5707 2182
rect 5713 2181 5714 2187
rect 96 2157 97 2163
rect 103 2162 1959 2163
rect 103 2158 111 2162
rect 115 2158 131 2162
rect 135 2158 299 2162
rect 303 2158 307 2162
rect 311 2158 499 2162
rect 503 2158 515 2162
rect 519 2158 715 2162
rect 719 2158 731 2162
rect 735 2158 931 2162
rect 935 2158 947 2162
rect 951 2158 1155 2162
rect 1159 2158 1171 2162
rect 1175 2158 1387 2162
rect 1391 2158 1403 2162
rect 1407 2158 1627 2162
rect 1631 2158 1643 2162
rect 1647 2158 1935 2162
rect 1939 2158 1959 2162
rect 103 2157 1959 2158
rect 1965 2157 1966 2163
rect 1958 2081 1959 2087
rect 1965 2086 3823 2087
rect 1965 2082 1975 2086
rect 1979 2082 2419 2086
rect 2423 2082 2435 2086
rect 2439 2082 2571 2086
rect 2575 2082 2611 2086
rect 2615 2082 2707 2086
rect 2711 2082 2795 2086
rect 2799 2082 2979 2086
rect 2983 2082 3155 2086
rect 3159 2082 3323 2086
rect 3327 2082 3499 2086
rect 3503 2082 3651 2086
rect 3655 2082 3799 2086
rect 3803 2082 3823 2086
rect 1965 2081 3823 2082
rect 3829 2081 3830 2087
rect 3810 2049 3811 2055
rect 3817 2054 5695 2055
rect 3817 2050 3839 2054
rect 3843 2050 3887 2054
rect 3891 2050 4071 2054
rect 4075 2050 4279 2054
rect 4283 2050 4287 2054
rect 4291 2050 4423 2054
rect 4427 2050 4487 2054
rect 4491 2050 4559 2054
rect 4563 2050 4687 2054
rect 4691 2050 4695 2054
rect 4699 2050 4839 2054
rect 4843 2050 4879 2054
rect 4883 2050 5063 2054
rect 5067 2050 5247 2054
rect 5251 2050 5439 2054
rect 5443 2050 5663 2054
rect 5667 2050 5695 2054
rect 3817 2049 5695 2050
rect 5701 2049 5702 2055
rect 84 2037 85 2043
rect 91 2042 1947 2043
rect 91 2038 111 2042
rect 115 2038 159 2042
rect 163 2038 327 2042
rect 331 2038 343 2042
rect 347 2038 527 2042
rect 531 2038 567 2042
rect 571 2038 743 2042
rect 747 2038 807 2042
rect 811 2038 959 2042
rect 963 2038 1063 2042
rect 1067 2038 1183 2042
rect 1187 2038 1335 2042
rect 1339 2038 1415 2042
rect 1419 2038 1607 2042
rect 1611 2038 1655 2042
rect 1659 2038 1935 2042
rect 1939 2038 1947 2042
rect 91 2037 1947 2038
rect 1953 2037 1954 2043
rect 1946 1957 1947 1963
rect 1953 1962 3811 1963
rect 1953 1958 1975 1962
rect 1979 1958 2359 1962
rect 2363 1958 2447 1962
rect 2451 1958 2495 1962
rect 2499 1958 2631 1962
rect 2635 1958 2639 1962
rect 2643 1958 2767 1962
rect 2771 1958 2823 1962
rect 2827 1958 2903 1962
rect 2907 1958 3007 1962
rect 3011 1958 3039 1962
rect 3043 1958 3175 1962
rect 3179 1958 3183 1962
rect 3187 1958 3319 1962
rect 3323 1958 3351 1962
rect 3355 1958 3527 1962
rect 3531 1958 3679 1962
rect 3683 1958 3799 1962
rect 3803 1958 3811 1962
rect 1953 1957 3811 1958
rect 3817 1957 3818 1963
rect 96 1921 97 1927
rect 103 1926 1959 1927
rect 103 1922 111 1926
rect 115 1922 131 1926
rect 135 1922 315 1926
rect 319 1922 331 1926
rect 335 1922 499 1926
rect 503 1922 539 1926
rect 543 1922 667 1926
rect 671 1922 779 1926
rect 783 1922 843 1926
rect 847 1922 1027 1926
rect 1031 1922 1035 1926
rect 1039 1922 1219 1926
rect 1223 1922 1307 1926
rect 1311 1922 1411 1926
rect 1415 1922 1579 1926
rect 1583 1922 1603 1926
rect 1607 1922 1935 1926
rect 1939 1922 1959 1926
rect 103 1921 1959 1922
rect 1965 1921 1966 1927
rect 3822 1917 3823 1923
rect 3829 1922 5707 1923
rect 3829 1918 3839 1922
rect 3843 1918 3955 1922
rect 3959 1918 4195 1922
rect 4199 1918 4259 1922
rect 4263 1918 4395 1922
rect 4399 1918 4467 1922
rect 4471 1918 4531 1922
rect 4535 1918 4667 1922
rect 4671 1918 4771 1922
rect 4775 1918 4811 1922
rect 4815 1918 5091 1922
rect 5095 1918 5411 1922
rect 5415 1918 5663 1922
rect 5667 1918 5707 1922
rect 3829 1917 5707 1918
rect 5713 1917 5714 1923
rect 1958 1845 1959 1851
rect 1965 1850 3823 1851
rect 1965 1846 1975 1850
rect 1979 1846 2211 1850
rect 2215 1846 2331 1850
rect 2335 1846 2355 1850
rect 2359 1846 2467 1850
rect 2471 1846 2499 1850
rect 2503 1846 2603 1850
rect 2607 1846 2643 1850
rect 2647 1846 2739 1850
rect 2743 1846 2787 1850
rect 2791 1846 2875 1850
rect 2879 1846 2931 1850
rect 2935 1846 3011 1850
rect 3015 1846 3083 1850
rect 3087 1846 3147 1850
rect 3151 1846 3291 1850
rect 3295 1846 3799 1850
rect 3803 1846 3823 1850
rect 1965 1845 3823 1846
rect 3829 1845 3830 1851
rect 3810 1805 3811 1811
rect 3817 1810 5695 1811
rect 3817 1806 3839 1810
rect 3843 1806 3983 1810
rect 3987 1806 4223 1810
rect 4227 1806 4367 1810
rect 4371 1806 4495 1810
rect 4499 1806 4575 1810
rect 4579 1806 4783 1810
rect 4787 1806 4799 1810
rect 4803 1806 4983 1810
rect 4987 1806 5119 1810
rect 5123 1806 5175 1810
rect 5179 1806 5367 1810
rect 5371 1806 5439 1810
rect 5443 1806 5543 1810
rect 5547 1806 5663 1810
rect 5667 1806 5695 1810
rect 3817 1805 5695 1806
rect 5701 1805 5702 1811
rect 84 1797 85 1803
rect 91 1802 1947 1803
rect 91 1798 111 1802
rect 115 1798 359 1802
rect 363 1798 527 1802
rect 531 1798 535 1802
rect 539 1798 695 1802
rect 699 1798 855 1802
rect 859 1798 871 1802
rect 875 1798 1015 1802
rect 1019 1798 1055 1802
rect 1059 1798 1183 1802
rect 1187 1798 1247 1802
rect 1251 1798 1351 1802
rect 1355 1798 1439 1802
rect 1443 1798 1519 1802
rect 1523 1798 1631 1802
rect 1635 1798 1935 1802
rect 1939 1798 1947 1802
rect 91 1797 1947 1798
rect 1953 1797 1954 1803
rect 1946 1733 1947 1739
rect 1953 1738 3811 1739
rect 1953 1734 1975 1738
rect 1979 1734 2023 1738
rect 2027 1734 2215 1738
rect 2219 1734 2239 1738
rect 2243 1734 2383 1738
rect 2387 1734 2407 1738
rect 2411 1734 2527 1738
rect 2531 1734 2599 1738
rect 2603 1734 2671 1738
rect 2675 1734 2791 1738
rect 2795 1734 2815 1738
rect 2819 1734 2959 1738
rect 2963 1734 2975 1738
rect 2979 1734 3111 1738
rect 3115 1734 3151 1738
rect 3155 1734 3335 1738
rect 3339 1734 3519 1738
rect 3523 1734 3799 1738
rect 3803 1734 3811 1738
rect 1953 1733 3811 1734
rect 3817 1733 3818 1739
rect 3822 1677 3823 1683
rect 3829 1682 5707 1683
rect 3829 1678 3839 1682
rect 3843 1678 4339 1682
rect 4343 1678 4547 1682
rect 4551 1678 4603 1682
rect 4607 1678 4755 1682
rect 4759 1678 4787 1682
rect 4791 1678 4955 1682
rect 4959 1678 4971 1682
rect 4975 1678 5147 1682
rect 5151 1678 5155 1682
rect 5159 1678 5339 1682
rect 5343 1678 5515 1682
rect 5519 1678 5663 1682
rect 5667 1678 5707 1682
rect 3829 1677 5707 1678
rect 5713 1677 5714 1683
rect 96 1669 97 1675
rect 103 1674 1959 1675
rect 103 1670 111 1674
rect 115 1670 427 1674
rect 431 1670 507 1674
rect 511 1670 611 1674
rect 615 1670 667 1674
rect 671 1670 803 1674
rect 807 1670 827 1674
rect 831 1670 987 1674
rect 991 1670 995 1674
rect 999 1670 1155 1674
rect 1159 1670 1187 1674
rect 1191 1670 1323 1674
rect 1327 1670 1379 1674
rect 1383 1670 1491 1674
rect 1495 1670 1935 1674
rect 1939 1670 1959 1674
rect 103 1669 1959 1670
rect 1965 1669 1966 1675
rect 1958 1621 1959 1627
rect 1965 1626 3823 1627
rect 1965 1622 1975 1626
rect 1979 1622 1995 1626
rect 1999 1622 2163 1626
rect 2167 1622 2187 1626
rect 2191 1622 2371 1626
rect 2375 1622 2379 1626
rect 2383 1622 2571 1626
rect 2575 1622 2587 1626
rect 2591 1622 2763 1626
rect 2767 1622 2803 1626
rect 2807 1622 2947 1626
rect 2951 1622 3019 1626
rect 3023 1622 3123 1626
rect 3127 1622 3235 1626
rect 3239 1622 3307 1626
rect 3311 1622 3451 1626
rect 3455 1622 3491 1626
rect 3495 1622 3651 1626
rect 3655 1622 3799 1626
rect 3803 1622 3823 1626
rect 1965 1621 3823 1622
rect 3829 1621 3830 1627
rect 84 1549 85 1555
rect 91 1554 1947 1555
rect 91 1550 111 1554
rect 115 1550 359 1554
rect 363 1550 455 1554
rect 459 1550 631 1554
rect 635 1550 639 1554
rect 643 1550 831 1554
rect 835 1550 887 1554
rect 891 1550 1023 1554
rect 1027 1550 1135 1554
rect 1139 1550 1215 1554
rect 1219 1550 1367 1554
rect 1371 1550 1407 1554
rect 1411 1550 1599 1554
rect 1603 1550 1815 1554
rect 1819 1550 1935 1554
rect 1939 1550 1947 1554
rect 91 1549 1947 1550
rect 1953 1549 1954 1555
rect 3810 1549 3811 1555
rect 3817 1554 5695 1555
rect 3817 1550 3839 1554
rect 3843 1550 3887 1554
rect 3891 1550 4031 1554
rect 4035 1550 4199 1554
rect 4203 1550 4367 1554
rect 4371 1550 4527 1554
rect 4531 1550 4631 1554
rect 4635 1550 4695 1554
rect 4699 1550 4815 1554
rect 4819 1550 4863 1554
rect 4867 1550 4999 1554
rect 5003 1550 5031 1554
rect 5035 1550 5183 1554
rect 5187 1550 5207 1554
rect 5211 1550 5367 1554
rect 5371 1550 5383 1554
rect 5387 1550 5543 1554
rect 5547 1550 5663 1554
rect 5667 1550 5695 1554
rect 3817 1549 5695 1550
rect 5701 1549 5702 1555
rect 96 1437 97 1443
rect 103 1442 1959 1443
rect 103 1438 111 1442
rect 115 1438 131 1442
rect 135 1438 307 1442
rect 311 1438 331 1442
rect 335 1438 499 1442
rect 503 1438 603 1442
rect 607 1438 683 1442
rect 687 1438 859 1442
rect 863 1438 1027 1442
rect 1031 1438 1107 1442
rect 1111 1438 1187 1442
rect 1191 1438 1339 1442
rect 1343 1438 1491 1442
rect 1495 1438 1571 1442
rect 1575 1438 1651 1442
rect 1655 1438 1787 1442
rect 1791 1438 1935 1442
rect 1939 1438 1959 1442
rect 103 1437 1959 1438
rect 1965 1437 1966 1443
rect 3822 1433 3823 1439
rect 3829 1438 5707 1439
rect 3829 1434 3839 1438
rect 3843 1434 3859 1438
rect 3863 1434 4003 1438
rect 4007 1434 4171 1438
rect 4175 1434 4179 1438
rect 4183 1434 4339 1438
rect 4343 1434 4355 1438
rect 4359 1434 4499 1438
rect 4503 1434 4531 1438
rect 4535 1434 4667 1438
rect 4671 1434 4707 1438
rect 4711 1434 4835 1438
rect 4839 1434 4875 1438
rect 4879 1434 5003 1438
rect 5007 1434 5043 1438
rect 5047 1434 5179 1438
rect 5183 1434 5203 1438
rect 5207 1434 5355 1438
rect 5359 1434 5371 1438
rect 5375 1434 5515 1438
rect 5519 1434 5663 1438
rect 5667 1434 5707 1438
rect 3829 1433 5707 1434
rect 5713 1433 5714 1439
rect 84 1317 85 1323
rect 91 1322 1947 1323
rect 91 1318 111 1322
rect 115 1318 159 1322
rect 163 1318 335 1322
rect 339 1318 375 1322
rect 379 1318 527 1322
rect 531 1318 599 1322
rect 603 1318 711 1322
rect 715 1318 807 1322
rect 811 1318 887 1322
rect 891 1318 999 1322
rect 1003 1318 1055 1322
rect 1059 1318 1175 1322
rect 1179 1318 1215 1322
rect 1219 1318 1343 1322
rect 1347 1318 1367 1322
rect 1371 1318 1511 1322
rect 1515 1318 1519 1322
rect 1523 1318 1671 1322
rect 1675 1318 1679 1322
rect 1683 1318 1815 1322
rect 1819 1318 1935 1322
rect 1939 1318 1947 1322
rect 91 1317 1947 1318
rect 1953 1317 1954 1323
rect 3810 1321 3811 1327
rect 3817 1326 5695 1327
rect 3817 1322 3839 1326
rect 3843 1322 3887 1326
rect 3891 1322 4031 1326
rect 4035 1322 4175 1326
rect 4179 1322 4207 1326
rect 4211 1322 4383 1326
rect 4387 1322 4471 1326
rect 4475 1322 4559 1326
rect 4563 1322 4735 1326
rect 4739 1322 4751 1326
rect 4755 1322 4903 1326
rect 4907 1322 5023 1326
rect 5027 1322 5071 1326
rect 5075 1322 5231 1326
rect 5235 1322 5287 1326
rect 5291 1322 5399 1326
rect 5403 1322 5543 1326
rect 5547 1322 5663 1326
rect 5667 1322 5695 1326
rect 3817 1321 5695 1322
rect 5701 1321 5702 1327
rect 1946 1305 1947 1311
rect 1953 1310 3811 1311
rect 1953 1306 1975 1310
rect 1979 1306 2023 1310
rect 2027 1306 2191 1310
rect 2195 1306 2399 1310
rect 2403 1306 2615 1310
rect 2619 1306 2831 1310
rect 2835 1306 3047 1310
rect 3051 1306 3263 1310
rect 3267 1306 3271 1310
rect 3275 1306 3407 1310
rect 3411 1306 3479 1310
rect 3483 1306 3543 1310
rect 3547 1306 3679 1310
rect 3683 1306 3799 1310
rect 3803 1306 3811 1310
rect 1953 1305 3811 1306
rect 3817 1305 3818 1311
rect 96 1205 97 1211
rect 103 1210 1959 1211
rect 103 1206 111 1210
rect 115 1206 131 1210
rect 135 1206 347 1210
rect 351 1206 563 1210
rect 567 1206 571 1210
rect 575 1206 779 1210
rect 783 1206 971 1210
rect 975 1206 987 1210
rect 991 1206 1147 1210
rect 1151 1206 1195 1210
rect 1199 1206 1315 1210
rect 1319 1206 1395 1210
rect 1399 1206 1483 1210
rect 1487 1206 1603 1210
rect 1607 1206 1643 1210
rect 1647 1206 1787 1210
rect 1791 1206 1935 1210
rect 1939 1206 1959 1210
rect 103 1205 1959 1206
rect 1965 1205 1966 1211
rect 3822 1197 3823 1203
rect 3829 1202 5707 1203
rect 3829 1198 3839 1202
rect 3843 1198 3859 1202
rect 3863 1198 4147 1202
rect 4151 1198 4427 1202
rect 4431 1198 4443 1202
rect 4447 1198 4563 1202
rect 4567 1198 4699 1202
rect 4703 1198 4723 1202
rect 4727 1198 4835 1202
rect 4839 1198 4971 1202
rect 4975 1198 4995 1202
rect 4999 1198 5107 1202
rect 5111 1198 5243 1202
rect 5247 1198 5259 1202
rect 5263 1198 5379 1202
rect 5383 1198 5515 1202
rect 5519 1198 5663 1202
rect 5667 1198 5707 1202
rect 3829 1197 5707 1198
rect 5713 1197 5714 1203
rect 1958 1181 1959 1187
rect 1965 1186 3823 1187
rect 1965 1182 1975 1186
rect 1979 1182 1995 1186
rect 1999 1182 2227 1186
rect 2231 1182 2467 1186
rect 2471 1182 2691 1186
rect 2695 1182 2907 1186
rect 2911 1182 3107 1186
rect 3111 1182 3243 1186
rect 3247 1182 3299 1186
rect 3303 1182 3379 1186
rect 3383 1182 3483 1186
rect 3487 1182 3515 1186
rect 3519 1182 3651 1186
rect 3655 1182 3799 1186
rect 3803 1182 3823 1186
rect 1965 1181 3823 1182
rect 3829 1181 3830 1187
rect 84 1069 85 1075
rect 91 1074 1947 1075
rect 91 1070 111 1074
rect 115 1070 159 1074
rect 163 1070 375 1074
rect 379 1070 471 1074
rect 475 1070 591 1074
rect 595 1070 607 1074
rect 611 1070 743 1074
rect 747 1070 807 1074
rect 811 1070 887 1074
rect 891 1070 1015 1074
rect 1019 1070 1031 1074
rect 1035 1070 1223 1074
rect 1227 1070 1423 1074
rect 1427 1070 1631 1074
rect 1635 1070 1815 1074
rect 1819 1070 1935 1074
rect 1939 1070 1947 1074
rect 91 1069 1947 1070
rect 1953 1074 5702 1075
rect 1953 1070 1975 1074
rect 1979 1070 2023 1074
rect 2027 1070 2183 1074
rect 2187 1070 2255 1074
rect 2259 1070 2319 1074
rect 2323 1070 2455 1074
rect 2459 1070 2495 1074
rect 2499 1070 2599 1074
rect 2603 1070 2719 1074
rect 2723 1070 2743 1074
rect 2747 1070 2887 1074
rect 2891 1070 2935 1074
rect 2939 1070 3031 1074
rect 3035 1070 3135 1074
rect 3139 1070 3175 1074
rect 3179 1070 3319 1074
rect 3323 1070 3327 1074
rect 3331 1070 3463 1074
rect 3467 1070 3511 1074
rect 3515 1070 3679 1074
rect 3683 1070 3799 1074
rect 3803 1070 3839 1074
rect 3843 1070 4367 1074
rect 4371 1070 4455 1074
rect 4459 1070 4503 1074
rect 4507 1070 4591 1074
rect 4595 1070 4639 1074
rect 4643 1070 4727 1074
rect 4731 1070 4775 1074
rect 4779 1070 4863 1074
rect 4867 1070 4911 1074
rect 4915 1070 4999 1074
rect 5003 1070 5135 1074
rect 5139 1070 5271 1074
rect 5275 1070 5407 1074
rect 5411 1070 5543 1074
rect 5547 1070 5663 1074
rect 5667 1070 5702 1074
rect 1953 1069 5702 1070
rect 96 945 97 951
rect 103 950 1959 951
rect 103 946 111 950
rect 115 946 259 950
rect 263 946 395 950
rect 399 946 443 950
rect 447 946 531 950
rect 535 946 579 950
rect 583 946 667 950
rect 671 946 715 950
rect 719 946 803 950
rect 807 946 859 950
rect 863 946 939 950
rect 943 946 1003 950
rect 1007 946 1935 950
rect 1939 946 1959 950
rect 103 945 1959 946
rect 1965 950 5714 951
rect 1965 946 1975 950
rect 1979 946 1995 950
rect 1999 946 2131 950
rect 2135 946 2155 950
rect 2159 946 2267 950
rect 2271 946 2291 950
rect 2295 946 2403 950
rect 2407 946 2427 950
rect 2431 946 2539 950
rect 2543 946 2571 950
rect 2575 946 2675 950
rect 2679 946 2715 950
rect 2719 946 2811 950
rect 2815 946 2859 950
rect 2863 946 2947 950
rect 2951 946 3003 950
rect 3007 946 3083 950
rect 3087 946 3147 950
rect 3151 946 3219 950
rect 3223 946 3291 950
rect 3295 946 3355 950
rect 3359 946 3435 950
rect 3439 946 3491 950
rect 3495 946 3799 950
rect 3803 946 3839 950
rect 3843 946 4019 950
rect 4023 946 4155 950
rect 4159 946 4291 950
rect 4295 946 4339 950
rect 4343 946 4427 950
rect 4431 946 4475 950
rect 4479 946 4563 950
rect 4567 946 4611 950
rect 4615 946 4699 950
rect 4703 946 4747 950
rect 4751 946 4883 950
rect 4887 946 5663 950
rect 5667 946 5714 950
rect 1965 945 5714 946
rect 1946 833 1947 839
rect 1953 838 3811 839
rect 1953 834 1975 838
rect 1979 834 2023 838
rect 2027 834 2159 838
rect 2163 834 2167 838
rect 2171 834 2295 838
rect 2299 834 2335 838
rect 2339 834 2431 838
rect 2435 834 2495 838
rect 2499 834 2567 838
rect 2571 834 2655 838
rect 2659 834 2703 838
rect 2707 834 2823 838
rect 2827 834 2839 838
rect 2843 834 2975 838
rect 2979 834 2991 838
rect 2995 834 3111 838
rect 3115 834 3247 838
rect 3251 834 3383 838
rect 3387 834 3519 838
rect 3523 834 3799 838
rect 3803 834 3811 838
rect 1953 833 3811 834
rect 3817 833 3818 839
rect 84 821 85 827
rect 91 826 1947 827
rect 91 822 111 826
rect 115 822 239 826
rect 243 822 287 826
rect 291 822 423 826
rect 427 822 439 826
rect 443 822 559 826
rect 563 822 647 826
rect 651 822 695 826
rect 699 822 831 826
rect 835 822 855 826
rect 859 822 967 826
rect 971 822 1063 826
rect 1067 822 1935 826
rect 1939 822 1947 826
rect 91 821 1947 822
rect 1953 821 1954 827
rect 3810 817 3811 823
rect 3817 822 5695 823
rect 3817 818 3839 822
rect 3843 818 3887 822
rect 3891 818 4023 822
rect 4027 818 4047 822
rect 4051 818 4159 822
rect 4163 818 4183 822
rect 4187 818 4295 822
rect 4299 818 4319 822
rect 4323 818 4431 822
rect 4435 818 4455 822
rect 4459 818 4567 822
rect 4571 818 4591 822
rect 4595 818 4703 822
rect 4707 818 4727 822
rect 4731 818 4839 822
rect 4843 818 5663 822
rect 5667 818 5695 822
rect 3817 817 5695 818
rect 5701 817 5702 823
rect 3822 705 3823 711
rect 3829 710 5707 711
rect 3829 706 3839 710
rect 3843 706 3859 710
rect 3863 706 3995 710
rect 3999 706 4131 710
rect 4135 706 4267 710
rect 4271 706 4403 710
rect 4407 706 4539 710
rect 4543 706 4675 710
rect 4679 706 4811 710
rect 4815 706 4947 710
rect 4951 706 5083 710
rect 5087 706 5663 710
rect 5667 706 5707 710
rect 3829 705 5707 706
rect 5713 705 5714 711
rect 1958 698 3830 699
rect 1958 695 1975 698
rect 96 689 97 695
rect 103 694 1959 695
rect 103 690 111 694
rect 115 690 131 694
rect 135 690 211 694
rect 215 690 347 694
rect 351 690 411 694
rect 415 690 587 694
rect 591 690 619 694
rect 623 690 827 694
rect 831 690 1035 694
rect 1039 690 1067 694
rect 1071 690 1315 694
rect 1319 690 1563 694
rect 1567 690 1787 694
rect 1791 690 1935 694
rect 1939 690 1959 694
rect 103 689 1959 690
rect 1965 694 1975 695
rect 1979 694 1995 698
rect 1999 694 2139 698
rect 2143 694 2299 698
rect 2303 694 2307 698
rect 2311 694 2467 698
rect 2471 694 2627 698
rect 2631 694 2635 698
rect 2639 694 2795 698
rect 2799 694 2963 698
rect 2967 694 2979 698
rect 2983 694 3323 698
rect 3327 694 3651 698
rect 3655 694 3799 698
rect 3803 694 3830 698
rect 1965 693 3830 694
rect 1965 689 1966 693
rect 1946 581 1947 587
rect 1953 586 3811 587
rect 1953 582 1975 586
rect 1979 582 2023 586
rect 2027 582 2327 586
rect 2331 582 2335 586
rect 2339 582 2527 586
rect 2531 582 2663 586
rect 2667 582 2711 586
rect 2715 582 2887 586
rect 2891 582 3007 586
rect 3011 582 3063 586
rect 3067 582 3231 586
rect 3235 582 3351 586
rect 3355 582 3407 586
rect 3411 582 3583 586
rect 3587 582 3679 586
rect 3683 582 3799 586
rect 3803 582 3811 586
rect 1953 581 3811 582
rect 3817 581 3818 587
rect 1946 579 1954 581
rect 84 573 85 579
rect 91 578 1947 579
rect 91 574 111 578
rect 115 574 159 578
rect 163 574 375 578
rect 379 574 407 578
rect 411 574 615 578
rect 619 574 671 578
rect 675 574 855 578
rect 859 574 935 578
rect 939 574 1095 578
rect 1099 574 1191 578
rect 1195 574 1343 578
rect 1347 574 1447 578
rect 1451 574 1591 578
rect 1595 574 1711 578
rect 1715 574 1815 578
rect 1819 574 1935 578
rect 1939 574 1947 578
rect 91 573 1947 574
rect 1953 573 1954 579
rect 3810 579 3818 581
rect 3810 573 3811 579
rect 3817 578 5695 579
rect 3817 574 3839 578
rect 3843 574 3887 578
rect 3891 574 4023 578
rect 4027 574 4047 578
rect 4051 574 4159 578
rect 4163 574 4207 578
rect 4211 574 4295 578
rect 4299 574 4367 578
rect 4371 574 4431 578
rect 4435 574 4527 578
rect 4531 574 4567 578
rect 4571 574 4687 578
rect 4691 574 4703 578
rect 4707 574 4839 578
rect 4843 574 4975 578
rect 4979 574 5111 578
rect 5115 574 5663 578
rect 5667 574 5695 578
rect 3817 573 5695 574
rect 5701 573 5702 579
rect 1958 469 1959 475
rect 1965 474 3823 475
rect 1965 470 1975 474
rect 1979 470 2171 474
rect 2175 470 2307 474
rect 2311 470 2315 474
rect 2319 470 2459 474
rect 2463 470 2499 474
rect 2503 470 2603 474
rect 2607 470 2683 474
rect 2687 470 2747 474
rect 2751 470 2859 474
rect 2863 470 2891 474
rect 2895 470 3035 474
rect 3039 470 3203 474
rect 3207 470 3379 474
rect 3383 470 3555 474
rect 3559 470 3799 474
rect 3803 470 3823 474
rect 1965 469 3823 470
rect 3829 469 3830 475
rect 1958 467 1966 469
rect 96 461 97 467
rect 103 466 1959 467
rect 103 462 111 466
rect 115 462 131 466
rect 135 462 195 466
rect 199 462 379 466
rect 383 462 427 466
rect 431 462 643 466
rect 647 462 659 466
rect 663 462 883 466
rect 887 462 907 466
rect 911 462 1099 466
rect 1103 462 1163 466
rect 1167 462 1323 466
rect 1327 462 1419 466
rect 1423 462 1547 466
rect 1551 462 1683 466
rect 1687 462 1935 466
rect 1939 462 1959 466
rect 103 461 1959 462
rect 1965 461 1966 467
rect 3822 453 3823 459
rect 3829 458 5707 459
rect 3829 454 3839 458
rect 3843 454 3931 458
rect 3935 454 4019 458
rect 4023 454 4131 458
rect 4135 454 4179 458
rect 4183 454 4331 458
rect 4335 454 4339 458
rect 4343 454 4499 458
rect 4503 454 4523 458
rect 4527 454 4659 458
rect 4663 454 4723 458
rect 4727 454 4923 458
rect 4927 454 5663 458
rect 5667 454 5707 458
rect 3829 453 5707 454
rect 5713 453 5714 459
rect 1946 353 1947 359
rect 1953 358 3811 359
rect 1953 354 1975 358
rect 1979 354 2023 358
rect 2027 354 2175 358
rect 2179 354 2199 358
rect 2203 354 2343 358
rect 2347 354 2367 358
rect 2371 354 2487 358
rect 2491 354 2591 358
rect 2595 354 2631 358
rect 2635 354 2775 358
rect 2779 354 2847 358
rect 2851 354 2919 358
rect 2923 354 3063 358
rect 3067 354 3119 358
rect 3123 354 3407 358
rect 3411 354 3679 358
rect 3683 354 3799 358
rect 3803 354 3811 358
rect 1953 353 3811 354
rect 3817 353 3818 359
rect 84 341 85 347
rect 91 346 1947 347
rect 91 342 111 346
rect 115 342 223 346
rect 227 342 351 346
rect 355 342 455 346
rect 459 342 575 346
rect 579 342 687 346
rect 691 342 799 346
rect 803 342 911 346
rect 915 342 1015 346
rect 1019 342 1127 346
rect 1131 342 1231 346
rect 1235 342 1351 346
rect 1355 342 1455 346
rect 1459 342 1575 346
rect 1579 342 1935 346
rect 1939 342 1947 346
rect 91 341 1947 342
rect 1953 341 1954 347
rect 3810 341 3811 347
rect 3817 346 5695 347
rect 3817 342 3839 346
rect 3843 342 3887 346
rect 3891 342 3959 346
rect 3963 342 4135 346
rect 4139 342 4159 346
rect 4163 342 4359 346
rect 4363 342 4383 346
rect 4387 342 4551 346
rect 4555 342 4615 346
rect 4619 342 4751 346
rect 4755 342 4823 346
rect 4827 342 4951 346
rect 4955 342 5015 346
rect 5019 342 5199 346
rect 5203 342 5383 346
rect 5387 342 5543 346
rect 5547 342 5663 346
rect 5667 342 5695 346
rect 3817 341 5695 342
rect 5701 341 5702 347
rect 3822 222 5714 223
rect 3822 219 3839 222
rect 1958 213 1959 219
rect 1965 218 3823 219
rect 1965 214 1975 218
rect 1979 214 1995 218
rect 1999 214 2147 218
rect 2151 214 2171 218
rect 2175 214 2339 218
rect 2343 214 2363 218
rect 2367 214 2547 218
rect 2551 214 2563 218
rect 2567 214 2723 218
rect 2727 214 2819 218
rect 2823 214 2891 218
rect 2895 214 3051 218
rect 3055 214 3091 218
rect 3095 214 3203 218
rect 3207 214 3355 218
rect 3359 214 3379 218
rect 3383 214 3515 218
rect 3519 214 3651 218
rect 3655 214 3799 218
rect 3803 214 3823 218
rect 1965 213 3823 214
rect 3829 218 3839 219
rect 3843 218 3859 222
rect 3863 218 4107 222
rect 4111 218 4291 222
rect 4295 218 4355 222
rect 4359 218 4427 222
rect 4431 218 4563 222
rect 4567 218 4587 222
rect 4591 218 4699 222
rect 4703 218 4795 222
rect 4799 218 4835 222
rect 4839 218 4971 222
rect 4975 218 4987 222
rect 4991 218 5107 222
rect 5111 218 5171 222
rect 5175 218 5243 222
rect 5247 218 5355 222
rect 5359 218 5379 222
rect 5383 218 5515 222
rect 5519 218 5663 222
rect 5667 218 5714 222
rect 3829 217 5714 218
rect 3829 213 3830 217
rect 96 193 97 199
rect 103 198 1959 199
rect 103 194 111 198
rect 115 194 131 198
rect 135 194 267 198
rect 271 194 323 198
rect 327 194 403 198
rect 407 194 539 198
rect 543 194 547 198
rect 551 194 675 198
rect 679 194 771 198
rect 775 194 811 198
rect 815 194 947 198
rect 951 194 987 198
rect 991 194 1083 198
rect 1087 194 1203 198
rect 1207 194 1227 198
rect 1231 194 1371 198
rect 1375 194 1427 198
rect 1431 194 1515 198
rect 1519 194 1651 198
rect 1655 194 1787 198
rect 1791 194 1935 198
rect 1939 194 1959 198
rect 103 193 1959 194
rect 1965 193 1966 199
rect 3810 110 5702 111
rect 3810 107 3839 110
rect 1946 101 1947 107
rect 1953 106 3811 107
rect 1953 102 1975 106
rect 1979 102 2023 106
rect 2027 102 2199 106
rect 2203 102 2391 106
rect 2395 102 2575 106
rect 2579 102 2751 106
rect 2755 102 2919 106
rect 2923 102 3079 106
rect 3083 102 3231 106
rect 3235 102 3383 106
rect 3387 102 3543 106
rect 3547 102 3679 106
rect 3683 102 3799 106
rect 3803 102 3811 106
rect 1953 101 3811 102
rect 3817 106 3839 107
rect 3843 106 4319 110
rect 4323 106 4455 110
rect 4459 106 4591 110
rect 4595 106 4727 110
rect 4731 106 4863 110
rect 4867 106 4999 110
rect 5003 106 5135 110
rect 5139 106 5271 110
rect 5275 106 5407 110
rect 5411 106 5543 110
rect 5547 106 5663 110
rect 5667 106 5702 110
rect 3817 105 5702 106
rect 3817 101 3818 105
rect 84 81 85 87
rect 91 86 1947 87
rect 91 82 111 86
rect 115 82 159 86
rect 163 82 295 86
rect 299 82 431 86
rect 435 82 567 86
rect 571 82 703 86
rect 707 82 839 86
rect 843 82 975 86
rect 979 82 1111 86
rect 1115 82 1255 86
rect 1259 82 1399 86
rect 1403 82 1543 86
rect 1547 82 1679 86
rect 1683 82 1815 86
rect 1819 82 1935 86
rect 1939 82 1947 86
rect 91 81 1947 82
rect 1953 81 1954 87
<< m5c >>
rect 85 5729 91 5735
rect 1947 5729 1953 5735
rect 1947 5669 1953 5675
rect 3811 5669 3817 5675
rect 97 5601 103 5607
rect 1959 5601 1965 5607
rect 3823 5605 3829 5611
rect 5707 5605 5713 5611
rect 1959 5557 1965 5563
rect 3823 5557 3829 5563
rect 3811 5493 3817 5499
rect 5695 5493 5701 5499
rect 85 5477 91 5483
rect 1947 5477 1953 5483
rect 1947 5433 1953 5439
rect 3811 5433 3817 5439
rect 3823 5381 3829 5387
rect 5707 5381 5713 5387
rect 97 5365 103 5371
rect 1959 5365 1965 5371
rect 1959 5285 1965 5291
rect 3823 5285 3829 5291
rect 85 5253 91 5259
rect 1947 5253 1953 5259
rect 3811 5241 3817 5247
rect 5695 5241 5701 5247
rect 1947 5169 1953 5175
rect 3811 5169 3817 5175
rect 97 5125 103 5131
rect 1959 5125 1965 5131
rect 3823 5129 3829 5135
rect 5707 5129 5713 5135
rect 1959 5057 1965 5063
rect 3823 5057 3829 5063
rect 85 5001 91 5007
rect 1947 5001 1953 5007
rect 3811 5001 3817 5007
rect 5695 5001 5701 5007
rect 1947 4937 1953 4943
rect 3811 4937 3817 4943
rect 97 4881 103 4887
rect 1959 4881 1965 4887
rect 3823 4877 3829 4883
rect 5707 4877 5713 4883
rect 1959 4797 1965 4803
rect 3823 4797 3829 4803
rect 85 4765 91 4771
rect 1947 4765 1953 4771
rect 3811 4745 3817 4751
rect 5695 4745 5701 4751
rect 1947 4655 1953 4661
rect 97 4645 103 4651
rect 1959 4645 1965 4651
rect 3811 4645 3817 4651
rect 3823 4613 3829 4619
rect 5707 4613 5713 4619
rect 85 4533 91 4539
rect 1947 4533 1953 4539
rect 1959 4533 1965 4539
rect 3823 4533 3829 4539
rect 3811 4485 3817 4491
rect 5695 4485 5701 4491
rect 1947 4427 1953 4433
rect 97 4417 103 4423
rect 1959 4417 1965 4423
rect 3811 4417 3817 4423
rect 3823 4353 3829 4359
rect 5707 4353 5713 4359
rect 85 4305 91 4311
rect 1947 4305 1953 4311
rect 1959 4297 1965 4303
rect 3823 4297 3829 4303
rect 3811 4221 3817 4227
rect 5695 4221 5701 4227
rect 1947 4191 1953 4197
rect 97 4181 103 4187
rect 1959 4181 1965 4187
rect 3811 4181 3817 4187
rect 3823 4105 3829 4111
rect 5707 4105 5713 4111
rect 1959 4069 1965 4075
rect 3823 4069 3829 4075
rect 85 4053 91 4059
rect 1947 4053 1953 4059
rect 3811 3985 3817 3991
rect 5695 3985 5701 3991
rect 1947 3951 1953 3957
rect 97 3941 103 3947
rect 1959 3941 1965 3947
rect 3811 3937 3817 3943
rect 3823 3853 3829 3859
rect 5707 3853 5713 3859
rect 85 3829 91 3835
rect 1947 3829 1953 3835
rect 1959 3813 1965 3819
rect 3823 3813 3829 3819
rect 3811 3717 3817 3723
rect 5695 3717 5701 3723
rect 1947 3703 1953 3709
rect 97 3693 103 3699
rect 1959 3693 1965 3699
rect 3811 3693 3817 3699
rect 3823 3601 3829 3607
rect 5707 3601 5713 3607
rect 1959 3569 1965 3575
rect 3823 3569 3829 3575
rect 3811 3489 3817 3495
rect 5695 3489 5701 3495
rect 1947 3421 1953 3427
rect 3811 3421 3817 3427
rect 3823 3369 3829 3375
rect 5707 3369 5713 3375
rect 1959 3309 1965 3315
rect 3823 3309 3829 3315
rect 85 3293 91 3299
rect 1947 3293 1953 3299
rect 3811 3245 3817 3251
rect 5695 3245 5701 3251
rect 1947 3193 1953 3199
rect 3811 3193 3817 3199
rect 97 3153 103 3159
rect 1959 3153 1965 3159
rect 3823 3129 3829 3135
rect 5707 3129 5713 3135
rect 1959 3061 1965 3067
rect 3823 3061 3829 3067
rect 85 3041 91 3047
rect 1947 3041 1953 3047
rect 3811 3017 3817 3023
rect 5695 3017 5701 3023
rect 1947 2941 1953 2947
rect 3811 2941 3817 2947
rect 97 2929 103 2935
rect 1959 2929 1965 2935
rect 3823 2905 3829 2911
rect 5707 2905 5713 2911
rect 1959 2829 1965 2835
rect 3823 2829 3829 2835
rect 85 2785 91 2791
rect 1947 2785 1953 2791
rect 3811 2785 3817 2791
rect 5695 2785 5701 2791
rect 1947 2717 1953 2723
rect 3811 2717 3817 2723
rect 3823 2669 3829 2675
rect 5707 2669 5713 2675
rect 97 2653 103 2659
rect 1959 2653 1965 2659
rect 1959 2605 1965 2611
rect 3823 2605 3829 2611
rect 3811 2553 3817 2559
rect 5695 2553 5701 2559
rect 85 2529 91 2535
rect 1947 2529 1953 2535
rect 1947 2485 1953 2491
rect 3811 2485 3817 2491
rect 3823 2425 3829 2431
rect 5707 2425 5713 2431
rect 97 2409 103 2415
rect 1959 2409 1965 2415
rect 1959 2365 1965 2371
rect 3823 2365 3829 2371
rect 85 2289 91 2295
rect 1947 2289 1953 2295
rect 3811 2293 3817 2299
rect 5695 2293 5701 2299
rect 1947 2225 1953 2231
rect 3811 2225 3817 2231
rect 3823 2181 3829 2187
rect 5707 2181 5713 2187
rect 97 2157 103 2163
rect 1959 2157 1965 2163
rect 1959 2081 1965 2087
rect 3823 2081 3829 2087
rect 3811 2049 3817 2055
rect 5695 2049 5701 2055
rect 85 2037 91 2043
rect 1947 2037 1953 2043
rect 1947 1957 1953 1963
rect 3811 1957 3817 1963
rect 97 1921 103 1927
rect 1959 1921 1965 1927
rect 3823 1917 3829 1923
rect 5707 1917 5713 1923
rect 1959 1845 1965 1851
rect 3823 1845 3829 1851
rect 3811 1805 3817 1811
rect 5695 1805 5701 1811
rect 85 1797 91 1803
rect 1947 1797 1953 1803
rect 1947 1733 1953 1739
rect 3811 1733 3817 1739
rect 3823 1677 3829 1683
rect 5707 1677 5713 1683
rect 97 1669 103 1675
rect 1959 1669 1965 1675
rect 1959 1621 1965 1627
rect 3823 1621 3829 1627
rect 85 1549 91 1555
rect 1947 1549 1953 1555
rect 3811 1549 3817 1555
rect 5695 1549 5701 1555
rect 97 1437 103 1443
rect 1959 1437 1965 1443
rect 3823 1433 3829 1439
rect 5707 1433 5713 1439
rect 85 1317 91 1323
rect 1947 1317 1953 1323
rect 3811 1321 3817 1327
rect 5695 1321 5701 1327
rect 1947 1305 1953 1311
rect 3811 1305 3817 1311
rect 97 1205 103 1211
rect 1959 1205 1965 1211
rect 3823 1197 3829 1203
rect 5707 1197 5713 1203
rect 1959 1181 1965 1187
rect 3823 1181 3829 1187
rect 85 1069 91 1075
rect 1947 1069 1953 1075
rect 97 945 103 951
rect 1959 945 1965 951
rect 1947 833 1953 839
rect 3811 833 3817 839
rect 85 821 91 827
rect 1947 821 1953 827
rect 3811 817 3817 823
rect 5695 817 5701 823
rect 3823 705 3829 711
rect 5707 705 5713 711
rect 97 689 103 695
rect 1959 689 1965 695
rect 1947 581 1953 587
rect 3811 581 3817 587
rect 85 573 91 579
rect 1947 573 1953 579
rect 3811 573 3817 579
rect 5695 573 5701 579
rect 1959 469 1965 475
rect 3823 469 3829 475
rect 97 461 103 467
rect 1959 461 1965 467
rect 3823 453 3829 459
rect 5707 453 5713 459
rect 1947 353 1953 359
rect 3811 353 3817 359
rect 85 341 91 347
rect 1947 341 1953 347
rect 3811 341 3817 347
rect 5695 341 5701 347
rect 1959 213 1965 219
rect 3823 213 3829 219
rect 97 193 103 199
rect 1959 193 1965 199
rect 1947 101 1953 107
rect 3811 101 3817 107
rect 85 81 91 87
rect 1947 81 1953 87
<< m5 >>
rect 84 5735 92 5760
rect 84 5729 85 5735
rect 91 5729 92 5735
rect 84 5483 92 5729
rect 84 5477 85 5483
rect 91 5477 92 5483
rect 84 5259 92 5477
rect 84 5253 85 5259
rect 91 5253 92 5259
rect 84 5007 92 5253
rect 84 5001 85 5007
rect 91 5001 92 5007
rect 84 4771 92 5001
rect 84 4765 85 4771
rect 91 4765 92 4771
rect 84 4539 92 4765
rect 84 4533 85 4539
rect 91 4533 92 4539
rect 84 4311 92 4533
rect 84 4305 85 4311
rect 91 4305 92 4311
rect 84 4059 92 4305
rect 84 4053 85 4059
rect 91 4053 92 4059
rect 84 3835 92 4053
rect 84 3829 85 3835
rect 91 3829 92 3835
rect 84 3299 92 3829
rect 84 3293 85 3299
rect 91 3293 92 3299
rect 84 3047 92 3293
rect 84 3041 85 3047
rect 91 3041 92 3047
rect 84 2791 92 3041
rect 84 2785 85 2791
rect 91 2785 92 2791
rect 84 2535 92 2785
rect 84 2529 85 2535
rect 91 2529 92 2535
rect 84 2295 92 2529
rect 84 2289 85 2295
rect 91 2289 92 2295
rect 84 2043 92 2289
rect 84 2037 85 2043
rect 91 2037 92 2043
rect 84 1803 92 2037
rect 84 1797 85 1803
rect 91 1797 92 1803
rect 84 1555 92 1797
rect 84 1549 85 1555
rect 91 1549 92 1555
rect 84 1323 92 1549
rect 84 1317 85 1323
rect 91 1317 92 1323
rect 84 1075 92 1317
rect 84 1069 85 1075
rect 91 1069 92 1075
rect 84 827 92 1069
rect 84 821 85 827
rect 91 821 92 827
rect 84 579 92 821
rect 84 573 85 579
rect 91 573 92 579
rect 84 347 92 573
rect 84 341 85 347
rect 91 341 92 347
rect 84 87 92 341
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 5607 104 5760
rect 96 5601 97 5607
rect 103 5601 104 5607
rect 96 5371 104 5601
rect 96 5365 97 5371
rect 103 5365 104 5371
rect 96 5131 104 5365
rect 96 5125 97 5131
rect 103 5125 104 5131
rect 96 4887 104 5125
rect 96 4881 97 4887
rect 103 4881 104 4887
rect 96 4651 104 4881
rect 96 4645 97 4651
rect 103 4645 104 4651
rect 96 4423 104 4645
rect 96 4417 97 4423
rect 103 4417 104 4423
rect 96 4187 104 4417
rect 96 4181 97 4187
rect 103 4181 104 4187
rect 96 3947 104 4181
rect 96 3941 97 3947
rect 103 3941 104 3947
rect 96 3699 104 3941
rect 96 3693 97 3699
rect 103 3693 104 3699
rect 96 3159 104 3693
rect 96 3153 97 3159
rect 103 3153 104 3159
rect 96 2935 104 3153
rect 96 2929 97 2935
rect 103 2929 104 2935
rect 96 2659 104 2929
rect 96 2653 97 2659
rect 103 2653 104 2659
rect 96 2415 104 2653
rect 96 2409 97 2415
rect 103 2409 104 2415
rect 96 2163 104 2409
rect 96 2157 97 2163
rect 103 2157 104 2163
rect 96 1927 104 2157
rect 96 1921 97 1927
rect 103 1921 104 1927
rect 96 1675 104 1921
rect 96 1669 97 1675
rect 103 1669 104 1675
rect 96 1443 104 1669
rect 96 1437 97 1443
rect 103 1437 104 1443
rect 96 1211 104 1437
rect 96 1205 97 1211
rect 103 1205 104 1211
rect 96 951 104 1205
rect 96 945 97 951
rect 103 945 104 951
rect 96 695 104 945
rect 96 689 97 695
rect 103 689 104 695
rect 96 467 104 689
rect 96 461 97 467
rect 103 461 104 467
rect 96 199 104 461
rect 96 193 97 199
rect 103 193 104 199
rect 96 72 104 193
rect 1946 5735 1954 5760
rect 1946 5729 1947 5735
rect 1953 5729 1954 5735
rect 1946 5675 1954 5729
rect 1946 5669 1947 5675
rect 1953 5669 1954 5675
rect 1946 5483 1954 5669
rect 1946 5477 1947 5483
rect 1953 5477 1954 5483
rect 1946 5439 1954 5477
rect 1946 5433 1947 5439
rect 1953 5433 1954 5439
rect 1946 5259 1954 5433
rect 1946 5253 1947 5259
rect 1953 5253 1954 5259
rect 1946 5175 1954 5253
rect 1946 5169 1947 5175
rect 1953 5169 1954 5175
rect 1946 5007 1954 5169
rect 1946 5001 1947 5007
rect 1953 5001 1954 5007
rect 1946 4943 1954 5001
rect 1946 4937 1947 4943
rect 1953 4937 1954 4943
rect 1946 4771 1954 4937
rect 1946 4765 1947 4771
rect 1953 4765 1954 4771
rect 1946 4661 1954 4765
rect 1946 4655 1947 4661
rect 1953 4655 1954 4661
rect 1946 4539 1954 4655
rect 1946 4533 1947 4539
rect 1953 4533 1954 4539
rect 1946 4433 1954 4533
rect 1946 4427 1947 4433
rect 1953 4427 1954 4433
rect 1946 4311 1954 4427
rect 1946 4305 1947 4311
rect 1953 4305 1954 4311
rect 1946 4197 1954 4305
rect 1946 4191 1947 4197
rect 1953 4191 1954 4197
rect 1946 4059 1954 4191
rect 1946 4053 1947 4059
rect 1953 4053 1954 4059
rect 1946 3957 1954 4053
rect 1946 3951 1947 3957
rect 1953 3951 1954 3957
rect 1946 3835 1954 3951
rect 1946 3829 1947 3835
rect 1953 3829 1954 3835
rect 1946 3709 1954 3829
rect 1946 3703 1947 3709
rect 1953 3703 1954 3709
rect 1946 3427 1954 3703
rect 1946 3421 1947 3427
rect 1953 3421 1954 3427
rect 1946 3299 1954 3421
rect 1946 3293 1947 3299
rect 1953 3293 1954 3299
rect 1946 3199 1954 3293
rect 1946 3193 1947 3199
rect 1953 3193 1954 3199
rect 1946 3047 1954 3193
rect 1946 3041 1947 3047
rect 1953 3041 1954 3047
rect 1946 2947 1954 3041
rect 1946 2941 1947 2947
rect 1953 2941 1954 2947
rect 1946 2791 1954 2941
rect 1946 2785 1947 2791
rect 1953 2785 1954 2791
rect 1946 2723 1954 2785
rect 1946 2717 1947 2723
rect 1953 2717 1954 2723
rect 1946 2535 1954 2717
rect 1946 2529 1947 2535
rect 1953 2529 1954 2535
rect 1946 2491 1954 2529
rect 1946 2485 1947 2491
rect 1953 2485 1954 2491
rect 1946 2295 1954 2485
rect 1946 2289 1947 2295
rect 1953 2289 1954 2295
rect 1946 2231 1954 2289
rect 1946 2225 1947 2231
rect 1953 2225 1954 2231
rect 1946 2043 1954 2225
rect 1946 2037 1947 2043
rect 1953 2037 1954 2043
rect 1946 1963 1954 2037
rect 1946 1957 1947 1963
rect 1953 1957 1954 1963
rect 1946 1803 1954 1957
rect 1946 1797 1947 1803
rect 1953 1797 1954 1803
rect 1946 1739 1954 1797
rect 1946 1733 1947 1739
rect 1953 1733 1954 1739
rect 1946 1555 1954 1733
rect 1946 1549 1947 1555
rect 1953 1549 1954 1555
rect 1946 1323 1954 1549
rect 1946 1317 1947 1323
rect 1953 1317 1954 1323
rect 1946 1311 1954 1317
rect 1946 1305 1947 1311
rect 1953 1305 1954 1311
rect 1946 1075 1954 1305
rect 1946 1069 1947 1075
rect 1953 1069 1954 1075
rect 1946 839 1954 1069
rect 1946 833 1947 839
rect 1953 833 1954 839
rect 1946 827 1954 833
rect 1946 821 1947 827
rect 1953 821 1954 827
rect 1946 587 1954 821
rect 1946 581 1947 587
rect 1953 581 1954 587
rect 1946 579 1954 581
rect 1946 573 1947 579
rect 1953 573 1954 579
rect 1946 359 1954 573
rect 1946 353 1947 359
rect 1953 353 1954 359
rect 1946 347 1954 353
rect 1946 341 1947 347
rect 1953 341 1954 347
rect 1946 107 1954 341
rect 1946 101 1947 107
rect 1953 101 1954 107
rect 1946 87 1954 101
rect 1946 81 1947 87
rect 1953 81 1954 87
rect 1946 72 1954 81
rect 1958 5607 1966 5760
rect 1958 5601 1959 5607
rect 1965 5601 1966 5607
rect 1958 5563 1966 5601
rect 1958 5557 1959 5563
rect 1965 5557 1966 5563
rect 1958 5371 1966 5557
rect 1958 5365 1959 5371
rect 1965 5365 1966 5371
rect 1958 5291 1966 5365
rect 1958 5285 1959 5291
rect 1965 5285 1966 5291
rect 1958 5131 1966 5285
rect 1958 5125 1959 5131
rect 1965 5125 1966 5131
rect 1958 5063 1966 5125
rect 1958 5057 1959 5063
rect 1965 5057 1966 5063
rect 1958 4887 1966 5057
rect 1958 4881 1959 4887
rect 1965 4881 1966 4887
rect 1958 4803 1966 4881
rect 1958 4797 1959 4803
rect 1965 4797 1966 4803
rect 1958 4651 1966 4797
rect 1958 4645 1959 4651
rect 1965 4645 1966 4651
rect 1958 4539 1966 4645
rect 1958 4533 1959 4539
rect 1965 4533 1966 4539
rect 1958 4423 1966 4533
rect 1958 4417 1959 4423
rect 1965 4417 1966 4423
rect 1958 4303 1966 4417
rect 1958 4297 1959 4303
rect 1965 4297 1966 4303
rect 1958 4187 1966 4297
rect 1958 4181 1959 4187
rect 1965 4181 1966 4187
rect 1958 4075 1966 4181
rect 1958 4069 1959 4075
rect 1965 4069 1966 4075
rect 1958 3947 1966 4069
rect 1958 3941 1959 3947
rect 1965 3941 1966 3947
rect 1958 3819 1966 3941
rect 1958 3813 1959 3819
rect 1965 3813 1966 3819
rect 1958 3699 1966 3813
rect 1958 3693 1959 3699
rect 1965 3693 1966 3699
rect 1958 3575 1966 3693
rect 1958 3569 1959 3575
rect 1965 3569 1966 3575
rect 1958 3315 1966 3569
rect 1958 3309 1959 3315
rect 1965 3309 1966 3315
rect 1958 3159 1966 3309
rect 1958 3153 1959 3159
rect 1965 3153 1966 3159
rect 1958 3067 1966 3153
rect 1958 3061 1959 3067
rect 1965 3061 1966 3067
rect 1958 2935 1966 3061
rect 1958 2929 1959 2935
rect 1965 2929 1966 2935
rect 1958 2835 1966 2929
rect 1958 2829 1959 2835
rect 1965 2829 1966 2835
rect 1958 2659 1966 2829
rect 1958 2653 1959 2659
rect 1965 2653 1966 2659
rect 1958 2611 1966 2653
rect 1958 2605 1959 2611
rect 1965 2605 1966 2611
rect 1958 2415 1966 2605
rect 1958 2409 1959 2415
rect 1965 2409 1966 2415
rect 1958 2371 1966 2409
rect 1958 2365 1959 2371
rect 1965 2365 1966 2371
rect 1958 2163 1966 2365
rect 1958 2157 1959 2163
rect 1965 2157 1966 2163
rect 1958 2087 1966 2157
rect 1958 2081 1959 2087
rect 1965 2081 1966 2087
rect 1958 1927 1966 2081
rect 1958 1921 1959 1927
rect 1965 1921 1966 1927
rect 1958 1851 1966 1921
rect 1958 1845 1959 1851
rect 1965 1845 1966 1851
rect 1958 1675 1966 1845
rect 1958 1669 1959 1675
rect 1965 1669 1966 1675
rect 1958 1627 1966 1669
rect 1958 1621 1959 1627
rect 1965 1621 1966 1627
rect 1958 1443 1966 1621
rect 1958 1437 1959 1443
rect 1965 1437 1966 1443
rect 1958 1211 1966 1437
rect 1958 1205 1959 1211
rect 1965 1205 1966 1211
rect 1958 1187 1966 1205
rect 1958 1181 1959 1187
rect 1965 1181 1966 1187
rect 1958 951 1966 1181
rect 1958 945 1959 951
rect 1965 945 1966 951
rect 1958 695 1966 945
rect 1958 689 1959 695
rect 1965 689 1966 695
rect 1958 475 1966 689
rect 1958 469 1959 475
rect 1965 469 1966 475
rect 1958 467 1966 469
rect 1958 461 1959 467
rect 1965 461 1966 467
rect 1958 219 1966 461
rect 1958 213 1959 219
rect 1965 213 1966 219
rect 1958 199 1966 213
rect 1958 193 1959 199
rect 1965 193 1966 199
rect 1958 72 1966 193
rect 3810 5675 3818 5760
rect 3810 5669 3811 5675
rect 3817 5669 3818 5675
rect 3810 5499 3818 5669
rect 3810 5493 3811 5499
rect 3817 5493 3818 5499
rect 3810 5439 3818 5493
rect 3810 5433 3811 5439
rect 3817 5433 3818 5439
rect 3810 5247 3818 5433
rect 3810 5241 3811 5247
rect 3817 5241 3818 5247
rect 3810 5175 3818 5241
rect 3810 5169 3811 5175
rect 3817 5169 3818 5175
rect 3810 5007 3818 5169
rect 3810 5001 3811 5007
rect 3817 5001 3818 5007
rect 3810 4943 3818 5001
rect 3810 4937 3811 4943
rect 3817 4937 3818 4943
rect 3810 4751 3818 4937
rect 3810 4745 3811 4751
rect 3817 4745 3818 4751
rect 3810 4651 3818 4745
rect 3810 4645 3811 4651
rect 3817 4645 3818 4651
rect 3810 4491 3818 4645
rect 3810 4485 3811 4491
rect 3817 4485 3818 4491
rect 3810 4423 3818 4485
rect 3810 4417 3811 4423
rect 3817 4417 3818 4423
rect 3810 4227 3818 4417
rect 3810 4221 3811 4227
rect 3817 4221 3818 4227
rect 3810 4187 3818 4221
rect 3810 4181 3811 4187
rect 3817 4181 3818 4187
rect 3810 3991 3818 4181
rect 3810 3985 3811 3991
rect 3817 3985 3818 3991
rect 3810 3943 3818 3985
rect 3810 3937 3811 3943
rect 3817 3937 3818 3943
rect 3810 3723 3818 3937
rect 3810 3717 3811 3723
rect 3817 3717 3818 3723
rect 3810 3699 3818 3717
rect 3810 3693 3811 3699
rect 3817 3693 3818 3699
rect 3810 3495 3818 3693
rect 3810 3489 3811 3495
rect 3817 3489 3818 3495
rect 3810 3427 3818 3489
rect 3810 3421 3811 3427
rect 3817 3421 3818 3427
rect 3810 3251 3818 3421
rect 3810 3245 3811 3251
rect 3817 3245 3818 3251
rect 3810 3199 3818 3245
rect 3810 3193 3811 3199
rect 3817 3193 3818 3199
rect 3810 3023 3818 3193
rect 3810 3017 3811 3023
rect 3817 3017 3818 3023
rect 3810 2947 3818 3017
rect 3810 2941 3811 2947
rect 3817 2941 3818 2947
rect 3810 2791 3818 2941
rect 3810 2785 3811 2791
rect 3817 2785 3818 2791
rect 3810 2723 3818 2785
rect 3810 2717 3811 2723
rect 3817 2717 3818 2723
rect 3810 2559 3818 2717
rect 3810 2553 3811 2559
rect 3817 2553 3818 2559
rect 3810 2491 3818 2553
rect 3810 2485 3811 2491
rect 3817 2485 3818 2491
rect 3810 2299 3818 2485
rect 3810 2293 3811 2299
rect 3817 2293 3818 2299
rect 3810 2231 3818 2293
rect 3810 2225 3811 2231
rect 3817 2225 3818 2231
rect 3810 2055 3818 2225
rect 3810 2049 3811 2055
rect 3817 2049 3818 2055
rect 3810 1963 3818 2049
rect 3810 1957 3811 1963
rect 3817 1957 3818 1963
rect 3810 1811 3818 1957
rect 3810 1805 3811 1811
rect 3817 1805 3818 1811
rect 3810 1739 3818 1805
rect 3810 1733 3811 1739
rect 3817 1733 3818 1739
rect 3810 1555 3818 1733
rect 3810 1549 3811 1555
rect 3817 1549 3818 1555
rect 3810 1327 3818 1549
rect 3810 1321 3811 1327
rect 3817 1321 3818 1327
rect 3810 1311 3818 1321
rect 3810 1305 3811 1311
rect 3817 1305 3818 1311
rect 3810 839 3818 1305
rect 3810 833 3811 839
rect 3817 833 3818 839
rect 3810 823 3818 833
rect 3810 817 3811 823
rect 3817 817 3818 823
rect 3810 587 3818 817
rect 3810 581 3811 587
rect 3817 581 3818 587
rect 3810 579 3818 581
rect 3810 573 3811 579
rect 3817 573 3818 579
rect 3810 359 3818 573
rect 3810 353 3811 359
rect 3817 353 3818 359
rect 3810 347 3818 353
rect 3810 341 3811 347
rect 3817 341 3818 347
rect 3810 107 3818 341
rect 3810 101 3811 107
rect 3817 101 3818 107
rect 3810 72 3818 101
rect 3822 5611 3830 5760
rect 3822 5605 3823 5611
rect 3829 5605 3830 5611
rect 3822 5563 3830 5605
rect 3822 5557 3823 5563
rect 3829 5557 3830 5563
rect 3822 5387 3830 5557
rect 3822 5381 3823 5387
rect 3829 5381 3830 5387
rect 3822 5291 3830 5381
rect 3822 5285 3823 5291
rect 3829 5285 3830 5291
rect 3822 5135 3830 5285
rect 3822 5129 3823 5135
rect 3829 5129 3830 5135
rect 3822 5063 3830 5129
rect 3822 5057 3823 5063
rect 3829 5057 3830 5063
rect 3822 4883 3830 5057
rect 3822 4877 3823 4883
rect 3829 4877 3830 4883
rect 3822 4803 3830 4877
rect 3822 4797 3823 4803
rect 3829 4797 3830 4803
rect 3822 4619 3830 4797
rect 3822 4613 3823 4619
rect 3829 4613 3830 4619
rect 3822 4539 3830 4613
rect 3822 4533 3823 4539
rect 3829 4533 3830 4539
rect 3822 4359 3830 4533
rect 3822 4353 3823 4359
rect 3829 4353 3830 4359
rect 3822 4303 3830 4353
rect 3822 4297 3823 4303
rect 3829 4297 3830 4303
rect 3822 4111 3830 4297
rect 3822 4105 3823 4111
rect 3829 4105 3830 4111
rect 3822 4075 3830 4105
rect 3822 4069 3823 4075
rect 3829 4069 3830 4075
rect 3822 3859 3830 4069
rect 3822 3853 3823 3859
rect 3829 3853 3830 3859
rect 3822 3819 3830 3853
rect 3822 3813 3823 3819
rect 3829 3813 3830 3819
rect 3822 3607 3830 3813
rect 3822 3601 3823 3607
rect 3829 3601 3830 3607
rect 3822 3575 3830 3601
rect 3822 3569 3823 3575
rect 3829 3569 3830 3575
rect 3822 3375 3830 3569
rect 3822 3369 3823 3375
rect 3829 3369 3830 3375
rect 3822 3315 3830 3369
rect 3822 3309 3823 3315
rect 3829 3309 3830 3315
rect 3822 3135 3830 3309
rect 3822 3129 3823 3135
rect 3829 3129 3830 3135
rect 3822 3067 3830 3129
rect 3822 3061 3823 3067
rect 3829 3061 3830 3067
rect 3822 2911 3830 3061
rect 3822 2905 3823 2911
rect 3829 2905 3830 2911
rect 3822 2835 3830 2905
rect 3822 2829 3823 2835
rect 3829 2829 3830 2835
rect 3822 2675 3830 2829
rect 3822 2669 3823 2675
rect 3829 2669 3830 2675
rect 3822 2611 3830 2669
rect 3822 2605 3823 2611
rect 3829 2605 3830 2611
rect 3822 2431 3830 2605
rect 3822 2425 3823 2431
rect 3829 2425 3830 2431
rect 3822 2371 3830 2425
rect 3822 2365 3823 2371
rect 3829 2365 3830 2371
rect 3822 2187 3830 2365
rect 3822 2181 3823 2187
rect 3829 2181 3830 2187
rect 3822 2087 3830 2181
rect 3822 2081 3823 2087
rect 3829 2081 3830 2087
rect 3822 1923 3830 2081
rect 3822 1917 3823 1923
rect 3829 1917 3830 1923
rect 3822 1851 3830 1917
rect 3822 1845 3823 1851
rect 3829 1845 3830 1851
rect 3822 1683 3830 1845
rect 3822 1677 3823 1683
rect 3829 1677 3830 1683
rect 3822 1627 3830 1677
rect 3822 1621 3823 1627
rect 3829 1621 3830 1627
rect 3822 1439 3830 1621
rect 3822 1433 3823 1439
rect 3829 1433 3830 1439
rect 3822 1203 3830 1433
rect 3822 1197 3823 1203
rect 3829 1197 3830 1203
rect 3822 1187 3830 1197
rect 3822 1181 3823 1187
rect 3829 1181 3830 1187
rect 3822 711 3830 1181
rect 3822 705 3823 711
rect 3829 705 3830 711
rect 3822 475 3830 705
rect 3822 469 3823 475
rect 3829 469 3830 475
rect 3822 459 3830 469
rect 3822 453 3823 459
rect 3829 453 3830 459
rect 3822 219 3830 453
rect 3822 213 3823 219
rect 3829 213 3830 219
rect 3822 72 3830 213
rect 5694 5499 5702 5760
rect 5694 5493 5695 5499
rect 5701 5493 5702 5499
rect 5694 5247 5702 5493
rect 5694 5241 5695 5247
rect 5701 5241 5702 5247
rect 5694 5007 5702 5241
rect 5694 5001 5695 5007
rect 5701 5001 5702 5007
rect 5694 4751 5702 5001
rect 5694 4745 5695 4751
rect 5701 4745 5702 4751
rect 5694 4491 5702 4745
rect 5694 4485 5695 4491
rect 5701 4485 5702 4491
rect 5694 4227 5702 4485
rect 5694 4221 5695 4227
rect 5701 4221 5702 4227
rect 5694 3991 5702 4221
rect 5694 3985 5695 3991
rect 5701 3985 5702 3991
rect 5694 3723 5702 3985
rect 5694 3717 5695 3723
rect 5701 3717 5702 3723
rect 5694 3495 5702 3717
rect 5694 3489 5695 3495
rect 5701 3489 5702 3495
rect 5694 3251 5702 3489
rect 5694 3245 5695 3251
rect 5701 3245 5702 3251
rect 5694 3023 5702 3245
rect 5694 3017 5695 3023
rect 5701 3017 5702 3023
rect 5694 2791 5702 3017
rect 5694 2785 5695 2791
rect 5701 2785 5702 2791
rect 5694 2559 5702 2785
rect 5694 2553 5695 2559
rect 5701 2553 5702 2559
rect 5694 2299 5702 2553
rect 5694 2293 5695 2299
rect 5701 2293 5702 2299
rect 5694 2055 5702 2293
rect 5694 2049 5695 2055
rect 5701 2049 5702 2055
rect 5694 1811 5702 2049
rect 5694 1805 5695 1811
rect 5701 1805 5702 1811
rect 5694 1555 5702 1805
rect 5694 1549 5695 1555
rect 5701 1549 5702 1555
rect 5694 1327 5702 1549
rect 5694 1321 5695 1327
rect 5701 1321 5702 1327
rect 5694 823 5702 1321
rect 5694 817 5695 823
rect 5701 817 5702 823
rect 5694 579 5702 817
rect 5694 573 5695 579
rect 5701 573 5702 579
rect 5694 347 5702 573
rect 5694 341 5695 347
rect 5701 341 5702 347
rect 5694 72 5702 341
rect 5706 5611 5714 5760
rect 5706 5605 5707 5611
rect 5713 5605 5714 5611
rect 5706 5387 5714 5605
rect 5706 5381 5707 5387
rect 5713 5381 5714 5387
rect 5706 5135 5714 5381
rect 5706 5129 5707 5135
rect 5713 5129 5714 5135
rect 5706 4883 5714 5129
rect 5706 4877 5707 4883
rect 5713 4877 5714 4883
rect 5706 4619 5714 4877
rect 5706 4613 5707 4619
rect 5713 4613 5714 4619
rect 5706 4359 5714 4613
rect 5706 4353 5707 4359
rect 5713 4353 5714 4359
rect 5706 4111 5714 4353
rect 5706 4105 5707 4111
rect 5713 4105 5714 4111
rect 5706 3859 5714 4105
rect 5706 3853 5707 3859
rect 5713 3853 5714 3859
rect 5706 3607 5714 3853
rect 5706 3601 5707 3607
rect 5713 3601 5714 3607
rect 5706 3375 5714 3601
rect 5706 3369 5707 3375
rect 5713 3369 5714 3375
rect 5706 3135 5714 3369
rect 5706 3129 5707 3135
rect 5713 3129 5714 3135
rect 5706 2911 5714 3129
rect 5706 2905 5707 2911
rect 5713 2905 5714 2911
rect 5706 2675 5714 2905
rect 5706 2669 5707 2675
rect 5713 2669 5714 2675
rect 5706 2431 5714 2669
rect 5706 2425 5707 2431
rect 5713 2425 5714 2431
rect 5706 2187 5714 2425
rect 5706 2181 5707 2187
rect 5713 2181 5714 2187
rect 5706 1923 5714 2181
rect 5706 1917 5707 1923
rect 5713 1917 5714 1923
rect 5706 1683 5714 1917
rect 5706 1677 5707 1683
rect 5713 1677 5714 1683
rect 5706 1439 5714 1677
rect 5706 1433 5707 1439
rect 5713 1433 5714 1439
rect 5706 1203 5714 1433
rect 5706 1197 5707 1203
rect 5713 1197 5714 1203
rect 5706 711 5714 1197
rect 5706 705 5707 711
rect 5713 705 5714 711
rect 5706 459 5714 705
rect 5706 453 5707 459
rect 5713 453 5714 459
rect 5706 72 5714 453
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__265
timestamp 1731220455
transform 1 0 5656 0 1 5520
box 7 3 12 24
use welltap_svt  __well_tap__264
timestamp 1731220455
transform 1 0 3832 0 1 5520
box 7 3 12 24
use welltap_svt  __well_tap__263
timestamp 1731220455
transform 1 0 5656 0 -1 5472
box 7 3 12 24
use welltap_svt  __well_tap__262
timestamp 1731220455
transform 1 0 3832 0 -1 5472
box 7 3 12 24
use welltap_svt  __well_tap__261
timestamp 1731220455
transform 1 0 5656 0 1 5296
box 7 3 12 24
use welltap_svt  __well_tap__260
timestamp 1731220455
transform 1 0 3832 0 1 5296
box 7 3 12 24
use welltap_svt  __well_tap__259
timestamp 1731220455
transform 1 0 5656 0 -1 5220
box 7 3 12 24
use welltap_svt  __well_tap__258
timestamp 1731220455
transform 1 0 3832 0 -1 5220
box 7 3 12 24
use welltap_svt  __well_tap__257
timestamp 1731220455
transform 1 0 5656 0 1 5044
box 7 3 12 24
use welltap_svt  __well_tap__256
timestamp 1731220455
transform 1 0 3832 0 1 5044
box 7 3 12 24
use welltap_svt  __well_tap__255
timestamp 1731220455
transform 1 0 5656 0 -1 4980
box 7 3 12 24
use welltap_svt  __well_tap__254
timestamp 1731220455
transform 1 0 3832 0 -1 4980
box 7 3 12 24
use welltap_svt  __well_tap__253
timestamp 1731220455
transform 1 0 5656 0 1 4792
box 7 3 12 24
use welltap_svt  __well_tap__252
timestamp 1731220455
transform 1 0 3832 0 1 4792
box 7 3 12 24
use welltap_svt  __well_tap__251
timestamp 1731220455
transform 1 0 5656 0 -1 4724
box 7 3 12 24
use welltap_svt  __well_tap__250
timestamp 1731220455
transform 1 0 3832 0 -1 4724
box 7 3 12 24
use welltap_svt  __well_tap__249
timestamp 1731220455
transform 1 0 5656 0 1 4528
box 7 3 12 24
use welltap_svt  __well_tap__248
timestamp 1731220455
transform 1 0 3832 0 1 4528
box 7 3 12 24
use welltap_svt  __well_tap__247
timestamp 1731220455
transform 1 0 5656 0 -1 4464
box 7 3 12 24
use welltap_svt  __well_tap__246
timestamp 1731220455
transform 1 0 3832 0 -1 4464
box 7 3 12 24
use welltap_svt  __well_tap__245
timestamp 1731220455
transform 1 0 5656 0 1 4268
box 7 3 12 24
use welltap_svt  __well_tap__244
timestamp 1731220455
transform 1 0 3832 0 1 4268
box 7 3 12 24
use welltap_svt  __well_tap__243
timestamp 1731220455
transform 1 0 5656 0 -1 4200
box 7 3 12 24
use welltap_svt  __well_tap__242
timestamp 1731220455
transform 1 0 3832 0 -1 4200
box 7 3 12 24
use welltap_svt  __well_tap__241
timestamp 1731220455
transform 1 0 5656 0 1 4020
box 7 3 12 24
use welltap_svt  __well_tap__240
timestamp 1731220455
transform 1 0 3832 0 1 4020
box 7 3 12 24
use welltap_svt  __well_tap__239
timestamp 1731220455
transform 1 0 5656 0 -1 3964
box 7 3 12 24
use welltap_svt  __well_tap__238
timestamp 1731220455
transform 1 0 3832 0 -1 3964
box 7 3 12 24
use welltap_svt  __well_tap__237
timestamp 1731220455
transform 1 0 5656 0 1 3768
box 7 3 12 24
use welltap_svt  __well_tap__236
timestamp 1731220455
transform 1 0 3832 0 1 3768
box 7 3 12 24
use welltap_svt  __well_tap__235
timestamp 1731220455
transform 1 0 5656 0 -1 3696
box 7 3 12 24
use welltap_svt  __well_tap__234
timestamp 1731220455
transform 1 0 3832 0 -1 3696
box 7 3 12 24
use welltap_svt  __well_tap__233
timestamp 1731220455
transform 1 0 5656 0 1 3516
box 7 3 12 24
use welltap_svt  __well_tap__232
timestamp 1731220455
transform 1 0 3832 0 1 3516
box 7 3 12 24
use welltap_svt  __well_tap__231
timestamp 1731220455
transform 1 0 5656 0 -1 3468
box 7 3 12 24
use welltap_svt  __well_tap__230
timestamp 1731220455
transform 1 0 3832 0 -1 3468
box 7 3 12 24
use welltap_svt  __well_tap__229
timestamp 1731220455
transform 1 0 5656 0 1 3284
box 7 3 12 24
use welltap_svt  __well_tap__228
timestamp 1731220455
transform 1 0 3832 0 1 3284
box 7 3 12 24
use welltap_svt  __well_tap__227
timestamp 1731220455
transform 1 0 5656 0 -1 3224
box 7 3 12 24
use welltap_svt  __well_tap__226
timestamp 1731220455
transform 1 0 3832 0 -1 3224
box 7 3 12 24
use welltap_svt  __well_tap__225
timestamp 1731220455
transform 1 0 5656 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__224
timestamp 1731220455
transform 1 0 3832 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__223
timestamp 1731220455
transform 1 0 5656 0 -1 2996
box 7 3 12 24
use welltap_svt  __well_tap__222
timestamp 1731220455
transform 1 0 3832 0 -1 2996
box 7 3 12 24
use welltap_svt  __well_tap__221
timestamp 1731220455
transform 1 0 5656 0 1 2820
box 7 3 12 24
use welltap_svt  __well_tap__220
timestamp 1731220455
transform 1 0 3832 0 1 2820
box 7 3 12 24
use welltap_svt  __well_tap__219
timestamp 1731220455
transform 1 0 5656 0 -1 2764
box 7 3 12 24
use welltap_svt  __well_tap__218
timestamp 1731220455
transform 1 0 3832 0 -1 2764
box 7 3 12 24
use welltap_svt  __well_tap__217
timestamp 1731220455
transform 1 0 5656 0 1 2584
box 7 3 12 24
use welltap_svt  __well_tap__216
timestamp 1731220455
transform 1 0 3832 0 1 2584
box 7 3 12 24
use welltap_svt  __well_tap__215
timestamp 1731220455
transform 1 0 5656 0 -1 2532
box 7 3 12 24
use welltap_svt  __well_tap__214
timestamp 1731220455
transform 1 0 3832 0 -1 2532
box 7 3 12 24
use welltap_svt  __well_tap__213
timestamp 1731220455
transform 1 0 5656 0 1 2340
box 7 3 12 24
use welltap_svt  __well_tap__212
timestamp 1731220455
transform 1 0 3832 0 1 2340
box 7 3 12 24
use welltap_svt  __well_tap__211
timestamp 1731220455
transform 1 0 5656 0 -1 2272
box 7 3 12 24
use welltap_svt  __well_tap__210
timestamp 1731220455
transform 1 0 3832 0 -1 2272
box 7 3 12 24
use welltap_svt  __well_tap__209
timestamp 1731220455
transform 1 0 5656 0 1 2096
box 7 3 12 24
use welltap_svt  __well_tap__208
timestamp 1731220455
transform 1 0 3832 0 1 2096
box 7 3 12 24
use welltap_svt  __well_tap__207
timestamp 1731220455
transform 1 0 5656 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__206
timestamp 1731220455
transform 1 0 3832 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__205
timestamp 1731220455
transform 1 0 5656 0 1 1832
box 7 3 12 24
use welltap_svt  __well_tap__204
timestamp 1731220455
transform 1 0 3832 0 1 1832
box 7 3 12 24
use welltap_svt  __well_tap__203
timestamp 1731220455
transform 1 0 5656 0 -1 1784
box 7 3 12 24
use welltap_svt  __well_tap__202
timestamp 1731220455
transform 1 0 3832 0 -1 1784
box 7 3 12 24
use welltap_svt  __well_tap__201
timestamp 1731220455
transform 1 0 5656 0 1 1592
box 7 3 12 24
use welltap_svt  __well_tap__200
timestamp 1731220455
transform 1 0 3832 0 1 1592
box 7 3 12 24
use welltap_svt  __well_tap__199
timestamp 1731220455
transform 1 0 5656 0 -1 1528
box 7 3 12 24
use welltap_svt  __well_tap__198
timestamp 1731220455
transform 1 0 3832 0 -1 1528
box 7 3 12 24
use welltap_svt  __well_tap__197
timestamp 1731220455
transform 1 0 5656 0 1 1348
box 7 3 12 24
use welltap_svt  __well_tap__196
timestamp 1731220455
transform 1 0 3832 0 1 1348
box 7 3 12 24
use welltap_svt  __well_tap__195
timestamp 1731220455
transform 1 0 5656 0 -1 1300
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220455
transform 1 0 3832 0 -1 1300
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220455
transform 1 0 5656 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220455
transform 1 0 3832 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220455
transform 1 0 5656 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220455
transform 1 0 3832 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220455
transform 1 0 5656 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220455
transform 1 0 3832 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220455
transform 1 0 5656 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220455
transform 1 0 3832 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220455
transform 1 0 5656 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220455
transform 1 0 3832 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220455
transform 1 0 5656 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220455
transform 1 0 3832 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220455
transform 1 0 5656 0 1 368
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220455
transform 1 0 3832 0 1 368
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220455
transform 1 0 5656 0 -1 320
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220455
transform 1 0 3832 0 -1 320
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220455
transform 1 0 5656 0 1 132
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220455
transform 1 0 3832 0 1 132
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220455
transform 1 0 3792 0 -1 5648
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220455
transform 1 0 1968 0 -1 5648
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220455
transform 1 0 3792 0 1 5472
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220455
transform 1 0 1968 0 1 5472
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220455
transform 1 0 3792 0 -1 5412
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220455
transform 1 0 1968 0 -1 5412
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220455
transform 1 0 3792 0 1 5200
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220455
transform 1 0 1968 0 1 5200
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220455
transform 1 0 3792 0 -1 5148
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220455
transform 1 0 1968 0 -1 5148
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220455
transform 1 0 3792 0 1 4972
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220455
transform 1 0 1968 0 1 4972
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220455
transform 1 0 3792 0 -1 4916
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220455
transform 1 0 1968 0 -1 4916
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220455
transform 1 0 3792 0 1 4712
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220455
transform 1 0 1968 0 1 4712
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220455
transform 1 0 3792 0 -1 4624
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220455
transform 1 0 1968 0 -1 4624
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220455
transform 1 0 3792 0 1 4448
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220455
transform 1 0 1968 0 1 4448
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220455
transform 1 0 3792 0 -1 4396
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220455
transform 1 0 1968 0 -1 4396
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220455
transform 1 0 3792 0 1 4212
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220455
transform 1 0 1968 0 1 4212
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220455
transform 1 0 3792 0 -1 4160
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220455
transform 1 0 1968 0 -1 4160
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220455
transform 1 0 3792 0 1 3984
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220455
transform 1 0 1968 0 1 3984
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220455
transform 1 0 3792 0 -1 3916
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220455
transform 1 0 1968 0 -1 3916
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220455
transform 1 0 3792 0 1 3728
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220455
transform 1 0 1968 0 1 3728
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220455
transform 1 0 3792 0 -1 3672
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220455
transform 1 0 1968 0 -1 3672
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220455
transform 1 0 3792 0 1 3484
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220455
transform 1 0 1968 0 1 3484
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220455
transform 1 0 3792 0 -1 3400
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220455
transform 1 0 1968 0 -1 3400
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220455
transform 1 0 3792 0 1 3224
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220455
transform 1 0 1968 0 1 3224
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220455
transform 1 0 3792 0 -1 3172
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220455
transform 1 0 1968 0 -1 3172
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220455
transform 1 0 3792 0 1 2976
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220455
transform 1 0 1968 0 1 2976
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220455
transform 1 0 3792 0 -1 2920
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220455
transform 1 0 1968 0 -1 2920
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220455
transform 1 0 3792 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220455
transform 1 0 1968 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220455
transform 1 0 3792 0 -1 2696
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220455
transform 1 0 1968 0 -1 2696
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220455
transform 1 0 3792 0 1 2520
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220455
transform 1 0 1968 0 1 2520
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220455
transform 1 0 3792 0 -1 2464
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220455
transform 1 0 1968 0 -1 2464
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220455
transform 1 0 3792 0 1 2280
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220455
transform 1 0 1968 0 1 2280
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220455
transform 1 0 3792 0 -1 2204
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220455
transform 1 0 1968 0 -1 2204
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220455
transform 1 0 3792 0 1 1996
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220455
transform 1 0 1968 0 1 1996
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220455
transform 1 0 3792 0 -1 1936
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220455
transform 1 0 1968 0 -1 1936
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220455
transform 1 0 3792 0 1 1760
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220455
transform 1 0 1968 0 1 1760
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220455
transform 1 0 3792 0 -1 1712
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220455
transform 1 0 1968 0 -1 1712
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220455
transform 1 0 3792 0 1 1536
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220455
transform 1 0 1968 0 1 1536
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220455
transform 1 0 3792 0 -1 1284
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220455
transform 1 0 1968 0 -1 1284
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220455
transform 1 0 3792 0 1 1096
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220455
transform 1 0 1968 0 1 1096
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220455
transform 1 0 3792 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220455
transform 1 0 1968 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220455
transform 1 0 3792 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220455
transform 1 0 1968 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220455
transform 1 0 3792 0 -1 812
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220455
transform 1 0 1968 0 -1 812
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220455
transform 1 0 3792 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220455
transform 1 0 1968 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220455
transform 1 0 3792 0 -1 560
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220455
transform 1 0 1968 0 -1 560
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220455
transform 1 0 3792 0 1 384
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220455
transform 1 0 1968 0 1 384
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220455
transform 1 0 3792 0 -1 332
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220455
transform 1 0 1968 0 -1 332
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220455
transform 1 0 3792 0 1 128
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220455
transform 1 0 1968 0 1 128
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220455
transform 1 0 1928 0 -1 5708
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220455
transform 1 0 104 0 -1 5708
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220455
transform 1 0 1928 0 1 5516
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220455
transform 1 0 104 0 1 5516
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220455
transform 1 0 1928 0 -1 5456
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220455
transform 1 0 104 0 -1 5456
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220455
transform 1 0 1928 0 1 5280
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220455
transform 1 0 104 0 1 5280
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220455
transform 1 0 1928 0 -1 5232
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220455
transform 1 0 104 0 -1 5232
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220455
transform 1 0 1928 0 1 5040
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220455
transform 1 0 104 0 1 5040
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220455
transform 1 0 1928 0 -1 4980
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220455
transform 1 0 104 0 -1 4980
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220455
transform 1 0 1928 0 1 4796
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220455
transform 1 0 104 0 1 4796
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220455
transform 1 0 1928 0 -1 4744
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220455
transform 1 0 104 0 -1 4744
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220455
transform 1 0 1928 0 1 4560
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220455
transform 1 0 104 0 1 4560
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220455
transform 1 0 1928 0 -1 4512
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220455
transform 1 0 104 0 -1 4512
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220455
transform 1 0 1928 0 1 4332
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220455
transform 1 0 104 0 1 4332
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220455
transform 1 0 1928 0 -1 4284
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220455
transform 1 0 104 0 -1 4284
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220455
transform 1 0 1928 0 1 4096
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220455
transform 1 0 104 0 1 4096
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220455
transform 1 0 1928 0 -1 4032
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220455
transform 1 0 104 0 -1 4032
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220455
transform 1 0 1928 0 1 3856
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220455
transform 1 0 104 0 1 3856
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220455
transform 1 0 1928 0 -1 3808
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220455
transform 1 0 104 0 -1 3808
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220455
transform 1 0 1928 0 1 3608
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220455
transform 1 0 104 0 1 3608
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220455
transform 1 0 1928 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220455
transform 1 0 104 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220455
transform 1 0 1928 0 1 3068
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220455
transform 1 0 104 0 1 3068
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220455
transform 1 0 1928 0 -1 3020
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220455
transform 1 0 104 0 -1 3020
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220455
transform 1 0 1928 0 1 2844
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220455
transform 1 0 104 0 1 2844
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220455
transform 1 0 1928 0 -1 2764
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220455
transform 1 0 104 0 -1 2764
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220455
transform 1 0 1928 0 1 2568
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220455
transform 1 0 104 0 1 2568
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220455
transform 1 0 1928 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220455
transform 1 0 104 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220455
transform 1 0 1928 0 1 2324
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220455
transform 1 0 104 0 1 2324
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220455
transform 1 0 1928 0 -1 2268
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220455
transform 1 0 104 0 -1 2268
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220455
transform 1 0 1928 0 1 2072
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220455
transform 1 0 104 0 1 2072
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220455
transform 1 0 1928 0 -1 2016
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220455
transform 1 0 104 0 -1 2016
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220455
transform 1 0 1928 0 1 1836
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220455
transform 1 0 104 0 1 1836
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220455
transform 1 0 1928 0 -1 1776
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220455
transform 1 0 104 0 -1 1776
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220455
transform 1 0 1928 0 1 1584
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220455
transform 1 0 104 0 1 1584
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220455
transform 1 0 1928 0 -1 1528
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220455
transform 1 0 104 0 -1 1528
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220455
transform 1 0 1928 0 1 1352
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220455
transform 1 0 104 0 1 1352
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220455
transform 1 0 1928 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220455
transform 1 0 104 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220455
transform 1 0 1928 0 1 1120
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220455
transform 1 0 104 0 1 1120
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220455
transform 1 0 1928 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220455
transform 1 0 104 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220455
transform 1 0 1928 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220455
transform 1 0 104 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220455
transform 1 0 1928 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220455
transform 1 0 104 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220455
transform 1 0 1928 0 1 604
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220455
transform 1 0 104 0 1 604
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220455
transform 1 0 1928 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220455
transform 1 0 104 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220455
transform 1 0 1928 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220455
transform 1 0 104 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220455
transform 1 0 1928 0 -1 320
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220455
transform 1 0 104 0 -1 320
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220455
transform 1 0 1928 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220455
transform 1 0 104 0 1 108
box 7 3 12 24
use _0_0std_0_0cells_0_0FAX1  tst_5999_6
timestamp 1731220455
transform 1 0 5512 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5998_6
timestamp 1731220455
transform 1 0 5376 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5997_6
timestamp 1731220455
transform 1 0 5512 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5996_6
timestamp 1731220455
transform 1 0 5352 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5995_6
timestamp 1731220455
transform 1 0 5168 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5994_6
timestamp 1731220455
transform 1 0 5240 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5993_6
timestamp 1731220455
transform 1 0 5104 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5992_6
timestamp 1731220455
transform 1 0 4968 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5991_6
timestamp 1731220455
transform 1 0 4832 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5990_6
timestamp 1731220455
transform 1 0 4696 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5989_6
timestamp 1731220455
transform 1 0 4560 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5988_6
timestamp 1731220455
transform 1 0 4424 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5987_6
timestamp 1731220455
transform 1 0 4288 0 1 108
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5986_6
timestamp 1731220455
transform 1 0 4984 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5985_6
timestamp 1731220455
transform 1 0 4792 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5984_6
timestamp 1731220455
transform 1 0 4584 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5983_6
timestamp 1731220455
transform 1 0 4352 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5982_6
timestamp 1731220455
transform 1 0 4104 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5981_6
timestamp 1731220455
transform 1 0 4920 0 1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5980_6
timestamp 1731220455
transform 1 0 4720 0 1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5979_6
timestamp 1731220455
transform 1 0 4520 0 1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5978_6
timestamp 1731220455
transform 1 0 4328 0 1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5977_6
timestamp 1731220455
transform 1 0 4496 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5976_6
timestamp 1731220455
transform 1 0 4656 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5975_6
timestamp 1731220455
transform 1 0 5080 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5974_6
timestamp 1731220455
transform 1 0 4944 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5973_6
timestamp 1731220455
transform 1 0 4808 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5972_6
timestamp 1731220455
transform 1 0 4808 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5971_6
timestamp 1731220455
transform 1 0 4672 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5970_6
timestamp 1731220455
transform 1 0 4536 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5969_6
timestamp 1731220455
transform 1 0 4400 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5968_6
timestamp 1731220455
transform 1 0 4336 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5967_6
timestamp 1731220455
transform 1 0 4176 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5966_6
timestamp 1731220455
transform 1 0 4016 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5965_6
timestamp 1731220455
transform 1 0 4128 0 1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5964_6
timestamp 1731220455
transform 1 0 3928 0 1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5963_6
timestamp 1731220455
transform 1 0 3856 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5962_6
timestamp 1731220455
transform 1 0 3648 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5961_6
timestamp 1731220455
transform 1 0 3648 0 1 104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5960_6
timestamp 1731220455
transform 1 0 3512 0 1 104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5959_6
timestamp 1731220455
transform 1 0 3352 0 1 104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5958_6
timestamp 1731220455
transform 1 0 3200 0 1 104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5957_6
timestamp 1731220455
transform 1 0 3048 0 1 104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5956_6
timestamp 1731220455
transform 1 0 2888 0 1 104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5955_6
timestamp 1731220455
transform 1 0 2720 0 1 104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5954_6
timestamp 1731220455
transform 1 0 2544 0 1 104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5953_6
timestamp 1731220455
transform 1 0 3376 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5952_6
timestamp 1731220455
transform 1 0 3088 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5951_6
timestamp 1731220455
transform 1 0 2816 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5950_6
timestamp 1731220455
transform 1 0 2744 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5949_6
timestamp 1731220455
transform 1 0 2600 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5948_6
timestamp 1731220455
transform 1 0 3032 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5947_6
timestamp 1731220455
transform 1 0 2888 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5946_6
timestamp 1731220455
transform 1 0 2856 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5945_6
timestamp 1731220455
transform 1 0 3032 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5944_6
timestamp 1731220455
transform 1 0 3200 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5943_6
timestamp 1731220455
transform 1 0 3552 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5942_6
timestamp 1731220455
transform 1 0 3376 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5941_6
timestamp 1731220455
transform 1 0 3320 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5940_6
timestamp 1731220455
transform 1 0 3648 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5939_6
timestamp 1731220455
transform 1 0 3856 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5938_6
timestamp 1731220455
transform 1 0 3992 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5937_6
timestamp 1731220455
transform 1 0 4264 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5936_6
timestamp 1731220455
transform 1 0 4128 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5935_6
timestamp 1731220455
transform 1 0 3992 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5934_6
timestamp 1731220455
transform 1 0 3856 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5933_6
timestamp 1731220455
transform 1 0 4128 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5932_6
timestamp 1731220455
transform 1 0 4264 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5931_6
timestamp 1731220455
transform 1 0 4672 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5930_6
timestamp 1731220455
transform 1 0 4536 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5929_6
timestamp 1731220455
transform 1 0 4400 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5928_6
timestamp 1731220455
transform 1 0 4288 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5927_6
timestamp 1731220455
transform 1 0 4152 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5926_6
timestamp 1731220455
transform 1 0 4016 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5925_6
timestamp 1731220455
transform 1 0 4696 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5924_6
timestamp 1731220455
transform 1 0 4560 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5923_6
timestamp 1731220455
transform 1 0 4424 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5922_6
timestamp 1731220455
transform 1 0 4336 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5921_6
timestamp 1731220455
transform 1 0 4472 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5920_6
timestamp 1731220455
transform 1 0 4608 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5919_6
timestamp 1731220455
transform 1 0 4880 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5918_6
timestamp 1731220455
transform 1 0 4744 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5917_6
timestamp 1731220455
transform 1 0 4696 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5916_6
timestamp 1731220455
transform 1 0 4560 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5915_6
timestamp 1731220455
transform 1 0 4424 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5914_6
timestamp 1731220455
transform 1 0 4440 0 -1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5913_6
timestamp 1731220455
transform 1 0 4144 0 -1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5912_6
timestamp 1731220455
transform 1 0 4720 0 -1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5911_6
timestamp 1731220455
transform 1 0 4704 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5910_6
timestamp 1731220455
transform 1 0 4872 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5909_6
timestamp 1731220455
transform 1 0 5040 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5908_6
timestamp 1731220455
transform 1 0 5200 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5907_6
timestamp 1731220455
transform 1 0 5256 0 -1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5906_6
timestamp 1731220455
transform 1 0 4992 0 -1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5905_6
timestamp 1731220455
transform 1 0 4968 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5904_6
timestamp 1731220455
transform 1 0 4832 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5903_6
timestamp 1731220455
transform 1 0 5104 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5902_6
timestamp 1731220455
transform 1 0 5240 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5901_6
timestamp 1731220455
transform 1 0 5376 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5900_6
timestamp 1731220455
transform 1 0 5512 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5899_6
timestamp 1731220455
transform 1 0 5512 0 -1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5898_6
timestamp 1731220455
transform 1 0 5368 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5897_6
timestamp 1731220455
transform 1 0 5512 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5896_6
timestamp 1731220455
transform 1 0 5512 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5895_6
timestamp 1731220455
transform 1 0 5512 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5894_6
timestamp 1731220455
transform 1 0 5512 0 -1 1808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5893_6
timestamp 1731220455
transform 1 0 5336 0 -1 1808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5892_6
timestamp 1731220455
transform 1 0 5408 0 1 1808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5891_6
timestamp 1731220455
transform 1 0 5144 0 -1 1808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5890_6
timestamp 1731220455
transform 1 0 4952 0 -1 1808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5889_6
timestamp 1731220455
transform 1 0 4968 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5888_6
timestamp 1731220455
transform 1 0 5152 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5887_6
timestamp 1731220455
transform 1 0 5336 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5886_6
timestamp 1731220455
transform 1 0 5352 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5885_6
timestamp 1731220455
transform 1 0 5176 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5884_6
timestamp 1731220455
transform 1 0 5000 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5883_6
timestamp 1731220455
transform 1 0 4832 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5882_6
timestamp 1731220455
transform 1 0 4664 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5881_6
timestamp 1731220455
transform 1 0 4496 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5880_6
timestamp 1731220455
transform 1 0 4784 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5879_6
timestamp 1731220455
transform 1 0 4600 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5878_6
timestamp 1731220455
transform 1 0 4544 0 -1 1808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5877_6
timestamp 1731220455
transform 1 0 4336 0 -1 1808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5876_6
timestamp 1731220455
transform 1 0 4752 0 -1 1808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5875_6
timestamp 1731220455
transform 1 0 5088 0 1 1808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5874_6
timestamp 1731220455
transform 1 0 4768 0 1 1808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5873_6
timestamp 1731220455
transform 1 0 4464 0 1 1808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5872_6
timestamp 1731220455
transform 1 0 4192 0 1 1808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5871_6
timestamp 1731220455
transform 1 0 3952 0 1 1808
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5870_6
timestamp 1731220455
transform 1 0 4256 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5869_6
timestamp 1731220455
transform 1 0 4392 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5868_6
timestamp 1731220455
transform 1 0 4528 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5867_6
timestamp 1731220455
transform 1 0 4664 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5866_6
timestamp 1731220455
transform 1 0 4808 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5865_6
timestamp 1731220455
transform 1 0 4656 0 1 2072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5864_6
timestamp 1731220455
transform 1 0 4848 0 1 2072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5863_6
timestamp 1731220455
transform 1 0 5032 0 1 2072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5862_6
timestamp 1731220455
transform 1 0 5216 0 1 2072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5861_6
timestamp 1731220455
transform 1 0 5408 0 1 2072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5860_6
timestamp 1731220455
transform 1 0 5328 0 -1 2296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5859_6
timestamp 1731220455
transform 1 0 5504 0 -1 2296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5858_6
timestamp 1731220455
transform 1 0 5512 0 1 2316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5857_6
timestamp 1731220455
transform 1 0 5512 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5856_6
timestamp 1731220455
transform 1 0 5512 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5855_6
timestamp 1731220455
transform 1 0 5512 0 -1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5854_6
timestamp 1731220455
transform 1 0 5512 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5853_6
timestamp 1731220455
transform 1 0 5504 0 -1 3020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5852_6
timestamp 1731220455
transform 1 0 5512 0 1 3020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5851_6
timestamp 1731220455
transform 1 0 5376 0 1 3020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5850_6
timestamp 1731220455
transform 1 0 5216 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5849_6
timestamp 1731220455
transform 1 0 5200 0 -1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5848_6
timestamp 1731220455
transform 1 0 5272 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5847_6
timestamp 1731220455
transform 1 0 5320 0 1 2316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5846_6
timestamp 1731220455
transform 1 0 5136 0 1 2316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5845_6
timestamp 1731220455
transform 1 0 5152 0 -1 2296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5844_6
timestamp 1731220455
transform 1 0 4984 0 -1 2296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5843_6
timestamp 1731220455
transform 1 0 4808 0 -1 2296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5842_6
timestamp 1731220455
transform 1 0 4624 0 -1 2296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5841_6
timestamp 1731220455
transform 1 0 4432 0 -1 2296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5840_6
timestamp 1731220455
transform 1 0 4960 0 1 2316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5839_6
timestamp 1731220455
transform 1 0 4792 0 1 2316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5838_6
timestamp 1731220455
transform 1 0 4632 0 1 2316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5837_6
timestamp 1731220455
transform 1 0 4488 0 1 2316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5836_6
timestamp 1731220455
transform 1 0 5016 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5835_6
timestamp 1731220455
transform 1 0 4768 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5834_6
timestamp 1731220455
transform 1 0 4528 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5833_6
timestamp 1731220455
transform 1 0 4304 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5832_6
timestamp 1731220455
transform 1 0 5200 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5831_6
timestamp 1731220455
transform 1 0 4864 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5830_6
timestamp 1731220455
transform 1 0 4552 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5829_6
timestamp 1731220455
transform 1 0 4272 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5828_6
timestamp 1731220455
transform 1 0 4024 0 1 2560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5827_6
timestamp 1731220455
transform 1 0 4864 0 -1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5826_6
timestamp 1731220455
transform 1 0 4536 0 -1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5825_6
timestamp 1731220455
transform 1 0 4224 0 -1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5824_6
timestamp 1731220455
transform 1 0 3936 0 -1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5823_6
timestamp 1731220455
transform 1 0 4032 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5822_6
timestamp 1731220455
transform 1 0 4312 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5821_6
timestamp 1731220455
transform 1 0 4600 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5820_6
timestamp 1731220455
transform 1 0 4904 0 1 2796
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5819_6
timestamp 1731220455
transform 1 0 4752 0 -1 3020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5818_6
timestamp 1731220455
transform 1 0 4536 0 -1 3020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5817_6
timestamp 1731220455
transform 1 0 4336 0 -1 3020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5816_6
timestamp 1731220455
transform 1 0 5248 0 -1 3020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5815_6
timestamp 1731220455
transform 1 0 4992 0 -1 3020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5814_6
timestamp 1731220455
transform 1 0 4832 0 1 3020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5813_6
timestamp 1731220455
transform 1 0 4696 0 1 3020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5812_6
timestamp 1731220455
transform 1 0 4968 0 1 3020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5811_6
timestamp 1731220455
transform 1 0 5104 0 1 3020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5810_6
timestamp 1731220455
transform 1 0 5240 0 1 3020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5809_6
timestamp 1731220455
transform 1 0 5320 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5808_6
timestamp 1731220455
transform 1 0 5184 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5807_6
timestamp 1731220455
transform 1 0 5048 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5806_6
timestamp 1731220455
transform 1 0 4912 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5805_6
timestamp 1731220455
transform 1 0 4776 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5804_6
timestamp 1731220455
transform 1 0 4944 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5803_6
timestamp 1731220455
transform 1 0 4784 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5802_6
timestamp 1731220455
transform 1 0 4624 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5801_6
timestamp 1731220455
transform 1 0 4464 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5800_6
timestamp 1731220455
transform 1 0 4312 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5799_6
timestamp 1731220455
transform 1 0 5352 0 -1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5798_6
timestamp 1731220455
transform 1 0 5216 0 -1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5797_6
timestamp 1731220455
transform 1 0 5080 0 -1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5796_6
timestamp 1731220455
transform 1 0 4944 0 -1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5795_6
timestamp 1731220455
transform 1 0 4808 0 -1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5794_6
timestamp 1731220455
transform 1 0 4672 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5793_6
timestamp 1731220455
transform 1 0 4536 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5792_6
timestamp 1731220455
transform 1 0 4400 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5791_6
timestamp 1731220455
transform 1 0 4808 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5790_6
timestamp 1731220455
transform 1 0 4944 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5789_6
timestamp 1731220455
transform 1 0 5160 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5788_6
timestamp 1731220455
transform 1 0 4904 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5787_6
timestamp 1731220455
transform 1 0 4664 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5786_6
timestamp 1731220455
transform 1 0 4440 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5785_6
timestamp 1731220455
transform 1 0 4240 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5784_6
timestamp 1731220455
transform 1 0 4496 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5783_6
timestamp 1731220455
transform 1 0 4672 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5782_6
timestamp 1731220455
transform 1 0 4872 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5781_6
timestamp 1731220455
transform 1 0 5312 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5780_6
timestamp 1731220455
transform 1 0 5088 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5779_6
timestamp 1731220455
transform 1 0 5080 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5778_6
timestamp 1731220455
transform 1 0 4936 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5777_6
timestamp 1731220455
transform 1 0 4800 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5776_6
timestamp 1731220455
transform 1 0 5224 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5775_6
timestamp 1731220455
transform 1 0 5376 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5774_6
timestamp 1731220455
transform 1 0 5344 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5773_6
timestamp 1731220455
transform 1 0 5208 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5772_6
timestamp 1731220455
transform 1 0 5072 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5771_6
timestamp 1731220455
transform 1 0 4936 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5770_6
timestamp 1731220455
transform 1 0 5192 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5769_6
timestamp 1731220455
transform 1 0 5056 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5768_6
timestamp 1731220455
transform 1 0 4920 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5767_6
timestamp 1731220455
transform 1 0 4784 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5766_6
timestamp 1731220455
transform 1 0 5064 0 1 4244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5765_6
timestamp 1731220455
transform 1 0 4872 0 1 4244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5764_6
timestamp 1731220455
transform 1 0 4688 0 1 4244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5763_6
timestamp 1731220455
transform 1 0 4512 0 1 4244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5762_6
timestamp 1731220455
transform 1 0 4992 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5761_6
timestamp 1731220455
transform 1 0 4744 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5760_6
timestamp 1731220455
transform 1 0 4504 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5759_6
timestamp 1731220455
transform 1 0 4280 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5758_6
timestamp 1731220455
transform 1 0 4624 0 1 4504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5757_6
timestamp 1731220455
transform 1 0 4328 0 1 4504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5756_6
timestamp 1731220455
transform 1 0 4032 0 1 4504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5755_6
timestamp 1731220455
transform 1 0 4088 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5754_6
timestamp 1731220455
transform 1 0 4344 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5753_6
timestamp 1731220455
transform 1 0 4616 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5752_6
timestamp 1731220455
transform 1 0 4912 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5751_6
timestamp 1731220455
transform 1 0 4872 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5750_6
timestamp 1731220455
transform 1 0 4672 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5749_6
timestamp 1731220455
transform 1 0 4480 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5748_6
timestamp 1731220455
transform 1 0 5088 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5747_6
timestamp 1731220455
transform 1 0 5224 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5746_6
timestamp 1731220455
transform 1 0 4928 0 1 4504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5745_6
timestamp 1731220455
transform 1 0 5232 0 1 4504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5744_6
timestamp 1731220455
transform 1 0 5248 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5743_6
timestamp 1731220455
transform 1 0 5264 0 1 4244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5742_6
timestamp 1731220455
transform 1 0 5328 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5741_6
timestamp 1731220455
transform 1 0 5480 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5740_6
timestamp 1731220455
transform 1 0 5416 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5739_6
timestamp 1731220455
transform 1 0 5488 0 -1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5738_6
timestamp 1731220455
transform 1 0 5512 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5737_6
timestamp 1731220455
transform 1 0 5512 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5736_6
timestamp 1731220455
transform 1 0 5464 0 -1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5735_6
timestamp 1731220455
transform 1 0 5464 0 1 4244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5734_6
timestamp 1731220455
transform 1 0 5512 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5733_6
timestamp 1731220455
transform 1 0 5512 0 1 4504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5732_6
timestamp 1731220455
transform 1 0 5512 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5731_6
timestamp 1731220455
transform 1 0 5512 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5730_6
timestamp 1731220455
transform 1 0 5512 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5729_6
timestamp 1731220455
transform 1 0 5512 0 1 5020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5728_6
timestamp 1731220455
transform 1 0 5464 0 -1 5244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5727_6
timestamp 1731220455
transform 1 0 5416 0 1 5272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5726_6
timestamp 1731220455
transform 1 0 5376 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5725_6
timestamp 1731220455
transform 1 0 5240 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5724_6
timestamp 1731220455
transform 1 0 5312 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5723_6
timestamp 1731220455
transform 1 0 5104 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5722_6
timestamp 1731220455
transform 1 0 4968 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5721_6
timestamp 1731220455
transform 1 0 4832 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5720_6
timestamp 1731220455
transform 1 0 4880 0 1 5020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5719_6
timestamp 1731220455
transform 1 0 5192 0 1 5020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5718_6
timestamp 1731220455
transform 1 0 5120 0 -1 5244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5717_6
timestamp 1731220455
transform 1 0 5288 0 -1 5244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5716_6
timestamp 1731220455
transform 1 0 5168 0 1 5272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5715_6
timestamp 1731220455
transform 1 0 4928 0 1 5272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5714_6
timestamp 1731220455
transform 1 0 4832 0 -1 5496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5713_6
timestamp 1731220455
transform 1 0 4696 0 -1 5496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5712_6
timestamp 1731220455
transform 1 0 5056 0 1 5496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5711_6
timestamp 1731220455
transform 1 0 4920 0 1 5496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5710_6
timestamp 1731220455
transform 1 0 4784 0 1 5496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5709_6
timestamp 1731220455
transform 1 0 4648 0 1 5496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5708_6
timestamp 1731220455
transform 1 0 4512 0 1 5496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5707_6
timestamp 1731220455
transform 1 0 4376 0 1 5496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5706_6
timestamp 1731220455
transform 1 0 4240 0 1 5496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5705_6
timestamp 1731220455
transform 1 0 4424 0 -1 5496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5704_6
timestamp 1731220455
transform 1 0 4560 0 -1 5496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5703_6
timestamp 1731220455
transform 1 0 4480 0 1 5272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5702_6
timestamp 1731220455
transform 1 0 4280 0 1 5272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5701_6
timestamp 1731220455
transform 1 0 4696 0 1 5272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5700_6
timestamp 1731220455
transform 1 0 4960 0 -1 5244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5699_6
timestamp 1731220455
transform 1 0 4808 0 -1 5244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5698_6
timestamp 1731220455
transform 1 0 4672 0 -1 5244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5697_6
timestamp 1731220455
transform 1 0 4576 0 1 5020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5696_6
timestamp 1731220455
transform 1 0 4272 0 1 5020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5695_6
timestamp 1731220455
transform 1 0 3976 0 1 5020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5694_6
timestamp 1731220455
transform 1 0 4536 0 -1 5244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5693_6
timestamp 1731220455
transform 1 0 4400 0 -1 5244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5692_6
timestamp 1731220455
transform 1 0 4264 0 -1 5244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5691_6
timestamp 1731220455
transform 1 0 4128 0 -1 5244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5690_6
timestamp 1731220455
transform 1 0 3992 0 -1 5244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5689_6
timestamp 1731220455
transform 1 0 3856 0 -1 5244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5688_6
timestamp 1731220455
transform 1 0 3648 0 -1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5687_6
timestamp 1731220455
transform 1 0 3512 0 -1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5686_6
timestamp 1731220455
transform 1 0 3648 0 1 4948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5685_6
timestamp 1731220455
transform 1 0 3512 0 1 4948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5684_6
timestamp 1731220455
transform 1 0 3376 0 1 4948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5683_6
timestamp 1731220455
transform 1 0 3240 0 1 4948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5682_6
timestamp 1731220455
transform 1 0 3104 0 1 4948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5681_6
timestamp 1731220455
transform 1 0 3104 0 -1 4940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5680_6
timestamp 1731220455
transform 1 0 3240 0 -1 4940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5679_6
timestamp 1731220455
transform 1 0 3648 0 -1 4940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5678_6
timestamp 1731220455
transform 1 0 3512 0 -1 4940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5677_6
timestamp 1731220455
transform 1 0 3376 0 -1 4940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5676_6
timestamp 1731220455
transform 1 0 3240 0 1 4688
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5675_6
timestamp 1731220455
transform 1 0 3104 0 1 4688
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5674_6
timestamp 1731220455
transform 1 0 3376 0 1 4688
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5673_6
timestamp 1731220455
transform 1 0 3512 0 1 4688
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5672_6
timestamp 1731220455
transform 1 0 3648 0 1 4688
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5671_6
timestamp 1731220455
transform 1 0 3648 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5670_6
timestamp 1731220455
transform 1 0 3496 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5669_6
timestamp 1731220455
transform 1 0 3320 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5668_6
timestamp 1731220455
transform 1 0 3152 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5667_6
timestamp 1731220455
transform 1 0 2976 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5666_6
timestamp 1731220455
transform 1 0 3576 0 1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5665_6
timestamp 1731220455
transform 1 0 3352 0 1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5664_6
timestamp 1731220455
transform 1 0 3128 0 1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5663_6
timestamp 1731220455
transform 1 0 2912 0 1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5662_6
timestamp 1731220455
transform 1 0 3376 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5661_6
timestamp 1731220455
transform 1 0 3168 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5660_6
timestamp 1731220455
transform 1 0 2960 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5659_6
timestamp 1731220455
transform 1 0 2752 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5658_6
timestamp 1731220455
transform 1 0 2664 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5657_6
timestamp 1731220455
transform 1 0 2872 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5656_6
timestamp 1731220455
transform 1 0 3288 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5655_6
timestamp 1731220455
transform 1 0 3080 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5654_6
timestamp 1731220455
transform 1 0 3008 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5653_6
timestamp 1731220455
transform 1 0 2768 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5652_6
timestamp 1731220455
transform 1 0 2520 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5651_6
timestamp 1731220455
transform 1 0 3248 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5650_6
timestamp 1731220455
transform 1 0 3488 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5649_6
timestamp 1731220455
transform 1 0 3448 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5648_6
timestamp 1731220455
transform 1 0 3160 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5647_6
timestamp 1731220455
transform 1 0 2872 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5646_6
timestamp 1731220455
transform 1 0 2584 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5645_6
timestamp 1731220455
transform 1 0 2280 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5644_6
timestamp 1731220455
transform 1 0 3184 0 -1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5643_6
timestamp 1731220455
transform 1 0 3048 0 -1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5642_6
timestamp 1731220455
transform 1 0 2912 0 -1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5641_6
timestamp 1731220455
transform 1 0 2776 0 -1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5640_6
timestamp 1731220455
transform 1 0 2640 0 -1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5639_6
timestamp 1731220455
transform 1 0 2760 0 1 3704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5638_6
timestamp 1731220455
transform 1 0 2920 0 1 3704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5637_6
timestamp 1731220455
transform 1 0 3080 0 1 3704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5636_6
timestamp 1731220455
transform 1 0 3240 0 1 3704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5635_6
timestamp 1731220455
transform 1 0 3408 0 1 3704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5634_6
timestamp 1731220455
transform 1 0 3304 0 -1 3696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5633_6
timestamp 1731220455
transform 1 0 3120 0 -1 3696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5632_6
timestamp 1731220455
transform 1 0 2936 0 -1 3696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5631_6
timestamp 1731220455
transform 1 0 3488 0 -1 3696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5630_6
timestamp 1731220455
transform 1 0 3648 0 -1 3696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5629_6
timestamp 1731220455
transform 1 0 3856 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5628_6
timestamp 1731220455
transform 1 0 3992 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5627_6
timestamp 1731220455
transform 1 0 4128 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5626_6
timestamp 1731220455
transform 1 0 4264 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5625_6
timestamp 1731220455
transform 1 0 4264 0 -1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5624_6
timestamp 1731220455
transform 1 0 4672 0 -1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5623_6
timestamp 1731220455
transform 1 0 4536 0 -1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5622_6
timestamp 1731220455
transform 1 0 4400 0 -1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5621_6
timestamp 1731220455
transform 1 0 4128 0 -1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5620_6
timestamp 1731220455
transform 1 0 3992 0 -1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5619_6
timestamp 1731220455
transform 1 0 3856 0 -1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5618_6
timestamp 1731220455
transform 1 0 4152 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5617_6
timestamp 1731220455
transform 1 0 3992 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5616_6
timestamp 1731220455
transform 1 0 3856 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5615_6
timestamp 1731220455
transform 1 0 3648 0 1 3200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5614_6
timestamp 1731220455
transform 1 0 3424 0 1 3200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5613_6
timestamp 1731220455
transform 1 0 3648 0 -1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5612_6
timestamp 1731220455
transform 1 0 3472 0 -1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5611_6
timestamp 1731220455
transform 1 0 3400 0 1 2952
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5610_6
timestamp 1731220455
transform 1 0 3600 0 1 2952
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5609_6
timestamp 1731220455
transform 1 0 3640 0 -1 2944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5608_6
timestamp 1731220455
transform 1 0 3496 0 -1 2944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5607_6
timestamp 1731220455
transform 1 0 3360 0 -1 2944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5606_6
timestamp 1731220455
transform 1 0 3224 0 -1 2944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5605_6
timestamp 1731220455
transform 1 0 3088 0 -1 2944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5604_6
timestamp 1731220455
transform 1 0 3000 0 1 2952
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5603_6
timestamp 1731220455
transform 1 0 3200 0 1 2952
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5602_6
timestamp 1731220455
transform 1 0 3280 0 -1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5601_6
timestamp 1731220455
transform 1 0 3096 0 -1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5600_6
timestamp 1731220455
transform 1 0 2920 0 -1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5599_6
timestamp 1731220455
transform 1 0 2952 0 1 3200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5598_6
timestamp 1731220455
transform 1 0 3184 0 1 3200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5597_6
timestamp 1731220455
transform 1 0 2952 0 -1 3424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5596_6
timestamp 1731220455
transform 1 0 2544 0 -1 3424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5595_6
timestamp 1731220455
transform 1 0 2408 0 -1 3424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5594_6
timestamp 1731220455
transform 1 0 2272 0 -1 3424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5593_6
timestamp 1731220455
transform 1 0 2136 0 -1 3424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5592_6
timestamp 1731220455
transform 1 0 2536 0 1 3200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5591_6
timestamp 1731220455
transform 1 0 2360 0 1 3200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5590_6
timestamp 1731220455
transform 1 0 2200 0 1 3200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5589_6
timestamp 1731220455
transform 1 0 2056 0 1 3200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5588_6
timestamp 1731220455
transform 1 0 2424 0 -1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5587_6
timestamp 1731220455
transform 1 0 2272 0 -1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5586_6
timestamp 1731220455
transform 1 0 2128 0 -1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5585_6
timestamp 1731220455
transform 1 0 1992 0 -1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5584_6
timestamp 1731220455
transform 1 0 1784 0 1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5583_6
timestamp 1731220455
transform 1 0 1592 0 1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5582_6
timestamp 1731220455
transform 1 0 1504 0 -1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5581_6
timestamp 1731220455
transform 1 0 1648 0 -1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5580_6
timestamp 1731220455
transform 1 0 1784 0 -1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5579_6
timestamp 1731220455
transform 1 0 1784 0 1 2820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5578_6
timestamp 1731220455
transform 1 0 1608 0 1 2820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5577_6
timestamp 1731220455
transform 1 0 1408 0 1 2820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5576_6
timestamp 1731220455
transform 1 0 1216 0 1 2820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5575_6
timestamp 1731220455
transform 1 0 1016 0 1 2820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5574_6
timestamp 1731220455
transform 1 0 1360 0 -1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5573_6
timestamp 1731220455
transform 1 0 1216 0 -1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5572_6
timestamp 1731220455
transform 1 0 1072 0 -1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5571_6
timestamp 1731220455
transform 1 0 928 0 -1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5570_6
timestamp 1731220455
transform 1 0 776 0 -1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5569_6
timestamp 1731220455
transform 1 0 616 0 -1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5568_6
timestamp 1731220455
transform 1 0 1384 0 1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5567_6
timestamp 1731220455
transform 1 0 1184 0 1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5566_6
timestamp 1731220455
transform 1 0 992 0 1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5565_6
timestamp 1731220455
transform 1 0 808 0 1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5564_6
timestamp 1731220455
transform 1 0 1488 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5563_6
timestamp 1731220455
transform 1 0 1352 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5562_6
timestamp 1731220455
transform 1 0 1216 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5561_6
timestamp 1731220455
transform 1 0 1080 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5560_6
timestamp 1731220455
transform 1 0 944 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5559_6
timestamp 1731220455
transform 1 0 808 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5558_6
timestamp 1731220455
transform 1 0 672 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5557_6
timestamp 1731220455
transform 1 0 536 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5556_6
timestamp 1731220455
transform 1 0 400 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5555_6
timestamp 1731220455
transform 1 0 264 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5554_6
timestamp 1731220455
transform 1 0 128 0 -1 3296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5553_6
timestamp 1731220455
transform 1 0 288 0 1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5552_6
timestamp 1731220455
transform 1 0 456 0 1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5551_6
timestamp 1731220455
transform 1 0 624 0 1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5550_6
timestamp 1731220455
transform 1 0 456 0 -1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5549_6
timestamp 1731220455
transform 1 0 296 0 -1 3044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5548_6
timestamp 1731220455
transform 1 0 152 0 1 2820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5547_6
timestamp 1731220455
transform 1 0 376 0 1 2820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5546_6
timestamp 1731220455
transform 1 0 592 0 1 2820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5545_6
timestamp 1731220455
transform 1 0 808 0 1 2820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5544_6
timestamp 1731220455
transform 1 0 800 0 -1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5543_6
timestamp 1731220455
transform 1 0 664 0 -1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5542_6
timestamp 1731220455
transform 1 0 528 0 -1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5541_6
timestamp 1731220455
transform 1 0 392 0 -1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5540_6
timestamp 1731220455
transform 1 0 256 0 -1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5539_6
timestamp 1731220455
transform 1 0 536 0 1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5538_6
timestamp 1731220455
transform 1 0 696 0 1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5537_6
timestamp 1731220455
transform 1 0 880 0 1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5536_6
timestamp 1731220455
transform 1 0 1088 0 1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5535_6
timestamp 1731220455
transform 1 0 1560 0 1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5534_6
timestamp 1731220455
transform 1 0 1320 0 1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5533_6
timestamp 1731220455
transform 1 0 1296 0 -1 2532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5532_6
timestamp 1731220455
transform 1 0 1128 0 -1 2532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5531_6
timestamp 1731220455
transform 1 0 968 0 -1 2532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5530_6
timestamp 1731220455
transform 1 0 816 0 -1 2532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5529_6
timestamp 1731220455
transform 1 0 664 0 -1 2532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5528_6
timestamp 1731220455
transform 1 0 1264 0 1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5527_6
timestamp 1731220455
transform 1 0 1056 0 1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5526_6
timestamp 1731220455
transform 1 0 856 0 1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5525_6
timestamp 1731220455
transform 1 0 672 0 1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5524_6
timestamp 1731220455
transform 1 0 504 0 1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5523_6
timestamp 1731220455
transform 1 0 352 0 1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5522_6
timestamp 1731220455
transform 1 0 944 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5521_6
timestamp 1731220455
transform 1 0 728 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5520_6
timestamp 1731220455
transform 1 0 512 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5519_6
timestamp 1731220455
transform 1 0 304 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5518_6
timestamp 1731220455
transform 1 0 128 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5517_6
timestamp 1731220455
transform 1 0 928 0 1 2048
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5516_6
timestamp 1731220455
transform 1 0 712 0 1 2048
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5515_6
timestamp 1731220455
transform 1 0 496 0 1 2048
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5514_6
timestamp 1731220455
transform 1 0 296 0 1 2048
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5513_6
timestamp 1731220455
transform 1 0 128 0 1 2048
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5512_6
timestamp 1731220455
transform 1 0 128 0 -1 2040
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5511_6
timestamp 1731220455
transform 1 0 312 0 -1 2040
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5510_6
timestamp 1731220455
transform 1 0 536 0 -1 2040
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5509_6
timestamp 1731220455
transform 1 0 1032 0 -1 2040
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5508_6
timestamp 1731220455
transform 1 0 776 0 -1 2040
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5507_6
timestamp 1731220455
transform 1 0 664 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5506_6
timestamp 1731220455
transform 1 0 496 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5505_6
timestamp 1731220455
transform 1 0 328 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5504_6
timestamp 1731220455
transform 1 0 840 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5503_6
timestamp 1731220455
transform 1 0 1024 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5502_6
timestamp 1731220455
transform 1 0 984 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5501_6
timestamp 1731220455
transform 1 0 824 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5500_6
timestamp 1731220455
transform 1 0 664 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5499_6
timestamp 1731220455
transform 1 0 504 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5498_6
timestamp 1731220455
transform 1 0 800 0 1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5497_6
timestamp 1731220455
transform 1 0 608 0 1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5496_6
timestamp 1731220455
transform 1 0 424 0 1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5495_6
timestamp 1731220455
transform 1 0 328 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5494_6
timestamp 1731220455
transform 1 0 600 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5493_6
timestamp 1731220455
transform 1 0 496 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5492_6
timestamp 1731220455
transform 1 0 304 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5491_6
timestamp 1731220455
transform 1 0 128 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5490_6
timestamp 1731220455
transform 1 0 128 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5489_6
timestamp 1731220455
transform 1 0 344 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5488_6
timestamp 1731220455
transform 1 0 344 0 1 1096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5487_6
timestamp 1731220455
transform 1 0 128 0 1 1096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5486_6
timestamp 1731220455
transform 1 0 560 0 1 1096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5485_6
timestamp 1731220455
transform 1 0 440 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5484_6
timestamp 1731220455
transform 1 0 576 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5483_6
timestamp 1731220455
transform 1 0 528 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5482_6
timestamp 1731220455
transform 1 0 392 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5481_6
timestamp 1731220455
transform 1 0 256 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5480_6
timestamp 1731220455
transform 1 0 208 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5479_6
timestamp 1731220455
transform 1 0 408 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5478_6
timestamp 1731220455
transform 1 0 584 0 1 580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5477_6
timestamp 1731220455
transform 1 0 344 0 1 580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5476_6
timestamp 1731220455
transform 1 0 128 0 1 580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5475_6
timestamp 1731220455
transform 1 0 128 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5474_6
timestamp 1731220455
transform 1 0 376 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5473_6
timestamp 1731220455
transform 1 0 192 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5472_6
timestamp 1731220455
transform 1 0 424 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5471_6
timestamp 1731220455
transform 1 0 320 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5470_6
timestamp 1731220455
transform 1 0 264 0 1 84
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5469_6
timestamp 1731220455
transform 1 0 128 0 1 84
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5468_6
timestamp 1731220455
transform 1 0 400 0 1 84
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5467_6
timestamp 1731220455
transform 1 0 536 0 1 84
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5466_6
timestamp 1731220455
transform 1 0 672 0 1 84
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5465_6
timestamp 1731220455
transform 1 0 1080 0 1 84
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5464_6
timestamp 1731220455
transform 1 0 944 0 1 84
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5463_6
timestamp 1731220455
transform 1 0 808 0 1 84
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5462_6
timestamp 1731220455
transform 1 0 768 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5461_6
timestamp 1731220455
transform 1 0 544 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5460_6
timestamp 1731220455
transform 1 0 880 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5459_6
timestamp 1731220455
transform 1 0 656 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5458_6
timestamp 1731220455
transform 1 0 640 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5457_6
timestamp 1731220455
transform 1 0 904 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5456_6
timestamp 1731220455
transform 1 0 1160 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5455_6
timestamp 1731220455
transform 1 0 1312 0 1 580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5454_6
timestamp 1731220455
transform 1 0 1064 0 1 580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5453_6
timestamp 1731220455
transform 1 0 824 0 1 580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5452_6
timestamp 1731220455
transform 1 0 824 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5451_6
timestamp 1731220455
transform 1 0 616 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5450_6
timestamp 1731220455
transform 1 0 1032 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5449_6
timestamp 1731220455
transform 1 0 936 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5448_6
timestamp 1731220455
transform 1 0 800 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5447_6
timestamp 1731220455
transform 1 0 664 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5446_6
timestamp 1731220455
transform 1 0 712 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5445_6
timestamp 1731220455
transform 1 0 856 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5444_6
timestamp 1731220455
transform 1 0 1000 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5443_6
timestamp 1731220455
transform 1 0 1192 0 1 1096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5442_6
timestamp 1731220455
transform 1 0 984 0 1 1096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5441_6
timestamp 1731220455
transform 1 0 776 0 1 1096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5440_6
timestamp 1731220455
transform 1 0 568 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5439_6
timestamp 1731220455
transform 1 0 776 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5438_6
timestamp 1731220455
transform 1 0 968 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5437_6
timestamp 1731220455
transform 1 0 1024 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5436_6
timestamp 1731220455
transform 1 0 856 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5435_6
timestamp 1731220455
transform 1 0 680 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5434_6
timestamp 1731220455
transform 1 0 856 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5433_6
timestamp 1731220455
transform 1 0 1104 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5432_6
timestamp 1731220455
transform 1 0 992 0 1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5431_6
timestamp 1731220455
transform 1 0 1184 0 1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5430_6
timestamp 1731220455
transform 1 0 1376 0 1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5429_6
timestamp 1731220455
transform 1 0 1320 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5428_6
timestamp 1731220455
transform 1 0 1152 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5427_6
timestamp 1731220455
transform 1 0 1488 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5426_6
timestamp 1731220455
transform 1 0 1408 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5425_6
timestamp 1731220455
transform 1 0 1216 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5424_6
timestamp 1731220455
transform 1 0 1600 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5423_6
timestamp 1731220455
transform 1 0 1576 0 -1 2040
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5422_6
timestamp 1731220455
transform 1 0 1304 0 -1 2040
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5421_6
timestamp 1731220455
transform 1 0 1624 0 1 2048
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5420_6
timestamp 1731220455
transform 1 0 1384 0 1 2048
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5419_6
timestamp 1731220455
transform 1 0 1152 0 1 2048
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5418_6
timestamp 1731220455
transform 1 0 1168 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5417_6
timestamp 1731220455
transform 1 0 1400 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5416_6
timestamp 1731220455
transform 1 0 1640 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5415_6
timestamp 1731220455
transform 1 0 1696 0 1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5414_6
timestamp 1731220455
transform 1 0 1480 0 1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5413_6
timestamp 1731220455
transform 1 0 1464 0 -1 2532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5412_6
timestamp 1731220455
transform 1 0 1632 0 -1 2532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5411_6
timestamp 1731220455
transform 1 0 1784 0 -1 2532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5410_6
timestamp 1731220455
transform 1 0 1784 0 1 2544
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5409_6
timestamp 1731220455
transform 1 0 1992 0 1 2496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5408_6
timestamp 1731220455
transform 1 0 1992 0 -1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5407_6
timestamp 1731220455
transform 1 0 2264 0 -1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5406_6
timestamp 1731220455
transform 1 0 2128 0 -1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5405_6
timestamp 1731220455
transform 1 0 2008 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5404_6
timestamp 1731220455
transform 1 0 2248 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5403_6
timestamp 1731220455
transform 1 0 2400 0 -1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5402_6
timestamp 1731220455
transform 1 0 2672 0 -1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5401_6
timestamp 1731220455
transform 1 0 2536 0 -1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5400_6
timestamp 1731220455
transform 1 0 2416 0 1 2496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5399_6
timestamp 1731220455
transform 1 0 2200 0 1 2496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5398_6
timestamp 1731220455
transform 1 0 2288 0 -1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5397_6
timestamp 1731220455
transform 1 0 2536 0 -1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5396_6
timestamp 1731220455
transform 1 0 2536 0 1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5395_6
timestamp 1731220455
transform 1 0 2328 0 1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5394_6
timestamp 1731220455
transform 1 0 2736 0 1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5393_6
timestamp 1731220455
transform 1 0 2704 0 -1 2228
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5392_6
timestamp 1731220455
transform 1 0 2568 0 -1 2228
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5391_6
timestamp 1731220455
transform 1 0 2432 0 -1 2228
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5390_6
timestamp 1731220455
transform 1 0 2416 0 1 1972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5389_6
timestamp 1731220455
transform 1 0 2792 0 1 1972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5388_6
timestamp 1731220455
transform 1 0 2608 0 1 1972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5387_6
timestamp 1731220455
transform 1 0 2600 0 -1 1960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5386_6
timestamp 1731220455
transform 1 0 2464 0 -1 1960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5385_6
timestamp 1731220455
transform 1 0 2328 0 -1 1960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5384_6
timestamp 1731220455
transform 1 0 2208 0 1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5383_6
timestamp 1731220455
transform 1 0 2352 0 1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5382_6
timestamp 1731220455
transform 1 0 2496 0 1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5381_6
timestamp 1731220455
transform 1 0 2568 0 -1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5380_6
timestamp 1731220455
transform 1 0 2376 0 -1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5379_6
timestamp 1731220455
transform 1 0 2184 0 -1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5378_6
timestamp 1731220455
transform 1 0 1992 0 -1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5377_6
timestamp 1731220455
transform 1 0 2800 0 1 1512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5376_6
timestamp 1731220455
transform 1 0 2584 0 1 1512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5375_6
timestamp 1731220455
transform 1 0 2368 0 1 1512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5374_6
timestamp 1731220455
transform 1 0 2160 0 1 1512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5373_6
timestamp 1731220455
transform 1 0 1992 0 1 1512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5372_6
timestamp 1731220455
transform 1 0 1784 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5371_6
timestamp 1731220455
transform 1 0 1568 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5370_6
timestamp 1731220455
transform 1 0 1336 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5369_6
timestamp 1731220455
transform 1 0 1784 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5368_6
timestamp 1731220455
transform 1 0 1648 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5367_6
timestamp 1731220455
transform 1 0 1488 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5366_6
timestamp 1731220455
transform 1 0 1336 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5365_6
timestamp 1731220455
transform 1 0 1184 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5364_6
timestamp 1731220455
transform 1 0 1144 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5363_6
timestamp 1731220455
transform 1 0 1312 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5362_6
timestamp 1731220455
transform 1 0 1480 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5361_6
timestamp 1731220455
transform 1 0 1784 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5360_6
timestamp 1731220455
transform 1 0 1640 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5359_6
timestamp 1731220455
transform 1 0 1600 0 1 1096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5358_6
timestamp 1731220455
transform 1 0 1392 0 1 1096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5357_6
timestamp 1731220455
transform 1 0 1784 0 1 1096
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5356_6
timestamp 1731220455
transform 1 0 1992 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5355_6
timestamp 1731220455
transform 1 0 2224 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5354_6
timestamp 1731220455
transform 1 0 2464 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5353_6
timestamp 1731220455
transform 1 0 2424 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5352_6
timestamp 1731220455
transform 1 0 2288 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5351_6
timestamp 1731220455
transform 1 0 2152 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5350_6
timestamp 1731220455
transform 1 0 2568 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5349_6
timestamp 1731220455
transform 1 0 2712 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5348_6
timestamp 1731220455
transform 1 0 2672 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5347_6
timestamp 1731220455
transform 1 0 2536 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5346_6
timestamp 1731220455
transform 1 0 2400 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5345_6
timestamp 1731220455
transform 1 0 2264 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5344_6
timestamp 1731220455
transform 1 0 2128 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5343_6
timestamp 1731220455
transform 1 0 1992 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5342_6
timestamp 1731220455
transform 1 0 2136 0 -1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5341_6
timestamp 1731220455
transform 1 0 1992 0 -1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5340_6
timestamp 1731220455
transform 1 0 1992 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5339_6
timestamp 1731220455
transform 1 0 1784 0 1 580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5338_6
timestamp 1731220455
transform 1 0 1560 0 1 580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5337_6
timestamp 1731220455
transform 1 0 1416 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5336_6
timestamp 1731220455
transform 1 0 1680 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5335_6
timestamp 1731220455
transform 1 0 1544 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5334_6
timestamp 1731220455
transform 1 0 1320 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5333_6
timestamp 1731220455
transform 1 0 1096 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5332_6
timestamp 1731220455
transform 1 0 984 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5331_6
timestamp 1731220455
transform 1 0 1200 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5330_6
timestamp 1731220455
transform 1 0 1424 0 -1 344
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5329_6
timestamp 1731220455
transform 1 0 1368 0 1 84
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5328_6
timestamp 1731220455
transform 1 0 1224 0 1 84
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5327_6
timestamp 1731220455
transform 1 0 1512 0 1 84
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5326_6
timestamp 1731220455
transform 1 0 1648 0 1 84
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5325_6
timestamp 1731220455
transform 1 0 1784 0 1 84
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5324_6
timestamp 1731220455
transform 1 0 1992 0 1 104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5323_6
timestamp 1731220455
transform 1 0 2360 0 1 104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5322_6
timestamp 1731220455
transform 1 0 2168 0 1 104
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5321_6
timestamp 1731220455
transform 1 0 2144 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5320_6
timestamp 1731220455
transform 1 0 1992 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5319_6
timestamp 1731220455
transform 1 0 2336 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5318_6
timestamp 1731220455
transform 1 0 2560 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5317_6
timestamp 1731220455
transform 1 0 2456 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5316_6
timestamp 1731220455
transform 1 0 2312 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5315_6
timestamp 1731220455
transform 1 0 2168 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5314_6
timestamp 1731220455
transform 1 0 2304 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5313_6
timestamp 1731220455
transform 1 0 2496 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5312_6
timestamp 1731220455
transform 1 0 2680 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5311_6
timestamp 1731220455
transform 1 0 2976 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5310_6
timestamp 1731220455
transform 1 0 2632 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5309_6
timestamp 1731220455
transform 1 0 2296 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5308_6
timestamp 1731220455
transform 1 0 2304 0 -1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5307_6
timestamp 1731220455
transform 1 0 2464 0 -1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5306_6
timestamp 1731220455
transform 1 0 2624 0 -1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5305_6
timestamp 1731220455
transform 1 0 2960 0 -1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5304_6
timestamp 1731220455
transform 1 0 2792 0 -1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5303_6
timestamp 1731220455
transform 1 0 2808 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5302_6
timestamp 1731220455
transform 1 0 2944 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5301_6
timestamp 1731220455
transform 1 0 3080 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5300_6
timestamp 1731220455
transform 1 0 3488 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5299_6
timestamp 1731220455
transform 1 0 3352 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5298_6
timestamp 1731220455
transform 1 0 3216 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5297_6
timestamp 1731220455
transform 1 0 3144 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5296_6
timestamp 1731220455
transform 1 0 3000 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5295_6
timestamp 1731220455
transform 1 0 2856 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5294_6
timestamp 1731220455
transform 1 0 3432 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5293_6
timestamp 1731220455
transform 1 0 3288 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5292_6
timestamp 1731220455
transform 1 0 3104 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5291_6
timestamp 1731220455
transform 1 0 2904 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5290_6
timestamp 1731220455
transform 1 0 2688 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5289_6
timestamp 1731220455
transform 1 0 3648 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5288_6
timestamp 1731220455
transform 1 0 3480 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5287_6
timestamp 1731220455
transform 1 0 3296 0 1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5286_6
timestamp 1731220455
transform 1 0 3240 0 -1 1308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5285_6
timestamp 1731220455
transform 1 0 3376 0 -1 1308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5284_6
timestamp 1731220455
transform 1 0 3512 0 -1 1308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5283_6
timestamp 1731220455
transform 1 0 3648 0 -1 1308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5282_6
timestamp 1731220455
transform 1 0 3856 0 -1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5281_6
timestamp 1731220455
transform 1 0 3856 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5280_6
timestamp 1731220455
transform 1 0 4000 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5279_6
timestamp 1731220455
transform 1 0 4176 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5278_6
timestamp 1731220455
transform 1 0 4528 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5277_6
timestamp 1731220455
transform 1 0 4352 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5276_6
timestamp 1731220455
transform 1 0 4336 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5275_6
timestamp 1731220455
transform 1 0 4168 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5274_6
timestamp 1731220455
transform 1 0 4000 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5273_6
timestamp 1731220455
transform 1 0 3856 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5272_6
timestamp 1731220455
transform 1 0 3648 0 1 1512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5271_6
timestamp 1731220455
transform 1 0 3448 0 1 1512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5270_6
timestamp 1731220455
transform 1 0 3232 0 1 1512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5269_6
timestamp 1731220455
transform 1 0 3016 0 1 1512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5268_6
timestamp 1731220455
transform 1 0 3488 0 -1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5267_6
timestamp 1731220455
transform 1 0 3304 0 -1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5266_6
timestamp 1731220455
transform 1 0 3120 0 -1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5265_6
timestamp 1731220455
transform 1 0 2944 0 -1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5264_6
timestamp 1731220455
transform 1 0 2760 0 -1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5263_6
timestamp 1731220455
transform 1 0 3080 0 1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5262_6
timestamp 1731220455
transform 1 0 2928 0 1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5261_6
timestamp 1731220455
transform 1 0 2784 0 1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5260_6
timestamp 1731220455
transform 1 0 2640 0 1 1736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5259_6
timestamp 1731220455
transform 1 0 2736 0 -1 1960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5258_6
timestamp 1731220455
transform 1 0 2872 0 -1 1960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5257_6
timestamp 1731220455
transform 1 0 3288 0 -1 1960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5256_6
timestamp 1731220455
transform 1 0 3144 0 -1 1960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5255_6
timestamp 1731220455
transform 1 0 3008 0 -1 1960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5254_6
timestamp 1731220455
transform 1 0 2976 0 1 1972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5253_6
timestamp 1731220455
transform 1 0 3152 0 1 1972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5252_6
timestamp 1731220455
transform 1 0 3320 0 1 1972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5251_6
timestamp 1731220455
transform 1 0 3496 0 1 1972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5250_6
timestamp 1731220455
transform 1 0 3648 0 1 1972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5249_6
timestamp 1731220455
transform 1 0 3856 0 1 2072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5248_6
timestamp 1731220455
transform 1 0 4040 0 1 2072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5247_6
timestamp 1731220455
transform 1 0 4248 0 1 2072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5246_6
timestamp 1731220455
transform 1 0 4456 0 1 2072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5245_6
timestamp 1731220455
transform 1 0 4240 0 -1 2296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5244_6
timestamp 1731220455
transform 1 0 4040 0 -1 2296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5243_6
timestamp 1731220455
transform 1 0 3856 0 -1 2296
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5242_6
timestamp 1731220455
transform 1 0 3648 0 1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5241_6
timestamp 1731220455
transform 1 0 3488 0 1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5240_6
timestamp 1731220455
transform 1 0 3304 0 1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5239_6
timestamp 1731220455
transform 1 0 3120 0 1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5238_6
timestamp 1731220455
transform 1 0 2928 0 1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5237_6
timestamp 1731220455
transform 1 0 3640 0 -1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5236_6
timestamp 1731220455
transform 1 0 3424 0 -1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5235_6
timestamp 1731220455
transform 1 0 3208 0 -1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5234_6
timestamp 1731220455
transform 1 0 2992 0 -1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5233_6
timestamp 1731220455
transform 1 0 2768 0 -1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5232_6
timestamp 1731220455
transform 1 0 3400 0 1 2496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5231_6
timestamp 1731220455
transform 1 0 3208 0 1 2496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5230_6
timestamp 1731220455
transform 1 0 3016 0 1 2496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5229_6
timestamp 1731220455
transform 1 0 2824 0 1 2496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5228_6
timestamp 1731220455
transform 1 0 2624 0 1 2496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5227_6
timestamp 1731220455
transform 1 0 3352 0 -1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5226_6
timestamp 1731220455
transform 1 0 3216 0 -1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5225_6
timestamp 1731220455
transform 1 0 3080 0 -1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5224_6
timestamp 1731220455
transform 1 0 2944 0 -1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5223_6
timestamp 1731220455
transform 1 0 2808 0 -1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5222_6
timestamp 1731220455
transform 1 0 2728 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5221_6
timestamp 1731220455
transform 1 0 2488 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5220_6
timestamp 1731220455
transform 1 0 2968 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5219_6
timestamp 1731220455
transform 1 0 2952 0 -1 2944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5218_6
timestamp 1731220455
transform 1 0 2816 0 -1 2944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5217_6
timestamp 1731220455
transform 1 0 2808 0 1 2952
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5216_6
timestamp 1731220455
transform 1 0 2752 0 -1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5215_6
timestamp 1731220455
transform 1 0 2584 0 -1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5214_6
timestamp 1731220455
transform 1 0 2736 0 1 3200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5213_6
timestamp 1731220455
transform 1 0 2680 0 -1 3424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5212_6
timestamp 1731220455
transform 1 0 2816 0 -1 3424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5211_6
timestamp 1731220455
transform 1 0 2712 0 1 3460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5210_6
timestamp 1731220455
transform 1 0 2576 0 1 3460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5209_6
timestamp 1731220455
transform 1 0 2440 0 1 3460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5208_6
timestamp 1731220455
transform 1 0 2304 0 1 3460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5207_6
timestamp 1731220455
transform 1 0 2752 0 -1 3696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5206_6
timestamp 1731220455
transform 1 0 2560 0 -1 3696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5205_6
timestamp 1731220455
transform 1 0 2376 0 -1 3696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5204_6
timestamp 1731220455
transform 1 0 2192 0 -1 3696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5203_6
timestamp 1731220455
transform 1 0 2016 0 -1 3696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5202_6
timestamp 1731220455
transform 1 0 2600 0 1 3704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5201_6
timestamp 1731220455
transform 1 0 2440 0 1 3704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5200_6
timestamp 1731220455
transform 1 0 2280 0 1 3704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5199_6
timestamp 1731220455
transform 1 0 2128 0 1 3704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5198_6
timestamp 1731220455
transform 1 0 1992 0 1 3704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5197_6
timestamp 1731220455
transform 1 0 1784 0 -1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5196_6
timestamp 1731220455
transform 1 0 1784 0 1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5195_6
timestamp 1731220455
transform 1 0 1648 0 1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5194_6
timestamp 1731220455
transform 1 0 1488 0 1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5193_6
timestamp 1731220455
transform 1 0 1328 0 1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5192_6
timestamp 1731220455
transform 1 0 1472 0 -1 4056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5191_6
timestamp 1731220455
transform 1 0 1640 0 -1 4056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5190_6
timestamp 1731220455
transform 1 0 1784 0 -1 4056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5189_6
timestamp 1731220455
transform 1 0 1992 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5188_6
timestamp 1731220455
transform 1 0 1992 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5187_6
timestamp 1731220455
transform 1 0 2256 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5186_6
timestamp 1731220455
transform 1 0 2456 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5185_6
timestamp 1731220455
transform 1 0 2240 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5184_6
timestamp 1731220455
transform 1 0 2016 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5183_6
timestamp 1731220455
transform 1 0 2088 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5182_6
timestamp 1731220455
transform 1 0 2312 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5181_6
timestamp 1731220455
transform 1 0 2536 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5180_6
timestamp 1731220455
transform 1 0 2688 0 1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5179_6
timestamp 1731220455
transform 1 0 2456 0 1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5178_6
timestamp 1731220455
transform 1 0 2224 0 1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5177_6
timestamp 1731220455
transform 1 0 1992 0 1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5176_6
timestamp 1731220455
transform 1 0 2800 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5175_6
timestamp 1731220455
transform 1 0 2624 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5174_6
timestamp 1731220455
transform 1 0 2448 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5173_6
timestamp 1731220455
transform 1 0 2280 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5172_6
timestamp 1731220455
transform 1 0 2128 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5171_6
timestamp 1731220455
transform 1 0 1992 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5170_6
timestamp 1731220455
transform 1 0 1784 0 1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5169_6
timestamp 1731220455
transform 1 0 1512 0 1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5168_6
timestamp 1731220455
transform 1 0 1376 0 -1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5167_6
timestamp 1731220455
transform 1 0 1784 0 -1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5166_6
timestamp 1731220455
transform 1 0 1592 0 -1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5165_6
timestamp 1731220455
transform 1 0 1496 0 1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5164_6
timestamp 1731220455
transform 1 0 1704 0 1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5163_6
timestamp 1731220455
transform 1 0 1672 0 -1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5162_6
timestamp 1731220455
transform 1 0 1488 0 -1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5161_6
timestamp 1731220455
transform 1 0 1312 0 -1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5160_6
timestamp 1731220455
transform 1 0 1528 0 1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5159_6
timestamp 1731220455
transform 1 0 1312 0 1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5158_6
timestamp 1731220455
transform 1 0 1304 0 -1 4056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5157_6
timestamp 1731220455
transform 1 0 1136 0 -1 4056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5156_6
timestamp 1731220455
transform 1 0 960 0 -1 4056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5155_6
timestamp 1731220455
transform 1 0 824 0 1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5154_6
timestamp 1731220455
transform 1 0 1000 0 1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5153_6
timestamp 1731220455
transform 1 0 1168 0 1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5152_6
timestamp 1731220455
transform 1 0 1232 0 -1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5151_6
timestamp 1731220455
transform 1 0 1520 0 -1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5150_6
timestamp 1731220455
transform 1 0 1512 0 1 3584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5149_6
timestamp 1731220455
transform 1 0 1376 0 1 3584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5148_6
timestamp 1731220455
transform 1 0 1240 0 1 3584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5147_6
timestamp 1731220455
transform 1 0 1104 0 1 3584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5146_6
timestamp 1731220455
transform 1 0 968 0 1 3584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5145_6
timestamp 1731220455
transform 1 0 832 0 1 3584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5144_6
timestamp 1731220455
transform 1 0 696 0 1 3584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5143_6
timestamp 1731220455
transform 1 0 560 0 1 3584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5142_6
timestamp 1731220455
transform 1 0 424 0 1 3584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5141_6
timestamp 1731220455
transform 1 0 288 0 1 3584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5140_6
timestamp 1731220455
transform 1 0 152 0 1 3584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5139_6
timestamp 1731220455
transform 1 0 960 0 -1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5138_6
timestamp 1731220455
transform 1 0 704 0 -1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5137_6
timestamp 1731220455
transform 1 0 480 0 -1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5136_6
timestamp 1731220455
transform 1 0 280 0 -1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5135_6
timestamp 1731220455
transform 1 0 640 0 1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5134_6
timestamp 1731220455
transform 1 0 448 0 1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5133_6
timestamp 1731220455
transform 1 0 248 0 1 3832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5132_6
timestamp 1731220455
transform 1 0 200 0 -1 4056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5131_6
timestamp 1731220455
transform 1 0 392 0 -1 4056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5130_6
timestamp 1731220455
transform 1 0 776 0 -1 4056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5129_6
timestamp 1731220455
transform 1 0 584 0 -1 4056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5128_6
timestamp 1731220455
transform 1 0 512 0 1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5127_6
timestamp 1731220455
transform 1 0 344 0 1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5126_6
timestamp 1731220455
transform 1 0 696 0 1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5125_6
timestamp 1731220455
transform 1 0 1096 0 1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5124_6
timestamp 1731220455
transform 1 0 888 0 1 4072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5123_6
timestamp 1731220455
transform 1 0 792 0 -1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5122_6
timestamp 1731220455
transform 1 0 624 0 -1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5121_6
timestamp 1731220455
transform 1 0 960 0 -1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5120_6
timestamp 1731220455
transform 1 0 1136 0 -1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5119_6
timestamp 1731220455
transform 1 0 1296 0 1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5118_6
timestamp 1731220455
transform 1 0 1104 0 1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5117_6
timestamp 1731220455
transform 1 0 912 0 1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5116_6
timestamp 1731220455
transform 1 0 736 0 1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5115_6
timestamp 1731220455
transform 1 0 568 0 1 4308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5114_6
timestamp 1731220455
transform 1 0 1168 0 -1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5113_6
timestamp 1731220455
transform 1 0 968 0 -1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5112_6
timestamp 1731220455
transform 1 0 776 0 -1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5111_6
timestamp 1731220455
transform 1 0 592 0 -1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5110_6
timestamp 1731220455
transform 1 0 416 0 -1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5109_6
timestamp 1731220455
transform 1 0 1216 0 1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5108_6
timestamp 1731220455
transform 1 0 928 0 1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5107_6
timestamp 1731220455
transform 1 0 664 0 1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5106_6
timestamp 1731220455
transform 1 0 424 0 1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5105_6
timestamp 1731220455
transform 1 0 208 0 1 4536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5104_6
timestamp 1731220455
transform 1 0 672 0 -1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5103_6
timestamp 1731220455
transform 1 0 536 0 -1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5102_6
timestamp 1731220455
transform 1 0 400 0 -1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5101_6
timestamp 1731220455
transform 1 0 264 0 -1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5100_6
timestamp 1731220455
transform 1 0 128 0 -1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_599_6
timestamp 1731220455
transform 1 0 128 0 1 4772
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_598_6
timestamp 1731220455
transform 1 0 264 0 1 4772
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_597_6
timestamp 1731220455
transform 1 0 672 0 1 4772
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_596_6
timestamp 1731220455
transform 1 0 536 0 1 4772
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_595_6
timestamp 1731220455
transform 1 0 400 0 1 4772
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_594_6
timestamp 1731220455
transform 1 0 264 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_593_6
timestamp 1731220455
transform 1 0 128 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_592_6
timestamp 1731220455
transform 1 0 672 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_591_6
timestamp 1731220455
transform 1 0 536 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_590_6
timestamp 1731220455
transform 1 0 400 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_589_6
timestamp 1731220455
transform 1 0 264 0 1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_588_6
timestamp 1731220455
transform 1 0 400 0 1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_587_6
timestamp 1731220455
transform 1 0 536 0 1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_586_6
timestamp 1731220455
transform 1 0 944 0 1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_585_6
timestamp 1731220455
transform 1 0 808 0 1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_584_6
timestamp 1731220455
transform 1 0 672 0 1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_583_6
timestamp 1731220455
transform 1 0 560 0 -1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_582_6
timestamp 1731220455
transform 1 0 424 0 -1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_581_6
timestamp 1731220455
transform 1 0 696 0 -1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_580_6
timestamp 1731220455
transform 1 0 832 0 -1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_579_6
timestamp 1731220455
transform 1 0 968 0 -1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_578_6
timestamp 1731220455
transform 1 0 1376 0 -1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_577_6
timestamp 1731220455
transform 1 0 1240 0 -1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_576_6
timestamp 1731220455
transform 1 0 1104 0 -1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_575_6
timestamp 1731220455
transform 1 0 696 0 1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_574_6
timestamp 1731220455
transform 1 0 560 0 1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_573_6
timestamp 1731220455
transform 1 0 424 0 1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_572_6
timestamp 1731220455
transform 1 0 832 0 1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_571_6
timestamp 1731220455
transform 1 0 968 0 1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_570_6
timestamp 1731220455
transform 1 0 1104 0 1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_569_6
timestamp 1731220455
transform 1 0 1240 0 1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_568_6
timestamp 1731220455
transform 1 0 1376 0 1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_567_6
timestamp 1731220455
transform 1 0 1376 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_566_6
timestamp 1731220455
transform 1 0 1512 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_565_6
timestamp 1731220455
transform 1 0 1648 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_564_6
timestamp 1731220455
transform 1 0 1784 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_563_6
timestamp 1731220455
transform 1 0 1992 0 1 5448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_562_6
timestamp 1731220455
transform 1 0 2128 0 1 5448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_561_6
timestamp 1731220455
transform 1 0 2264 0 1 5448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_560_6
timestamp 1731220455
transform 1 0 2704 0 1 5448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_559_6
timestamp 1731220455
transform 1 0 2552 0 1 5448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_558_6
timestamp 1731220455
transform 1 0 2400 0 1 5448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_557_6
timestamp 1731220455
transform 1 0 2344 0 -1 5672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_556_6
timestamp 1731220455
transform 1 0 2208 0 -1 5672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_555_6
timestamp 1731220455
transform 1 0 2072 0 -1 5672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_554_6
timestamp 1731220455
transform 1 0 2480 0 -1 5672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_553_6
timestamp 1731220455
transform 1 0 2616 0 -1 5672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_552_6
timestamp 1731220455
transform 1 0 2752 0 -1 5672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_551_6
timestamp 1731220455
transform 1 0 2888 0 -1 5672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_550_6
timestamp 1731220455
transform 1 0 3024 0 -1 5672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_549_6
timestamp 1731220455
transform 1 0 3160 0 -1 5672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_548_6
timestamp 1731220455
transform 1 0 3296 0 -1 5672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_547_6
timestamp 1731220455
transform 1 0 3432 0 -1 5672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_546_6
timestamp 1731220455
transform 1 0 3568 0 -1 5672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_545_6
timestamp 1731220455
transform 1 0 3480 0 1 5448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_544_6
timestamp 1731220455
transform 1 0 3320 0 1 5448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_543_6
timestamp 1731220455
transform 1 0 3160 0 1 5448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_542_6
timestamp 1731220455
transform 1 0 3008 0 1 5448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_541_6
timestamp 1731220455
transform 1 0 2856 0 1 5448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_540_6
timestamp 1731220455
transform 1 0 3208 0 -1 5436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_539_6
timestamp 1731220455
transform 1 0 3072 0 -1 5436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_538_6
timestamp 1731220455
transform 1 0 2936 0 -1 5436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_537_6
timestamp 1731220455
transform 1 0 2800 0 -1 5436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_536_6
timestamp 1731220455
transform 1 0 2968 0 1 5176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_535_6
timestamp 1731220455
transform 1 0 2712 0 1 5176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_534_6
timestamp 1731220455
transform 1 0 2464 0 1 5176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_533_6
timestamp 1731220455
transform 1 0 2216 0 1 5176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_532_6
timestamp 1731220455
transform 1 0 3360 0 -1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_531_6
timestamp 1731220455
transform 1 0 3216 0 -1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_530_6
timestamp 1731220455
transform 1 0 3080 0 -1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_529_6
timestamp 1731220455
transform 1 0 2944 0 -1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_528_6
timestamp 1731220455
transform 1 0 2808 0 -1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_527_6
timestamp 1731220455
transform 1 0 2672 0 -1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_526_6
timestamp 1731220455
transform 1 0 2536 0 -1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_525_6
timestamp 1731220455
transform 1 0 2400 0 -1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_524_6
timestamp 1731220455
transform 1 0 2264 0 -1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_523_6
timestamp 1731220455
transform 1 0 2128 0 -1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_522_6
timestamp 1731220455
transform 1 0 1992 0 -1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_521_6
timestamp 1731220455
transform 1 0 1992 0 1 5176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_520_6
timestamp 1731220455
transform 1 0 1784 0 -1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_519_6
timestamp 1731220455
transform 1 0 1648 0 -1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_518_6
timestamp 1731220455
transform 1 0 1512 0 -1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_517_6
timestamp 1731220455
transform 1 0 1784 0 1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_516_6
timestamp 1731220455
transform 1 0 1648 0 1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_515_6
timestamp 1731220455
transform 1 0 1512 0 1 5256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_514_6
timestamp 1731220455
transform 1 0 1240 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_513_6
timestamp 1731220455
transform 1 0 1104 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_512_6
timestamp 1731220455
transform 1 0 968 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_511_6
timestamp 1731220455
transform 1 0 832 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_510_6
timestamp 1731220455
transform 1 0 1160 0 1 5492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_59_6
timestamp 1731220455
transform 1 0 1024 0 1 5492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_58_6
timestamp 1731220455
transform 1 0 888 0 1 5492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_57_6
timestamp 1731220455
transform 1 0 752 0 1 5492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_56_6
timestamp 1731220455
transform 1 0 944 0 -1 5732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_55_6
timestamp 1731220455
transform 1 0 808 0 -1 5732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_54_6
timestamp 1731220455
transform 1 0 672 0 -1 5732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_53_6
timestamp 1731220455
transform 1 0 536 0 -1 5732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_52_6
timestamp 1731220455
transform 1 0 400 0 -1 5732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_51_6
timestamp 1731220455
transform 1 0 264 0 -1 5732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_50_6
timestamp 1731220455
transform 1 0 128 0 -1 5732
box 3 5 132 108
<< end >>
