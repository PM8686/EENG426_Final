magic
tech sky130l
timestamp 1730254555
<< m1 >>
rect 8 32 12 36
rect 32 32 36 36
rect 56 32 60 36
rect 80 32 84 36
rect 104 32 108 36
rect 8 4 12 8
<< labels >>
rlabel m1 s 8 32 12 36 6 in_50_6
port 1 nsew signal input
rlabel m1 s 32 32 36 36 6 in_51_6
port 2 nsew signal input
rlabel m1 s 56 32 60 36 6 in_52_6
port 3 nsew signal input
rlabel m1 s 8 4 12 8 6 out
port 4 nsew signal output
rlabel m1 s 80 32 84 36 6 Vdd
port 5 nsew power input
rlabel m1 s 104 32 108 36 6 GND
port 6 nsew ground input
<< properties >>
string LEFsite CoreSite
string LEFclass CORE
string FIXED_BBOX 0 0 120 40
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
