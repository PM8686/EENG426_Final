magic
tech sky130l
timestamp 1729040465
<< ndiffusion >>
rect 8 11 13 16
rect 8 8 9 11
rect 12 8 13 11
rect 8 6 13 8
rect 15 6 20 16
rect 22 14 27 16
rect 22 11 23 14
rect 26 11 27 14
rect 22 6 27 11
rect 33 15 38 16
rect 33 12 34 15
rect 37 12 38 15
rect 33 10 38 12
rect 40 14 47 16
rect 40 11 41 14
rect 44 11 47 14
rect 40 10 47 11
rect 43 6 47 10
rect 49 11 54 16
rect 49 8 50 11
rect 53 8 54 11
rect 49 6 54 8
rect 60 14 65 16
rect 60 11 61 14
rect 64 11 65 14
rect 60 6 65 11
rect 67 11 72 16
rect 67 8 68 11
rect 71 8 72 11
rect 67 6 72 8
<< ndc >>
rect 9 8 12 11
rect 23 11 26 14
rect 34 12 37 15
rect 41 11 44 14
rect 50 8 53 11
rect 61 11 64 14
rect 68 8 71 11
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
rect 38 10 40 16
rect 47 6 49 16
rect 65 6 67 16
<< pdiffusion >>
rect 8 35 13 38
rect 8 32 9 35
rect 12 32 13 35
rect 8 23 13 32
rect 15 31 19 38
rect 15 30 20 31
rect 15 27 16 30
rect 19 27 20 30
rect 15 23 20 27
rect 22 27 27 31
rect 22 24 23 27
rect 26 24 27 27
rect 22 23 27 24
rect 33 28 38 38
rect 33 25 34 28
rect 37 25 38 28
rect 33 23 38 25
rect 40 23 47 38
rect 49 37 54 38
rect 49 34 50 37
rect 53 34 54 37
rect 49 23 54 34
rect 60 35 65 38
rect 60 32 61 35
rect 64 32 65 35
rect 60 23 65 32
rect 67 28 72 38
rect 67 25 68 28
rect 71 25 72 28
rect 67 23 72 25
<< pdc >>
rect 9 32 12 35
rect 16 27 19 30
rect 23 24 26 27
rect 34 25 37 28
rect 50 34 53 37
rect 61 32 64 35
rect 68 25 71 28
<< ptransistor >>
rect 13 23 15 38
rect 20 23 22 31
rect 38 23 40 38
rect 47 23 49 38
rect 65 23 67 38
<< polysilicon >>
rect 9 45 15 46
rect 9 42 10 45
rect 13 42 15 45
rect 9 41 15 42
rect 32 45 40 46
rect 32 42 33 45
rect 36 42 40 45
rect 32 41 40 42
rect 43 45 49 46
rect 43 42 44 45
rect 47 42 49 45
rect 43 41 49 42
rect 13 38 15 41
rect 20 38 28 39
rect 38 38 40 41
rect 47 38 49 41
rect 65 38 67 40
rect 20 35 24 38
rect 27 35 28 38
rect 20 34 28 35
rect 20 31 22 34
rect 13 16 15 23
rect 20 16 22 23
rect 38 16 40 23
rect 47 16 49 23
rect 65 22 67 23
rect 65 21 80 22
rect 65 20 76 21
rect 65 16 67 20
rect 75 18 76 20
rect 79 18 80 21
rect 75 17 80 18
rect 38 8 40 10
rect 13 4 15 6
rect 20 4 22 6
rect 47 4 49 6
rect 65 4 67 6
<< pc >>
rect 10 42 13 45
rect 33 42 36 45
rect 44 42 47 45
rect 24 35 27 38
rect 76 18 79 21
<< m1 >>
rect 8 45 13 46
rect 8 42 10 45
rect 8 40 13 42
rect 16 42 20 44
rect 19 40 20 42
rect 24 42 33 45
rect 36 42 37 45
rect 24 41 37 42
rect 8 32 9 35
rect 12 32 13 35
rect 16 30 19 39
rect 24 38 28 41
rect 40 40 44 45
rect 47 42 48 45
rect 51 42 54 43
rect 27 35 28 38
rect 51 37 54 39
rect 24 34 28 35
rect 49 34 50 37
rect 53 34 54 37
rect 60 32 61 35
rect 64 32 65 35
rect 56 28 60 29
rect 16 26 19 27
rect 23 27 26 28
rect 33 25 34 28
rect 37 25 38 28
rect 59 25 60 28
rect 67 25 68 28
rect 71 25 72 28
rect 23 21 26 24
rect 23 17 26 18
rect 34 21 37 22
rect 34 15 37 18
rect 56 15 60 25
rect 75 18 76 21
rect 79 18 80 21
rect 8 11 12 12
rect 22 11 23 14
rect 26 11 27 14
rect 34 11 37 12
rect 41 14 44 15
rect 56 14 64 15
rect 8 8 9 11
rect 8 7 12 8
rect 8 4 9 7
rect 8 3 12 4
rect 41 7 44 11
rect 41 3 44 4
rect 50 11 53 12
rect 50 7 53 8
rect 56 11 61 14
rect 56 10 64 11
rect 68 11 71 12
rect 56 4 60 10
rect 68 7 71 8
rect 50 3 53 4
rect 68 3 71 4
<< m2c >>
rect 16 39 19 42
rect 9 32 12 35
rect 51 39 54 42
rect 61 32 64 35
rect 34 25 37 28
rect 56 25 59 28
rect 68 25 71 28
rect 23 18 26 21
rect 34 18 37 21
rect 76 18 79 21
rect 23 11 26 14
rect 9 4 12 7
rect 41 4 44 7
rect 50 4 53 7
rect 61 11 64 14
rect 68 4 71 7
<< m2 >>
rect 15 42 55 43
rect 15 39 16 42
rect 19 39 51 42
rect 54 39 55 42
rect 15 38 55 39
rect 8 35 65 36
rect 8 32 9 35
rect 12 32 61 35
rect 64 32 65 35
rect 8 31 65 32
rect 33 28 72 29
rect 33 25 34 28
rect 37 25 56 28
rect 59 25 68 28
rect 71 25 72 28
rect 33 24 72 25
rect 22 21 80 22
rect 22 18 23 21
rect 26 18 34 21
rect 37 18 76 21
rect 79 18 80 21
rect 22 17 80 18
rect 22 14 65 15
rect 22 11 23 14
rect 26 11 61 14
rect 64 11 65 14
rect 22 10 65 11
rect 8 7 46 8
rect 8 4 9 7
rect 12 4 41 7
rect 44 4 46 7
rect 8 3 46 4
rect 49 7 72 8
rect 49 4 50 7
rect 53 4 68 7
rect 71 4 72 7
rect 49 3 72 4
<< labels >>
rlabel pdiffusion 23 24 23 24 3 _S
rlabel polysilicon 21 17 21 17 3 S
rlabel polysilicon 21 22 21 22 3 S
rlabel pdiffusion 16 24 16 24 3 Vdd
rlabel polysilicon 14 17 14 17 3 A
rlabel polysilicon 14 22 14 22 3 A
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 24 9 24 3 #5
rlabel ndiffusion 50 7 50 7 3 #10
rlabel polysilicon 48 17 48 17 3 B
rlabel polysilicon 48 22 48 22 3 B
rlabel pdiffusion 50 24 50 24 3 Vdd
rlabel ndiffusion 41 11 41 11 3 GND
rlabel polysilicon 39 17 39 17 3 S
rlabel polysilicon 39 22 39 22 3 S
rlabel ndiffusion 34 11 34 11 3 _S
rlabel ndiffusion 68 7 68 7 3 #10
rlabel polysilicon 66 17 66 17 3 _S
rlabel polysilicon 66 22 66 22 3 _S
rlabel pdiffusion 61 24 61 24 3 #5
rlabel m1 9 41 9 41 3 A
port 6 e
rlabel m2 9 5 9 5 3 GND
rlabel ndiffusion 61 7 61 7 3 Y
rlabel pdiffusion 34 24 34 24 3 Y
rlabel pdiffusion 68 24 68 24 3 Y
rlabel ndiffusion 23 7 23 7 3 Y
rlabel m1 57 5 57 5 3 Y
rlabel m2c 17 41 17 41 3 Vdd
rlabel m1 41 41 41 41 3 B
rlabel m1 25 41 25 41 3 S
<< end >>
