magic
tech TSMC180
timestamp 1734145863
<< ndiffusion >>
rect 6 10 12 12
rect 6 8 7 10
rect 9 8 12 10
rect 6 7 12 8
rect 14 11 20 12
rect 14 9 17 11
rect 19 9 20 11
rect 14 7 20 9
<< ndcontact >>
rect 7 8 9 10
rect 17 9 19 11
<< ntransistor >>
rect 12 7 14 12
<< pdiffusion >>
rect 6 35 12 36
rect 6 33 7 35
rect 9 33 12 35
rect 6 28 12 33
rect 14 31 20 36
rect 14 29 17 31
rect 19 29 20 31
rect 14 28 20 29
<< pdcontact >>
rect 7 33 9 35
rect 17 29 19 31
<< ptransistor >>
rect 12 28 14 36
<< polysilicon >>
rect 17 43 21 44
rect 17 42 18 43
rect 12 41 18 42
rect 20 41 21 43
rect 12 40 21 41
rect 12 36 14 40
rect 12 12 14 28
rect 12 4 14 7
<< polycontact >>
rect 18 41 20 43
<< m1 >>
rect 18 44 21 50
rect 17 43 21 44
rect 17 41 18 43
rect 20 41 21 43
rect 17 40 21 41
rect 6 35 11 37
rect 6 33 7 35
rect 9 33 11 35
rect 6 32 11 33
rect 16 31 20 32
rect 16 29 17 31
rect 19 29 20 31
rect 16 28 20 29
rect 17 19 20 28
rect 17 16 27 19
rect 17 12 20 16
rect 16 11 20 12
rect 5 10 10 11
rect 5 8 7 10
rect 9 8 10 10
rect 16 9 17 11
rect 19 9 20 11
rect 16 8 20 9
rect 5 6 10 8
<< labels >>
rlabel ndiffusion 15 8 15 8 3 Y
rlabel pdiffusion 15 29 15 29 3 Y
rlabel polysilicon 13 13 13 13 3 A
rlabel polysilicon 13 26 13 26 3 A
rlabel pdiffusion 7 29 7 29 3 Vdd
rlabel m1 25 17 25 17 3 Y
rlabel m1 19 48 19 48 3 A
rlabel pdcontact 8 34 9 35 3 Vdd
rlabel ndcontact 7 8 8 9 2 GND
<< end >>
