magic
tech sky130l
timestamp 1730589753
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 10 20 12
rect 15 7 16 10
rect 19 7 20 10
rect 15 6 20 7
<< ndc >>
rect 9 7 12 10
rect 16 7 19 10
<< ntransistor >>
rect 13 6 15 12
<< pdiffusion >>
rect 8 28 13 29
rect 8 25 9 28
rect 12 25 13 28
rect 8 19 13 25
rect 15 28 20 29
rect 15 25 16 28
rect 19 25 20 28
rect 15 19 20 25
<< pdc >>
rect 9 25 12 28
rect 16 25 19 28
<< ptransistor >>
rect 13 19 15 29
<< polysilicon >>
rect 13 36 20 37
rect 13 33 16 36
rect 19 33 20 36
rect 13 32 20 33
rect 13 29 15 32
rect 13 12 15 19
rect 13 4 15 6
<< pc >>
rect 16 33 19 36
<< m1 >>
rect 7 37 12 38
rect 7 34 8 37
rect 11 34 12 37
rect 7 33 12 34
rect 8 28 12 33
rect 8 25 9 28
rect 8 24 12 25
rect 16 36 20 37
rect 19 33 20 36
rect 16 28 20 33
rect 19 25 20 28
rect 16 24 20 25
rect 8 10 12 11
rect 16 10 20 11
rect 8 8 9 10
rect 7 7 9 8
rect 12 7 13 10
rect 19 7 20 10
rect 7 4 8 7
rect 11 4 12 7
rect 16 4 20 7
rect 7 3 12 4
<< m2c >>
rect 8 34 11 37
rect 8 4 11 7
<< m2 >>
rect 7 37 12 38
rect 7 34 8 37
rect 11 34 12 37
rect 7 33 12 34
rect 7 7 12 8
rect 7 4 8 7
rect 11 4 12 7
rect 7 3 12 4
<< labels >>
rlabel m1 s 19 7 20 10 6 Y
port 1 nsew signal output
rlabel m1 s 16 7 19 10 6 Y
port 1 nsew signal output
rlabel m1 s 16 10 20 11 6 Y
port 1 nsew signal output
rlabel m1 s 16 4 20 7 6 Y
port 1 nsew signal output
rlabel m1 s 9 25 12 28 6 Vdd
port 2 nsew power input
rlabel m1 s 8 24 12 25 6 Vdd
port 2 nsew power input
rlabel m1 s 8 25 9 28 6 Vdd
port 2 nsew power input
rlabel m1 s 8 28 12 36 6 Vdd
port 2 nsew power input
rlabel m1 s 9 7 12 10 6 GND
port 3 nsew ground input
rlabel m1 s 8 4 12 7 6 GND
port 3 nsew ground input
rlabel m1 s 8 7 9 10 6 GND
port 3 nsew ground input
rlabel m1 s 8 10 12 11 6 GND
port 3 nsew ground input
rlabel space 0 0 24 40 3 prboundary
rlabel ndiffusion 16 7 16 7 3 Y
rlabel ndiffusion 16 8 16 8 3 Y
rlabel ndiffusion 16 11 16 11 3 Y
rlabel ndiffusion 13 8 13 8 3 GND
rlabel pdiffusion 16 20 16 20 3 x
rlabel pdiffusion 16 26 16 26 3 x
rlabel pdiffusion 16 29 16 29 3 x
rlabel pdiffusion 13 26 13 26 3 Vdd
rlabel polysilicon 14 5 14 5 3 x
rlabel ntransistor 14 7 14 7 3 x
rlabel polysilicon 14 13 14 13 3 x
rlabel ptransistor 14 20 14 20 3 x
rlabel polysilicon 14 30 14 30 3 x
rlabel polysilicon 14 33 14 33 3 x
rlabel polysilicon 14 34 14 34 3 x
rlabel polysilicon 14 37 14 37 3 x
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel m1 20 8 20 8 3 Y
port 1 e default output
rlabel m1 20 26 20 26 3 x
rlabel m1 20 34 20 34 3 x
rlabel ndc 17 8 17 8 3 Y
port 1 e default output
rlabel m1 17 11 17 11 3 Y
port 1 e default output
rlabel m1 17 25 17 25 3 x
rlabel pdc 17 26 17 26 3 x
rlabel m1 17 29 17 29 3 x
rlabel pc 17 34 17 34 3 x
rlabel m1 17 37 17 37 3 x
rlabel m1 17 5 17 5 3 Y
port 1 e
rlabel ndc 10 8 10 8 3 GND
rlabel pdc 10 26 10 26 3 Vdd
rlabel m2c 9 5 9 5 3 GND
rlabel m1 9 8 9 8 3 GND
rlabel m1 9 11 9 11 3 GND
rlabel m1 9 25 9 25 3 Vdd
rlabel m1 9 26 9 26 3 Vdd
rlabel m1 9 29 9 29 3 Vdd
<< properties >>
string LEFsite CoreSite
string LEFclass CORE
string FIXED_BBOX 0 0 24 40
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
