magic
tech TSMC180
timestamp 1734150802
<< ppdiff >>
rect 6 3 11 8
<< nndiff >>
rect 6 13 11 18
<< m1 >>
rect 6 17 9 20
rect 6 10 9 13
<< labels >>
rlabel space 0 0 18 30 6 prboundary
rlabel m1 7 11 7 11 3 GND
port 1 e
rlabel m1 7 18 7 18 3 Vdd
port 2 e
rlabel ppdiff 7 4 7 4 3 GND
rlabel nndiff 7 13 7 13 3 Vdd
<< end >>
