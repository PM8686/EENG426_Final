magic
tech sky130l
timestamp 1731220505
<< m1 >>
rect 2624 5627 2628 5687
rect 584 5551 588 5611
rect 1464 5551 1468 5611
rect 3072 5475 3076 5583
rect 2136 5403 2140 5471
rect 2656 5395 2660 5455
rect 880 5211 884 5259
rect 832 5067 836 5127
rect 1384 5067 1388 5127
rect 2664 5055 2668 5111
rect 4280 5071 4284 5127
rect 5080 5071 5084 5127
rect 5504 4923 5508 4983
rect 4064 4807 4068 4863
rect 3504 4655 3508 4715
rect 5200 4675 5204 4735
rect 264 4571 268 4631
rect 5648 4619 5652 4735
rect 3304 4531 3308 4587
rect 824 4339 828 4399
rect 2896 4391 2900 4451
rect 4608 4415 4612 4475
rect 4792 4415 4796 4475
rect 5208 4415 5212 4475
rect 1240 4227 1244 4275
rect 4264 4167 4268 4227
rect 4616 4167 4620 4227
rect 4888 4167 4892 4227
rect 640 4091 644 4151
rect 5648 4095 5652 4227
rect 528 3999 532 4047
rect 2248 4035 2252 4091
rect 3104 4035 3108 4083
rect 1432 3863 1436 3923
rect 1696 3863 1700 3923
rect 2248 3895 2252 3955
rect 2424 3895 2428 3955
rect 2768 3895 2772 3955
rect 5272 3883 5276 3943
rect 4256 3783 4260 3839
rect 5480 3783 5484 3831
rect 888 3627 892 3687
rect 4368 3623 4372 3683
rect 1104 3367 1108 3427
rect 2680 3287 2684 3343
rect 4320 3143 4324 3203
rect 1776 3035 1780 3091
rect 264 2899 268 2959
rect 4272 2891 4276 2951
rect 768 2799 772 2859
rect 4360 2783 4364 2839
rect 1176 2667 1180 2727
rect 4152 2639 4156 2771
rect 856 2443 860 2503
rect 280 2339 284 2439
rect 4440 2379 4444 2487
rect 296 2199 300 2259
rect 2408 2207 2412 2267
rect 496 1959 500 2019
rect 5120 1923 5124 1983
rect 1232 1463 1236 1523
rect 4448 1459 4452 1519
rect 2992 1359 2996 1415
rect 3152 1359 3156 1415
rect 2136 1223 2140 1283
rect 2984 1223 2988 1347
rect 3592 1223 3596 1283
rect 5648 1235 5652 1519
rect 3240 1123 3244 1179
rect 5176 883 5180 939
rect 4496 751 4500 811
rect 3648 643 3652 703
rect 336 383 340 479
rect 608 383 612 455
rect 944 391 948 447
rect 800 191 804 319
rect 992 259 996 319
<< m2c >>
rect 2608 5687 2612 5691
rect 2624 5687 2628 5691
rect 2760 5687 2764 5691
rect 2912 5687 2916 5691
rect 3072 5687 3076 5691
rect 3240 5687 3244 5691
rect 3416 5687 3420 5691
rect 3592 5687 3596 5691
rect 256 5671 260 5675
rect 496 5671 500 5675
rect 760 5671 764 5675
rect 1032 5671 1036 5675
rect 1304 5671 1308 5675
rect 1576 5671 1580 5675
rect 1848 5671 1852 5675
rect 2624 5623 2628 5627
rect 552 5611 556 5615
rect 584 5611 588 5615
rect 744 5611 748 5615
rect 952 5611 956 5615
rect 1184 5611 1188 5615
rect 1424 5611 1428 5615
rect 1464 5611 1468 5615
rect 1680 5611 1684 5615
rect 1912 5611 1916 5615
rect 584 5547 588 5551
rect 4232 5587 4236 5591
rect 4368 5587 4372 5591
rect 4504 5587 4508 5591
rect 4640 5587 4644 5591
rect 4776 5587 4780 5591
rect 4912 5587 4916 5591
rect 5048 5587 5052 5591
rect 5184 5587 5188 5591
rect 5320 5587 5324 5591
rect 1464 5547 1468 5551
rect 3072 5583 3076 5587
rect 2120 5515 2124 5519
rect 2328 5515 2332 5519
rect 2560 5515 2564 5519
rect 2784 5515 2788 5519
rect 2992 5515 2996 5519
rect 3200 5515 3204 5519
rect 3400 5515 3404 5519
rect 3600 5515 3604 5519
rect 3776 5515 3780 5519
rect 4400 5495 4404 5499
rect 4608 5495 4612 5499
rect 4816 5495 4820 5499
rect 5024 5495 5028 5499
rect 5232 5495 5236 5499
rect 2136 5471 2140 5475
rect 3072 5471 3076 5475
rect 2120 5455 2124 5459
rect 912 5447 916 5451
rect 1048 5447 1052 5451
rect 1184 5447 1188 5451
rect 1320 5447 1324 5451
rect 1456 5448 1460 5452
rect 2264 5455 2268 5459
rect 2440 5455 2444 5459
rect 2624 5455 2628 5459
rect 2656 5455 2660 5459
rect 2816 5457 2820 5461
rect 3008 5455 3012 5459
rect 3208 5455 3212 5459
rect 3408 5457 3412 5461
rect 2136 5399 2140 5403
rect 2656 5391 2660 5395
rect 1000 5367 1004 5371
rect 1136 5367 1140 5371
rect 1280 5367 1284 5371
rect 1432 5367 1436 5371
rect 1592 5367 1596 5371
rect 1760 5367 1764 5371
rect 1912 5367 1916 5371
rect 3984 5307 3988 5311
rect 4120 5307 4124 5311
rect 4256 5307 4260 5311
rect 4400 5307 4404 5311
rect 4560 5307 4564 5311
rect 4728 5307 4732 5311
rect 4904 5307 4908 5311
rect 5088 5309 5092 5313
rect 2176 5267 2180 5271
rect 2584 5267 2588 5271
rect 2984 5267 2988 5271
rect 3392 5267 3396 5271
rect 3776 5267 3780 5271
rect 880 5259 884 5263
rect 4096 5243 4100 5247
rect 4296 5243 4300 5247
rect 4496 5243 4500 5247
rect 4704 5243 4708 5247
rect 4920 5243 4924 5247
rect 5136 5243 5140 5247
rect 880 5207 884 5211
rect 2336 5207 2340 5211
rect 2688 5207 2692 5211
rect 3040 5207 3044 5211
rect 3400 5207 3404 5211
rect 3760 5207 3764 5211
rect 712 5199 716 5203
rect 864 5199 868 5203
rect 1024 5199 1028 5203
rect 1192 5199 1196 5203
rect 1368 5199 1372 5203
rect 1552 5199 1556 5203
rect 1744 5199 1748 5203
rect 1912 5199 1916 5203
rect 464 5127 468 5131
rect 632 5127 636 5131
rect 808 5127 812 5131
rect 832 5127 836 5131
rect 992 5127 996 5131
rect 1176 5127 1180 5131
rect 1360 5127 1364 5131
rect 1384 5127 1388 5131
rect 1544 5127 1548 5131
rect 1728 5127 1732 5131
rect 1912 5127 1916 5131
rect 4280 5127 4284 5131
rect 832 5063 836 5067
rect 1384 5063 1388 5067
rect 2664 5111 2668 5115
rect 4280 5067 4284 5071
rect 5080 5127 5084 5131
rect 5080 5067 5084 5071
rect 4224 5059 4228 5063
rect 4472 5061 4476 5065
rect 4720 5059 4724 5063
rect 4968 5059 4972 5063
rect 5224 5059 5228 5063
rect 2664 5051 2668 5055
rect 2392 5043 2396 5047
rect 2640 5043 2644 5047
rect 2880 5045 2884 5049
rect 3120 5043 3124 5047
rect 3360 5045 3364 5049
rect 3600 5043 3604 5047
rect 4080 4983 4084 4987
rect 4320 4983 4324 4987
rect 4544 4983 4548 4987
rect 4752 4983 4756 4987
rect 4952 4983 4956 4987
rect 5136 4983 5140 4987
rect 5312 4983 5316 4987
rect 5488 4983 5492 4987
rect 5504 4983 5508 4987
rect 5640 4983 5644 4987
rect 256 4959 260 4963
rect 448 4959 452 4963
rect 680 4959 684 4963
rect 936 4959 940 4963
rect 1208 4959 1212 4963
rect 1496 4959 1500 4963
rect 1784 4959 1788 4963
rect 2280 4951 2284 4955
rect 2416 4951 2420 4955
rect 2552 4951 2556 4955
rect 2696 4951 2700 4955
rect 2840 4951 2844 4955
rect 2992 4951 2996 4955
rect 3144 4951 3148 4955
rect 3296 4951 3300 4955
rect 3448 4951 3452 4955
rect 5504 4919 5508 4923
rect 256 4875 260 4879
rect 392 4875 396 4879
rect 528 4875 532 4879
rect 664 4875 668 4879
rect 800 4875 804 4879
rect 4064 4863 4068 4867
rect 4064 4803 4068 4807
rect 3984 4795 3988 4799
rect 4200 4795 4204 4799
rect 4424 4795 4428 4799
rect 4632 4795 4636 4799
rect 4824 4795 4828 4799
rect 5000 4795 5004 4799
rect 5168 4795 5172 4799
rect 5336 4795 5340 4799
rect 5496 4795 5500 4799
rect 5640 4795 5644 4799
rect 2552 4779 2556 4783
rect 2696 4779 2700 4783
rect 2848 4779 2852 4783
rect 3000 4779 3004 4783
rect 3152 4779 3156 4783
rect 3304 4779 3308 4783
rect 5040 4735 5044 4739
rect 5184 4735 5188 4739
rect 5200 4735 5204 4739
rect 5336 4735 5340 4739
rect 5496 4735 5500 4739
rect 5640 4735 5644 4739
rect 5648 4735 5652 4739
rect 2120 4715 2124 4719
rect 2256 4715 2260 4719
rect 2392 4715 2396 4719
rect 2528 4715 2532 4719
rect 2664 4715 2668 4719
rect 2800 4715 2804 4719
rect 2936 4715 2940 4719
rect 3072 4715 3076 4719
rect 3208 4715 3212 4719
rect 3344 4715 3348 4719
rect 3496 4715 3500 4719
rect 3504 4715 3508 4719
rect 3640 4715 3644 4719
rect 3776 4715 3780 4719
rect 256 4699 260 4703
rect 392 4699 396 4703
rect 528 4699 532 4703
rect 664 4699 668 4703
rect 800 4699 804 4703
rect 5200 4671 5204 4675
rect 3504 4651 3508 4655
rect 256 4631 260 4635
rect 264 4631 268 4635
rect 392 4631 396 4635
rect 528 4631 532 4635
rect 664 4631 668 4635
rect 800 4631 804 4635
rect 5648 4615 5652 4619
rect 264 4567 268 4571
rect 3304 4587 3308 4591
rect 4896 4547 4900 4551
rect 5080 4547 5084 4551
rect 5272 4547 5276 4551
rect 5464 4547 5468 4551
rect 5640 4547 5644 4551
rect 3304 4527 3308 4531
rect 2448 4519 2452 4523
rect 2704 4519 2708 4523
rect 2952 4519 2956 4523
rect 3200 4521 3204 4525
rect 3440 4521 3444 4525
rect 3688 4521 3692 4525
rect 4584 4475 4588 4479
rect 4608 4475 4612 4479
rect 4768 4475 4772 4479
rect 4792 4475 4796 4479
rect 4976 4475 4980 4479
rect 5192 4475 5196 4479
rect 5208 4475 5212 4479
rect 5424 4475 5428 4479
rect 5640 4475 5644 4479
rect 464 4459 468 4463
rect 640 4459 644 4463
rect 816 4459 820 4463
rect 1000 4459 1004 4463
rect 1184 4459 1188 4463
rect 1368 4459 1372 4463
rect 1552 4459 1556 4463
rect 1744 4459 1748 4463
rect 1912 4459 1916 4463
rect 2640 4451 2644 4455
rect 2880 4451 2884 4455
rect 2896 4451 2900 4455
rect 3112 4451 3116 4455
rect 3344 4451 3348 4455
rect 3568 4451 3572 4455
rect 3776 4451 3780 4455
rect 664 4399 668 4403
rect 808 4399 812 4403
rect 824 4399 828 4403
rect 960 4399 964 4403
rect 1120 4399 1124 4403
rect 1280 4399 1284 4403
rect 1440 4399 1444 4403
rect 1600 4399 1604 4403
rect 1768 4399 1772 4403
rect 1912 4399 1916 4403
rect 4608 4411 4612 4415
rect 4792 4411 4796 4415
rect 5208 4411 5212 4415
rect 2896 4387 2900 4391
rect 824 4335 828 4339
rect 3984 4287 3988 4291
rect 4120 4287 4124 4291
rect 4256 4287 4260 4291
rect 4408 4287 4412 4291
rect 4608 4287 4612 4291
rect 4840 4287 4844 4291
rect 5104 4287 5108 4291
rect 5376 4287 5380 4291
rect 5640 4287 5644 4291
rect 1240 4275 1244 4279
rect 2120 4275 2124 4279
rect 2504 4275 2508 4279
rect 2928 4275 2932 4279
rect 3360 4275 3364 4279
rect 3776 4275 3780 4279
rect 3984 4227 3988 4231
rect 4120 4227 4124 4231
rect 4256 4227 4260 4231
rect 4264 4227 4268 4231
rect 4400 4227 4404 4231
rect 4600 4227 4604 4231
rect 4616 4227 4620 4231
rect 4832 4227 4836 4231
rect 4888 4227 4892 4231
rect 5096 4227 5100 4231
rect 5368 4227 5372 4231
rect 5640 4227 5644 4231
rect 5648 4227 5652 4231
rect 1240 4223 1244 4227
rect 752 4215 756 4219
rect 896 4215 900 4219
rect 1048 4215 1052 4219
rect 1208 4215 1212 4219
rect 1376 4217 1380 4221
rect 1544 4215 1548 4219
rect 1720 4215 1724 4219
rect 2120 4187 2124 4191
rect 2288 4187 2292 4191
rect 2480 4187 2484 4191
rect 2680 4187 2684 4191
rect 2880 4187 2884 4191
rect 3080 4187 3084 4191
rect 4264 4163 4268 4167
rect 4616 4163 4620 4167
rect 4888 4163 4892 4167
rect 616 4151 620 4155
rect 640 4151 644 4155
rect 800 4151 804 4155
rect 992 4151 996 4155
rect 1200 4151 1204 4155
rect 1424 4151 1428 4155
rect 1648 4151 1652 4155
rect 1880 4151 1884 4155
rect 640 4087 644 4091
rect 2248 4091 2252 4095
rect 5648 4091 5652 4095
rect 528 4047 532 4051
rect 2248 4031 2252 4035
rect 3104 4083 3108 4087
rect 3104 4031 3108 4035
rect 2200 4023 2204 4027
rect 2384 4025 2388 4029
rect 2568 4023 2572 4027
rect 2744 4023 2748 4027
rect 2912 4025 2916 4029
rect 3080 4023 3084 4027
rect 3256 4025 3260 4029
rect 4688 4023 4692 4027
rect 4824 4023 4828 4027
rect 4960 4023 4964 4027
rect 5096 4023 5100 4027
rect 5232 4023 5236 4027
rect 5368 4023 5372 4027
rect 5504 4023 5508 4027
rect 5640 4023 5644 4027
rect 528 3995 532 3999
rect 256 3987 260 3991
rect 464 3987 468 3991
rect 720 3989 724 3993
rect 1000 3987 1004 3991
rect 1304 3987 1308 3991
rect 1616 3987 1620 3991
rect 1912 3987 1916 3991
rect 2224 3955 2228 3959
rect 2248 3955 2252 3959
rect 2408 3955 2412 3959
rect 2424 3955 2428 3959
rect 2584 3955 2588 3959
rect 2760 3955 2764 3959
rect 2768 3955 2772 3959
rect 2928 3955 2932 3959
rect 3096 3955 3100 3959
rect 3272 3955 3276 3959
rect 3448 3955 3452 3959
rect 256 3923 260 3927
rect 440 3923 444 3927
rect 664 3923 668 3927
rect 904 3923 908 3927
rect 1152 3925 1156 3929
rect 1408 3923 1412 3927
rect 1432 3923 1436 3927
rect 1672 3923 1676 3927
rect 1696 3923 1700 3927
rect 1912 3923 1916 3927
rect 1432 3859 1436 3863
rect 2248 3891 2252 3895
rect 2424 3891 2428 3895
rect 4456 3943 4460 3947
rect 4640 3943 4644 3947
rect 4832 3943 4836 3947
rect 5024 3943 5028 3947
rect 5224 3943 5228 3947
rect 5272 3943 5276 3947
rect 5424 3943 5428 3947
rect 5624 3943 5628 3947
rect 2768 3891 2772 3895
rect 5272 3879 5276 3883
rect 1696 3859 1700 3863
rect 4256 3839 4260 3843
rect 2416 3783 2420 3787
rect 2648 3783 2652 3787
rect 2864 3783 2868 3787
rect 3072 3783 3076 3787
rect 3280 3783 3284 3787
rect 3480 3783 3484 3787
rect 3688 3785 3692 3789
rect 4256 3779 4260 3783
rect 5480 3831 5484 3835
rect 5480 3779 5484 3783
rect 4176 3771 4180 3775
rect 4392 3771 4396 3775
rect 4608 3771 4612 3775
rect 4824 3771 4828 3775
rect 5032 3771 5036 3775
rect 5240 3771 5244 3775
rect 5448 3771 5452 3775
rect 5640 3771 5644 3775
rect 392 3751 396 3755
rect 600 3751 604 3755
rect 832 3751 836 3755
rect 1088 3751 1092 3755
rect 1360 3751 1364 3755
rect 1640 3753 1644 3757
rect 1912 3751 1916 3755
rect 2504 3719 2508 3723
rect 2744 3719 2748 3723
rect 2968 3719 2972 3723
rect 3184 3719 3188 3723
rect 3392 3719 3396 3723
rect 3592 3719 3596 3723
rect 3776 3719 3780 3723
rect 728 3687 732 3691
rect 872 3687 876 3691
rect 888 3687 892 3691
rect 1024 3687 1028 3691
rect 1184 3687 1188 3691
rect 1352 3687 1356 3691
rect 1520 3687 1524 3691
rect 1688 3687 1692 3691
rect 1856 3687 1860 3691
rect 3984 3683 3988 3687
rect 4152 3683 4156 3687
rect 4344 3683 4348 3687
rect 4368 3683 4372 3687
rect 4536 3683 4540 3687
rect 4728 3683 4732 3687
rect 888 3623 892 3627
rect 4368 3619 4372 3623
rect 1464 3587 1468 3591
rect 2536 3547 2540 3551
rect 2672 3547 2676 3551
rect 2808 3547 2812 3551
rect 3984 3519 3988 3523
rect 4120 3519 4124 3523
rect 4256 3519 4260 3523
rect 4392 3519 4396 3523
rect 4528 3519 4532 3523
rect 4664 3519 4668 3523
rect 4800 3519 4804 3523
rect 4936 3519 4940 3523
rect 5072 3519 5076 3523
rect 5208 3519 5212 3523
rect 904 3511 908 3515
rect 1040 3511 1044 3515
rect 1176 3511 1180 3515
rect 1312 3511 1316 3515
rect 1448 3511 1452 3515
rect 1584 3511 1588 3515
rect 1720 3511 1724 3515
rect 1856 3511 1860 3515
rect 4928 3451 4932 3455
rect 5064 3451 5068 3455
rect 5200 3451 5204 3455
rect 5336 3451 5340 3455
rect 5472 3451 5476 3455
rect 2696 3447 2700 3451
rect 2920 3447 2924 3451
rect 3144 3447 3148 3451
rect 3360 3447 3364 3451
rect 3576 3447 3580 3451
rect 3776 3447 3780 3451
rect 824 3427 828 3431
rect 960 3427 964 3431
rect 1096 3427 1100 3431
rect 1104 3427 1108 3431
rect 1232 3427 1236 3431
rect 1368 3427 1372 3431
rect 1504 3427 1508 3431
rect 1640 3427 1644 3431
rect 1776 3427 1780 3431
rect 1912 3427 1916 3431
rect 1104 3363 1108 3367
rect 2680 3343 2684 3347
rect 3984 3289 3988 3293
rect 4264 3287 4268 3291
rect 4552 3287 4556 3291
rect 4816 3287 4820 3291
rect 5064 3287 5068 3291
rect 5304 3287 5308 3291
rect 5552 3289 5556 3293
rect 2680 3283 2684 3287
rect 2656 3275 2660 3279
rect 2840 3277 2844 3281
rect 3024 3275 3028 3279
rect 3208 3275 3212 3279
rect 3392 3275 3396 3279
rect 880 3259 884 3263
rect 1016 3259 1020 3263
rect 1160 3259 1164 3263
rect 1312 3261 1316 3265
rect 1464 3259 1468 3263
rect 1616 3259 1620 3263
rect 1776 3259 1780 3263
rect 1912 3259 1916 3263
rect 2120 3215 2124 3219
rect 2352 3215 2356 3219
rect 2600 3215 2604 3219
rect 2840 3215 2844 3219
rect 3072 3215 3076 3219
rect 3304 3215 3308 3219
rect 3544 3215 3548 3219
rect 4008 3203 4012 3207
rect 4280 3203 4284 3207
rect 4320 3203 4324 3207
rect 4536 3203 4540 3207
rect 4784 3203 4788 3207
rect 5032 3203 5036 3207
rect 5288 3203 5292 3207
rect 488 3199 492 3203
rect 744 3199 748 3203
rect 1024 3199 1028 3203
rect 1320 3199 1324 3203
rect 1624 3199 1628 3203
rect 1912 3199 1916 3203
rect 4320 3139 4324 3143
rect 1776 3091 1780 3095
rect 2608 3051 2612 3055
rect 2904 3051 2908 3055
rect 3200 3051 3204 3055
rect 3496 3051 3500 3055
rect 3776 3051 3780 3055
rect 4056 3035 4060 3039
rect 4256 3035 4260 3039
rect 4456 3035 4460 3039
rect 4648 3035 4652 3039
rect 4840 3035 4844 3039
rect 5040 3035 5044 3039
rect 1776 3031 1780 3035
rect 256 3023 260 3027
rect 432 3023 436 3027
rect 632 3023 636 3027
rect 832 3023 836 3027
rect 1024 3023 1028 3027
rect 1216 3023 1220 3027
rect 1400 3023 1404 3027
rect 1576 3023 1580 3027
rect 1752 3023 1756 3027
rect 1912 3023 1916 3027
rect 2288 2983 2292 2987
rect 2448 2983 2452 2987
rect 2616 2983 2620 2987
rect 2800 2983 2804 2987
rect 3000 2983 3004 2987
rect 3216 2983 3220 2987
rect 3432 2983 3436 2987
rect 3656 2983 3660 2987
rect 256 2959 260 2963
rect 264 2959 268 2963
rect 392 2959 396 2963
rect 528 2959 532 2963
rect 664 2959 668 2963
rect 800 2959 804 2963
rect 4096 2951 4100 2955
rect 4256 2951 4260 2955
rect 4272 2951 4276 2955
rect 4432 2951 4436 2955
rect 4616 2951 4620 2955
rect 4816 2951 4820 2955
rect 5024 2951 5028 2955
rect 5232 2951 5236 2955
rect 5448 2951 5452 2955
rect 5640 2951 5644 2955
rect 264 2895 268 2899
rect 4272 2887 4276 2891
rect 768 2859 772 2863
rect 4360 2839 4364 2843
rect 2120 2815 2124 2819
rect 2256 2815 2260 2819
rect 2392 2815 2396 2819
rect 2528 2815 2532 2819
rect 2664 2815 2668 2819
rect 2808 2815 2812 2819
rect 2960 2815 2964 2819
rect 3120 2815 3124 2819
rect 3280 2815 3284 2819
rect 3440 2815 3444 2819
rect 768 2795 772 2799
rect 352 2791 356 2795
rect 488 2791 492 2795
rect 624 2791 628 2795
rect 760 2791 764 2795
rect 896 2791 900 2795
rect 4360 2779 4364 2783
rect 3984 2771 3988 2775
rect 4136 2771 4140 2775
rect 4152 2771 4156 2775
rect 4336 2773 4340 2777
rect 4560 2771 4564 2775
rect 4816 2771 4820 2775
rect 5088 2771 5092 2775
rect 5376 2771 5380 2775
rect 5640 2771 5644 2775
rect 2120 2751 2124 2755
rect 2256 2751 2260 2755
rect 2400 2751 2404 2755
rect 2560 2751 2564 2755
rect 2720 2751 2724 2755
rect 2880 2751 2884 2755
rect 3040 2751 3044 2755
rect 3200 2751 3204 2755
rect 472 2727 476 2731
rect 672 2727 676 2731
rect 896 2727 900 2731
rect 1136 2727 1140 2731
rect 1176 2727 1180 2731
rect 1392 2727 1396 2731
rect 1664 2727 1668 2731
rect 1912 2727 1916 2731
rect 4064 2699 4068 2703
rect 1176 2663 1180 2667
rect 4320 2699 4324 2703
rect 4624 2699 4628 2703
rect 4960 2699 4964 2703
rect 5312 2701 5316 2705
rect 5640 2699 5644 2703
rect 4152 2635 4156 2639
rect 2824 2579 2828 2583
rect 2960 2579 2964 2583
rect 3096 2579 3100 2583
rect 512 2563 516 2567
rect 664 2563 668 2567
rect 824 2563 828 2567
rect 992 2565 996 2569
rect 1160 2563 1164 2567
rect 1328 2563 1332 2567
rect 1496 2563 1500 2567
rect 1664 2563 1668 2567
rect 1840 2563 1844 2567
rect 4016 2535 4020 2539
rect 4192 2535 4196 2539
rect 4392 2535 4396 2539
rect 4616 2535 4620 2539
rect 4856 2535 4860 2539
rect 5120 2535 5124 2539
rect 5392 2535 5396 2539
rect 5640 2535 5644 2539
rect 2704 2519 2708 2523
rect 2856 2519 2860 2523
rect 3008 2519 3012 2523
rect 3160 2519 3164 2523
rect 3320 2519 3324 2523
rect 424 2503 428 2507
rect 632 2503 636 2507
rect 832 2503 836 2507
rect 856 2503 860 2507
rect 1016 2503 1020 2507
rect 1192 2503 1196 2507
rect 1368 2503 1372 2507
rect 1536 2503 1540 2507
rect 1704 2503 1708 2507
rect 1872 2503 1876 2507
rect 4440 2487 4444 2491
rect 3984 2471 3988 2475
rect 4184 2471 4188 2475
rect 4416 2471 4420 2475
rect 280 2439 284 2443
rect 856 2439 860 2443
rect 4664 2471 4668 2475
rect 4920 2471 4924 2475
rect 5184 2471 5188 2475
rect 5448 2471 5452 2475
rect 4440 2375 4444 2379
rect 2120 2339 2124 2343
rect 2400 2339 2404 2343
rect 2696 2339 2700 2343
rect 2984 2339 2988 2343
rect 3272 2339 3276 2343
rect 3560 2339 3564 2343
rect 256 2335 260 2339
rect 280 2335 284 2339
rect 528 2335 532 2339
rect 816 2335 820 2339
rect 1096 2335 1100 2339
rect 1376 2335 1380 2339
rect 1656 2335 1660 2339
rect 1912 2335 1916 2339
rect 3984 2307 3988 2311
rect 4216 2307 4220 2311
rect 4464 2307 4468 2311
rect 4704 2307 4708 2311
rect 4936 2307 4940 2311
rect 5168 2307 5172 2311
rect 5408 2307 5412 2311
rect 5640 2307 5644 2311
rect 2120 2267 2124 2271
rect 2256 2267 2260 2271
rect 2392 2267 2396 2271
rect 2408 2267 2412 2271
rect 2544 2267 2548 2271
rect 2704 2267 2708 2271
rect 2864 2267 2868 2271
rect 3024 2267 3028 2271
rect 3176 2267 3180 2271
rect 3328 2267 3332 2271
rect 3480 2267 3484 2271
rect 3640 2267 3644 2271
rect 3776 2267 3780 2271
rect 256 2259 260 2263
rect 296 2259 300 2263
rect 520 2259 524 2263
rect 808 2259 812 2263
rect 1096 2259 1100 2263
rect 1392 2259 1396 2263
rect 4688 2223 4692 2227
rect 4824 2223 4828 2227
rect 4960 2223 4964 2227
rect 5096 2223 5100 2227
rect 5232 2223 5236 2227
rect 5368 2223 5372 2227
rect 5504 2223 5508 2227
rect 5640 2223 5644 2227
rect 2408 2203 2412 2207
rect 296 2195 300 2199
rect 2256 2095 2260 2099
rect 2456 2095 2460 2099
rect 2656 2095 2660 2099
rect 2856 2095 2860 2099
rect 3048 2095 3052 2099
rect 3240 2095 3244 2099
rect 3424 2095 3428 2099
rect 3608 2095 3612 2099
rect 3776 2095 3780 2099
rect 256 2083 260 2087
rect 528 2083 532 2087
rect 856 2083 860 2087
rect 1208 2083 1212 2087
rect 1568 2083 1572 2087
rect 1912 2083 1916 2087
rect 5080 2043 5084 2047
rect 5216 2043 5220 2047
rect 5352 2043 5356 2047
rect 2120 2027 2124 2031
rect 2376 2027 2380 2031
rect 2648 2027 2652 2031
rect 2896 2027 2900 2031
rect 3128 2027 3132 2031
rect 3352 2027 3356 2031
rect 3576 2027 3580 2031
rect 3776 2027 3780 2031
rect 320 2019 324 2023
rect 480 2019 484 2023
rect 496 2019 500 2023
rect 656 2019 660 2023
rect 848 2019 852 2023
rect 1056 2019 1060 2023
rect 1264 2019 1268 2023
rect 1480 2019 1484 2023
rect 1704 2019 1708 2023
rect 1912 2019 1916 2023
rect 4824 1983 4828 1987
rect 4960 1983 4964 1987
rect 5104 1983 5108 1987
rect 5120 1983 5124 1987
rect 5256 1983 5260 1987
rect 5416 1983 5420 1987
rect 5584 1983 5588 1987
rect 496 1955 500 1959
rect 5120 1919 5124 1923
rect 320 1847 324 1851
rect 512 1847 516 1851
rect 720 1847 724 1851
rect 944 1847 948 1851
rect 1176 1847 1180 1851
rect 1408 1847 1412 1851
rect 1648 1847 1652 1851
rect 1896 1849 1900 1853
rect 2120 1851 2124 1855
rect 2440 1851 2444 1855
rect 2744 1851 2748 1855
rect 3024 1851 3028 1855
rect 3288 1851 3292 1855
rect 3544 1851 3548 1855
rect 3776 1851 3780 1855
rect 4400 1819 4404 1823
rect 4624 1819 4628 1823
rect 4856 1819 4860 1823
rect 5104 1821 5108 1825
rect 5360 1819 5364 1823
rect 5624 1819 5628 1823
rect 2208 1787 2212 1791
rect 2488 1787 2492 1791
rect 2760 1787 2764 1791
rect 3024 1787 3028 1791
rect 3280 1787 3284 1791
rect 3536 1787 3540 1791
rect 3776 1787 3780 1791
rect 256 1771 260 1775
rect 400 1771 404 1775
rect 576 1771 580 1775
rect 752 1771 756 1775
rect 928 1771 932 1775
rect 1104 1771 1108 1775
rect 1280 1771 1284 1775
rect 1456 1771 1460 1775
rect 1632 1771 1636 1775
rect 1808 1771 1812 1775
rect 3984 1751 3988 1755
rect 4184 1751 4188 1755
rect 4440 1751 4444 1755
rect 4720 1751 4724 1755
rect 5024 1751 5028 1755
rect 5344 1751 5348 1755
rect 5640 1751 5644 1755
rect 1000 1603 1004 1607
rect 1136 1603 1140 1607
rect 1272 1603 1276 1607
rect 1408 1603 1412 1607
rect 1544 1603 1548 1607
rect 1680 1603 1684 1607
rect 2208 1591 2212 1595
rect 2344 1591 2348 1595
rect 2480 1591 2484 1595
rect 2616 1591 2620 1595
rect 2752 1591 2756 1595
rect 2896 1591 2900 1595
rect 3040 1591 3044 1595
rect 3984 1583 3988 1587
rect 4120 1583 4124 1587
rect 4264 1583 4268 1587
rect 4448 1583 4452 1587
rect 4656 1583 4660 1587
rect 4888 1583 4892 1587
rect 5136 1583 5140 1587
rect 5400 1583 5404 1587
rect 5640 1583 5644 1587
rect 2240 1527 2244 1531
rect 2376 1527 2380 1531
rect 2512 1527 2516 1531
rect 2648 1527 2652 1531
rect 2784 1527 2788 1531
rect 2920 1527 2924 1531
rect 3056 1527 3060 1531
rect 3192 1527 3196 1531
rect 3328 1527 3332 1531
rect 256 1523 260 1527
rect 488 1523 492 1527
rect 728 1523 732 1527
rect 968 1523 972 1527
rect 1208 1523 1212 1527
rect 1232 1523 1236 1527
rect 1448 1523 1452 1527
rect 3984 1519 3988 1523
rect 4208 1519 4212 1523
rect 4440 1519 4444 1523
rect 4448 1519 4452 1523
rect 4672 1519 4676 1523
rect 4912 1519 4916 1523
rect 5160 1519 5164 1523
rect 5408 1519 5412 1523
rect 5640 1520 5644 1524
rect 5648 1519 5652 1523
rect 1232 1459 1236 1463
rect 4448 1455 4452 1459
rect 2992 1415 2996 1419
rect 2992 1355 2996 1359
rect 3152 1415 3156 1419
rect 3152 1355 3156 1359
rect 3984 1355 3988 1359
rect 4208 1355 4212 1359
rect 4448 1355 4452 1359
rect 4672 1355 4676 1359
rect 4896 1355 4900 1359
rect 5112 1355 5116 1359
rect 5328 1355 5332 1359
rect 5544 1355 5548 1359
rect 256 1347 260 1351
rect 456 1347 460 1351
rect 680 1347 684 1351
rect 904 1347 908 1351
rect 1128 1347 1132 1351
rect 2224 1347 2228 1351
rect 2368 1347 2372 1351
rect 2512 1347 2516 1351
rect 2664 1347 2668 1351
rect 2816 1347 2820 1351
rect 2976 1347 2980 1351
rect 2984 1347 2988 1351
rect 3136 1347 3140 1351
rect 3296 1347 3300 1351
rect 256 1287 260 1291
rect 464 1287 468 1291
rect 704 1287 708 1291
rect 944 1287 948 1291
rect 1184 1287 1188 1291
rect 2120 1283 2124 1287
rect 2136 1283 2140 1287
rect 2272 1283 2276 1287
rect 2464 1283 2468 1287
rect 2672 1283 2676 1287
rect 2888 1283 2892 1287
rect 2136 1219 2140 1223
rect 3984 1295 3988 1299
rect 4216 1295 4220 1299
rect 4488 1295 4492 1299
rect 4768 1295 4772 1299
rect 5064 1295 5068 1299
rect 5360 1295 5364 1299
rect 5640 1295 5644 1299
rect 3112 1283 3116 1287
rect 3336 1283 3340 1287
rect 3568 1283 3572 1287
rect 3592 1283 3596 1287
rect 3776 1283 3780 1287
rect 2984 1219 2988 1223
rect 5648 1231 5652 1235
rect 3592 1219 3596 1223
rect 3240 1179 3244 1183
rect 3240 1119 3244 1123
rect 256 1111 260 1115
rect 400 1111 404 1115
rect 568 1111 572 1115
rect 728 1111 732 1115
rect 888 1111 892 1115
rect 1048 1113 1052 1117
rect 1200 1111 1204 1115
rect 1344 1111 1348 1115
rect 1488 1111 1492 1115
rect 1632 1111 1636 1115
rect 1776 1111 1780 1115
rect 1912 1111 1916 1115
rect 2848 1111 2852 1115
rect 3024 1111 3028 1115
rect 3208 1111 3212 1115
rect 3400 1111 3404 1115
rect 3592 1111 3596 1115
rect 3776 1111 3780 1115
rect 4136 1111 4140 1115
rect 4336 1111 4340 1115
rect 4560 1111 4564 1115
rect 4816 1111 4820 1115
rect 5088 1111 5092 1115
rect 5376 1111 5380 1115
rect 5640 1111 5644 1115
rect 272 1043 276 1047
rect 512 1043 516 1047
rect 736 1043 740 1047
rect 952 1043 956 1047
rect 1152 1043 1156 1047
rect 1336 1043 1340 1047
rect 1520 1043 1524 1047
rect 1704 1043 1708 1047
rect 1888 1043 1892 1047
rect 2656 1039 2660 1043
rect 2848 1039 2852 1043
rect 3048 1039 3052 1043
rect 3248 1039 3252 1043
rect 3456 1039 3460 1043
rect 3672 1039 3676 1043
rect 4192 1039 4196 1043
rect 4488 1039 4492 1043
rect 4784 1039 4788 1043
rect 5072 1039 5076 1043
rect 5360 1039 5364 1043
rect 5640 1041 5644 1045
rect 5176 939 5180 943
rect 5176 879 5180 883
rect 320 871 324 875
rect 544 871 548 875
rect 792 871 796 875
rect 1056 872 1060 876
rect 2120 875 2124 879
rect 2344 875 2348 879
rect 2592 875 2596 879
rect 2832 875 2836 879
rect 3064 875 3068 879
rect 3296 875 3300 879
rect 3536 875 3540 879
rect 1344 871 1348 875
rect 1640 871 1644 875
rect 1912 871 1916 875
rect 4056 871 4060 875
rect 4280 871 4284 875
rect 4504 871 4508 875
rect 4720 871 4724 875
rect 4936 871 4940 875
rect 5152 871 5156 875
rect 5368 873 5372 877
rect 5592 871 5596 875
rect 2320 815 2324 819
rect 2536 815 2540 819
rect 2760 815 2764 819
rect 2984 815 2988 819
rect 3208 815 3212 819
rect 3432 815 3436 819
rect 3656 815 3660 819
rect 3984 811 3988 815
rect 4208 811 4212 815
rect 4440 811 4444 815
rect 4496 811 4500 815
rect 4672 811 4676 815
rect 4896 811 4900 815
rect 5128 811 5132 815
rect 5360 811 5364 815
rect 5592 811 5596 815
rect 320 787 324 791
rect 544 787 548 791
rect 760 787 764 791
rect 976 787 980 791
rect 1184 787 1188 791
rect 1392 787 1396 791
rect 1608 787 1612 791
rect 4496 747 4500 751
rect 3648 703 3652 707
rect 3984 647 3988 651
rect 4208 647 4212 651
rect 4448 647 4452 651
rect 4680 647 4684 651
rect 4904 647 4908 651
rect 5128 647 5132 651
rect 5352 647 5356 651
rect 5584 647 5588 651
rect 3648 639 3652 643
rect 3504 635 3508 639
rect 3640 635 3644 639
rect 3776 635 3780 639
rect 256 615 260 619
rect 400 615 404 619
rect 568 615 572 619
rect 736 615 740 619
rect 896 615 900 619
rect 1048 615 1052 619
rect 1200 615 1204 619
rect 1344 615 1348 619
rect 1488 615 1492 619
rect 1632 615 1636 619
rect 1776 615 1780 619
rect 1912 615 1916 619
rect 3984 579 3988 583
rect 4240 579 4244 583
rect 4504 579 4508 583
rect 4744 579 4748 583
rect 4976 579 4980 583
rect 5192 579 5196 583
rect 5408 579 5412 583
rect 5624 579 5628 583
rect 3368 567 3372 571
rect 3504 567 3508 571
rect 3640 567 3644 571
rect 3776 567 3780 571
rect 256 543 260 547
rect 472 543 476 547
rect 696 543 700 547
rect 904 543 908 547
rect 1096 543 1100 547
rect 1272 543 1276 547
rect 1440 543 1444 547
rect 1608 543 1612 547
rect 1768 543 1772 547
rect 1912 543 1916 547
rect 336 479 340 483
rect 608 455 612 459
rect 944 447 948 451
rect 4016 399 4020 403
rect 4296 399 4300 403
rect 4560 399 4564 403
rect 4808 399 4812 403
rect 5032 399 5036 403
rect 5248 399 5252 403
rect 5456 399 5460 403
rect 5640 399 5644 403
rect 944 387 948 391
rect 320 379 324 383
rect 336 379 340 383
rect 600 379 604 383
rect 608 379 612 383
rect 880 379 884 383
rect 1168 379 1172 383
rect 1456 381 1460 385
rect 2120 383 2124 387
rect 2280 383 2284 387
rect 2472 383 2476 387
rect 2664 383 2668 387
rect 2864 383 2868 387
rect 3056 383 3060 387
rect 3256 383 3260 387
rect 3456 383 3460 387
rect 3656 383 3660 387
rect 4104 335 4108 339
rect 4296 335 4300 339
rect 4520 335 4524 339
rect 4776 335 4780 339
rect 5064 335 5068 339
rect 5360 335 5364 339
rect 5640 335 5644 339
rect 408 319 412 323
rect 600 319 604 323
rect 792 319 796 323
rect 800 319 804 323
rect 984 319 988 323
rect 992 319 996 323
rect 1176 319 1180 323
rect 2120 299 2124 303
rect 2256 299 2260 303
rect 2392 299 2396 303
rect 2528 299 2532 303
rect 2664 299 2668 303
rect 2800 299 2804 303
rect 2936 299 2940 303
rect 3072 299 3076 303
rect 3208 299 3212 303
rect 3344 299 3348 303
rect 3480 299 3484 303
rect 3616 299 3620 303
rect 992 255 996 259
rect 800 187 804 191
rect 256 119 260 123
rect 392 119 396 123
rect 528 119 532 123
rect 664 119 668 123
rect 800 121 804 125
rect 936 119 940 123
rect 1072 119 1076 123
rect 1208 119 1212 123
rect 3984 119 3988 123
rect 4120 119 4124 123
rect 4256 119 4260 123
rect 4392 119 4396 123
rect 4560 119 4564 123
rect 4752 119 4756 123
rect 4968 119 4972 123
rect 5192 119 5196 123
rect 5640 121 5644 125
rect 2120 103 2124 107
rect 2256 103 2260 107
rect 2392 103 2396 107
rect 2528 103 2532 107
rect 2664 103 2668 107
rect 2800 103 2804 107
rect 2936 103 2940 107
rect 3072 103 3076 107
rect 3208 103 3212 107
rect 3344 103 3348 107
rect 3480 103 3484 107
rect 3616 103 3620 107
rect 3752 103 3756 107
<< m2 >>
rect 1678 5747 1684 5748
rect 1678 5746 1679 5747
rect 1432 5744 1679 5746
rect 1432 5742 1434 5744
rect 1678 5743 1679 5744
rect 1683 5743 1684 5747
rect 1678 5742 1684 5743
rect 1277 5740 1434 5742
rect 378 5739 384 5740
rect 378 5735 379 5739
rect 383 5735 384 5739
rect 378 5734 384 5735
rect 642 5739 648 5740
rect 642 5735 643 5739
rect 647 5735 648 5739
rect 642 5734 648 5735
rect 914 5739 920 5740
rect 914 5735 915 5739
rect 919 5735 920 5739
rect 914 5734 920 5735
rect 1458 5739 1464 5740
rect 1458 5735 1459 5739
rect 1463 5735 1464 5739
rect 1458 5734 1464 5735
rect 1730 5739 1736 5740
rect 1730 5735 1731 5739
rect 1735 5735 1736 5739
rect 1730 5734 1736 5735
rect 1974 5693 1980 5694
rect 3798 5693 3804 5694
rect 110 5692 116 5693
rect 1934 5692 1940 5693
rect 110 5688 111 5692
rect 115 5688 116 5692
rect 110 5687 116 5688
rect 130 5691 136 5692
rect 130 5687 131 5691
rect 135 5687 136 5691
rect 130 5686 136 5687
rect 370 5691 376 5692
rect 370 5687 371 5691
rect 375 5687 376 5691
rect 370 5686 376 5687
rect 634 5691 640 5692
rect 634 5687 635 5691
rect 639 5687 640 5691
rect 634 5686 640 5687
rect 906 5691 912 5692
rect 906 5687 907 5691
rect 911 5687 912 5691
rect 906 5686 912 5687
rect 1178 5691 1184 5692
rect 1178 5687 1179 5691
rect 1183 5687 1184 5691
rect 1178 5686 1184 5687
rect 1450 5691 1456 5692
rect 1450 5687 1451 5691
rect 1455 5687 1456 5691
rect 1450 5686 1456 5687
rect 1722 5691 1728 5692
rect 1722 5687 1723 5691
rect 1727 5687 1728 5691
rect 1934 5688 1935 5692
rect 1939 5688 1940 5692
rect 1974 5689 1975 5693
rect 1979 5689 1980 5693
rect 1974 5688 1980 5689
rect 2510 5692 2516 5693
rect 2662 5692 2668 5693
rect 2814 5692 2820 5693
rect 2974 5692 2980 5693
rect 3142 5692 3148 5693
rect 3318 5692 3324 5693
rect 3494 5692 3500 5693
rect 2510 5688 2511 5692
rect 2515 5688 2516 5692
rect 1934 5687 1940 5688
rect 2510 5687 2516 5688
rect 2607 5691 2613 5692
rect 2607 5687 2608 5691
rect 2612 5690 2613 5691
rect 2623 5691 2629 5692
rect 2623 5690 2624 5691
rect 2612 5688 2624 5690
rect 2612 5687 2613 5688
rect 1722 5686 1728 5687
rect 2607 5686 2613 5687
rect 2623 5687 2624 5688
rect 2628 5687 2629 5691
rect 2662 5688 2663 5692
rect 2667 5688 2668 5692
rect 2662 5687 2668 5688
rect 2754 5691 2765 5692
rect 2754 5687 2755 5691
rect 2759 5687 2760 5691
rect 2764 5687 2765 5691
rect 2814 5688 2815 5692
rect 2819 5688 2820 5692
rect 2814 5687 2820 5688
rect 2906 5691 2917 5692
rect 2906 5687 2907 5691
rect 2911 5687 2912 5691
rect 2916 5687 2917 5691
rect 2974 5688 2975 5692
rect 2979 5688 2980 5692
rect 2974 5687 2980 5688
rect 3070 5691 3077 5692
rect 3070 5687 3071 5691
rect 3076 5687 3077 5691
rect 3142 5688 3143 5692
rect 3147 5688 3148 5692
rect 3142 5687 3148 5688
rect 3238 5691 3245 5692
rect 3238 5687 3239 5691
rect 3244 5687 3245 5691
rect 3318 5688 3319 5692
rect 3323 5688 3324 5692
rect 3318 5687 3324 5688
rect 3414 5691 3421 5692
rect 3414 5687 3415 5691
rect 3420 5687 3421 5691
rect 3494 5688 3495 5692
rect 3499 5688 3500 5692
rect 3494 5687 3500 5688
rect 3590 5691 3597 5692
rect 3590 5687 3591 5691
rect 3596 5687 3597 5691
rect 3798 5689 3799 5693
rect 3803 5689 3804 5693
rect 3798 5688 3804 5689
rect 2623 5686 2629 5687
rect 2754 5686 2765 5687
rect 2906 5686 2917 5687
rect 3070 5686 3077 5687
rect 3238 5686 3245 5687
rect 3414 5686 3421 5687
rect 3590 5686 3597 5687
rect 2482 5677 2488 5678
rect 158 5676 164 5677
rect 398 5676 404 5677
rect 662 5676 668 5677
rect 934 5676 940 5677
rect 1206 5676 1212 5677
rect 1478 5676 1484 5677
rect 1750 5676 1756 5677
rect 1974 5676 1980 5677
rect 110 5675 116 5676
rect 110 5671 111 5675
rect 115 5671 116 5675
rect 158 5672 159 5676
rect 163 5672 164 5676
rect 158 5671 164 5672
rect 255 5675 261 5676
rect 255 5671 256 5675
rect 260 5674 261 5675
rect 378 5675 384 5676
rect 378 5674 379 5675
rect 260 5672 379 5674
rect 260 5671 261 5672
rect 110 5670 116 5671
rect 255 5670 261 5671
rect 378 5671 379 5672
rect 383 5671 384 5675
rect 398 5672 399 5676
rect 403 5672 404 5676
rect 398 5671 404 5672
rect 495 5675 501 5676
rect 495 5671 496 5675
rect 500 5674 501 5675
rect 642 5675 648 5676
rect 642 5674 643 5675
rect 500 5672 643 5674
rect 500 5671 501 5672
rect 378 5670 384 5671
rect 495 5670 501 5671
rect 642 5671 643 5672
rect 647 5671 648 5675
rect 662 5672 663 5676
rect 667 5672 668 5676
rect 662 5671 668 5672
rect 759 5675 765 5676
rect 759 5671 760 5675
rect 764 5674 765 5675
rect 914 5675 920 5676
rect 914 5674 915 5675
rect 764 5672 915 5674
rect 764 5671 765 5672
rect 642 5670 648 5671
rect 759 5670 765 5671
rect 914 5671 915 5672
rect 919 5671 920 5675
rect 934 5672 935 5676
rect 939 5672 940 5676
rect 934 5671 940 5672
rect 1030 5675 1037 5676
rect 1030 5671 1031 5675
rect 1036 5671 1037 5675
rect 1206 5672 1207 5676
rect 1211 5672 1212 5676
rect 1206 5671 1212 5672
rect 1303 5675 1309 5676
rect 1303 5671 1304 5675
rect 1308 5674 1309 5675
rect 1458 5675 1464 5676
rect 1458 5674 1459 5675
rect 1308 5672 1459 5674
rect 1308 5671 1309 5672
rect 914 5670 920 5671
rect 1030 5670 1037 5671
rect 1303 5670 1309 5671
rect 1458 5671 1459 5672
rect 1463 5671 1464 5675
rect 1478 5672 1479 5676
rect 1483 5672 1484 5676
rect 1478 5671 1484 5672
rect 1575 5675 1581 5676
rect 1575 5671 1576 5675
rect 1580 5674 1581 5675
rect 1730 5675 1736 5676
rect 1730 5674 1731 5675
rect 1580 5672 1731 5674
rect 1580 5671 1581 5672
rect 1458 5670 1464 5671
rect 1575 5670 1581 5671
rect 1730 5671 1731 5672
rect 1735 5671 1736 5675
rect 1750 5672 1751 5676
rect 1755 5672 1756 5676
rect 1750 5671 1756 5672
rect 1846 5675 1853 5676
rect 1846 5671 1847 5675
rect 1852 5671 1853 5675
rect 1730 5670 1736 5671
rect 1846 5670 1853 5671
rect 1934 5675 1940 5676
rect 1934 5671 1935 5675
rect 1939 5671 1940 5675
rect 1974 5672 1975 5676
rect 1979 5672 1980 5676
rect 2482 5673 2483 5677
rect 2487 5673 2488 5677
rect 2482 5672 2488 5673
rect 2634 5677 2640 5678
rect 2634 5673 2635 5677
rect 2639 5673 2640 5677
rect 2634 5672 2640 5673
rect 2786 5677 2792 5678
rect 2786 5673 2787 5677
rect 2791 5673 2792 5677
rect 2786 5672 2792 5673
rect 2946 5677 2952 5678
rect 2946 5673 2947 5677
rect 2951 5673 2952 5677
rect 2946 5672 2952 5673
rect 3114 5677 3120 5678
rect 3114 5673 3115 5677
rect 3119 5673 3120 5677
rect 3114 5672 3120 5673
rect 3290 5677 3296 5678
rect 3290 5673 3291 5677
rect 3295 5673 3296 5677
rect 3290 5672 3296 5673
rect 3466 5677 3472 5678
rect 3466 5673 3467 5677
rect 3471 5673 3472 5677
rect 3466 5672 3472 5673
rect 3798 5676 3804 5677
rect 3798 5672 3799 5676
rect 3803 5672 3804 5676
rect 1974 5671 1980 5672
rect 3210 5671 3216 5672
rect 1934 5670 1940 5671
rect 3210 5667 3211 5671
rect 3215 5670 3216 5671
rect 3414 5671 3420 5672
rect 3798 5671 3804 5672
rect 3414 5670 3415 5671
rect 3215 5668 3415 5670
rect 3215 5667 3216 5668
rect 3210 5666 3216 5667
rect 3414 5667 3415 5668
rect 3419 5667 3420 5671
rect 3414 5666 3420 5667
rect 4202 5655 4208 5656
rect 4202 5651 4203 5655
rect 4207 5651 4208 5655
rect 4202 5650 4208 5651
rect 4250 5655 4256 5656
rect 4250 5651 4251 5655
rect 4255 5651 4256 5655
rect 4250 5650 4256 5651
rect 4386 5655 4392 5656
rect 4386 5651 4387 5655
rect 4391 5651 4392 5655
rect 4386 5650 4392 5651
rect 4522 5655 4528 5656
rect 4522 5651 4523 5655
rect 4527 5651 4528 5655
rect 4522 5650 4528 5651
rect 4658 5655 4664 5656
rect 4658 5651 4659 5655
rect 4663 5651 4664 5655
rect 4658 5650 4664 5651
rect 4794 5655 4800 5656
rect 4794 5651 4795 5655
rect 4799 5651 4800 5655
rect 4794 5650 4800 5651
rect 4930 5655 4936 5656
rect 4930 5651 4931 5655
rect 4935 5651 4936 5655
rect 4930 5650 4936 5651
rect 5066 5655 5072 5656
rect 5066 5651 5067 5655
rect 5071 5651 5072 5655
rect 5066 5650 5072 5651
rect 5202 5655 5208 5656
rect 5202 5651 5203 5655
rect 5207 5651 5208 5655
rect 5202 5650 5208 5651
rect 2623 5627 2629 5628
rect 2580 5618 2582 5625
rect 2623 5623 2624 5627
rect 2628 5626 2629 5627
rect 3210 5627 3216 5628
rect 2628 5624 2641 5626
rect 2885 5624 2930 5626
rect 3045 5624 3114 5626
rect 2628 5623 2629 5624
rect 2623 5622 2629 5623
rect 2906 5619 2912 5620
rect 2906 5618 2907 5619
rect 110 5617 116 5618
rect 1934 5617 1940 5618
rect 110 5613 111 5617
rect 115 5613 116 5617
rect 110 5612 116 5613
rect 454 5616 460 5617
rect 646 5616 652 5617
rect 854 5616 860 5617
rect 1086 5616 1092 5617
rect 1326 5616 1332 5617
rect 1582 5616 1588 5617
rect 1814 5616 1820 5617
rect 454 5612 455 5616
rect 459 5612 460 5616
rect 454 5611 460 5612
rect 551 5615 557 5616
rect 551 5611 552 5615
rect 556 5614 557 5615
rect 583 5615 589 5616
rect 583 5614 584 5615
rect 556 5612 584 5614
rect 556 5611 557 5612
rect 551 5610 557 5611
rect 583 5611 584 5612
rect 588 5611 589 5615
rect 646 5612 647 5616
rect 651 5612 652 5616
rect 646 5611 652 5612
rect 743 5615 752 5616
rect 743 5611 744 5615
rect 751 5611 752 5615
rect 854 5612 855 5616
rect 859 5612 860 5616
rect 854 5611 860 5612
rect 951 5615 957 5616
rect 951 5611 952 5615
rect 956 5614 957 5615
rect 966 5615 972 5616
rect 966 5614 967 5615
rect 956 5612 967 5614
rect 956 5611 957 5612
rect 583 5610 589 5611
rect 743 5610 752 5611
rect 951 5610 957 5611
rect 966 5611 967 5612
rect 971 5611 972 5615
rect 1086 5612 1087 5616
rect 1091 5612 1092 5616
rect 1086 5611 1092 5612
rect 1178 5615 1189 5616
rect 1178 5611 1179 5615
rect 1183 5611 1184 5615
rect 1188 5611 1189 5615
rect 1326 5612 1327 5616
rect 1331 5612 1332 5616
rect 1326 5611 1332 5612
rect 1423 5615 1429 5616
rect 1423 5611 1424 5615
rect 1428 5614 1429 5615
rect 1463 5615 1469 5616
rect 1463 5614 1464 5615
rect 1428 5612 1464 5614
rect 1428 5611 1429 5612
rect 966 5610 972 5611
rect 1178 5610 1189 5611
rect 1423 5610 1429 5611
rect 1463 5611 1464 5612
rect 1468 5611 1469 5615
rect 1582 5612 1583 5616
rect 1587 5612 1588 5616
rect 1582 5611 1588 5612
rect 1678 5615 1685 5616
rect 1678 5611 1679 5615
rect 1684 5611 1685 5615
rect 1814 5612 1815 5616
rect 1819 5612 1820 5616
rect 1814 5611 1820 5612
rect 1911 5615 1917 5616
rect 1911 5611 1912 5615
rect 1916 5614 1917 5615
rect 1926 5615 1932 5616
rect 1926 5614 1927 5615
rect 1916 5612 1927 5614
rect 1916 5611 1917 5612
rect 1463 5610 1469 5611
rect 1678 5610 1685 5611
rect 1911 5610 1917 5611
rect 1926 5611 1927 5612
rect 1931 5611 1932 5615
rect 1934 5613 1935 5617
rect 1939 5613 1940 5617
rect 2580 5616 2907 5618
rect 2906 5615 2907 5616
rect 2911 5615 2912 5619
rect 2928 5618 2930 5624
rect 3070 5619 3076 5620
rect 3070 5618 3071 5619
rect 2928 5616 3071 5618
rect 2906 5614 2912 5615
rect 3070 5615 3071 5616
rect 3075 5615 3076 5619
rect 3112 5618 3114 5624
rect 3210 5623 3211 5627
rect 3215 5623 3216 5627
rect 3774 5627 3780 5628
rect 3774 5626 3775 5627
rect 3210 5622 3216 5623
rect 3238 5619 3244 5620
rect 3238 5618 3239 5619
rect 3112 5616 3239 5618
rect 3070 5614 3076 5615
rect 3238 5615 3239 5616
rect 3243 5615 3244 5619
rect 3388 5618 3390 5625
rect 3565 5624 3775 5626
rect 3774 5623 3775 5624
rect 3779 5623 3780 5627
rect 3774 5622 3780 5623
rect 3590 5619 3596 5620
rect 3590 5618 3591 5619
rect 3388 5616 3591 5618
rect 3238 5614 3244 5615
rect 3590 5615 3591 5616
rect 3595 5615 3596 5619
rect 3590 5614 3596 5615
rect 1934 5612 1940 5613
rect 1926 5610 1932 5611
rect 3838 5608 3844 5609
rect 5662 5608 5668 5609
rect 3838 5604 3839 5608
rect 3843 5604 3844 5608
rect 3838 5603 3844 5604
rect 4106 5607 4112 5608
rect 4106 5603 4107 5607
rect 4111 5603 4112 5607
rect 4106 5602 4112 5603
rect 4242 5607 4248 5608
rect 4242 5603 4243 5607
rect 4247 5603 4248 5607
rect 4242 5602 4248 5603
rect 4378 5607 4384 5608
rect 4378 5603 4379 5607
rect 4383 5603 4384 5607
rect 4378 5602 4384 5603
rect 4514 5607 4520 5608
rect 4514 5603 4515 5607
rect 4519 5603 4520 5607
rect 4514 5602 4520 5603
rect 4650 5607 4656 5608
rect 4650 5603 4651 5607
rect 4655 5603 4656 5607
rect 4650 5602 4656 5603
rect 4786 5607 4792 5608
rect 4786 5603 4787 5607
rect 4791 5603 4792 5607
rect 4786 5602 4792 5603
rect 4922 5607 4928 5608
rect 4922 5603 4923 5607
rect 4927 5603 4928 5607
rect 4922 5602 4928 5603
rect 5058 5607 5064 5608
rect 5058 5603 5059 5607
rect 5063 5603 5064 5607
rect 5058 5602 5064 5603
rect 5194 5607 5200 5608
rect 5194 5603 5195 5607
rect 5199 5603 5200 5607
rect 5662 5604 5663 5608
rect 5667 5604 5668 5608
rect 5662 5603 5668 5604
rect 5194 5602 5200 5603
rect 426 5601 432 5602
rect 110 5600 116 5601
rect 110 5596 111 5600
rect 115 5596 116 5600
rect 426 5597 427 5601
rect 431 5597 432 5601
rect 426 5596 432 5597
rect 618 5601 624 5602
rect 618 5597 619 5601
rect 623 5597 624 5601
rect 618 5596 624 5597
rect 826 5601 832 5602
rect 826 5597 827 5601
rect 831 5597 832 5601
rect 826 5596 832 5597
rect 1058 5601 1064 5602
rect 1058 5597 1059 5601
rect 1063 5597 1064 5601
rect 1058 5596 1064 5597
rect 1298 5601 1304 5602
rect 1298 5597 1299 5601
rect 1303 5597 1304 5601
rect 1298 5596 1304 5597
rect 1554 5601 1560 5602
rect 1554 5597 1555 5601
rect 1559 5597 1560 5601
rect 1554 5596 1560 5597
rect 1786 5601 1792 5602
rect 1786 5597 1787 5601
rect 1791 5597 1792 5601
rect 1786 5596 1792 5597
rect 1934 5600 1940 5601
rect 1934 5596 1935 5600
rect 1939 5596 1940 5600
rect 110 5595 116 5596
rect 1934 5595 1940 5596
rect 2778 5595 2784 5596
rect 2778 5594 2779 5595
rect 2436 5592 2779 5594
rect 1926 5587 1932 5588
rect 1926 5583 1927 5587
rect 1931 5586 1932 5587
rect 2436 5586 2438 5592
rect 2778 5591 2779 5592
rect 2783 5591 2784 5595
rect 4134 5592 4140 5593
rect 4270 5592 4276 5593
rect 4406 5592 4412 5593
rect 4542 5592 4548 5593
rect 4678 5592 4684 5593
rect 4814 5592 4820 5593
rect 4950 5592 4956 5593
rect 5086 5592 5092 5593
rect 5222 5592 5228 5593
rect 2778 5590 2784 5591
rect 3838 5591 3844 5592
rect 1931 5584 2001 5586
rect 2301 5584 2438 5586
rect 2754 5587 2760 5588
rect 1931 5583 1932 5584
rect 1926 5582 1932 5583
rect 2442 5583 2448 5584
rect 2442 5579 2443 5583
rect 2447 5579 2448 5583
rect 2754 5583 2755 5587
rect 2759 5583 2760 5587
rect 3071 5587 3077 5588
rect 3071 5586 3072 5587
rect 2965 5584 3072 5586
rect 2754 5582 2760 5583
rect 3071 5583 3072 5584
rect 3076 5583 3077 5587
rect 3838 5587 3839 5591
rect 3843 5587 3844 5591
rect 4134 5588 4135 5592
rect 4139 5588 4140 5592
rect 4134 5587 4140 5588
rect 4231 5591 4237 5592
rect 4231 5587 4232 5591
rect 4236 5590 4237 5591
rect 4250 5591 4256 5592
rect 4250 5590 4251 5591
rect 4236 5588 4251 5590
rect 4236 5587 4237 5588
rect 3838 5586 3844 5587
rect 4231 5586 4237 5587
rect 4250 5587 4251 5588
rect 4255 5587 4256 5591
rect 4270 5588 4271 5592
rect 4275 5588 4276 5592
rect 4270 5587 4276 5588
rect 4367 5591 4373 5592
rect 4367 5587 4368 5591
rect 4372 5590 4373 5591
rect 4386 5591 4392 5592
rect 4386 5590 4387 5591
rect 4372 5588 4387 5590
rect 4372 5587 4373 5588
rect 4250 5586 4256 5587
rect 4367 5586 4373 5587
rect 4386 5587 4387 5588
rect 4391 5587 4392 5591
rect 4406 5588 4407 5592
rect 4411 5588 4412 5592
rect 4406 5587 4412 5588
rect 4503 5591 4509 5592
rect 4503 5587 4504 5591
rect 4508 5590 4509 5591
rect 4522 5591 4528 5592
rect 4522 5590 4523 5591
rect 4508 5588 4523 5590
rect 4508 5587 4509 5588
rect 4386 5586 4392 5587
rect 4503 5586 4509 5587
rect 4522 5587 4523 5588
rect 4527 5587 4528 5591
rect 4542 5588 4543 5592
rect 4547 5588 4548 5592
rect 4542 5587 4548 5588
rect 4639 5591 4645 5592
rect 4639 5587 4640 5591
rect 4644 5590 4645 5591
rect 4658 5591 4664 5592
rect 4658 5590 4659 5591
rect 4644 5588 4659 5590
rect 4644 5587 4645 5588
rect 4522 5586 4528 5587
rect 4639 5586 4645 5587
rect 4658 5587 4659 5588
rect 4663 5587 4664 5591
rect 4678 5588 4679 5592
rect 4683 5588 4684 5592
rect 4678 5587 4684 5588
rect 4775 5591 4781 5592
rect 4775 5587 4776 5591
rect 4780 5590 4781 5591
rect 4794 5591 4800 5592
rect 4794 5590 4795 5591
rect 4780 5588 4795 5590
rect 4780 5587 4781 5588
rect 4658 5586 4664 5587
rect 4775 5586 4781 5587
rect 4794 5587 4795 5588
rect 4799 5587 4800 5591
rect 4814 5588 4815 5592
rect 4819 5588 4820 5592
rect 4814 5587 4820 5588
rect 4911 5591 4917 5592
rect 4911 5587 4912 5591
rect 4916 5590 4917 5591
rect 4930 5591 4936 5592
rect 4930 5590 4931 5591
rect 4916 5588 4931 5590
rect 4916 5587 4917 5588
rect 4794 5586 4800 5587
rect 4911 5586 4917 5587
rect 4930 5587 4931 5588
rect 4935 5587 4936 5591
rect 4950 5588 4951 5592
rect 4955 5588 4956 5592
rect 4950 5587 4956 5588
rect 5047 5591 5053 5592
rect 5047 5587 5048 5591
rect 5052 5590 5053 5591
rect 5066 5591 5072 5592
rect 5066 5590 5067 5591
rect 5052 5588 5067 5590
rect 5052 5587 5053 5588
rect 4930 5586 4936 5587
rect 5047 5586 5053 5587
rect 5066 5587 5067 5588
rect 5071 5587 5072 5591
rect 5086 5588 5087 5592
rect 5091 5588 5092 5592
rect 5086 5587 5092 5588
rect 5183 5591 5189 5592
rect 5183 5587 5184 5591
rect 5188 5590 5189 5591
rect 5202 5591 5208 5592
rect 5202 5590 5203 5591
rect 5188 5588 5203 5590
rect 5188 5587 5189 5588
rect 5066 5586 5072 5587
rect 5183 5586 5189 5587
rect 5202 5587 5203 5588
rect 5207 5587 5208 5591
rect 5222 5588 5223 5592
rect 5227 5588 5228 5592
rect 5222 5587 5228 5588
rect 5314 5591 5325 5592
rect 5314 5587 5315 5591
rect 5319 5587 5320 5591
rect 5324 5587 5325 5591
rect 5202 5586 5208 5587
rect 5314 5586 5325 5587
rect 5662 5591 5668 5592
rect 5662 5587 5663 5591
rect 5667 5587 5668 5591
rect 5662 5586 5668 5587
rect 3071 5582 3077 5583
rect 3082 5583 3088 5584
rect 2442 5578 2448 5579
rect 3082 5579 3083 5583
rect 3087 5579 3088 5583
rect 3082 5578 3088 5579
rect 3282 5583 3288 5584
rect 3282 5579 3283 5583
rect 3287 5579 3288 5583
rect 3282 5578 3288 5579
rect 3482 5583 3488 5584
rect 3482 5579 3483 5583
rect 3487 5579 3488 5583
rect 3482 5578 3488 5579
rect 3658 5583 3664 5584
rect 3658 5579 3659 5583
rect 3663 5579 3664 5583
rect 3658 5578 3664 5579
rect 4202 5559 4208 5560
rect 4202 5555 4203 5559
rect 4207 5558 4208 5559
rect 4398 5559 4404 5560
rect 4398 5558 4399 5559
rect 4207 5556 4399 5558
rect 4207 5555 4208 5556
rect 4202 5554 4208 5555
rect 4398 5555 4399 5556
rect 4403 5555 4404 5559
rect 4398 5554 4404 5555
rect 583 5551 589 5552
rect 524 5542 526 5549
rect 583 5547 584 5551
rect 588 5550 589 5551
rect 746 5551 752 5552
rect 588 5548 625 5550
rect 588 5547 589 5548
rect 583 5546 589 5547
rect 746 5547 747 5551
rect 751 5550 752 5551
rect 966 5551 972 5552
rect 751 5548 833 5550
rect 751 5547 752 5548
rect 746 5546 752 5547
rect 966 5547 967 5551
rect 971 5550 972 5551
rect 1318 5551 1324 5552
rect 971 5548 1065 5550
rect 971 5547 972 5548
rect 966 5546 972 5547
rect 1318 5547 1319 5551
rect 1323 5547 1324 5551
rect 1318 5546 1324 5547
rect 1463 5551 1469 5552
rect 1463 5547 1464 5551
rect 1468 5550 1469 5551
rect 1846 5551 1852 5552
rect 1468 5548 1561 5550
rect 1468 5547 1469 5548
rect 1463 5546 1469 5547
rect 1846 5547 1847 5551
rect 1851 5547 1852 5551
rect 1846 5546 1852 5547
rect 1030 5543 1036 5544
rect 1030 5542 1031 5543
rect 524 5540 1031 5542
rect 1030 5539 1031 5540
rect 1035 5539 1036 5543
rect 1030 5538 1036 5539
rect 1974 5536 1980 5537
rect 3798 5536 3804 5537
rect 1974 5532 1975 5536
rect 1979 5532 1980 5536
rect 1974 5531 1980 5532
rect 1994 5535 2000 5536
rect 1994 5531 1995 5535
rect 1999 5531 2000 5535
rect 1994 5530 2000 5531
rect 2202 5535 2208 5536
rect 2202 5531 2203 5535
rect 2207 5531 2208 5535
rect 2202 5530 2208 5531
rect 2434 5535 2440 5536
rect 2434 5531 2435 5535
rect 2439 5531 2440 5535
rect 2434 5530 2440 5531
rect 2658 5535 2664 5536
rect 2658 5531 2659 5535
rect 2663 5531 2664 5535
rect 2658 5530 2664 5531
rect 2866 5535 2872 5536
rect 2866 5531 2867 5535
rect 2871 5531 2872 5535
rect 2866 5530 2872 5531
rect 3074 5535 3080 5536
rect 3074 5531 3075 5535
rect 3079 5531 3080 5535
rect 3074 5530 3080 5531
rect 3274 5535 3280 5536
rect 3274 5531 3275 5535
rect 3279 5531 3280 5535
rect 3274 5530 3280 5531
rect 3474 5535 3480 5536
rect 3474 5531 3475 5535
rect 3479 5531 3480 5535
rect 3474 5530 3480 5531
rect 3650 5535 3656 5536
rect 3650 5531 3651 5535
rect 3655 5531 3656 5535
rect 3798 5532 3799 5536
rect 3803 5532 3804 5536
rect 3798 5531 3804 5532
rect 3650 5530 3656 5531
rect 2022 5520 2028 5521
rect 2230 5520 2236 5521
rect 2462 5520 2468 5521
rect 2686 5520 2692 5521
rect 2894 5520 2900 5521
rect 3102 5520 3108 5521
rect 3302 5520 3308 5521
rect 3502 5520 3508 5521
rect 3678 5520 3684 5521
rect 882 5519 888 5520
rect 882 5515 883 5519
rect 887 5515 888 5519
rect 1974 5519 1980 5520
rect 882 5514 888 5515
rect 930 5515 936 5516
rect 930 5511 931 5515
rect 935 5511 936 5515
rect 930 5510 936 5511
rect 1066 5515 1072 5516
rect 1066 5511 1067 5515
rect 1071 5511 1072 5515
rect 1066 5510 1072 5511
rect 1202 5515 1208 5516
rect 1202 5511 1203 5515
rect 1207 5511 1208 5515
rect 1202 5510 1208 5511
rect 1426 5515 1432 5516
rect 1426 5511 1427 5515
rect 1431 5511 1432 5515
rect 1974 5515 1975 5519
rect 1979 5515 1980 5519
rect 2022 5516 2023 5520
rect 2027 5516 2028 5520
rect 2022 5515 2028 5516
rect 2119 5519 2128 5520
rect 2119 5515 2120 5519
rect 2127 5515 2128 5519
rect 2230 5516 2231 5520
rect 2235 5516 2236 5520
rect 2230 5515 2236 5516
rect 2327 5519 2333 5520
rect 2327 5515 2328 5519
rect 2332 5518 2333 5519
rect 2442 5519 2448 5520
rect 2442 5518 2443 5519
rect 2332 5516 2443 5518
rect 2332 5515 2333 5516
rect 1974 5514 1980 5515
rect 2119 5514 2128 5515
rect 2327 5514 2333 5515
rect 2442 5515 2443 5516
rect 2447 5515 2448 5519
rect 2462 5516 2463 5520
rect 2467 5516 2468 5520
rect 2462 5515 2468 5516
rect 2558 5519 2565 5520
rect 2558 5515 2559 5519
rect 2564 5515 2565 5519
rect 2686 5516 2687 5520
rect 2691 5516 2692 5520
rect 2686 5515 2692 5516
rect 2778 5519 2789 5520
rect 2778 5515 2779 5519
rect 2783 5515 2784 5519
rect 2788 5515 2789 5519
rect 2894 5516 2895 5520
rect 2899 5516 2900 5520
rect 2894 5515 2900 5516
rect 2991 5519 2997 5520
rect 2991 5515 2992 5519
rect 2996 5518 2997 5519
rect 3082 5519 3088 5520
rect 3082 5518 3083 5519
rect 2996 5516 3083 5518
rect 2996 5515 2997 5516
rect 2442 5514 2448 5515
rect 2558 5514 2565 5515
rect 2778 5514 2789 5515
rect 2991 5514 2997 5515
rect 3082 5515 3083 5516
rect 3087 5515 3088 5519
rect 3102 5516 3103 5520
rect 3107 5516 3108 5520
rect 3102 5515 3108 5516
rect 3199 5519 3205 5520
rect 3199 5515 3200 5519
rect 3204 5518 3205 5519
rect 3282 5519 3288 5520
rect 3282 5518 3283 5519
rect 3204 5516 3283 5518
rect 3204 5515 3205 5516
rect 3082 5514 3088 5515
rect 3199 5514 3205 5515
rect 3282 5515 3283 5516
rect 3287 5515 3288 5519
rect 3302 5516 3303 5520
rect 3307 5516 3308 5520
rect 3302 5515 3308 5516
rect 3399 5519 3405 5520
rect 3399 5515 3400 5519
rect 3404 5518 3405 5519
rect 3482 5519 3488 5520
rect 3482 5518 3483 5519
rect 3404 5516 3483 5518
rect 3404 5515 3405 5516
rect 3282 5514 3288 5515
rect 3399 5514 3405 5515
rect 3482 5515 3483 5516
rect 3487 5515 3488 5519
rect 3502 5516 3503 5520
rect 3507 5516 3508 5520
rect 3502 5515 3508 5516
rect 3599 5519 3605 5520
rect 3599 5515 3600 5519
rect 3604 5518 3605 5519
rect 3658 5519 3664 5520
rect 3658 5518 3659 5519
rect 3604 5516 3659 5518
rect 3604 5515 3605 5516
rect 3482 5514 3488 5515
rect 3599 5514 3605 5515
rect 3658 5515 3659 5516
rect 3663 5515 3664 5519
rect 3678 5516 3679 5520
rect 3683 5516 3684 5520
rect 3678 5515 3684 5516
rect 3774 5519 3781 5520
rect 3774 5515 3775 5519
rect 3780 5515 3781 5519
rect 3658 5514 3664 5515
rect 3774 5514 3781 5515
rect 3798 5519 3804 5520
rect 3798 5515 3799 5519
rect 3803 5515 3804 5519
rect 3798 5514 3804 5515
rect 1426 5510 1432 5511
rect 3838 5501 3844 5502
rect 5662 5501 5668 5502
rect 3838 5497 3839 5501
rect 3843 5497 3844 5501
rect 3838 5496 3844 5497
rect 4302 5500 4308 5501
rect 4510 5500 4516 5501
rect 4718 5500 4724 5501
rect 4926 5500 4932 5501
rect 5134 5500 5140 5501
rect 4302 5496 4303 5500
rect 4307 5496 4308 5500
rect 4302 5495 4308 5496
rect 4398 5499 4405 5500
rect 4398 5495 4399 5499
rect 4404 5495 4405 5499
rect 4510 5496 4511 5500
rect 4515 5496 4516 5500
rect 4510 5495 4516 5496
rect 4602 5499 4613 5500
rect 4602 5495 4603 5499
rect 4607 5495 4608 5499
rect 4612 5495 4613 5499
rect 4718 5496 4719 5500
rect 4723 5496 4724 5500
rect 4718 5495 4724 5496
rect 4815 5499 4824 5500
rect 4815 5495 4816 5499
rect 4823 5495 4824 5499
rect 4926 5496 4927 5500
rect 4931 5496 4932 5500
rect 4926 5495 4932 5496
rect 5022 5499 5029 5500
rect 5022 5495 5023 5499
rect 5028 5495 5029 5499
rect 5134 5496 5135 5500
rect 5139 5496 5140 5500
rect 5134 5495 5140 5496
rect 5230 5499 5237 5500
rect 5230 5495 5231 5499
rect 5236 5495 5237 5499
rect 5662 5497 5663 5501
rect 5667 5497 5668 5501
rect 5662 5496 5668 5497
rect 4398 5494 4405 5495
rect 4602 5494 4613 5495
rect 4815 5494 4824 5495
rect 5022 5494 5029 5495
rect 5230 5494 5237 5495
rect 4274 5485 4280 5486
rect 3838 5484 3844 5485
rect 3838 5480 3839 5484
rect 3843 5480 3844 5484
rect 4274 5481 4275 5485
rect 4279 5481 4280 5485
rect 4274 5480 4280 5481
rect 4482 5485 4488 5486
rect 4482 5481 4483 5485
rect 4487 5481 4488 5485
rect 4482 5480 4488 5481
rect 4690 5485 4696 5486
rect 4690 5481 4691 5485
rect 4695 5481 4696 5485
rect 4690 5480 4696 5481
rect 4898 5485 4904 5486
rect 4898 5481 4899 5485
rect 4903 5481 4904 5485
rect 4898 5480 4904 5481
rect 5106 5485 5112 5486
rect 5106 5481 5107 5485
rect 5111 5481 5112 5485
rect 5106 5480 5112 5481
rect 5662 5484 5668 5485
rect 5662 5480 5663 5484
rect 5667 5480 5668 5484
rect 3838 5479 3844 5480
rect 5662 5479 5668 5480
rect 2135 5475 2141 5476
rect 2135 5471 2136 5475
rect 2140 5474 2141 5475
rect 3071 5475 3077 5476
rect 2140 5472 2814 5474
rect 2140 5471 2141 5472
rect 2135 5470 2141 5471
rect 110 5468 116 5469
rect 1934 5468 1940 5469
rect 110 5464 111 5468
rect 115 5464 116 5468
rect 110 5463 116 5464
rect 786 5467 792 5468
rect 786 5463 787 5467
rect 791 5463 792 5467
rect 786 5462 792 5463
rect 922 5467 928 5468
rect 922 5463 923 5467
rect 927 5463 928 5467
rect 922 5462 928 5463
rect 1058 5467 1064 5468
rect 1058 5463 1059 5467
rect 1063 5463 1064 5467
rect 1058 5462 1064 5463
rect 1194 5467 1200 5468
rect 1194 5463 1195 5467
rect 1199 5463 1200 5467
rect 1194 5462 1200 5463
rect 1330 5467 1336 5468
rect 1330 5463 1331 5467
rect 1335 5463 1336 5467
rect 1934 5464 1935 5468
rect 1939 5464 1940 5468
rect 2812 5466 2814 5472
rect 3071 5471 3072 5475
rect 3076 5474 3077 5475
rect 3076 5472 3410 5474
rect 3076 5471 3077 5472
rect 3071 5470 3077 5471
rect 2812 5464 2818 5466
rect 1934 5463 1940 5464
rect 1330 5462 1336 5463
rect 2816 5462 2818 5464
rect 3408 5462 3410 5472
rect 1974 5461 1980 5462
rect 2815 5461 2821 5462
rect 3407 5461 3413 5462
rect 1974 5457 1975 5461
rect 1979 5457 1980 5461
rect 1974 5456 1980 5457
rect 2022 5460 2028 5461
rect 2166 5460 2172 5461
rect 2342 5460 2348 5461
rect 2526 5460 2532 5461
rect 2718 5460 2724 5461
rect 2022 5456 2023 5460
rect 2027 5456 2028 5460
rect 2022 5455 2028 5456
rect 2114 5459 2125 5460
rect 2114 5455 2115 5459
rect 2119 5455 2120 5459
rect 2124 5455 2125 5459
rect 2166 5456 2167 5460
rect 2171 5456 2172 5460
rect 2166 5455 2172 5456
rect 2263 5459 2269 5460
rect 2263 5455 2264 5459
rect 2268 5458 2269 5459
rect 2278 5459 2284 5460
rect 2278 5458 2279 5459
rect 2268 5456 2279 5458
rect 2268 5455 2269 5456
rect 2114 5454 2125 5455
rect 2263 5454 2269 5455
rect 2278 5455 2279 5456
rect 2283 5455 2284 5459
rect 2342 5456 2343 5460
rect 2347 5456 2348 5460
rect 2342 5455 2348 5456
rect 2439 5459 2448 5460
rect 2439 5455 2440 5459
rect 2447 5455 2448 5459
rect 2526 5456 2527 5460
rect 2531 5456 2532 5460
rect 2526 5455 2532 5456
rect 2623 5459 2629 5460
rect 2623 5455 2624 5459
rect 2628 5458 2629 5459
rect 2655 5459 2661 5460
rect 2655 5458 2656 5459
rect 2628 5456 2656 5458
rect 2628 5455 2629 5456
rect 2278 5454 2284 5455
rect 2439 5454 2448 5455
rect 2623 5454 2629 5455
rect 2655 5455 2656 5456
rect 2660 5455 2661 5459
rect 2718 5456 2719 5460
rect 2723 5456 2724 5460
rect 2815 5457 2816 5461
rect 2820 5457 2821 5461
rect 2815 5456 2821 5457
rect 2910 5460 2916 5461
rect 3110 5460 3116 5461
rect 3310 5460 3316 5461
rect 2910 5456 2911 5460
rect 2915 5456 2916 5460
rect 2718 5455 2724 5456
rect 2910 5455 2916 5456
rect 3007 5459 3016 5460
rect 3007 5455 3008 5459
rect 3015 5455 3016 5459
rect 3110 5456 3111 5460
rect 3115 5456 3116 5460
rect 3110 5455 3116 5456
rect 3207 5459 3216 5460
rect 3207 5455 3208 5459
rect 3215 5455 3216 5459
rect 3310 5456 3311 5460
rect 3315 5456 3316 5460
rect 3407 5457 3408 5461
rect 3412 5457 3413 5461
rect 3407 5456 3413 5457
rect 3798 5461 3804 5462
rect 3798 5457 3799 5461
rect 3803 5457 3804 5461
rect 3798 5456 3804 5457
rect 3310 5455 3316 5456
rect 2655 5454 2661 5455
rect 3007 5454 3016 5455
rect 3207 5454 3216 5455
rect 814 5452 820 5453
rect 950 5452 956 5453
rect 1086 5452 1092 5453
rect 1222 5452 1228 5453
rect 1358 5452 1364 5453
rect 1455 5452 1461 5453
rect 110 5451 116 5452
rect 110 5447 111 5451
rect 115 5447 116 5451
rect 814 5448 815 5452
rect 819 5448 820 5452
rect 814 5447 820 5448
rect 911 5451 917 5452
rect 911 5447 912 5451
rect 916 5450 917 5451
rect 930 5451 936 5452
rect 930 5450 931 5451
rect 916 5448 931 5450
rect 916 5447 917 5448
rect 110 5446 116 5447
rect 911 5446 917 5447
rect 930 5447 931 5448
rect 935 5447 936 5451
rect 950 5448 951 5452
rect 955 5448 956 5452
rect 950 5447 956 5448
rect 1047 5451 1053 5452
rect 1047 5447 1048 5451
rect 1052 5450 1053 5451
rect 1066 5451 1072 5452
rect 1066 5450 1067 5451
rect 1052 5448 1067 5450
rect 1052 5447 1053 5448
rect 930 5446 936 5447
rect 1047 5446 1053 5447
rect 1066 5447 1067 5448
rect 1071 5447 1072 5451
rect 1086 5448 1087 5452
rect 1091 5448 1092 5452
rect 1086 5447 1092 5448
rect 1183 5451 1189 5452
rect 1183 5447 1184 5451
rect 1188 5450 1189 5451
rect 1202 5451 1208 5452
rect 1202 5450 1203 5451
rect 1188 5448 1203 5450
rect 1188 5447 1189 5448
rect 1066 5446 1072 5447
rect 1183 5446 1189 5447
rect 1202 5447 1203 5448
rect 1207 5447 1208 5451
rect 1222 5448 1223 5452
rect 1227 5448 1228 5452
rect 1222 5447 1228 5448
rect 1318 5451 1325 5452
rect 1318 5447 1319 5451
rect 1324 5447 1325 5451
rect 1358 5448 1359 5452
rect 1363 5448 1364 5452
rect 1358 5447 1364 5448
rect 1454 5451 1456 5452
rect 1454 5447 1455 5451
rect 1460 5448 1461 5452
rect 1459 5447 1461 5448
rect 1934 5451 1940 5452
rect 1934 5447 1935 5451
rect 1939 5447 1940 5451
rect 1202 5446 1208 5447
rect 1318 5446 1325 5447
rect 1454 5446 1460 5447
rect 1934 5446 1940 5447
rect 1994 5445 2000 5446
rect 1974 5444 1980 5445
rect 1974 5440 1975 5444
rect 1979 5440 1980 5444
rect 1994 5441 1995 5445
rect 1999 5441 2000 5445
rect 1994 5440 2000 5441
rect 2138 5445 2144 5446
rect 2138 5441 2139 5445
rect 2143 5441 2144 5445
rect 2138 5440 2144 5441
rect 2314 5445 2320 5446
rect 2314 5441 2315 5445
rect 2319 5441 2320 5445
rect 2314 5440 2320 5441
rect 2498 5445 2504 5446
rect 2498 5441 2499 5445
rect 2503 5441 2504 5445
rect 2498 5440 2504 5441
rect 2690 5445 2696 5446
rect 2690 5441 2691 5445
rect 2695 5441 2696 5445
rect 2690 5440 2696 5441
rect 2882 5445 2888 5446
rect 2882 5441 2883 5445
rect 2887 5441 2888 5445
rect 2882 5440 2888 5441
rect 3082 5445 3088 5446
rect 3082 5441 3083 5445
rect 3087 5441 3088 5445
rect 3082 5440 3088 5441
rect 3282 5445 3288 5446
rect 3282 5441 3283 5445
rect 3287 5441 3288 5445
rect 3282 5440 3288 5441
rect 3798 5444 3804 5445
rect 3798 5440 3799 5444
rect 3803 5440 3804 5444
rect 1974 5439 1980 5440
rect 3798 5439 3804 5440
rect 4558 5435 4564 5436
rect 4373 5432 4461 5434
rect 4459 5426 4461 5432
rect 4558 5431 4559 5435
rect 4563 5431 4564 5435
rect 4818 5435 4824 5436
rect 4558 5430 4564 5431
rect 4602 5427 4608 5428
rect 4602 5426 4603 5427
rect 4459 5424 4603 5426
rect 4602 5423 4603 5424
rect 4607 5423 4608 5427
rect 4788 5426 4790 5433
rect 4818 5431 4819 5435
rect 4823 5434 4824 5435
rect 5314 5435 5320 5436
rect 5314 5434 5315 5435
rect 4823 5432 4905 5434
rect 5205 5432 5315 5434
rect 4823 5431 4824 5432
rect 4818 5430 4824 5431
rect 5314 5431 5315 5432
rect 5319 5431 5320 5435
rect 5314 5430 5320 5431
rect 5230 5427 5236 5428
rect 5230 5426 5231 5427
rect 4788 5424 5231 5426
rect 4602 5422 4608 5423
rect 5230 5423 5231 5424
rect 5235 5423 5236 5427
rect 5230 5422 5236 5423
rect 1250 5419 1256 5420
rect 1250 5415 1251 5419
rect 1255 5418 1256 5419
rect 1454 5419 1460 5420
rect 1454 5418 1455 5419
rect 1255 5416 1455 5418
rect 1255 5415 1256 5416
rect 1250 5414 1256 5415
rect 1454 5415 1455 5416
rect 1459 5415 1460 5419
rect 1454 5414 1460 5415
rect 2135 5403 2141 5404
rect 2135 5402 2136 5403
rect 2092 5400 2136 5402
rect 2092 5393 2094 5400
rect 2135 5399 2136 5400
rect 2140 5399 2141 5403
rect 2135 5398 2141 5399
rect 2122 5395 2128 5396
rect 2122 5391 2123 5395
rect 2127 5394 2128 5395
rect 2278 5395 2284 5396
rect 2127 5392 2145 5394
rect 2127 5391 2128 5392
rect 2122 5390 2128 5391
rect 2278 5391 2279 5395
rect 2283 5394 2284 5395
rect 2558 5395 2564 5396
rect 2283 5392 2321 5394
rect 2283 5391 2284 5392
rect 2278 5390 2284 5391
rect 2558 5391 2559 5395
rect 2563 5391 2564 5395
rect 2558 5390 2564 5391
rect 2655 5395 2661 5396
rect 2655 5391 2656 5395
rect 2660 5394 2661 5395
rect 2978 5395 2984 5396
rect 2660 5392 2697 5394
rect 2660 5391 2661 5392
rect 2655 5390 2661 5391
rect 2978 5391 2979 5395
rect 2983 5391 2984 5395
rect 2978 5390 2984 5391
rect 3010 5395 3016 5396
rect 3010 5391 3011 5395
rect 3015 5394 3016 5395
rect 3210 5395 3216 5396
rect 3015 5392 3089 5394
rect 3015 5391 3016 5392
rect 3010 5390 3016 5391
rect 3210 5391 3211 5395
rect 3215 5394 3216 5395
rect 3215 5392 3289 5394
rect 3215 5391 3216 5392
rect 3210 5390 3216 5391
rect 4722 5383 4728 5384
rect 4722 5382 4723 5383
rect 4596 5380 4723 5382
rect 3786 5379 3792 5380
rect 3786 5375 3787 5379
rect 3791 5378 3792 5379
rect 4596 5378 4598 5380
rect 4722 5379 4723 5380
rect 4727 5379 4728 5383
rect 4722 5378 4728 5379
rect 4930 5379 4936 5380
rect 4930 5378 4931 5379
rect 3791 5376 3865 5378
rect 4533 5376 4598 5378
rect 4877 5376 4931 5378
rect 3791 5375 3792 5376
rect 3786 5374 3792 5375
rect 4002 5375 4008 5376
rect 110 5373 116 5374
rect 1934 5373 1940 5374
rect 110 5369 111 5373
rect 115 5369 116 5373
rect 110 5368 116 5369
rect 902 5372 908 5373
rect 1038 5372 1044 5373
rect 1182 5372 1188 5373
rect 1334 5372 1340 5373
rect 1494 5372 1500 5373
rect 1662 5372 1668 5373
rect 1814 5372 1820 5373
rect 902 5368 903 5372
rect 907 5368 908 5372
rect 902 5367 908 5368
rect 999 5371 1008 5372
rect 999 5367 1000 5371
rect 1007 5367 1008 5371
rect 1038 5368 1039 5372
rect 1043 5368 1044 5372
rect 1038 5367 1044 5368
rect 1134 5371 1141 5372
rect 1134 5367 1135 5371
rect 1140 5367 1141 5371
rect 1182 5368 1183 5372
rect 1187 5368 1188 5372
rect 1182 5367 1188 5368
rect 1274 5371 1285 5372
rect 1274 5367 1275 5371
rect 1279 5367 1280 5371
rect 1284 5367 1285 5371
rect 1334 5368 1335 5372
rect 1339 5368 1340 5372
rect 1334 5367 1340 5368
rect 1426 5371 1437 5372
rect 1426 5367 1427 5371
rect 1431 5367 1432 5371
rect 1436 5367 1437 5371
rect 1494 5368 1495 5372
rect 1499 5368 1500 5372
rect 1494 5367 1500 5368
rect 1591 5371 1600 5372
rect 1591 5367 1592 5371
rect 1599 5367 1600 5371
rect 1662 5368 1663 5372
rect 1667 5368 1668 5372
rect 1662 5367 1668 5368
rect 1758 5371 1765 5372
rect 1758 5367 1759 5371
rect 1764 5367 1765 5371
rect 1814 5368 1815 5372
rect 1819 5368 1820 5372
rect 1814 5367 1820 5368
rect 1906 5371 1917 5372
rect 1906 5367 1907 5371
rect 1911 5367 1912 5371
rect 1916 5367 1917 5371
rect 1934 5369 1935 5373
rect 1939 5369 1940 5373
rect 4002 5371 4003 5375
rect 4007 5371 4008 5375
rect 4002 5370 4008 5371
rect 4138 5375 4144 5376
rect 4138 5371 4139 5375
rect 4143 5371 4144 5375
rect 4138 5370 4144 5371
rect 4282 5375 4288 5376
rect 4282 5371 4283 5375
rect 4287 5371 4288 5375
rect 4282 5370 4288 5371
rect 4698 5375 4704 5376
rect 4698 5371 4699 5375
rect 4703 5371 4704 5375
rect 4930 5375 4931 5376
rect 4935 5375 4936 5379
rect 4930 5374 4936 5375
rect 5022 5379 5028 5380
rect 5022 5375 5023 5379
rect 5027 5375 5028 5379
rect 5022 5374 5028 5375
rect 4698 5370 4704 5371
rect 1934 5368 1940 5369
rect 999 5366 1008 5367
rect 1134 5366 1141 5367
rect 1274 5366 1285 5367
rect 1426 5366 1437 5367
rect 1591 5366 1600 5367
rect 1758 5366 1765 5367
rect 1906 5366 1917 5367
rect 874 5357 880 5358
rect 110 5356 116 5357
rect 110 5352 111 5356
rect 115 5352 116 5356
rect 874 5353 875 5357
rect 879 5353 880 5357
rect 874 5352 880 5353
rect 1010 5357 1016 5358
rect 1010 5353 1011 5357
rect 1015 5353 1016 5357
rect 1010 5352 1016 5353
rect 1154 5357 1160 5358
rect 1154 5353 1155 5357
rect 1159 5353 1160 5357
rect 1154 5352 1160 5353
rect 1306 5357 1312 5358
rect 1306 5353 1307 5357
rect 1311 5353 1312 5357
rect 1306 5352 1312 5353
rect 1466 5357 1472 5358
rect 1466 5353 1467 5357
rect 1471 5353 1472 5357
rect 1466 5352 1472 5353
rect 1634 5357 1640 5358
rect 1634 5353 1635 5357
rect 1639 5353 1640 5357
rect 1634 5352 1640 5353
rect 1786 5357 1792 5358
rect 1786 5353 1787 5357
rect 1791 5353 1792 5357
rect 1786 5352 1792 5353
rect 1934 5356 1940 5357
rect 1934 5352 1935 5356
rect 1939 5352 1940 5356
rect 110 5351 116 5352
rect 1934 5351 1940 5352
rect 3758 5343 3764 5344
rect 3758 5342 3759 5343
rect 3619 5340 3759 5342
rect 2442 5339 2448 5340
rect 2146 5335 2152 5336
rect 2146 5331 2147 5335
rect 2151 5331 2152 5335
rect 2442 5335 2443 5339
rect 2447 5338 2448 5339
rect 3619 5338 3621 5340
rect 3758 5339 3759 5340
rect 3763 5339 3764 5343
rect 3758 5338 3764 5339
rect 2447 5336 2465 5338
rect 3365 5336 3621 5338
rect 2447 5335 2448 5336
rect 2442 5334 2448 5335
rect 2866 5335 2872 5336
rect 2146 5330 2152 5331
rect 2866 5331 2867 5335
rect 2871 5331 2872 5335
rect 2866 5330 2872 5331
rect 3658 5335 3664 5336
rect 3658 5331 3659 5335
rect 3663 5331 3664 5335
rect 3658 5330 3664 5331
rect 3838 5328 3844 5329
rect 5662 5328 5668 5329
rect 3838 5324 3839 5328
rect 3843 5324 3844 5328
rect 3838 5323 3844 5324
rect 3858 5327 3864 5328
rect 3858 5323 3859 5327
rect 3863 5323 3864 5327
rect 3858 5322 3864 5323
rect 3994 5327 4000 5328
rect 3994 5323 3995 5327
rect 3999 5323 4000 5327
rect 3994 5322 4000 5323
rect 4130 5327 4136 5328
rect 4130 5323 4131 5327
rect 4135 5323 4136 5327
rect 4130 5322 4136 5323
rect 4274 5327 4280 5328
rect 4274 5323 4275 5327
rect 4279 5323 4280 5327
rect 4274 5322 4280 5323
rect 4434 5327 4440 5328
rect 4434 5323 4435 5327
rect 4439 5323 4440 5327
rect 4434 5322 4440 5323
rect 4602 5327 4608 5328
rect 4602 5323 4603 5327
rect 4607 5323 4608 5327
rect 4602 5322 4608 5323
rect 4778 5327 4784 5328
rect 4778 5323 4779 5327
rect 4783 5323 4784 5327
rect 4778 5322 4784 5323
rect 4962 5327 4968 5328
rect 4962 5323 4963 5327
rect 4967 5323 4968 5327
rect 5662 5324 5663 5328
rect 5667 5324 5668 5328
rect 5662 5323 5668 5324
rect 4962 5322 4968 5323
rect 4930 5319 4936 5320
rect 2146 5315 2152 5316
rect 2146 5311 2147 5315
rect 2151 5314 2152 5315
rect 2582 5315 2588 5316
rect 2582 5314 2583 5315
rect 2151 5312 2583 5314
rect 2151 5311 2152 5312
rect 2146 5310 2152 5311
rect 2582 5311 2583 5312
rect 2587 5311 2588 5315
rect 4930 5315 4931 5319
rect 4935 5318 4936 5319
rect 4935 5316 5090 5318
rect 4935 5315 4936 5316
rect 4930 5314 4936 5315
rect 5088 5314 5090 5316
rect 5087 5313 5093 5314
rect 3886 5312 3892 5313
rect 4022 5312 4028 5313
rect 4158 5312 4164 5313
rect 4302 5312 4308 5313
rect 4462 5312 4468 5313
rect 4630 5312 4636 5313
rect 4806 5312 4812 5313
rect 4990 5312 4996 5313
rect 2582 5310 2588 5311
rect 3838 5311 3844 5312
rect 1002 5307 1008 5308
rect 972 5298 974 5305
rect 1002 5303 1003 5307
rect 1007 5306 1008 5307
rect 1250 5307 1256 5308
rect 1007 5304 1017 5306
rect 1007 5303 1008 5304
rect 1002 5302 1008 5303
rect 1250 5303 1251 5307
rect 1255 5303 1256 5307
rect 1550 5307 1556 5308
rect 1250 5302 1256 5303
rect 1274 5299 1280 5300
rect 1274 5298 1275 5299
rect 972 5296 1275 5298
rect 1274 5295 1275 5296
rect 1279 5295 1280 5299
rect 1404 5298 1406 5305
rect 1550 5303 1551 5307
rect 1555 5303 1556 5307
rect 1550 5302 1556 5303
rect 1594 5307 1600 5308
rect 1594 5303 1595 5307
rect 1599 5306 1600 5307
rect 2114 5307 2120 5308
rect 2114 5306 2115 5307
rect 1599 5304 1641 5306
rect 1885 5304 2115 5306
rect 1599 5303 1600 5304
rect 1594 5302 1600 5303
rect 2114 5303 2115 5304
rect 2119 5303 2120 5307
rect 3838 5307 3839 5311
rect 3843 5307 3844 5311
rect 3886 5308 3887 5312
rect 3891 5308 3892 5312
rect 3886 5307 3892 5308
rect 3983 5311 3989 5312
rect 3983 5307 3984 5311
rect 3988 5310 3989 5311
rect 4002 5311 4008 5312
rect 4002 5310 4003 5311
rect 3988 5308 4003 5310
rect 3988 5307 3989 5308
rect 3838 5306 3844 5307
rect 3983 5306 3989 5307
rect 4002 5307 4003 5308
rect 4007 5307 4008 5311
rect 4022 5308 4023 5312
rect 4027 5308 4028 5312
rect 4022 5307 4028 5308
rect 4119 5311 4125 5312
rect 4119 5307 4120 5311
rect 4124 5310 4125 5311
rect 4138 5311 4144 5312
rect 4138 5310 4139 5311
rect 4124 5308 4139 5310
rect 4124 5307 4125 5308
rect 4002 5306 4008 5307
rect 4119 5306 4125 5307
rect 4138 5307 4139 5308
rect 4143 5307 4144 5311
rect 4158 5308 4159 5312
rect 4163 5308 4164 5312
rect 4158 5307 4164 5308
rect 4255 5311 4261 5312
rect 4255 5307 4256 5311
rect 4260 5310 4261 5311
rect 4282 5311 4288 5312
rect 4282 5310 4283 5311
rect 4260 5308 4283 5310
rect 4260 5307 4261 5308
rect 4138 5306 4144 5307
rect 4255 5306 4261 5307
rect 4282 5307 4283 5308
rect 4287 5307 4288 5311
rect 4302 5308 4303 5312
rect 4307 5308 4308 5312
rect 4302 5307 4308 5308
rect 4394 5311 4405 5312
rect 4394 5307 4395 5311
rect 4399 5307 4400 5311
rect 4404 5307 4405 5311
rect 4462 5308 4463 5312
rect 4467 5308 4468 5312
rect 4462 5307 4468 5308
rect 4558 5311 4565 5312
rect 4558 5307 4559 5311
rect 4564 5307 4565 5311
rect 4630 5308 4631 5312
rect 4635 5308 4636 5312
rect 4630 5307 4636 5308
rect 4722 5311 4733 5312
rect 4722 5307 4723 5311
rect 4727 5307 4728 5311
rect 4732 5307 4733 5311
rect 4806 5308 4807 5312
rect 4811 5308 4812 5312
rect 4806 5307 4812 5308
rect 4898 5311 4909 5312
rect 4898 5307 4899 5311
rect 4903 5307 4904 5311
rect 4908 5307 4909 5311
rect 4990 5308 4991 5312
rect 4995 5308 4996 5312
rect 5087 5309 5088 5313
rect 5092 5309 5093 5313
rect 5087 5308 5093 5309
rect 5662 5311 5668 5312
rect 4990 5307 4996 5308
rect 5662 5307 5663 5311
rect 5667 5307 5668 5311
rect 4282 5306 4288 5307
rect 4394 5306 4405 5307
rect 4558 5306 4565 5307
rect 4722 5306 4733 5307
rect 4898 5306 4909 5307
rect 5662 5306 5668 5307
rect 2114 5302 2120 5303
rect 1758 5299 1764 5300
rect 1758 5298 1759 5299
rect 1404 5296 1759 5298
rect 1274 5294 1280 5295
rect 1758 5295 1759 5296
rect 1763 5295 1764 5299
rect 1758 5294 1764 5295
rect 1974 5288 1980 5289
rect 3798 5288 3804 5289
rect 1974 5284 1975 5288
rect 1979 5284 1980 5288
rect 1974 5283 1980 5284
rect 2050 5287 2056 5288
rect 2050 5283 2051 5287
rect 2055 5283 2056 5287
rect 2050 5282 2056 5283
rect 2458 5287 2464 5288
rect 2458 5283 2459 5287
rect 2463 5283 2464 5287
rect 2458 5282 2464 5283
rect 2858 5287 2864 5288
rect 2858 5283 2859 5287
rect 2863 5283 2864 5287
rect 2858 5282 2864 5283
rect 3266 5287 3272 5288
rect 3266 5283 3267 5287
rect 3271 5283 3272 5287
rect 3266 5282 3272 5283
rect 3650 5287 3656 5288
rect 3650 5283 3651 5287
rect 3655 5283 3656 5287
rect 3798 5284 3799 5288
rect 3803 5284 3804 5288
rect 3798 5283 3804 5284
rect 3650 5282 3656 5283
rect 4066 5279 4072 5280
rect 862 5275 868 5276
rect 862 5274 863 5275
rect 736 5272 863 5274
rect 736 5270 738 5272
rect 862 5271 863 5272
rect 867 5271 868 5275
rect 4066 5275 4067 5279
rect 4071 5278 4072 5279
rect 4390 5279 4396 5280
rect 4390 5278 4391 5279
rect 4071 5276 4391 5278
rect 4071 5275 4072 5276
rect 4066 5274 4072 5275
rect 4390 5275 4391 5276
rect 4395 5275 4396 5279
rect 4390 5274 4396 5275
rect 2078 5272 2084 5273
rect 2486 5272 2492 5273
rect 2886 5272 2892 5273
rect 3294 5272 3300 5273
rect 3678 5272 3684 5273
rect 862 5270 868 5271
rect 1134 5271 1140 5272
rect 685 5268 738 5270
rect 994 5267 1000 5268
rect 832 5262 834 5265
rect 879 5263 885 5264
rect 879 5262 880 5263
rect 832 5260 880 5262
rect 879 5259 880 5260
rect 884 5259 885 5263
rect 994 5263 995 5267
rect 999 5263 1000 5267
rect 1134 5267 1135 5271
rect 1139 5267 1140 5271
rect 1542 5271 1548 5272
rect 1542 5270 1543 5271
rect 1525 5268 1543 5270
rect 1134 5266 1140 5267
rect 1250 5267 1256 5268
rect 994 5262 1000 5263
rect 1250 5263 1251 5267
rect 1255 5263 1256 5267
rect 1542 5267 1543 5268
rect 1547 5267 1548 5271
rect 1778 5271 1784 5272
rect 1778 5270 1779 5271
rect 1717 5268 1779 5270
rect 1542 5266 1548 5267
rect 1778 5267 1779 5268
rect 1783 5267 1784 5271
rect 1906 5271 1912 5272
rect 1906 5270 1907 5271
rect 1885 5268 1907 5270
rect 1778 5266 1784 5267
rect 1906 5267 1907 5268
rect 1911 5267 1912 5271
rect 1906 5266 1912 5267
rect 1974 5271 1980 5272
rect 1974 5267 1975 5271
rect 1979 5267 1980 5271
rect 2078 5268 2079 5272
rect 2083 5268 2084 5272
rect 2078 5267 2084 5268
rect 2175 5271 2181 5272
rect 2175 5267 2176 5271
rect 2180 5270 2181 5271
rect 2198 5271 2204 5272
rect 2198 5270 2199 5271
rect 2180 5268 2199 5270
rect 2180 5267 2181 5268
rect 1974 5266 1980 5267
rect 2175 5266 2181 5267
rect 2198 5267 2199 5268
rect 2203 5267 2204 5271
rect 2486 5268 2487 5272
rect 2491 5268 2492 5272
rect 2486 5267 2492 5268
rect 2582 5271 2589 5272
rect 2582 5267 2583 5271
rect 2588 5267 2589 5271
rect 2886 5268 2887 5272
rect 2891 5268 2892 5272
rect 2886 5267 2892 5268
rect 2978 5271 2989 5272
rect 2978 5267 2979 5271
rect 2983 5267 2984 5271
rect 2988 5267 2989 5271
rect 3294 5268 3295 5272
rect 3299 5268 3300 5272
rect 3294 5267 3300 5268
rect 3391 5271 3397 5272
rect 3391 5267 3392 5271
rect 3396 5270 3397 5271
rect 3658 5271 3664 5272
rect 3658 5270 3659 5271
rect 3396 5268 3659 5270
rect 3396 5267 3397 5268
rect 2198 5266 2204 5267
rect 2582 5266 2589 5267
rect 2978 5266 2989 5267
rect 3391 5266 3397 5267
rect 3658 5267 3659 5268
rect 3663 5267 3664 5271
rect 3678 5268 3679 5272
rect 3683 5268 3684 5272
rect 3678 5267 3684 5268
rect 3775 5271 3781 5272
rect 3775 5267 3776 5271
rect 3780 5270 3781 5271
rect 3786 5271 3792 5272
rect 3786 5270 3787 5271
rect 3780 5268 3787 5270
rect 3780 5267 3781 5268
rect 3658 5266 3664 5267
rect 3775 5266 3781 5267
rect 3786 5267 3787 5268
rect 3791 5267 3792 5271
rect 3786 5266 3792 5267
rect 3798 5271 3804 5272
rect 3798 5267 3799 5271
rect 3803 5267 3804 5271
rect 3798 5266 3804 5267
rect 1250 5262 1256 5263
rect 879 5258 885 5259
rect 3838 5249 3844 5250
rect 5662 5249 5668 5250
rect 3838 5245 3839 5249
rect 3843 5245 3844 5249
rect 3838 5244 3844 5245
rect 3998 5248 4004 5249
rect 4198 5248 4204 5249
rect 4398 5248 4404 5249
rect 4606 5248 4612 5249
rect 4822 5248 4828 5249
rect 5038 5248 5044 5249
rect 3998 5244 3999 5248
rect 4003 5244 4004 5248
rect 3998 5243 4004 5244
rect 4095 5247 4104 5248
rect 4095 5243 4096 5247
rect 4103 5243 4104 5247
rect 4198 5244 4199 5248
rect 4203 5244 4204 5248
rect 4198 5243 4204 5244
rect 4295 5247 4304 5248
rect 4295 5243 4296 5247
rect 4303 5243 4304 5247
rect 4398 5244 4399 5248
rect 4403 5244 4404 5248
rect 4398 5243 4404 5244
rect 4490 5247 4501 5248
rect 4490 5243 4491 5247
rect 4495 5243 4496 5247
rect 4500 5243 4501 5247
rect 4606 5244 4607 5248
rect 4611 5244 4612 5248
rect 4606 5243 4612 5244
rect 4698 5247 4709 5248
rect 4698 5243 4699 5247
rect 4703 5243 4704 5247
rect 4708 5243 4709 5247
rect 4822 5244 4823 5248
rect 4827 5244 4828 5248
rect 4822 5243 4828 5244
rect 4919 5247 4928 5248
rect 4919 5243 4920 5247
rect 4927 5243 4928 5247
rect 5038 5244 5039 5248
rect 5043 5244 5044 5248
rect 5038 5243 5044 5244
rect 5134 5247 5141 5248
rect 5134 5243 5135 5247
rect 5140 5243 5141 5247
rect 5662 5245 5663 5249
rect 5667 5245 5668 5249
rect 5662 5244 5668 5245
rect 4095 5242 4104 5243
rect 4295 5242 4304 5243
rect 4490 5242 4501 5243
rect 4698 5242 4709 5243
rect 4919 5242 4928 5243
rect 5134 5242 5141 5243
rect 994 5239 1000 5240
rect 994 5235 995 5239
rect 999 5238 1000 5239
rect 1366 5239 1372 5240
rect 1366 5238 1367 5239
rect 999 5236 1367 5238
rect 999 5235 1000 5236
rect 994 5234 1000 5235
rect 1366 5235 1367 5236
rect 1371 5235 1372 5239
rect 1366 5234 1372 5235
rect 3970 5233 3976 5234
rect 3838 5232 3844 5233
rect 3838 5228 3839 5232
rect 3843 5228 3844 5232
rect 3970 5229 3971 5233
rect 3975 5229 3976 5233
rect 3970 5228 3976 5229
rect 4170 5233 4176 5234
rect 4170 5229 4171 5233
rect 4175 5229 4176 5233
rect 4170 5228 4176 5229
rect 4370 5233 4376 5234
rect 4370 5229 4371 5233
rect 4375 5229 4376 5233
rect 4370 5228 4376 5229
rect 4578 5233 4584 5234
rect 4578 5229 4579 5233
rect 4583 5229 4584 5233
rect 4578 5228 4584 5229
rect 4794 5233 4800 5234
rect 4794 5229 4795 5233
rect 4799 5229 4800 5233
rect 4794 5228 4800 5229
rect 5010 5233 5016 5234
rect 5010 5229 5011 5233
rect 5015 5229 5016 5233
rect 5010 5228 5016 5229
rect 5662 5232 5668 5233
rect 5662 5228 5663 5232
rect 5667 5228 5668 5232
rect 3838 5227 3844 5228
rect 5662 5227 5668 5228
rect 110 5220 116 5221
rect 1934 5220 1940 5221
rect 110 5216 111 5220
rect 115 5216 116 5220
rect 110 5215 116 5216
rect 586 5219 592 5220
rect 586 5215 587 5219
rect 591 5215 592 5219
rect 586 5214 592 5215
rect 738 5219 744 5220
rect 738 5215 739 5219
rect 743 5215 744 5219
rect 738 5214 744 5215
rect 898 5219 904 5220
rect 898 5215 899 5219
rect 903 5215 904 5219
rect 898 5214 904 5215
rect 1066 5219 1072 5220
rect 1066 5215 1067 5219
rect 1071 5215 1072 5219
rect 1066 5214 1072 5215
rect 1242 5219 1248 5220
rect 1242 5215 1243 5219
rect 1247 5215 1248 5219
rect 1242 5214 1248 5215
rect 1426 5219 1432 5220
rect 1426 5215 1427 5219
rect 1431 5215 1432 5219
rect 1426 5214 1432 5215
rect 1618 5219 1624 5220
rect 1618 5215 1619 5219
rect 1623 5215 1624 5219
rect 1618 5214 1624 5215
rect 1786 5219 1792 5220
rect 1786 5215 1787 5219
rect 1791 5215 1792 5219
rect 1934 5216 1935 5220
rect 1939 5216 1940 5220
rect 1934 5215 1940 5216
rect 1786 5214 1792 5215
rect 1974 5213 1980 5214
rect 3798 5213 3804 5214
rect 879 5211 885 5212
rect 879 5207 880 5211
rect 884 5210 885 5211
rect 1778 5211 1784 5212
rect 884 5208 1026 5210
rect 884 5207 885 5208
rect 879 5206 885 5207
rect 614 5204 620 5205
rect 766 5204 772 5205
rect 926 5204 932 5205
rect 1024 5204 1026 5208
rect 1778 5207 1779 5211
rect 1783 5210 1784 5211
rect 1783 5208 1914 5210
rect 1974 5209 1975 5213
rect 1979 5209 1980 5213
rect 1974 5208 1980 5209
rect 2238 5212 2244 5213
rect 2590 5212 2596 5213
rect 2942 5212 2948 5213
rect 3302 5212 3308 5213
rect 3662 5212 3668 5213
rect 2238 5208 2239 5212
rect 2243 5208 2244 5212
rect 1783 5207 1784 5208
rect 1778 5206 1784 5207
rect 1094 5204 1100 5205
rect 1270 5204 1276 5205
rect 1454 5204 1460 5205
rect 1646 5204 1652 5205
rect 1814 5204 1820 5205
rect 1912 5204 1914 5208
rect 2238 5207 2244 5208
rect 2334 5211 2341 5212
rect 2334 5207 2335 5211
rect 2340 5207 2341 5211
rect 2590 5208 2591 5212
rect 2595 5208 2596 5212
rect 2590 5207 2596 5208
rect 2687 5211 2693 5212
rect 2687 5207 2688 5211
rect 2692 5210 2693 5211
rect 2866 5211 2872 5212
rect 2866 5210 2867 5211
rect 2692 5208 2867 5210
rect 2692 5207 2693 5208
rect 2334 5206 2341 5207
rect 2687 5206 2693 5207
rect 2866 5207 2867 5208
rect 2871 5207 2872 5211
rect 2942 5208 2943 5212
rect 2947 5208 2948 5212
rect 2942 5207 2948 5208
rect 3038 5211 3045 5212
rect 3038 5207 3039 5211
rect 3044 5207 3045 5211
rect 3302 5208 3303 5212
rect 3307 5208 3308 5212
rect 3302 5207 3308 5208
rect 3399 5211 3405 5212
rect 3399 5207 3400 5211
rect 3404 5210 3405 5211
rect 3594 5211 3600 5212
rect 3594 5210 3595 5211
rect 3404 5208 3595 5210
rect 3404 5207 3405 5208
rect 2866 5206 2872 5207
rect 3038 5206 3045 5207
rect 3399 5206 3405 5207
rect 3594 5207 3595 5208
rect 3599 5207 3600 5211
rect 3662 5208 3663 5212
rect 3667 5208 3668 5212
rect 3662 5207 3668 5208
rect 3758 5211 3765 5212
rect 3758 5207 3759 5211
rect 3764 5207 3765 5211
rect 3798 5209 3799 5213
rect 3803 5209 3804 5213
rect 3798 5208 3804 5209
rect 3594 5206 3600 5207
rect 3758 5206 3765 5207
rect 110 5203 116 5204
rect 110 5199 111 5203
rect 115 5199 116 5203
rect 614 5200 615 5204
rect 619 5200 620 5204
rect 614 5199 620 5200
rect 710 5203 717 5204
rect 710 5199 711 5203
rect 716 5199 717 5203
rect 766 5200 767 5204
rect 771 5200 772 5204
rect 766 5199 772 5200
rect 862 5203 869 5204
rect 862 5199 863 5203
rect 868 5199 869 5203
rect 926 5200 927 5204
rect 931 5200 932 5204
rect 926 5199 932 5200
rect 1023 5203 1029 5204
rect 1023 5199 1024 5203
rect 1028 5199 1029 5203
rect 1094 5200 1095 5204
rect 1099 5200 1100 5204
rect 1094 5199 1100 5200
rect 1191 5203 1197 5204
rect 1191 5199 1192 5203
rect 1196 5202 1197 5203
rect 1250 5203 1256 5204
rect 1250 5202 1251 5203
rect 1196 5200 1251 5202
rect 1196 5199 1197 5200
rect 110 5198 116 5199
rect 710 5198 717 5199
rect 862 5198 869 5199
rect 1023 5198 1029 5199
rect 1191 5198 1197 5199
rect 1250 5199 1251 5200
rect 1255 5199 1256 5203
rect 1270 5200 1271 5204
rect 1275 5200 1276 5204
rect 1270 5199 1276 5200
rect 1366 5203 1373 5204
rect 1366 5199 1367 5203
rect 1372 5199 1373 5203
rect 1454 5200 1455 5204
rect 1459 5200 1460 5204
rect 1454 5199 1460 5200
rect 1550 5203 1557 5204
rect 1550 5199 1551 5203
rect 1556 5199 1557 5203
rect 1646 5200 1647 5204
rect 1651 5200 1652 5204
rect 1646 5199 1652 5200
rect 1743 5203 1752 5204
rect 1743 5199 1744 5203
rect 1751 5199 1752 5203
rect 1814 5200 1815 5204
rect 1819 5200 1820 5204
rect 1814 5199 1820 5200
rect 1911 5203 1917 5204
rect 1911 5199 1912 5203
rect 1916 5199 1917 5203
rect 1250 5198 1256 5199
rect 1366 5198 1373 5199
rect 1550 5198 1557 5199
rect 1743 5198 1752 5199
rect 1911 5198 1917 5199
rect 1934 5203 1940 5204
rect 1934 5199 1935 5203
rect 1939 5199 1940 5203
rect 1934 5198 1940 5199
rect 2210 5197 2216 5198
rect 1974 5196 1980 5197
rect 1974 5192 1975 5196
rect 1979 5192 1980 5196
rect 2210 5193 2211 5197
rect 2215 5193 2216 5197
rect 2210 5192 2216 5193
rect 2562 5197 2568 5198
rect 2562 5193 2563 5197
rect 2567 5193 2568 5197
rect 2562 5192 2568 5193
rect 2914 5197 2920 5198
rect 2914 5193 2915 5197
rect 2919 5193 2920 5197
rect 2914 5192 2920 5193
rect 3274 5197 3280 5198
rect 3274 5193 3275 5197
rect 3279 5193 3280 5197
rect 3274 5192 3280 5193
rect 3634 5197 3640 5198
rect 3634 5193 3635 5197
rect 3639 5193 3640 5197
rect 3634 5192 3640 5193
rect 3798 5196 3804 5197
rect 3798 5192 3799 5196
rect 3803 5192 3804 5196
rect 1974 5191 1980 5192
rect 3798 5191 3804 5192
rect 4066 5183 4072 5184
rect 4066 5179 4067 5183
rect 4071 5179 4072 5183
rect 4066 5178 4072 5179
rect 4098 5183 4104 5184
rect 4098 5179 4099 5183
rect 4103 5182 4104 5183
rect 4298 5183 4304 5184
rect 4103 5180 4177 5182
rect 4103 5179 4104 5180
rect 4098 5178 4104 5179
rect 4298 5179 4299 5183
rect 4303 5182 4304 5183
rect 4714 5183 4720 5184
rect 4714 5182 4715 5183
rect 4303 5180 4377 5182
rect 4677 5180 4715 5182
rect 4303 5179 4304 5180
rect 4298 5178 4304 5179
rect 4714 5179 4715 5180
rect 4719 5179 4720 5183
rect 4898 5183 4904 5184
rect 4898 5182 4899 5183
rect 4893 5180 4899 5182
rect 4714 5178 4720 5179
rect 4898 5179 4899 5180
rect 4903 5179 4904 5183
rect 4898 5178 4904 5179
rect 4922 5183 4928 5184
rect 4922 5179 4923 5183
rect 4927 5182 4928 5183
rect 4927 5180 5017 5182
rect 4927 5179 4928 5180
rect 4922 5178 4928 5179
rect 2198 5147 2204 5148
rect 2198 5143 2199 5147
rect 2203 5146 2204 5147
rect 2638 5147 2644 5148
rect 2203 5144 2217 5146
rect 2203 5143 2204 5144
rect 2198 5142 2204 5143
rect 2638 5143 2639 5147
rect 2643 5143 2644 5147
rect 3038 5147 3044 5148
rect 3013 5144 3022 5146
rect 2638 5142 2644 5143
rect 3020 5138 3022 5144
rect 3038 5143 3039 5147
rect 3043 5146 3044 5147
rect 3594 5147 3600 5148
rect 3043 5144 3281 5146
rect 3043 5143 3044 5144
rect 3038 5142 3044 5143
rect 3594 5143 3595 5147
rect 3599 5146 3600 5147
rect 3599 5144 3641 5146
rect 3599 5143 3600 5144
rect 3594 5142 3600 5143
rect 3114 5139 3120 5140
rect 3114 5138 3115 5139
rect 3020 5136 3115 5138
rect 3114 5135 3115 5136
rect 3119 5135 3120 5139
rect 3114 5134 3120 5135
rect 110 5133 116 5134
rect 1934 5133 1940 5134
rect 110 5129 111 5133
rect 115 5129 116 5133
rect 110 5128 116 5129
rect 366 5132 372 5133
rect 534 5132 540 5133
rect 710 5132 716 5133
rect 894 5132 900 5133
rect 1078 5132 1084 5133
rect 1262 5132 1268 5133
rect 1446 5132 1452 5133
rect 1630 5132 1636 5133
rect 1814 5132 1820 5133
rect 366 5128 367 5132
rect 371 5128 372 5132
rect 366 5127 372 5128
rect 463 5131 472 5132
rect 463 5127 464 5131
rect 471 5127 472 5131
rect 534 5128 535 5132
rect 539 5128 540 5132
rect 534 5127 540 5128
rect 630 5131 637 5132
rect 630 5127 631 5131
rect 636 5127 637 5131
rect 710 5128 711 5132
rect 715 5128 716 5132
rect 710 5127 716 5128
rect 807 5131 813 5132
rect 807 5127 808 5131
rect 812 5130 813 5131
rect 831 5131 837 5132
rect 831 5130 832 5131
rect 812 5128 832 5130
rect 812 5127 813 5128
rect 463 5126 472 5127
rect 630 5126 637 5127
rect 807 5126 813 5127
rect 831 5127 832 5128
rect 836 5127 837 5131
rect 894 5128 895 5132
rect 899 5128 900 5132
rect 894 5127 900 5128
rect 991 5131 997 5132
rect 991 5127 992 5131
rect 996 5130 997 5131
rect 1014 5131 1020 5132
rect 1014 5130 1015 5131
rect 996 5128 1015 5130
rect 996 5127 997 5128
rect 831 5126 837 5127
rect 991 5126 997 5127
rect 1014 5127 1015 5128
rect 1019 5127 1020 5131
rect 1078 5128 1079 5132
rect 1083 5128 1084 5132
rect 1078 5127 1084 5128
rect 1170 5131 1181 5132
rect 1170 5127 1171 5131
rect 1175 5127 1176 5131
rect 1180 5127 1181 5131
rect 1262 5128 1263 5132
rect 1267 5128 1268 5132
rect 1262 5127 1268 5128
rect 1359 5131 1365 5132
rect 1359 5127 1360 5131
rect 1364 5130 1365 5131
rect 1383 5131 1389 5132
rect 1383 5130 1384 5131
rect 1364 5128 1384 5130
rect 1364 5127 1365 5128
rect 1014 5126 1020 5127
rect 1170 5126 1181 5127
rect 1359 5126 1365 5127
rect 1383 5127 1384 5128
rect 1388 5127 1389 5131
rect 1446 5128 1447 5132
rect 1451 5128 1452 5132
rect 1446 5127 1452 5128
rect 1542 5131 1549 5132
rect 1542 5127 1543 5131
rect 1548 5127 1549 5131
rect 1630 5128 1631 5132
rect 1635 5128 1636 5132
rect 1630 5127 1636 5128
rect 1726 5131 1733 5132
rect 1726 5127 1727 5131
rect 1732 5127 1733 5131
rect 1814 5128 1815 5132
rect 1819 5128 1820 5132
rect 1814 5127 1820 5128
rect 1910 5131 1917 5132
rect 1910 5127 1911 5131
rect 1916 5127 1917 5131
rect 1934 5129 1935 5133
rect 1939 5129 1940 5133
rect 4279 5131 4285 5132
rect 4279 5130 4280 5131
rect 1934 5128 1940 5129
rect 4197 5128 4280 5130
rect 1383 5126 1389 5127
rect 1542 5126 1549 5127
rect 1726 5126 1733 5127
rect 1910 5126 1917 5127
rect 4279 5127 4280 5128
rect 4284 5127 4285 5131
rect 4490 5131 4496 5132
rect 4490 5130 4491 5131
rect 4445 5128 4491 5130
rect 4279 5126 4285 5127
rect 4490 5127 4491 5128
rect 4495 5127 4496 5131
rect 5079 5131 5085 5132
rect 5079 5130 5080 5131
rect 4941 5128 5080 5130
rect 4490 5126 4496 5127
rect 4602 5127 4608 5128
rect 4602 5123 4603 5127
rect 4607 5123 4608 5127
rect 5079 5127 5080 5128
rect 5084 5127 5085 5131
rect 5079 5126 5085 5127
rect 5134 5131 5140 5132
rect 5134 5127 5135 5131
rect 5139 5127 5140 5131
rect 5134 5126 5140 5127
rect 4602 5122 4608 5123
rect 3598 5119 3604 5120
rect 3598 5118 3599 5119
rect 338 5117 344 5118
rect 110 5116 116 5117
rect 110 5112 111 5116
rect 115 5112 116 5116
rect 338 5113 339 5117
rect 343 5113 344 5117
rect 338 5112 344 5113
rect 506 5117 512 5118
rect 506 5113 507 5117
rect 511 5113 512 5117
rect 506 5112 512 5113
rect 682 5117 688 5118
rect 682 5113 683 5117
rect 687 5113 688 5117
rect 682 5112 688 5113
rect 866 5117 872 5118
rect 866 5113 867 5117
rect 871 5113 872 5117
rect 866 5112 872 5113
rect 1050 5117 1056 5118
rect 1050 5113 1051 5117
rect 1055 5113 1056 5117
rect 1050 5112 1056 5113
rect 1234 5117 1240 5118
rect 1234 5113 1235 5117
rect 1239 5113 1240 5117
rect 1234 5112 1240 5113
rect 1418 5117 1424 5118
rect 1418 5113 1419 5117
rect 1423 5113 1424 5117
rect 1418 5112 1424 5113
rect 1602 5117 1608 5118
rect 1602 5113 1603 5117
rect 1607 5113 1608 5117
rect 1602 5112 1608 5113
rect 1786 5117 1792 5118
rect 1786 5113 1787 5117
rect 1791 5113 1792 5117
rect 1786 5112 1792 5113
rect 1934 5116 1940 5117
rect 3420 5116 3599 5118
rect 1934 5112 1935 5116
rect 1939 5112 1940 5116
rect 110 5111 116 5112
rect 434 5111 440 5112
rect 434 5107 435 5111
rect 439 5110 440 5111
rect 1170 5111 1176 5112
rect 1934 5111 1940 5112
rect 2334 5115 2340 5116
rect 2334 5111 2335 5115
rect 2339 5111 2340 5115
rect 2663 5115 2669 5116
rect 2663 5114 2664 5115
rect 2613 5112 2664 5114
rect 1170 5110 1171 5111
rect 439 5108 1171 5110
rect 439 5107 440 5108
rect 434 5106 440 5107
rect 1170 5107 1171 5108
rect 1175 5107 1176 5111
rect 2334 5110 2340 5111
rect 2663 5111 2664 5112
rect 2668 5111 2669 5115
rect 2663 5110 2669 5111
rect 2838 5115 2844 5116
rect 2838 5111 2839 5115
rect 2843 5111 2844 5115
rect 3226 5115 3232 5116
rect 3226 5114 3227 5115
rect 3093 5112 3227 5114
rect 2838 5110 2844 5111
rect 3226 5111 3227 5112
rect 3231 5111 3232 5115
rect 3420 5114 3422 5116
rect 3598 5115 3599 5116
rect 3603 5115 3604 5119
rect 3598 5114 3604 5115
rect 3333 5112 3422 5114
rect 3226 5110 3232 5111
rect 3482 5111 3488 5112
rect 1170 5106 1176 5107
rect 3482 5107 3483 5111
rect 3487 5107 3488 5111
rect 3482 5106 3488 5107
rect 3838 5080 3844 5081
rect 5662 5080 5668 5081
rect 3838 5076 3839 5080
rect 3843 5076 3844 5080
rect 3838 5075 3844 5076
rect 4098 5079 4104 5080
rect 4098 5075 4099 5079
rect 4103 5075 4104 5079
rect 4098 5074 4104 5075
rect 4346 5079 4352 5080
rect 4346 5075 4347 5079
rect 4351 5075 4352 5079
rect 4346 5074 4352 5075
rect 4594 5079 4600 5080
rect 4594 5075 4595 5079
rect 4599 5075 4600 5079
rect 4594 5074 4600 5075
rect 4842 5079 4848 5080
rect 4842 5075 4843 5079
rect 4847 5075 4848 5079
rect 4842 5074 4848 5075
rect 5098 5079 5104 5080
rect 5098 5075 5099 5079
rect 5103 5075 5104 5079
rect 5662 5076 5663 5080
rect 5667 5076 5668 5080
rect 5662 5075 5668 5076
rect 5098 5074 5104 5075
rect 4279 5071 4285 5072
rect 434 5067 440 5068
rect 434 5063 435 5067
rect 439 5063 440 5067
rect 434 5062 440 5063
rect 466 5067 472 5068
rect 466 5063 467 5067
rect 471 5066 472 5067
rect 702 5067 708 5068
rect 471 5064 513 5066
rect 471 5063 472 5064
rect 466 5062 472 5063
rect 702 5063 703 5067
rect 707 5063 708 5067
rect 702 5062 708 5063
rect 831 5067 837 5068
rect 831 5063 832 5067
rect 836 5066 837 5067
rect 1014 5067 1020 5068
rect 836 5064 873 5066
rect 836 5063 837 5064
rect 831 5062 837 5063
rect 1014 5063 1015 5067
rect 1019 5066 1020 5067
rect 1330 5067 1336 5068
rect 1019 5064 1057 5066
rect 1019 5063 1020 5064
rect 1014 5062 1020 5063
rect 1330 5063 1331 5067
rect 1335 5063 1336 5067
rect 1330 5062 1336 5063
rect 1383 5067 1389 5068
rect 1383 5063 1384 5067
rect 1388 5066 1389 5067
rect 1746 5067 1752 5068
rect 1388 5064 1425 5066
rect 1388 5063 1389 5064
rect 1383 5062 1389 5063
rect 1700 5058 1702 5065
rect 1746 5063 1747 5067
rect 1751 5066 1752 5067
rect 4279 5067 4280 5071
rect 4284 5070 4285 5071
rect 5079 5071 5085 5072
rect 4284 5068 4474 5070
rect 4284 5067 4285 5068
rect 4279 5066 4285 5067
rect 4472 5066 4474 5068
rect 5079 5067 5080 5071
rect 5084 5070 5085 5071
rect 5084 5068 5226 5070
rect 5084 5067 5085 5068
rect 5079 5066 5085 5067
rect 1751 5064 1793 5066
rect 4471 5065 4477 5066
rect 1974 5064 1980 5065
rect 3798 5064 3804 5065
rect 4126 5064 4132 5065
rect 4374 5064 4380 5065
rect 1751 5063 1752 5064
rect 1746 5062 1752 5063
rect 1974 5060 1975 5064
rect 1979 5060 1980 5064
rect 1910 5059 1916 5060
rect 1974 5059 1980 5060
rect 2266 5063 2272 5064
rect 2266 5059 2267 5063
rect 2271 5059 2272 5063
rect 1910 5058 1911 5059
rect 1700 5056 1911 5058
rect 1910 5055 1911 5056
rect 1915 5055 1916 5059
rect 2266 5058 2272 5059
rect 2514 5063 2520 5064
rect 2514 5059 2515 5063
rect 2519 5059 2520 5063
rect 2514 5058 2520 5059
rect 2754 5063 2760 5064
rect 2754 5059 2755 5063
rect 2759 5059 2760 5063
rect 2754 5058 2760 5059
rect 2994 5063 3000 5064
rect 2994 5059 2995 5063
rect 2999 5059 3000 5063
rect 2994 5058 3000 5059
rect 3234 5063 3240 5064
rect 3234 5059 3235 5063
rect 3239 5059 3240 5063
rect 3234 5058 3240 5059
rect 3474 5063 3480 5064
rect 3474 5059 3475 5063
rect 3479 5059 3480 5063
rect 3798 5060 3799 5064
rect 3803 5060 3804 5064
rect 3798 5059 3804 5060
rect 3838 5063 3844 5064
rect 3838 5059 3839 5063
rect 3843 5059 3844 5063
rect 4126 5060 4127 5064
rect 4131 5060 4132 5064
rect 4126 5059 4132 5060
rect 4222 5063 4229 5064
rect 4222 5059 4223 5063
rect 4228 5059 4229 5063
rect 4374 5060 4375 5064
rect 4379 5060 4380 5064
rect 4471 5061 4472 5065
rect 4476 5061 4477 5065
rect 4471 5060 4477 5061
rect 4622 5064 4628 5065
rect 4870 5064 4876 5065
rect 5126 5064 5132 5065
rect 5224 5064 5226 5068
rect 4622 5060 4623 5064
rect 4627 5060 4628 5064
rect 4374 5059 4380 5060
rect 4622 5059 4628 5060
rect 4714 5063 4725 5064
rect 4714 5059 4715 5063
rect 4719 5059 4720 5063
rect 4724 5059 4725 5063
rect 4870 5060 4871 5064
rect 4875 5060 4876 5064
rect 4870 5059 4876 5060
rect 4966 5063 4973 5064
rect 4966 5059 4967 5063
rect 4972 5059 4973 5063
rect 5126 5060 5127 5064
rect 5131 5060 5132 5064
rect 5126 5059 5132 5060
rect 5223 5063 5229 5064
rect 5223 5059 5224 5063
rect 5228 5059 5229 5063
rect 3474 5058 3480 5059
rect 3838 5058 3844 5059
rect 4222 5058 4229 5059
rect 4714 5058 4725 5059
rect 4966 5058 4973 5059
rect 5223 5058 5229 5059
rect 5662 5063 5668 5064
rect 5662 5059 5663 5063
rect 5667 5059 5668 5063
rect 5662 5058 5668 5059
rect 1910 5054 1916 5055
rect 2663 5055 2669 5056
rect 2663 5051 2664 5055
rect 2668 5054 2669 5055
rect 3226 5055 3232 5056
rect 2668 5052 2882 5054
rect 2668 5051 2669 5052
rect 2663 5050 2669 5051
rect 2880 5050 2882 5052
rect 3226 5051 3227 5055
rect 3231 5054 3232 5055
rect 3231 5052 3362 5054
rect 3231 5051 3232 5052
rect 3226 5050 3232 5051
rect 3360 5050 3362 5052
rect 2879 5049 2885 5050
rect 3359 5049 3365 5050
rect 2294 5048 2300 5049
rect 2542 5048 2548 5049
rect 2782 5048 2788 5049
rect 1974 5047 1980 5048
rect 1974 5043 1975 5047
rect 1979 5043 1980 5047
rect 2294 5044 2295 5048
rect 2299 5044 2300 5048
rect 2294 5043 2300 5044
rect 2390 5047 2397 5048
rect 2390 5043 2391 5047
rect 2396 5043 2397 5047
rect 2542 5044 2543 5048
rect 2547 5044 2548 5048
rect 2542 5043 2548 5044
rect 2638 5047 2645 5048
rect 2638 5043 2639 5047
rect 2644 5043 2645 5047
rect 2782 5044 2783 5048
rect 2787 5044 2788 5048
rect 2879 5045 2880 5049
rect 2884 5045 2885 5049
rect 2879 5044 2885 5045
rect 3022 5048 3028 5049
rect 3262 5048 3268 5049
rect 3022 5044 3023 5048
rect 3027 5044 3028 5048
rect 2782 5043 2788 5044
rect 3022 5043 3028 5044
rect 3114 5047 3125 5048
rect 3114 5043 3115 5047
rect 3119 5043 3120 5047
rect 3124 5043 3125 5047
rect 3262 5044 3263 5048
rect 3267 5044 3268 5048
rect 3359 5045 3360 5049
rect 3364 5045 3365 5049
rect 3359 5044 3365 5045
rect 3502 5048 3508 5049
rect 3502 5044 3503 5048
rect 3507 5044 3508 5048
rect 3262 5043 3268 5044
rect 3502 5043 3508 5044
rect 3598 5047 3605 5048
rect 3598 5043 3599 5047
rect 3604 5043 3605 5047
rect 1974 5042 1980 5043
rect 2390 5042 2397 5043
rect 2638 5042 2645 5043
rect 3114 5042 3125 5043
rect 3598 5042 3605 5043
rect 3798 5047 3804 5048
rect 3798 5043 3799 5047
rect 3803 5043 3804 5047
rect 3798 5042 3804 5043
rect 630 5031 636 5032
rect 226 5027 232 5028
rect 226 5023 227 5027
rect 231 5023 232 5027
rect 226 5022 232 5023
rect 330 5027 336 5028
rect 330 5023 331 5027
rect 335 5023 336 5027
rect 630 5027 631 5031
rect 635 5027 636 5031
rect 1726 5031 1732 5032
rect 630 5026 636 5027
rect 818 5027 824 5028
rect 330 5022 336 5023
rect 818 5023 819 5027
rect 823 5023 824 5027
rect 818 5022 824 5023
rect 1090 5027 1096 5028
rect 1090 5023 1091 5027
rect 1095 5023 1096 5027
rect 1090 5022 1096 5023
rect 1466 5027 1472 5028
rect 1466 5023 1467 5027
rect 1471 5023 1472 5027
rect 1726 5027 1727 5031
rect 1731 5027 1732 5031
rect 1726 5026 1732 5027
rect 1466 5022 1472 5023
rect 1466 4995 1472 4996
rect 226 4991 232 4992
rect 226 4987 227 4991
rect 231 4990 232 4991
rect 1206 4991 1212 4992
rect 1206 4990 1207 4991
rect 231 4988 1207 4990
rect 231 4987 232 4988
rect 226 4986 232 4987
rect 1206 4987 1207 4988
rect 1211 4987 1212 4991
rect 1466 4991 1467 4995
rect 1471 4994 1472 4995
rect 1782 4995 1788 4996
rect 1782 4994 1783 4995
rect 1471 4992 1783 4994
rect 1471 4991 1472 4992
rect 1466 4990 1472 4991
rect 1782 4991 1783 4992
rect 1787 4991 1788 4995
rect 1782 4990 1788 4991
rect 1206 4986 1212 4987
rect 3838 4989 3844 4990
rect 5662 4989 5668 4990
rect 3838 4985 3839 4989
rect 3843 4985 3844 4989
rect 3838 4984 3844 4985
rect 3982 4988 3988 4989
rect 4222 4988 4228 4989
rect 4446 4988 4452 4989
rect 4654 4988 4660 4989
rect 4854 4988 4860 4989
rect 5038 4988 5044 4989
rect 5214 4988 5220 4989
rect 5390 4988 5396 4989
rect 5542 4988 5548 4989
rect 3982 4984 3983 4988
rect 3987 4984 3988 4988
rect 3982 4983 3988 4984
rect 4079 4987 4088 4988
rect 4079 4983 4080 4987
rect 4087 4983 4088 4987
rect 4222 4984 4223 4988
rect 4227 4984 4228 4988
rect 4222 4983 4228 4984
rect 4318 4987 4325 4988
rect 4318 4983 4319 4987
rect 4324 4983 4325 4987
rect 4446 4984 4447 4988
rect 4451 4984 4452 4988
rect 4446 4983 4452 4984
rect 4543 4987 4549 4988
rect 4543 4983 4544 4987
rect 4548 4986 4549 4987
rect 4602 4987 4608 4988
rect 4602 4986 4603 4987
rect 4548 4984 4603 4986
rect 4548 4983 4549 4984
rect 4079 4982 4088 4983
rect 4318 4982 4325 4983
rect 4543 4982 4549 4983
rect 4602 4983 4603 4984
rect 4607 4983 4608 4987
rect 4654 4984 4655 4988
rect 4659 4984 4660 4988
rect 4654 4983 4660 4984
rect 4750 4987 4757 4988
rect 4750 4983 4751 4987
rect 4756 4983 4757 4987
rect 4854 4984 4855 4988
rect 4859 4984 4860 4988
rect 4854 4983 4860 4984
rect 4950 4987 4957 4988
rect 4950 4983 4951 4987
rect 4956 4983 4957 4987
rect 5038 4984 5039 4988
rect 5043 4984 5044 4988
rect 5038 4983 5044 4984
rect 5135 4987 5141 4988
rect 5135 4983 5136 4987
rect 5140 4986 5141 4987
rect 5150 4987 5156 4988
rect 5150 4986 5151 4987
rect 5140 4984 5151 4986
rect 5140 4983 5141 4984
rect 4602 4982 4608 4983
rect 4750 4982 4757 4983
rect 4950 4982 4957 4983
rect 5135 4982 5141 4983
rect 5150 4983 5151 4984
rect 5155 4983 5156 4987
rect 5214 4984 5215 4988
rect 5219 4984 5220 4988
rect 5214 4983 5220 4984
rect 5311 4987 5320 4988
rect 5311 4983 5312 4987
rect 5319 4983 5320 4987
rect 5390 4984 5391 4988
rect 5395 4984 5396 4988
rect 5390 4983 5396 4984
rect 5487 4987 5493 4988
rect 5487 4983 5488 4987
rect 5492 4986 5493 4987
rect 5503 4987 5509 4988
rect 5503 4986 5504 4987
rect 5492 4984 5504 4986
rect 5492 4983 5493 4984
rect 5150 4982 5156 4983
rect 5311 4982 5320 4983
rect 5487 4982 5493 4983
rect 5503 4983 5504 4984
rect 5508 4983 5509 4987
rect 5542 4984 5543 4988
rect 5547 4984 5548 4988
rect 5542 4983 5548 4984
rect 5634 4987 5645 4988
rect 5634 4983 5635 4987
rect 5639 4983 5640 4987
rect 5644 4983 5645 4987
rect 5662 4985 5663 4989
rect 5667 4985 5668 4989
rect 5662 4984 5668 4985
rect 5503 4982 5509 4983
rect 5634 4982 5645 4983
rect 110 4980 116 4981
rect 1934 4980 1940 4981
rect 110 4976 111 4980
rect 115 4976 116 4980
rect 110 4975 116 4976
rect 130 4979 136 4980
rect 130 4975 131 4979
rect 135 4975 136 4979
rect 130 4974 136 4975
rect 322 4979 328 4980
rect 322 4975 323 4979
rect 327 4975 328 4979
rect 322 4974 328 4975
rect 554 4979 560 4980
rect 554 4975 555 4979
rect 559 4975 560 4979
rect 554 4974 560 4975
rect 810 4979 816 4980
rect 810 4975 811 4979
rect 815 4975 816 4979
rect 810 4974 816 4975
rect 1082 4979 1088 4980
rect 1082 4975 1083 4979
rect 1087 4975 1088 4979
rect 1082 4974 1088 4975
rect 1370 4979 1376 4980
rect 1370 4975 1371 4979
rect 1375 4975 1376 4979
rect 1370 4974 1376 4975
rect 1658 4979 1664 4980
rect 1658 4975 1659 4979
rect 1663 4975 1664 4979
rect 1934 4976 1935 4980
rect 1939 4976 1940 4980
rect 1934 4975 1940 4976
rect 1658 4974 1664 4975
rect 3954 4973 3960 4974
rect 3838 4972 3844 4973
rect 1330 4971 1336 4972
rect 1330 4967 1331 4971
rect 1335 4970 1336 4971
rect 1335 4968 1498 4970
rect 1335 4967 1336 4968
rect 1330 4966 1336 4967
rect 158 4964 164 4965
rect 350 4964 356 4965
rect 582 4964 588 4965
rect 838 4964 844 4965
rect 1110 4964 1116 4965
rect 1398 4964 1404 4965
rect 1496 4964 1498 4968
rect 3838 4968 3839 4972
rect 3843 4968 3844 4972
rect 3954 4969 3955 4973
rect 3959 4969 3960 4973
rect 3954 4968 3960 4969
rect 4194 4973 4200 4974
rect 4194 4969 4195 4973
rect 4199 4969 4200 4973
rect 4194 4968 4200 4969
rect 4418 4973 4424 4974
rect 4418 4969 4419 4973
rect 4423 4969 4424 4973
rect 4418 4968 4424 4969
rect 4626 4973 4632 4974
rect 4626 4969 4627 4973
rect 4631 4969 4632 4973
rect 4626 4968 4632 4969
rect 4826 4973 4832 4974
rect 4826 4969 4827 4973
rect 4831 4969 4832 4973
rect 4826 4968 4832 4969
rect 5010 4973 5016 4974
rect 5010 4969 5011 4973
rect 5015 4969 5016 4973
rect 5010 4968 5016 4969
rect 5186 4973 5192 4974
rect 5186 4969 5187 4973
rect 5191 4969 5192 4973
rect 5186 4968 5192 4969
rect 5362 4973 5368 4974
rect 5362 4969 5363 4973
rect 5367 4969 5368 4973
rect 5362 4968 5368 4969
rect 5514 4973 5520 4974
rect 5514 4969 5515 4973
rect 5519 4969 5520 4973
rect 5514 4968 5520 4969
rect 5662 4972 5668 4973
rect 5662 4968 5663 4972
rect 5667 4968 5668 4972
rect 3838 4967 3844 4968
rect 5662 4967 5668 4968
rect 1686 4964 1692 4965
rect 110 4963 116 4964
rect 110 4959 111 4963
rect 115 4959 116 4963
rect 158 4960 159 4964
rect 163 4960 164 4964
rect 158 4959 164 4960
rect 255 4963 261 4964
rect 255 4959 256 4963
rect 260 4962 261 4963
rect 330 4963 336 4964
rect 330 4962 331 4963
rect 260 4960 331 4962
rect 260 4959 261 4960
rect 110 4958 116 4959
rect 255 4958 261 4959
rect 330 4959 331 4960
rect 335 4959 336 4963
rect 350 4960 351 4964
rect 355 4960 356 4964
rect 350 4959 356 4960
rect 446 4963 453 4964
rect 446 4959 447 4963
rect 452 4959 453 4963
rect 582 4960 583 4964
rect 587 4960 588 4964
rect 582 4959 588 4960
rect 679 4963 685 4964
rect 679 4959 680 4963
rect 684 4962 685 4963
rect 818 4963 824 4964
rect 818 4962 819 4963
rect 684 4960 819 4962
rect 684 4959 685 4960
rect 330 4958 336 4959
rect 446 4958 453 4959
rect 679 4958 685 4959
rect 818 4959 819 4960
rect 823 4959 824 4963
rect 838 4960 839 4964
rect 843 4960 844 4964
rect 838 4959 844 4960
rect 935 4963 941 4964
rect 935 4959 936 4963
rect 940 4962 941 4963
rect 1090 4963 1096 4964
rect 1090 4962 1091 4963
rect 940 4960 1091 4962
rect 940 4959 941 4960
rect 818 4958 824 4959
rect 935 4958 941 4959
rect 1090 4959 1091 4960
rect 1095 4959 1096 4963
rect 1110 4960 1111 4964
rect 1115 4960 1116 4964
rect 1110 4959 1116 4960
rect 1206 4963 1213 4964
rect 1206 4959 1207 4963
rect 1212 4959 1213 4963
rect 1398 4960 1399 4964
rect 1403 4960 1404 4964
rect 1398 4959 1404 4960
rect 1495 4963 1501 4964
rect 1495 4959 1496 4963
rect 1500 4959 1501 4963
rect 1686 4960 1687 4964
rect 1691 4960 1692 4964
rect 1686 4959 1692 4960
rect 1782 4963 1789 4964
rect 1782 4959 1783 4963
rect 1788 4959 1789 4963
rect 1090 4958 1096 4959
rect 1206 4958 1213 4959
rect 1495 4958 1501 4959
rect 1782 4958 1789 4959
rect 1934 4963 1940 4964
rect 1934 4959 1935 4963
rect 1939 4959 1940 4963
rect 1934 4958 1940 4959
rect 1974 4957 1980 4958
rect 3798 4957 3804 4958
rect 1974 4953 1975 4957
rect 1979 4953 1980 4957
rect 1974 4952 1980 4953
rect 2182 4956 2188 4957
rect 2318 4956 2324 4957
rect 2454 4956 2460 4957
rect 2598 4956 2604 4957
rect 2742 4956 2748 4957
rect 2894 4956 2900 4957
rect 3046 4956 3052 4957
rect 3198 4956 3204 4957
rect 3350 4956 3356 4957
rect 2182 4952 2183 4956
rect 2187 4952 2188 4956
rect 2182 4951 2188 4952
rect 2279 4955 2288 4956
rect 2279 4951 2280 4955
rect 2287 4951 2288 4955
rect 2318 4952 2319 4956
rect 2323 4952 2324 4956
rect 2318 4951 2324 4952
rect 2415 4955 2424 4956
rect 2415 4951 2416 4955
rect 2423 4951 2424 4955
rect 2454 4952 2455 4956
rect 2459 4952 2460 4956
rect 2454 4951 2460 4952
rect 2551 4955 2560 4956
rect 2551 4951 2552 4955
rect 2559 4951 2560 4955
rect 2598 4952 2599 4956
rect 2603 4952 2604 4956
rect 2598 4951 2604 4952
rect 2690 4955 2701 4956
rect 2690 4951 2691 4955
rect 2695 4951 2696 4955
rect 2700 4951 2701 4955
rect 2742 4952 2743 4956
rect 2747 4952 2748 4956
rect 2742 4951 2748 4952
rect 2838 4955 2845 4956
rect 2838 4951 2839 4955
rect 2844 4951 2845 4955
rect 2894 4952 2895 4956
rect 2899 4952 2900 4956
rect 2894 4951 2900 4952
rect 2986 4955 2997 4956
rect 2986 4951 2987 4955
rect 2991 4951 2992 4955
rect 2996 4951 2997 4955
rect 3046 4952 3047 4956
rect 3051 4952 3052 4956
rect 3046 4951 3052 4952
rect 3142 4955 3149 4956
rect 3142 4951 3143 4955
rect 3148 4951 3149 4955
rect 3198 4952 3199 4956
rect 3203 4952 3204 4956
rect 3198 4951 3204 4952
rect 3294 4955 3301 4956
rect 3294 4951 3295 4955
rect 3300 4951 3301 4955
rect 3350 4952 3351 4956
rect 3355 4952 3356 4956
rect 3350 4951 3356 4952
rect 3447 4955 3453 4956
rect 3447 4951 3448 4955
rect 3452 4954 3453 4955
rect 3482 4955 3488 4956
rect 3482 4954 3483 4955
rect 3452 4952 3483 4954
rect 3452 4951 3453 4952
rect 2279 4950 2288 4951
rect 2415 4950 2424 4951
rect 2551 4950 2560 4951
rect 2690 4950 2701 4951
rect 2838 4950 2845 4951
rect 2986 4950 2997 4951
rect 3142 4950 3149 4951
rect 3294 4950 3301 4951
rect 3447 4950 3453 4951
rect 3482 4951 3483 4952
rect 3487 4951 3488 4955
rect 3798 4953 3799 4957
rect 3803 4953 3804 4957
rect 3798 4952 3804 4953
rect 3482 4950 3488 4951
rect 2154 4941 2160 4942
rect 1974 4940 1980 4941
rect 1974 4936 1975 4940
rect 1979 4936 1980 4940
rect 2154 4937 2155 4941
rect 2159 4937 2160 4941
rect 2154 4936 2160 4937
rect 2290 4941 2296 4942
rect 2290 4937 2291 4941
rect 2295 4937 2296 4941
rect 2290 4936 2296 4937
rect 2426 4941 2432 4942
rect 2426 4937 2427 4941
rect 2431 4937 2432 4941
rect 2426 4936 2432 4937
rect 2570 4941 2576 4942
rect 2570 4937 2571 4941
rect 2575 4937 2576 4941
rect 2570 4936 2576 4937
rect 2714 4941 2720 4942
rect 2714 4937 2715 4941
rect 2719 4937 2720 4941
rect 2714 4936 2720 4937
rect 2866 4941 2872 4942
rect 2866 4937 2867 4941
rect 2871 4937 2872 4941
rect 2866 4936 2872 4937
rect 3018 4941 3024 4942
rect 3018 4937 3019 4941
rect 3023 4937 3024 4941
rect 3018 4936 3024 4937
rect 3170 4941 3176 4942
rect 3170 4937 3171 4941
rect 3175 4937 3176 4941
rect 3170 4936 3176 4937
rect 3322 4941 3328 4942
rect 3322 4937 3323 4941
rect 3327 4937 3328 4941
rect 3322 4936 3328 4937
rect 3798 4940 3804 4941
rect 3798 4936 3799 4940
rect 3803 4936 3804 4940
rect 1974 4935 1980 4936
rect 3798 4935 3804 4936
rect 4214 4923 4220 4924
rect 4052 4914 4054 4921
rect 4214 4919 4215 4923
rect 4219 4919 4220 4923
rect 4214 4918 4220 4919
rect 4426 4923 4432 4924
rect 4426 4919 4427 4923
rect 4431 4919 4432 4923
rect 4966 4923 4972 4924
rect 4966 4922 4967 4923
rect 4426 4918 4432 4919
rect 4318 4915 4324 4916
rect 4318 4914 4319 4915
rect 4052 4912 4319 4914
rect 4318 4911 4319 4912
rect 4323 4911 4324 4915
rect 4724 4914 4726 4921
rect 4925 4920 4967 4922
rect 4966 4919 4967 4920
rect 4971 4919 4972 4923
rect 5150 4923 5156 4924
rect 4966 4918 4972 4919
rect 4950 4915 4956 4916
rect 4950 4914 4951 4915
rect 4724 4912 4951 4914
rect 4318 4910 4324 4911
rect 4950 4911 4951 4912
rect 4955 4911 4956 4915
rect 5108 4914 5110 4921
rect 5150 4919 5151 4923
rect 5155 4922 5156 4923
rect 5314 4923 5320 4924
rect 5155 4920 5193 4922
rect 5155 4919 5156 4920
rect 5150 4918 5156 4919
rect 5314 4919 5315 4923
rect 5319 4922 5320 4923
rect 5503 4923 5509 4924
rect 5319 4920 5369 4922
rect 5319 4919 5320 4920
rect 5314 4918 5320 4919
rect 5503 4919 5504 4923
rect 5508 4922 5509 4923
rect 5508 4920 5521 4922
rect 5508 4919 5509 4920
rect 5503 4918 5509 4919
rect 5494 4915 5500 4916
rect 5494 4914 5495 4915
rect 5108 4912 5495 4914
rect 4950 4910 4956 4911
rect 5494 4911 5495 4912
rect 5499 4911 5500 4915
rect 5494 4910 5500 4911
rect 2282 4891 2288 4892
rect 2252 4882 2254 4889
rect 2282 4887 2283 4891
rect 2287 4890 2288 4891
rect 2418 4891 2424 4892
rect 2287 4888 2297 4890
rect 2287 4887 2288 4888
rect 2282 4886 2288 4887
rect 2418 4887 2419 4891
rect 2423 4890 2424 4891
rect 2554 4891 2560 4892
rect 2423 4888 2433 4890
rect 2423 4887 2424 4888
rect 2418 4886 2424 4887
rect 2554 4887 2555 4891
rect 2559 4890 2560 4891
rect 2850 4891 2856 4892
rect 2559 4888 2577 4890
rect 2559 4887 2560 4888
rect 2554 4886 2560 4887
rect 2390 4883 2396 4884
rect 2390 4882 2391 4883
rect 110 4881 116 4882
rect 1934 4881 1940 4882
rect 110 4877 111 4881
rect 115 4877 116 4881
rect 110 4876 116 4877
rect 158 4880 164 4881
rect 294 4880 300 4881
rect 430 4880 436 4881
rect 566 4880 572 4881
rect 702 4880 708 4881
rect 158 4876 159 4880
rect 163 4876 164 4880
rect 158 4875 164 4876
rect 250 4879 261 4880
rect 250 4875 251 4879
rect 255 4875 256 4879
rect 260 4875 261 4879
rect 294 4876 295 4880
rect 299 4876 300 4880
rect 294 4875 300 4876
rect 386 4879 397 4880
rect 386 4875 387 4879
rect 391 4875 392 4879
rect 396 4875 397 4879
rect 430 4876 431 4880
rect 435 4876 436 4880
rect 430 4875 436 4876
rect 527 4879 536 4880
rect 527 4875 528 4879
rect 535 4875 536 4879
rect 566 4876 567 4880
rect 571 4876 572 4880
rect 566 4875 572 4876
rect 663 4879 672 4880
rect 663 4875 664 4879
rect 671 4875 672 4879
rect 702 4876 703 4880
rect 707 4876 708 4880
rect 702 4875 708 4876
rect 798 4879 805 4880
rect 798 4875 799 4879
rect 804 4875 805 4879
rect 1934 4877 1935 4881
rect 1939 4877 1940 4881
rect 2252 4880 2391 4882
rect 2390 4879 2391 4880
rect 2395 4879 2396 4883
rect 2812 4882 2814 4889
rect 2850 4887 2851 4891
rect 2855 4890 2856 4891
rect 3002 4891 3008 4892
rect 2855 4888 2873 4890
rect 2855 4887 2856 4888
rect 2850 4886 2856 4887
rect 3002 4887 3003 4891
rect 3007 4890 3008 4891
rect 3142 4891 3148 4892
rect 3007 4888 3025 4890
rect 3007 4887 3008 4888
rect 3002 4886 3008 4887
rect 3142 4887 3143 4891
rect 3147 4890 3148 4891
rect 3294 4891 3300 4892
rect 3147 4888 3177 4890
rect 3147 4887 3148 4888
rect 3142 4886 3148 4887
rect 3294 4887 3295 4891
rect 3299 4890 3300 4891
rect 3299 4888 3329 4890
rect 3299 4887 3300 4888
rect 3294 4886 3300 4887
rect 2986 4883 2992 4884
rect 2986 4882 2987 4883
rect 2812 4880 2987 4882
rect 2390 4878 2396 4879
rect 2986 4879 2987 4880
rect 2991 4879 2992 4883
rect 2986 4878 2992 4879
rect 1934 4876 1940 4877
rect 250 4874 261 4875
rect 386 4874 397 4875
rect 527 4874 536 4875
rect 663 4874 672 4875
rect 798 4874 805 4875
rect 4630 4871 4636 4872
rect 4630 4870 4631 4871
rect 4459 4868 4631 4870
rect 4063 4867 4069 4868
rect 4063 4866 4064 4867
rect 130 4865 136 4866
rect 110 4864 116 4865
rect 110 4860 111 4864
rect 115 4860 116 4864
rect 130 4861 131 4865
rect 135 4861 136 4865
rect 130 4860 136 4861
rect 266 4865 272 4866
rect 266 4861 267 4865
rect 271 4861 272 4865
rect 266 4860 272 4861
rect 402 4865 408 4866
rect 402 4861 403 4865
rect 407 4861 408 4865
rect 402 4860 408 4861
rect 538 4865 544 4866
rect 538 4861 539 4865
rect 543 4861 544 4865
rect 538 4860 544 4861
rect 674 4865 680 4866
rect 674 4861 675 4865
rect 679 4861 680 4865
rect 674 4860 680 4861
rect 1934 4864 1940 4865
rect 3957 4864 4064 4866
rect 1934 4860 1935 4864
rect 1939 4860 1940 4864
rect 4063 4863 4064 4864
rect 4068 4863 4069 4867
rect 4063 4862 4069 4863
rect 4082 4867 4088 4868
rect 4082 4863 4083 4867
rect 4087 4863 4088 4867
rect 4459 4866 4461 4868
rect 4630 4867 4631 4868
rect 4635 4867 4636 4871
rect 4630 4866 4636 4867
rect 4750 4867 4756 4868
rect 4397 4864 4461 4866
rect 4082 4862 4088 4863
rect 4602 4863 4608 4864
rect 110 4859 116 4860
rect 1934 4859 1940 4860
rect 4602 4859 4603 4863
rect 4607 4859 4608 4863
rect 4750 4863 4751 4867
rect 4755 4863 4756 4867
rect 5330 4867 5336 4868
rect 5330 4866 5331 4867
rect 5309 4864 5331 4866
rect 4750 4862 4756 4863
rect 4882 4863 4888 4864
rect 4602 4858 4608 4859
rect 4882 4859 4883 4863
rect 4887 4859 4888 4863
rect 4882 4858 4888 4859
rect 5050 4863 5056 4864
rect 5050 4859 5051 4863
rect 5055 4859 5056 4863
rect 5330 4863 5331 4864
rect 5335 4863 5336 4867
rect 5634 4867 5640 4868
rect 5634 4866 5635 4867
rect 5613 4864 5635 4866
rect 5330 4862 5336 4863
rect 5378 4863 5384 4864
rect 5050 4858 5056 4859
rect 5378 4859 5379 4863
rect 5383 4859 5384 4863
rect 5634 4863 5635 4864
rect 5639 4863 5640 4867
rect 5634 4862 5640 4863
rect 5378 4858 5384 4859
rect 2690 4855 2696 4856
rect 2690 4854 2691 4855
rect 2564 4852 2691 4854
rect 2564 4850 2566 4852
rect 2690 4851 2691 4852
rect 2695 4851 2696 4855
rect 3302 4855 3308 4856
rect 3302 4854 3303 4855
rect 3176 4852 3303 4854
rect 2690 4850 2696 4851
rect 3018 4851 3024 4852
rect 3018 4850 3019 4851
rect 2525 4848 2566 4850
rect 2973 4848 3019 4850
rect 2578 4847 2584 4848
rect 2578 4843 2579 4847
rect 2583 4843 2584 4847
rect 2578 4842 2584 4843
rect 2730 4847 2736 4848
rect 2730 4843 2731 4847
rect 2735 4843 2736 4847
rect 3018 4847 3019 4848
rect 3023 4847 3024 4851
rect 3176 4850 3178 4852
rect 3302 4851 3303 4852
rect 3307 4851 3308 4855
rect 3302 4850 3308 4851
rect 3125 4848 3178 4850
rect 3018 4846 3024 4847
rect 2730 4842 2736 4843
rect 3272 4842 3274 4845
rect 3342 4843 3348 4844
rect 3342 4842 3343 4843
rect 3272 4840 3343 4842
rect 3342 4839 3343 4840
rect 3347 4839 3348 4843
rect 3342 4838 3348 4839
rect 3838 4816 3844 4817
rect 5662 4816 5668 4817
rect 446 4815 452 4816
rect 229 4812 261 4814
rect 365 4812 406 4814
rect 259 4806 261 4812
rect 386 4807 392 4808
rect 386 4806 387 4807
rect 259 4804 387 4806
rect 386 4803 387 4804
rect 391 4803 392 4807
rect 404 4806 406 4812
rect 446 4811 447 4815
rect 451 4811 452 4815
rect 446 4810 452 4811
rect 530 4815 536 4816
rect 530 4811 531 4815
rect 535 4814 536 4815
rect 666 4815 672 4816
rect 535 4812 545 4814
rect 535 4811 536 4812
rect 530 4810 536 4811
rect 666 4811 667 4815
rect 671 4814 672 4815
rect 671 4812 681 4814
rect 3838 4812 3839 4816
rect 3843 4812 3844 4816
rect 671 4811 672 4812
rect 3838 4811 3844 4812
rect 3858 4815 3864 4816
rect 3858 4811 3859 4815
rect 3863 4811 3864 4815
rect 666 4810 672 4811
rect 3858 4810 3864 4811
rect 4074 4815 4080 4816
rect 4074 4811 4075 4815
rect 4079 4811 4080 4815
rect 4074 4810 4080 4811
rect 4298 4815 4304 4816
rect 4298 4811 4299 4815
rect 4303 4811 4304 4815
rect 4298 4810 4304 4811
rect 4506 4815 4512 4816
rect 4506 4811 4507 4815
rect 4511 4811 4512 4815
rect 4506 4810 4512 4811
rect 4698 4815 4704 4816
rect 4698 4811 4699 4815
rect 4703 4811 4704 4815
rect 4698 4810 4704 4811
rect 4874 4815 4880 4816
rect 4874 4811 4875 4815
rect 4879 4811 4880 4815
rect 4874 4810 4880 4811
rect 5042 4815 5048 4816
rect 5042 4811 5043 4815
rect 5047 4811 5048 4815
rect 5042 4810 5048 4811
rect 5210 4815 5216 4816
rect 5210 4811 5211 4815
rect 5215 4811 5216 4815
rect 5210 4810 5216 4811
rect 5370 4815 5376 4816
rect 5370 4811 5371 4815
rect 5375 4811 5376 4815
rect 5370 4810 5376 4811
rect 5514 4815 5520 4816
rect 5514 4811 5515 4815
rect 5519 4811 5520 4815
rect 5662 4812 5663 4816
rect 5667 4812 5668 4816
rect 5662 4811 5668 4812
rect 5514 4810 5520 4811
rect 798 4807 804 4808
rect 798 4806 799 4807
rect 404 4804 799 4806
rect 386 4802 392 4803
rect 798 4803 799 4804
rect 803 4803 804 4807
rect 798 4802 804 4803
rect 4063 4807 4069 4808
rect 4063 4803 4064 4807
rect 4068 4806 4069 4807
rect 4068 4804 4202 4806
rect 4068 4803 4069 4804
rect 4063 4802 4069 4803
rect 1974 4800 1980 4801
rect 3798 4800 3804 4801
rect 3886 4800 3892 4801
rect 4102 4800 4108 4801
rect 4200 4800 4202 4804
rect 4326 4800 4332 4801
rect 4534 4800 4540 4801
rect 4726 4800 4732 4801
rect 4902 4800 4908 4801
rect 5070 4800 5076 4801
rect 5238 4800 5244 4801
rect 5398 4800 5404 4801
rect 5542 4800 5548 4801
rect 1974 4796 1975 4800
rect 1979 4796 1980 4800
rect 1974 4795 1980 4796
rect 2426 4799 2432 4800
rect 2426 4795 2427 4799
rect 2431 4795 2432 4799
rect 2426 4794 2432 4795
rect 2570 4799 2576 4800
rect 2570 4795 2571 4799
rect 2575 4795 2576 4799
rect 2570 4794 2576 4795
rect 2722 4799 2728 4800
rect 2722 4795 2723 4799
rect 2727 4795 2728 4799
rect 2722 4794 2728 4795
rect 2874 4799 2880 4800
rect 2874 4795 2875 4799
rect 2879 4795 2880 4799
rect 2874 4794 2880 4795
rect 3026 4799 3032 4800
rect 3026 4795 3027 4799
rect 3031 4795 3032 4799
rect 3026 4794 3032 4795
rect 3178 4799 3184 4800
rect 3178 4795 3179 4799
rect 3183 4795 3184 4799
rect 3798 4796 3799 4800
rect 3803 4796 3804 4800
rect 3798 4795 3804 4796
rect 3838 4799 3844 4800
rect 3838 4795 3839 4799
rect 3843 4795 3844 4799
rect 3886 4796 3887 4800
rect 3891 4796 3892 4800
rect 3886 4795 3892 4796
rect 3982 4799 3989 4800
rect 3982 4795 3983 4799
rect 3988 4795 3989 4799
rect 4102 4796 4103 4800
rect 4107 4796 4108 4800
rect 4102 4795 4108 4796
rect 4199 4799 4205 4800
rect 4199 4795 4200 4799
rect 4204 4795 4205 4799
rect 4326 4796 4327 4800
rect 4331 4796 4332 4800
rect 4326 4795 4332 4796
rect 4423 4799 4432 4800
rect 4423 4795 4424 4799
rect 4431 4795 4432 4799
rect 4534 4796 4535 4800
rect 4539 4796 4540 4800
rect 4534 4795 4540 4796
rect 4630 4799 4637 4800
rect 4630 4795 4631 4799
rect 4636 4795 4637 4799
rect 4726 4796 4727 4800
rect 4731 4796 4732 4800
rect 4726 4795 4732 4796
rect 4823 4799 4829 4800
rect 4823 4795 4824 4799
rect 4828 4798 4829 4799
rect 4882 4799 4888 4800
rect 4882 4798 4883 4799
rect 4828 4796 4883 4798
rect 4828 4795 4829 4796
rect 3178 4794 3184 4795
rect 3838 4794 3844 4795
rect 3982 4794 3989 4795
rect 4199 4794 4205 4795
rect 4423 4794 4432 4795
rect 4630 4794 4637 4795
rect 4823 4794 4829 4795
rect 4882 4795 4883 4796
rect 4887 4795 4888 4799
rect 4902 4796 4903 4800
rect 4907 4796 4908 4800
rect 4902 4795 4908 4796
rect 4999 4799 5005 4800
rect 4999 4795 5000 4799
rect 5004 4798 5005 4799
rect 5050 4799 5056 4800
rect 5050 4798 5051 4799
rect 5004 4796 5051 4798
rect 5004 4795 5005 4796
rect 4882 4794 4888 4795
rect 4999 4794 5005 4795
rect 5050 4795 5051 4796
rect 5055 4795 5056 4799
rect 5070 4796 5071 4800
rect 5075 4796 5076 4800
rect 5070 4795 5076 4796
rect 5166 4799 5173 4800
rect 5166 4795 5167 4799
rect 5172 4795 5173 4799
rect 5238 4796 5239 4800
rect 5243 4796 5244 4800
rect 5238 4795 5244 4796
rect 5335 4799 5341 4800
rect 5335 4795 5336 4799
rect 5340 4798 5341 4799
rect 5378 4799 5384 4800
rect 5378 4798 5379 4799
rect 5340 4796 5379 4798
rect 5340 4795 5341 4796
rect 5050 4794 5056 4795
rect 5166 4794 5173 4795
rect 5335 4794 5341 4795
rect 5378 4795 5379 4796
rect 5383 4795 5384 4799
rect 5398 4796 5399 4800
rect 5403 4796 5404 4800
rect 5398 4795 5404 4796
rect 5494 4799 5501 4800
rect 5494 4795 5495 4799
rect 5500 4795 5501 4799
rect 5542 4796 5543 4800
rect 5547 4796 5548 4800
rect 5542 4795 5548 4796
rect 5638 4799 5645 4800
rect 5638 4795 5639 4799
rect 5644 4795 5645 4799
rect 5378 4794 5384 4795
rect 5494 4794 5501 4795
rect 5638 4794 5645 4795
rect 5662 4799 5668 4800
rect 5662 4795 5663 4799
rect 5667 4795 5668 4799
rect 5662 4794 5668 4795
rect 3018 4791 3024 4792
rect 3018 4787 3019 4791
rect 3023 4790 3024 4791
rect 3023 4788 3154 4790
rect 3023 4787 3024 4788
rect 3018 4786 3024 4787
rect 2454 4784 2460 4785
rect 2598 4784 2604 4785
rect 2750 4784 2756 4785
rect 2902 4784 2908 4785
rect 3054 4784 3060 4785
rect 3152 4784 3154 4788
rect 3206 4784 3212 4785
rect 1974 4783 1980 4784
rect 1974 4779 1975 4783
rect 1979 4779 1980 4783
rect 2454 4780 2455 4784
rect 2459 4780 2460 4784
rect 2454 4779 2460 4780
rect 2551 4783 2557 4784
rect 2551 4779 2552 4783
rect 2556 4782 2557 4783
rect 2578 4783 2584 4784
rect 2578 4782 2579 4783
rect 2556 4780 2579 4782
rect 2556 4779 2557 4780
rect 1974 4778 1980 4779
rect 2551 4778 2557 4779
rect 2578 4779 2579 4780
rect 2583 4779 2584 4783
rect 2598 4780 2599 4784
rect 2603 4780 2604 4784
rect 2598 4779 2604 4780
rect 2695 4783 2701 4784
rect 2695 4779 2696 4783
rect 2700 4782 2701 4783
rect 2730 4783 2736 4784
rect 2730 4782 2731 4783
rect 2700 4780 2731 4782
rect 2700 4779 2701 4780
rect 2578 4778 2584 4779
rect 2695 4778 2701 4779
rect 2730 4779 2731 4780
rect 2735 4779 2736 4783
rect 2750 4780 2751 4784
rect 2755 4780 2756 4784
rect 2750 4779 2756 4780
rect 2847 4783 2856 4784
rect 2847 4779 2848 4783
rect 2855 4779 2856 4783
rect 2902 4780 2903 4784
rect 2907 4780 2908 4784
rect 2902 4779 2908 4780
rect 2999 4783 3008 4784
rect 2999 4779 3000 4783
rect 3007 4779 3008 4783
rect 3054 4780 3055 4784
rect 3059 4780 3060 4784
rect 3054 4779 3060 4780
rect 3151 4783 3157 4784
rect 3151 4779 3152 4783
rect 3156 4779 3157 4783
rect 3206 4780 3207 4784
rect 3211 4780 3212 4784
rect 3206 4779 3212 4780
rect 3302 4783 3309 4784
rect 3302 4779 3303 4783
rect 3308 4779 3309 4783
rect 2730 4778 2736 4779
rect 2847 4778 2856 4779
rect 2999 4778 3008 4779
rect 3151 4778 3157 4779
rect 3302 4778 3309 4779
rect 3798 4783 3804 4784
rect 3798 4779 3799 4783
rect 3803 4779 3804 4783
rect 3798 4778 3804 4779
rect 250 4771 256 4772
rect 250 4770 251 4771
rect 229 4768 251 4770
rect 250 4767 251 4768
rect 255 4767 256 4771
rect 250 4766 256 4767
rect 274 4767 280 4768
rect 274 4763 275 4767
rect 279 4763 280 4767
rect 274 4762 280 4763
rect 410 4767 416 4768
rect 410 4763 411 4767
rect 415 4763 416 4767
rect 410 4762 416 4763
rect 546 4767 552 4768
rect 546 4763 547 4767
rect 551 4763 552 4767
rect 546 4762 552 4763
rect 682 4767 688 4768
rect 682 4763 683 4767
rect 687 4763 688 4767
rect 682 4762 688 4763
rect 4602 4755 4608 4756
rect 4602 4751 4603 4755
rect 4607 4754 4608 4755
rect 4607 4752 5042 4754
rect 4607 4751 4608 4752
rect 4602 4750 4608 4751
rect 3838 4741 3844 4742
rect 3838 4737 3839 4741
rect 3843 4737 3844 4741
rect 3838 4736 3844 4737
rect 4942 4740 4948 4741
rect 5040 4740 5042 4752
rect 5662 4741 5668 4742
rect 5086 4740 5092 4741
rect 5238 4740 5244 4741
rect 5398 4740 5404 4741
rect 5542 4740 5548 4741
rect 4942 4736 4943 4740
rect 4947 4736 4948 4740
rect 4942 4735 4948 4736
rect 5039 4739 5045 4740
rect 5039 4735 5040 4739
rect 5044 4735 5045 4739
rect 5086 4736 5087 4740
rect 5091 4736 5092 4740
rect 5086 4735 5092 4736
rect 5183 4739 5189 4740
rect 5183 4735 5184 4739
rect 5188 4738 5189 4739
rect 5199 4739 5205 4740
rect 5199 4738 5200 4739
rect 5188 4736 5200 4738
rect 5188 4735 5189 4736
rect 5039 4734 5045 4735
rect 5183 4734 5189 4735
rect 5199 4735 5200 4736
rect 5204 4735 5205 4739
rect 5238 4736 5239 4740
rect 5243 4736 5244 4740
rect 5238 4735 5244 4736
rect 5330 4739 5341 4740
rect 5330 4735 5331 4739
rect 5335 4735 5336 4739
rect 5340 4735 5341 4739
rect 5398 4736 5399 4740
rect 5403 4736 5404 4740
rect 5398 4735 5404 4736
rect 5490 4739 5501 4740
rect 5490 4735 5491 4739
rect 5495 4735 5496 4739
rect 5500 4735 5501 4739
rect 5542 4736 5543 4740
rect 5547 4736 5548 4740
rect 5542 4735 5548 4736
rect 5639 4739 5645 4740
rect 5639 4735 5640 4739
rect 5644 4738 5645 4739
rect 5647 4739 5653 4740
rect 5647 4738 5648 4739
rect 5644 4736 5648 4738
rect 5644 4735 5645 4736
rect 5199 4734 5205 4735
rect 5330 4734 5341 4735
rect 5490 4734 5501 4735
rect 5639 4734 5645 4735
rect 5647 4735 5648 4736
rect 5652 4735 5653 4739
rect 5662 4737 5663 4741
rect 5667 4737 5668 4741
rect 5662 4736 5668 4737
rect 5647 4734 5653 4735
rect 4914 4725 4920 4726
rect 3838 4724 3844 4725
rect 1974 4721 1980 4722
rect 3798 4721 3804 4722
rect 110 4720 116 4721
rect 1934 4720 1940 4721
rect 110 4716 111 4720
rect 115 4716 116 4720
rect 110 4715 116 4716
rect 130 4719 136 4720
rect 130 4715 131 4719
rect 135 4715 136 4719
rect 130 4714 136 4715
rect 266 4719 272 4720
rect 266 4715 267 4719
rect 271 4715 272 4719
rect 266 4714 272 4715
rect 402 4719 408 4720
rect 402 4715 403 4719
rect 407 4715 408 4719
rect 402 4714 408 4715
rect 538 4719 544 4720
rect 538 4715 539 4719
rect 543 4715 544 4719
rect 538 4714 544 4715
rect 674 4719 680 4720
rect 674 4715 675 4719
rect 679 4715 680 4719
rect 1934 4716 1935 4720
rect 1939 4716 1940 4720
rect 1974 4717 1975 4721
rect 1979 4717 1980 4721
rect 1974 4716 1980 4717
rect 2022 4720 2028 4721
rect 2158 4720 2164 4721
rect 2294 4720 2300 4721
rect 2430 4720 2436 4721
rect 2566 4720 2572 4721
rect 2702 4720 2708 4721
rect 2838 4720 2844 4721
rect 2974 4720 2980 4721
rect 3110 4720 3116 4721
rect 3246 4720 3252 4721
rect 3398 4720 3404 4721
rect 3542 4720 3548 4721
rect 3678 4720 3684 4721
rect 2022 4716 2023 4720
rect 2027 4716 2028 4720
rect 1934 4715 1940 4716
rect 2022 4715 2028 4716
rect 2119 4719 2128 4720
rect 2119 4715 2120 4719
rect 2127 4715 2128 4719
rect 2158 4716 2159 4720
rect 2163 4716 2164 4720
rect 2158 4715 2164 4716
rect 2255 4719 2264 4720
rect 2255 4715 2256 4719
rect 2263 4715 2264 4719
rect 2294 4716 2295 4720
rect 2299 4716 2300 4720
rect 2294 4715 2300 4716
rect 2391 4719 2400 4720
rect 2391 4715 2392 4719
rect 2399 4715 2400 4719
rect 2430 4716 2431 4720
rect 2435 4716 2436 4720
rect 2430 4715 2436 4716
rect 2527 4719 2536 4720
rect 2527 4715 2528 4719
rect 2535 4715 2536 4719
rect 2566 4716 2567 4720
rect 2571 4716 2572 4720
rect 2566 4715 2572 4716
rect 2663 4719 2672 4720
rect 2663 4715 2664 4719
rect 2671 4715 2672 4719
rect 2702 4716 2703 4720
rect 2707 4716 2708 4720
rect 2702 4715 2708 4716
rect 2799 4719 2808 4720
rect 2799 4715 2800 4719
rect 2807 4715 2808 4719
rect 2838 4716 2839 4720
rect 2843 4716 2844 4720
rect 2838 4715 2844 4716
rect 2935 4719 2944 4720
rect 2935 4715 2936 4719
rect 2943 4715 2944 4719
rect 2974 4716 2975 4720
rect 2979 4716 2980 4720
rect 2974 4715 2980 4716
rect 3071 4719 3080 4720
rect 3071 4715 3072 4719
rect 3079 4715 3080 4719
rect 3110 4716 3111 4720
rect 3115 4716 3116 4720
rect 3110 4715 3116 4716
rect 3207 4719 3216 4720
rect 3207 4715 3208 4719
rect 3215 4715 3216 4719
rect 3246 4716 3247 4720
rect 3251 4716 3252 4720
rect 3246 4715 3252 4716
rect 3342 4719 3349 4720
rect 3342 4715 3343 4719
rect 3348 4715 3349 4719
rect 3398 4716 3399 4720
rect 3403 4716 3404 4720
rect 3398 4715 3404 4716
rect 3495 4719 3501 4720
rect 3495 4715 3496 4719
rect 3500 4718 3501 4719
rect 3503 4719 3509 4720
rect 3503 4718 3504 4719
rect 3500 4716 3504 4718
rect 3500 4715 3501 4716
rect 674 4714 680 4715
rect 2119 4714 2128 4715
rect 2255 4714 2264 4715
rect 2391 4714 2400 4715
rect 2527 4714 2536 4715
rect 2663 4714 2672 4715
rect 2799 4714 2808 4715
rect 2935 4714 2944 4715
rect 3071 4714 3080 4715
rect 3207 4714 3216 4715
rect 3342 4714 3349 4715
rect 3495 4714 3501 4715
rect 3503 4715 3504 4716
rect 3508 4715 3509 4719
rect 3542 4716 3543 4720
rect 3547 4716 3548 4720
rect 3542 4715 3548 4716
rect 3638 4719 3645 4720
rect 3638 4715 3639 4719
rect 3644 4715 3645 4719
rect 3678 4716 3679 4720
rect 3683 4716 3684 4720
rect 3678 4715 3684 4716
rect 3770 4719 3781 4720
rect 3770 4715 3771 4719
rect 3775 4715 3776 4719
rect 3780 4715 3781 4719
rect 3798 4717 3799 4721
rect 3803 4717 3804 4721
rect 3838 4720 3839 4724
rect 3843 4720 3844 4724
rect 4914 4721 4915 4725
rect 4919 4721 4920 4725
rect 4914 4720 4920 4721
rect 5058 4725 5064 4726
rect 5058 4721 5059 4725
rect 5063 4721 5064 4725
rect 5058 4720 5064 4721
rect 5210 4725 5216 4726
rect 5210 4721 5211 4725
rect 5215 4721 5216 4725
rect 5210 4720 5216 4721
rect 5370 4725 5376 4726
rect 5370 4721 5371 4725
rect 5375 4721 5376 4725
rect 5370 4720 5376 4721
rect 5514 4725 5520 4726
rect 5514 4721 5515 4725
rect 5519 4721 5520 4725
rect 5514 4720 5520 4721
rect 5662 4724 5668 4725
rect 5662 4720 5663 4724
rect 5667 4720 5668 4724
rect 3838 4719 3844 4720
rect 5662 4719 5668 4720
rect 3798 4716 3804 4717
rect 3503 4714 3509 4715
rect 3638 4714 3645 4715
rect 3770 4714 3781 4715
rect 1994 4705 2000 4706
rect 158 4704 164 4705
rect 294 4704 300 4705
rect 430 4704 436 4705
rect 566 4704 572 4705
rect 702 4704 708 4705
rect 1974 4704 1980 4705
rect 110 4703 116 4704
rect 110 4699 111 4703
rect 115 4699 116 4703
rect 158 4700 159 4704
rect 163 4700 164 4704
rect 158 4699 164 4700
rect 255 4703 261 4704
rect 255 4699 256 4703
rect 260 4702 261 4703
rect 274 4703 280 4704
rect 274 4702 275 4703
rect 260 4700 275 4702
rect 260 4699 261 4700
rect 110 4698 116 4699
rect 255 4698 261 4699
rect 274 4699 275 4700
rect 279 4699 280 4703
rect 294 4700 295 4704
rect 299 4700 300 4704
rect 294 4699 300 4700
rect 391 4703 397 4704
rect 391 4699 392 4703
rect 396 4702 397 4703
rect 410 4703 416 4704
rect 410 4702 411 4703
rect 396 4700 411 4702
rect 396 4699 397 4700
rect 274 4698 280 4699
rect 391 4698 397 4699
rect 410 4699 411 4700
rect 415 4699 416 4703
rect 430 4700 431 4704
rect 435 4700 436 4704
rect 430 4699 436 4700
rect 527 4703 533 4704
rect 527 4699 528 4703
rect 532 4702 533 4703
rect 546 4703 552 4704
rect 546 4702 547 4703
rect 532 4700 547 4702
rect 532 4699 533 4700
rect 410 4698 416 4699
rect 527 4698 533 4699
rect 546 4699 547 4700
rect 551 4699 552 4703
rect 566 4700 567 4704
rect 571 4700 572 4704
rect 566 4699 572 4700
rect 663 4703 669 4704
rect 663 4699 664 4703
rect 668 4702 669 4703
rect 682 4703 688 4704
rect 682 4702 683 4703
rect 668 4700 683 4702
rect 668 4699 669 4700
rect 546 4698 552 4699
rect 663 4698 669 4699
rect 682 4699 683 4700
rect 687 4699 688 4703
rect 702 4700 703 4704
rect 707 4700 708 4704
rect 702 4699 708 4700
rect 799 4703 808 4704
rect 799 4699 800 4703
rect 807 4699 808 4703
rect 682 4698 688 4699
rect 799 4698 808 4699
rect 1934 4703 1940 4704
rect 1934 4699 1935 4703
rect 1939 4699 1940 4703
rect 1974 4700 1975 4704
rect 1979 4700 1980 4704
rect 1994 4701 1995 4705
rect 1999 4701 2000 4705
rect 1994 4700 2000 4701
rect 2130 4705 2136 4706
rect 2130 4701 2131 4705
rect 2135 4701 2136 4705
rect 2130 4700 2136 4701
rect 2266 4705 2272 4706
rect 2266 4701 2267 4705
rect 2271 4701 2272 4705
rect 2266 4700 2272 4701
rect 2402 4705 2408 4706
rect 2402 4701 2403 4705
rect 2407 4701 2408 4705
rect 2402 4700 2408 4701
rect 2538 4705 2544 4706
rect 2538 4701 2539 4705
rect 2543 4701 2544 4705
rect 2538 4700 2544 4701
rect 2674 4705 2680 4706
rect 2674 4701 2675 4705
rect 2679 4701 2680 4705
rect 2674 4700 2680 4701
rect 2810 4705 2816 4706
rect 2810 4701 2811 4705
rect 2815 4701 2816 4705
rect 2810 4700 2816 4701
rect 2946 4705 2952 4706
rect 2946 4701 2947 4705
rect 2951 4701 2952 4705
rect 2946 4700 2952 4701
rect 3082 4705 3088 4706
rect 3082 4701 3083 4705
rect 3087 4701 3088 4705
rect 3082 4700 3088 4701
rect 3218 4705 3224 4706
rect 3218 4701 3219 4705
rect 3223 4701 3224 4705
rect 3218 4700 3224 4701
rect 3370 4705 3376 4706
rect 3370 4701 3371 4705
rect 3375 4701 3376 4705
rect 3370 4700 3376 4701
rect 3514 4705 3520 4706
rect 3514 4701 3515 4705
rect 3519 4701 3520 4705
rect 3514 4700 3520 4701
rect 3650 4705 3656 4706
rect 3650 4701 3651 4705
rect 3655 4701 3656 4705
rect 3650 4700 3656 4701
rect 3798 4704 3804 4705
rect 3798 4700 3799 4704
rect 3803 4700 3804 4704
rect 1974 4699 1980 4700
rect 3798 4699 3804 4700
rect 1934 4698 1940 4699
rect 5166 4675 5172 4676
rect 5166 4674 5167 4675
rect 5012 4666 5014 4673
rect 5157 4672 5167 4674
rect 5166 4671 5167 4672
rect 5171 4671 5172 4675
rect 5166 4670 5172 4671
rect 5199 4675 5205 4676
rect 5199 4671 5200 4675
rect 5204 4674 5205 4675
rect 5462 4675 5468 4676
rect 5204 4672 5217 4674
rect 5204 4671 5205 4672
rect 5199 4670 5205 4671
rect 5462 4671 5463 4675
rect 5467 4671 5468 4675
rect 5638 4675 5644 4676
rect 5638 4674 5639 4675
rect 5613 4672 5639 4674
rect 5462 4670 5468 4671
rect 5638 4671 5639 4672
rect 5643 4671 5644 4675
rect 5638 4670 5644 4671
rect 5490 4667 5496 4668
rect 5490 4666 5491 4667
rect 5012 4664 5491 4666
rect 5490 4663 5491 4664
rect 5495 4663 5496 4667
rect 5490 4662 5496 4663
rect 2122 4655 2128 4656
rect 2092 4646 2094 4653
rect 2122 4651 2123 4655
rect 2127 4654 2128 4655
rect 2258 4655 2264 4656
rect 2127 4652 2137 4654
rect 2127 4651 2128 4652
rect 2122 4650 2128 4651
rect 2258 4651 2259 4655
rect 2263 4654 2264 4655
rect 2394 4655 2400 4656
rect 2263 4652 2273 4654
rect 2263 4651 2264 4652
rect 2258 4650 2264 4651
rect 2394 4651 2395 4655
rect 2399 4654 2400 4655
rect 2530 4655 2536 4656
rect 2399 4652 2409 4654
rect 2399 4651 2400 4652
rect 2394 4650 2400 4651
rect 2530 4651 2531 4655
rect 2535 4654 2536 4655
rect 2666 4655 2672 4656
rect 2535 4652 2545 4654
rect 2535 4651 2536 4652
rect 2530 4650 2536 4651
rect 2666 4651 2667 4655
rect 2671 4654 2672 4655
rect 2802 4655 2808 4656
rect 2671 4652 2681 4654
rect 2671 4651 2672 4652
rect 2666 4650 2672 4651
rect 2802 4651 2803 4655
rect 2807 4654 2808 4655
rect 2938 4655 2944 4656
rect 2807 4652 2817 4654
rect 2807 4651 2808 4652
rect 2802 4650 2808 4651
rect 2938 4651 2939 4655
rect 2943 4654 2944 4655
rect 3074 4655 3080 4656
rect 2943 4652 2953 4654
rect 2943 4651 2944 4652
rect 2938 4650 2944 4651
rect 3074 4651 3075 4655
rect 3079 4654 3080 4655
rect 3210 4655 3216 4656
rect 3079 4652 3089 4654
rect 3079 4651 3080 4652
rect 3074 4650 3080 4651
rect 3210 4651 3211 4655
rect 3215 4654 3216 4655
rect 3503 4655 3509 4656
rect 3215 4652 3225 4654
rect 3215 4651 3216 4652
rect 3210 4650 3216 4651
rect 2442 4647 2448 4648
rect 2442 4646 2443 4647
rect 2092 4644 2443 4646
rect 2442 4643 2443 4644
rect 2447 4643 2448 4647
rect 3468 4646 3470 4653
rect 3503 4651 3504 4655
rect 3508 4654 3509 4655
rect 3982 4655 3988 4656
rect 3982 4654 3983 4655
rect 3508 4652 3521 4654
rect 3749 4652 3983 4654
rect 3508 4651 3509 4652
rect 3503 4650 3509 4651
rect 3982 4651 3983 4652
rect 3987 4651 3988 4655
rect 3982 4650 3988 4651
rect 3770 4647 3776 4648
rect 3770 4646 3771 4647
rect 3468 4644 3771 4646
rect 2442 4642 2448 4643
rect 3770 4643 3771 4644
rect 3775 4643 3776 4647
rect 3770 4642 3776 4643
rect 110 4637 116 4638
rect 1934 4637 1940 4638
rect 110 4633 111 4637
rect 115 4633 116 4637
rect 110 4632 116 4633
rect 158 4636 164 4637
rect 294 4636 300 4637
rect 430 4636 436 4637
rect 566 4636 572 4637
rect 702 4636 708 4637
rect 158 4632 159 4636
rect 163 4632 164 4636
rect 158 4631 164 4632
rect 255 4635 261 4636
rect 255 4631 256 4635
rect 260 4634 261 4635
rect 263 4635 269 4636
rect 263 4634 264 4635
rect 260 4632 264 4634
rect 260 4631 261 4632
rect 255 4630 261 4631
rect 263 4631 264 4632
rect 268 4631 269 4635
rect 294 4632 295 4636
rect 299 4632 300 4636
rect 294 4631 300 4632
rect 391 4635 400 4636
rect 391 4631 392 4635
rect 399 4631 400 4635
rect 430 4632 431 4636
rect 435 4632 436 4636
rect 430 4631 436 4632
rect 527 4635 536 4636
rect 527 4631 528 4635
rect 535 4631 536 4635
rect 566 4632 567 4636
rect 571 4632 572 4636
rect 566 4631 572 4632
rect 663 4635 672 4636
rect 663 4631 664 4635
rect 671 4631 672 4635
rect 702 4632 703 4636
rect 707 4632 708 4636
rect 702 4631 708 4632
rect 794 4635 805 4636
rect 794 4631 795 4635
rect 799 4631 800 4635
rect 804 4631 805 4635
rect 1934 4633 1935 4637
rect 1939 4633 1940 4637
rect 1934 4632 1940 4633
rect 263 4630 269 4631
rect 391 4630 400 4631
rect 527 4630 536 4631
rect 663 4630 672 4631
rect 794 4630 805 4631
rect 130 4621 136 4622
rect 110 4620 116 4621
rect 110 4616 111 4620
rect 115 4616 116 4620
rect 130 4617 131 4621
rect 135 4617 136 4621
rect 130 4616 136 4617
rect 266 4621 272 4622
rect 266 4617 267 4621
rect 271 4617 272 4621
rect 266 4616 272 4617
rect 402 4621 408 4622
rect 402 4617 403 4621
rect 407 4617 408 4621
rect 402 4616 408 4617
rect 538 4621 544 4622
rect 538 4617 539 4621
rect 543 4617 544 4621
rect 538 4616 544 4617
rect 674 4621 680 4622
rect 674 4617 675 4621
rect 679 4617 680 4621
rect 674 4616 680 4617
rect 1934 4620 1940 4621
rect 1934 4616 1935 4620
rect 1939 4616 1940 4620
rect 5647 4619 5653 4620
rect 5647 4618 5648 4619
rect 5613 4616 5648 4618
rect 110 4615 116 4616
rect 1934 4615 1940 4616
rect 4866 4615 4872 4616
rect 4866 4611 4867 4615
rect 4871 4611 4872 4615
rect 4866 4610 4872 4611
rect 4962 4615 4968 4616
rect 4962 4611 4963 4615
rect 4967 4611 4968 4615
rect 4962 4610 4968 4611
rect 5154 4615 5160 4616
rect 5154 4611 5155 4615
rect 5159 4611 5160 4615
rect 5154 4610 5160 4611
rect 5346 4615 5352 4616
rect 5346 4611 5347 4615
rect 5351 4611 5352 4615
rect 5647 4615 5648 4616
rect 5652 4615 5653 4619
rect 5647 4614 5653 4615
rect 5346 4610 5352 4611
rect 2566 4591 2572 4592
rect 2566 4590 2567 4591
rect 2421 4588 2567 4590
rect 2566 4587 2567 4588
rect 2571 4587 2572 4591
rect 2566 4586 2572 4587
rect 2638 4591 2644 4592
rect 2638 4587 2639 4591
rect 2643 4587 2644 4591
rect 3066 4591 3072 4592
rect 3066 4590 3067 4591
rect 2925 4588 3067 4590
rect 2638 4586 2644 4587
rect 3066 4587 3067 4588
rect 3071 4587 3072 4591
rect 3303 4591 3309 4592
rect 3303 4590 3304 4591
rect 3173 4588 3304 4590
rect 3066 4586 3072 4587
rect 3303 4587 3304 4588
rect 3308 4587 3309 4591
rect 3466 4591 3472 4592
rect 3466 4590 3467 4591
rect 3413 4588 3467 4590
rect 3303 4586 3309 4587
rect 3466 4587 3467 4588
rect 3471 4587 3472 4591
rect 3466 4586 3472 4587
rect 3638 4591 3644 4592
rect 3638 4587 3639 4591
rect 3643 4587 3644 4591
rect 3638 4586 3644 4587
rect 263 4571 269 4572
rect 228 4562 230 4569
rect 263 4567 264 4571
rect 268 4570 269 4571
rect 394 4571 400 4572
rect 268 4568 273 4570
rect 268 4567 269 4568
rect 263 4566 269 4567
rect 394 4567 395 4571
rect 399 4570 400 4571
rect 530 4571 536 4572
rect 399 4568 409 4570
rect 399 4567 400 4568
rect 394 4566 400 4567
rect 530 4567 531 4571
rect 535 4570 536 4571
rect 666 4571 672 4572
rect 535 4568 545 4570
rect 535 4567 536 4568
rect 530 4566 536 4567
rect 666 4567 667 4571
rect 671 4570 672 4571
rect 671 4568 681 4570
rect 3838 4568 3844 4569
rect 5662 4568 5668 4569
rect 671 4567 672 4568
rect 666 4566 672 4567
rect 3838 4564 3839 4568
rect 3843 4564 3844 4568
rect 802 4563 808 4564
rect 3838 4563 3844 4564
rect 4770 4567 4776 4568
rect 4770 4563 4771 4567
rect 4775 4563 4776 4567
rect 802 4562 803 4563
rect 228 4560 803 4562
rect 802 4559 803 4560
rect 807 4559 808 4563
rect 4770 4562 4776 4563
rect 4954 4567 4960 4568
rect 4954 4563 4955 4567
rect 4959 4563 4960 4567
rect 4954 4562 4960 4563
rect 5146 4567 5152 4568
rect 5146 4563 5147 4567
rect 5151 4563 5152 4567
rect 5146 4562 5152 4563
rect 5338 4567 5344 4568
rect 5338 4563 5339 4567
rect 5343 4563 5344 4567
rect 5338 4562 5344 4563
rect 5514 4567 5520 4568
rect 5514 4563 5515 4567
rect 5519 4563 5520 4567
rect 5662 4564 5663 4568
rect 5667 4564 5668 4568
rect 5662 4563 5668 4564
rect 5514 4562 5520 4563
rect 802 4558 808 4559
rect 4798 4552 4804 4553
rect 4982 4552 4988 4553
rect 5174 4552 5180 4553
rect 5366 4552 5372 4553
rect 5542 4552 5548 4553
rect 3838 4551 3844 4552
rect 3838 4547 3839 4551
rect 3843 4547 3844 4551
rect 4798 4548 4799 4552
rect 4803 4548 4804 4552
rect 4798 4547 4804 4548
rect 4895 4551 4901 4552
rect 4895 4547 4896 4551
rect 4900 4550 4901 4551
rect 4962 4551 4968 4552
rect 4962 4550 4963 4551
rect 4900 4548 4963 4550
rect 4900 4547 4901 4548
rect 3838 4546 3844 4547
rect 4895 4546 4901 4547
rect 4962 4547 4963 4548
rect 4967 4547 4968 4551
rect 4982 4548 4983 4552
rect 4987 4548 4988 4552
rect 4982 4547 4988 4548
rect 5079 4551 5085 4552
rect 5079 4547 5080 4551
rect 5084 4550 5085 4551
rect 5154 4551 5160 4552
rect 5154 4550 5155 4551
rect 5084 4548 5155 4550
rect 5084 4547 5085 4548
rect 4962 4546 4968 4547
rect 5079 4546 5085 4547
rect 5154 4547 5155 4548
rect 5159 4547 5160 4551
rect 5174 4548 5175 4552
rect 5179 4548 5180 4552
rect 5174 4547 5180 4548
rect 5271 4551 5277 4552
rect 5271 4547 5272 4551
rect 5276 4550 5277 4551
rect 5346 4551 5352 4552
rect 5346 4550 5347 4551
rect 5276 4548 5347 4550
rect 5276 4547 5277 4548
rect 5154 4546 5160 4547
rect 5271 4546 5277 4547
rect 5346 4547 5347 4548
rect 5351 4547 5352 4551
rect 5366 4548 5367 4552
rect 5371 4548 5372 4552
rect 5366 4547 5372 4548
rect 5462 4551 5469 4552
rect 5462 4547 5463 4551
rect 5468 4547 5469 4551
rect 5542 4548 5543 4552
rect 5547 4548 5548 4552
rect 5542 4547 5548 4548
rect 5639 4551 5648 4552
rect 5639 4547 5640 4551
rect 5647 4547 5648 4551
rect 5346 4546 5352 4547
rect 5462 4546 5469 4547
rect 5639 4546 5648 4547
rect 5662 4551 5668 4552
rect 5662 4547 5663 4551
rect 5667 4547 5668 4551
rect 5662 4546 5668 4547
rect 1974 4540 1980 4541
rect 3798 4540 3804 4541
rect 1974 4536 1975 4540
rect 1979 4536 1980 4540
rect 794 4535 800 4536
rect 1974 4535 1980 4536
rect 2322 4539 2328 4540
rect 2322 4535 2323 4539
rect 2327 4535 2328 4539
rect 794 4534 795 4535
rect 516 4532 795 4534
rect 516 4530 518 4532
rect 794 4531 795 4532
rect 799 4531 800 4535
rect 2322 4534 2328 4535
rect 2578 4539 2584 4540
rect 2578 4535 2579 4539
rect 2583 4535 2584 4539
rect 2578 4534 2584 4535
rect 2826 4539 2832 4540
rect 2826 4535 2827 4539
rect 2831 4535 2832 4539
rect 2826 4534 2832 4535
rect 3074 4539 3080 4540
rect 3074 4535 3075 4539
rect 3079 4535 3080 4539
rect 3074 4534 3080 4535
rect 3314 4539 3320 4540
rect 3314 4535 3315 4539
rect 3319 4535 3320 4539
rect 3314 4534 3320 4535
rect 3562 4539 3568 4540
rect 3562 4535 3563 4539
rect 3567 4535 3568 4539
rect 3798 4536 3799 4540
rect 3803 4536 3804 4540
rect 3798 4535 3804 4536
rect 3562 4534 3568 4535
rect 794 4530 800 4531
rect 1418 4531 1424 4532
rect 1418 4530 1419 4531
rect 437 4528 518 4530
rect 1341 4528 1419 4530
rect 522 4527 528 4528
rect 522 4523 523 4527
rect 527 4523 528 4527
rect 522 4522 528 4523
rect 698 4527 704 4528
rect 698 4523 699 4527
rect 703 4523 704 4527
rect 698 4522 704 4523
rect 882 4527 888 4528
rect 882 4523 883 4527
rect 887 4523 888 4527
rect 882 4522 888 4523
rect 1066 4527 1072 4528
rect 1066 4523 1067 4527
rect 1071 4523 1072 4527
rect 1418 4527 1419 4528
rect 1423 4527 1424 4531
rect 2566 4531 2572 4532
rect 1418 4526 1424 4527
rect 1434 4527 1440 4528
rect 1066 4522 1072 4523
rect 1434 4523 1435 4527
rect 1439 4523 1440 4527
rect 1434 4522 1440 4523
rect 1626 4527 1632 4528
rect 1626 4523 1627 4527
rect 1631 4523 1632 4527
rect 1626 4522 1632 4523
rect 1794 4527 1800 4528
rect 1794 4523 1795 4527
rect 1799 4523 1800 4527
rect 2566 4527 2567 4531
rect 2571 4530 2572 4531
rect 3066 4531 3072 4532
rect 2571 4528 2706 4530
rect 2571 4527 2572 4528
rect 2566 4526 2572 4527
rect 2350 4524 2356 4525
rect 2606 4524 2612 4525
rect 2704 4524 2706 4528
rect 3066 4527 3067 4531
rect 3071 4530 3072 4531
rect 3303 4531 3309 4532
rect 3071 4528 3202 4530
rect 3071 4527 3072 4528
rect 3066 4526 3072 4527
rect 3200 4526 3202 4528
rect 3303 4527 3304 4531
rect 3308 4530 3309 4531
rect 3466 4531 3472 4532
rect 3308 4528 3442 4530
rect 3308 4527 3309 4528
rect 3303 4526 3309 4527
rect 3440 4526 3442 4528
rect 3466 4527 3467 4531
rect 3471 4530 3472 4531
rect 3471 4528 3690 4530
rect 3471 4527 3472 4528
rect 3466 4526 3472 4527
rect 3688 4526 3690 4528
rect 3199 4525 3205 4526
rect 3439 4525 3445 4526
rect 3687 4525 3693 4526
rect 2854 4524 2860 4525
rect 3102 4524 3108 4525
rect 1794 4522 1800 4523
rect 1974 4523 1980 4524
rect 1974 4519 1975 4523
rect 1979 4519 1980 4523
rect 2350 4520 2351 4524
rect 2355 4520 2356 4524
rect 2350 4519 2356 4520
rect 2442 4523 2453 4524
rect 2442 4519 2443 4523
rect 2447 4519 2448 4523
rect 2452 4519 2453 4523
rect 2606 4520 2607 4524
rect 2611 4520 2612 4524
rect 2606 4519 2612 4520
rect 2703 4523 2709 4524
rect 2703 4519 2704 4523
rect 2708 4519 2709 4523
rect 2854 4520 2855 4524
rect 2859 4520 2860 4524
rect 2854 4519 2860 4520
rect 2950 4523 2957 4524
rect 2950 4519 2951 4523
rect 2956 4519 2957 4523
rect 3102 4520 3103 4524
rect 3107 4520 3108 4524
rect 3199 4521 3200 4525
rect 3204 4521 3205 4525
rect 3199 4520 3205 4521
rect 3342 4524 3348 4525
rect 3342 4520 3343 4524
rect 3347 4520 3348 4524
rect 3439 4521 3440 4525
rect 3444 4521 3445 4525
rect 3439 4520 3445 4521
rect 3590 4524 3596 4525
rect 3590 4520 3591 4524
rect 3595 4520 3596 4524
rect 3687 4521 3688 4525
rect 3692 4521 3693 4525
rect 3687 4520 3693 4521
rect 3798 4523 3804 4524
rect 3102 4519 3108 4520
rect 3342 4519 3348 4520
rect 3590 4519 3596 4520
rect 3798 4519 3799 4523
rect 3803 4519 3804 4523
rect 1974 4518 1980 4519
rect 2442 4518 2453 4519
rect 2703 4518 2709 4519
rect 2950 4518 2957 4519
rect 3798 4518 3804 4519
rect 3838 4481 3844 4482
rect 5662 4481 5668 4482
rect 110 4480 116 4481
rect 1934 4480 1940 4481
rect 110 4476 111 4480
rect 115 4476 116 4480
rect 110 4475 116 4476
rect 338 4479 344 4480
rect 338 4475 339 4479
rect 343 4475 344 4479
rect 338 4474 344 4475
rect 514 4479 520 4480
rect 514 4475 515 4479
rect 519 4475 520 4479
rect 514 4474 520 4475
rect 690 4479 696 4480
rect 690 4475 691 4479
rect 695 4475 696 4479
rect 690 4474 696 4475
rect 874 4479 880 4480
rect 874 4475 875 4479
rect 879 4475 880 4479
rect 874 4474 880 4475
rect 1058 4479 1064 4480
rect 1058 4475 1059 4479
rect 1063 4475 1064 4479
rect 1058 4474 1064 4475
rect 1242 4479 1248 4480
rect 1242 4475 1243 4479
rect 1247 4475 1248 4479
rect 1242 4474 1248 4475
rect 1426 4479 1432 4480
rect 1426 4475 1427 4479
rect 1431 4475 1432 4479
rect 1426 4474 1432 4475
rect 1618 4479 1624 4480
rect 1618 4475 1619 4479
rect 1623 4475 1624 4479
rect 1618 4474 1624 4475
rect 1786 4479 1792 4480
rect 1786 4475 1787 4479
rect 1791 4475 1792 4479
rect 1934 4476 1935 4480
rect 1939 4476 1940 4480
rect 3838 4477 3839 4481
rect 3843 4477 3844 4481
rect 3838 4476 3844 4477
rect 4486 4480 4492 4481
rect 4670 4480 4676 4481
rect 4878 4480 4884 4481
rect 5094 4480 5100 4481
rect 5326 4480 5332 4481
rect 5542 4480 5548 4481
rect 4486 4476 4487 4480
rect 4491 4476 4492 4480
rect 1934 4475 1940 4476
rect 4486 4475 4492 4476
rect 4583 4479 4589 4480
rect 4583 4475 4584 4479
rect 4588 4478 4589 4479
rect 4607 4479 4613 4480
rect 4607 4478 4608 4479
rect 4588 4476 4608 4478
rect 4588 4475 4589 4476
rect 1786 4474 1792 4475
rect 4583 4474 4589 4475
rect 4607 4475 4608 4476
rect 4612 4475 4613 4479
rect 4670 4476 4671 4480
rect 4675 4476 4676 4480
rect 4670 4475 4676 4476
rect 4767 4479 4773 4480
rect 4767 4475 4768 4479
rect 4772 4478 4773 4479
rect 4791 4479 4797 4480
rect 4791 4478 4792 4479
rect 4772 4476 4792 4478
rect 4772 4475 4773 4476
rect 4607 4474 4613 4475
rect 4767 4474 4773 4475
rect 4791 4475 4792 4476
rect 4796 4475 4797 4479
rect 4878 4476 4879 4480
rect 4883 4476 4884 4480
rect 4878 4475 4884 4476
rect 4975 4479 4984 4480
rect 4975 4475 4976 4479
rect 4983 4475 4984 4479
rect 5094 4476 5095 4480
rect 5099 4476 5100 4480
rect 5094 4475 5100 4476
rect 5191 4479 5197 4480
rect 5191 4475 5192 4479
rect 5196 4478 5197 4479
rect 5207 4479 5213 4480
rect 5207 4478 5208 4479
rect 5196 4476 5208 4478
rect 5196 4475 5197 4476
rect 4791 4474 4797 4475
rect 4975 4474 4984 4475
rect 5191 4474 5197 4475
rect 5207 4475 5208 4476
rect 5212 4475 5213 4479
rect 5326 4476 5327 4480
rect 5331 4476 5332 4480
rect 5326 4475 5332 4476
rect 5422 4479 5429 4480
rect 5422 4475 5423 4479
rect 5428 4475 5429 4479
rect 5542 4476 5543 4480
rect 5547 4476 5548 4480
rect 5542 4475 5548 4476
rect 5634 4479 5645 4480
rect 5634 4475 5635 4479
rect 5639 4475 5640 4479
rect 5644 4475 5645 4479
rect 5662 4477 5663 4481
rect 5667 4477 5668 4481
rect 5662 4476 5668 4477
rect 5207 4474 5213 4475
rect 5422 4474 5429 4475
rect 5634 4474 5645 4475
rect 4458 4465 4464 4466
rect 366 4464 372 4465
rect 542 4464 548 4465
rect 718 4464 724 4465
rect 902 4464 908 4465
rect 1086 4464 1092 4465
rect 1270 4464 1276 4465
rect 1454 4464 1460 4465
rect 1646 4464 1652 4465
rect 1814 4464 1820 4465
rect 3838 4464 3844 4465
rect 110 4463 116 4464
rect 110 4459 111 4463
rect 115 4459 116 4463
rect 366 4460 367 4464
rect 371 4460 372 4464
rect 366 4459 372 4460
rect 463 4463 469 4464
rect 463 4459 464 4463
rect 468 4462 469 4463
rect 522 4463 528 4464
rect 522 4462 523 4463
rect 468 4460 523 4462
rect 468 4459 469 4460
rect 110 4458 116 4459
rect 463 4458 469 4459
rect 522 4459 523 4460
rect 527 4459 528 4463
rect 542 4460 543 4464
rect 547 4460 548 4464
rect 542 4459 548 4460
rect 639 4463 645 4464
rect 639 4459 640 4463
rect 644 4462 645 4463
rect 698 4463 704 4464
rect 698 4462 699 4463
rect 644 4460 699 4462
rect 644 4459 645 4460
rect 522 4458 528 4459
rect 639 4458 645 4459
rect 698 4459 699 4460
rect 703 4459 704 4463
rect 718 4460 719 4464
rect 723 4460 724 4464
rect 718 4459 724 4460
rect 815 4463 821 4464
rect 815 4459 816 4463
rect 820 4462 821 4463
rect 882 4463 888 4464
rect 882 4462 883 4463
rect 820 4460 883 4462
rect 820 4459 821 4460
rect 698 4458 704 4459
rect 815 4458 821 4459
rect 882 4459 883 4460
rect 887 4459 888 4463
rect 902 4460 903 4464
rect 907 4460 908 4464
rect 902 4459 908 4460
rect 999 4463 1005 4464
rect 999 4459 1000 4463
rect 1004 4462 1005 4463
rect 1066 4463 1072 4464
rect 1066 4462 1067 4463
rect 1004 4460 1067 4462
rect 1004 4459 1005 4460
rect 882 4458 888 4459
rect 999 4458 1005 4459
rect 1066 4459 1067 4460
rect 1071 4459 1072 4463
rect 1086 4460 1087 4464
rect 1091 4460 1092 4464
rect 1086 4459 1092 4460
rect 1178 4463 1189 4464
rect 1178 4459 1179 4463
rect 1183 4459 1184 4463
rect 1188 4459 1189 4463
rect 1270 4460 1271 4464
rect 1275 4460 1276 4464
rect 1270 4459 1276 4460
rect 1367 4463 1373 4464
rect 1367 4459 1368 4463
rect 1372 4462 1373 4463
rect 1434 4463 1440 4464
rect 1434 4462 1435 4463
rect 1372 4460 1435 4462
rect 1372 4459 1373 4460
rect 1066 4458 1072 4459
rect 1178 4458 1189 4459
rect 1367 4458 1373 4459
rect 1434 4459 1435 4460
rect 1439 4459 1440 4463
rect 1454 4460 1455 4464
rect 1459 4460 1460 4464
rect 1454 4459 1460 4460
rect 1551 4463 1557 4464
rect 1551 4459 1552 4463
rect 1556 4462 1557 4463
rect 1626 4463 1632 4464
rect 1626 4462 1627 4463
rect 1556 4460 1627 4462
rect 1556 4459 1557 4460
rect 1434 4458 1440 4459
rect 1551 4458 1557 4459
rect 1626 4459 1627 4460
rect 1631 4459 1632 4463
rect 1646 4460 1647 4464
rect 1651 4460 1652 4464
rect 1646 4459 1652 4460
rect 1743 4463 1749 4464
rect 1743 4459 1744 4463
rect 1748 4462 1749 4463
rect 1794 4463 1800 4464
rect 1794 4462 1795 4463
rect 1748 4460 1795 4462
rect 1748 4459 1749 4460
rect 1626 4458 1632 4459
rect 1743 4458 1749 4459
rect 1794 4459 1795 4460
rect 1799 4459 1800 4463
rect 1814 4460 1815 4464
rect 1819 4460 1820 4464
rect 1814 4459 1820 4460
rect 1910 4463 1917 4464
rect 1910 4459 1911 4463
rect 1916 4459 1917 4463
rect 1794 4458 1800 4459
rect 1910 4458 1917 4459
rect 1934 4463 1940 4464
rect 1934 4459 1935 4463
rect 1939 4459 1940 4463
rect 3838 4460 3839 4464
rect 3843 4460 3844 4464
rect 4458 4461 4459 4465
rect 4463 4461 4464 4465
rect 4458 4460 4464 4461
rect 4642 4465 4648 4466
rect 4642 4461 4643 4465
rect 4647 4461 4648 4465
rect 4642 4460 4648 4461
rect 4850 4465 4856 4466
rect 4850 4461 4851 4465
rect 4855 4461 4856 4465
rect 4850 4460 4856 4461
rect 5066 4465 5072 4466
rect 5066 4461 5067 4465
rect 5071 4461 5072 4465
rect 5066 4460 5072 4461
rect 5298 4465 5304 4466
rect 5298 4461 5299 4465
rect 5303 4461 5304 4465
rect 5298 4460 5304 4461
rect 5514 4465 5520 4466
rect 5514 4461 5515 4465
rect 5519 4461 5520 4465
rect 5514 4460 5520 4461
rect 5662 4464 5668 4465
rect 5662 4460 5663 4464
rect 5667 4460 5668 4464
rect 3838 4459 3844 4460
rect 5662 4459 5668 4460
rect 1934 4458 1940 4459
rect 1974 4457 1980 4458
rect 3798 4457 3804 4458
rect 1974 4453 1975 4457
rect 1979 4453 1980 4457
rect 1974 4452 1980 4453
rect 2542 4456 2548 4457
rect 2782 4456 2788 4457
rect 3014 4456 3020 4457
rect 3246 4456 3252 4457
rect 3470 4456 3476 4457
rect 3678 4456 3684 4457
rect 2542 4452 2543 4456
rect 2547 4452 2548 4456
rect 2542 4451 2548 4452
rect 2638 4455 2645 4456
rect 2638 4451 2639 4455
rect 2644 4451 2645 4455
rect 2782 4452 2783 4456
rect 2787 4452 2788 4456
rect 2782 4451 2788 4452
rect 2879 4455 2885 4456
rect 2879 4451 2880 4455
rect 2884 4454 2885 4455
rect 2895 4455 2901 4456
rect 2895 4454 2896 4455
rect 2884 4452 2896 4454
rect 2884 4451 2885 4452
rect 2638 4450 2645 4451
rect 2879 4450 2885 4451
rect 2895 4451 2896 4452
rect 2900 4451 2901 4455
rect 3014 4452 3015 4456
rect 3019 4452 3020 4456
rect 3014 4451 3020 4452
rect 3111 4455 3117 4456
rect 3111 4451 3112 4455
rect 3116 4454 3117 4455
rect 3126 4455 3132 4456
rect 3126 4454 3127 4455
rect 3116 4452 3127 4454
rect 3116 4451 3117 4452
rect 2895 4450 2901 4451
rect 3111 4450 3117 4451
rect 3126 4451 3127 4452
rect 3131 4451 3132 4455
rect 3246 4452 3247 4456
rect 3251 4452 3252 4456
rect 3246 4451 3252 4452
rect 3343 4455 3352 4456
rect 3343 4451 3344 4455
rect 3351 4451 3352 4455
rect 3470 4452 3471 4456
rect 3475 4452 3476 4456
rect 3470 4451 3476 4452
rect 3567 4455 3576 4456
rect 3567 4451 3568 4455
rect 3575 4451 3576 4455
rect 3678 4452 3679 4456
rect 3683 4452 3684 4456
rect 3678 4451 3684 4452
rect 3770 4455 3781 4456
rect 3770 4451 3771 4455
rect 3775 4451 3776 4455
rect 3780 4451 3781 4455
rect 3798 4453 3799 4457
rect 3803 4453 3804 4457
rect 3798 4452 3804 4453
rect 3126 4450 3132 4451
rect 3343 4450 3352 4451
rect 3567 4450 3576 4451
rect 3770 4450 3781 4451
rect 2514 4441 2520 4442
rect 1974 4440 1980 4441
rect 1974 4436 1975 4440
rect 1979 4436 1980 4440
rect 2514 4437 2515 4441
rect 2519 4437 2520 4441
rect 2514 4436 2520 4437
rect 2754 4441 2760 4442
rect 2754 4437 2755 4441
rect 2759 4437 2760 4441
rect 2754 4436 2760 4437
rect 2986 4441 2992 4442
rect 2986 4437 2987 4441
rect 2991 4437 2992 4441
rect 2986 4436 2992 4437
rect 3218 4441 3224 4442
rect 3218 4437 3219 4441
rect 3223 4437 3224 4441
rect 3218 4436 3224 4437
rect 3442 4441 3448 4442
rect 3442 4437 3443 4441
rect 3447 4437 3448 4441
rect 3442 4436 3448 4437
rect 3650 4441 3656 4442
rect 3650 4437 3651 4441
rect 3655 4437 3656 4441
rect 3650 4436 3656 4437
rect 3798 4440 3804 4441
rect 3798 4436 3799 4440
rect 3803 4436 3804 4440
rect 1974 4435 1980 4436
rect 3798 4435 3804 4436
rect 4550 4415 4556 4416
rect 4550 4411 4551 4415
rect 4555 4411 4556 4415
rect 4550 4410 4556 4411
rect 4607 4415 4613 4416
rect 4607 4411 4608 4415
rect 4612 4414 4613 4415
rect 4791 4415 4797 4416
rect 4612 4412 4649 4414
rect 4612 4411 4613 4412
rect 4607 4410 4613 4411
rect 4791 4411 4792 4415
rect 4796 4414 4797 4415
rect 4978 4415 4984 4416
rect 4796 4412 4857 4414
rect 4796 4411 4797 4412
rect 4791 4410 4797 4411
rect 4978 4411 4979 4415
rect 4983 4414 4984 4415
rect 5207 4415 5213 4416
rect 4983 4412 5073 4414
rect 4983 4411 4984 4412
rect 4978 4410 4984 4411
rect 5207 4411 5208 4415
rect 5212 4414 5213 4415
rect 5642 4415 5648 4416
rect 5642 4414 5643 4415
rect 5212 4412 5305 4414
rect 5613 4412 5643 4414
rect 5212 4411 5213 4412
rect 5207 4410 5213 4411
rect 5642 4411 5643 4412
rect 5647 4411 5648 4415
rect 5642 4410 5648 4411
rect 110 4405 116 4406
rect 1934 4405 1940 4406
rect 110 4401 111 4405
rect 115 4401 116 4405
rect 110 4400 116 4401
rect 566 4404 572 4405
rect 710 4404 716 4405
rect 862 4404 868 4405
rect 1022 4404 1028 4405
rect 1182 4404 1188 4405
rect 1342 4404 1348 4405
rect 1502 4404 1508 4405
rect 1670 4404 1676 4405
rect 1814 4404 1820 4405
rect 566 4400 567 4404
rect 571 4400 572 4404
rect 566 4399 572 4400
rect 663 4403 672 4404
rect 663 4399 664 4403
rect 671 4399 672 4403
rect 710 4400 711 4404
rect 715 4400 716 4404
rect 710 4399 716 4400
rect 807 4403 813 4404
rect 807 4399 808 4403
rect 812 4402 813 4403
rect 823 4403 829 4404
rect 823 4402 824 4403
rect 812 4400 824 4402
rect 812 4399 813 4400
rect 663 4398 672 4399
rect 807 4398 813 4399
rect 823 4399 824 4400
rect 828 4399 829 4403
rect 862 4400 863 4404
rect 867 4400 868 4404
rect 862 4399 868 4400
rect 959 4403 968 4404
rect 959 4399 960 4403
rect 967 4399 968 4403
rect 1022 4400 1023 4404
rect 1027 4400 1028 4404
rect 1022 4399 1028 4400
rect 1119 4403 1128 4404
rect 1119 4399 1120 4403
rect 1127 4399 1128 4403
rect 1182 4400 1183 4404
rect 1187 4400 1188 4404
rect 1182 4399 1188 4400
rect 1278 4403 1285 4404
rect 1278 4399 1279 4403
rect 1284 4399 1285 4403
rect 1342 4400 1343 4404
rect 1347 4400 1348 4404
rect 1342 4399 1348 4400
rect 1434 4403 1445 4404
rect 1434 4399 1435 4403
rect 1439 4399 1440 4403
rect 1444 4399 1445 4403
rect 1502 4400 1503 4404
rect 1507 4400 1508 4404
rect 1502 4399 1508 4400
rect 1594 4403 1605 4404
rect 1594 4399 1595 4403
rect 1599 4399 1600 4403
rect 1604 4399 1605 4403
rect 1670 4400 1671 4404
rect 1675 4400 1676 4404
rect 1670 4399 1676 4400
rect 1767 4403 1776 4404
rect 1767 4399 1768 4403
rect 1775 4399 1776 4403
rect 1814 4400 1815 4404
rect 1819 4400 1820 4404
rect 1814 4399 1820 4400
rect 1911 4403 1917 4404
rect 1911 4399 1912 4403
rect 1916 4402 1917 4403
rect 1926 4403 1932 4404
rect 1926 4402 1927 4403
rect 1916 4400 1927 4402
rect 1916 4399 1917 4400
rect 823 4398 829 4399
rect 959 4398 968 4399
rect 1119 4398 1128 4399
rect 1278 4398 1285 4399
rect 1434 4398 1445 4399
rect 1594 4398 1605 4399
rect 1767 4398 1776 4399
rect 1911 4398 1917 4399
rect 1926 4399 1927 4400
rect 1931 4399 1932 4403
rect 1934 4401 1935 4405
rect 1939 4401 1940 4405
rect 1934 4400 1940 4401
rect 1926 4398 1932 4399
rect 2950 4399 2956 4400
rect 2950 4398 2951 4399
rect 2852 4396 2951 4398
rect 538 4389 544 4390
rect 110 4388 116 4389
rect 110 4384 111 4388
rect 115 4384 116 4388
rect 538 4385 539 4389
rect 543 4385 544 4389
rect 538 4384 544 4385
rect 682 4389 688 4390
rect 682 4385 683 4389
rect 687 4385 688 4389
rect 682 4384 688 4385
rect 834 4389 840 4390
rect 834 4385 835 4389
rect 839 4385 840 4389
rect 834 4384 840 4385
rect 994 4389 1000 4390
rect 994 4385 995 4389
rect 999 4385 1000 4389
rect 994 4384 1000 4385
rect 1154 4389 1160 4390
rect 1154 4385 1155 4389
rect 1159 4385 1160 4389
rect 1154 4384 1160 4385
rect 1314 4389 1320 4390
rect 1314 4385 1315 4389
rect 1319 4385 1320 4389
rect 1314 4384 1320 4385
rect 1474 4389 1480 4390
rect 1474 4385 1475 4389
rect 1479 4385 1480 4389
rect 1474 4384 1480 4385
rect 1642 4389 1648 4390
rect 1642 4385 1643 4389
rect 1647 4385 1648 4389
rect 1642 4384 1648 4385
rect 1786 4389 1792 4390
rect 2852 4389 2854 4396
rect 2950 4395 2951 4396
rect 2955 4395 2956 4399
rect 2950 4394 2956 4395
rect 2895 4391 2901 4392
rect 1786 4385 1787 4389
rect 1791 4385 1792 4389
rect 1786 4384 1792 4385
rect 1934 4388 1940 4389
rect 1934 4384 1935 4388
rect 1939 4384 1940 4388
rect 110 4383 116 4384
rect 1934 4383 1940 4384
rect 2612 4382 2614 4389
rect 2895 4387 2896 4391
rect 2900 4390 2901 4391
rect 3126 4391 3132 4392
rect 2900 4388 2993 4390
rect 2900 4387 2901 4388
rect 2895 4386 2901 4387
rect 3126 4387 3127 4391
rect 3131 4390 3132 4391
rect 3346 4391 3352 4392
rect 3131 4388 3225 4390
rect 3131 4387 3132 4388
rect 3126 4386 3132 4387
rect 3346 4387 3347 4391
rect 3351 4390 3352 4391
rect 3570 4391 3576 4392
rect 3351 4388 3449 4390
rect 3351 4387 3352 4388
rect 3346 4386 3352 4387
rect 3570 4387 3571 4391
rect 3575 4390 3576 4391
rect 3575 4388 3657 4390
rect 3575 4387 3576 4388
rect 3570 4386 3576 4387
rect 2926 4383 2932 4384
rect 2926 4382 2927 4383
rect 2612 4380 2927 4382
rect 2926 4379 2927 4380
rect 2931 4379 2932 4383
rect 2926 4378 2932 4379
rect 3778 4359 3784 4360
rect 3778 4355 3779 4359
rect 3783 4358 3784 4359
rect 5634 4359 5640 4360
rect 5634 4358 5635 4359
rect 3783 4356 3865 4358
rect 5613 4356 5635 4358
rect 3783 4355 3784 4356
rect 3778 4354 3784 4355
rect 4002 4355 4008 4356
rect 3358 4351 3364 4352
rect 3358 4350 3359 4351
rect 3236 4348 3359 4350
rect 1926 4347 1932 4348
rect 1926 4343 1927 4347
rect 1931 4346 1932 4347
rect 3236 4346 3238 4348
rect 3358 4347 3359 4348
rect 3363 4347 3364 4351
rect 4002 4351 4003 4355
rect 4007 4351 4008 4355
rect 4002 4350 4008 4351
rect 4138 4355 4144 4356
rect 4138 4351 4139 4355
rect 4143 4351 4144 4355
rect 4138 4350 4144 4351
rect 4378 4355 4384 4356
rect 4378 4351 4379 4355
rect 4383 4351 4384 4355
rect 4378 4350 4384 4351
rect 4490 4355 4496 4356
rect 4490 4351 4491 4355
rect 4495 4351 4496 4355
rect 4490 4350 4496 4351
rect 4722 4355 4728 4356
rect 4722 4351 4723 4355
rect 4727 4351 4728 4355
rect 4722 4350 4728 4351
rect 4986 4355 4992 4356
rect 4986 4351 4987 4355
rect 4991 4351 4992 4355
rect 4986 4350 4992 4351
rect 5258 4355 5264 4356
rect 5258 4351 5259 4355
rect 5263 4351 5264 4355
rect 5634 4355 5635 4356
rect 5639 4355 5640 4359
rect 5634 4354 5640 4355
rect 5258 4350 5264 4351
rect 3358 4346 3364 4347
rect 3770 4347 3776 4348
rect 3770 4346 3771 4347
rect 1931 4344 2001 4346
rect 2901 4344 3238 4346
rect 3749 4344 3771 4346
rect 1931 4343 1932 4344
rect 1926 4342 1932 4343
rect 2386 4343 2392 4344
rect 666 4339 672 4340
rect 636 4330 638 4337
rect 666 4335 667 4339
rect 671 4338 672 4339
rect 823 4339 829 4340
rect 671 4336 689 4338
rect 671 4335 672 4336
rect 666 4334 672 4335
rect 823 4335 824 4339
rect 828 4338 829 4339
rect 962 4339 968 4340
rect 828 4336 841 4338
rect 828 4335 829 4336
rect 823 4334 829 4335
rect 962 4335 963 4339
rect 967 4338 968 4339
rect 1122 4339 1128 4340
rect 967 4336 1001 4338
rect 967 4335 968 4336
rect 962 4334 968 4335
rect 1122 4335 1123 4339
rect 1127 4338 1128 4339
rect 1542 4339 1548 4340
rect 1127 4336 1161 4338
rect 1413 4336 1461 4338
rect 1127 4335 1128 4336
rect 1122 4334 1128 4335
rect 1174 4331 1180 4332
rect 1174 4330 1175 4331
rect 636 4328 1175 4330
rect 1174 4327 1175 4328
rect 1179 4327 1180 4331
rect 1459 4330 1461 4336
rect 1542 4335 1543 4339
rect 1547 4335 1548 4339
rect 1770 4339 1776 4340
rect 1542 4334 1548 4335
rect 1594 4331 1600 4332
rect 1594 4330 1595 4331
rect 1459 4328 1595 4330
rect 1174 4326 1180 4327
rect 1594 4327 1595 4328
rect 1599 4327 1600 4331
rect 1740 4330 1742 4337
rect 1770 4335 1771 4339
rect 1775 4338 1776 4339
rect 2386 4339 2387 4343
rect 2391 4339 2392 4343
rect 2386 4338 2392 4339
rect 3242 4343 3248 4344
rect 3242 4339 3243 4343
rect 3247 4339 3248 4343
rect 3770 4343 3771 4344
rect 3775 4343 3776 4347
rect 3770 4342 3776 4343
rect 3242 4338 3248 4339
rect 1775 4336 1793 4338
rect 1775 4335 1776 4336
rect 1770 4334 1776 4335
rect 1910 4331 1916 4332
rect 1910 4330 1911 4331
rect 1740 4328 1911 4330
rect 1594 4326 1600 4327
rect 1910 4327 1911 4328
rect 1915 4327 1916 4331
rect 1910 4326 1916 4327
rect 3838 4308 3844 4309
rect 5662 4308 5668 4309
rect 3838 4304 3839 4308
rect 3843 4304 3844 4308
rect 3838 4303 3844 4304
rect 3858 4307 3864 4308
rect 3858 4303 3859 4307
rect 3863 4303 3864 4307
rect 3858 4302 3864 4303
rect 3994 4307 4000 4308
rect 3994 4303 3995 4307
rect 3999 4303 4000 4307
rect 3994 4302 4000 4303
rect 4130 4307 4136 4308
rect 4130 4303 4131 4307
rect 4135 4303 4136 4307
rect 4130 4302 4136 4303
rect 4282 4307 4288 4308
rect 4282 4303 4283 4307
rect 4287 4303 4288 4307
rect 4282 4302 4288 4303
rect 4482 4307 4488 4308
rect 4482 4303 4483 4307
rect 4487 4303 4488 4307
rect 4482 4302 4488 4303
rect 4714 4307 4720 4308
rect 4714 4303 4715 4307
rect 4719 4303 4720 4307
rect 4714 4302 4720 4303
rect 4978 4307 4984 4308
rect 4978 4303 4979 4307
rect 4983 4303 4984 4307
rect 4978 4302 4984 4303
rect 5250 4307 5256 4308
rect 5250 4303 5251 4307
rect 5255 4303 5256 4307
rect 5250 4302 5256 4303
rect 5514 4307 5520 4308
rect 5514 4303 5515 4307
rect 5519 4303 5520 4307
rect 5662 4304 5663 4308
rect 5667 4304 5668 4308
rect 5662 4303 5668 4304
rect 5514 4302 5520 4303
rect 1046 4299 1052 4300
rect 1046 4298 1047 4299
rect 772 4296 1047 4298
rect 772 4286 774 4296
rect 1046 4295 1047 4296
rect 1051 4295 1052 4299
rect 1046 4294 1052 4295
rect 1974 4296 1980 4297
rect 3798 4296 3804 4297
rect 1974 4292 1975 4296
rect 1979 4292 1980 4296
rect 1206 4291 1212 4292
rect 1206 4290 1207 4291
rect 1024 4288 1207 4290
rect 1024 4286 1026 4288
rect 1206 4287 1207 4288
rect 1211 4287 1212 4291
rect 1714 4291 1720 4292
rect 1974 4291 1980 4292
rect 1994 4295 2000 4296
rect 1994 4291 1995 4295
rect 1999 4291 2000 4295
rect 1714 4290 1715 4291
rect 1592 4288 1715 4290
rect 1206 4286 1212 4287
rect 1278 4287 1284 4288
rect 725 4284 774 4286
rect 1021 4284 1026 4286
rect 778 4283 784 4284
rect 778 4279 779 4283
rect 783 4279 784 4283
rect 1278 4283 1279 4287
rect 1283 4283 1284 4287
rect 1592 4286 1594 4288
rect 1714 4287 1715 4288
rect 1719 4287 1720 4291
rect 1994 4290 2000 4291
rect 2378 4295 2384 4296
rect 2378 4291 2379 4295
rect 2383 4291 2384 4295
rect 2378 4290 2384 4291
rect 2802 4295 2808 4296
rect 2802 4291 2803 4295
rect 2807 4291 2808 4295
rect 2802 4290 2808 4291
rect 3234 4295 3240 4296
rect 3234 4291 3235 4295
rect 3239 4291 3240 4295
rect 3234 4290 3240 4291
rect 3650 4295 3656 4296
rect 3650 4291 3651 4295
rect 3655 4291 3656 4295
rect 3798 4292 3799 4296
rect 3803 4292 3804 4296
rect 3886 4292 3892 4293
rect 4022 4292 4028 4293
rect 4158 4292 4164 4293
rect 4310 4292 4316 4293
rect 4510 4292 4516 4293
rect 4742 4292 4748 4293
rect 5006 4292 5012 4293
rect 5278 4292 5284 4293
rect 5542 4292 5548 4293
rect 3798 4291 3804 4292
rect 3838 4291 3844 4292
rect 3650 4290 3656 4291
rect 1714 4286 1720 4287
rect 3838 4287 3839 4291
rect 3843 4287 3844 4291
rect 3886 4288 3887 4292
rect 3891 4288 3892 4292
rect 3886 4287 3892 4288
rect 3983 4291 3989 4292
rect 3983 4287 3984 4291
rect 3988 4290 3989 4291
rect 4002 4291 4008 4292
rect 4002 4290 4003 4291
rect 3988 4288 4003 4290
rect 3988 4287 3989 4288
rect 3838 4286 3844 4287
rect 3983 4286 3989 4287
rect 4002 4287 4003 4288
rect 4007 4287 4008 4291
rect 4022 4288 4023 4292
rect 4027 4288 4028 4292
rect 4022 4287 4028 4288
rect 4119 4291 4125 4292
rect 4119 4287 4120 4291
rect 4124 4290 4125 4291
rect 4138 4291 4144 4292
rect 4138 4290 4139 4291
rect 4124 4288 4139 4290
rect 4124 4287 4125 4288
rect 4002 4286 4008 4287
rect 4119 4286 4125 4287
rect 4138 4287 4139 4288
rect 4143 4287 4144 4291
rect 4158 4288 4159 4292
rect 4163 4288 4164 4292
rect 4158 4287 4164 4288
rect 4254 4291 4261 4292
rect 4254 4287 4255 4291
rect 4260 4287 4261 4291
rect 4310 4288 4311 4292
rect 4315 4288 4316 4292
rect 4310 4287 4316 4288
rect 4407 4291 4413 4292
rect 4407 4287 4408 4291
rect 4412 4290 4413 4291
rect 4490 4291 4496 4292
rect 4490 4290 4491 4291
rect 4412 4288 4491 4290
rect 4412 4287 4413 4288
rect 4138 4286 4144 4287
rect 4254 4286 4261 4287
rect 4407 4286 4413 4287
rect 4490 4287 4491 4288
rect 4495 4287 4496 4291
rect 4510 4288 4511 4292
rect 4515 4288 4516 4292
rect 4510 4287 4516 4288
rect 4607 4291 4613 4292
rect 4607 4287 4608 4291
rect 4612 4290 4613 4291
rect 4722 4291 4728 4292
rect 4722 4290 4723 4291
rect 4612 4288 4723 4290
rect 4612 4287 4613 4288
rect 4490 4286 4496 4287
rect 4607 4286 4613 4287
rect 4722 4287 4723 4288
rect 4727 4287 4728 4291
rect 4742 4288 4743 4292
rect 4747 4288 4748 4292
rect 4742 4287 4748 4288
rect 4839 4291 4845 4292
rect 4839 4287 4840 4291
rect 4844 4290 4845 4291
rect 4986 4291 4992 4292
rect 4986 4290 4987 4291
rect 4844 4288 4987 4290
rect 4844 4287 4845 4288
rect 4722 4286 4728 4287
rect 4839 4286 4845 4287
rect 4986 4287 4987 4288
rect 4991 4287 4992 4291
rect 5006 4288 5007 4292
rect 5011 4288 5012 4292
rect 5006 4287 5012 4288
rect 5103 4291 5109 4292
rect 5103 4287 5104 4291
rect 5108 4290 5109 4291
rect 5258 4291 5264 4292
rect 5258 4290 5259 4291
rect 5108 4288 5259 4290
rect 5108 4287 5109 4288
rect 4986 4286 4992 4287
rect 5103 4286 5109 4287
rect 5258 4287 5259 4288
rect 5263 4287 5264 4291
rect 5278 4288 5279 4292
rect 5283 4288 5284 4292
rect 5278 4287 5284 4288
rect 5375 4291 5381 4292
rect 5375 4287 5376 4291
rect 5380 4287 5381 4291
rect 5542 4288 5543 4292
rect 5547 4288 5548 4292
rect 5542 4287 5548 4288
rect 5638 4291 5645 4292
rect 5638 4287 5639 4291
rect 5644 4287 5645 4291
rect 5258 4286 5264 4287
rect 5375 4286 5381 4287
rect 5638 4286 5645 4287
rect 5662 4291 5668 4292
rect 5662 4287 5663 4291
rect 5667 4287 5668 4291
rect 5662 4286 5668 4287
rect 1517 4284 1594 4286
rect 1278 4282 1284 4283
rect 778 4278 784 4279
rect 1176 4278 1178 4281
rect 1239 4279 1245 4280
rect 1239 4278 1240 4279
rect 1176 4276 1240 4278
rect 1239 4275 1240 4276
rect 1244 4275 1245 4279
rect 1688 4278 1690 4281
rect 2022 4280 2028 4281
rect 2406 4280 2412 4281
rect 2830 4280 2836 4281
rect 3262 4280 3268 4281
rect 3678 4280 3684 4281
rect 1878 4279 1884 4280
rect 1878 4278 1879 4279
rect 1688 4276 1879 4278
rect 1239 4274 1245 4275
rect 1878 4275 1879 4276
rect 1883 4275 1884 4279
rect 1878 4274 1884 4275
rect 1974 4279 1980 4280
rect 1974 4275 1975 4279
rect 1979 4275 1980 4279
rect 2022 4276 2023 4280
rect 2027 4276 2028 4280
rect 2022 4275 2028 4276
rect 2119 4279 2125 4280
rect 2119 4275 2120 4279
rect 2124 4278 2125 4279
rect 2386 4279 2392 4280
rect 2386 4278 2387 4279
rect 2124 4276 2387 4278
rect 2124 4275 2125 4276
rect 1974 4274 1980 4275
rect 2119 4274 2125 4275
rect 2386 4275 2387 4276
rect 2391 4275 2392 4279
rect 2406 4276 2407 4280
rect 2411 4276 2412 4280
rect 2406 4275 2412 4276
rect 2502 4279 2509 4280
rect 2502 4275 2503 4279
rect 2508 4275 2509 4279
rect 2830 4276 2831 4280
rect 2835 4276 2836 4280
rect 2830 4275 2836 4276
rect 2926 4279 2933 4280
rect 2926 4275 2927 4279
rect 2932 4275 2933 4279
rect 3262 4276 3263 4280
rect 3267 4276 3268 4280
rect 3262 4275 3268 4276
rect 3358 4279 3365 4280
rect 3358 4275 3359 4279
rect 3364 4275 3365 4279
rect 3678 4276 3679 4280
rect 3683 4276 3684 4280
rect 3678 4275 3684 4276
rect 3775 4279 3784 4280
rect 3775 4275 3776 4279
rect 3783 4275 3784 4279
rect 2386 4274 2392 4275
rect 2502 4274 2509 4275
rect 2926 4274 2933 4275
rect 3358 4274 3365 4275
rect 3775 4274 3784 4275
rect 3798 4279 3804 4280
rect 3798 4275 3799 4279
rect 3803 4275 3804 4279
rect 3798 4274 3804 4275
rect 4550 4279 4556 4280
rect 4550 4275 4551 4279
rect 4555 4275 4556 4279
rect 4550 4274 4556 4275
rect 5376 4274 5378 4286
rect 4552 4272 5378 4274
rect 110 4236 116 4237
rect 1934 4236 1940 4237
rect 110 4232 111 4236
rect 115 4232 116 4236
rect 110 4231 116 4232
rect 626 4235 632 4236
rect 626 4231 627 4235
rect 631 4231 632 4235
rect 626 4230 632 4231
rect 770 4235 776 4236
rect 770 4231 771 4235
rect 775 4231 776 4235
rect 770 4230 776 4231
rect 922 4235 928 4236
rect 922 4231 923 4235
rect 927 4231 928 4235
rect 922 4230 928 4231
rect 1082 4235 1088 4236
rect 1082 4231 1083 4235
rect 1087 4231 1088 4235
rect 1082 4230 1088 4231
rect 1250 4235 1256 4236
rect 1250 4231 1251 4235
rect 1255 4231 1256 4235
rect 1250 4230 1256 4231
rect 1418 4235 1424 4236
rect 1418 4231 1419 4235
rect 1423 4231 1424 4235
rect 1418 4230 1424 4231
rect 1594 4235 1600 4236
rect 1594 4231 1595 4235
rect 1599 4231 1600 4235
rect 1934 4232 1935 4236
rect 1939 4232 1940 4236
rect 1934 4231 1940 4232
rect 3838 4233 3844 4234
rect 5662 4233 5668 4234
rect 1594 4230 1600 4231
rect 3838 4229 3839 4233
rect 3843 4229 3844 4233
rect 3838 4228 3844 4229
rect 3886 4232 3892 4233
rect 4022 4232 4028 4233
rect 4158 4232 4164 4233
rect 4302 4232 4308 4233
rect 4502 4232 4508 4233
rect 4734 4232 4740 4233
rect 4998 4232 5004 4233
rect 5270 4232 5276 4233
rect 5542 4232 5548 4233
rect 3886 4228 3887 4232
rect 3891 4228 3892 4232
rect 1239 4227 1245 4228
rect 3886 4227 3892 4228
rect 3983 4231 3992 4232
rect 3983 4227 3984 4231
rect 3991 4227 3992 4231
rect 4022 4228 4023 4232
rect 4027 4228 4028 4232
rect 4022 4227 4028 4228
rect 4119 4231 4128 4232
rect 4119 4227 4120 4231
rect 4127 4227 4128 4231
rect 4158 4228 4159 4232
rect 4163 4228 4164 4232
rect 4158 4227 4164 4228
rect 4255 4231 4261 4232
rect 4255 4227 4256 4231
rect 4260 4230 4261 4231
rect 4263 4231 4269 4232
rect 4263 4230 4264 4231
rect 4260 4228 4264 4230
rect 4260 4227 4261 4228
rect 1239 4223 1240 4227
rect 1244 4226 1245 4227
rect 3983 4226 3992 4227
rect 4119 4226 4128 4227
rect 4255 4226 4261 4227
rect 4263 4227 4264 4228
rect 4268 4227 4269 4231
rect 4302 4228 4303 4232
rect 4307 4228 4308 4232
rect 4302 4227 4308 4228
rect 4399 4231 4405 4232
rect 4399 4227 4400 4231
rect 4404 4230 4405 4231
rect 4446 4231 4452 4232
rect 4446 4230 4447 4231
rect 4404 4228 4447 4230
rect 4404 4227 4405 4228
rect 4263 4226 4269 4227
rect 4399 4226 4405 4227
rect 4446 4227 4447 4228
rect 4451 4227 4452 4231
rect 4502 4228 4503 4232
rect 4507 4228 4508 4232
rect 4502 4227 4508 4228
rect 4599 4231 4605 4232
rect 4599 4227 4600 4231
rect 4604 4230 4605 4231
rect 4615 4231 4621 4232
rect 4615 4230 4616 4231
rect 4604 4228 4616 4230
rect 4604 4227 4605 4228
rect 4446 4226 4452 4227
rect 4599 4226 4605 4227
rect 4615 4227 4616 4228
rect 4620 4227 4621 4231
rect 4734 4228 4735 4232
rect 4739 4228 4740 4232
rect 4734 4227 4740 4228
rect 4831 4231 4837 4232
rect 4831 4227 4832 4231
rect 4836 4230 4837 4231
rect 4887 4231 4893 4232
rect 4887 4230 4888 4231
rect 4836 4228 4888 4230
rect 4836 4227 4837 4228
rect 4615 4226 4621 4227
rect 4831 4226 4837 4227
rect 4887 4227 4888 4228
rect 4892 4227 4893 4231
rect 4998 4228 4999 4232
rect 5003 4228 5004 4232
rect 4998 4227 5004 4228
rect 5095 4231 5104 4232
rect 5095 4227 5096 4231
rect 5103 4227 5104 4231
rect 5270 4228 5271 4232
rect 5275 4228 5276 4232
rect 5270 4227 5276 4228
rect 5366 4231 5373 4232
rect 5366 4227 5367 4231
rect 5372 4227 5373 4231
rect 5542 4228 5543 4232
rect 5547 4228 5548 4232
rect 5542 4227 5548 4228
rect 5639 4231 5645 4232
rect 5639 4227 5640 4231
rect 5644 4230 5645 4231
rect 5647 4231 5653 4232
rect 5647 4230 5648 4231
rect 5644 4228 5648 4230
rect 5644 4227 5645 4228
rect 4887 4226 4893 4227
rect 5095 4226 5104 4227
rect 5366 4226 5373 4227
rect 5639 4226 5645 4227
rect 5647 4227 5648 4228
rect 5652 4227 5653 4231
rect 5662 4229 5663 4233
rect 5667 4229 5668 4233
rect 5662 4228 5668 4229
rect 5647 4226 5653 4227
rect 1244 4224 1378 4226
rect 1244 4223 1245 4224
rect 1239 4222 1245 4223
rect 1376 4222 1378 4224
rect 1375 4221 1381 4222
rect 654 4220 660 4221
rect 798 4220 804 4221
rect 950 4220 956 4221
rect 1110 4220 1116 4221
rect 1278 4220 1284 4221
rect 110 4219 116 4220
rect 110 4215 111 4219
rect 115 4215 116 4219
rect 654 4216 655 4220
rect 659 4216 660 4220
rect 654 4215 660 4216
rect 751 4219 757 4220
rect 751 4215 752 4219
rect 756 4218 757 4219
rect 778 4219 784 4220
rect 778 4218 779 4219
rect 756 4216 779 4218
rect 756 4215 757 4216
rect 110 4214 116 4215
rect 751 4214 757 4215
rect 778 4215 779 4216
rect 783 4215 784 4219
rect 798 4216 799 4220
rect 803 4216 804 4220
rect 798 4215 804 4216
rect 894 4219 901 4220
rect 894 4215 895 4219
rect 900 4215 901 4219
rect 950 4216 951 4220
rect 955 4216 956 4220
rect 950 4215 956 4216
rect 1046 4219 1053 4220
rect 1046 4215 1047 4219
rect 1052 4215 1053 4219
rect 1110 4216 1111 4220
rect 1115 4216 1116 4220
rect 1110 4215 1116 4216
rect 1206 4219 1213 4220
rect 1206 4215 1207 4219
rect 1212 4215 1213 4219
rect 1278 4216 1279 4220
rect 1283 4216 1284 4220
rect 1375 4217 1376 4221
rect 1380 4217 1381 4221
rect 1375 4216 1381 4217
rect 1446 4220 1452 4221
rect 1622 4220 1628 4221
rect 1446 4216 1447 4220
rect 1451 4216 1452 4220
rect 1278 4215 1284 4216
rect 1446 4215 1452 4216
rect 1542 4219 1549 4220
rect 1542 4215 1543 4219
rect 1548 4215 1549 4219
rect 1622 4216 1623 4220
rect 1627 4216 1628 4220
rect 1622 4215 1628 4216
rect 1714 4219 1725 4220
rect 1714 4215 1715 4219
rect 1719 4215 1720 4219
rect 1724 4215 1725 4219
rect 778 4214 784 4215
rect 894 4214 901 4215
rect 1046 4214 1053 4215
rect 1206 4214 1213 4215
rect 1542 4214 1549 4215
rect 1714 4214 1725 4215
rect 1934 4219 1940 4220
rect 1934 4215 1935 4219
rect 1939 4215 1940 4219
rect 3858 4217 3864 4218
rect 1934 4214 1940 4215
rect 3838 4216 3844 4217
rect 3838 4212 3839 4216
rect 3843 4212 3844 4216
rect 3858 4213 3859 4217
rect 3863 4213 3864 4217
rect 3858 4212 3864 4213
rect 3994 4217 4000 4218
rect 3994 4213 3995 4217
rect 3999 4213 4000 4217
rect 3994 4212 4000 4213
rect 4130 4217 4136 4218
rect 4130 4213 4131 4217
rect 4135 4213 4136 4217
rect 4130 4212 4136 4213
rect 4274 4217 4280 4218
rect 4274 4213 4275 4217
rect 4279 4213 4280 4217
rect 4274 4212 4280 4213
rect 4474 4217 4480 4218
rect 4474 4213 4475 4217
rect 4479 4213 4480 4217
rect 4474 4212 4480 4213
rect 4706 4217 4712 4218
rect 4706 4213 4707 4217
rect 4711 4213 4712 4217
rect 4706 4212 4712 4213
rect 4970 4217 4976 4218
rect 4970 4213 4971 4217
rect 4975 4213 4976 4217
rect 4970 4212 4976 4213
rect 5242 4217 5248 4218
rect 5242 4213 5243 4217
rect 5247 4213 5248 4217
rect 5242 4212 5248 4213
rect 5514 4217 5520 4218
rect 5514 4213 5515 4217
rect 5519 4213 5520 4217
rect 5514 4212 5520 4213
rect 5662 4216 5668 4217
rect 5662 4212 5663 4216
rect 5667 4212 5668 4216
rect 3838 4211 3844 4212
rect 5662 4211 5668 4212
rect 1974 4193 1980 4194
rect 3798 4193 3804 4194
rect 1974 4189 1975 4193
rect 1979 4189 1980 4193
rect 1974 4188 1980 4189
rect 2022 4192 2028 4193
rect 2190 4192 2196 4193
rect 2382 4192 2388 4193
rect 2582 4192 2588 4193
rect 2782 4192 2788 4193
rect 2982 4192 2988 4193
rect 2022 4188 2023 4192
rect 2027 4188 2028 4192
rect 2022 4187 2028 4188
rect 2119 4191 2128 4192
rect 2119 4187 2120 4191
rect 2127 4187 2128 4191
rect 2190 4188 2191 4192
rect 2195 4188 2196 4192
rect 2190 4187 2196 4188
rect 2286 4191 2293 4192
rect 2286 4187 2287 4191
rect 2292 4187 2293 4191
rect 2382 4188 2383 4192
rect 2387 4188 2388 4192
rect 2382 4187 2388 4188
rect 2478 4191 2485 4192
rect 2478 4187 2479 4191
rect 2484 4187 2485 4191
rect 2582 4188 2583 4192
rect 2587 4188 2588 4192
rect 2582 4187 2588 4188
rect 2679 4191 2688 4192
rect 2679 4187 2680 4191
rect 2687 4187 2688 4191
rect 2782 4188 2783 4192
rect 2787 4188 2788 4192
rect 2782 4187 2788 4188
rect 2879 4191 2888 4192
rect 2879 4187 2880 4191
rect 2887 4187 2888 4191
rect 2982 4188 2983 4192
rect 2987 4188 2988 4192
rect 2982 4187 2988 4188
rect 3079 4191 3085 4192
rect 3079 4187 3080 4191
rect 3084 4190 3085 4191
rect 3242 4191 3248 4192
rect 3242 4190 3243 4191
rect 3084 4188 3243 4190
rect 3084 4187 3085 4188
rect 2119 4186 2128 4187
rect 2286 4186 2293 4187
rect 2478 4186 2485 4187
rect 2679 4186 2688 4187
rect 2879 4186 2888 4187
rect 3079 4186 3085 4187
rect 3242 4187 3243 4188
rect 3247 4187 3248 4191
rect 3798 4189 3799 4193
rect 3803 4189 3804 4193
rect 3798 4188 3804 4189
rect 3242 4186 3248 4187
rect 1994 4177 2000 4178
rect 1974 4176 1980 4177
rect 1974 4172 1975 4176
rect 1979 4172 1980 4176
rect 1994 4173 1995 4177
rect 1999 4173 2000 4177
rect 1994 4172 2000 4173
rect 2162 4177 2168 4178
rect 2162 4173 2163 4177
rect 2167 4173 2168 4177
rect 2162 4172 2168 4173
rect 2354 4177 2360 4178
rect 2354 4173 2355 4177
rect 2359 4173 2360 4177
rect 2354 4172 2360 4173
rect 2554 4177 2560 4178
rect 2554 4173 2555 4177
rect 2559 4173 2560 4177
rect 2554 4172 2560 4173
rect 2754 4177 2760 4178
rect 2754 4173 2755 4177
rect 2759 4173 2760 4177
rect 2754 4172 2760 4173
rect 2954 4177 2960 4178
rect 2954 4173 2955 4177
rect 2959 4173 2960 4177
rect 2954 4172 2960 4173
rect 3798 4176 3804 4177
rect 3798 4172 3799 4176
rect 3803 4172 3804 4176
rect 1974 4171 1980 4172
rect 3798 4171 3804 4172
rect 3986 4167 3992 4168
rect 3956 4158 3958 4165
rect 3986 4163 3987 4167
rect 3991 4166 3992 4167
rect 4122 4167 4128 4168
rect 3991 4164 4001 4166
rect 3991 4163 3992 4164
rect 3986 4162 3992 4163
rect 4122 4163 4123 4167
rect 4127 4166 4128 4167
rect 4263 4167 4269 4168
rect 4127 4164 4137 4166
rect 4127 4163 4128 4164
rect 4122 4162 4128 4163
rect 4263 4163 4264 4167
rect 4268 4166 4269 4167
rect 4446 4167 4452 4168
rect 4268 4164 4281 4166
rect 4268 4163 4269 4164
rect 4263 4162 4269 4163
rect 4446 4163 4447 4167
rect 4451 4166 4452 4167
rect 4615 4167 4621 4168
rect 4451 4164 4481 4166
rect 4451 4163 4452 4164
rect 4446 4162 4452 4163
rect 4615 4163 4616 4167
rect 4620 4166 4621 4167
rect 4887 4167 4893 4168
rect 4620 4164 4713 4166
rect 4620 4163 4621 4164
rect 4615 4162 4621 4163
rect 4887 4163 4888 4167
rect 4892 4166 4893 4167
rect 5098 4167 5104 4168
rect 4892 4164 4977 4166
rect 4892 4163 4893 4164
rect 4887 4162 4893 4163
rect 5098 4163 5099 4167
rect 5103 4166 5104 4167
rect 5638 4167 5644 4168
rect 5638 4166 5639 4167
rect 5103 4164 5249 4166
rect 5613 4164 5639 4166
rect 5103 4163 5104 4164
rect 5098 4162 5104 4163
rect 5638 4163 5639 4164
rect 5643 4163 5644 4167
rect 5638 4162 5644 4163
rect 4254 4159 4260 4160
rect 4254 4158 4255 4159
rect 110 4157 116 4158
rect 1934 4157 1940 4158
rect 110 4153 111 4157
rect 115 4153 116 4157
rect 110 4152 116 4153
rect 518 4156 524 4157
rect 702 4156 708 4157
rect 894 4156 900 4157
rect 1102 4156 1108 4157
rect 1326 4156 1332 4157
rect 1550 4156 1556 4157
rect 1782 4156 1788 4157
rect 518 4152 519 4156
rect 523 4152 524 4156
rect 518 4151 524 4152
rect 615 4155 621 4156
rect 615 4151 616 4155
rect 620 4154 621 4155
rect 639 4155 645 4156
rect 639 4154 640 4155
rect 620 4152 640 4154
rect 620 4151 621 4152
rect 615 4150 621 4151
rect 639 4151 640 4152
rect 644 4151 645 4155
rect 702 4152 703 4156
rect 707 4152 708 4156
rect 702 4151 708 4152
rect 799 4155 808 4156
rect 799 4151 800 4155
rect 807 4151 808 4155
rect 894 4152 895 4156
rect 899 4152 900 4156
rect 894 4151 900 4152
rect 991 4155 1000 4156
rect 991 4151 992 4155
rect 999 4151 1000 4155
rect 1102 4152 1103 4156
rect 1107 4152 1108 4156
rect 1102 4151 1108 4152
rect 1199 4155 1208 4156
rect 1199 4151 1200 4155
rect 1207 4151 1208 4155
rect 1326 4152 1327 4156
rect 1331 4152 1332 4156
rect 1326 4151 1332 4152
rect 1418 4155 1429 4156
rect 1418 4151 1419 4155
rect 1423 4151 1424 4155
rect 1428 4151 1429 4155
rect 1550 4152 1551 4156
rect 1555 4152 1556 4156
rect 1550 4151 1556 4152
rect 1647 4155 1656 4156
rect 1647 4151 1648 4155
rect 1655 4151 1656 4155
rect 1782 4152 1783 4156
rect 1787 4152 1788 4156
rect 1782 4151 1788 4152
rect 1878 4155 1885 4156
rect 1878 4151 1879 4155
rect 1884 4151 1885 4155
rect 1934 4153 1935 4157
rect 1939 4153 1940 4157
rect 3956 4156 4255 4158
rect 4254 4155 4255 4156
rect 4259 4155 4260 4159
rect 4254 4154 4260 4155
rect 1934 4152 1940 4153
rect 639 4150 645 4151
rect 799 4150 808 4151
rect 991 4150 1000 4151
rect 1199 4150 1208 4151
rect 1418 4150 1429 4151
rect 1647 4150 1656 4151
rect 1878 4150 1885 4151
rect 490 4141 496 4142
rect 110 4140 116 4141
rect 110 4136 111 4140
rect 115 4136 116 4140
rect 490 4137 491 4141
rect 495 4137 496 4141
rect 490 4136 496 4137
rect 674 4141 680 4142
rect 674 4137 675 4141
rect 679 4137 680 4141
rect 674 4136 680 4137
rect 866 4141 872 4142
rect 866 4137 867 4141
rect 871 4137 872 4141
rect 866 4136 872 4137
rect 1074 4141 1080 4142
rect 1074 4137 1075 4141
rect 1079 4137 1080 4141
rect 1074 4136 1080 4137
rect 1298 4141 1304 4142
rect 1298 4137 1299 4141
rect 1303 4137 1304 4141
rect 1298 4136 1304 4137
rect 1522 4141 1528 4142
rect 1522 4137 1523 4141
rect 1527 4137 1528 4141
rect 1522 4136 1528 4137
rect 1754 4141 1760 4142
rect 1754 4137 1755 4141
rect 1759 4137 1760 4141
rect 1754 4136 1760 4137
rect 1934 4140 1940 4141
rect 1934 4136 1935 4140
rect 1939 4136 1940 4140
rect 110 4135 116 4136
rect 1934 4135 1940 4136
rect 586 4127 592 4128
rect 586 4123 587 4127
rect 591 4126 592 4127
rect 1418 4127 1424 4128
rect 1418 4126 1419 4127
rect 591 4124 1419 4126
rect 591 4123 592 4124
rect 586 4122 592 4123
rect 1418 4123 1419 4124
rect 1423 4123 1424 4127
rect 2122 4127 2128 4128
rect 1418 4122 1424 4123
rect 2092 4118 2094 4125
rect 2122 4123 2123 4127
rect 2127 4126 2128 4127
rect 2502 4127 2508 4128
rect 2502 4126 2503 4127
rect 2127 4124 2169 4126
rect 2453 4124 2503 4126
rect 2127 4123 2128 4124
rect 2122 4122 2128 4123
rect 2502 4123 2503 4124
rect 2507 4123 2508 4127
rect 2502 4122 2508 4123
rect 2566 4127 2572 4128
rect 2566 4123 2567 4127
rect 2571 4123 2572 4127
rect 2566 4122 2572 4123
rect 2682 4127 2688 4128
rect 2682 4123 2683 4127
rect 2687 4126 2688 4127
rect 2882 4127 2888 4128
rect 2687 4124 2761 4126
rect 2687 4123 2688 4124
rect 2682 4122 2688 4123
rect 2882 4123 2883 4127
rect 2887 4126 2888 4127
rect 2887 4124 2961 4126
rect 2887 4123 2888 4124
rect 2882 4122 2888 4123
rect 2478 4119 2484 4120
rect 2478 4118 2479 4119
rect 2092 4116 2479 4118
rect 2478 4115 2479 4116
rect 2483 4115 2484 4119
rect 2478 4114 2484 4115
rect 5090 4103 5096 4104
rect 5090 4102 5091 4103
rect 4700 4100 5091 4102
rect 3078 4099 3084 4100
rect 3078 4098 3079 4099
rect 2936 4096 3079 4098
rect 2247 4095 2253 4096
rect 2247 4094 2248 4095
rect 2173 4092 2248 4094
rect 586 4091 592 4092
rect 586 4087 587 4091
rect 591 4087 592 4091
rect 586 4086 592 4087
rect 639 4091 645 4092
rect 639 4087 640 4091
rect 644 4090 645 4091
rect 886 4091 892 4092
rect 644 4088 681 4090
rect 644 4087 645 4088
rect 639 4086 645 4087
rect 886 4087 887 4091
rect 891 4087 892 4091
rect 886 4086 892 4087
rect 994 4091 1000 4092
rect 994 4087 995 4091
rect 999 4090 1000 4091
rect 1202 4091 1208 4092
rect 999 4088 1081 4090
rect 999 4087 1000 4088
rect 994 4086 1000 4087
rect 1202 4087 1203 4091
rect 1207 4090 1208 4091
rect 1614 4091 1620 4092
rect 1207 4088 1305 4090
rect 1207 4087 1208 4088
rect 1202 4086 1208 4087
rect 1614 4087 1615 4091
rect 1619 4087 1620 4091
rect 1614 4086 1620 4087
rect 1650 4091 1656 4092
rect 1650 4087 1651 4091
rect 1655 4090 1656 4091
rect 2247 4091 2248 4092
rect 2252 4091 2253 4095
rect 2247 4090 2253 4091
rect 2286 4095 2292 4096
rect 2286 4091 2287 4095
rect 2291 4091 2292 4095
rect 2746 4095 2752 4096
rect 2746 4094 2747 4095
rect 2717 4092 2747 4094
rect 2286 4090 2292 4091
rect 2538 4091 2544 4092
rect 1655 4088 1761 4090
rect 1655 4087 1656 4088
rect 1650 4086 1656 4087
rect 2538 4087 2539 4091
rect 2543 4087 2544 4091
rect 2746 4091 2747 4092
rect 2751 4091 2752 4095
rect 2936 4094 2938 4096
rect 3078 4095 3079 4096
rect 3083 4095 3084 4099
rect 3078 4094 3084 4095
rect 4700 4094 4702 4100
rect 5090 4099 5091 4100
rect 5095 4099 5096 4103
rect 5090 4098 5096 4099
rect 5230 4099 5236 4100
rect 5230 4098 5231 4099
rect 5100 4096 5231 4098
rect 5100 4094 5102 4096
rect 5230 4095 5231 4096
rect 5235 4095 5236 4099
rect 5230 4094 5236 4095
rect 5422 4095 5428 4096
rect 2885 4092 2938 4094
rect 4661 4092 4702 4094
rect 5069 4092 5102 4094
rect 2746 4090 2752 4091
rect 3138 4091 3144 4092
rect 2538 4086 2544 4087
rect 3048 4086 3050 4089
rect 3103 4087 3109 4088
rect 3103 4086 3104 4087
rect 3048 4084 3104 4086
rect 3103 4083 3104 4084
rect 3108 4083 3109 4087
rect 3138 4087 3139 4091
rect 3143 4087 3144 4091
rect 3138 4086 3144 4087
rect 4706 4091 4712 4092
rect 4706 4087 4707 4091
rect 4711 4087 4712 4091
rect 4706 4086 4712 4087
rect 4842 4091 4848 4092
rect 4842 4087 4843 4091
rect 4847 4087 4848 4091
rect 4842 4086 4848 4087
rect 5202 4091 5208 4092
rect 5202 4087 5203 4091
rect 5207 4087 5208 4091
rect 5202 4086 5208 4087
rect 5338 4091 5344 4092
rect 5338 4087 5339 4091
rect 5343 4087 5344 4091
rect 5422 4091 5423 4095
rect 5427 4091 5428 4095
rect 5647 4095 5653 4096
rect 5647 4094 5648 4095
rect 5613 4092 5648 4094
rect 5422 4090 5428 4091
rect 5647 4091 5648 4092
rect 5652 4091 5653 4095
rect 5647 4090 5653 4091
rect 5338 4086 5344 4087
rect 3103 4082 3109 4083
rect 462 4063 468 4064
rect 462 4062 463 4063
rect 259 4060 463 4062
rect 259 4058 261 4060
rect 462 4059 463 4060
rect 467 4059 468 4063
rect 2538 4063 2544 4064
rect 462 4058 468 4059
rect 794 4059 800 4060
rect 794 4058 795 4059
rect 229 4056 261 4058
rect 693 4056 795 4058
rect 794 4055 795 4056
rect 799 4055 800 4059
rect 794 4054 800 4055
rect 802 4059 808 4060
rect 802 4055 803 4059
rect 807 4058 808 4059
rect 1906 4059 1912 4060
rect 1906 4058 1907 4059
rect 807 4056 881 4058
rect 1885 4056 1907 4058
rect 807 4055 808 4056
rect 802 4054 808 4055
rect 1186 4055 1192 4056
rect 432 4050 434 4053
rect 527 4051 533 4052
rect 527 4050 528 4051
rect 432 4048 528 4050
rect 527 4047 528 4048
rect 532 4047 533 4051
rect 1186 4051 1187 4055
rect 1191 4051 1192 4055
rect 1186 4050 1192 4051
rect 1586 4055 1592 4056
rect 1586 4051 1587 4055
rect 1591 4051 1592 4055
rect 1906 4055 1907 4056
rect 1911 4055 1912 4059
rect 2538 4059 2539 4063
rect 2543 4062 2544 4063
rect 2738 4063 2744 4064
rect 2738 4062 2739 4063
rect 2543 4060 2739 4062
rect 2543 4059 2544 4060
rect 2538 4058 2544 4059
rect 2738 4059 2739 4060
rect 2743 4059 2744 4063
rect 2738 4058 2744 4059
rect 5202 4063 5208 4064
rect 5202 4059 5203 4063
rect 5207 4062 5208 4063
rect 5366 4063 5372 4064
rect 5366 4062 5367 4063
rect 5207 4060 5367 4062
rect 5207 4059 5208 4060
rect 5202 4058 5208 4059
rect 5366 4059 5367 4060
rect 5371 4059 5372 4063
rect 5366 4058 5372 4059
rect 1906 4054 1912 4055
rect 5338 4055 5344 4056
rect 1586 4050 1592 4051
rect 5338 4051 5339 4055
rect 5343 4054 5344 4055
rect 5498 4055 5504 4056
rect 5498 4054 5499 4055
rect 5343 4052 5499 4054
rect 5343 4051 5344 4052
rect 5338 4050 5344 4051
rect 5498 4051 5499 4052
rect 5503 4051 5504 4055
rect 5498 4050 5504 4051
rect 527 4046 533 4047
rect 1974 4044 1980 4045
rect 3798 4044 3804 4045
rect 1974 4040 1975 4044
rect 1979 4040 1980 4044
rect 1974 4039 1980 4040
rect 2074 4043 2080 4044
rect 2074 4039 2075 4043
rect 2079 4039 2080 4043
rect 2074 4038 2080 4039
rect 2258 4043 2264 4044
rect 2258 4039 2259 4043
rect 2263 4039 2264 4043
rect 2258 4038 2264 4039
rect 2442 4043 2448 4044
rect 2442 4039 2443 4043
rect 2447 4039 2448 4043
rect 2442 4038 2448 4039
rect 2618 4043 2624 4044
rect 2618 4039 2619 4043
rect 2623 4039 2624 4043
rect 2618 4038 2624 4039
rect 2786 4043 2792 4044
rect 2786 4039 2787 4043
rect 2791 4039 2792 4043
rect 2786 4038 2792 4039
rect 2954 4043 2960 4044
rect 2954 4039 2955 4043
rect 2959 4039 2960 4043
rect 2954 4038 2960 4039
rect 3130 4043 3136 4044
rect 3130 4039 3131 4043
rect 3135 4039 3136 4043
rect 3798 4040 3799 4044
rect 3803 4040 3804 4044
rect 3798 4039 3804 4040
rect 3838 4044 3844 4045
rect 5662 4044 5668 4045
rect 3838 4040 3839 4044
rect 3843 4040 3844 4044
rect 3838 4039 3844 4040
rect 4562 4043 4568 4044
rect 4562 4039 4563 4043
rect 4567 4039 4568 4043
rect 3130 4038 3136 4039
rect 4562 4038 4568 4039
rect 4698 4043 4704 4044
rect 4698 4039 4699 4043
rect 4703 4039 4704 4043
rect 4698 4038 4704 4039
rect 4834 4043 4840 4044
rect 4834 4039 4835 4043
rect 4839 4039 4840 4043
rect 4834 4038 4840 4039
rect 4970 4043 4976 4044
rect 4970 4039 4971 4043
rect 4975 4039 4976 4043
rect 4970 4038 4976 4039
rect 5106 4043 5112 4044
rect 5106 4039 5107 4043
rect 5111 4039 5112 4043
rect 5106 4038 5112 4039
rect 5242 4043 5248 4044
rect 5242 4039 5243 4043
rect 5247 4039 5248 4043
rect 5242 4038 5248 4039
rect 5378 4043 5384 4044
rect 5378 4039 5379 4043
rect 5383 4039 5384 4043
rect 5378 4038 5384 4039
rect 5514 4043 5520 4044
rect 5514 4039 5515 4043
rect 5519 4039 5520 4043
rect 5662 4040 5663 4044
rect 5667 4040 5668 4044
rect 5662 4039 5668 4040
rect 5514 4038 5520 4039
rect 1586 4035 1592 4036
rect 1586 4031 1587 4035
rect 1591 4034 1592 4035
rect 1914 4035 1920 4036
rect 1914 4034 1915 4035
rect 1591 4032 1915 4034
rect 1591 4031 1592 4032
rect 1586 4030 1592 4031
rect 1914 4031 1915 4032
rect 1919 4031 1920 4035
rect 1914 4030 1920 4031
rect 2247 4035 2253 4036
rect 2247 4031 2248 4035
rect 2252 4034 2253 4035
rect 2746 4035 2752 4036
rect 2252 4032 2386 4034
rect 2252 4031 2253 4032
rect 2247 4030 2253 4031
rect 2384 4030 2386 4032
rect 2746 4031 2747 4035
rect 2751 4034 2752 4035
rect 3103 4035 3109 4036
rect 2751 4032 2914 4034
rect 2751 4031 2752 4032
rect 2746 4030 2752 4031
rect 2912 4030 2914 4032
rect 3103 4031 3104 4035
rect 3108 4034 3109 4035
rect 3108 4032 3258 4034
rect 3108 4031 3109 4032
rect 3103 4030 3109 4031
rect 3256 4030 3258 4032
rect 2383 4029 2389 4030
rect 2911 4029 2917 4030
rect 3255 4029 3261 4030
rect 2102 4028 2108 4029
rect 2286 4028 2292 4029
rect 1974 4027 1980 4028
rect 1974 4023 1975 4027
rect 1979 4023 1980 4027
rect 2102 4024 2103 4028
rect 2107 4024 2108 4028
rect 2102 4023 2108 4024
rect 2194 4027 2205 4028
rect 2194 4023 2195 4027
rect 2199 4023 2200 4027
rect 2204 4023 2205 4027
rect 2286 4024 2287 4028
rect 2291 4024 2292 4028
rect 2383 4025 2384 4029
rect 2388 4025 2389 4029
rect 2383 4024 2389 4025
rect 2470 4028 2476 4029
rect 2646 4028 2652 4029
rect 2814 4028 2820 4029
rect 2470 4024 2471 4028
rect 2475 4024 2476 4028
rect 2286 4023 2292 4024
rect 2470 4023 2476 4024
rect 2566 4027 2573 4028
rect 2566 4023 2567 4027
rect 2572 4023 2573 4027
rect 2646 4024 2647 4028
rect 2651 4024 2652 4028
rect 2646 4023 2652 4024
rect 2742 4027 2749 4028
rect 2742 4023 2743 4027
rect 2748 4023 2749 4027
rect 2814 4024 2815 4028
rect 2819 4024 2820 4028
rect 2911 4025 2912 4029
rect 2916 4025 2917 4029
rect 2911 4024 2917 4025
rect 2982 4028 2988 4029
rect 3158 4028 3164 4029
rect 2982 4024 2983 4028
rect 2987 4024 2988 4028
rect 2814 4023 2820 4024
rect 2982 4023 2988 4024
rect 3078 4027 3085 4028
rect 3078 4023 3079 4027
rect 3084 4023 3085 4027
rect 3158 4024 3159 4028
rect 3163 4024 3164 4028
rect 3255 4025 3256 4029
rect 3260 4025 3261 4029
rect 4590 4028 4596 4029
rect 4726 4028 4732 4029
rect 4862 4028 4868 4029
rect 4998 4028 5004 4029
rect 5134 4028 5140 4029
rect 5270 4028 5276 4029
rect 5406 4028 5412 4029
rect 5542 4028 5548 4029
rect 3255 4024 3261 4025
rect 3798 4027 3804 4028
rect 3158 4023 3164 4024
rect 3798 4023 3799 4027
rect 3803 4023 3804 4027
rect 1974 4022 1980 4023
rect 2194 4022 2205 4023
rect 2566 4022 2573 4023
rect 2742 4022 2749 4023
rect 3078 4022 3085 4023
rect 3798 4022 3804 4023
rect 3838 4027 3844 4028
rect 3838 4023 3839 4027
rect 3843 4023 3844 4027
rect 4590 4024 4591 4028
rect 4595 4024 4596 4028
rect 4590 4023 4596 4024
rect 4687 4027 4693 4028
rect 4687 4023 4688 4027
rect 4692 4026 4693 4027
rect 4706 4027 4712 4028
rect 4706 4026 4707 4027
rect 4692 4024 4707 4026
rect 4692 4023 4693 4024
rect 3838 4022 3844 4023
rect 4687 4022 4693 4023
rect 4706 4023 4707 4024
rect 4711 4023 4712 4027
rect 4726 4024 4727 4028
rect 4731 4024 4732 4028
rect 4726 4023 4732 4024
rect 4823 4027 4829 4028
rect 4823 4023 4824 4027
rect 4828 4026 4829 4027
rect 4842 4027 4848 4028
rect 4842 4026 4843 4027
rect 4828 4024 4843 4026
rect 4828 4023 4829 4024
rect 4706 4022 4712 4023
rect 4823 4022 4829 4023
rect 4842 4023 4843 4024
rect 4847 4023 4848 4027
rect 4862 4024 4863 4028
rect 4867 4024 4868 4028
rect 4862 4023 4868 4024
rect 4958 4027 4965 4028
rect 4958 4023 4959 4027
rect 4964 4023 4965 4027
rect 4998 4024 4999 4028
rect 5003 4024 5004 4028
rect 4998 4023 5004 4024
rect 5090 4027 5101 4028
rect 5090 4023 5091 4027
rect 5095 4023 5096 4027
rect 5100 4023 5101 4027
rect 5134 4024 5135 4028
rect 5139 4024 5140 4028
rect 5134 4023 5140 4024
rect 5230 4027 5237 4028
rect 5230 4023 5231 4027
rect 5236 4023 5237 4027
rect 5270 4024 5271 4028
rect 5275 4024 5276 4028
rect 5270 4023 5276 4024
rect 5366 4027 5373 4028
rect 5366 4023 5367 4027
rect 5372 4023 5373 4027
rect 5406 4024 5407 4028
rect 5411 4024 5412 4028
rect 5406 4023 5412 4024
rect 5498 4027 5509 4028
rect 5498 4023 5499 4027
rect 5503 4023 5504 4027
rect 5508 4023 5509 4027
rect 5542 4024 5543 4028
rect 5547 4024 5548 4028
rect 5542 4023 5548 4024
rect 5638 4027 5645 4028
rect 5638 4023 5639 4027
rect 5644 4023 5645 4027
rect 4842 4022 4848 4023
rect 4958 4022 4965 4023
rect 5090 4022 5101 4023
rect 5230 4022 5237 4023
rect 5366 4022 5373 4023
rect 5498 4022 5509 4023
rect 5638 4022 5645 4023
rect 5662 4027 5668 4028
rect 5662 4023 5663 4027
rect 5667 4023 5668 4027
rect 5662 4022 5668 4023
rect 110 4008 116 4009
rect 1934 4008 1940 4009
rect 110 4004 111 4008
rect 115 4004 116 4008
rect 110 4003 116 4004
rect 130 4007 136 4008
rect 130 4003 131 4007
rect 135 4003 136 4007
rect 130 4002 136 4003
rect 338 4007 344 4008
rect 338 4003 339 4007
rect 343 4003 344 4007
rect 338 4002 344 4003
rect 594 4007 600 4008
rect 594 4003 595 4007
rect 599 4003 600 4007
rect 594 4002 600 4003
rect 874 4007 880 4008
rect 874 4003 875 4007
rect 879 4003 880 4007
rect 874 4002 880 4003
rect 1178 4007 1184 4008
rect 1178 4003 1179 4007
rect 1183 4003 1184 4007
rect 1178 4002 1184 4003
rect 1490 4007 1496 4008
rect 1490 4003 1491 4007
rect 1495 4003 1496 4007
rect 1490 4002 1496 4003
rect 1786 4007 1792 4008
rect 1786 4003 1787 4007
rect 1791 4003 1792 4007
rect 1934 4004 1935 4008
rect 1939 4004 1940 4008
rect 1934 4003 1940 4004
rect 1786 4002 1792 4003
rect 527 3999 533 4000
rect 527 3995 528 3999
rect 532 3998 533 3999
rect 794 3999 800 4000
rect 532 3996 722 3998
rect 532 3995 533 3996
rect 527 3994 533 3995
rect 720 3994 722 3996
rect 794 3995 795 3999
rect 799 3998 800 3999
rect 799 3996 1306 3998
rect 799 3995 800 3996
rect 794 3994 800 3995
rect 719 3993 725 3994
rect 158 3992 164 3993
rect 366 3992 372 3993
rect 622 3992 628 3993
rect 110 3991 116 3992
rect 110 3987 111 3991
rect 115 3987 116 3991
rect 158 3988 159 3992
rect 163 3988 164 3992
rect 158 3987 164 3988
rect 254 3991 261 3992
rect 254 3987 255 3991
rect 260 3987 261 3991
rect 366 3988 367 3992
rect 371 3988 372 3992
rect 366 3987 372 3988
rect 462 3991 469 3992
rect 462 3987 463 3991
rect 468 3987 469 3991
rect 622 3988 623 3992
rect 627 3988 628 3992
rect 719 3989 720 3993
rect 724 3989 725 3993
rect 719 3988 725 3989
rect 902 3992 908 3993
rect 1206 3992 1212 3993
rect 1304 3992 1306 3996
rect 1518 3992 1524 3993
rect 1814 3992 1820 3993
rect 902 3988 903 3992
rect 907 3988 908 3992
rect 622 3987 628 3988
rect 902 3987 908 3988
rect 999 3991 1005 3992
rect 999 3987 1000 3991
rect 1004 3990 1005 3991
rect 1186 3991 1192 3992
rect 1186 3990 1187 3991
rect 1004 3988 1187 3990
rect 1004 3987 1005 3988
rect 110 3986 116 3987
rect 254 3986 261 3987
rect 462 3986 469 3987
rect 999 3986 1005 3987
rect 1186 3987 1187 3988
rect 1191 3987 1192 3991
rect 1206 3988 1207 3992
rect 1211 3988 1212 3992
rect 1206 3987 1212 3988
rect 1303 3991 1309 3992
rect 1303 3987 1304 3991
rect 1308 3987 1309 3991
rect 1518 3988 1519 3992
rect 1523 3988 1524 3992
rect 1518 3987 1524 3988
rect 1614 3991 1621 3992
rect 1614 3987 1615 3991
rect 1620 3987 1621 3991
rect 1814 3988 1815 3992
rect 1819 3988 1820 3992
rect 1814 3987 1820 3988
rect 1911 3991 1920 3992
rect 1911 3987 1912 3991
rect 1919 3987 1920 3991
rect 1186 3986 1192 3987
rect 1303 3986 1309 3987
rect 1614 3986 1621 3987
rect 1911 3986 1920 3987
rect 1934 3991 1940 3992
rect 1934 3987 1935 3991
rect 1939 3987 1940 3991
rect 1934 3986 1940 3987
rect 1974 3961 1980 3962
rect 3798 3961 3804 3962
rect 1974 3957 1975 3961
rect 1979 3957 1980 3961
rect 1974 3956 1980 3957
rect 2126 3960 2132 3961
rect 2310 3960 2316 3961
rect 2486 3960 2492 3961
rect 2662 3960 2668 3961
rect 2830 3960 2836 3961
rect 2998 3960 3004 3961
rect 3174 3960 3180 3961
rect 3350 3960 3356 3961
rect 2126 3956 2127 3960
rect 2131 3956 2132 3960
rect 2126 3955 2132 3956
rect 2223 3959 2229 3960
rect 2223 3955 2224 3959
rect 2228 3958 2229 3959
rect 2247 3959 2253 3960
rect 2247 3958 2248 3959
rect 2228 3956 2248 3958
rect 2228 3955 2229 3956
rect 2223 3954 2229 3955
rect 2247 3955 2248 3956
rect 2252 3955 2253 3959
rect 2310 3956 2311 3960
rect 2315 3956 2316 3960
rect 2310 3955 2316 3956
rect 2407 3959 2413 3960
rect 2407 3955 2408 3959
rect 2412 3958 2413 3959
rect 2423 3959 2429 3960
rect 2423 3958 2424 3959
rect 2412 3956 2424 3958
rect 2412 3955 2413 3956
rect 2247 3954 2253 3955
rect 2407 3954 2413 3955
rect 2423 3955 2424 3956
rect 2428 3955 2429 3959
rect 2486 3956 2487 3960
rect 2491 3956 2492 3960
rect 2486 3955 2492 3956
rect 2578 3959 2589 3960
rect 2578 3955 2579 3959
rect 2583 3955 2584 3959
rect 2588 3955 2589 3959
rect 2662 3956 2663 3960
rect 2667 3956 2668 3960
rect 2662 3955 2668 3956
rect 2759 3959 2765 3960
rect 2759 3955 2760 3959
rect 2764 3958 2765 3959
rect 2767 3959 2773 3960
rect 2767 3958 2768 3959
rect 2764 3956 2768 3958
rect 2764 3955 2765 3956
rect 2423 3954 2429 3955
rect 2578 3954 2589 3955
rect 2759 3954 2765 3955
rect 2767 3955 2768 3956
rect 2772 3955 2773 3959
rect 2830 3956 2831 3960
rect 2835 3956 2836 3960
rect 2830 3955 2836 3956
rect 2926 3959 2933 3960
rect 2926 3955 2927 3959
rect 2932 3955 2933 3959
rect 2998 3956 2999 3960
rect 3003 3956 3004 3960
rect 2998 3955 3004 3956
rect 3095 3959 3101 3960
rect 3095 3955 3096 3959
rect 3100 3958 3101 3959
rect 3138 3959 3144 3960
rect 3138 3958 3139 3959
rect 3100 3956 3139 3958
rect 3100 3955 3101 3956
rect 2767 3954 2773 3955
rect 2926 3954 2933 3955
rect 3095 3954 3101 3955
rect 3138 3955 3139 3956
rect 3143 3955 3144 3959
rect 3174 3956 3175 3960
rect 3179 3956 3180 3960
rect 3174 3955 3180 3956
rect 3266 3959 3277 3960
rect 3266 3955 3267 3959
rect 3271 3955 3272 3959
rect 3276 3955 3277 3959
rect 3350 3956 3351 3960
rect 3355 3956 3356 3960
rect 3350 3955 3356 3956
rect 3446 3959 3453 3960
rect 3446 3955 3447 3959
rect 3452 3955 3453 3959
rect 3798 3957 3799 3961
rect 3803 3957 3804 3961
rect 3798 3956 3804 3957
rect 3138 3954 3144 3955
rect 3266 3954 3277 3955
rect 3446 3954 3453 3955
rect 3838 3949 3844 3950
rect 5662 3949 5668 3950
rect 2098 3945 2104 3946
rect 1974 3944 1980 3945
rect 362 3943 368 3944
rect 362 3939 363 3943
rect 367 3942 368 3943
rect 367 3940 1154 3942
rect 367 3939 368 3940
rect 362 3938 368 3939
rect 1152 3930 1154 3940
rect 1974 3940 1975 3944
rect 1979 3940 1980 3944
rect 2098 3941 2099 3945
rect 2103 3941 2104 3945
rect 2098 3940 2104 3941
rect 2282 3945 2288 3946
rect 2282 3941 2283 3945
rect 2287 3941 2288 3945
rect 2282 3940 2288 3941
rect 2458 3945 2464 3946
rect 2458 3941 2459 3945
rect 2463 3941 2464 3945
rect 2458 3940 2464 3941
rect 2634 3945 2640 3946
rect 2634 3941 2635 3945
rect 2639 3941 2640 3945
rect 2634 3940 2640 3941
rect 2802 3945 2808 3946
rect 2802 3941 2803 3945
rect 2807 3941 2808 3945
rect 2802 3940 2808 3941
rect 2970 3945 2976 3946
rect 2970 3941 2971 3945
rect 2975 3941 2976 3945
rect 2970 3940 2976 3941
rect 3146 3945 3152 3946
rect 3146 3941 3147 3945
rect 3151 3941 3152 3945
rect 3146 3940 3152 3941
rect 3322 3945 3328 3946
rect 3838 3945 3839 3949
rect 3843 3945 3844 3949
rect 3322 3941 3323 3945
rect 3327 3941 3328 3945
rect 3322 3940 3328 3941
rect 3798 3944 3804 3945
rect 3838 3944 3844 3945
rect 4358 3948 4364 3949
rect 4542 3948 4548 3949
rect 4734 3948 4740 3949
rect 4926 3948 4932 3949
rect 5126 3948 5132 3949
rect 5326 3948 5332 3949
rect 5526 3948 5532 3949
rect 4358 3944 4359 3948
rect 4363 3944 4364 3948
rect 3798 3940 3799 3944
rect 3803 3940 3804 3944
rect 4358 3943 4364 3944
rect 4455 3947 4461 3948
rect 4455 3943 4456 3947
rect 4460 3946 4461 3947
rect 4470 3947 4476 3948
rect 4470 3946 4471 3947
rect 4460 3944 4471 3946
rect 4460 3943 4461 3944
rect 4455 3942 4461 3943
rect 4470 3943 4471 3944
rect 4475 3943 4476 3947
rect 4542 3944 4543 3948
rect 4547 3944 4548 3948
rect 4542 3943 4548 3944
rect 4639 3947 4648 3948
rect 4639 3943 4640 3947
rect 4647 3943 4648 3947
rect 4734 3944 4735 3948
rect 4739 3944 4740 3948
rect 4734 3943 4740 3944
rect 4826 3947 4837 3948
rect 4826 3943 4827 3947
rect 4831 3943 4832 3947
rect 4836 3943 4837 3947
rect 4926 3944 4927 3948
rect 4931 3944 4932 3948
rect 4926 3943 4932 3944
rect 5022 3947 5029 3948
rect 5022 3943 5023 3947
rect 5028 3943 5029 3947
rect 5126 3944 5127 3948
rect 5131 3944 5132 3948
rect 5126 3943 5132 3944
rect 5223 3947 5229 3948
rect 5223 3943 5224 3947
rect 5228 3946 5229 3947
rect 5271 3947 5277 3948
rect 5271 3946 5272 3947
rect 5228 3944 5272 3946
rect 5228 3943 5229 3944
rect 4470 3942 4476 3943
rect 4639 3942 4648 3943
rect 4826 3942 4837 3943
rect 5022 3942 5029 3943
rect 5223 3942 5229 3943
rect 5271 3943 5272 3944
rect 5276 3943 5277 3947
rect 5326 3944 5327 3948
rect 5331 3944 5332 3948
rect 5326 3943 5332 3944
rect 5422 3947 5429 3948
rect 5422 3943 5423 3947
rect 5428 3943 5429 3947
rect 5526 3944 5527 3948
rect 5531 3944 5532 3948
rect 5526 3943 5532 3944
rect 5618 3947 5629 3948
rect 5618 3943 5619 3947
rect 5623 3943 5624 3947
rect 5628 3943 5629 3947
rect 5662 3945 5663 3949
rect 5667 3945 5668 3949
rect 5662 3944 5668 3945
rect 5271 3942 5277 3943
rect 5422 3942 5429 3943
rect 5618 3942 5629 3943
rect 1974 3939 1980 3940
rect 3798 3939 3804 3940
rect 4330 3933 4336 3934
rect 3838 3932 3844 3933
rect 110 3929 116 3930
rect 1151 3929 1157 3930
rect 1934 3929 1940 3930
rect 110 3925 111 3929
rect 115 3925 116 3929
rect 110 3924 116 3925
rect 158 3928 164 3929
rect 342 3928 348 3929
rect 566 3928 572 3929
rect 806 3928 812 3929
rect 1054 3928 1060 3929
rect 158 3924 159 3928
rect 163 3924 164 3928
rect 158 3923 164 3924
rect 255 3927 261 3928
rect 255 3923 256 3927
rect 260 3926 261 3927
rect 274 3927 280 3928
rect 274 3926 275 3927
rect 260 3924 275 3926
rect 260 3923 261 3924
rect 255 3922 261 3923
rect 274 3923 275 3924
rect 279 3923 280 3927
rect 342 3924 343 3928
rect 347 3924 348 3928
rect 342 3923 348 3924
rect 438 3927 445 3928
rect 438 3923 439 3927
rect 444 3923 445 3927
rect 566 3924 567 3928
rect 571 3924 572 3928
rect 566 3923 572 3924
rect 663 3927 669 3928
rect 663 3923 664 3927
rect 668 3926 669 3927
rect 694 3927 700 3928
rect 694 3926 695 3927
rect 668 3924 695 3926
rect 668 3923 669 3924
rect 274 3922 280 3923
rect 438 3922 445 3923
rect 663 3922 669 3923
rect 694 3923 695 3924
rect 699 3923 700 3927
rect 806 3924 807 3928
rect 811 3924 812 3928
rect 806 3923 812 3924
rect 903 3927 909 3928
rect 903 3923 904 3927
rect 908 3926 909 3927
rect 942 3927 948 3928
rect 942 3926 943 3927
rect 908 3924 943 3926
rect 908 3923 909 3924
rect 694 3922 700 3923
rect 903 3922 909 3923
rect 942 3923 943 3924
rect 947 3923 948 3927
rect 1054 3924 1055 3928
rect 1059 3924 1060 3928
rect 1151 3925 1152 3929
rect 1156 3925 1157 3929
rect 1151 3924 1157 3925
rect 1310 3928 1316 3929
rect 1574 3928 1580 3929
rect 1814 3928 1820 3929
rect 1310 3924 1311 3928
rect 1315 3924 1316 3928
rect 1054 3923 1060 3924
rect 1310 3923 1316 3924
rect 1407 3927 1413 3928
rect 1407 3923 1408 3927
rect 1412 3926 1413 3927
rect 1431 3927 1437 3928
rect 1431 3926 1432 3927
rect 1412 3924 1432 3926
rect 1412 3923 1413 3924
rect 942 3922 948 3923
rect 1407 3922 1413 3923
rect 1431 3923 1432 3924
rect 1436 3923 1437 3927
rect 1574 3924 1575 3928
rect 1579 3924 1580 3928
rect 1574 3923 1580 3924
rect 1671 3927 1677 3928
rect 1671 3923 1672 3927
rect 1676 3926 1677 3927
rect 1695 3927 1701 3928
rect 1695 3926 1696 3927
rect 1676 3924 1696 3926
rect 1676 3923 1677 3924
rect 1431 3922 1437 3923
rect 1671 3922 1677 3923
rect 1695 3923 1696 3924
rect 1700 3923 1701 3927
rect 1814 3924 1815 3928
rect 1819 3924 1820 3928
rect 1814 3923 1820 3924
rect 1906 3927 1917 3928
rect 1906 3923 1907 3927
rect 1911 3923 1912 3927
rect 1916 3923 1917 3927
rect 1934 3925 1935 3929
rect 1939 3925 1940 3929
rect 3838 3928 3839 3932
rect 3843 3928 3844 3932
rect 4330 3929 4331 3933
rect 4335 3929 4336 3933
rect 4330 3928 4336 3929
rect 4514 3933 4520 3934
rect 4514 3929 4515 3933
rect 4519 3929 4520 3933
rect 4514 3928 4520 3929
rect 4706 3933 4712 3934
rect 4706 3929 4707 3933
rect 4711 3929 4712 3933
rect 4706 3928 4712 3929
rect 4898 3933 4904 3934
rect 4898 3929 4899 3933
rect 4903 3929 4904 3933
rect 4898 3928 4904 3929
rect 5098 3933 5104 3934
rect 5098 3929 5099 3933
rect 5103 3929 5104 3933
rect 5098 3928 5104 3929
rect 5298 3933 5304 3934
rect 5298 3929 5299 3933
rect 5303 3929 5304 3933
rect 5298 3928 5304 3929
rect 5498 3933 5504 3934
rect 5498 3929 5499 3933
rect 5503 3929 5504 3933
rect 5498 3928 5504 3929
rect 5662 3932 5668 3933
rect 5662 3928 5663 3932
rect 5667 3928 5668 3932
rect 3838 3927 3844 3928
rect 5662 3927 5668 3928
rect 1934 3924 1940 3925
rect 1695 3922 1701 3923
rect 1906 3922 1917 3923
rect 2730 3923 2736 3924
rect 2730 3919 2731 3923
rect 2735 3922 2736 3923
rect 3266 3923 3272 3924
rect 3266 3922 3267 3923
rect 2735 3920 3267 3922
rect 2735 3919 2736 3920
rect 2730 3918 2736 3919
rect 3266 3919 3267 3920
rect 3271 3919 3272 3923
rect 3266 3918 3272 3919
rect 4426 3915 4432 3916
rect 130 3913 136 3914
rect 110 3912 116 3913
rect 110 3908 111 3912
rect 115 3908 116 3912
rect 130 3909 131 3913
rect 135 3909 136 3913
rect 130 3908 136 3909
rect 314 3913 320 3914
rect 314 3909 315 3913
rect 319 3909 320 3913
rect 314 3908 320 3909
rect 538 3913 544 3914
rect 538 3909 539 3913
rect 543 3909 544 3913
rect 538 3908 544 3909
rect 778 3913 784 3914
rect 778 3909 779 3913
rect 783 3909 784 3913
rect 778 3908 784 3909
rect 1026 3913 1032 3914
rect 1026 3909 1027 3913
rect 1031 3909 1032 3913
rect 1026 3908 1032 3909
rect 1282 3913 1288 3914
rect 1282 3909 1283 3913
rect 1287 3909 1288 3913
rect 1282 3908 1288 3909
rect 1546 3913 1552 3914
rect 1546 3909 1547 3913
rect 1551 3909 1552 3913
rect 1546 3908 1552 3909
rect 1786 3913 1792 3914
rect 1786 3909 1787 3913
rect 1791 3909 1792 3913
rect 1786 3908 1792 3909
rect 1934 3912 1940 3913
rect 1934 3908 1935 3912
rect 1939 3908 1940 3912
rect 4426 3911 4427 3915
rect 4431 3914 4432 3915
rect 4826 3915 4832 3916
rect 4826 3914 4827 3915
rect 4431 3912 4827 3914
rect 4431 3911 4432 3912
rect 4426 3910 4432 3911
rect 4826 3911 4827 3912
rect 4831 3911 4832 3915
rect 4826 3910 4832 3911
rect 110 3907 116 3908
rect 1934 3907 1940 3908
rect 2194 3895 2200 3896
rect 2194 3891 2195 3895
rect 2199 3891 2200 3895
rect 2194 3890 2200 3891
rect 2247 3895 2253 3896
rect 2247 3891 2248 3895
rect 2252 3894 2253 3895
rect 2423 3895 2429 3896
rect 2252 3892 2289 3894
rect 2252 3891 2253 3892
rect 2247 3890 2253 3891
rect 2423 3891 2424 3895
rect 2428 3894 2429 3895
rect 2730 3895 2736 3896
rect 2428 3892 2465 3894
rect 2428 3891 2429 3892
rect 2423 3890 2429 3891
rect 2730 3891 2731 3895
rect 2735 3891 2736 3895
rect 2730 3890 2736 3891
rect 2767 3895 2773 3896
rect 2767 3891 2768 3895
rect 2772 3894 2773 3895
rect 2926 3895 2932 3896
rect 2772 3892 2809 3894
rect 2772 3891 2773 3892
rect 2767 3890 2773 3891
rect 2926 3891 2927 3895
rect 2931 3894 2932 3895
rect 3282 3895 3288 3896
rect 2931 3892 2977 3894
rect 2931 3891 2932 3892
rect 2926 3890 2932 3891
rect 3244 3886 3246 3893
rect 3282 3891 3283 3895
rect 3287 3894 3288 3895
rect 3287 3892 3329 3894
rect 3287 3891 3288 3892
rect 3282 3890 3288 3891
rect 3446 3887 3452 3888
rect 3446 3886 3447 3887
rect 3244 3884 3447 3886
rect 3446 3883 3447 3884
rect 3451 3883 3452 3887
rect 3446 3882 3452 3883
rect 4426 3883 4432 3884
rect 4426 3879 4427 3883
rect 4431 3879 4432 3883
rect 4426 3878 4432 3879
rect 4470 3883 4476 3884
rect 4470 3879 4471 3883
rect 4475 3882 4476 3883
rect 4958 3883 4964 3884
rect 4475 3880 4521 3882
rect 4475 3879 4476 3880
rect 4470 3878 4476 3879
rect 4804 3874 4806 3881
rect 4958 3879 4959 3883
rect 4963 3879 4964 3883
rect 4958 3878 4964 3879
rect 5034 3883 5040 3884
rect 5034 3879 5035 3883
rect 5039 3882 5040 3883
rect 5271 3883 5277 3884
rect 5039 3880 5105 3882
rect 5039 3879 5040 3880
rect 5034 3878 5040 3879
rect 5271 3879 5272 3883
rect 5276 3882 5277 3883
rect 5638 3883 5644 3884
rect 5638 3882 5639 3883
rect 5276 3880 5305 3882
rect 5597 3880 5639 3882
rect 5276 3879 5277 3880
rect 5271 3878 5277 3879
rect 5638 3879 5639 3880
rect 5643 3879 5644 3883
rect 5638 3878 5644 3879
rect 5022 3875 5028 3876
rect 5022 3874 5023 3875
rect 4804 3872 5023 3874
rect 5022 3871 5023 3872
rect 5027 3871 5028 3875
rect 5022 3870 5028 3871
rect 254 3863 260 3864
rect 254 3862 255 3863
rect 229 3860 255 3862
rect 254 3859 255 3860
rect 259 3859 260 3863
rect 254 3858 260 3859
rect 274 3863 280 3864
rect 274 3859 275 3863
rect 279 3862 280 3863
rect 438 3863 444 3864
rect 279 3860 321 3862
rect 279 3859 280 3860
rect 274 3858 280 3859
rect 438 3859 439 3863
rect 443 3862 444 3863
rect 694 3863 700 3864
rect 443 3860 545 3862
rect 443 3859 444 3860
rect 438 3858 444 3859
rect 694 3859 695 3863
rect 699 3862 700 3863
rect 942 3863 948 3864
rect 699 3860 785 3862
rect 699 3859 700 3860
rect 694 3858 700 3859
rect 942 3859 943 3863
rect 947 3862 948 3863
rect 1378 3863 1384 3864
rect 947 3860 1033 3862
rect 947 3859 948 3860
rect 942 3858 948 3859
rect 1378 3859 1379 3863
rect 1383 3859 1384 3863
rect 1378 3858 1384 3859
rect 1431 3863 1437 3864
rect 1431 3859 1432 3863
rect 1436 3862 1437 3863
rect 1695 3863 1701 3864
rect 1436 3860 1553 3862
rect 1436 3859 1437 3860
rect 1431 3858 1437 3859
rect 1695 3859 1696 3863
rect 1700 3862 1701 3863
rect 2578 3863 2584 3864
rect 1700 3860 1793 3862
rect 1700 3859 1701 3860
rect 1695 3858 1701 3859
rect 2578 3859 2579 3863
rect 2583 3859 2584 3863
rect 2578 3858 2584 3859
rect 2440 3856 2582 3858
rect 2440 3854 2442 3856
rect 2938 3855 2944 3856
rect 2938 3854 2939 3855
rect 2389 3852 2442 3854
rect 2837 3852 2939 3854
rect 2530 3851 2536 3852
rect 2530 3847 2531 3851
rect 2535 3847 2536 3851
rect 2938 3851 2939 3852
rect 2943 3851 2944 3855
rect 3390 3855 3396 3856
rect 2938 3850 2944 3851
rect 2954 3851 2960 3852
rect 2530 3846 2536 3847
rect 2954 3847 2955 3851
rect 2959 3847 2960 3851
rect 2954 3846 2960 3847
rect 3162 3851 3168 3852
rect 3162 3847 3163 3851
rect 3167 3847 3168 3851
rect 3390 3851 3391 3855
rect 3395 3851 3396 3855
rect 3390 3850 3396 3851
rect 3570 3851 3576 3852
rect 3162 3846 3168 3847
rect 3570 3847 3571 3851
rect 3575 3847 3576 3851
rect 3570 3846 3576 3847
rect 5446 3847 5452 3848
rect 5446 3846 5447 3847
rect 5299 3844 5447 3846
rect 4255 3843 4261 3844
rect 4255 3842 4256 3843
rect 4149 3840 4256 3842
rect 4255 3839 4256 3840
rect 4260 3839 4261 3843
rect 4474 3843 4480 3844
rect 4474 3842 4475 3843
rect 4365 3840 4475 3842
rect 4255 3838 4261 3839
rect 4474 3839 4475 3840
rect 4479 3839 4480 3843
rect 4634 3843 4640 3844
rect 4634 3842 4635 3843
rect 4581 3840 4635 3842
rect 4474 3838 4480 3839
rect 4634 3839 4635 3840
rect 4639 3839 4640 3843
rect 4634 3838 4640 3839
rect 4642 3843 4648 3844
rect 4642 3839 4643 3843
rect 4647 3842 4648 3843
rect 5098 3843 5104 3844
rect 5098 3842 5099 3843
rect 4647 3840 4705 3842
rect 5005 3840 5099 3842
rect 4647 3839 4648 3840
rect 4642 3838 4648 3839
rect 5098 3839 5099 3840
rect 5103 3839 5104 3843
rect 5299 3842 5301 3844
rect 5446 3843 5447 3844
rect 5451 3843 5452 3847
rect 5446 3842 5452 3843
rect 5618 3843 5624 3844
rect 5618 3842 5619 3843
rect 5213 3840 5301 3842
rect 5613 3840 5619 3842
rect 5098 3838 5104 3839
rect 5618 3839 5619 3840
rect 5623 3839 5624 3843
rect 5618 3838 5624 3839
rect 5416 3834 5418 3837
rect 5479 3835 5485 3836
rect 5479 3834 5480 3835
rect 5416 3832 5480 3834
rect 5479 3831 5480 3832
rect 5484 3831 5485 3835
rect 5479 3830 5485 3831
rect 362 3823 368 3824
rect 362 3819 363 3823
rect 367 3819 368 3823
rect 1854 3823 1860 3824
rect 362 3818 368 3819
rect 482 3819 488 3820
rect 482 3815 483 3819
rect 487 3815 488 3819
rect 482 3814 488 3815
rect 714 3819 720 3820
rect 714 3815 715 3819
rect 719 3815 720 3819
rect 714 3814 720 3815
rect 970 3819 976 3820
rect 970 3815 971 3819
rect 975 3815 976 3819
rect 970 3814 976 3815
rect 1242 3819 1248 3820
rect 1242 3815 1243 3819
rect 1247 3815 1248 3819
rect 1242 3814 1248 3815
rect 1610 3819 1616 3820
rect 1610 3815 1611 3819
rect 1615 3815 1616 3819
rect 1854 3819 1855 3823
rect 1859 3819 1860 3823
rect 1854 3818 1860 3819
rect 1610 3814 1616 3815
rect 1974 3804 1980 3805
rect 3798 3804 3804 3805
rect 1974 3800 1975 3804
rect 1979 3800 1980 3804
rect 1974 3799 1980 3800
rect 2290 3803 2296 3804
rect 2290 3799 2291 3803
rect 2295 3799 2296 3803
rect 2290 3798 2296 3799
rect 2522 3803 2528 3804
rect 2522 3799 2523 3803
rect 2527 3799 2528 3803
rect 2522 3798 2528 3799
rect 2738 3803 2744 3804
rect 2738 3799 2739 3803
rect 2743 3799 2744 3803
rect 2738 3798 2744 3799
rect 2946 3803 2952 3804
rect 2946 3799 2947 3803
rect 2951 3799 2952 3803
rect 2946 3798 2952 3799
rect 3154 3803 3160 3804
rect 3154 3799 3155 3803
rect 3159 3799 3160 3803
rect 3154 3798 3160 3799
rect 3354 3803 3360 3804
rect 3354 3799 3355 3803
rect 3359 3799 3360 3803
rect 3354 3798 3360 3799
rect 3562 3803 3568 3804
rect 3562 3799 3563 3803
rect 3567 3799 3568 3803
rect 3798 3800 3799 3804
rect 3803 3800 3804 3804
rect 3798 3799 3804 3800
rect 3562 3798 3568 3799
rect 1610 3795 1616 3796
rect 1610 3791 1611 3795
rect 1615 3794 1616 3795
rect 1910 3795 1916 3796
rect 1910 3794 1911 3795
rect 1615 3792 1911 3794
rect 1615 3791 1616 3792
rect 1610 3790 1616 3791
rect 1910 3791 1911 3792
rect 1915 3791 1916 3795
rect 1910 3790 1916 3791
rect 2938 3795 2944 3796
rect 2938 3791 2939 3795
rect 2943 3794 2944 3795
rect 2943 3792 3690 3794
rect 2943 3791 2944 3792
rect 2938 3790 2944 3791
rect 3688 3790 3690 3792
rect 3838 3792 3844 3793
rect 5662 3792 5668 3793
rect 3687 3789 3693 3790
rect 2318 3788 2324 3789
rect 2550 3788 2556 3789
rect 2766 3788 2772 3789
rect 2974 3788 2980 3789
rect 3182 3788 3188 3789
rect 3382 3788 3388 3789
rect 3590 3788 3596 3789
rect 1974 3787 1980 3788
rect 1974 3783 1975 3787
rect 1979 3783 1980 3787
rect 2318 3784 2319 3788
rect 2323 3784 2324 3788
rect 2318 3783 2324 3784
rect 2415 3787 2421 3788
rect 2415 3783 2416 3787
rect 2420 3786 2421 3787
rect 2530 3787 2536 3788
rect 2530 3786 2531 3787
rect 2420 3784 2531 3786
rect 2420 3783 2421 3784
rect 1974 3782 1980 3783
rect 2415 3782 2421 3783
rect 2530 3783 2531 3784
rect 2535 3783 2536 3787
rect 2550 3784 2551 3788
rect 2555 3784 2556 3788
rect 2550 3783 2556 3784
rect 2646 3787 2653 3788
rect 2646 3783 2647 3787
rect 2652 3783 2653 3787
rect 2766 3784 2767 3788
rect 2771 3784 2772 3788
rect 2766 3783 2772 3784
rect 2863 3787 2869 3788
rect 2863 3783 2864 3787
rect 2868 3786 2869 3787
rect 2954 3787 2960 3788
rect 2954 3786 2955 3787
rect 2868 3784 2955 3786
rect 2868 3783 2869 3784
rect 2530 3782 2536 3783
rect 2646 3782 2653 3783
rect 2863 3782 2869 3783
rect 2954 3783 2955 3784
rect 2959 3783 2960 3787
rect 2974 3784 2975 3788
rect 2979 3784 2980 3788
rect 2974 3783 2980 3784
rect 3071 3787 3077 3788
rect 3071 3783 3072 3787
rect 3076 3786 3077 3787
rect 3162 3787 3168 3788
rect 3162 3786 3163 3787
rect 3076 3784 3163 3786
rect 3076 3783 3077 3784
rect 2954 3782 2960 3783
rect 3071 3782 3077 3783
rect 3162 3783 3163 3784
rect 3167 3783 3168 3787
rect 3182 3784 3183 3788
rect 3187 3784 3188 3788
rect 3182 3783 3188 3784
rect 3279 3787 3288 3788
rect 3279 3783 3280 3787
rect 3287 3783 3288 3787
rect 3382 3784 3383 3788
rect 3387 3784 3388 3788
rect 3382 3783 3388 3784
rect 3479 3787 3485 3788
rect 3479 3783 3480 3787
rect 3484 3786 3485 3787
rect 3570 3787 3576 3788
rect 3570 3786 3571 3787
rect 3484 3784 3571 3786
rect 3484 3783 3485 3784
rect 3162 3782 3168 3783
rect 3279 3782 3288 3783
rect 3479 3782 3485 3783
rect 3570 3783 3571 3784
rect 3575 3783 3576 3787
rect 3590 3784 3591 3788
rect 3595 3784 3596 3788
rect 3687 3785 3688 3789
rect 3692 3785 3693 3789
rect 3838 3788 3839 3792
rect 3843 3788 3844 3792
rect 3687 3784 3693 3785
rect 3798 3787 3804 3788
rect 3838 3787 3844 3788
rect 4050 3791 4056 3792
rect 4050 3787 4051 3791
rect 4055 3787 4056 3791
rect 3590 3783 3596 3784
rect 3798 3783 3799 3787
rect 3803 3783 3804 3787
rect 4050 3786 4056 3787
rect 4266 3791 4272 3792
rect 4266 3787 4267 3791
rect 4271 3787 4272 3791
rect 4266 3786 4272 3787
rect 4482 3791 4488 3792
rect 4482 3787 4483 3791
rect 4487 3787 4488 3791
rect 4482 3786 4488 3787
rect 4698 3791 4704 3792
rect 4698 3787 4699 3791
rect 4703 3787 4704 3791
rect 4698 3786 4704 3787
rect 4906 3791 4912 3792
rect 4906 3787 4907 3791
rect 4911 3787 4912 3791
rect 4906 3786 4912 3787
rect 5114 3791 5120 3792
rect 5114 3787 5115 3791
rect 5119 3787 5120 3791
rect 5114 3786 5120 3787
rect 5322 3791 5328 3792
rect 5322 3787 5323 3791
rect 5327 3787 5328 3791
rect 5322 3786 5328 3787
rect 5514 3791 5520 3792
rect 5514 3787 5515 3791
rect 5519 3787 5520 3791
rect 5662 3788 5663 3792
rect 5667 3788 5668 3792
rect 5662 3787 5668 3788
rect 5514 3786 5520 3787
rect 3570 3782 3576 3783
rect 3798 3782 3804 3783
rect 4255 3783 4261 3784
rect 4255 3779 4256 3783
rect 4260 3782 4261 3783
rect 4474 3783 4480 3784
rect 4260 3780 4394 3782
rect 4260 3779 4261 3780
rect 4255 3778 4261 3779
rect 4078 3776 4084 3777
rect 4294 3776 4300 3777
rect 4392 3776 4394 3780
rect 4474 3779 4475 3783
rect 4479 3782 4480 3783
rect 4634 3783 4640 3784
rect 4479 3780 4611 3782
rect 4479 3779 4480 3780
rect 4474 3778 4480 3779
rect 4510 3776 4516 3777
rect 4609 3776 4611 3780
rect 4634 3779 4635 3783
rect 4639 3782 4640 3783
rect 5098 3783 5104 3784
rect 4639 3780 4826 3782
rect 4639 3779 4640 3780
rect 4634 3778 4640 3779
rect 4726 3776 4732 3777
rect 4824 3776 4826 3780
rect 5098 3779 5099 3783
rect 5103 3782 5104 3783
rect 5479 3783 5485 3784
rect 5103 3780 5242 3782
rect 5103 3779 5104 3780
rect 5098 3778 5104 3779
rect 4934 3776 4940 3777
rect 5142 3776 5148 3777
rect 5240 3776 5242 3780
rect 5479 3779 5480 3783
rect 5484 3782 5485 3783
rect 5484 3780 5643 3782
rect 5484 3779 5485 3780
rect 5479 3778 5485 3779
rect 5350 3776 5356 3777
rect 5542 3776 5548 3777
rect 5641 3776 5643 3780
rect 3838 3775 3844 3776
rect 110 3772 116 3773
rect 1934 3772 1940 3773
rect 110 3768 111 3772
rect 115 3768 116 3772
rect 110 3767 116 3768
rect 266 3771 272 3772
rect 266 3767 267 3771
rect 271 3767 272 3771
rect 266 3766 272 3767
rect 474 3771 480 3772
rect 474 3767 475 3771
rect 479 3767 480 3771
rect 474 3766 480 3767
rect 706 3771 712 3772
rect 706 3767 707 3771
rect 711 3767 712 3771
rect 706 3766 712 3767
rect 962 3771 968 3772
rect 962 3767 963 3771
rect 967 3767 968 3771
rect 962 3766 968 3767
rect 1234 3771 1240 3772
rect 1234 3767 1235 3771
rect 1239 3767 1240 3771
rect 1234 3766 1240 3767
rect 1514 3771 1520 3772
rect 1514 3767 1515 3771
rect 1519 3767 1520 3771
rect 1514 3766 1520 3767
rect 1786 3771 1792 3772
rect 1786 3767 1787 3771
rect 1791 3767 1792 3771
rect 1934 3768 1935 3772
rect 1939 3768 1940 3772
rect 3838 3771 3839 3775
rect 3843 3771 3844 3775
rect 4078 3772 4079 3776
rect 4083 3772 4084 3776
rect 4078 3771 4084 3772
rect 4170 3775 4181 3776
rect 4170 3771 4171 3775
rect 4175 3771 4176 3775
rect 4180 3771 4181 3775
rect 4294 3772 4295 3776
rect 4299 3772 4300 3776
rect 4294 3771 4300 3772
rect 4391 3775 4397 3776
rect 4391 3771 4392 3775
rect 4396 3771 4397 3775
rect 4510 3772 4511 3776
rect 4515 3772 4516 3776
rect 4510 3771 4516 3772
rect 4607 3775 4613 3776
rect 4607 3771 4608 3775
rect 4612 3771 4613 3775
rect 4726 3772 4727 3776
rect 4731 3772 4732 3776
rect 4726 3771 4732 3772
rect 4823 3775 4829 3776
rect 4823 3771 4824 3775
rect 4828 3771 4829 3775
rect 4934 3772 4935 3776
rect 4939 3772 4940 3776
rect 4934 3771 4940 3772
rect 5031 3775 5040 3776
rect 5031 3771 5032 3775
rect 5039 3771 5040 3775
rect 5142 3772 5143 3776
rect 5147 3772 5148 3776
rect 5142 3771 5148 3772
rect 5239 3775 5245 3776
rect 5239 3771 5240 3775
rect 5244 3771 5245 3775
rect 5350 3772 5351 3776
rect 5355 3772 5356 3776
rect 5350 3771 5356 3772
rect 5446 3775 5453 3776
rect 5446 3771 5447 3775
rect 5452 3771 5453 3775
rect 5542 3772 5543 3776
rect 5547 3772 5548 3776
rect 5542 3771 5548 3772
rect 5639 3775 5645 3776
rect 5639 3771 5640 3775
rect 5644 3771 5645 3775
rect 3838 3770 3844 3771
rect 4170 3770 4181 3771
rect 4391 3770 4397 3771
rect 4607 3770 4613 3771
rect 4823 3770 4829 3771
rect 5031 3770 5040 3771
rect 5239 3770 5245 3771
rect 5446 3770 5453 3771
rect 5639 3770 5645 3771
rect 5662 3775 5668 3776
rect 5662 3771 5663 3775
rect 5667 3771 5668 3775
rect 5662 3770 5668 3771
rect 1934 3767 1940 3768
rect 1786 3766 1792 3767
rect 1378 3763 1384 3764
rect 1378 3759 1379 3763
rect 1383 3762 1384 3763
rect 1383 3760 1642 3762
rect 1383 3759 1384 3760
rect 1378 3758 1384 3759
rect 1640 3758 1642 3760
rect 1639 3757 1645 3758
rect 294 3756 300 3757
rect 502 3756 508 3757
rect 734 3756 740 3757
rect 990 3756 996 3757
rect 1262 3756 1268 3757
rect 1542 3756 1548 3757
rect 110 3755 116 3756
rect 110 3751 111 3755
rect 115 3751 116 3755
rect 294 3752 295 3756
rect 299 3752 300 3756
rect 294 3751 300 3752
rect 391 3755 397 3756
rect 391 3751 392 3755
rect 396 3754 397 3755
rect 482 3755 488 3756
rect 482 3754 483 3755
rect 396 3752 483 3754
rect 396 3751 397 3752
rect 110 3750 116 3751
rect 391 3750 397 3751
rect 482 3751 483 3752
rect 487 3751 488 3755
rect 502 3752 503 3756
rect 507 3752 508 3756
rect 502 3751 508 3752
rect 599 3755 605 3756
rect 599 3751 600 3755
rect 604 3754 605 3755
rect 714 3755 720 3756
rect 714 3754 715 3755
rect 604 3752 715 3754
rect 604 3751 605 3752
rect 482 3750 488 3751
rect 599 3750 605 3751
rect 714 3751 715 3752
rect 719 3751 720 3755
rect 734 3752 735 3756
rect 739 3752 740 3756
rect 734 3751 740 3752
rect 831 3755 837 3756
rect 831 3751 832 3755
rect 836 3754 837 3755
rect 970 3755 976 3756
rect 970 3754 971 3755
rect 836 3752 971 3754
rect 836 3751 837 3752
rect 714 3750 720 3751
rect 831 3750 837 3751
rect 970 3751 971 3752
rect 975 3751 976 3755
rect 990 3752 991 3756
rect 995 3752 996 3756
rect 990 3751 996 3752
rect 1087 3755 1093 3756
rect 1087 3751 1088 3755
rect 1092 3754 1093 3755
rect 1242 3755 1248 3756
rect 1242 3754 1243 3755
rect 1092 3752 1243 3754
rect 1092 3751 1093 3752
rect 970 3750 976 3751
rect 1087 3750 1093 3751
rect 1242 3751 1243 3752
rect 1247 3751 1248 3755
rect 1262 3752 1263 3756
rect 1267 3752 1268 3756
rect 1262 3751 1268 3752
rect 1359 3755 1365 3756
rect 1359 3751 1360 3755
rect 1364 3751 1365 3755
rect 1542 3752 1543 3756
rect 1547 3752 1548 3756
rect 1639 3753 1640 3757
rect 1644 3753 1645 3757
rect 1639 3752 1645 3753
rect 1814 3756 1820 3757
rect 1814 3752 1815 3756
rect 1819 3752 1820 3756
rect 1542 3751 1548 3752
rect 1814 3751 1820 3752
rect 1910 3755 1917 3756
rect 1910 3751 1911 3755
rect 1916 3751 1917 3755
rect 1242 3750 1248 3751
rect 1359 3750 1365 3751
rect 1910 3750 1917 3751
rect 1934 3755 1940 3756
rect 1934 3751 1935 3755
rect 1939 3751 1940 3755
rect 1934 3750 1940 3751
rect 698 3739 704 3740
rect 698 3735 699 3739
rect 703 3738 704 3739
rect 1360 3738 1362 3750
rect 703 3736 1362 3738
rect 703 3735 704 3736
rect 698 3734 704 3735
rect 1974 3725 1980 3726
rect 3798 3725 3804 3726
rect 1974 3721 1975 3725
rect 1979 3721 1980 3725
rect 1974 3720 1980 3721
rect 2406 3724 2412 3725
rect 2646 3724 2652 3725
rect 2870 3724 2876 3725
rect 3086 3724 3092 3725
rect 3294 3724 3300 3725
rect 3494 3724 3500 3725
rect 3678 3724 3684 3725
rect 2406 3720 2407 3724
rect 2411 3720 2412 3724
rect 2406 3719 2412 3720
rect 2502 3723 2509 3724
rect 2502 3719 2503 3723
rect 2508 3719 2509 3723
rect 2646 3720 2647 3724
rect 2651 3720 2652 3724
rect 2646 3719 2652 3720
rect 2742 3723 2749 3724
rect 2742 3719 2743 3723
rect 2748 3719 2749 3723
rect 2870 3720 2871 3724
rect 2875 3720 2876 3724
rect 2870 3719 2876 3720
rect 2967 3723 2976 3724
rect 2967 3719 2968 3723
rect 2975 3719 2976 3723
rect 3086 3720 3087 3724
rect 3091 3720 3092 3724
rect 3086 3719 3092 3720
rect 3183 3723 3192 3724
rect 3183 3719 3184 3723
rect 3191 3719 3192 3723
rect 3294 3720 3295 3724
rect 3299 3720 3300 3724
rect 3294 3719 3300 3720
rect 3390 3723 3397 3724
rect 3390 3719 3391 3723
rect 3396 3719 3397 3723
rect 3494 3720 3495 3724
rect 3499 3720 3500 3724
rect 3494 3719 3500 3720
rect 3590 3723 3597 3724
rect 3590 3719 3591 3723
rect 3596 3719 3597 3723
rect 3678 3720 3679 3724
rect 3683 3720 3684 3724
rect 3678 3719 3684 3720
rect 3770 3723 3781 3724
rect 3770 3719 3771 3723
rect 3775 3719 3776 3723
rect 3780 3719 3781 3723
rect 3798 3721 3799 3725
rect 3803 3721 3804 3725
rect 3798 3720 3804 3721
rect 2502 3718 2509 3719
rect 2742 3718 2749 3719
rect 2967 3718 2976 3719
rect 3183 3718 3192 3719
rect 3390 3718 3397 3719
rect 3590 3718 3597 3719
rect 3770 3718 3781 3719
rect 2378 3709 2384 3710
rect 1974 3708 1980 3709
rect 1974 3704 1975 3708
rect 1979 3704 1980 3708
rect 2378 3705 2379 3709
rect 2383 3705 2384 3709
rect 2378 3704 2384 3705
rect 2618 3709 2624 3710
rect 2618 3705 2619 3709
rect 2623 3705 2624 3709
rect 2618 3704 2624 3705
rect 2842 3709 2848 3710
rect 2842 3705 2843 3709
rect 2847 3705 2848 3709
rect 2842 3704 2848 3705
rect 3058 3709 3064 3710
rect 3058 3705 3059 3709
rect 3063 3705 3064 3709
rect 3058 3704 3064 3705
rect 3266 3709 3272 3710
rect 3266 3705 3267 3709
rect 3271 3705 3272 3709
rect 3266 3704 3272 3705
rect 3466 3709 3472 3710
rect 3466 3705 3467 3709
rect 3471 3705 3472 3709
rect 3466 3704 3472 3705
rect 3650 3709 3656 3710
rect 3650 3705 3651 3709
rect 3655 3705 3656 3709
rect 3650 3704 3656 3705
rect 3798 3708 3804 3709
rect 3798 3704 3799 3708
rect 3803 3704 3804 3708
rect 1974 3703 1980 3704
rect 3798 3703 3804 3704
rect 110 3693 116 3694
rect 1934 3693 1940 3694
rect 110 3689 111 3693
rect 115 3689 116 3693
rect 110 3688 116 3689
rect 630 3692 636 3693
rect 774 3692 780 3693
rect 926 3692 932 3693
rect 1086 3692 1092 3693
rect 1254 3692 1260 3693
rect 1422 3692 1428 3693
rect 1590 3692 1596 3693
rect 1758 3692 1764 3693
rect 630 3688 631 3692
rect 635 3688 636 3692
rect 630 3687 636 3688
rect 727 3691 736 3692
rect 727 3687 728 3691
rect 735 3687 736 3691
rect 774 3688 775 3692
rect 779 3688 780 3692
rect 774 3687 780 3688
rect 871 3691 877 3692
rect 871 3687 872 3691
rect 876 3690 877 3691
rect 887 3691 893 3692
rect 887 3690 888 3691
rect 876 3688 888 3690
rect 876 3687 877 3688
rect 727 3686 736 3687
rect 871 3686 877 3687
rect 887 3687 888 3688
rect 892 3687 893 3691
rect 926 3688 927 3692
rect 931 3688 932 3692
rect 926 3687 932 3688
rect 1023 3691 1032 3692
rect 1023 3687 1024 3691
rect 1031 3687 1032 3691
rect 1086 3688 1087 3692
rect 1091 3688 1092 3692
rect 1086 3687 1092 3688
rect 1183 3691 1192 3692
rect 1183 3687 1184 3691
rect 1191 3687 1192 3691
rect 1254 3688 1255 3692
rect 1259 3688 1260 3692
rect 1254 3687 1260 3688
rect 1346 3691 1357 3692
rect 1346 3687 1347 3691
rect 1351 3687 1352 3691
rect 1356 3687 1357 3691
rect 1422 3688 1423 3692
rect 1427 3688 1428 3692
rect 1422 3687 1428 3688
rect 1519 3691 1528 3692
rect 1519 3687 1520 3691
rect 1527 3687 1528 3691
rect 1590 3688 1591 3692
rect 1595 3688 1596 3692
rect 1590 3687 1596 3688
rect 1687 3691 1696 3692
rect 1687 3687 1688 3691
rect 1695 3687 1696 3691
rect 1758 3688 1759 3692
rect 1763 3688 1764 3692
rect 1758 3687 1764 3688
rect 1854 3691 1861 3692
rect 1854 3687 1855 3691
rect 1860 3687 1861 3691
rect 1934 3689 1935 3693
rect 1939 3689 1940 3693
rect 1934 3688 1940 3689
rect 3838 3689 3844 3690
rect 5662 3689 5668 3690
rect 887 3686 893 3687
rect 1023 3686 1032 3687
rect 1183 3686 1192 3687
rect 1346 3686 1357 3687
rect 1519 3686 1528 3687
rect 1687 3686 1696 3687
rect 1854 3686 1861 3687
rect 2938 3687 2944 3688
rect 2938 3683 2939 3687
rect 2943 3686 2944 3687
rect 3590 3687 3596 3688
rect 3590 3686 3591 3687
rect 2943 3684 3591 3686
rect 2943 3683 2944 3684
rect 2938 3682 2944 3683
rect 3590 3683 3591 3684
rect 3595 3683 3596 3687
rect 3838 3685 3839 3689
rect 3843 3685 3844 3689
rect 3838 3684 3844 3685
rect 3886 3688 3892 3689
rect 4054 3688 4060 3689
rect 4246 3688 4252 3689
rect 4438 3688 4444 3689
rect 4630 3688 4636 3689
rect 3886 3684 3887 3688
rect 3891 3684 3892 3688
rect 3886 3683 3892 3684
rect 3982 3687 3989 3688
rect 3982 3683 3983 3687
rect 3988 3683 3989 3687
rect 4054 3684 4055 3688
rect 4059 3684 4060 3688
rect 4054 3683 4060 3684
rect 4151 3687 4157 3688
rect 4151 3683 4152 3687
rect 4156 3686 4157 3687
rect 4182 3687 4188 3688
rect 4182 3686 4183 3687
rect 4156 3684 4183 3686
rect 4156 3683 4157 3684
rect 3590 3682 3596 3683
rect 3982 3682 3989 3683
rect 4151 3682 4157 3683
rect 4182 3683 4183 3684
rect 4187 3683 4188 3687
rect 4246 3684 4247 3688
rect 4251 3684 4252 3688
rect 4246 3683 4252 3684
rect 4343 3687 4349 3688
rect 4343 3683 4344 3687
rect 4348 3686 4349 3687
rect 4367 3687 4373 3688
rect 4367 3686 4368 3687
rect 4348 3684 4368 3686
rect 4348 3683 4349 3684
rect 4182 3682 4188 3683
rect 4343 3682 4349 3683
rect 4367 3683 4368 3684
rect 4372 3683 4373 3687
rect 4438 3684 4439 3688
rect 4443 3684 4444 3688
rect 4438 3683 4444 3684
rect 4535 3687 4541 3688
rect 4535 3683 4536 3687
rect 4540 3686 4541 3687
rect 4566 3687 4572 3688
rect 4566 3686 4567 3687
rect 4540 3684 4567 3686
rect 4540 3683 4541 3684
rect 4367 3682 4373 3683
rect 4535 3682 4541 3683
rect 4566 3683 4567 3684
rect 4571 3683 4572 3687
rect 4630 3684 4631 3688
rect 4635 3684 4636 3688
rect 4630 3683 4636 3684
rect 4722 3687 4733 3688
rect 4722 3683 4723 3687
rect 4727 3683 4728 3687
rect 4732 3683 4733 3687
rect 5662 3685 5663 3689
rect 5667 3685 5668 3689
rect 5662 3684 5668 3685
rect 4566 3682 4572 3683
rect 4722 3682 4733 3683
rect 602 3677 608 3678
rect 110 3676 116 3677
rect 110 3672 111 3676
rect 115 3672 116 3676
rect 602 3673 603 3677
rect 607 3673 608 3677
rect 602 3672 608 3673
rect 746 3677 752 3678
rect 746 3673 747 3677
rect 751 3673 752 3677
rect 746 3672 752 3673
rect 898 3677 904 3678
rect 898 3673 899 3677
rect 903 3673 904 3677
rect 898 3672 904 3673
rect 1058 3677 1064 3678
rect 1058 3673 1059 3677
rect 1063 3673 1064 3677
rect 1058 3672 1064 3673
rect 1226 3677 1232 3678
rect 1226 3673 1227 3677
rect 1231 3673 1232 3677
rect 1226 3672 1232 3673
rect 1394 3677 1400 3678
rect 1394 3673 1395 3677
rect 1399 3673 1400 3677
rect 1394 3672 1400 3673
rect 1562 3677 1568 3678
rect 1562 3673 1563 3677
rect 1567 3673 1568 3677
rect 1562 3672 1568 3673
rect 1730 3677 1736 3678
rect 1730 3673 1731 3677
rect 1735 3673 1736 3677
rect 1730 3672 1736 3673
rect 1934 3676 1940 3677
rect 1934 3672 1935 3676
rect 1939 3672 1940 3676
rect 3858 3673 3864 3674
rect 110 3671 116 3672
rect 1934 3671 1940 3672
rect 3838 3672 3844 3673
rect 3838 3668 3839 3672
rect 3843 3668 3844 3672
rect 3858 3669 3859 3673
rect 3863 3669 3864 3673
rect 3858 3668 3864 3669
rect 4026 3673 4032 3674
rect 4026 3669 4027 3673
rect 4031 3669 4032 3673
rect 4026 3668 4032 3669
rect 4218 3673 4224 3674
rect 4218 3669 4219 3673
rect 4223 3669 4224 3673
rect 4218 3668 4224 3669
rect 4410 3673 4416 3674
rect 4410 3669 4411 3673
rect 4415 3669 4416 3673
rect 4410 3668 4416 3669
rect 4602 3673 4608 3674
rect 4602 3669 4603 3673
rect 4607 3669 4608 3673
rect 4602 3668 4608 3669
rect 5662 3672 5668 3673
rect 5662 3668 5663 3672
rect 5667 3668 5668 3672
rect 3838 3667 3844 3668
rect 5662 3667 5668 3668
rect 2638 3659 2644 3660
rect 2476 3650 2478 3657
rect 2638 3655 2639 3659
rect 2643 3655 2644 3659
rect 2638 3654 2644 3655
rect 2938 3659 2944 3660
rect 2938 3655 2939 3659
rect 2943 3655 2944 3659
rect 2938 3654 2944 3655
rect 2970 3659 2976 3660
rect 2970 3655 2971 3659
rect 2975 3658 2976 3659
rect 3186 3659 3192 3660
rect 2975 3656 3065 3658
rect 2975 3655 2976 3656
rect 2970 3654 2976 3655
rect 3186 3655 3187 3659
rect 3191 3658 3192 3659
rect 3982 3659 3988 3660
rect 3982 3658 3983 3659
rect 3191 3656 3273 3658
rect 3565 3656 3621 3658
rect 3749 3656 3983 3658
rect 3191 3655 3192 3656
rect 3186 3654 3192 3655
rect 2742 3651 2748 3652
rect 2742 3650 2743 3651
rect 2476 3648 2743 3650
rect 2742 3647 2743 3648
rect 2747 3647 2748 3651
rect 3619 3650 3621 3656
rect 3982 3655 3983 3656
rect 3987 3655 3988 3659
rect 3982 3654 3988 3655
rect 3770 3651 3776 3652
rect 3770 3650 3771 3651
rect 3619 3648 3771 3650
rect 2742 3646 2748 3647
rect 3770 3647 3771 3648
rect 3775 3647 3776 3651
rect 3770 3646 3776 3647
rect 698 3627 704 3628
rect 698 3623 699 3627
rect 703 3623 704 3627
rect 698 3622 704 3623
rect 730 3627 736 3628
rect 730 3623 731 3627
rect 735 3626 736 3627
rect 887 3627 893 3628
rect 735 3624 753 3626
rect 735 3623 736 3624
rect 730 3622 736 3623
rect 887 3623 888 3627
rect 892 3626 893 3627
rect 1026 3627 1032 3628
rect 892 3624 905 3626
rect 892 3623 893 3624
rect 887 3622 893 3623
rect 1026 3623 1027 3627
rect 1031 3626 1032 3627
rect 1186 3627 1192 3628
rect 1031 3624 1065 3626
rect 1031 3623 1032 3624
rect 1026 3622 1032 3623
rect 1186 3623 1187 3627
rect 1191 3626 1192 3627
rect 1522 3627 1528 3628
rect 1191 3624 1233 3626
rect 1191 3623 1192 3624
rect 1186 3622 1192 3623
rect 1492 3618 1494 3625
rect 1522 3623 1523 3627
rect 1527 3626 1528 3627
rect 1690 3627 1696 3628
rect 1527 3624 1569 3626
rect 1527 3623 1528 3624
rect 1522 3622 1528 3623
rect 1690 3623 1691 3627
rect 1695 3626 1696 3627
rect 1695 3624 1737 3626
rect 1695 3623 1696 3624
rect 1690 3622 1696 3623
rect 3954 3623 3960 3624
rect 1850 3619 1856 3620
rect 1850 3618 1851 3619
rect 1492 3616 1851 3618
rect 1850 3615 1851 3616
rect 1855 3615 1856 3619
rect 1850 3614 1856 3615
rect 2502 3619 2508 3620
rect 2502 3615 2503 3619
rect 2507 3615 2508 3619
rect 3954 3619 3955 3623
rect 3959 3619 3960 3623
rect 4170 3623 4176 3624
rect 4170 3622 4171 3623
rect 4125 3620 4171 3622
rect 3954 3618 3960 3619
rect 4170 3619 4171 3620
rect 4175 3619 4176 3623
rect 4170 3618 4176 3619
rect 4182 3623 4188 3624
rect 4182 3619 4183 3623
rect 4187 3622 4188 3623
rect 4367 3623 4373 3624
rect 4187 3620 4225 3622
rect 4187 3619 4188 3620
rect 4182 3618 4188 3619
rect 4367 3619 4368 3623
rect 4372 3622 4373 3623
rect 4566 3623 4572 3624
rect 4372 3620 4417 3622
rect 4372 3619 4373 3620
rect 4367 3618 4373 3619
rect 4566 3619 4567 3623
rect 4571 3622 4572 3623
rect 4571 3620 4609 3622
rect 4571 3619 4572 3620
rect 4566 3618 4572 3619
rect 2502 3614 2508 3615
rect 2554 3615 2560 3616
rect 2554 3611 2555 3615
rect 2559 3611 2560 3615
rect 2554 3610 2560 3611
rect 2690 3615 2696 3616
rect 2690 3611 2691 3615
rect 2695 3611 2696 3615
rect 2690 3610 2696 3611
rect 4722 3599 4728 3600
rect 4722 3598 4723 3599
rect 4672 3596 4723 3598
rect 1346 3591 1352 3592
rect 1346 3590 1347 3591
rect 916 3588 1347 3590
rect 916 3582 918 3588
rect 1346 3587 1347 3588
rect 1351 3587 1352 3591
rect 1346 3586 1352 3587
rect 1370 3591 1376 3592
rect 1370 3587 1371 3591
rect 1375 3590 1376 3591
rect 1463 3591 1469 3592
rect 1463 3590 1464 3591
rect 1375 3588 1464 3590
rect 1375 3587 1376 3588
rect 1370 3586 1376 3587
rect 1463 3587 1464 3588
rect 1468 3587 1469 3591
rect 1463 3586 1469 3587
rect 3778 3591 3784 3592
rect 3778 3587 3779 3591
rect 3783 3590 3784 3591
rect 4672 3590 4674 3596
rect 4722 3595 4723 3596
rect 4727 3595 4728 3599
rect 4722 3594 4728 3595
rect 3783 3588 3865 3590
rect 4637 3588 4674 3590
rect 3783 3587 3784 3588
rect 3778 3586 3784 3587
rect 4002 3587 4008 3588
rect 4002 3583 4003 3587
rect 4007 3583 4008 3587
rect 4002 3582 4008 3583
rect 4138 3587 4144 3588
rect 4138 3583 4139 3587
rect 4143 3583 4144 3587
rect 4138 3582 4144 3583
rect 4274 3587 4280 3588
rect 4274 3583 4275 3587
rect 4279 3583 4280 3587
rect 4274 3582 4280 3583
rect 4410 3587 4416 3588
rect 4410 3583 4411 3587
rect 4415 3583 4416 3587
rect 4410 3582 4416 3583
rect 4682 3587 4688 3588
rect 4682 3583 4683 3587
rect 4687 3583 4688 3587
rect 4682 3582 4688 3583
rect 4818 3587 4824 3588
rect 4818 3583 4819 3587
rect 4823 3583 4824 3587
rect 4818 3582 4824 3583
rect 4954 3587 4960 3588
rect 4954 3583 4955 3587
rect 4959 3583 4960 3587
rect 4954 3582 4960 3583
rect 5090 3587 5096 3588
rect 5090 3583 5091 3587
rect 5095 3583 5096 3587
rect 5090 3582 5096 3583
rect 877 3580 918 3582
rect 922 3579 928 3580
rect 922 3575 923 3579
rect 927 3575 928 3579
rect 922 3574 928 3575
rect 1058 3579 1064 3580
rect 1058 3575 1059 3579
rect 1063 3575 1064 3579
rect 1058 3574 1064 3575
rect 1194 3579 1200 3580
rect 1194 3575 1195 3579
rect 1199 3575 1200 3579
rect 1194 3574 1200 3575
rect 1330 3579 1336 3580
rect 1330 3575 1331 3579
rect 1335 3575 1336 3579
rect 1330 3574 1336 3575
rect 1602 3579 1608 3580
rect 1602 3575 1603 3579
rect 1607 3575 1608 3579
rect 1602 3574 1608 3575
rect 1738 3579 1744 3580
rect 1738 3575 1739 3579
rect 1743 3575 1744 3579
rect 1738 3574 1744 3575
rect 1974 3568 1980 3569
rect 3798 3568 3804 3569
rect 1974 3564 1975 3568
rect 1979 3564 1980 3568
rect 1974 3563 1980 3564
rect 2410 3567 2416 3568
rect 2410 3563 2411 3567
rect 2415 3563 2416 3567
rect 2410 3562 2416 3563
rect 2546 3567 2552 3568
rect 2546 3563 2547 3567
rect 2551 3563 2552 3567
rect 2546 3562 2552 3563
rect 2682 3567 2688 3568
rect 2682 3563 2683 3567
rect 2687 3563 2688 3567
rect 3798 3564 3799 3568
rect 3803 3564 3804 3568
rect 3798 3563 3804 3564
rect 2682 3562 2688 3563
rect 2438 3552 2444 3553
rect 2574 3552 2580 3553
rect 2710 3552 2716 3553
rect 1974 3551 1980 3552
rect 1974 3547 1975 3551
rect 1979 3547 1980 3551
rect 2438 3548 2439 3552
rect 2443 3548 2444 3552
rect 2438 3547 2444 3548
rect 2535 3551 2541 3552
rect 2535 3547 2536 3551
rect 2540 3550 2541 3551
rect 2554 3551 2560 3552
rect 2554 3550 2555 3551
rect 2540 3548 2555 3550
rect 2540 3547 2541 3548
rect 1974 3546 1980 3547
rect 2535 3546 2541 3547
rect 2554 3547 2555 3548
rect 2559 3547 2560 3551
rect 2574 3548 2575 3552
rect 2579 3548 2580 3552
rect 2574 3547 2580 3548
rect 2671 3551 2677 3552
rect 2671 3547 2672 3551
rect 2676 3550 2677 3551
rect 2690 3551 2696 3552
rect 2690 3550 2691 3551
rect 2676 3548 2691 3550
rect 2676 3547 2677 3548
rect 2554 3546 2560 3547
rect 2671 3546 2677 3547
rect 2690 3547 2691 3548
rect 2695 3547 2696 3551
rect 2710 3548 2711 3552
rect 2715 3548 2716 3552
rect 2710 3547 2716 3548
rect 2806 3551 2813 3552
rect 2806 3547 2807 3551
rect 2812 3547 2813 3551
rect 2690 3546 2696 3547
rect 2806 3546 2813 3547
rect 3798 3551 3804 3552
rect 3798 3547 3799 3551
rect 3803 3547 3804 3551
rect 3798 3546 3804 3547
rect 3838 3540 3844 3541
rect 5662 3540 5668 3541
rect 3838 3536 3839 3540
rect 3843 3536 3844 3540
rect 3838 3535 3844 3536
rect 3858 3539 3864 3540
rect 3858 3535 3859 3539
rect 3863 3535 3864 3539
rect 3858 3534 3864 3535
rect 3994 3539 4000 3540
rect 3994 3535 3995 3539
rect 3999 3535 4000 3539
rect 3994 3534 4000 3535
rect 4130 3539 4136 3540
rect 4130 3535 4131 3539
rect 4135 3535 4136 3539
rect 4130 3534 4136 3535
rect 4266 3539 4272 3540
rect 4266 3535 4267 3539
rect 4271 3535 4272 3539
rect 4266 3534 4272 3535
rect 4402 3539 4408 3540
rect 4402 3535 4403 3539
rect 4407 3535 4408 3539
rect 4402 3534 4408 3535
rect 4538 3539 4544 3540
rect 4538 3535 4539 3539
rect 4543 3535 4544 3539
rect 4538 3534 4544 3535
rect 4674 3539 4680 3540
rect 4674 3535 4675 3539
rect 4679 3535 4680 3539
rect 4674 3534 4680 3535
rect 4810 3539 4816 3540
rect 4810 3535 4811 3539
rect 4815 3535 4816 3539
rect 4810 3534 4816 3535
rect 4946 3539 4952 3540
rect 4946 3535 4947 3539
rect 4951 3535 4952 3539
rect 4946 3534 4952 3535
rect 5082 3539 5088 3540
rect 5082 3535 5083 3539
rect 5087 3535 5088 3539
rect 5662 3536 5663 3540
rect 5667 3536 5668 3540
rect 5662 3535 5668 3536
rect 5082 3534 5088 3535
rect 110 3532 116 3533
rect 1934 3532 1940 3533
rect 110 3528 111 3532
rect 115 3528 116 3532
rect 110 3527 116 3528
rect 778 3531 784 3532
rect 778 3527 779 3531
rect 783 3527 784 3531
rect 778 3526 784 3527
rect 914 3531 920 3532
rect 914 3527 915 3531
rect 919 3527 920 3531
rect 914 3526 920 3527
rect 1050 3531 1056 3532
rect 1050 3527 1051 3531
rect 1055 3527 1056 3531
rect 1050 3526 1056 3527
rect 1186 3531 1192 3532
rect 1186 3527 1187 3531
rect 1191 3527 1192 3531
rect 1186 3526 1192 3527
rect 1322 3531 1328 3532
rect 1322 3527 1323 3531
rect 1327 3527 1328 3531
rect 1322 3526 1328 3527
rect 1458 3531 1464 3532
rect 1458 3527 1459 3531
rect 1463 3527 1464 3531
rect 1458 3526 1464 3527
rect 1594 3531 1600 3532
rect 1594 3527 1595 3531
rect 1599 3527 1600 3531
rect 1594 3526 1600 3527
rect 1730 3531 1736 3532
rect 1730 3527 1731 3531
rect 1735 3527 1736 3531
rect 1934 3528 1935 3532
rect 1939 3528 1940 3532
rect 1934 3527 1940 3528
rect 1730 3526 1736 3527
rect 3886 3524 3892 3525
rect 4022 3524 4028 3525
rect 4158 3524 4164 3525
rect 4294 3524 4300 3525
rect 4430 3524 4436 3525
rect 4566 3524 4572 3525
rect 4702 3524 4708 3525
rect 4838 3524 4844 3525
rect 4974 3524 4980 3525
rect 5110 3524 5116 3525
rect 3838 3523 3844 3524
rect 3838 3519 3839 3523
rect 3843 3519 3844 3523
rect 3886 3520 3887 3524
rect 3891 3520 3892 3524
rect 3886 3519 3892 3520
rect 3983 3523 3989 3524
rect 3983 3519 3984 3523
rect 3988 3522 3989 3523
rect 4002 3523 4008 3524
rect 4002 3522 4003 3523
rect 3988 3520 4003 3522
rect 3988 3519 3989 3520
rect 3838 3518 3844 3519
rect 3983 3518 3989 3519
rect 4002 3519 4003 3520
rect 4007 3519 4008 3523
rect 4022 3520 4023 3524
rect 4027 3520 4028 3524
rect 4022 3519 4028 3520
rect 4119 3523 4125 3524
rect 4119 3519 4120 3523
rect 4124 3522 4125 3523
rect 4138 3523 4144 3524
rect 4138 3522 4139 3523
rect 4124 3520 4139 3522
rect 4124 3519 4125 3520
rect 4002 3518 4008 3519
rect 4119 3518 4125 3519
rect 4138 3519 4139 3520
rect 4143 3519 4144 3523
rect 4158 3520 4159 3524
rect 4163 3520 4164 3524
rect 4158 3519 4164 3520
rect 4255 3523 4261 3524
rect 4255 3519 4256 3523
rect 4260 3522 4261 3523
rect 4274 3523 4280 3524
rect 4274 3522 4275 3523
rect 4260 3520 4275 3522
rect 4260 3519 4261 3520
rect 4138 3518 4144 3519
rect 4255 3518 4261 3519
rect 4274 3519 4275 3520
rect 4279 3519 4280 3523
rect 4294 3520 4295 3524
rect 4299 3520 4300 3524
rect 4294 3519 4300 3520
rect 4391 3523 4397 3524
rect 4391 3519 4392 3523
rect 4396 3522 4397 3523
rect 4410 3523 4416 3524
rect 4410 3522 4411 3523
rect 4396 3520 4411 3522
rect 4396 3519 4397 3520
rect 4274 3518 4280 3519
rect 4391 3518 4397 3519
rect 4410 3519 4411 3520
rect 4415 3519 4416 3523
rect 4430 3520 4431 3524
rect 4435 3520 4436 3524
rect 4430 3519 4436 3520
rect 4526 3523 4533 3524
rect 4526 3519 4527 3523
rect 4532 3519 4533 3523
rect 4566 3520 4567 3524
rect 4571 3520 4572 3524
rect 4566 3519 4572 3520
rect 4663 3523 4669 3524
rect 4663 3519 4664 3523
rect 4668 3522 4669 3523
rect 4682 3523 4688 3524
rect 4682 3522 4683 3523
rect 4668 3520 4683 3522
rect 4668 3519 4669 3520
rect 4410 3518 4416 3519
rect 4526 3518 4533 3519
rect 4663 3518 4669 3519
rect 4682 3519 4683 3520
rect 4687 3519 4688 3523
rect 4702 3520 4703 3524
rect 4707 3520 4708 3524
rect 4702 3519 4708 3520
rect 4799 3523 4805 3524
rect 4799 3519 4800 3523
rect 4804 3522 4805 3523
rect 4818 3523 4824 3524
rect 4818 3522 4819 3523
rect 4804 3520 4819 3522
rect 4804 3519 4805 3520
rect 4682 3518 4688 3519
rect 4799 3518 4805 3519
rect 4818 3519 4819 3520
rect 4823 3519 4824 3523
rect 4838 3520 4839 3524
rect 4843 3520 4844 3524
rect 4838 3519 4844 3520
rect 4935 3523 4941 3524
rect 4935 3519 4936 3523
rect 4940 3522 4941 3523
rect 4954 3523 4960 3524
rect 4954 3522 4955 3523
rect 4940 3520 4955 3522
rect 4940 3519 4941 3520
rect 4818 3518 4824 3519
rect 4935 3518 4941 3519
rect 4954 3519 4955 3520
rect 4959 3519 4960 3523
rect 4974 3520 4975 3524
rect 4979 3520 4980 3524
rect 4974 3519 4980 3520
rect 5071 3523 5077 3524
rect 5071 3519 5072 3523
rect 5076 3522 5077 3523
rect 5090 3523 5096 3524
rect 5090 3522 5091 3523
rect 5076 3520 5091 3522
rect 5076 3519 5077 3520
rect 4954 3518 4960 3519
rect 5071 3518 5077 3519
rect 5090 3519 5091 3520
rect 5095 3519 5096 3523
rect 5110 3520 5111 3524
rect 5115 3520 5116 3524
rect 5110 3519 5116 3520
rect 5206 3523 5213 3524
rect 5206 3519 5207 3523
rect 5212 3519 5213 3523
rect 5090 3518 5096 3519
rect 5206 3518 5213 3519
rect 5662 3523 5668 3524
rect 5662 3519 5663 3523
rect 5667 3519 5668 3523
rect 5662 3518 5668 3519
rect 806 3516 812 3517
rect 942 3516 948 3517
rect 1078 3516 1084 3517
rect 1214 3516 1220 3517
rect 1350 3516 1356 3517
rect 1486 3516 1492 3517
rect 1622 3516 1628 3517
rect 1758 3516 1764 3517
rect 110 3515 116 3516
rect 110 3511 111 3515
rect 115 3511 116 3515
rect 806 3512 807 3516
rect 811 3512 812 3516
rect 806 3511 812 3512
rect 903 3515 909 3516
rect 903 3511 904 3515
rect 908 3514 909 3515
rect 922 3515 928 3516
rect 922 3514 923 3515
rect 908 3512 923 3514
rect 908 3511 909 3512
rect 110 3510 116 3511
rect 903 3510 909 3511
rect 922 3511 923 3512
rect 927 3511 928 3515
rect 942 3512 943 3516
rect 947 3512 948 3516
rect 942 3511 948 3512
rect 1039 3515 1045 3516
rect 1039 3511 1040 3515
rect 1044 3514 1045 3515
rect 1058 3515 1064 3516
rect 1058 3514 1059 3515
rect 1044 3512 1059 3514
rect 1044 3511 1045 3512
rect 922 3510 928 3511
rect 1039 3510 1045 3511
rect 1058 3511 1059 3512
rect 1063 3511 1064 3515
rect 1078 3512 1079 3516
rect 1083 3512 1084 3516
rect 1078 3511 1084 3512
rect 1175 3515 1181 3516
rect 1175 3511 1176 3515
rect 1180 3514 1181 3515
rect 1194 3515 1200 3516
rect 1194 3514 1195 3515
rect 1180 3512 1195 3514
rect 1180 3511 1181 3512
rect 1058 3510 1064 3511
rect 1175 3510 1181 3511
rect 1194 3511 1195 3512
rect 1199 3511 1200 3515
rect 1214 3512 1215 3516
rect 1219 3512 1220 3516
rect 1214 3511 1220 3512
rect 1311 3515 1317 3516
rect 1311 3511 1312 3515
rect 1316 3514 1317 3515
rect 1330 3515 1336 3516
rect 1330 3514 1331 3515
rect 1316 3512 1331 3514
rect 1316 3511 1317 3512
rect 1194 3510 1200 3511
rect 1311 3510 1317 3511
rect 1330 3511 1331 3512
rect 1335 3511 1336 3515
rect 1350 3512 1351 3516
rect 1355 3512 1356 3516
rect 1350 3511 1356 3512
rect 1446 3515 1453 3516
rect 1446 3511 1447 3515
rect 1452 3511 1453 3515
rect 1486 3512 1487 3516
rect 1491 3512 1492 3516
rect 1486 3511 1492 3512
rect 1583 3515 1589 3516
rect 1583 3511 1584 3515
rect 1588 3514 1589 3515
rect 1602 3515 1608 3516
rect 1602 3514 1603 3515
rect 1588 3512 1603 3514
rect 1588 3511 1589 3512
rect 1330 3510 1336 3511
rect 1446 3510 1453 3511
rect 1583 3510 1589 3511
rect 1602 3511 1603 3512
rect 1607 3511 1608 3515
rect 1622 3512 1623 3516
rect 1627 3512 1628 3516
rect 1622 3511 1628 3512
rect 1719 3515 1725 3516
rect 1719 3511 1720 3515
rect 1724 3514 1725 3515
rect 1738 3515 1744 3516
rect 1738 3514 1739 3515
rect 1724 3512 1739 3514
rect 1724 3511 1725 3512
rect 1602 3510 1608 3511
rect 1719 3510 1725 3511
rect 1738 3511 1739 3512
rect 1743 3511 1744 3515
rect 1758 3512 1759 3516
rect 1763 3512 1764 3516
rect 1758 3511 1764 3512
rect 1850 3515 1861 3516
rect 1850 3511 1851 3515
rect 1855 3511 1856 3515
rect 1860 3511 1861 3515
rect 1738 3510 1744 3511
rect 1850 3510 1861 3511
rect 1934 3515 1940 3516
rect 1934 3511 1935 3515
rect 1939 3511 1940 3515
rect 1934 3510 1940 3511
rect 4898 3487 4904 3488
rect 4898 3483 4899 3487
rect 4903 3486 4904 3487
rect 5206 3487 5212 3488
rect 5206 3486 5207 3487
rect 4903 3484 5207 3486
rect 4903 3483 4904 3484
rect 4898 3482 4904 3483
rect 5206 3483 5207 3484
rect 5211 3483 5212 3487
rect 5206 3482 5212 3483
rect 3838 3457 3844 3458
rect 5662 3457 5668 3458
rect 1974 3453 1980 3454
rect 3798 3453 3804 3454
rect 1974 3449 1975 3453
rect 1979 3449 1980 3453
rect 1974 3448 1980 3449
rect 2598 3452 2604 3453
rect 2822 3452 2828 3453
rect 3046 3452 3052 3453
rect 3262 3452 3268 3453
rect 3478 3452 3484 3453
rect 3678 3452 3684 3453
rect 2598 3448 2599 3452
rect 2603 3448 2604 3452
rect 2598 3447 2604 3448
rect 2695 3451 2704 3452
rect 2695 3447 2696 3451
rect 2703 3447 2704 3451
rect 2822 3448 2823 3452
rect 2827 3448 2828 3452
rect 2822 3447 2828 3448
rect 2914 3451 2925 3452
rect 2914 3447 2915 3451
rect 2919 3447 2920 3451
rect 2924 3447 2925 3451
rect 3046 3448 3047 3452
rect 3051 3448 3052 3452
rect 3046 3447 3052 3448
rect 3143 3451 3152 3452
rect 3143 3447 3144 3451
rect 3151 3447 3152 3451
rect 3262 3448 3263 3452
rect 3267 3448 3268 3452
rect 3262 3447 3268 3448
rect 3359 3451 3368 3452
rect 3359 3447 3360 3451
rect 3367 3447 3368 3451
rect 3478 3448 3479 3452
rect 3483 3448 3484 3452
rect 3478 3447 3484 3448
rect 3575 3451 3581 3452
rect 3575 3447 3576 3451
rect 3580 3450 3581 3451
rect 3598 3451 3604 3452
rect 3598 3450 3599 3451
rect 3580 3448 3599 3450
rect 3580 3447 3581 3448
rect 2695 3446 2704 3447
rect 2914 3446 2925 3447
rect 3143 3446 3152 3447
rect 3359 3446 3368 3447
rect 3575 3446 3581 3447
rect 3598 3447 3599 3448
rect 3603 3447 3604 3451
rect 3678 3448 3679 3452
rect 3683 3448 3684 3452
rect 3678 3447 3684 3448
rect 3775 3451 3784 3452
rect 3775 3447 3776 3451
rect 3783 3447 3784 3451
rect 3798 3449 3799 3453
rect 3803 3449 3804 3453
rect 3838 3453 3839 3457
rect 3843 3453 3844 3457
rect 3838 3452 3844 3453
rect 4830 3456 4836 3457
rect 4966 3456 4972 3457
rect 5102 3456 5108 3457
rect 5238 3456 5244 3457
rect 5374 3456 5380 3457
rect 4830 3452 4831 3456
rect 4835 3452 4836 3456
rect 4830 3451 4836 3452
rect 4927 3455 4936 3456
rect 4927 3451 4928 3455
rect 4935 3451 4936 3455
rect 4966 3452 4967 3456
rect 4971 3452 4972 3456
rect 4966 3451 4972 3452
rect 5063 3455 5072 3456
rect 5063 3451 5064 3455
rect 5071 3451 5072 3455
rect 5102 3452 5103 3456
rect 5107 3452 5108 3456
rect 5102 3451 5108 3452
rect 5199 3455 5208 3456
rect 5199 3451 5200 3455
rect 5207 3451 5208 3455
rect 5238 3452 5239 3456
rect 5243 3452 5244 3456
rect 5238 3451 5244 3452
rect 5335 3455 5344 3456
rect 5335 3451 5336 3455
rect 5343 3451 5344 3455
rect 5374 3452 5375 3456
rect 5379 3452 5380 3456
rect 5374 3451 5380 3452
rect 5470 3455 5477 3456
rect 5470 3451 5471 3455
rect 5476 3451 5477 3455
rect 5662 3453 5663 3457
rect 5667 3453 5668 3457
rect 5662 3452 5668 3453
rect 4927 3450 4936 3451
rect 5063 3450 5072 3451
rect 5199 3450 5208 3451
rect 5335 3450 5344 3451
rect 5470 3450 5477 3451
rect 3798 3448 3804 3449
rect 3598 3446 3604 3447
rect 3775 3446 3784 3447
rect 4802 3441 4808 3442
rect 3838 3440 3844 3441
rect 2570 3437 2576 3438
rect 1974 3436 1980 3437
rect 110 3433 116 3434
rect 1934 3433 1940 3434
rect 110 3429 111 3433
rect 115 3429 116 3433
rect 110 3428 116 3429
rect 726 3432 732 3433
rect 862 3432 868 3433
rect 998 3432 1004 3433
rect 1134 3432 1140 3433
rect 1270 3432 1276 3433
rect 1406 3432 1412 3433
rect 1542 3432 1548 3433
rect 1678 3432 1684 3433
rect 1814 3432 1820 3433
rect 726 3428 727 3432
rect 731 3428 732 3432
rect 726 3427 732 3428
rect 823 3431 832 3432
rect 823 3427 824 3431
rect 831 3427 832 3431
rect 862 3428 863 3432
rect 867 3428 868 3432
rect 862 3427 868 3428
rect 959 3431 968 3432
rect 959 3427 960 3431
rect 967 3427 968 3431
rect 998 3428 999 3432
rect 1003 3428 1004 3432
rect 998 3427 1004 3428
rect 1095 3431 1101 3432
rect 1095 3427 1096 3431
rect 1100 3430 1101 3431
rect 1103 3431 1109 3432
rect 1103 3430 1104 3431
rect 1100 3428 1104 3430
rect 1100 3427 1101 3428
rect 823 3426 832 3427
rect 959 3426 968 3427
rect 1095 3426 1101 3427
rect 1103 3427 1104 3428
rect 1108 3427 1109 3431
rect 1134 3428 1135 3432
rect 1139 3428 1140 3432
rect 1134 3427 1140 3428
rect 1231 3431 1240 3432
rect 1231 3427 1232 3431
rect 1239 3427 1240 3431
rect 1270 3428 1271 3432
rect 1275 3428 1276 3432
rect 1270 3427 1276 3428
rect 1367 3431 1376 3432
rect 1367 3427 1368 3431
rect 1375 3427 1376 3431
rect 1406 3428 1407 3432
rect 1411 3428 1412 3432
rect 1406 3427 1412 3428
rect 1503 3431 1512 3432
rect 1503 3427 1504 3431
rect 1511 3427 1512 3431
rect 1542 3428 1543 3432
rect 1547 3428 1548 3432
rect 1542 3427 1548 3428
rect 1639 3431 1648 3432
rect 1639 3427 1640 3431
rect 1647 3427 1648 3431
rect 1678 3428 1679 3432
rect 1683 3428 1684 3432
rect 1678 3427 1684 3428
rect 1775 3431 1784 3432
rect 1775 3427 1776 3431
rect 1783 3427 1784 3431
rect 1814 3428 1815 3432
rect 1819 3428 1820 3432
rect 1814 3427 1820 3428
rect 1906 3431 1917 3432
rect 1906 3427 1907 3431
rect 1911 3427 1912 3431
rect 1916 3427 1917 3431
rect 1934 3429 1935 3433
rect 1939 3429 1940 3433
rect 1974 3432 1975 3436
rect 1979 3432 1980 3436
rect 2570 3433 2571 3437
rect 2575 3433 2576 3437
rect 2570 3432 2576 3433
rect 2794 3437 2800 3438
rect 2794 3433 2795 3437
rect 2799 3433 2800 3437
rect 2794 3432 2800 3433
rect 3018 3437 3024 3438
rect 3018 3433 3019 3437
rect 3023 3433 3024 3437
rect 3018 3432 3024 3433
rect 3234 3437 3240 3438
rect 3234 3433 3235 3437
rect 3239 3433 3240 3437
rect 3234 3432 3240 3433
rect 3450 3437 3456 3438
rect 3450 3433 3451 3437
rect 3455 3433 3456 3437
rect 3450 3432 3456 3433
rect 3650 3437 3656 3438
rect 3650 3433 3651 3437
rect 3655 3433 3656 3437
rect 3650 3432 3656 3433
rect 3798 3436 3804 3437
rect 3798 3432 3799 3436
rect 3803 3432 3804 3436
rect 3838 3436 3839 3440
rect 3843 3436 3844 3440
rect 4802 3437 4803 3441
rect 4807 3437 4808 3441
rect 4802 3436 4808 3437
rect 4938 3441 4944 3442
rect 4938 3437 4939 3441
rect 4943 3437 4944 3441
rect 4938 3436 4944 3437
rect 5074 3441 5080 3442
rect 5074 3437 5075 3441
rect 5079 3437 5080 3441
rect 5074 3436 5080 3437
rect 5210 3441 5216 3442
rect 5210 3437 5211 3441
rect 5215 3437 5216 3441
rect 5210 3436 5216 3437
rect 5346 3441 5352 3442
rect 5346 3437 5347 3441
rect 5351 3437 5352 3441
rect 5346 3436 5352 3437
rect 5662 3440 5668 3441
rect 5662 3436 5663 3440
rect 5667 3436 5668 3440
rect 3838 3435 3844 3436
rect 5662 3435 5668 3436
rect 1974 3431 1980 3432
rect 3798 3431 3804 3432
rect 1934 3428 1940 3429
rect 1103 3426 1109 3427
rect 1231 3426 1240 3427
rect 1367 3426 1376 3427
rect 1503 3426 1512 3427
rect 1639 3426 1648 3427
rect 1775 3426 1784 3427
rect 1906 3426 1917 3427
rect 698 3417 704 3418
rect 110 3416 116 3417
rect 110 3412 111 3416
rect 115 3412 116 3416
rect 698 3413 699 3417
rect 703 3413 704 3417
rect 698 3412 704 3413
rect 834 3417 840 3418
rect 834 3413 835 3417
rect 839 3413 840 3417
rect 834 3412 840 3413
rect 970 3417 976 3418
rect 970 3413 971 3417
rect 975 3413 976 3417
rect 970 3412 976 3413
rect 1106 3417 1112 3418
rect 1106 3413 1107 3417
rect 1111 3413 1112 3417
rect 1106 3412 1112 3413
rect 1242 3417 1248 3418
rect 1242 3413 1243 3417
rect 1247 3413 1248 3417
rect 1242 3412 1248 3413
rect 1378 3417 1384 3418
rect 1378 3413 1379 3417
rect 1383 3413 1384 3417
rect 1378 3412 1384 3413
rect 1514 3417 1520 3418
rect 1514 3413 1515 3417
rect 1519 3413 1520 3417
rect 1514 3412 1520 3413
rect 1650 3417 1656 3418
rect 1650 3413 1651 3417
rect 1655 3413 1656 3417
rect 1650 3412 1656 3413
rect 1786 3417 1792 3418
rect 1786 3413 1787 3417
rect 1791 3413 1792 3417
rect 1786 3412 1792 3413
rect 1934 3416 1940 3417
rect 1934 3412 1935 3416
rect 1939 3412 1940 3416
rect 110 3411 116 3412
rect 1934 3411 1940 3412
rect 4898 3391 4904 3392
rect 2806 3387 2812 3388
rect 2669 3384 2781 3386
rect 2779 3378 2781 3384
rect 2806 3383 2807 3387
rect 2811 3383 2812 3387
rect 2806 3382 2812 3383
rect 3114 3387 3120 3388
rect 3114 3383 3115 3387
rect 3119 3383 3120 3387
rect 3114 3382 3120 3383
rect 3146 3387 3152 3388
rect 3146 3383 3147 3387
rect 3151 3386 3152 3387
rect 3362 3387 3368 3388
rect 3151 3384 3241 3386
rect 3151 3383 3152 3384
rect 3146 3382 3152 3383
rect 3362 3383 3363 3387
rect 3367 3386 3368 3387
rect 3598 3387 3604 3388
rect 3367 3384 3457 3386
rect 3367 3383 3368 3384
rect 3362 3382 3368 3383
rect 3598 3383 3599 3387
rect 3603 3386 3604 3387
rect 4898 3387 4899 3391
rect 4903 3387 4904 3391
rect 4898 3386 4904 3387
rect 4930 3391 4936 3392
rect 4930 3387 4931 3391
rect 4935 3390 4936 3391
rect 5066 3391 5072 3392
rect 4935 3388 4945 3390
rect 4935 3387 4936 3388
rect 4930 3386 4936 3387
rect 5066 3387 5067 3391
rect 5071 3390 5072 3391
rect 5202 3391 5208 3392
rect 5071 3388 5081 3390
rect 5071 3387 5072 3388
rect 5066 3386 5072 3387
rect 5202 3387 5203 3391
rect 5207 3390 5208 3391
rect 5338 3391 5344 3392
rect 5207 3388 5217 3390
rect 5207 3387 5208 3388
rect 5202 3386 5208 3387
rect 5338 3387 5339 3391
rect 5343 3390 5344 3391
rect 5343 3388 5353 3390
rect 5343 3387 5344 3388
rect 5338 3386 5344 3387
rect 3603 3384 3657 3386
rect 3603 3383 3604 3384
rect 3598 3382 3604 3383
rect 2914 3379 2920 3380
rect 2914 3378 2915 3379
rect 2779 3376 2915 3378
rect 2914 3375 2915 3376
rect 2919 3375 2920 3379
rect 2914 3374 2920 3375
rect 826 3367 832 3368
rect 796 3358 798 3365
rect 826 3363 827 3367
rect 831 3366 832 3367
rect 962 3367 968 3368
rect 831 3364 841 3366
rect 831 3363 832 3364
rect 826 3362 832 3363
rect 962 3363 963 3367
rect 967 3366 968 3367
rect 1103 3367 1109 3368
rect 967 3364 977 3366
rect 967 3363 968 3364
rect 962 3362 968 3363
rect 1103 3363 1104 3367
rect 1108 3366 1109 3367
rect 1234 3367 1240 3368
rect 1108 3364 1113 3366
rect 1108 3363 1109 3364
rect 1103 3362 1109 3363
rect 1234 3363 1235 3367
rect 1239 3366 1240 3367
rect 1446 3367 1452 3368
rect 1239 3364 1249 3366
rect 1239 3363 1240 3364
rect 1234 3362 1240 3363
rect 1446 3363 1447 3367
rect 1451 3363 1452 3367
rect 1446 3362 1452 3363
rect 1506 3367 1512 3368
rect 1506 3363 1507 3367
rect 1511 3366 1512 3367
rect 1642 3367 1648 3368
rect 1511 3364 1521 3366
rect 1511 3363 1512 3364
rect 1506 3362 1512 3363
rect 1642 3363 1643 3367
rect 1647 3366 1648 3367
rect 1778 3367 1784 3368
rect 1647 3364 1657 3366
rect 1647 3363 1648 3364
rect 1642 3362 1648 3363
rect 1778 3363 1779 3367
rect 1783 3366 1784 3367
rect 1783 3364 1793 3366
rect 1783 3363 1784 3364
rect 1778 3362 1784 3363
rect 4262 3363 4268 3364
rect 4262 3362 4263 3363
rect 4136 3360 4263 3362
rect 874 3359 880 3360
rect 874 3358 875 3359
rect 796 3356 875 3358
rect 874 3355 875 3356
rect 879 3355 880 3359
rect 4136 3358 4138 3360
rect 4262 3359 4263 3360
rect 4267 3359 4268 3363
rect 5302 3363 5308 3364
rect 5302 3362 5303 3363
rect 4262 3358 4268 3359
rect 5120 3360 5303 3362
rect 5120 3358 5122 3360
rect 5302 3359 5303 3360
rect 5307 3359 5308 3363
rect 5302 3358 5308 3359
rect 5470 3359 5476 3360
rect 3957 3356 4138 3358
rect 5037 3356 5122 3358
rect 874 3354 880 3355
rect 4146 3355 4152 3356
rect 4146 3351 4147 3355
rect 4151 3351 4152 3355
rect 4146 3350 4152 3351
rect 4522 3355 4528 3356
rect 4522 3351 4523 3355
rect 4527 3351 4528 3355
rect 4522 3350 4528 3351
rect 4698 3355 4704 3356
rect 4698 3351 4699 3355
rect 4703 3351 4704 3355
rect 5470 3355 5471 3359
rect 5475 3355 5476 3359
rect 5470 3354 5476 3355
rect 4698 3350 4704 3351
rect 5272 3350 5274 3353
rect 5418 3351 5424 3352
rect 5418 3350 5419 3351
rect 5272 3348 5419 3350
rect 2679 3347 2685 3348
rect 2679 3346 2680 3347
rect 2629 3344 2680 3346
rect 2679 3343 2680 3344
rect 2684 3343 2685 3347
rect 2679 3342 2685 3343
rect 2698 3347 2704 3348
rect 2698 3343 2699 3347
rect 2703 3346 2704 3347
rect 3070 3347 3076 3348
rect 3070 3346 3071 3347
rect 2703 3344 2721 3346
rect 2997 3344 3071 3346
rect 2703 3343 2704 3344
rect 2698 3342 2704 3343
rect 3070 3343 3071 3344
rect 3075 3343 3076 3347
rect 5418 3347 5419 3348
rect 5423 3347 5424 3351
rect 5418 3346 5424 3347
rect 3070 3342 3076 3343
rect 3090 3343 3096 3344
rect 1158 3339 1164 3340
rect 1158 3338 1159 3339
rect 892 3336 1159 3338
rect 892 3330 894 3336
rect 1158 3335 1159 3336
rect 1163 3335 1164 3339
rect 3090 3339 3091 3343
rect 3095 3339 3096 3343
rect 3090 3338 3096 3339
rect 3274 3343 3280 3344
rect 3274 3339 3275 3343
rect 3279 3339 3280 3343
rect 3274 3338 3280 3339
rect 1158 3334 1164 3335
rect 1462 3335 1468 3336
rect 1462 3334 1463 3335
rect 1336 3332 1463 3334
rect 1018 3331 1024 3332
rect 1018 3330 1019 3331
rect 853 3328 894 3330
rect 989 3328 1019 3330
rect 1018 3327 1019 3328
rect 1023 3327 1024 3331
rect 1336 3330 1338 3332
rect 1462 3331 1463 3332
rect 1467 3331 1468 3335
rect 1906 3335 1912 3336
rect 1906 3334 1907 3335
rect 1462 3330 1468 3331
rect 1652 3332 1907 3334
rect 1652 3330 1654 3332
rect 1906 3331 1907 3332
rect 1911 3331 1912 3335
rect 1906 3330 1912 3331
rect 1285 3328 1338 3330
rect 1589 3328 1654 3330
rect 1018 3326 1024 3327
rect 1130 3327 1136 3328
rect 1130 3323 1131 3327
rect 1135 3323 1136 3327
rect 1130 3322 1136 3323
rect 1434 3327 1440 3328
rect 1434 3323 1435 3327
rect 1439 3323 1440 3327
rect 1434 3322 1440 3323
rect 1658 3327 1664 3328
rect 1658 3323 1659 3327
rect 1663 3323 1664 3327
rect 1658 3322 1664 3323
rect 1794 3327 1800 3328
rect 1794 3323 1795 3327
rect 1799 3323 1800 3327
rect 1794 3322 1800 3323
rect 3838 3308 3844 3309
rect 5662 3308 5668 3309
rect 3838 3304 3839 3308
rect 3843 3304 3844 3308
rect 3114 3303 3120 3304
rect 3838 3303 3844 3304
rect 3858 3307 3864 3308
rect 3858 3303 3859 3307
rect 3863 3303 3864 3307
rect 3114 3299 3115 3303
rect 3119 3302 3120 3303
rect 3858 3302 3864 3303
rect 4138 3307 4144 3308
rect 4138 3303 4139 3307
rect 4143 3303 4144 3307
rect 4138 3302 4144 3303
rect 4426 3307 4432 3308
rect 4426 3303 4427 3307
rect 4431 3303 4432 3307
rect 4426 3302 4432 3303
rect 4690 3307 4696 3308
rect 4690 3303 4691 3307
rect 4695 3303 4696 3307
rect 4690 3302 4696 3303
rect 4938 3307 4944 3308
rect 4938 3303 4939 3307
rect 4943 3303 4944 3307
rect 4938 3302 4944 3303
rect 5178 3307 5184 3308
rect 5178 3303 5179 3307
rect 5183 3303 5184 3307
rect 5178 3302 5184 3303
rect 5426 3307 5432 3308
rect 5426 3303 5427 3307
rect 5431 3303 5432 3307
rect 5662 3304 5663 3308
rect 5667 3304 5668 3308
rect 5662 3303 5668 3304
rect 5426 3302 5432 3303
rect 3119 3300 3834 3302
rect 3119 3299 3120 3300
rect 3114 3298 3120 3299
rect 3832 3298 3834 3300
rect 5418 3299 5424 3300
rect 1974 3296 1980 3297
rect 3798 3296 3804 3297
rect 3832 3296 3986 3298
rect 1974 3292 1975 3296
rect 1979 3292 1980 3296
rect 1974 3291 1980 3292
rect 2530 3295 2536 3296
rect 2530 3291 2531 3295
rect 2535 3291 2536 3295
rect 2530 3290 2536 3291
rect 2714 3295 2720 3296
rect 2714 3291 2715 3295
rect 2719 3291 2720 3295
rect 2714 3290 2720 3291
rect 2898 3295 2904 3296
rect 2898 3291 2899 3295
rect 2903 3291 2904 3295
rect 2898 3290 2904 3291
rect 3082 3295 3088 3296
rect 3082 3291 3083 3295
rect 3087 3291 3088 3295
rect 3082 3290 3088 3291
rect 3266 3295 3272 3296
rect 3266 3291 3267 3295
rect 3271 3291 3272 3295
rect 3798 3292 3799 3296
rect 3803 3292 3804 3296
rect 3984 3294 3986 3296
rect 5418 3295 5419 3299
rect 5423 3298 5424 3299
rect 5423 3296 5554 3298
rect 5423 3295 5424 3296
rect 5418 3294 5424 3295
rect 5552 3294 5554 3296
rect 3983 3293 3989 3294
rect 5551 3293 5557 3294
rect 3886 3292 3892 3293
rect 3798 3291 3804 3292
rect 3838 3291 3844 3292
rect 3266 3290 3272 3291
rect 2679 3287 2685 3288
rect 2679 3283 2680 3287
rect 2684 3286 2685 3287
rect 3838 3287 3839 3291
rect 3843 3287 3844 3291
rect 3886 3288 3887 3292
rect 3891 3288 3892 3292
rect 3983 3289 3984 3293
rect 3988 3289 3989 3293
rect 3983 3288 3989 3289
rect 4166 3292 4172 3293
rect 4454 3292 4460 3293
rect 4718 3292 4724 3293
rect 4966 3292 4972 3293
rect 5206 3292 5212 3293
rect 5454 3292 5460 3293
rect 4166 3288 4167 3292
rect 4171 3288 4172 3292
rect 3886 3287 3892 3288
rect 4166 3287 4172 3288
rect 4262 3291 4269 3292
rect 4262 3287 4263 3291
rect 4268 3287 4269 3291
rect 4454 3288 4455 3292
rect 4459 3288 4460 3292
rect 4454 3287 4460 3288
rect 4551 3291 4557 3292
rect 4551 3287 4552 3291
rect 4556 3290 4557 3291
rect 4698 3291 4704 3292
rect 4698 3290 4699 3291
rect 4556 3288 4699 3290
rect 4556 3287 4557 3288
rect 3838 3286 3844 3287
rect 4262 3286 4269 3287
rect 4551 3286 4557 3287
rect 4698 3287 4699 3288
rect 4703 3287 4704 3291
rect 4718 3288 4719 3292
rect 4723 3288 4724 3292
rect 4718 3287 4724 3288
rect 4815 3291 4824 3292
rect 4815 3287 4816 3291
rect 4823 3287 4824 3291
rect 4966 3288 4967 3292
rect 4971 3288 4972 3292
rect 4966 3287 4972 3288
rect 5058 3291 5069 3292
rect 5058 3287 5059 3291
rect 5063 3287 5064 3291
rect 5068 3287 5069 3291
rect 5206 3288 5207 3292
rect 5211 3288 5212 3292
rect 5206 3287 5212 3288
rect 5302 3291 5309 3292
rect 5302 3287 5303 3291
rect 5308 3287 5309 3291
rect 5454 3288 5455 3292
rect 5459 3288 5460 3292
rect 5551 3289 5552 3293
rect 5556 3289 5557 3293
rect 5551 3288 5557 3289
rect 5662 3291 5668 3292
rect 5454 3287 5460 3288
rect 5662 3287 5663 3291
rect 5667 3287 5668 3291
rect 4698 3286 4704 3287
rect 4815 3286 4824 3287
rect 5058 3286 5069 3287
rect 5302 3286 5309 3287
rect 5662 3286 5668 3287
rect 2684 3284 2842 3286
rect 2684 3283 2685 3284
rect 2679 3282 2685 3283
rect 2840 3282 2842 3284
rect 2839 3281 2845 3282
rect 110 3280 116 3281
rect 1934 3280 1940 3281
rect 2558 3280 2564 3281
rect 2742 3280 2748 3281
rect 110 3276 111 3280
rect 115 3276 116 3280
rect 110 3275 116 3276
rect 754 3279 760 3280
rect 754 3275 755 3279
rect 759 3275 760 3279
rect 754 3274 760 3275
rect 890 3279 896 3280
rect 890 3275 891 3279
rect 895 3275 896 3279
rect 890 3274 896 3275
rect 1034 3279 1040 3280
rect 1034 3275 1035 3279
rect 1039 3275 1040 3279
rect 1034 3274 1040 3275
rect 1186 3279 1192 3280
rect 1186 3275 1187 3279
rect 1191 3275 1192 3279
rect 1186 3274 1192 3275
rect 1338 3279 1344 3280
rect 1338 3275 1339 3279
rect 1343 3275 1344 3279
rect 1338 3274 1344 3275
rect 1490 3279 1496 3280
rect 1490 3275 1491 3279
rect 1495 3275 1496 3279
rect 1490 3274 1496 3275
rect 1650 3279 1656 3280
rect 1650 3275 1651 3279
rect 1655 3275 1656 3279
rect 1650 3274 1656 3275
rect 1786 3279 1792 3280
rect 1786 3275 1787 3279
rect 1791 3275 1792 3279
rect 1934 3276 1935 3280
rect 1939 3276 1940 3280
rect 1934 3275 1940 3276
rect 1974 3279 1980 3280
rect 1974 3275 1975 3279
rect 1979 3275 1980 3279
rect 2558 3276 2559 3280
rect 2563 3276 2564 3280
rect 2558 3275 2564 3276
rect 2654 3279 2661 3280
rect 2654 3275 2655 3279
rect 2660 3275 2661 3279
rect 2742 3276 2743 3280
rect 2747 3276 2748 3280
rect 2839 3277 2840 3281
rect 2844 3277 2845 3281
rect 2839 3276 2845 3277
rect 2926 3280 2932 3281
rect 3110 3280 3116 3281
rect 3294 3280 3300 3281
rect 2926 3276 2927 3280
rect 2931 3276 2932 3280
rect 2742 3275 2748 3276
rect 2926 3275 2932 3276
rect 3023 3279 3029 3280
rect 3023 3275 3024 3279
rect 3028 3278 3029 3279
rect 3090 3279 3096 3280
rect 3090 3278 3091 3279
rect 3028 3276 3091 3278
rect 3028 3275 3029 3276
rect 1786 3274 1792 3275
rect 1974 3274 1980 3275
rect 2654 3274 2661 3275
rect 3023 3274 3029 3275
rect 3090 3275 3091 3276
rect 3095 3275 3096 3279
rect 3110 3276 3111 3280
rect 3115 3276 3116 3280
rect 3110 3275 3116 3276
rect 3207 3279 3213 3280
rect 3207 3275 3208 3279
rect 3212 3278 3213 3279
rect 3274 3279 3280 3280
rect 3274 3278 3275 3279
rect 3212 3276 3275 3278
rect 3212 3275 3213 3276
rect 3090 3274 3096 3275
rect 3207 3274 3213 3275
rect 3274 3275 3275 3276
rect 3279 3275 3280 3279
rect 3294 3276 3295 3280
rect 3299 3276 3300 3280
rect 3294 3275 3300 3276
rect 3391 3279 3397 3280
rect 3391 3275 3392 3279
rect 3396 3278 3397 3279
rect 3402 3279 3408 3280
rect 3402 3278 3403 3279
rect 3396 3276 3403 3278
rect 3396 3275 3397 3276
rect 3274 3274 3280 3275
rect 3391 3274 3397 3275
rect 3402 3275 3403 3276
rect 3407 3275 3408 3279
rect 3402 3274 3408 3275
rect 3798 3279 3804 3280
rect 3798 3275 3799 3279
rect 3803 3275 3804 3279
rect 3798 3274 3804 3275
rect 1018 3271 1024 3272
rect 1018 3267 1019 3271
rect 1023 3270 1024 3271
rect 1023 3268 1314 3270
rect 1023 3267 1024 3268
rect 1018 3266 1024 3267
rect 1312 3266 1314 3268
rect 1311 3265 1317 3266
rect 782 3264 788 3265
rect 918 3264 924 3265
rect 1062 3264 1068 3265
rect 1214 3264 1220 3265
rect 110 3263 116 3264
rect 110 3259 111 3263
rect 115 3259 116 3263
rect 782 3260 783 3264
rect 787 3260 788 3264
rect 782 3259 788 3260
rect 874 3263 885 3264
rect 874 3259 875 3263
rect 879 3259 880 3263
rect 884 3259 885 3263
rect 918 3260 919 3264
rect 923 3260 924 3264
rect 918 3259 924 3260
rect 1010 3263 1021 3264
rect 1010 3259 1011 3263
rect 1015 3259 1016 3263
rect 1020 3259 1021 3263
rect 1062 3260 1063 3264
rect 1067 3260 1068 3264
rect 1062 3259 1068 3260
rect 1158 3263 1165 3264
rect 1158 3259 1159 3263
rect 1164 3259 1165 3263
rect 1214 3260 1215 3264
rect 1219 3260 1220 3264
rect 1311 3261 1312 3265
rect 1316 3261 1317 3265
rect 1311 3260 1317 3261
rect 1366 3264 1372 3265
rect 1518 3264 1524 3265
rect 1678 3264 1684 3265
rect 1814 3264 1820 3265
rect 1366 3260 1367 3264
rect 1371 3260 1372 3264
rect 1214 3259 1220 3260
rect 1366 3259 1372 3260
rect 1462 3263 1469 3264
rect 1462 3259 1463 3263
rect 1468 3259 1469 3263
rect 1518 3260 1519 3264
rect 1523 3260 1524 3264
rect 1518 3259 1524 3260
rect 1615 3263 1621 3264
rect 1615 3259 1616 3263
rect 1620 3262 1621 3263
rect 1658 3263 1664 3264
rect 1658 3262 1659 3263
rect 1620 3260 1659 3262
rect 1620 3259 1621 3260
rect 110 3258 116 3259
rect 874 3258 885 3259
rect 1010 3258 1021 3259
rect 1158 3258 1165 3259
rect 1462 3258 1469 3259
rect 1615 3258 1621 3259
rect 1658 3259 1659 3260
rect 1663 3259 1664 3263
rect 1678 3260 1679 3264
rect 1683 3260 1684 3264
rect 1678 3259 1684 3260
rect 1775 3263 1781 3264
rect 1775 3259 1776 3263
rect 1780 3262 1781 3263
rect 1794 3263 1800 3264
rect 1794 3262 1795 3263
rect 1780 3260 1795 3262
rect 1780 3259 1781 3260
rect 1658 3258 1664 3259
rect 1775 3258 1781 3259
rect 1794 3259 1795 3260
rect 1799 3259 1800 3263
rect 1814 3260 1815 3264
rect 1819 3260 1820 3264
rect 1814 3259 1820 3260
rect 1910 3263 1917 3264
rect 1910 3259 1911 3263
rect 1916 3259 1917 3263
rect 1794 3258 1800 3259
rect 1910 3258 1917 3259
rect 1934 3263 1940 3264
rect 1934 3259 1935 3263
rect 1939 3259 1940 3263
rect 1934 3258 1940 3259
rect 1974 3221 1980 3222
rect 3798 3221 3804 3222
rect 1130 3219 1136 3220
rect 1130 3215 1131 3219
rect 1135 3218 1136 3219
rect 1434 3219 1440 3220
rect 1135 3216 1322 3218
rect 1135 3215 1136 3216
rect 1130 3214 1136 3215
rect 110 3205 116 3206
rect 110 3201 111 3205
rect 115 3201 116 3205
rect 110 3200 116 3201
rect 390 3204 396 3205
rect 646 3204 652 3205
rect 926 3204 932 3205
rect 1222 3204 1228 3205
rect 1320 3204 1322 3216
rect 1434 3215 1435 3219
rect 1439 3218 1440 3219
rect 1439 3216 1626 3218
rect 1974 3217 1975 3221
rect 1979 3217 1980 3221
rect 1974 3216 1980 3217
rect 2022 3220 2028 3221
rect 2254 3220 2260 3221
rect 2502 3220 2508 3221
rect 2742 3220 2748 3221
rect 2974 3220 2980 3221
rect 3206 3220 3212 3221
rect 3446 3220 3452 3221
rect 2022 3216 2023 3220
rect 2027 3216 2028 3220
rect 1439 3215 1440 3216
rect 1434 3214 1440 3215
rect 1526 3204 1532 3205
rect 1624 3204 1626 3216
rect 2022 3215 2028 3216
rect 2119 3219 2125 3220
rect 2119 3215 2120 3219
rect 2124 3218 2125 3219
rect 2142 3219 2148 3220
rect 2142 3218 2143 3219
rect 2124 3216 2143 3218
rect 2124 3215 2125 3216
rect 2119 3214 2125 3215
rect 2142 3215 2143 3216
rect 2147 3215 2148 3219
rect 2254 3216 2255 3220
rect 2259 3216 2260 3220
rect 2254 3215 2260 3216
rect 2346 3219 2357 3220
rect 2346 3215 2347 3219
rect 2351 3215 2352 3219
rect 2356 3215 2357 3219
rect 2502 3216 2503 3220
rect 2507 3216 2508 3220
rect 2502 3215 2508 3216
rect 2594 3219 2605 3220
rect 2594 3215 2595 3219
rect 2599 3215 2600 3219
rect 2604 3215 2605 3219
rect 2742 3216 2743 3220
rect 2747 3216 2748 3220
rect 2742 3215 2748 3216
rect 2839 3219 2845 3220
rect 2839 3215 2840 3219
rect 2844 3218 2845 3219
rect 2854 3219 2860 3220
rect 2854 3218 2855 3219
rect 2844 3216 2855 3218
rect 2844 3215 2845 3216
rect 2142 3214 2148 3215
rect 2346 3214 2357 3215
rect 2594 3214 2605 3215
rect 2839 3214 2845 3215
rect 2854 3215 2855 3216
rect 2859 3215 2860 3219
rect 2974 3216 2975 3220
rect 2979 3216 2980 3220
rect 2974 3215 2980 3216
rect 3070 3219 3077 3220
rect 3070 3215 3071 3219
rect 3076 3215 3077 3219
rect 3206 3216 3207 3220
rect 3211 3216 3212 3220
rect 3206 3215 3212 3216
rect 3298 3219 3309 3220
rect 3298 3215 3299 3219
rect 3303 3215 3304 3219
rect 3308 3215 3309 3219
rect 3446 3216 3447 3220
rect 3451 3216 3452 3220
rect 3446 3215 3452 3216
rect 3542 3219 3549 3220
rect 3542 3215 3543 3219
rect 3548 3215 3549 3219
rect 3798 3217 3799 3221
rect 3803 3217 3804 3221
rect 3798 3216 3804 3217
rect 2854 3214 2860 3215
rect 3070 3214 3077 3215
rect 3298 3214 3309 3215
rect 3542 3214 3549 3215
rect 3838 3209 3844 3210
rect 5662 3209 5668 3210
rect 1934 3205 1940 3206
rect 1994 3205 2000 3206
rect 1814 3204 1820 3205
rect 390 3200 391 3204
rect 395 3200 396 3204
rect 390 3199 396 3200
rect 487 3203 496 3204
rect 487 3199 488 3203
rect 495 3199 496 3203
rect 646 3200 647 3204
rect 651 3200 652 3204
rect 646 3199 652 3200
rect 742 3203 749 3204
rect 742 3199 743 3203
rect 748 3199 749 3203
rect 926 3200 927 3204
rect 931 3200 932 3204
rect 926 3199 932 3200
rect 1018 3203 1029 3204
rect 1018 3199 1019 3203
rect 1023 3199 1024 3203
rect 1028 3199 1029 3203
rect 1222 3200 1223 3204
rect 1227 3200 1228 3204
rect 1222 3199 1228 3200
rect 1319 3203 1325 3204
rect 1319 3199 1320 3203
rect 1324 3199 1325 3203
rect 1526 3200 1527 3204
rect 1531 3200 1532 3204
rect 1526 3199 1532 3200
rect 1623 3203 1629 3204
rect 1623 3199 1624 3203
rect 1628 3199 1629 3203
rect 1814 3200 1815 3204
rect 1819 3200 1820 3204
rect 1814 3199 1820 3200
rect 1911 3203 1917 3204
rect 1911 3199 1912 3203
rect 1916 3202 1917 3203
rect 1926 3203 1932 3204
rect 1926 3202 1927 3203
rect 1916 3200 1927 3202
rect 1916 3199 1917 3200
rect 487 3198 496 3199
rect 742 3198 749 3199
rect 1018 3198 1029 3199
rect 1319 3198 1325 3199
rect 1623 3198 1629 3199
rect 1911 3198 1917 3199
rect 1926 3199 1927 3200
rect 1931 3199 1932 3203
rect 1934 3201 1935 3205
rect 1939 3201 1940 3205
rect 1934 3200 1940 3201
rect 1974 3204 1980 3205
rect 1974 3200 1975 3204
rect 1979 3200 1980 3204
rect 1994 3201 1995 3205
rect 1999 3201 2000 3205
rect 1994 3200 2000 3201
rect 2226 3205 2232 3206
rect 2226 3201 2227 3205
rect 2231 3201 2232 3205
rect 2226 3200 2232 3201
rect 2474 3205 2480 3206
rect 2474 3201 2475 3205
rect 2479 3201 2480 3205
rect 2474 3200 2480 3201
rect 2714 3205 2720 3206
rect 2714 3201 2715 3205
rect 2719 3201 2720 3205
rect 2714 3200 2720 3201
rect 2946 3205 2952 3206
rect 2946 3201 2947 3205
rect 2951 3201 2952 3205
rect 2946 3200 2952 3201
rect 3178 3205 3184 3206
rect 3178 3201 3179 3205
rect 3183 3201 3184 3205
rect 3178 3200 3184 3201
rect 3418 3205 3424 3206
rect 3838 3205 3839 3209
rect 3843 3205 3844 3209
rect 3418 3201 3419 3205
rect 3423 3201 3424 3205
rect 3418 3200 3424 3201
rect 3798 3204 3804 3205
rect 3838 3204 3844 3205
rect 3910 3208 3916 3209
rect 4182 3208 4188 3209
rect 4438 3208 4444 3209
rect 4686 3208 4692 3209
rect 4934 3208 4940 3209
rect 5190 3208 5196 3209
rect 3910 3204 3911 3208
rect 3915 3204 3916 3208
rect 3798 3200 3799 3204
rect 3803 3200 3804 3204
rect 3910 3203 3916 3204
rect 4007 3207 4013 3208
rect 4007 3203 4008 3207
rect 4012 3206 4013 3207
rect 4146 3207 4152 3208
rect 4146 3206 4147 3207
rect 4012 3204 4147 3206
rect 4012 3203 4013 3204
rect 4007 3202 4013 3203
rect 4146 3203 4147 3204
rect 4151 3203 4152 3207
rect 4182 3204 4183 3208
rect 4187 3204 4188 3208
rect 4182 3203 4188 3204
rect 4279 3207 4285 3208
rect 4279 3203 4280 3207
rect 4284 3206 4285 3207
rect 4319 3207 4325 3208
rect 4319 3206 4320 3207
rect 4284 3204 4320 3206
rect 4284 3203 4285 3204
rect 4146 3202 4152 3203
rect 4279 3202 4285 3203
rect 4319 3203 4320 3204
rect 4324 3203 4325 3207
rect 4438 3204 4439 3208
rect 4443 3204 4444 3208
rect 4438 3203 4444 3204
rect 4534 3207 4541 3208
rect 4534 3203 4535 3207
rect 4540 3203 4541 3207
rect 4686 3204 4687 3208
rect 4691 3204 4692 3208
rect 4686 3203 4692 3204
rect 4778 3207 4789 3208
rect 4778 3203 4779 3207
rect 4783 3203 4784 3207
rect 4788 3203 4789 3207
rect 4934 3204 4935 3208
rect 4939 3204 4940 3208
rect 4934 3203 4940 3204
rect 5030 3207 5037 3208
rect 5030 3203 5031 3207
rect 5036 3203 5037 3207
rect 5190 3204 5191 3208
rect 5195 3204 5196 3208
rect 5190 3203 5196 3204
rect 5286 3207 5293 3208
rect 5286 3203 5287 3207
rect 5292 3203 5293 3207
rect 5662 3205 5663 3209
rect 5667 3205 5668 3209
rect 5662 3204 5668 3205
rect 4319 3202 4325 3203
rect 4534 3202 4541 3203
rect 4778 3202 4789 3203
rect 5030 3202 5037 3203
rect 5286 3202 5293 3203
rect 1974 3199 1980 3200
rect 3798 3199 3804 3200
rect 1926 3198 1932 3199
rect 3882 3193 3888 3194
rect 3838 3192 3844 3193
rect 362 3189 368 3190
rect 110 3188 116 3189
rect 110 3184 111 3188
rect 115 3184 116 3188
rect 362 3185 363 3189
rect 367 3185 368 3189
rect 362 3184 368 3185
rect 618 3189 624 3190
rect 618 3185 619 3189
rect 623 3185 624 3189
rect 618 3184 624 3185
rect 898 3189 904 3190
rect 898 3185 899 3189
rect 903 3185 904 3189
rect 898 3184 904 3185
rect 1194 3189 1200 3190
rect 1194 3185 1195 3189
rect 1199 3185 1200 3189
rect 1194 3184 1200 3185
rect 1498 3189 1504 3190
rect 1498 3185 1499 3189
rect 1503 3185 1504 3189
rect 1498 3184 1504 3185
rect 1786 3189 1792 3190
rect 1786 3185 1787 3189
rect 1791 3185 1792 3189
rect 1786 3184 1792 3185
rect 1934 3188 1940 3189
rect 1934 3184 1935 3188
rect 1939 3184 1940 3188
rect 3838 3188 3839 3192
rect 3843 3188 3844 3192
rect 3882 3189 3883 3193
rect 3887 3189 3888 3193
rect 3882 3188 3888 3189
rect 4154 3193 4160 3194
rect 4154 3189 4155 3193
rect 4159 3189 4160 3193
rect 4154 3188 4160 3189
rect 4410 3193 4416 3194
rect 4410 3189 4411 3193
rect 4415 3189 4416 3193
rect 4410 3188 4416 3189
rect 4658 3193 4664 3194
rect 4658 3189 4659 3193
rect 4663 3189 4664 3193
rect 4658 3188 4664 3189
rect 4906 3193 4912 3194
rect 4906 3189 4907 3193
rect 4911 3189 4912 3193
rect 4906 3188 4912 3189
rect 5162 3193 5168 3194
rect 5162 3189 5163 3193
rect 5167 3189 5168 3193
rect 5162 3188 5168 3189
rect 5662 3192 5668 3193
rect 5662 3188 5663 3192
rect 5667 3188 5668 3192
rect 3838 3187 3844 3188
rect 5662 3187 5668 3188
rect 110 3183 116 3184
rect 1934 3183 1940 3184
rect 1926 3155 1932 3156
rect 1926 3151 1927 3155
rect 1931 3154 1932 3155
rect 2142 3155 2148 3156
rect 1931 3152 2001 3154
rect 1931 3151 1932 3152
rect 1926 3150 1932 3151
rect 2142 3151 2143 3155
rect 2147 3154 2148 3155
rect 2654 3155 2660 3156
rect 2654 3154 2655 3155
rect 2147 3152 2233 3154
rect 2573 3152 2655 3154
rect 2147 3151 2148 3152
rect 2142 3150 2148 3151
rect 2654 3151 2655 3152
rect 2659 3151 2660 3155
rect 2854 3155 2860 3156
rect 2654 3150 2660 3151
rect 2812 3146 2814 3153
rect 2854 3151 2855 3155
rect 2859 3154 2860 3155
rect 3402 3155 3408 3156
rect 2859 3152 2953 3154
rect 2859 3151 2860 3152
rect 2854 3150 2860 3151
rect 2898 3147 2904 3148
rect 2898 3146 2899 3147
rect 2812 3144 2899 3146
rect 2898 3143 2899 3144
rect 2903 3143 2904 3147
rect 3276 3146 3278 3153
rect 3402 3151 3403 3155
rect 3407 3154 3408 3155
rect 3407 3152 3425 3154
rect 3407 3151 3408 3152
rect 3402 3150 3408 3151
rect 3542 3147 3548 3148
rect 3542 3146 3543 3147
rect 3276 3144 3543 3146
rect 2898 3142 2904 3143
rect 3542 3143 3543 3144
rect 3547 3143 3548 3147
rect 3542 3142 3548 3143
rect 4050 3143 4056 3144
rect 4050 3142 4051 3143
rect 3981 3140 4051 3142
rect 1010 3139 1016 3140
rect 1010 3138 1011 3139
rect 460 3130 462 3137
rect 717 3136 902 3138
rect 997 3136 1011 3138
rect 742 3131 748 3132
rect 742 3130 743 3131
rect 460 3128 743 3130
rect 742 3127 743 3128
rect 747 3127 748 3131
rect 900 3130 902 3136
rect 1010 3135 1011 3136
rect 1015 3135 1016 3139
rect 1010 3134 1016 3135
rect 1026 3139 1032 3140
rect 1026 3135 1027 3139
rect 1031 3138 1032 3139
rect 1574 3139 1580 3140
rect 1031 3136 1201 3138
rect 1031 3135 1032 3136
rect 1026 3134 1032 3135
rect 1574 3135 1575 3139
rect 1579 3135 1580 3139
rect 1910 3139 1916 3140
rect 1910 3138 1911 3139
rect 1885 3136 1911 3138
rect 1574 3134 1580 3135
rect 1910 3135 1911 3136
rect 1915 3135 1916 3139
rect 4050 3139 4051 3140
rect 4055 3139 4056 3143
rect 4319 3143 4325 3144
rect 4050 3138 4056 3139
rect 1910 3134 1916 3135
rect 4252 3134 4254 3141
rect 4319 3139 4320 3143
rect 4324 3142 4325 3143
rect 4818 3143 4824 3144
rect 4324 3140 4417 3142
rect 4757 3140 4814 3142
rect 4324 3139 4325 3140
rect 4319 3138 4325 3139
rect 4778 3135 4784 3136
rect 4778 3134 4779 3135
rect 4252 3132 4779 3134
rect 1018 3131 1024 3132
rect 1018 3130 1019 3131
rect 900 3128 1019 3130
rect 742 3126 748 3127
rect 1018 3127 1019 3128
rect 1023 3127 1024 3131
rect 4778 3131 4779 3132
rect 4783 3131 4784 3135
rect 4812 3134 4814 3140
rect 4818 3139 4819 3143
rect 4823 3142 4824 3143
rect 5030 3143 5036 3144
rect 4823 3140 4913 3142
rect 4823 3139 4824 3140
rect 4818 3138 4824 3139
rect 5030 3139 5031 3143
rect 5035 3142 5036 3143
rect 5035 3140 5169 3142
rect 5035 3139 5036 3140
rect 5030 3138 5036 3139
rect 5286 3135 5292 3136
rect 5286 3134 5287 3135
rect 4812 3132 5287 3134
rect 4778 3130 4784 3131
rect 5286 3131 5287 3132
rect 5291 3131 5292 3135
rect 5286 3130 5292 3131
rect 1018 3126 1024 3127
rect 2594 3123 2600 3124
rect 2594 3122 2595 3123
rect 2581 3120 2595 3122
rect 2594 3119 2595 3120
rect 2599 3119 2600 3123
rect 3298 3123 3304 3124
rect 3298 3122 3299 3123
rect 3173 3120 3299 3122
rect 2594 3118 2600 3119
rect 2874 3119 2880 3120
rect 2874 3115 2875 3119
rect 2879 3115 2880 3119
rect 3298 3119 3299 3120
rect 3303 3119 3304 3123
rect 3298 3118 3304 3119
rect 3378 3119 3384 3120
rect 2874 3114 2880 3115
rect 3378 3115 3379 3119
rect 3383 3115 3384 3119
rect 3378 3114 3384 3115
rect 3658 3119 3664 3120
rect 3658 3115 3659 3119
rect 3663 3115 3664 3119
rect 3658 3114 3664 3115
rect 4094 3107 4100 3108
rect 4094 3106 4095 3107
rect 4029 3104 4095 3106
rect 4094 3103 4095 3104
rect 4099 3103 4100 3107
rect 4534 3107 4540 3108
rect 4094 3102 4100 3103
rect 4226 3103 4232 3104
rect 430 3099 436 3100
rect 430 3098 431 3099
rect 259 3096 431 3098
rect 259 3094 261 3096
rect 430 3095 431 3096
rect 435 3095 436 3099
rect 4226 3099 4227 3103
rect 4231 3099 4232 3103
rect 4226 3098 4232 3099
rect 4338 3103 4344 3104
rect 4338 3099 4339 3103
rect 4343 3099 4344 3103
rect 4534 3103 4535 3107
rect 4539 3103 4540 3107
rect 4534 3102 4540 3103
rect 4722 3103 4728 3104
rect 4338 3098 4344 3099
rect 4722 3099 4723 3103
rect 4727 3099 4728 3103
rect 4722 3098 4728 3099
rect 4922 3103 4928 3104
rect 4922 3099 4923 3103
rect 4927 3099 4928 3103
rect 4922 3098 4928 3099
rect 430 3094 436 3095
rect 490 3095 496 3096
rect 229 3092 261 3094
rect 490 3091 491 3095
rect 495 3094 496 3095
rect 1266 3095 1272 3096
rect 1266 3094 1267 3095
rect 495 3092 513 3094
rect 1189 3092 1267 3094
rect 495 3091 496 3092
rect 490 3090 496 3091
rect 802 3091 808 3092
rect 400 3086 402 3089
rect 498 3087 504 3088
rect 498 3086 499 3087
rect 400 3084 499 3086
rect 498 3083 499 3084
rect 503 3083 504 3087
rect 802 3087 803 3091
rect 807 3087 808 3091
rect 802 3086 808 3087
rect 906 3091 912 3092
rect 906 3087 907 3091
rect 911 3087 912 3091
rect 1266 3091 1267 3092
rect 1271 3091 1272 3095
rect 1775 3095 1781 3096
rect 1775 3094 1776 3095
rect 1725 3092 1776 3094
rect 1266 3090 1272 3091
rect 1282 3091 1288 3092
rect 906 3086 912 3087
rect 1282 3087 1283 3091
rect 1287 3087 1288 3091
rect 1282 3086 1288 3087
rect 1458 3091 1464 3092
rect 1458 3087 1459 3091
rect 1463 3087 1464 3091
rect 1775 3091 1776 3092
rect 1780 3091 1781 3095
rect 2346 3095 2352 3096
rect 2346 3094 2347 3095
rect 1885 3092 2347 3094
rect 1775 3090 1781 3091
rect 2346 3091 2347 3092
rect 2351 3091 2352 3095
rect 2346 3090 2352 3091
rect 1458 3086 1464 3087
rect 498 3082 504 3083
rect 2874 3079 2880 3080
rect 2874 3075 2875 3079
rect 2879 3078 2880 3079
rect 3214 3079 3220 3080
rect 3214 3078 3215 3079
rect 2879 3076 3215 3078
rect 2879 3075 2880 3076
rect 2874 3074 2880 3075
rect 3214 3075 3215 3076
rect 3219 3075 3220 3079
rect 3214 3074 3220 3075
rect 1974 3072 1980 3073
rect 3798 3072 3804 3073
rect 1974 3068 1975 3072
rect 1979 3068 1980 3072
rect 1974 3067 1980 3068
rect 2482 3071 2488 3072
rect 2482 3067 2483 3071
rect 2487 3067 2488 3071
rect 2482 3066 2488 3067
rect 2778 3071 2784 3072
rect 2778 3067 2779 3071
rect 2783 3067 2784 3071
rect 2778 3066 2784 3067
rect 3074 3071 3080 3072
rect 3074 3067 3075 3071
rect 3079 3067 3080 3071
rect 3074 3066 3080 3067
rect 3370 3071 3376 3072
rect 3370 3067 3371 3071
rect 3375 3067 3376 3071
rect 3370 3066 3376 3067
rect 3650 3071 3656 3072
rect 3650 3067 3651 3071
rect 3655 3067 3656 3071
rect 3798 3068 3799 3072
rect 3803 3068 3804 3072
rect 3798 3067 3804 3068
rect 3650 3066 3656 3067
rect 2510 3056 2516 3057
rect 2806 3056 2812 3057
rect 3102 3056 3108 3057
rect 3398 3056 3404 3057
rect 3678 3056 3684 3057
rect 3838 3056 3844 3057
rect 5662 3056 5668 3057
rect 1974 3055 1980 3056
rect 1974 3051 1975 3055
rect 1979 3051 1980 3055
rect 2510 3052 2511 3056
rect 2515 3052 2516 3056
rect 2510 3051 2516 3052
rect 2606 3055 2613 3056
rect 2606 3051 2607 3055
rect 2612 3051 2613 3055
rect 2806 3052 2807 3056
rect 2811 3052 2812 3056
rect 2806 3051 2812 3052
rect 2898 3055 2909 3056
rect 2898 3051 2899 3055
rect 2903 3051 2904 3055
rect 2908 3051 2909 3055
rect 3102 3052 3103 3056
rect 3107 3052 3108 3056
rect 3102 3051 3108 3052
rect 3199 3055 3205 3056
rect 3199 3051 3200 3055
rect 3204 3054 3205 3055
rect 3378 3055 3384 3056
rect 3378 3054 3379 3055
rect 3204 3052 3379 3054
rect 3204 3051 3205 3052
rect 1974 3050 1980 3051
rect 2606 3050 2613 3051
rect 2898 3050 2909 3051
rect 3199 3050 3205 3051
rect 3378 3051 3379 3052
rect 3383 3051 3384 3055
rect 3398 3052 3399 3056
rect 3403 3052 3404 3056
rect 3398 3051 3404 3052
rect 3495 3055 3501 3056
rect 3495 3051 3496 3055
rect 3500 3054 3501 3055
rect 3658 3055 3664 3056
rect 3658 3054 3659 3055
rect 3500 3052 3659 3054
rect 3500 3051 3501 3052
rect 3378 3050 3384 3051
rect 3495 3050 3501 3051
rect 3658 3051 3659 3052
rect 3663 3051 3664 3055
rect 3678 3052 3679 3056
rect 3683 3052 3684 3056
rect 3678 3051 3684 3052
rect 3770 3055 3781 3056
rect 3770 3051 3771 3055
rect 3775 3051 3776 3055
rect 3780 3051 3781 3055
rect 3658 3050 3664 3051
rect 3770 3050 3781 3051
rect 3798 3055 3804 3056
rect 3798 3051 3799 3055
rect 3803 3051 3804 3055
rect 3838 3052 3839 3056
rect 3843 3052 3844 3056
rect 3838 3051 3844 3052
rect 3930 3055 3936 3056
rect 3930 3051 3931 3055
rect 3935 3051 3936 3055
rect 3798 3050 3804 3051
rect 3930 3050 3936 3051
rect 4130 3055 4136 3056
rect 4130 3051 4131 3055
rect 4135 3051 4136 3055
rect 4130 3050 4136 3051
rect 4330 3055 4336 3056
rect 4330 3051 4331 3055
rect 4335 3051 4336 3055
rect 4330 3050 4336 3051
rect 4522 3055 4528 3056
rect 4522 3051 4523 3055
rect 4527 3051 4528 3055
rect 4522 3050 4528 3051
rect 4714 3055 4720 3056
rect 4714 3051 4715 3055
rect 4719 3051 4720 3055
rect 4714 3050 4720 3051
rect 4914 3055 4920 3056
rect 4914 3051 4915 3055
rect 4919 3051 4920 3055
rect 5662 3052 5663 3056
rect 5667 3052 5668 3056
rect 5662 3051 5668 3052
rect 4914 3050 4920 3051
rect 110 3044 116 3045
rect 1934 3044 1940 3045
rect 110 3040 111 3044
rect 115 3040 116 3044
rect 110 3039 116 3040
rect 130 3043 136 3044
rect 130 3039 131 3043
rect 135 3039 136 3043
rect 130 3038 136 3039
rect 306 3043 312 3044
rect 306 3039 307 3043
rect 311 3039 312 3043
rect 306 3038 312 3039
rect 506 3043 512 3044
rect 506 3039 507 3043
rect 511 3039 512 3043
rect 506 3038 512 3039
rect 706 3043 712 3044
rect 706 3039 707 3043
rect 711 3039 712 3043
rect 706 3038 712 3039
rect 898 3043 904 3044
rect 898 3039 899 3043
rect 903 3039 904 3043
rect 898 3038 904 3039
rect 1090 3043 1096 3044
rect 1090 3039 1091 3043
rect 1095 3039 1096 3043
rect 1090 3038 1096 3039
rect 1274 3043 1280 3044
rect 1274 3039 1275 3043
rect 1279 3039 1280 3043
rect 1274 3038 1280 3039
rect 1450 3043 1456 3044
rect 1450 3039 1451 3043
rect 1455 3039 1456 3043
rect 1450 3038 1456 3039
rect 1626 3043 1632 3044
rect 1626 3039 1627 3043
rect 1631 3039 1632 3043
rect 1626 3038 1632 3039
rect 1786 3043 1792 3044
rect 1786 3039 1787 3043
rect 1791 3039 1792 3043
rect 1934 3040 1935 3044
rect 1939 3040 1940 3044
rect 3958 3040 3964 3041
rect 4158 3040 4164 3041
rect 4358 3040 4364 3041
rect 4550 3040 4556 3041
rect 4742 3040 4748 3041
rect 4942 3040 4948 3041
rect 1934 3039 1940 3040
rect 3838 3039 3844 3040
rect 1786 3038 1792 3039
rect 498 3035 504 3036
rect 498 3031 499 3035
rect 503 3034 504 3035
rect 1266 3035 1272 3036
rect 503 3032 634 3034
rect 503 3031 504 3032
rect 498 3030 504 3031
rect 158 3028 164 3029
rect 334 3028 340 3029
rect 534 3028 540 3029
rect 632 3028 634 3032
rect 1266 3031 1267 3035
rect 1271 3034 1272 3035
rect 1775 3035 1781 3036
rect 1271 3032 1754 3034
rect 1271 3031 1272 3032
rect 1266 3030 1272 3031
rect 734 3028 740 3029
rect 926 3028 932 3029
rect 1118 3028 1124 3029
rect 1302 3028 1308 3029
rect 1478 3028 1484 3029
rect 1654 3028 1660 3029
rect 1752 3028 1754 3032
rect 1775 3031 1776 3035
rect 1780 3034 1781 3035
rect 3838 3035 3839 3039
rect 3843 3035 3844 3039
rect 3958 3036 3959 3040
rect 3963 3036 3964 3040
rect 3958 3035 3964 3036
rect 4050 3039 4061 3040
rect 4050 3035 4051 3039
rect 4055 3035 4056 3039
rect 4060 3035 4061 3039
rect 4158 3036 4159 3040
rect 4163 3036 4164 3040
rect 4158 3035 4164 3036
rect 4255 3039 4261 3040
rect 4255 3035 4256 3039
rect 4260 3038 4261 3039
rect 4338 3039 4344 3040
rect 4338 3038 4339 3039
rect 4260 3036 4339 3038
rect 4260 3035 4261 3036
rect 3838 3034 3844 3035
rect 4050 3034 4061 3035
rect 4255 3034 4261 3035
rect 4338 3035 4339 3036
rect 4343 3035 4344 3039
rect 4358 3036 4359 3040
rect 4363 3036 4364 3040
rect 4358 3035 4364 3036
rect 4455 3039 4461 3040
rect 4455 3035 4456 3039
rect 4460 3038 4461 3039
rect 4466 3039 4472 3040
rect 4466 3038 4467 3039
rect 4460 3036 4467 3038
rect 4460 3035 4461 3036
rect 4338 3034 4344 3035
rect 4455 3034 4461 3035
rect 4466 3035 4467 3036
rect 4471 3035 4472 3039
rect 4550 3036 4551 3040
rect 4555 3036 4556 3040
rect 4550 3035 4556 3036
rect 4647 3039 4653 3040
rect 4647 3035 4648 3039
rect 4652 3038 4653 3039
rect 4722 3039 4728 3040
rect 4722 3038 4723 3039
rect 4652 3036 4723 3038
rect 4652 3035 4653 3036
rect 4466 3034 4472 3035
rect 4647 3034 4653 3035
rect 4722 3035 4723 3036
rect 4727 3035 4728 3039
rect 4742 3036 4743 3040
rect 4747 3036 4748 3040
rect 4742 3035 4748 3036
rect 4839 3039 4845 3040
rect 4839 3035 4840 3039
rect 4844 3038 4845 3039
rect 4922 3039 4928 3040
rect 4922 3038 4923 3039
rect 4844 3036 4923 3038
rect 4844 3035 4845 3036
rect 4722 3034 4728 3035
rect 4839 3034 4845 3035
rect 4922 3035 4923 3036
rect 4927 3035 4928 3039
rect 4942 3036 4943 3040
rect 4947 3036 4948 3040
rect 4942 3035 4948 3036
rect 5038 3039 5045 3040
rect 5038 3035 5039 3039
rect 5044 3035 5045 3039
rect 4922 3034 4928 3035
rect 5038 3034 5045 3035
rect 5662 3039 5668 3040
rect 5662 3035 5663 3039
rect 5667 3035 5668 3039
rect 5662 3034 5668 3035
rect 1780 3032 1914 3034
rect 1780 3031 1781 3032
rect 1775 3030 1781 3031
rect 1814 3028 1820 3029
rect 1912 3028 1914 3032
rect 110 3027 116 3028
rect 110 3023 111 3027
rect 115 3023 116 3027
rect 158 3024 159 3028
rect 163 3024 164 3028
rect 158 3023 164 3024
rect 250 3027 261 3028
rect 250 3023 251 3027
rect 255 3023 256 3027
rect 260 3023 261 3027
rect 334 3024 335 3028
rect 339 3024 340 3028
rect 334 3023 340 3024
rect 430 3027 437 3028
rect 430 3023 431 3027
rect 436 3023 437 3027
rect 534 3024 535 3028
rect 539 3024 540 3028
rect 534 3023 540 3024
rect 631 3027 637 3028
rect 631 3023 632 3027
rect 636 3023 637 3027
rect 734 3024 735 3028
rect 739 3024 740 3028
rect 734 3023 740 3024
rect 831 3027 837 3028
rect 831 3023 832 3027
rect 836 3026 837 3027
rect 906 3027 912 3028
rect 906 3026 907 3027
rect 836 3024 907 3026
rect 836 3023 837 3024
rect 110 3022 116 3023
rect 250 3022 261 3023
rect 430 3022 437 3023
rect 631 3022 637 3023
rect 831 3022 837 3023
rect 906 3023 907 3024
rect 911 3023 912 3027
rect 926 3024 927 3028
rect 931 3024 932 3028
rect 926 3023 932 3024
rect 1023 3027 1032 3028
rect 1023 3023 1024 3027
rect 1031 3023 1032 3027
rect 1118 3024 1119 3028
rect 1123 3024 1124 3028
rect 1118 3023 1124 3024
rect 1215 3027 1221 3028
rect 1215 3023 1216 3027
rect 1220 3026 1221 3027
rect 1282 3027 1288 3028
rect 1282 3026 1283 3027
rect 1220 3024 1283 3026
rect 1220 3023 1221 3024
rect 906 3022 912 3023
rect 1023 3022 1032 3023
rect 1215 3022 1221 3023
rect 1282 3023 1283 3024
rect 1287 3023 1288 3027
rect 1302 3024 1303 3028
rect 1307 3024 1308 3028
rect 1302 3023 1308 3024
rect 1399 3027 1405 3028
rect 1399 3023 1400 3027
rect 1404 3026 1405 3027
rect 1458 3027 1464 3028
rect 1458 3026 1459 3027
rect 1404 3024 1459 3026
rect 1404 3023 1405 3024
rect 1282 3022 1288 3023
rect 1399 3022 1405 3023
rect 1458 3023 1459 3024
rect 1463 3023 1464 3027
rect 1478 3024 1479 3028
rect 1483 3024 1484 3028
rect 1478 3023 1484 3024
rect 1574 3027 1581 3028
rect 1574 3023 1575 3027
rect 1580 3023 1581 3027
rect 1654 3024 1655 3028
rect 1659 3024 1660 3028
rect 1654 3023 1660 3024
rect 1751 3027 1757 3028
rect 1751 3023 1752 3027
rect 1756 3023 1757 3027
rect 1814 3024 1815 3028
rect 1819 3024 1820 3028
rect 1814 3023 1820 3024
rect 1911 3027 1917 3028
rect 1911 3023 1912 3027
rect 1916 3023 1917 3027
rect 1458 3022 1464 3023
rect 1574 3022 1581 3023
rect 1751 3022 1757 3023
rect 1911 3022 1917 3023
rect 1934 3027 1940 3028
rect 1934 3023 1935 3027
rect 1939 3023 1940 3027
rect 1934 3022 1940 3023
rect 1974 2989 1980 2990
rect 3798 2989 3804 2990
rect 1974 2985 1975 2989
rect 1979 2985 1980 2989
rect 1974 2984 1980 2985
rect 2190 2988 2196 2989
rect 2350 2988 2356 2989
rect 2518 2988 2524 2989
rect 2702 2988 2708 2989
rect 2902 2988 2908 2989
rect 3118 2988 3124 2989
rect 3334 2988 3340 2989
rect 3558 2988 3564 2989
rect 2190 2984 2191 2988
rect 2195 2984 2196 2988
rect 2190 2983 2196 2984
rect 2286 2987 2293 2988
rect 2286 2983 2287 2987
rect 2292 2983 2293 2987
rect 2350 2984 2351 2988
rect 2355 2984 2356 2988
rect 2350 2983 2356 2984
rect 2446 2987 2453 2988
rect 2446 2983 2447 2987
rect 2452 2983 2453 2987
rect 2518 2984 2519 2988
rect 2523 2984 2524 2988
rect 2518 2983 2524 2984
rect 2615 2987 2621 2988
rect 2615 2983 2616 2987
rect 2620 2986 2621 2987
rect 2638 2987 2644 2988
rect 2638 2986 2639 2987
rect 2620 2984 2639 2986
rect 2620 2983 2621 2984
rect 2286 2982 2293 2983
rect 2446 2982 2453 2983
rect 2615 2982 2621 2983
rect 2638 2983 2639 2984
rect 2643 2983 2644 2987
rect 2702 2984 2703 2988
rect 2707 2984 2708 2988
rect 2702 2983 2708 2984
rect 2794 2987 2805 2988
rect 2794 2983 2795 2987
rect 2799 2983 2800 2987
rect 2804 2983 2805 2987
rect 2902 2984 2903 2988
rect 2907 2984 2908 2988
rect 2902 2983 2908 2984
rect 2999 2987 3008 2988
rect 2999 2983 3000 2987
rect 3007 2983 3008 2987
rect 3118 2984 3119 2988
rect 3123 2984 3124 2988
rect 3118 2983 3124 2984
rect 3214 2987 3221 2988
rect 3214 2983 3215 2987
rect 3220 2983 3221 2987
rect 3334 2984 3335 2988
rect 3339 2984 3340 2988
rect 3334 2983 3340 2984
rect 3426 2987 3437 2988
rect 3426 2983 3427 2987
rect 3431 2983 3432 2987
rect 3436 2983 3437 2987
rect 3558 2984 3559 2988
rect 3563 2984 3564 2988
rect 3558 2983 3564 2984
rect 3650 2987 3661 2988
rect 3650 2983 3651 2987
rect 3655 2983 3656 2987
rect 3660 2983 3661 2987
rect 3798 2985 3799 2989
rect 3803 2985 3804 2989
rect 3798 2984 3804 2985
rect 2638 2982 2644 2983
rect 2794 2982 2805 2983
rect 2999 2982 3008 2983
rect 3214 2982 3221 2983
rect 3426 2982 3437 2983
rect 3650 2982 3661 2983
rect 2162 2973 2168 2974
rect 1974 2972 1980 2973
rect 1974 2968 1975 2972
rect 1979 2968 1980 2972
rect 2162 2969 2163 2973
rect 2167 2969 2168 2973
rect 2162 2968 2168 2969
rect 2322 2973 2328 2974
rect 2322 2969 2323 2973
rect 2327 2969 2328 2973
rect 2322 2968 2328 2969
rect 2490 2973 2496 2974
rect 2490 2969 2491 2973
rect 2495 2969 2496 2973
rect 2490 2968 2496 2969
rect 2674 2973 2680 2974
rect 2674 2969 2675 2973
rect 2679 2969 2680 2973
rect 2674 2968 2680 2969
rect 2874 2973 2880 2974
rect 2874 2969 2875 2973
rect 2879 2969 2880 2973
rect 2874 2968 2880 2969
rect 3090 2973 3096 2974
rect 3090 2969 3091 2973
rect 3095 2969 3096 2973
rect 3090 2968 3096 2969
rect 3306 2973 3312 2974
rect 3306 2969 3307 2973
rect 3311 2969 3312 2973
rect 3306 2968 3312 2969
rect 3530 2973 3536 2974
rect 3530 2969 3531 2973
rect 3535 2969 3536 2973
rect 3530 2968 3536 2969
rect 3798 2972 3804 2973
rect 3798 2968 3799 2972
rect 3803 2968 3804 2972
rect 1974 2967 1980 2968
rect 3798 2967 3804 2968
rect 110 2965 116 2966
rect 1934 2965 1940 2966
rect 110 2961 111 2965
rect 115 2961 116 2965
rect 110 2960 116 2961
rect 158 2964 164 2965
rect 294 2964 300 2965
rect 430 2964 436 2965
rect 566 2964 572 2965
rect 702 2964 708 2965
rect 158 2960 159 2964
rect 163 2960 164 2964
rect 158 2959 164 2960
rect 255 2963 261 2964
rect 255 2959 256 2963
rect 260 2962 261 2963
rect 263 2963 269 2964
rect 263 2962 264 2963
rect 260 2960 264 2962
rect 260 2959 261 2960
rect 255 2958 261 2959
rect 263 2959 264 2960
rect 268 2959 269 2963
rect 294 2960 295 2964
rect 299 2960 300 2964
rect 294 2959 300 2960
rect 391 2963 400 2964
rect 391 2959 392 2963
rect 399 2959 400 2963
rect 430 2960 431 2964
rect 435 2960 436 2964
rect 430 2959 436 2960
rect 527 2963 536 2964
rect 527 2959 528 2963
rect 535 2959 536 2963
rect 566 2960 567 2964
rect 571 2960 572 2964
rect 566 2959 572 2960
rect 658 2963 669 2964
rect 658 2959 659 2963
rect 663 2959 664 2963
rect 668 2959 669 2963
rect 702 2960 703 2964
rect 707 2960 708 2964
rect 702 2959 708 2960
rect 799 2963 808 2964
rect 799 2959 800 2963
rect 807 2959 808 2963
rect 1934 2961 1935 2965
rect 1939 2961 1940 2965
rect 1934 2960 1940 2961
rect 263 2958 269 2959
rect 391 2958 400 2959
rect 527 2958 536 2959
rect 658 2958 669 2959
rect 799 2958 808 2959
rect 3838 2957 3844 2958
rect 5662 2957 5668 2958
rect 3838 2953 3839 2957
rect 3843 2953 3844 2957
rect 3838 2952 3844 2953
rect 3998 2956 4004 2957
rect 4158 2956 4164 2957
rect 4334 2956 4340 2957
rect 4518 2956 4524 2957
rect 4718 2956 4724 2957
rect 4926 2956 4932 2957
rect 5134 2956 5140 2957
rect 5350 2956 5356 2957
rect 5542 2956 5548 2957
rect 3998 2952 3999 2956
rect 4003 2952 4004 2956
rect 2258 2951 2264 2952
rect 130 2949 136 2950
rect 110 2948 116 2949
rect 110 2944 111 2948
rect 115 2944 116 2948
rect 130 2945 131 2949
rect 135 2945 136 2949
rect 130 2944 136 2945
rect 266 2949 272 2950
rect 266 2945 267 2949
rect 271 2945 272 2949
rect 266 2944 272 2945
rect 402 2949 408 2950
rect 402 2945 403 2949
rect 407 2945 408 2949
rect 402 2944 408 2945
rect 538 2949 544 2950
rect 538 2945 539 2949
rect 543 2945 544 2949
rect 538 2944 544 2945
rect 674 2949 680 2950
rect 674 2945 675 2949
rect 679 2945 680 2949
rect 674 2944 680 2945
rect 1934 2948 1940 2949
rect 1934 2944 1935 2948
rect 1939 2944 1940 2948
rect 2258 2947 2259 2951
rect 2263 2950 2264 2951
rect 2446 2951 2452 2952
rect 3998 2951 4004 2952
rect 4094 2955 4101 2956
rect 4094 2951 4095 2955
rect 4100 2951 4101 2955
rect 4158 2952 4159 2956
rect 4163 2952 4164 2956
rect 4158 2951 4164 2952
rect 4255 2955 4261 2956
rect 4255 2951 4256 2955
rect 4260 2954 4261 2955
rect 4271 2955 4277 2956
rect 4271 2954 4272 2955
rect 4260 2952 4272 2954
rect 4260 2951 4261 2952
rect 2446 2950 2447 2951
rect 2263 2948 2447 2950
rect 2263 2947 2264 2948
rect 2258 2946 2264 2947
rect 2446 2947 2447 2948
rect 2451 2947 2452 2951
rect 4094 2950 4101 2951
rect 4255 2950 4261 2951
rect 4271 2951 4272 2952
rect 4276 2951 4277 2955
rect 4334 2952 4335 2956
rect 4339 2952 4340 2956
rect 4334 2951 4340 2952
rect 4431 2955 4437 2956
rect 4431 2951 4432 2955
rect 4436 2954 4437 2955
rect 4442 2955 4448 2956
rect 4442 2954 4443 2955
rect 4436 2952 4443 2954
rect 4436 2951 4437 2952
rect 4271 2950 4277 2951
rect 4431 2950 4437 2951
rect 4442 2951 4443 2952
rect 4447 2951 4448 2955
rect 4518 2952 4519 2956
rect 4523 2952 4524 2956
rect 4518 2951 4524 2952
rect 4615 2955 4624 2956
rect 4615 2951 4616 2955
rect 4623 2951 4624 2955
rect 4718 2952 4719 2956
rect 4723 2952 4724 2956
rect 4718 2951 4724 2952
rect 4815 2955 4824 2956
rect 4815 2951 4816 2955
rect 4823 2951 4824 2955
rect 4926 2952 4927 2956
rect 4931 2952 4932 2956
rect 4926 2951 4932 2952
rect 5018 2955 5029 2956
rect 5018 2951 5019 2955
rect 5023 2951 5024 2955
rect 5028 2951 5029 2955
rect 5134 2952 5135 2956
rect 5139 2952 5140 2956
rect 5134 2951 5140 2952
rect 5231 2955 5237 2956
rect 5231 2951 5232 2955
rect 5236 2954 5237 2955
rect 5286 2955 5292 2956
rect 5286 2954 5287 2955
rect 5236 2952 5287 2954
rect 5236 2951 5237 2952
rect 4442 2950 4448 2951
rect 4615 2950 4624 2951
rect 4815 2950 4824 2951
rect 5018 2950 5029 2951
rect 5231 2950 5237 2951
rect 5286 2951 5287 2952
rect 5291 2951 5292 2955
rect 5350 2952 5351 2956
rect 5355 2952 5356 2956
rect 5350 2951 5356 2952
rect 5447 2955 5453 2956
rect 5447 2951 5448 2955
rect 5452 2954 5453 2955
rect 5482 2955 5488 2956
rect 5482 2954 5483 2955
rect 5452 2952 5483 2954
rect 5452 2951 5453 2952
rect 5286 2950 5292 2951
rect 5447 2950 5453 2951
rect 5482 2951 5483 2952
rect 5487 2951 5488 2955
rect 5542 2952 5543 2956
rect 5547 2952 5548 2956
rect 5542 2951 5548 2952
rect 5634 2955 5645 2956
rect 5634 2951 5635 2955
rect 5639 2951 5640 2955
rect 5644 2951 5645 2955
rect 5662 2953 5663 2957
rect 5667 2953 5668 2957
rect 5662 2952 5668 2953
rect 5482 2950 5488 2951
rect 5634 2950 5645 2951
rect 2446 2946 2452 2947
rect 110 2943 116 2944
rect 1934 2943 1940 2944
rect 3970 2941 3976 2942
rect 3838 2940 3844 2941
rect 3838 2936 3839 2940
rect 3843 2936 3844 2940
rect 3970 2937 3971 2941
rect 3975 2937 3976 2941
rect 3970 2936 3976 2937
rect 4130 2941 4136 2942
rect 4130 2937 4131 2941
rect 4135 2937 4136 2941
rect 4130 2936 4136 2937
rect 4306 2941 4312 2942
rect 4306 2937 4307 2941
rect 4311 2937 4312 2941
rect 4306 2936 4312 2937
rect 4490 2941 4496 2942
rect 4490 2937 4491 2941
rect 4495 2937 4496 2941
rect 4490 2936 4496 2937
rect 4690 2941 4696 2942
rect 4690 2937 4691 2941
rect 4695 2937 4696 2941
rect 4690 2936 4696 2937
rect 4898 2941 4904 2942
rect 4898 2937 4899 2941
rect 4903 2937 4904 2941
rect 4898 2936 4904 2937
rect 5106 2941 5112 2942
rect 5106 2937 5107 2941
rect 5111 2937 5112 2941
rect 5106 2936 5112 2937
rect 5322 2941 5328 2942
rect 5322 2937 5323 2941
rect 5327 2937 5328 2941
rect 5322 2936 5328 2937
rect 5514 2941 5520 2942
rect 5514 2937 5515 2941
rect 5519 2937 5520 2941
rect 5514 2936 5520 2937
rect 5662 2940 5668 2941
rect 5662 2936 5663 2940
rect 5667 2936 5668 2940
rect 3838 2935 3844 2936
rect 5662 2935 5668 2936
rect 2258 2923 2264 2924
rect 2258 2919 2259 2923
rect 2263 2919 2264 2923
rect 2606 2923 2612 2924
rect 2606 2922 2607 2923
rect 2258 2918 2264 2919
rect 2420 2914 2422 2921
rect 2589 2920 2607 2922
rect 2606 2919 2607 2920
rect 2611 2919 2612 2923
rect 2606 2918 2612 2919
rect 2638 2923 2644 2924
rect 2638 2919 2639 2923
rect 2643 2922 2644 2923
rect 2958 2923 2964 2924
rect 2643 2920 2681 2922
rect 2643 2919 2644 2920
rect 2638 2918 2644 2919
rect 2958 2919 2959 2923
rect 2963 2919 2964 2923
rect 2958 2918 2964 2919
rect 3002 2923 3008 2924
rect 3002 2919 3003 2923
rect 3007 2922 3008 2923
rect 3770 2923 3776 2924
rect 3770 2922 3771 2923
rect 3007 2920 3097 2922
rect 3007 2919 3008 2920
rect 3002 2918 3008 2919
rect 2794 2915 2800 2916
rect 2794 2914 2795 2915
rect 2420 2912 2795 2914
rect 2794 2911 2795 2912
rect 2799 2911 2800 2915
rect 3404 2914 3406 2921
rect 3629 2920 3771 2922
rect 3770 2919 3771 2920
rect 3775 2919 3776 2923
rect 3770 2918 3776 2919
rect 3650 2915 3656 2916
rect 3650 2914 3651 2915
rect 3404 2912 3651 2914
rect 2794 2910 2800 2911
rect 3650 2911 3651 2912
rect 3655 2911 3656 2915
rect 3650 2910 3656 2911
rect 250 2899 256 2900
rect 250 2898 251 2899
rect 229 2896 251 2898
rect 250 2895 251 2896
rect 255 2895 256 2899
rect 250 2894 256 2895
rect 263 2899 269 2900
rect 263 2895 264 2899
rect 268 2898 269 2899
rect 394 2899 400 2900
rect 268 2896 273 2898
rect 268 2895 269 2896
rect 263 2894 269 2895
rect 394 2895 395 2899
rect 399 2898 400 2899
rect 530 2899 536 2900
rect 399 2896 409 2898
rect 399 2895 400 2896
rect 394 2894 400 2895
rect 530 2895 531 2899
rect 535 2898 536 2899
rect 758 2899 764 2900
rect 535 2896 545 2898
rect 535 2895 536 2896
rect 530 2894 536 2895
rect 758 2895 759 2899
rect 763 2895 764 2899
rect 758 2894 764 2895
rect 3982 2891 3988 2892
rect 2286 2887 2292 2888
rect 2090 2883 2096 2884
rect 2090 2879 2091 2883
rect 2095 2879 2096 2883
rect 2090 2878 2096 2879
rect 2138 2883 2144 2884
rect 2138 2879 2139 2883
rect 2143 2879 2144 2883
rect 2286 2883 2287 2887
rect 2291 2883 2292 2887
rect 2718 2887 2724 2888
rect 2286 2882 2292 2883
rect 2410 2883 2416 2884
rect 2138 2878 2144 2879
rect 2410 2879 2411 2883
rect 2415 2879 2416 2883
rect 2410 2878 2416 2879
rect 2546 2883 2552 2884
rect 2546 2879 2547 2883
rect 2551 2879 2552 2883
rect 2718 2883 2719 2887
rect 2723 2883 2724 2887
rect 3146 2887 3152 2888
rect 3146 2886 3147 2887
rect 3093 2884 3147 2886
rect 2718 2882 2724 2883
rect 2842 2883 2848 2884
rect 2546 2878 2552 2879
rect 2842 2879 2843 2883
rect 2847 2879 2848 2883
rect 3146 2883 3147 2884
rect 3151 2883 3152 2887
rect 3306 2887 3312 2888
rect 3306 2886 3307 2887
rect 3253 2884 3307 2886
rect 3146 2882 3152 2883
rect 3306 2883 3307 2884
rect 3311 2883 3312 2887
rect 3426 2887 3432 2888
rect 3426 2886 3427 2887
rect 3413 2884 3427 2886
rect 3306 2882 3312 2883
rect 3426 2883 3427 2884
rect 3431 2883 3432 2887
rect 3982 2887 3983 2891
rect 3987 2887 3988 2891
rect 4271 2891 4277 2892
rect 3982 2886 3988 2887
rect 3426 2882 3432 2883
rect 4228 2882 4230 2889
rect 4271 2887 4272 2891
rect 4276 2890 4277 2891
rect 4466 2891 4472 2892
rect 4276 2888 4313 2890
rect 4276 2887 4277 2888
rect 4271 2886 4277 2887
rect 4466 2887 4467 2891
rect 4471 2890 4472 2891
rect 4618 2891 4624 2892
rect 4471 2888 4497 2890
rect 4471 2887 4472 2888
rect 4466 2886 4472 2887
rect 4618 2887 4619 2891
rect 4623 2890 4624 2891
rect 4818 2891 4824 2892
rect 4623 2888 4697 2890
rect 4623 2887 4624 2888
rect 4618 2886 4624 2887
rect 4818 2887 4819 2891
rect 4823 2890 4824 2891
rect 5286 2891 5292 2892
rect 4823 2888 4905 2890
rect 4823 2887 4824 2888
rect 4818 2886 4824 2887
rect 5018 2883 5024 2884
rect 5018 2882 5019 2883
rect 4228 2880 5019 2882
rect 2842 2878 2848 2879
rect 5018 2879 5019 2880
rect 5023 2879 5024 2883
rect 5204 2882 5206 2889
rect 5286 2887 5287 2891
rect 5291 2890 5292 2891
rect 5482 2891 5488 2892
rect 5291 2888 5329 2890
rect 5291 2887 5292 2888
rect 5286 2886 5292 2887
rect 5482 2887 5483 2891
rect 5487 2890 5488 2891
rect 5487 2888 5521 2890
rect 5487 2887 5488 2888
rect 5482 2886 5488 2887
rect 5374 2883 5380 2884
rect 5374 2882 5375 2883
rect 5204 2880 5375 2882
rect 5018 2878 5024 2879
rect 5374 2879 5375 2880
rect 5379 2879 5380 2883
rect 5374 2878 5380 2879
rect 658 2871 664 2872
rect 658 2867 659 2871
rect 663 2867 664 2871
rect 658 2866 664 2867
rect 364 2864 662 2866
rect 364 2862 366 2864
rect 767 2863 773 2864
rect 767 2862 768 2863
rect 325 2860 366 2862
rect 733 2860 768 2862
rect 370 2859 376 2860
rect 370 2855 371 2859
rect 375 2855 376 2859
rect 370 2854 376 2855
rect 506 2859 512 2860
rect 506 2855 507 2859
rect 511 2855 512 2859
rect 767 2859 768 2860
rect 772 2859 773 2863
rect 894 2863 900 2864
rect 894 2862 895 2863
rect 869 2860 895 2862
rect 767 2858 773 2859
rect 894 2859 895 2860
rect 899 2859 900 2863
rect 894 2858 900 2859
rect 506 2854 512 2855
rect 2090 2855 2096 2856
rect 2090 2851 2091 2855
rect 2095 2854 2096 2855
rect 2662 2855 2668 2856
rect 2662 2854 2663 2855
rect 2095 2852 2663 2854
rect 2095 2851 2096 2852
rect 2090 2850 2096 2851
rect 2662 2851 2663 2852
rect 2667 2851 2668 2855
rect 2662 2850 2668 2851
rect 4202 2843 4208 2844
rect 4202 2842 4203 2843
rect 4109 2840 4203 2842
rect 3954 2839 3960 2840
rect 1974 2836 1980 2837
rect 3798 2836 3804 2837
rect 1974 2832 1975 2836
rect 1979 2832 1980 2836
rect 1974 2831 1980 2832
rect 1994 2835 2000 2836
rect 1994 2831 1995 2835
rect 1999 2831 2000 2835
rect 1994 2830 2000 2831
rect 2130 2835 2136 2836
rect 2130 2831 2131 2835
rect 2135 2831 2136 2835
rect 2130 2830 2136 2831
rect 2266 2835 2272 2836
rect 2266 2831 2267 2835
rect 2271 2831 2272 2835
rect 2266 2830 2272 2831
rect 2402 2835 2408 2836
rect 2402 2831 2403 2835
rect 2407 2831 2408 2835
rect 2402 2830 2408 2831
rect 2538 2835 2544 2836
rect 2538 2831 2539 2835
rect 2543 2831 2544 2835
rect 2538 2830 2544 2831
rect 2682 2835 2688 2836
rect 2682 2831 2683 2835
rect 2687 2831 2688 2835
rect 2682 2830 2688 2831
rect 2834 2835 2840 2836
rect 2834 2831 2835 2835
rect 2839 2831 2840 2835
rect 2834 2830 2840 2831
rect 2994 2835 3000 2836
rect 2994 2831 2995 2835
rect 2999 2831 3000 2835
rect 2994 2830 3000 2831
rect 3154 2835 3160 2836
rect 3154 2831 3155 2835
rect 3159 2831 3160 2835
rect 3154 2830 3160 2831
rect 3314 2835 3320 2836
rect 3314 2831 3315 2835
rect 3319 2831 3320 2835
rect 3798 2832 3799 2836
rect 3803 2832 3804 2836
rect 3954 2835 3955 2839
rect 3959 2835 3960 2839
rect 4202 2839 4203 2840
rect 4207 2839 4208 2843
rect 4359 2843 4365 2844
rect 4359 2842 4360 2843
rect 4309 2840 4360 2842
rect 4202 2838 4208 2839
rect 4359 2839 4360 2840
rect 4364 2839 4365 2843
rect 4359 2838 4365 2839
rect 4442 2843 4448 2844
rect 4442 2839 4443 2843
rect 4447 2839 4448 2843
rect 5390 2843 5396 2844
rect 5390 2842 5391 2843
rect 5349 2840 5391 2842
rect 4442 2838 4448 2839
rect 4698 2839 4704 2840
rect 3954 2834 3960 2835
rect 4698 2835 4699 2839
rect 4703 2835 4704 2839
rect 4698 2834 4704 2835
rect 4970 2839 4976 2840
rect 4970 2835 4971 2839
rect 4975 2835 4976 2839
rect 5390 2839 5391 2840
rect 5395 2839 5396 2843
rect 5634 2843 5640 2844
rect 5634 2842 5635 2843
rect 5613 2840 5635 2842
rect 5390 2838 5396 2839
rect 5634 2839 5635 2840
rect 5639 2839 5640 2843
rect 5634 2838 5640 2839
rect 4970 2834 4976 2835
rect 3798 2831 3804 2832
rect 3314 2830 3320 2831
rect 3146 2827 3152 2828
rect 3146 2823 3147 2827
rect 3151 2826 3152 2827
rect 3306 2827 3312 2828
rect 3151 2824 3282 2826
rect 3151 2823 3152 2824
rect 3146 2822 3152 2823
rect 2022 2820 2028 2821
rect 2158 2820 2164 2821
rect 2294 2820 2300 2821
rect 2430 2820 2436 2821
rect 2566 2820 2572 2821
rect 2710 2820 2716 2821
rect 2862 2820 2868 2821
rect 3022 2820 3028 2821
rect 3182 2820 3188 2821
rect 3280 2820 3282 2824
rect 3306 2823 3307 2827
rect 3311 2826 3312 2827
rect 3311 2824 3442 2826
rect 3311 2823 3312 2824
rect 3306 2822 3312 2823
rect 3342 2820 3348 2821
rect 3440 2820 3442 2824
rect 1974 2819 1980 2820
rect 1974 2815 1975 2819
rect 1979 2815 1980 2819
rect 2022 2816 2023 2820
rect 2027 2816 2028 2820
rect 2022 2815 2028 2816
rect 2119 2819 2125 2820
rect 2119 2815 2120 2819
rect 2124 2818 2125 2819
rect 2138 2819 2144 2820
rect 2138 2818 2139 2819
rect 2124 2816 2139 2818
rect 2124 2815 2125 2816
rect 1974 2814 1980 2815
rect 2119 2814 2125 2815
rect 2138 2815 2139 2816
rect 2143 2815 2144 2819
rect 2158 2816 2159 2820
rect 2163 2816 2164 2820
rect 2158 2815 2164 2816
rect 2250 2819 2261 2820
rect 2250 2815 2251 2819
rect 2255 2815 2256 2819
rect 2260 2815 2261 2819
rect 2294 2816 2295 2820
rect 2299 2816 2300 2820
rect 2294 2815 2300 2816
rect 2391 2819 2397 2820
rect 2391 2815 2392 2819
rect 2396 2818 2397 2819
rect 2410 2819 2416 2820
rect 2410 2818 2411 2819
rect 2396 2816 2411 2818
rect 2396 2815 2397 2816
rect 2138 2814 2144 2815
rect 2250 2814 2261 2815
rect 2391 2814 2397 2815
rect 2410 2815 2411 2816
rect 2415 2815 2416 2819
rect 2430 2816 2431 2820
rect 2435 2816 2436 2820
rect 2430 2815 2436 2816
rect 2527 2819 2533 2820
rect 2527 2815 2528 2819
rect 2532 2818 2533 2819
rect 2546 2819 2552 2820
rect 2546 2818 2547 2819
rect 2532 2816 2547 2818
rect 2532 2815 2533 2816
rect 2410 2814 2416 2815
rect 2527 2814 2533 2815
rect 2546 2815 2547 2816
rect 2551 2815 2552 2819
rect 2566 2816 2567 2820
rect 2571 2816 2572 2820
rect 2566 2815 2572 2816
rect 2662 2819 2669 2820
rect 2662 2815 2663 2819
rect 2668 2815 2669 2819
rect 2710 2816 2711 2820
rect 2715 2816 2716 2820
rect 2710 2815 2716 2816
rect 2807 2819 2813 2820
rect 2807 2815 2808 2819
rect 2812 2818 2813 2819
rect 2842 2819 2848 2820
rect 2842 2818 2843 2819
rect 2812 2816 2843 2818
rect 2812 2815 2813 2816
rect 2546 2814 2552 2815
rect 2662 2814 2669 2815
rect 2807 2814 2813 2815
rect 2842 2815 2843 2816
rect 2847 2815 2848 2819
rect 2862 2816 2863 2820
rect 2867 2816 2868 2820
rect 2862 2815 2868 2816
rect 2958 2819 2965 2820
rect 2958 2815 2959 2819
rect 2964 2815 2965 2819
rect 3022 2816 3023 2820
rect 3027 2816 3028 2820
rect 3022 2815 3028 2816
rect 3118 2819 3125 2820
rect 3118 2815 3119 2819
rect 3124 2815 3125 2819
rect 3182 2816 3183 2820
rect 3187 2816 3188 2820
rect 3182 2815 3188 2816
rect 3279 2819 3285 2820
rect 3279 2815 3280 2819
rect 3284 2815 3285 2819
rect 3342 2816 3343 2820
rect 3347 2816 3348 2820
rect 3342 2815 3348 2816
rect 3439 2819 3445 2820
rect 3439 2815 3440 2819
rect 3444 2815 3445 2819
rect 2842 2814 2848 2815
rect 2958 2814 2965 2815
rect 3118 2814 3125 2815
rect 3279 2814 3285 2815
rect 3439 2814 3445 2815
rect 3798 2819 3804 2820
rect 3798 2815 3799 2819
rect 3803 2815 3804 2819
rect 3798 2814 3804 2815
rect 110 2812 116 2813
rect 1934 2812 1940 2813
rect 110 2808 111 2812
rect 115 2808 116 2812
rect 110 2807 116 2808
rect 226 2811 232 2812
rect 226 2807 227 2811
rect 231 2807 232 2811
rect 226 2806 232 2807
rect 362 2811 368 2812
rect 362 2807 363 2811
rect 367 2807 368 2811
rect 362 2806 368 2807
rect 498 2811 504 2812
rect 498 2807 499 2811
rect 503 2807 504 2811
rect 498 2806 504 2807
rect 634 2811 640 2812
rect 634 2807 635 2811
rect 639 2807 640 2811
rect 634 2806 640 2807
rect 770 2811 776 2812
rect 770 2807 771 2811
rect 775 2807 776 2811
rect 1934 2808 1935 2812
rect 1939 2808 1940 2812
rect 1934 2807 1940 2808
rect 770 2806 776 2807
rect 792 2800 891 2802
rect 767 2799 773 2800
rect 254 2796 260 2797
rect 390 2796 396 2797
rect 526 2796 532 2797
rect 662 2796 668 2797
rect 110 2795 116 2796
rect 110 2791 111 2795
rect 115 2791 116 2795
rect 254 2792 255 2796
rect 259 2792 260 2796
rect 254 2791 260 2792
rect 351 2795 357 2796
rect 351 2791 352 2795
rect 356 2794 357 2795
rect 370 2795 376 2796
rect 370 2794 371 2795
rect 356 2792 371 2794
rect 356 2791 357 2792
rect 110 2790 116 2791
rect 351 2790 357 2791
rect 370 2791 371 2792
rect 375 2791 376 2795
rect 390 2792 391 2796
rect 395 2792 396 2796
rect 390 2791 396 2792
rect 487 2795 493 2796
rect 487 2791 488 2795
rect 492 2794 493 2795
rect 506 2795 512 2796
rect 506 2794 507 2795
rect 492 2792 507 2794
rect 492 2791 493 2792
rect 370 2790 376 2791
rect 487 2790 493 2791
rect 506 2791 507 2792
rect 511 2791 512 2795
rect 526 2792 527 2796
rect 531 2792 532 2796
rect 526 2791 532 2792
rect 623 2795 629 2796
rect 623 2791 624 2795
rect 628 2794 629 2795
rect 628 2792 638 2794
rect 628 2791 629 2792
rect 506 2790 512 2791
rect 623 2790 629 2791
rect 636 2778 638 2792
rect 662 2792 663 2796
rect 667 2792 668 2796
rect 662 2791 668 2792
rect 758 2795 765 2796
rect 758 2791 759 2795
rect 764 2791 765 2795
rect 767 2795 768 2799
rect 772 2798 773 2799
rect 792 2798 794 2800
rect 772 2796 794 2798
rect 798 2796 804 2797
rect 772 2795 773 2796
rect 767 2794 773 2795
rect 798 2792 799 2796
rect 803 2792 804 2796
rect 889 2794 891 2800
rect 895 2795 901 2796
rect 895 2794 896 2795
rect 889 2792 896 2794
rect 798 2791 804 2792
rect 895 2791 896 2792
rect 900 2791 901 2795
rect 758 2790 765 2791
rect 895 2790 901 2791
rect 1934 2795 1940 2796
rect 1934 2791 1935 2795
rect 1939 2791 1940 2795
rect 1934 2790 1940 2791
rect 3838 2792 3844 2793
rect 5662 2792 5668 2793
rect 3838 2788 3839 2792
rect 3843 2788 3844 2792
rect 3838 2787 3844 2788
rect 3858 2791 3864 2792
rect 3858 2787 3859 2791
rect 3863 2787 3864 2791
rect 3858 2786 3864 2787
rect 4010 2791 4016 2792
rect 4010 2787 4011 2791
rect 4015 2787 4016 2791
rect 4010 2786 4016 2787
rect 4210 2791 4216 2792
rect 4210 2787 4211 2791
rect 4215 2787 4216 2791
rect 4210 2786 4216 2787
rect 4434 2791 4440 2792
rect 4434 2787 4435 2791
rect 4439 2787 4440 2791
rect 4434 2786 4440 2787
rect 4690 2791 4696 2792
rect 4690 2787 4691 2791
rect 4695 2787 4696 2791
rect 4690 2786 4696 2787
rect 4962 2791 4968 2792
rect 4962 2787 4963 2791
rect 4967 2787 4968 2791
rect 4962 2786 4968 2787
rect 5250 2791 5256 2792
rect 5250 2787 5251 2791
rect 5255 2787 5256 2791
rect 5250 2786 5256 2787
rect 5514 2791 5520 2792
rect 5514 2787 5515 2791
rect 5519 2787 5520 2791
rect 5662 2788 5663 2792
rect 5667 2788 5668 2792
rect 5662 2787 5668 2788
rect 5514 2786 5520 2787
rect 4202 2783 4208 2784
rect 918 2779 924 2780
rect 918 2778 919 2779
rect 636 2776 919 2778
rect 918 2775 919 2776
rect 923 2775 924 2779
rect 4202 2779 4203 2783
rect 4207 2782 4208 2783
rect 4359 2783 4365 2784
rect 4207 2780 4338 2782
rect 4207 2779 4208 2780
rect 4202 2778 4208 2779
rect 4336 2778 4338 2780
rect 4359 2779 4360 2783
rect 4364 2782 4365 2783
rect 4364 2780 5090 2782
rect 4364 2779 4365 2780
rect 4359 2778 4365 2779
rect 4335 2777 4341 2778
rect 3886 2776 3892 2777
rect 4038 2776 4044 2777
rect 4238 2776 4244 2777
rect 918 2774 924 2775
rect 3838 2775 3844 2776
rect 3838 2771 3839 2775
rect 3843 2771 3844 2775
rect 3886 2772 3887 2776
rect 3891 2772 3892 2776
rect 3886 2771 3892 2772
rect 3982 2775 3989 2776
rect 3982 2771 3983 2775
rect 3988 2771 3989 2775
rect 4038 2772 4039 2776
rect 4043 2772 4044 2776
rect 4038 2771 4044 2772
rect 4135 2775 4141 2776
rect 4135 2771 4136 2775
rect 4140 2774 4141 2775
rect 4151 2775 4157 2776
rect 4151 2774 4152 2775
rect 4140 2772 4152 2774
rect 4140 2771 4141 2772
rect 3838 2770 3844 2771
rect 3982 2770 3989 2771
rect 4135 2770 4141 2771
rect 4151 2771 4152 2772
rect 4156 2771 4157 2775
rect 4238 2772 4239 2776
rect 4243 2772 4244 2776
rect 4335 2773 4336 2777
rect 4340 2773 4341 2777
rect 4335 2772 4341 2773
rect 4462 2776 4468 2777
rect 4718 2776 4724 2777
rect 4990 2776 4996 2777
rect 5088 2776 5090 2780
rect 5278 2776 5284 2777
rect 5542 2776 5548 2777
rect 4462 2772 4463 2776
rect 4467 2772 4468 2776
rect 4238 2771 4244 2772
rect 4462 2771 4468 2772
rect 4559 2775 4565 2776
rect 4559 2771 4560 2775
rect 4564 2774 4565 2775
rect 4698 2775 4704 2776
rect 4698 2774 4699 2775
rect 4564 2772 4699 2774
rect 4564 2771 4565 2772
rect 4151 2770 4157 2771
rect 4559 2770 4565 2771
rect 4698 2771 4699 2772
rect 4703 2771 4704 2775
rect 4718 2772 4719 2776
rect 4723 2772 4724 2776
rect 4718 2771 4724 2772
rect 4815 2775 4821 2776
rect 4815 2771 4816 2775
rect 4820 2774 4821 2775
rect 4970 2775 4976 2776
rect 4970 2774 4971 2775
rect 4820 2772 4971 2774
rect 4820 2771 4821 2772
rect 4698 2770 4704 2771
rect 4815 2770 4821 2771
rect 4970 2771 4971 2772
rect 4975 2771 4976 2775
rect 4990 2772 4991 2776
rect 4995 2772 4996 2776
rect 4990 2771 4996 2772
rect 5087 2775 5093 2776
rect 5087 2771 5088 2775
rect 5092 2771 5093 2775
rect 5278 2772 5279 2776
rect 5283 2772 5284 2776
rect 5278 2771 5284 2772
rect 5374 2775 5381 2776
rect 5374 2771 5375 2775
rect 5380 2771 5381 2775
rect 5542 2772 5543 2776
rect 5547 2772 5548 2776
rect 5542 2771 5548 2772
rect 5639 2775 5648 2776
rect 5639 2771 5640 2775
rect 5647 2771 5648 2775
rect 4970 2770 4976 2771
rect 5087 2770 5093 2771
rect 5374 2770 5381 2771
rect 5639 2770 5648 2771
rect 5662 2775 5668 2776
rect 5662 2771 5663 2775
rect 5667 2771 5668 2775
rect 5662 2770 5668 2771
rect 1974 2757 1980 2758
rect 3798 2757 3804 2758
rect 1974 2753 1975 2757
rect 1979 2753 1980 2757
rect 1974 2752 1980 2753
rect 2022 2756 2028 2757
rect 2158 2756 2164 2757
rect 2302 2756 2308 2757
rect 2462 2756 2468 2757
rect 2622 2756 2628 2757
rect 2782 2756 2788 2757
rect 2942 2756 2948 2757
rect 3102 2756 3108 2757
rect 2022 2752 2023 2756
rect 2027 2752 2028 2756
rect 2022 2751 2028 2752
rect 2114 2755 2125 2756
rect 2114 2751 2115 2755
rect 2119 2751 2120 2755
rect 2124 2751 2125 2755
rect 2158 2752 2159 2756
rect 2163 2752 2164 2756
rect 2158 2751 2164 2752
rect 2255 2755 2264 2756
rect 2255 2751 2256 2755
rect 2263 2751 2264 2755
rect 2302 2752 2303 2756
rect 2307 2752 2308 2756
rect 2302 2751 2308 2752
rect 2399 2755 2408 2756
rect 2399 2751 2400 2755
rect 2407 2751 2408 2755
rect 2462 2752 2463 2756
rect 2467 2752 2468 2756
rect 2462 2751 2468 2752
rect 2558 2755 2565 2756
rect 2558 2751 2559 2755
rect 2564 2751 2565 2755
rect 2622 2752 2623 2756
rect 2627 2752 2628 2756
rect 2622 2751 2628 2752
rect 2718 2755 2725 2756
rect 2718 2751 2719 2755
rect 2724 2751 2725 2755
rect 2782 2752 2783 2756
rect 2787 2752 2788 2756
rect 2782 2751 2788 2752
rect 2874 2755 2885 2756
rect 2874 2751 2875 2755
rect 2879 2751 2880 2755
rect 2884 2751 2885 2755
rect 2942 2752 2943 2756
rect 2947 2752 2948 2756
rect 2942 2751 2948 2752
rect 3034 2755 3045 2756
rect 3034 2751 3035 2755
rect 3039 2751 3040 2755
rect 3044 2751 3045 2755
rect 3102 2752 3103 2756
rect 3107 2752 3108 2756
rect 3102 2751 3108 2752
rect 3198 2755 3205 2756
rect 3198 2751 3199 2755
rect 3204 2751 3205 2755
rect 3798 2753 3799 2757
rect 3803 2753 3804 2757
rect 3798 2752 3804 2753
rect 2114 2750 2125 2751
rect 2255 2750 2264 2751
rect 2399 2750 2408 2751
rect 2558 2750 2565 2751
rect 2718 2750 2725 2751
rect 2874 2750 2885 2751
rect 3034 2750 3045 2751
rect 3198 2750 3205 2751
rect 3954 2743 3960 2744
rect 1994 2741 2000 2742
rect 1974 2740 1980 2741
rect 1974 2736 1975 2740
rect 1979 2736 1980 2740
rect 1994 2737 1995 2741
rect 1999 2737 2000 2741
rect 1994 2736 2000 2737
rect 2130 2741 2136 2742
rect 2130 2737 2131 2741
rect 2135 2737 2136 2741
rect 2130 2736 2136 2737
rect 2274 2741 2280 2742
rect 2274 2737 2275 2741
rect 2279 2737 2280 2741
rect 2274 2736 2280 2737
rect 2434 2741 2440 2742
rect 2434 2737 2435 2741
rect 2439 2737 2440 2741
rect 2434 2736 2440 2737
rect 2594 2741 2600 2742
rect 2594 2737 2595 2741
rect 2599 2737 2600 2741
rect 2594 2736 2600 2737
rect 2754 2741 2760 2742
rect 2754 2737 2755 2741
rect 2759 2737 2760 2741
rect 2754 2736 2760 2737
rect 2914 2741 2920 2742
rect 2914 2737 2915 2741
rect 2919 2737 2920 2741
rect 2914 2736 2920 2737
rect 3074 2741 3080 2742
rect 3074 2737 3075 2741
rect 3079 2737 3080 2741
rect 3074 2736 3080 2737
rect 3798 2740 3804 2741
rect 3798 2736 3799 2740
rect 3803 2736 3804 2740
rect 3954 2739 3955 2743
rect 3959 2742 3960 2743
rect 4062 2743 4068 2744
rect 4062 2742 4063 2743
rect 3959 2740 4063 2742
rect 3959 2739 3960 2740
rect 3954 2738 3960 2739
rect 4062 2739 4063 2740
rect 4067 2739 4068 2743
rect 4062 2738 4068 2739
rect 1974 2735 1980 2736
rect 3798 2735 3804 2736
rect 110 2733 116 2734
rect 1934 2733 1940 2734
rect 110 2729 111 2733
rect 115 2729 116 2733
rect 110 2728 116 2729
rect 374 2732 380 2733
rect 574 2732 580 2733
rect 798 2732 804 2733
rect 1038 2732 1044 2733
rect 1294 2732 1300 2733
rect 1566 2732 1572 2733
rect 1814 2732 1820 2733
rect 374 2728 375 2732
rect 379 2728 380 2732
rect 374 2727 380 2728
rect 471 2731 480 2732
rect 471 2727 472 2731
rect 479 2727 480 2731
rect 574 2728 575 2732
rect 579 2728 580 2732
rect 574 2727 580 2728
rect 671 2731 680 2732
rect 671 2727 672 2731
rect 679 2727 680 2731
rect 798 2728 799 2732
rect 803 2728 804 2732
rect 798 2727 804 2728
rect 894 2731 901 2732
rect 894 2727 895 2731
rect 900 2727 901 2731
rect 1038 2728 1039 2732
rect 1043 2728 1044 2732
rect 1038 2727 1044 2728
rect 1135 2731 1141 2732
rect 1135 2727 1136 2731
rect 1140 2730 1141 2731
rect 1175 2731 1181 2732
rect 1175 2730 1176 2731
rect 1140 2728 1176 2730
rect 1140 2727 1141 2728
rect 471 2726 480 2727
rect 671 2726 680 2727
rect 894 2726 901 2727
rect 1135 2726 1141 2727
rect 1175 2727 1176 2728
rect 1180 2727 1181 2731
rect 1294 2728 1295 2732
rect 1299 2728 1300 2732
rect 1294 2727 1300 2728
rect 1386 2731 1397 2732
rect 1386 2727 1387 2731
rect 1391 2727 1392 2731
rect 1396 2727 1397 2731
rect 1566 2728 1567 2732
rect 1571 2728 1572 2732
rect 1566 2727 1572 2728
rect 1658 2731 1669 2732
rect 1658 2727 1659 2731
rect 1663 2727 1664 2731
rect 1668 2727 1669 2731
rect 1814 2728 1815 2732
rect 1819 2728 1820 2732
rect 1814 2727 1820 2728
rect 1910 2731 1917 2732
rect 1910 2727 1911 2731
rect 1916 2727 1917 2731
rect 1934 2729 1935 2733
rect 1939 2729 1940 2733
rect 1934 2728 1940 2729
rect 1175 2726 1181 2727
rect 1386 2726 1397 2727
rect 1658 2726 1669 2727
rect 1910 2726 1917 2727
rect 4362 2719 4368 2720
rect 346 2717 352 2718
rect 110 2716 116 2717
rect 110 2712 111 2716
rect 115 2712 116 2716
rect 346 2713 347 2717
rect 351 2713 352 2717
rect 346 2712 352 2713
rect 546 2717 552 2718
rect 546 2713 547 2717
rect 551 2713 552 2717
rect 546 2712 552 2713
rect 770 2717 776 2718
rect 770 2713 771 2717
rect 775 2713 776 2717
rect 770 2712 776 2713
rect 1010 2717 1016 2718
rect 1010 2713 1011 2717
rect 1015 2713 1016 2717
rect 1010 2712 1016 2713
rect 1266 2717 1272 2718
rect 1266 2713 1267 2717
rect 1271 2713 1272 2717
rect 1266 2712 1272 2713
rect 1538 2717 1544 2718
rect 1538 2713 1539 2717
rect 1543 2713 1544 2717
rect 1538 2712 1544 2713
rect 1786 2717 1792 2718
rect 1786 2713 1787 2717
rect 1791 2713 1792 2717
rect 1786 2712 1792 2713
rect 1934 2716 1940 2717
rect 1934 2712 1935 2716
rect 1939 2712 1940 2716
rect 4362 2715 4363 2719
rect 4367 2718 4368 2719
rect 4367 2716 5314 2718
rect 4367 2715 4368 2716
rect 4362 2714 4368 2715
rect 110 2711 116 2712
rect 1934 2711 1940 2712
rect 5312 2706 5314 2716
rect 3838 2705 3844 2706
rect 5311 2705 5317 2706
rect 5662 2705 5668 2706
rect 3838 2701 3839 2705
rect 3843 2701 3844 2705
rect 3838 2700 3844 2701
rect 3966 2704 3972 2705
rect 4222 2704 4228 2705
rect 4526 2704 4532 2705
rect 4862 2704 4868 2705
rect 5214 2704 5220 2705
rect 3966 2700 3967 2704
rect 3971 2700 3972 2704
rect 3966 2699 3972 2700
rect 4062 2703 4069 2704
rect 4062 2699 4063 2703
rect 4068 2699 4069 2703
rect 4222 2700 4223 2704
rect 4227 2700 4228 2704
rect 4222 2699 4228 2700
rect 4319 2703 4325 2704
rect 4319 2699 4320 2703
rect 4324 2702 4325 2703
rect 4422 2703 4428 2704
rect 4422 2702 4423 2703
rect 4324 2700 4423 2702
rect 4324 2699 4325 2700
rect 4062 2698 4069 2699
rect 4319 2698 4325 2699
rect 4422 2699 4423 2700
rect 4427 2699 4428 2703
rect 4526 2700 4527 2704
rect 4531 2700 4532 2704
rect 4526 2699 4532 2700
rect 4623 2703 4632 2704
rect 4623 2699 4624 2703
rect 4631 2699 4632 2703
rect 4862 2700 4863 2704
rect 4867 2700 4868 2704
rect 4862 2699 4868 2700
rect 4959 2703 4965 2704
rect 4959 2699 4960 2703
rect 4964 2702 4965 2703
rect 4982 2703 4988 2704
rect 4982 2702 4983 2703
rect 4964 2700 4983 2702
rect 4964 2699 4965 2700
rect 4422 2698 4428 2699
rect 4623 2698 4632 2699
rect 4959 2698 4965 2699
rect 4982 2699 4983 2700
rect 4987 2699 4988 2703
rect 5214 2700 5215 2704
rect 5219 2700 5220 2704
rect 5311 2701 5312 2705
rect 5316 2701 5317 2705
rect 5311 2700 5317 2701
rect 5542 2704 5548 2705
rect 5542 2700 5543 2704
rect 5547 2700 5548 2704
rect 5214 2699 5220 2700
rect 5542 2699 5548 2700
rect 5634 2703 5645 2704
rect 5634 2699 5635 2703
rect 5639 2699 5640 2703
rect 5644 2699 5645 2703
rect 5662 2701 5663 2705
rect 5667 2701 5668 2705
rect 5662 2700 5668 2701
rect 4982 2698 4988 2699
rect 5634 2698 5645 2699
rect 2250 2691 2256 2692
rect 2250 2690 2251 2691
rect 2092 2682 2094 2689
rect 2229 2688 2251 2690
rect 2250 2687 2251 2688
rect 2255 2687 2256 2691
rect 2250 2686 2256 2687
rect 2258 2691 2264 2692
rect 2258 2687 2259 2691
rect 2263 2690 2264 2691
rect 2402 2691 2408 2692
rect 2263 2688 2281 2690
rect 2263 2687 2264 2688
rect 2258 2686 2264 2687
rect 2402 2687 2403 2691
rect 2407 2690 2408 2691
rect 2822 2691 2828 2692
rect 2407 2688 2441 2690
rect 2407 2687 2408 2688
rect 2402 2686 2408 2687
rect 2558 2683 2564 2684
rect 2558 2682 2559 2683
rect 2092 2680 2559 2682
rect 2558 2679 2559 2680
rect 2563 2679 2564 2683
rect 2692 2682 2694 2689
rect 2822 2687 2823 2691
rect 2827 2687 2828 2691
rect 3118 2691 3124 2692
rect 2822 2686 2828 2687
rect 2874 2683 2880 2684
rect 2874 2682 2875 2683
rect 2692 2680 2875 2682
rect 2558 2678 2564 2679
rect 2874 2679 2875 2680
rect 2879 2679 2880 2683
rect 3012 2682 3014 2689
rect 3118 2687 3119 2691
rect 3123 2687 3124 2691
rect 3938 2689 3944 2690
rect 3118 2686 3124 2687
rect 3838 2688 3844 2689
rect 3838 2684 3839 2688
rect 3843 2684 3844 2688
rect 3938 2685 3939 2689
rect 3943 2685 3944 2689
rect 3938 2684 3944 2685
rect 4194 2689 4200 2690
rect 4194 2685 4195 2689
rect 4199 2685 4200 2689
rect 4194 2684 4200 2685
rect 4498 2689 4504 2690
rect 4498 2685 4499 2689
rect 4503 2685 4504 2689
rect 4498 2684 4504 2685
rect 4834 2689 4840 2690
rect 4834 2685 4835 2689
rect 4839 2685 4840 2689
rect 4834 2684 4840 2685
rect 5186 2689 5192 2690
rect 5186 2685 5187 2689
rect 5191 2685 5192 2689
rect 5186 2684 5192 2685
rect 5514 2689 5520 2690
rect 5514 2685 5515 2689
rect 5519 2685 5520 2689
rect 5514 2684 5520 2685
rect 5662 2688 5668 2689
rect 5662 2684 5663 2688
rect 5667 2684 5668 2688
rect 3198 2683 3204 2684
rect 3838 2683 3844 2684
rect 5662 2683 5668 2684
rect 3198 2682 3199 2683
rect 3012 2680 3199 2682
rect 2874 2678 2880 2679
rect 3198 2679 3199 2680
rect 3203 2679 3204 2683
rect 3198 2678 3204 2679
rect 474 2667 480 2668
rect 444 2658 446 2665
rect 474 2663 475 2667
rect 479 2666 480 2667
rect 674 2667 680 2668
rect 479 2664 553 2666
rect 479 2663 480 2664
rect 474 2662 480 2663
rect 674 2663 675 2667
rect 679 2666 680 2667
rect 918 2667 924 2668
rect 679 2664 777 2666
rect 679 2663 680 2664
rect 674 2662 680 2663
rect 918 2663 919 2667
rect 923 2666 924 2667
rect 1175 2667 1181 2668
rect 923 2664 1017 2666
rect 923 2663 924 2664
rect 918 2662 924 2663
rect 1175 2663 1176 2667
rect 1180 2666 1181 2667
rect 2114 2667 2120 2668
rect 2114 2666 2115 2667
rect 1180 2664 1273 2666
rect 1180 2663 1181 2664
rect 1175 2662 1181 2663
rect 506 2659 512 2660
rect 506 2658 507 2659
rect 444 2656 507 2658
rect 506 2655 507 2656
rect 511 2655 512 2659
rect 1636 2658 1638 2665
rect 1885 2664 2115 2666
rect 2114 2663 2115 2664
rect 2119 2663 2120 2667
rect 2114 2662 2120 2663
rect 1910 2659 1916 2660
rect 1910 2658 1911 2659
rect 1636 2656 1911 2658
rect 506 2654 512 2655
rect 1910 2655 1911 2656
rect 1915 2655 1916 2659
rect 1910 2654 1916 2655
rect 3034 2659 3040 2660
rect 3034 2655 3035 2659
rect 3039 2655 3040 2659
rect 3034 2654 3040 2655
rect 2940 2652 3038 2654
rect 2940 2650 2942 2652
rect 2933 2648 2942 2650
rect 1386 2647 1392 2648
rect 1386 2646 1387 2647
rect 1168 2644 1387 2646
rect 1158 2643 1164 2644
rect 1158 2642 1159 2643
rect 984 2640 1159 2642
rect 662 2639 668 2640
rect 662 2638 663 2639
rect 540 2636 663 2638
rect 540 2634 542 2636
rect 662 2635 663 2636
rect 667 2635 668 2639
rect 662 2634 668 2635
rect 854 2635 860 2636
rect 854 2634 855 2635
rect 485 2632 542 2634
rect 797 2632 855 2634
rect 634 2631 640 2632
rect 634 2627 635 2631
rect 639 2627 640 2631
rect 854 2631 855 2632
rect 859 2631 860 2635
rect 984 2634 986 2640
rect 1158 2639 1159 2640
rect 1163 2639 1164 2643
rect 1158 2638 1164 2639
rect 1168 2634 1170 2644
rect 1386 2643 1387 2644
rect 1391 2643 1392 2647
rect 1386 2642 1392 2643
rect 2794 2647 2800 2648
rect 2794 2643 2795 2647
rect 2799 2643 2800 2647
rect 2794 2642 2800 2643
rect 2978 2647 2984 2648
rect 2978 2643 2979 2647
rect 2983 2643 2984 2647
rect 2978 2642 2984 2643
rect 1494 2639 1500 2640
rect 1494 2638 1495 2639
rect 1364 2636 1495 2638
rect 1364 2634 1366 2636
rect 1494 2635 1495 2636
rect 1499 2635 1500 2639
rect 4151 2639 4157 2640
rect 1494 2634 1500 2635
rect 1658 2635 1664 2636
rect 1658 2634 1659 2635
rect 965 2632 986 2634
rect 1133 2632 1170 2634
rect 1301 2632 1366 2634
rect 1637 2632 1659 2634
rect 854 2630 860 2631
rect 1466 2631 1472 2632
rect 634 2626 640 2627
rect 1466 2627 1467 2631
rect 1471 2627 1472 2631
rect 1658 2631 1659 2632
rect 1663 2631 1664 2635
rect 1658 2630 1664 2631
rect 1722 2631 1728 2632
rect 1466 2626 1472 2627
rect 1722 2627 1723 2631
rect 1727 2627 1728 2631
rect 4036 2630 4038 2637
rect 4151 2635 4152 2639
rect 4156 2638 4157 2639
rect 4422 2639 4428 2640
rect 4156 2636 4201 2638
rect 4156 2635 4157 2636
rect 4151 2634 4157 2635
rect 4422 2635 4423 2639
rect 4427 2638 4428 2639
rect 4626 2639 4632 2640
rect 4427 2636 4505 2638
rect 4427 2635 4428 2636
rect 4422 2634 4428 2635
rect 4626 2635 4627 2639
rect 4631 2638 4632 2639
rect 4982 2639 4988 2640
rect 4631 2636 4841 2638
rect 4631 2635 4632 2636
rect 4626 2634 4632 2635
rect 4982 2635 4983 2639
rect 4987 2638 4988 2639
rect 5642 2639 5648 2640
rect 5642 2638 5643 2639
rect 4987 2636 5193 2638
rect 5613 2636 5643 2638
rect 4987 2635 4988 2636
rect 4982 2634 4988 2635
rect 5642 2635 5643 2636
rect 5647 2635 5648 2639
rect 5642 2634 5648 2635
rect 4186 2631 4192 2632
rect 4186 2630 4187 2631
rect 4036 2628 4187 2630
rect 1722 2626 1728 2627
rect 4186 2627 4187 2628
rect 4191 2627 4192 2631
rect 4186 2626 4192 2627
rect 4362 2607 4368 2608
rect 1466 2603 1472 2604
rect 1466 2599 1467 2603
rect 1471 2602 1472 2603
rect 1838 2603 1844 2604
rect 1838 2602 1839 2603
rect 1471 2600 1839 2602
rect 1471 2599 1472 2600
rect 1466 2598 1472 2599
rect 1838 2599 1839 2600
rect 1843 2599 1844 2603
rect 3986 2603 3992 2604
rect 1838 2598 1844 2599
rect 1974 2600 1980 2601
rect 3798 2600 3804 2601
rect 1974 2596 1975 2600
rect 1979 2596 1980 2600
rect 1974 2595 1980 2596
rect 2698 2599 2704 2600
rect 2698 2595 2699 2599
rect 2703 2595 2704 2599
rect 2698 2594 2704 2595
rect 2834 2599 2840 2600
rect 2834 2595 2835 2599
rect 2839 2595 2840 2599
rect 2834 2594 2840 2595
rect 2970 2599 2976 2600
rect 2970 2595 2971 2599
rect 2975 2595 2976 2599
rect 3798 2596 3799 2600
rect 3803 2596 3804 2600
rect 3986 2599 3987 2603
rect 3991 2599 3992 2603
rect 3986 2598 3992 2599
rect 4074 2603 4080 2604
rect 4074 2599 4075 2603
rect 4079 2599 4080 2603
rect 4362 2603 4363 2607
rect 4367 2603 4368 2607
rect 5442 2607 5448 2608
rect 5442 2606 5443 2607
rect 5365 2604 5443 2606
rect 4362 2602 4368 2603
rect 4498 2603 4504 2604
rect 4074 2598 4080 2599
rect 4498 2599 4499 2603
rect 4503 2599 4504 2603
rect 4498 2598 4504 2599
rect 4738 2603 4744 2604
rect 4738 2599 4739 2603
rect 4743 2599 4744 2603
rect 4738 2598 4744 2599
rect 5002 2603 5008 2604
rect 5002 2599 5003 2603
rect 5007 2599 5008 2603
rect 5442 2603 5443 2604
rect 5447 2603 5448 2607
rect 5634 2607 5640 2608
rect 5634 2606 5635 2607
rect 5613 2604 5635 2606
rect 5442 2602 5448 2603
rect 5634 2603 5635 2604
rect 5639 2603 5640 2607
rect 5634 2602 5640 2603
rect 5002 2598 5008 2599
rect 3798 2595 3804 2596
rect 2970 2594 2976 2595
rect 110 2584 116 2585
rect 1934 2584 1940 2585
rect 2726 2584 2732 2585
rect 2862 2584 2868 2585
rect 2998 2584 3004 2585
rect 110 2580 111 2584
rect 115 2580 116 2584
rect 110 2579 116 2580
rect 386 2583 392 2584
rect 386 2579 387 2583
rect 391 2579 392 2583
rect 386 2578 392 2579
rect 538 2583 544 2584
rect 538 2579 539 2583
rect 543 2579 544 2583
rect 538 2578 544 2579
rect 698 2583 704 2584
rect 698 2579 699 2583
rect 703 2579 704 2583
rect 698 2578 704 2579
rect 866 2583 872 2584
rect 866 2579 867 2583
rect 871 2579 872 2583
rect 866 2578 872 2579
rect 1034 2583 1040 2584
rect 1034 2579 1035 2583
rect 1039 2579 1040 2583
rect 1034 2578 1040 2579
rect 1202 2583 1208 2584
rect 1202 2579 1203 2583
rect 1207 2579 1208 2583
rect 1202 2578 1208 2579
rect 1370 2583 1376 2584
rect 1370 2579 1371 2583
rect 1375 2579 1376 2583
rect 1370 2578 1376 2579
rect 1538 2583 1544 2584
rect 1538 2579 1539 2583
rect 1543 2579 1544 2583
rect 1538 2578 1544 2579
rect 1714 2583 1720 2584
rect 1714 2579 1715 2583
rect 1719 2579 1720 2583
rect 1934 2580 1935 2584
rect 1939 2580 1940 2584
rect 1934 2579 1940 2580
rect 1974 2583 1980 2584
rect 1974 2579 1975 2583
rect 1979 2579 1980 2583
rect 2726 2580 2727 2584
rect 2731 2580 2732 2584
rect 2726 2579 2732 2580
rect 2822 2583 2829 2584
rect 2822 2579 2823 2583
rect 2828 2579 2829 2583
rect 2862 2580 2863 2584
rect 2867 2580 2868 2584
rect 2862 2579 2868 2580
rect 2959 2583 2965 2584
rect 2959 2579 2960 2583
rect 2964 2582 2965 2583
rect 2978 2583 2984 2584
rect 2978 2582 2979 2583
rect 2964 2580 2979 2582
rect 2964 2579 2965 2580
rect 1714 2578 1720 2579
rect 1974 2578 1980 2579
rect 2822 2578 2829 2579
rect 2959 2578 2965 2579
rect 2978 2579 2979 2580
rect 2983 2579 2984 2583
rect 2998 2580 2999 2584
rect 3003 2580 3004 2584
rect 2998 2579 3004 2580
rect 3094 2583 3101 2584
rect 3094 2579 3095 2583
rect 3100 2579 3101 2583
rect 2978 2578 2984 2579
rect 3094 2578 3101 2579
rect 3798 2583 3804 2584
rect 3798 2579 3799 2583
rect 3803 2579 3804 2583
rect 3798 2578 3804 2579
rect 854 2575 860 2576
rect 854 2571 855 2575
rect 859 2574 860 2575
rect 859 2572 994 2574
rect 859 2571 860 2572
rect 854 2570 860 2571
rect 992 2570 994 2572
rect 991 2569 997 2570
rect 414 2568 420 2569
rect 566 2568 572 2569
rect 726 2568 732 2569
rect 894 2568 900 2569
rect 110 2567 116 2568
rect 110 2563 111 2567
rect 115 2563 116 2567
rect 414 2564 415 2568
rect 419 2564 420 2568
rect 414 2563 420 2564
rect 506 2567 517 2568
rect 506 2563 507 2567
rect 511 2563 512 2567
rect 516 2563 517 2567
rect 566 2564 567 2568
rect 571 2564 572 2568
rect 566 2563 572 2564
rect 662 2567 669 2568
rect 662 2563 663 2567
rect 668 2563 669 2567
rect 726 2564 727 2568
rect 731 2564 732 2568
rect 726 2563 732 2564
rect 822 2567 829 2568
rect 822 2563 823 2567
rect 828 2563 829 2567
rect 894 2564 895 2568
rect 899 2564 900 2568
rect 991 2565 992 2569
rect 996 2565 997 2569
rect 991 2564 997 2565
rect 1062 2568 1068 2569
rect 1230 2568 1236 2569
rect 1398 2568 1404 2569
rect 1566 2568 1572 2569
rect 1742 2568 1748 2569
rect 1062 2564 1063 2568
rect 1067 2564 1068 2568
rect 894 2563 900 2564
rect 1062 2563 1068 2564
rect 1158 2567 1165 2568
rect 1158 2563 1159 2567
rect 1164 2563 1165 2567
rect 1230 2564 1231 2568
rect 1235 2564 1236 2568
rect 1230 2563 1236 2564
rect 1326 2567 1333 2568
rect 1326 2563 1327 2567
rect 1332 2563 1333 2567
rect 1398 2564 1399 2568
rect 1403 2564 1404 2568
rect 1398 2563 1404 2564
rect 1494 2567 1501 2568
rect 1494 2563 1495 2567
rect 1500 2563 1501 2567
rect 1566 2564 1567 2568
rect 1571 2564 1572 2568
rect 1566 2563 1572 2564
rect 1663 2567 1669 2568
rect 1663 2563 1664 2567
rect 1668 2566 1669 2567
rect 1722 2567 1728 2568
rect 1722 2566 1723 2567
rect 1668 2564 1723 2566
rect 1668 2563 1669 2564
rect 110 2562 116 2563
rect 506 2562 517 2563
rect 662 2562 669 2563
rect 822 2562 829 2563
rect 1158 2562 1165 2563
rect 1326 2562 1333 2563
rect 1494 2562 1501 2563
rect 1663 2562 1669 2563
rect 1722 2563 1723 2564
rect 1727 2563 1728 2567
rect 1742 2564 1743 2568
rect 1747 2564 1748 2568
rect 1742 2563 1748 2564
rect 1838 2567 1845 2568
rect 1838 2563 1839 2567
rect 1844 2563 1845 2567
rect 1722 2562 1728 2563
rect 1838 2562 1845 2563
rect 1934 2567 1940 2568
rect 1934 2563 1935 2567
rect 1939 2563 1940 2567
rect 1934 2562 1940 2563
rect 3838 2556 3844 2557
rect 5662 2556 5668 2557
rect 3838 2552 3839 2556
rect 3843 2552 3844 2556
rect 3838 2551 3844 2552
rect 3890 2555 3896 2556
rect 3890 2551 3891 2555
rect 3895 2551 3896 2555
rect 3890 2550 3896 2551
rect 4066 2555 4072 2556
rect 4066 2551 4067 2555
rect 4071 2551 4072 2555
rect 4066 2550 4072 2551
rect 4266 2555 4272 2556
rect 4266 2551 4267 2555
rect 4271 2551 4272 2555
rect 4266 2550 4272 2551
rect 4490 2555 4496 2556
rect 4490 2551 4491 2555
rect 4495 2551 4496 2555
rect 4490 2550 4496 2551
rect 4730 2555 4736 2556
rect 4730 2551 4731 2555
rect 4735 2551 4736 2555
rect 4730 2550 4736 2551
rect 4994 2555 5000 2556
rect 4994 2551 4995 2555
rect 4999 2551 5000 2555
rect 4994 2550 5000 2551
rect 5266 2555 5272 2556
rect 5266 2551 5267 2555
rect 5271 2551 5272 2555
rect 5266 2550 5272 2551
rect 5514 2555 5520 2556
rect 5514 2551 5515 2555
rect 5519 2551 5520 2555
rect 5662 2552 5663 2556
rect 5667 2552 5668 2556
rect 5662 2551 5668 2552
rect 5514 2550 5520 2551
rect 3918 2540 3924 2541
rect 4094 2540 4100 2541
rect 4294 2540 4300 2541
rect 4518 2540 4524 2541
rect 4758 2540 4764 2541
rect 5022 2540 5028 2541
rect 5294 2540 5300 2541
rect 5542 2540 5548 2541
rect 2794 2539 2800 2540
rect 2794 2535 2795 2539
rect 2799 2538 2800 2539
rect 3838 2539 3844 2540
rect 2799 2536 2858 2538
rect 2799 2535 2800 2536
rect 2794 2534 2800 2535
rect 1974 2525 1980 2526
rect 1974 2521 1975 2525
rect 1979 2521 1980 2525
rect 1974 2520 1980 2521
rect 2606 2524 2612 2525
rect 2758 2524 2764 2525
rect 2856 2524 2858 2536
rect 3838 2535 3839 2539
rect 3843 2535 3844 2539
rect 3918 2536 3919 2540
rect 3923 2536 3924 2540
rect 3918 2535 3924 2536
rect 4015 2539 4021 2540
rect 4015 2535 4016 2539
rect 4020 2538 4021 2539
rect 4074 2539 4080 2540
rect 4074 2538 4075 2539
rect 4020 2536 4075 2538
rect 4020 2535 4021 2536
rect 3838 2534 3844 2535
rect 4015 2534 4021 2535
rect 4074 2535 4075 2536
rect 4079 2535 4080 2539
rect 4094 2536 4095 2540
rect 4099 2536 4100 2540
rect 4094 2535 4100 2536
rect 4186 2539 4197 2540
rect 4186 2535 4187 2539
rect 4191 2535 4192 2539
rect 4196 2535 4197 2539
rect 4294 2536 4295 2540
rect 4299 2536 4300 2540
rect 4294 2535 4300 2536
rect 4391 2539 4397 2540
rect 4391 2535 4392 2539
rect 4396 2538 4397 2539
rect 4498 2539 4504 2540
rect 4498 2538 4499 2539
rect 4396 2536 4499 2538
rect 4396 2535 4397 2536
rect 4074 2534 4080 2535
rect 4186 2534 4197 2535
rect 4391 2534 4397 2535
rect 4498 2535 4499 2536
rect 4503 2535 4504 2539
rect 4518 2536 4519 2540
rect 4523 2536 4524 2540
rect 4518 2535 4524 2536
rect 4615 2539 4621 2540
rect 4615 2535 4616 2539
rect 4620 2538 4621 2539
rect 4738 2539 4744 2540
rect 4738 2538 4739 2539
rect 4620 2536 4739 2538
rect 4620 2535 4621 2536
rect 4498 2534 4504 2535
rect 4615 2534 4621 2535
rect 4738 2535 4739 2536
rect 4743 2535 4744 2539
rect 4758 2536 4759 2540
rect 4763 2536 4764 2540
rect 4758 2535 4764 2536
rect 4855 2539 4861 2540
rect 4855 2535 4856 2539
rect 4860 2538 4861 2539
rect 5002 2539 5008 2540
rect 5002 2538 5003 2539
rect 4860 2536 5003 2538
rect 4860 2535 4861 2536
rect 4738 2534 4744 2535
rect 4855 2534 4861 2535
rect 5002 2535 5003 2536
rect 5007 2535 5008 2539
rect 5022 2536 5023 2540
rect 5027 2536 5028 2540
rect 5022 2535 5028 2536
rect 5114 2539 5125 2540
rect 5114 2535 5115 2539
rect 5119 2535 5120 2539
rect 5124 2535 5125 2539
rect 5294 2536 5295 2540
rect 5299 2536 5300 2540
rect 5294 2535 5300 2536
rect 5390 2539 5397 2540
rect 5390 2535 5391 2539
rect 5396 2535 5397 2539
rect 5542 2536 5543 2540
rect 5547 2536 5548 2540
rect 5542 2535 5548 2536
rect 5634 2539 5645 2540
rect 5634 2535 5635 2539
rect 5639 2535 5640 2539
rect 5644 2535 5645 2539
rect 5002 2534 5008 2535
rect 5114 2534 5125 2535
rect 5390 2534 5397 2535
rect 5634 2534 5645 2535
rect 5662 2539 5668 2540
rect 5662 2535 5663 2539
rect 5667 2535 5668 2539
rect 5662 2534 5668 2535
rect 3798 2525 3804 2526
rect 2910 2524 2916 2525
rect 3062 2524 3068 2525
rect 3222 2524 3228 2525
rect 2606 2520 2607 2524
rect 2611 2520 2612 2524
rect 2606 2519 2612 2520
rect 2702 2523 2709 2524
rect 2702 2519 2703 2523
rect 2708 2519 2709 2523
rect 2758 2520 2759 2524
rect 2763 2520 2764 2524
rect 2758 2519 2764 2520
rect 2855 2523 2861 2524
rect 2855 2519 2856 2523
rect 2860 2519 2861 2523
rect 2910 2520 2911 2524
rect 2915 2520 2916 2524
rect 2910 2519 2916 2520
rect 3002 2523 3013 2524
rect 3002 2519 3003 2523
rect 3007 2519 3008 2523
rect 3012 2519 3013 2523
rect 3062 2520 3063 2524
rect 3067 2520 3068 2524
rect 3062 2519 3068 2520
rect 3159 2523 3168 2524
rect 3159 2519 3160 2523
rect 3167 2519 3168 2523
rect 3222 2520 3223 2524
rect 3227 2520 3228 2524
rect 3222 2519 3228 2520
rect 3318 2523 3325 2524
rect 3318 2519 3319 2523
rect 3324 2519 3325 2523
rect 3798 2521 3799 2525
rect 3803 2521 3804 2525
rect 3798 2520 3804 2521
rect 2702 2518 2709 2519
rect 2855 2518 2861 2519
rect 3002 2518 3013 2519
rect 3159 2518 3168 2519
rect 3318 2518 3325 2519
rect 110 2509 116 2510
rect 1934 2509 1940 2510
rect 2578 2509 2584 2510
rect 110 2505 111 2509
rect 115 2505 116 2509
rect 110 2504 116 2505
rect 326 2508 332 2509
rect 534 2508 540 2509
rect 734 2508 740 2509
rect 918 2508 924 2509
rect 1094 2508 1100 2509
rect 1270 2508 1276 2509
rect 1438 2508 1444 2509
rect 1606 2508 1612 2509
rect 1774 2508 1780 2509
rect 326 2504 327 2508
rect 331 2504 332 2508
rect 326 2503 332 2504
rect 423 2507 432 2508
rect 423 2503 424 2507
rect 431 2503 432 2507
rect 534 2504 535 2508
rect 539 2504 540 2508
rect 534 2503 540 2504
rect 631 2507 640 2508
rect 631 2503 632 2507
rect 639 2503 640 2507
rect 734 2504 735 2508
rect 739 2504 740 2508
rect 734 2503 740 2504
rect 831 2507 837 2508
rect 831 2503 832 2507
rect 836 2506 837 2507
rect 855 2507 861 2508
rect 855 2506 856 2507
rect 836 2504 856 2506
rect 836 2503 837 2504
rect 423 2502 432 2503
rect 631 2502 640 2503
rect 831 2502 837 2503
rect 855 2503 856 2504
rect 860 2503 861 2507
rect 918 2504 919 2508
rect 923 2504 924 2508
rect 918 2503 924 2504
rect 1015 2507 1021 2508
rect 1015 2503 1016 2507
rect 1020 2506 1021 2507
rect 1030 2507 1036 2508
rect 1030 2506 1031 2507
rect 1020 2504 1031 2506
rect 1020 2503 1021 2504
rect 855 2502 861 2503
rect 1015 2502 1021 2503
rect 1030 2503 1031 2504
rect 1035 2503 1036 2507
rect 1094 2504 1095 2508
rect 1099 2504 1100 2508
rect 1094 2503 1100 2504
rect 1186 2507 1197 2508
rect 1186 2503 1187 2507
rect 1191 2503 1192 2507
rect 1196 2503 1197 2507
rect 1270 2504 1271 2508
rect 1275 2504 1276 2508
rect 1270 2503 1276 2504
rect 1367 2507 1376 2508
rect 1367 2503 1368 2507
rect 1375 2503 1376 2507
rect 1438 2504 1439 2508
rect 1443 2504 1444 2508
rect 1438 2503 1444 2504
rect 1535 2507 1544 2508
rect 1535 2503 1536 2507
rect 1543 2503 1544 2507
rect 1606 2504 1607 2508
rect 1611 2504 1612 2508
rect 1606 2503 1612 2504
rect 1703 2507 1712 2508
rect 1703 2503 1704 2507
rect 1711 2503 1712 2507
rect 1774 2504 1775 2508
rect 1779 2504 1780 2508
rect 1774 2503 1780 2504
rect 1866 2507 1877 2508
rect 1866 2503 1867 2507
rect 1871 2503 1872 2507
rect 1876 2503 1877 2507
rect 1934 2505 1935 2509
rect 1939 2505 1940 2509
rect 1934 2504 1940 2505
rect 1974 2508 1980 2509
rect 1974 2504 1975 2508
rect 1979 2504 1980 2508
rect 2578 2505 2579 2509
rect 2583 2505 2584 2509
rect 2578 2504 2584 2505
rect 2730 2509 2736 2510
rect 2730 2505 2731 2509
rect 2735 2505 2736 2509
rect 2730 2504 2736 2505
rect 2882 2509 2888 2510
rect 2882 2505 2883 2509
rect 2887 2505 2888 2509
rect 2882 2504 2888 2505
rect 3034 2509 3040 2510
rect 3034 2505 3035 2509
rect 3039 2505 3040 2509
rect 3034 2504 3040 2505
rect 3194 2509 3200 2510
rect 3194 2505 3195 2509
rect 3199 2505 3200 2509
rect 3194 2504 3200 2505
rect 3798 2508 3804 2509
rect 3798 2504 3799 2508
rect 3803 2504 3804 2508
rect 1974 2503 1980 2504
rect 3798 2503 3804 2504
rect 1030 2502 1036 2503
rect 1186 2502 1197 2503
rect 1367 2502 1376 2503
rect 1535 2502 1544 2503
rect 1703 2502 1712 2503
rect 1866 2502 1877 2503
rect 298 2493 304 2494
rect 110 2492 116 2493
rect 110 2488 111 2492
rect 115 2488 116 2492
rect 298 2489 299 2493
rect 303 2489 304 2493
rect 298 2488 304 2489
rect 506 2493 512 2494
rect 506 2489 507 2493
rect 511 2489 512 2493
rect 506 2488 512 2489
rect 706 2493 712 2494
rect 706 2489 707 2493
rect 711 2489 712 2493
rect 706 2488 712 2489
rect 890 2493 896 2494
rect 890 2489 891 2493
rect 895 2489 896 2493
rect 890 2488 896 2489
rect 1066 2493 1072 2494
rect 1066 2489 1067 2493
rect 1071 2489 1072 2493
rect 1066 2488 1072 2489
rect 1242 2493 1248 2494
rect 1242 2489 1243 2493
rect 1247 2489 1248 2493
rect 1242 2488 1248 2489
rect 1410 2493 1416 2494
rect 1410 2489 1411 2493
rect 1415 2489 1416 2493
rect 1410 2488 1416 2489
rect 1578 2493 1584 2494
rect 1578 2489 1579 2493
rect 1583 2489 1584 2493
rect 1578 2488 1584 2489
rect 1746 2493 1752 2494
rect 1746 2489 1747 2493
rect 1751 2489 1752 2493
rect 1746 2488 1752 2489
rect 1934 2492 1940 2493
rect 1934 2488 1935 2492
rect 1939 2488 1940 2492
rect 110 2487 116 2488
rect 1934 2487 1940 2488
rect 4439 2491 4445 2492
rect 4439 2487 4440 2491
rect 4444 2490 4445 2491
rect 4444 2488 5186 2490
rect 4444 2487 4445 2488
rect 4439 2486 4445 2487
rect 3838 2477 3844 2478
rect 3838 2473 3839 2477
rect 3843 2473 3844 2477
rect 3838 2472 3844 2473
rect 3886 2476 3892 2477
rect 4086 2476 4092 2477
rect 4318 2476 4324 2477
rect 4566 2476 4572 2477
rect 4822 2476 4828 2477
rect 5086 2476 5092 2477
rect 5184 2476 5186 2488
rect 5662 2477 5668 2478
rect 5350 2476 5356 2477
rect 3886 2472 3887 2476
rect 3891 2472 3892 2476
rect 3886 2471 3892 2472
rect 3983 2475 3992 2476
rect 3983 2471 3984 2475
rect 3991 2471 3992 2475
rect 4086 2472 4087 2476
rect 4091 2472 4092 2476
rect 4086 2471 4092 2472
rect 4182 2475 4189 2476
rect 4182 2471 4183 2475
rect 4188 2471 4189 2475
rect 4318 2472 4319 2476
rect 4323 2472 4324 2476
rect 4318 2471 4324 2472
rect 4415 2475 4421 2476
rect 4415 2471 4416 2475
rect 4420 2474 4421 2475
rect 4438 2475 4444 2476
rect 4438 2474 4439 2475
rect 4420 2472 4439 2474
rect 4420 2471 4421 2472
rect 3983 2470 3992 2471
rect 4182 2470 4189 2471
rect 4415 2470 4421 2471
rect 4438 2471 4439 2472
rect 4443 2471 4444 2475
rect 4566 2472 4567 2476
rect 4571 2472 4572 2476
rect 4566 2471 4572 2472
rect 4663 2475 4669 2476
rect 4663 2471 4664 2475
rect 4668 2474 4669 2475
rect 4710 2475 4716 2476
rect 4710 2474 4711 2475
rect 4668 2472 4711 2474
rect 4668 2471 4669 2472
rect 4438 2470 4444 2471
rect 4663 2470 4669 2471
rect 4710 2471 4711 2472
rect 4715 2471 4716 2475
rect 4822 2472 4823 2476
rect 4827 2472 4828 2476
rect 4822 2471 4828 2472
rect 4919 2475 4925 2476
rect 4919 2471 4920 2475
rect 4924 2474 4925 2475
rect 4974 2475 4980 2476
rect 4974 2474 4975 2475
rect 4924 2472 4975 2474
rect 4924 2471 4925 2472
rect 4710 2470 4716 2471
rect 4919 2470 4925 2471
rect 4974 2471 4975 2472
rect 4979 2471 4980 2475
rect 5086 2472 5087 2476
rect 5091 2472 5092 2476
rect 5086 2471 5092 2472
rect 5183 2475 5189 2476
rect 5183 2471 5184 2475
rect 5188 2471 5189 2475
rect 5350 2472 5351 2476
rect 5355 2472 5356 2476
rect 5350 2471 5356 2472
rect 5442 2475 5453 2476
rect 5442 2471 5443 2475
rect 5447 2471 5448 2475
rect 5452 2471 5453 2475
rect 5662 2473 5663 2477
rect 5667 2473 5668 2477
rect 5662 2472 5668 2473
rect 4974 2470 4980 2471
rect 5183 2470 5189 2471
rect 5442 2470 5453 2471
rect 3858 2461 3864 2462
rect 3838 2460 3844 2461
rect 2690 2459 2696 2460
rect 2690 2458 2691 2459
rect 2677 2456 2691 2458
rect 2690 2455 2691 2456
rect 2695 2455 2696 2459
rect 2690 2454 2696 2455
rect 2702 2459 2708 2460
rect 2702 2455 2703 2459
rect 2707 2458 2708 2459
rect 3094 2459 3100 2460
rect 2707 2456 2737 2458
rect 2707 2455 2708 2456
rect 2702 2454 2708 2455
rect 2980 2450 2982 2457
rect 3094 2455 3095 2459
rect 3099 2455 3100 2459
rect 3094 2454 3100 2455
rect 3162 2459 3168 2460
rect 3162 2455 3163 2459
rect 3167 2458 3168 2459
rect 3167 2456 3201 2458
rect 3838 2456 3839 2460
rect 3843 2456 3844 2460
rect 3858 2457 3859 2461
rect 3863 2457 3864 2461
rect 3858 2456 3864 2457
rect 4058 2461 4064 2462
rect 4058 2457 4059 2461
rect 4063 2457 4064 2461
rect 4058 2456 4064 2457
rect 4290 2461 4296 2462
rect 4290 2457 4291 2461
rect 4295 2457 4296 2461
rect 4290 2456 4296 2457
rect 4538 2461 4544 2462
rect 4538 2457 4539 2461
rect 4543 2457 4544 2461
rect 4538 2456 4544 2457
rect 4794 2461 4800 2462
rect 4794 2457 4795 2461
rect 4799 2457 4800 2461
rect 4794 2456 4800 2457
rect 5058 2461 5064 2462
rect 5058 2457 5059 2461
rect 5063 2457 5064 2461
rect 5058 2456 5064 2457
rect 5322 2461 5328 2462
rect 5322 2457 5323 2461
rect 5327 2457 5328 2461
rect 5322 2456 5328 2457
rect 5662 2460 5668 2461
rect 5662 2456 5663 2460
rect 5667 2456 5668 2460
rect 3167 2455 3168 2456
rect 3838 2455 3844 2456
rect 5662 2455 5668 2456
rect 3162 2454 3168 2455
rect 3318 2451 3324 2452
rect 3318 2450 3319 2451
rect 2980 2448 3319 2450
rect 3318 2447 3319 2448
rect 3323 2447 3324 2451
rect 3318 2446 3324 2447
rect 279 2443 285 2444
rect 279 2439 280 2443
rect 284 2442 285 2443
rect 426 2443 432 2444
rect 284 2440 305 2442
rect 284 2439 285 2440
rect 279 2438 285 2439
rect 426 2439 427 2443
rect 431 2442 432 2443
rect 822 2443 828 2444
rect 822 2442 823 2443
rect 431 2440 513 2442
rect 805 2440 823 2442
rect 431 2439 432 2440
rect 426 2438 432 2439
rect 822 2439 823 2440
rect 827 2439 828 2443
rect 822 2438 828 2439
rect 855 2443 861 2444
rect 855 2439 856 2443
rect 860 2442 861 2443
rect 1030 2443 1036 2444
rect 860 2440 897 2442
rect 860 2439 861 2440
rect 855 2438 861 2439
rect 1030 2439 1031 2443
rect 1035 2442 1036 2443
rect 1326 2443 1332 2444
rect 1035 2440 1073 2442
rect 1035 2439 1036 2440
rect 1030 2438 1036 2439
rect 1326 2439 1327 2443
rect 1331 2439 1332 2443
rect 1326 2438 1332 2439
rect 1370 2443 1376 2444
rect 1370 2439 1371 2443
rect 1375 2442 1376 2443
rect 1538 2443 1544 2444
rect 1375 2440 1417 2442
rect 1375 2439 1376 2440
rect 1370 2438 1376 2439
rect 1538 2439 1539 2443
rect 1543 2442 1544 2443
rect 1706 2443 1712 2444
rect 1543 2440 1585 2442
rect 1543 2439 1544 2440
rect 1538 2438 1544 2439
rect 1706 2439 1707 2443
rect 1711 2442 1712 2443
rect 1711 2440 1753 2442
rect 1711 2439 1712 2440
rect 1706 2438 1712 2439
rect 1866 2415 1872 2416
rect 1866 2414 1867 2415
rect 1704 2412 1867 2414
rect 518 2407 524 2408
rect 518 2406 519 2407
rect 501 2404 519 2406
rect 226 2403 232 2404
rect 226 2399 227 2403
rect 231 2399 232 2403
rect 518 2403 519 2404
rect 523 2403 524 2407
rect 1186 2407 1192 2408
rect 1186 2406 1187 2407
rect 1069 2404 1187 2406
rect 518 2402 524 2403
rect 698 2403 704 2404
rect 226 2398 232 2399
rect 698 2399 699 2403
rect 703 2399 704 2403
rect 1186 2403 1187 2404
rect 1191 2403 1192 2407
rect 1704 2406 1706 2412
rect 1866 2411 1867 2412
rect 1871 2411 1872 2415
rect 2702 2415 2708 2416
rect 2702 2414 2703 2415
rect 2492 2412 2703 2414
rect 1866 2410 1872 2411
rect 1914 2411 1920 2412
rect 1914 2407 1915 2411
rect 1919 2410 1920 2411
rect 2492 2410 2494 2412
rect 2702 2411 2703 2412
rect 2707 2411 2708 2415
rect 2702 2410 2708 2411
rect 3002 2411 3008 2412
rect 3002 2410 3003 2411
rect 1919 2408 2001 2410
rect 2373 2408 2494 2410
rect 2957 2408 3003 2410
rect 1919 2407 1920 2408
rect 1914 2406 1920 2407
rect 2578 2407 2584 2408
rect 1629 2404 1706 2406
rect 1186 2402 1192 2403
rect 1258 2403 1264 2404
rect 698 2398 704 2399
rect 1258 2399 1259 2403
rect 1263 2399 1264 2403
rect 1258 2398 1264 2399
rect 1794 2403 1800 2404
rect 1794 2399 1795 2403
rect 1799 2399 1800 2403
rect 2578 2403 2579 2407
rect 2583 2403 2584 2407
rect 3002 2407 3003 2408
rect 3007 2407 3008 2411
rect 4210 2411 4216 2412
rect 4210 2410 4211 2411
rect 3002 2406 3008 2407
rect 3154 2407 3160 2408
rect 2578 2402 2584 2403
rect 3154 2403 3155 2407
rect 3159 2403 3160 2407
rect 3154 2402 3160 2403
rect 3442 2407 3448 2408
rect 3442 2403 3443 2407
rect 3447 2403 3448 2407
rect 3442 2402 3448 2403
rect 3956 2402 3958 2409
rect 4157 2408 4211 2410
rect 4210 2407 4211 2408
rect 4215 2407 4216 2411
rect 4210 2406 4216 2407
rect 4386 2411 4392 2412
rect 4386 2407 4387 2411
rect 4391 2407 4392 2411
rect 4386 2406 4392 2407
rect 4438 2411 4444 2412
rect 4438 2407 4439 2411
rect 4443 2410 4444 2411
rect 4710 2411 4716 2412
rect 4443 2408 4545 2410
rect 4443 2407 4444 2408
rect 4438 2406 4444 2407
rect 4710 2407 4711 2411
rect 4715 2410 4716 2411
rect 4974 2411 4980 2412
rect 4715 2408 4801 2410
rect 4715 2407 4716 2408
rect 4710 2406 4716 2407
rect 4974 2407 4975 2411
rect 4979 2410 4980 2411
rect 5406 2411 5412 2412
rect 4979 2408 5065 2410
rect 4979 2407 4980 2408
rect 4974 2406 4980 2407
rect 5406 2407 5407 2411
rect 5411 2407 5412 2411
rect 5406 2406 5412 2407
rect 4182 2403 4188 2404
rect 4182 2402 4183 2403
rect 3956 2400 4183 2402
rect 1794 2398 1800 2399
rect 4182 2399 4183 2400
rect 4187 2399 4188 2403
rect 4182 2398 4188 2399
rect 3790 2379 3796 2380
rect 226 2375 232 2376
rect 226 2371 227 2375
rect 231 2374 232 2375
rect 814 2375 820 2376
rect 814 2374 815 2375
rect 231 2372 815 2374
rect 231 2371 232 2372
rect 226 2370 232 2371
rect 814 2371 815 2372
rect 819 2371 820 2375
rect 3790 2375 3791 2379
rect 3795 2378 3796 2379
rect 4439 2379 4445 2380
rect 4439 2378 4440 2379
rect 3795 2376 3865 2378
rect 4437 2376 4440 2378
rect 3795 2375 3796 2376
rect 3790 2374 3796 2375
rect 4098 2375 4104 2376
rect 814 2370 820 2371
rect 4098 2371 4099 2375
rect 4103 2371 4104 2375
rect 4439 2375 4440 2376
rect 4444 2375 4445 2379
rect 5498 2379 5504 2380
rect 5498 2378 5499 2379
rect 5381 2376 5499 2378
rect 4439 2374 4445 2375
rect 4586 2375 4592 2376
rect 4098 2370 4104 2371
rect 4586 2371 4587 2375
rect 4591 2371 4592 2375
rect 4586 2370 4592 2371
rect 4818 2375 4824 2376
rect 4818 2371 4819 2375
rect 4823 2371 4824 2375
rect 4818 2370 4824 2371
rect 5050 2375 5056 2376
rect 5050 2371 5051 2375
rect 5055 2371 5056 2375
rect 5498 2375 5499 2376
rect 5503 2375 5504 2379
rect 5634 2379 5640 2380
rect 5634 2378 5635 2379
rect 5613 2376 5635 2378
rect 5498 2374 5504 2375
rect 5634 2375 5635 2376
rect 5639 2375 5640 2379
rect 5634 2374 5640 2375
rect 5050 2370 5056 2371
rect 1974 2360 1980 2361
rect 3798 2360 3804 2361
rect 110 2356 116 2357
rect 1934 2356 1940 2357
rect 110 2352 111 2356
rect 115 2352 116 2356
rect 110 2351 116 2352
rect 130 2355 136 2356
rect 130 2351 131 2355
rect 135 2351 136 2355
rect 130 2350 136 2351
rect 402 2355 408 2356
rect 402 2351 403 2355
rect 407 2351 408 2355
rect 402 2350 408 2351
rect 690 2355 696 2356
rect 690 2351 691 2355
rect 695 2351 696 2355
rect 690 2350 696 2351
rect 970 2355 976 2356
rect 970 2351 971 2355
rect 975 2351 976 2355
rect 970 2350 976 2351
rect 1250 2355 1256 2356
rect 1250 2351 1251 2355
rect 1255 2351 1256 2355
rect 1250 2350 1256 2351
rect 1530 2355 1536 2356
rect 1530 2351 1531 2355
rect 1535 2351 1536 2355
rect 1530 2350 1536 2351
rect 1786 2355 1792 2356
rect 1786 2351 1787 2355
rect 1791 2351 1792 2355
rect 1934 2352 1935 2356
rect 1939 2352 1940 2356
rect 1974 2356 1975 2360
rect 1979 2356 1980 2360
rect 1974 2355 1980 2356
rect 1994 2359 2000 2360
rect 1994 2355 1995 2359
rect 1999 2355 2000 2359
rect 1994 2354 2000 2355
rect 2274 2359 2280 2360
rect 2274 2355 2275 2359
rect 2279 2355 2280 2359
rect 2274 2354 2280 2355
rect 2570 2359 2576 2360
rect 2570 2355 2571 2359
rect 2575 2355 2576 2359
rect 2570 2354 2576 2355
rect 2858 2359 2864 2360
rect 2858 2355 2859 2359
rect 2863 2355 2864 2359
rect 2858 2354 2864 2355
rect 3146 2359 3152 2360
rect 3146 2355 3147 2359
rect 3151 2355 3152 2359
rect 3146 2354 3152 2355
rect 3434 2359 3440 2360
rect 3434 2355 3435 2359
rect 3439 2355 3440 2359
rect 3798 2356 3799 2360
rect 3803 2356 3804 2360
rect 3798 2355 3804 2356
rect 3434 2354 3440 2355
rect 1934 2351 1940 2352
rect 1786 2350 1792 2351
rect 2022 2344 2028 2345
rect 2302 2344 2308 2345
rect 2598 2344 2604 2345
rect 2886 2344 2892 2345
rect 3174 2344 3180 2345
rect 3462 2344 3468 2345
rect 1974 2343 1980 2344
rect 158 2340 164 2341
rect 430 2340 436 2341
rect 718 2340 724 2341
rect 998 2340 1004 2341
rect 1278 2340 1284 2341
rect 1558 2340 1564 2341
rect 1814 2340 1820 2341
rect 110 2339 116 2340
rect 110 2335 111 2339
rect 115 2335 116 2339
rect 158 2336 159 2340
rect 163 2336 164 2340
rect 158 2335 164 2336
rect 255 2339 261 2340
rect 255 2335 256 2339
rect 260 2338 261 2339
rect 279 2339 285 2340
rect 279 2338 280 2339
rect 260 2336 280 2338
rect 260 2335 261 2336
rect 110 2334 116 2335
rect 255 2334 261 2335
rect 279 2335 280 2336
rect 284 2335 285 2339
rect 430 2336 431 2340
rect 435 2336 436 2340
rect 430 2335 436 2336
rect 527 2339 533 2340
rect 527 2335 528 2339
rect 532 2338 533 2339
rect 698 2339 704 2340
rect 698 2338 699 2339
rect 532 2336 699 2338
rect 532 2335 533 2336
rect 279 2334 285 2335
rect 527 2334 533 2335
rect 698 2335 699 2336
rect 703 2335 704 2339
rect 718 2336 719 2340
rect 723 2336 724 2340
rect 718 2335 724 2336
rect 814 2339 821 2340
rect 814 2335 815 2339
rect 820 2335 821 2339
rect 998 2336 999 2340
rect 1003 2336 1004 2340
rect 998 2335 1004 2336
rect 1095 2339 1101 2340
rect 1095 2335 1096 2339
rect 1100 2338 1101 2339
rect 1258 2339 1264 2340
rect 1258 2338 1259 2339
rect 1100 2336 1259 2338
rect 1100 2335 1101 2336
rect 698 2334 704 2335
rect 814 2334 821 2335
rect 1095 2334 1101 2335
rect 1258 2335 1259 2336
rect 1263 2335 1264 2339
rect 1278 2336 1279 2340
rect 1283 2336 1284 2340
rect 1278 2335 1284 2336
rect 1374 2339 1381 2340
rect 1374 2335 1375 2339
rect 1380 2335 1381 2339
rect 1558 2336 1559 2340
rect 1563 2336 1564 2340
rect 1558 2335 1564 2336
rect 1655 2339 1661 2340
rect 1655 2335 1656 2339
rect 1660 2338 1661 2339
rect 1794 2339 1800 2340
rect 1794 2338 1795 2339
rect 1660 2336 1795 2338
rect 1660 2335 1661 2336
rect 1258 2334 1264 2335
rect 1374 2334 1381 2335
rect 1655 2334 1661 2335
rect 1794 2335 1795 2336
rect 1799 2335 1800 2339
rect 1814 2336 1815 2340
rect 1819 2336 1820 2340
rect 1814 2335 1820 2336
rect 1911 2339 1920 2340
rect 1911 2335 1912 2339
rect 1919 2335 1920 2339
rect 1794 2334 1800 2335
rect 1911 2334 1920 2335
rect 1934 2339 1940 2340
rect 1934 2335 1935 2339
rect 1939 2335 1940 2339
rect 1974 2339 1975 2343
rect 1979 2339 1980 2343
rect 2022 2340 2023 2344
rect 2027 2340 2028 2344
rect 2022 2339 2028 2340
rect 2114 2343 2125 2344
rect 2114 2339 2115 2343
rect 2119 2339 2120 2343
rect 2124 2339 2125 2343
rect 2302 2340 2303 2344
rect 2307 2340 2308 2344
rect 2302 2339 2308 2340
rect 2399 2343 2405 2344
rect 2399 2339 2400 2343
rect 2404 2342 2405 2343
rect 2578 2343 2584 2344
rect 2578 2342 2579 2343
rect 2404 2340 2579 2342
rect 2404 2339 2405 2340
rect 1974 2338 1980 2339
rect 2114 2338 2125 2339
rect 2399 2338 2405 2339
rect 2578 2339 2579 2340
rect 2583 2339 2584 2343
rect 2598 2340 2599 2344
rect 2603 2340 2604 2344
rect 2598 2339 2604 2340
rect 2690 2343 2701 2344
rect 2690 2339 2691 2343
rect 2695 2339 2696 2343
rect 2700 2339 2701 2343
rect 2886 2340 2887 2344
rect 2891 2340 2892 2344
rect 2886 2339 2892 2340
rect 2983 2343 2989 2344
rect 2983 2339 2984 2343
rect 2988 2342 2989 2343
rect 3154 2343 3160 2344
rect 3154 2342 3155 2343
rect 2988 2340 3155 2342
rect 2988 2339 2989 2340
rect 2578 2338 2584 2339
rect 2690 2338 2701 2339
rect 2983 2338 2989 2339
rect 3154 2339 3155 2340
rect 3159 2339 3160 2343
rect 3174 2340 3175 2344
rect 3179 2340 3180 2344
rect 3174 2339 3180 2340
rect 3271 2343 3277 2344
rect 3271 2339 3272 2343
rect 3276 2342 3277 2343
rect 3442 2343 3448 2344
rect 3442 2342 3443 2343
rect 3276 2340 3443 2342
rect 3276 2339 3277 2340
rect 3154 2338 3160 2339
rect 3271 2338 3277 2339
rect 3442 2339 3443 2340
rect 3447 2339 3448 2343
rect 3462 2340 3463 2344
rect 3467 2340 3468 2344
rect 3462 2339 3468 2340
rect 3558 2343 3565 2344
rect 3558 2339 3559 2343
rect 3564 2339 3565 2343
rect 3442 2338 3448 2339
rect 3558 2338 3565 2339
rect 3798 2343 3804 2344
rect 3798 2339 3799 2343
rect 3803 2339 3804 2343
rect 3798 2338 3804 2339
rect 1934 2334 1940 2335
rect 3838 2328 3844 2329
rect 5662 2328 5668 2329
rect 3838 2324 3839 2328
rect 3843 2324 3844 2328
rect 3838 2323 3844 2324
rect 3858 2327 3864 2328
rect 3858 2323 3859 2327
rect 3863 2323 3864 2327
rect 3858 2322 3864 2323
rect 4090 2327 4096 2328
rect 4090 2323 4091 2327
rect 4095 2323 4096 2327
rect 4090 2322 4096 2323
rect 4338 2327 4344 2328
rect 4338 2323 4339 2327
rect 4343 2323 4344 2327
rect 4338 2322 4344 2323
rect 4578 2327 4584 2328
rect 4578 2323 4579 2327
rect 4583 2323 4584 2327
rect 4578 2322 4584 2323
rect 4810 2327 4816 2328
rect 4810 2323 4811 2327
rect 4815 2323 4816 2327
rect 4810 2322 4816 2323
rect 5042 2327 5048 2328
rect 5042 2323 5043 2327
rect 5047 2323 5048 2327
rect 5042 2322 5048 2323
rect 5282 2327 5288 2328
rect 5282 2323 5283 2327
rect 5287 2323 5288 2327
rect 5282 2322 5288 2323
rect 5514 2327 5520 2328
rect 5514 2323 5515 2327
rect 5519 2323 5520 2327
rect 5662 2324 5663 2328
rect 5667 2324 5668 2328
rect 5662 2323 5668 2324
rect 5514 2322 5520 2323
rect 3886 2312 3892 2313
rect 4118 2312 4124 2313
rect 4366 2312 4372 2313
rect 4606 2312 4612 2313
rect 4838 2312 4844 2313
rect 5070 2312 5076 2313
rect 5310 2312 5316 2313
rect 5542 2312 5548 2313
rect 3838 2311 3844 2312
rect 3838 2307 3839 2311
rect 3843 2307 3844 2311
rect 3886 2308 3887 2312
rect 3891 2308 3892 2312
rect 3886 2307 3892 2308
rect 3983 2311 3989 2312
rect 3983 2307 3984 2311
rect 3988 2310 3989 2311
rect 4098 2311 4104 2312
rect 4098 2310 4099 2311
rect 3988 2308 4099 2310
rect 3988 2307 3989 2308
rect 3838 2306 3844 2307
rect 3983 2306 3989 2307
rect 4098 2307 4099 2308
rect 4103 2307 4104 2311
rect 4118 2308 4119 2312
rect 4123 2308 4124 2312
rect 4118 2307 4124 2308
rect 4210 2311 4221 2312
rect 4210 2307 4211 2311
rect 4215 2307 4216 2311
rect 4220 2307 4221 2311
rect 4366 2308 4367 2312
rect 4371 2308 4372 2312
rect 4366 2307 4372 2308
rect 4463 2311 4469 2312
rect 4463 2307 4464 2311
rect 4468 2310 4469 2311
rect 4586 2311 4592 2312
rect 4586 2310 4587 2311
rect 4468 2308 4587 2310
rect 4468 2307 4469 2308
rect 4098 2306 4104 2307
rect 4210 2306 4221 2307
rect 4463 2306 4469 2307
rect 4586 2307 4587 2308
rect 4591 2307 4592 2311
rect 4606 2308 4607 2312
rect 4611 2308 4612 2312
rect 4606 2307 4612 2308
rect 4703 2311 4709 2312
rect 4703 2307 4704 2311
rect 4708 2310 4709 2311
rect 4818 2311 4824 2312
rect 4818 2310 4819 2311
rect 4708 2308 4819 2310
rect 4708 2307 4709 2308
rect 4586 2306 4592 2307
rect 4703 2306 4709 2307
rect 4818 2307 4819 2308
rect 4823 2307 4824 2311
rect 4838 2308 4839 2312
rect 4843 2308 4844 2312
rect 4838 2307 4844 2308
rect 4935 2311 4941 2312
rect 4935 2307 4936 2311
rect 4940 2310 4941 2311
rect 5050 2311 5056 2312
rect 5050 2310 5051 2311
rect 4940 2308 5051 2310
rect 4940 2307 4941 2308
rect 4818 2306 4824 2307
rect 4935 2306 4941 2307
rect 5050 2307 5051 2308
rect 5055 2307 5056 2311
rect 5070 2308 5071 2312
rect 5075 2308 5076 2312
rect 5070 2307 5076 2308
rect 5166 2311 5173 2312
rect 5166 2307 5167 2311
rect 5172 2307 5173 2311
rect 5310 2308 5311 2312
rect 5315 2308 5316 2312
rect 5310 2307 5316 2308
rect 5406 2311 5413 2312
rect 5406 2307 5407 2311
rect 5412 2307 5413 2311
rect 5542 2308 5543 2312
rect 5547 2308 5548 2312
rect 5542 2307 5548 2308
rect 5634 2311 5645 2312
rect 5634 2307 5635 2311
rect 5639 2307 5640 2311
rect 5644 2307 5645 2311
rect 5050 2306 5056 2307
rect 5166 2306 5173 2307
rect 5406 2306 5413 2307
rect 5634 2306 5645 2307
rect 5662 2311 5668 2312
rect 5662 2307 5663 2311
rect 5667 2307 5668 2311
rect 5662 2306 5668 2307
rect 1974 2273 1980 2274
rect 3798 2273 3804 2274
rect 1974 2269 1975 2273
rect 1979 2269 1980 2273
rect 1974 2268 1980 2269
rect 2022 2272 2028 2273
rect 2158 2272 2164 2273
rect 2294 2272 2300 2273
rect 2446 2272 2452 2273
rect 2606 2272 2612 2273
rect 2766 2272 2772 2273
rect 2926 2272 2932 2273
rect 3078 2272 3084 2273
rect 3230 2272 3236 2273
rect 3382 2272 3388 2273
rect 3542 2272 3548 2273
rect 3678 2272 3684 2273
rect 2022 2268 2023 2272
rect 2027 2268 2028 2272
rect 2022 2267 2028 2268
rect 2119 2271 2128 2272
rect 2119 2267 2120 2271
rect 2127 2267 2128 2271
rect 2158 2268 2159 2272
rect 2163 2268 2164 2272
rect 2158 2267 2164 2268
rect 2255 2271 2264 2272
rect 2255 2267 2256 2271
rect 2263 2267 2264 2271
rect 2294 2268 2295 2272
rect 2299 2268 2300 2272
rect 2294 2267 2300 2268
rect 2391 2271 2397 2272
rect 2391 2267 2392 2271
rect 2396 2270 2397 2271
rect 2407 2271 2413 2272
rect 2407 2270 2408 2271
rect 2396 2268 2408 2270
rect 2396 2267 2397 2268
rect 2119 2266 2128 2267
rect 2255 2266 2264 2267
rect 2391 2266 2397 2267
rect 2407 2267 2408 2268
rect 2412 2267 2413 2271
rect 2446 2268 2447 2272
rect 2451 2268 2452 2272
rect 2446 2267 2452 2268
rect 2538 2271 2549 2272
rect 2538 2267 2539 2271
rect 2543 2267 2544 2271
rect 2548 2267 2549 2271
rect 2606 2268 2607 2272
rect 2611 2268 2612 2272
rect 2606 2267 2612 2268
rect 2702 2271 2709 2272
rect 2702 2267 2703 2271
rect 2708 2267 2709 2271
rect 2766 2268 2767 2272
rect 2771 2268 2772 2272
rect 2766 2267 2772 2268
rect 2858 2271 2869 2272
rect 2858 2267 2859 2271
rect 2863 2267 2864 2271
rect 2868 2267 2869 2271
rect 2926 2268 2927 2272
rect 2931 2268 2932 2272
rect 2926 2267 2932 2268
rect 3018 2271 3029 2272
rect 3018 2267 3019 2271
rect 3023 2267 3024 2271
rect 3028 2267 3029 2271
rect 3078 2268 3079 2272
rect 3083 2268 3084 2272
rect 3078 2267 3084 2268
rect 3174 2271 3181 2272
rect 3174 2267 3175 2271
rect 3180 2267 3181 2271
rect 3230 2268 3231 2272
rect 3235 2268 3236 2272
rect 3230 2267 3236 2268
rect 3326 2271 3333 2272
rect 3326 2267 3327 2271
rect 3332 2267 3333 2271
rect 3382 2268 3383 2272
rect 3387 2268 3388 2272
rect 3382 2267 3388 2268
rect 3478 2271 3485 2272
rect 3478 2267 3479 2271
rect 3484 2267 3485 2271
rect 3542 2268 3543 2272
rect 3547 2268 3548 2272
rect 3542 2267 3548 2268
rect 3639 2271 3648 2272
rect 3639 2267 3640 2271
rect 3647 2267 3648 2271
rect 3678 2268 3679 2272
rect 3683 2268 3684 2272
rect 3678 2267 3684 2268
rect 3775 2271 3781 2272
rect 3775 2267 3776 2271
rect 3780 2270 3781 2271
rect 3790 2271 3796 2272
rect 3790 2270 3791 2271
rect 3780 2268 3791 2270
rect 3780 2267 3781 2268
rect 2407 2266 2413 2267
rect 2538 2266 2549 2267
rect 2702 2266 2709 2267
rect 2858 2266 2869 2267
rect 3018 2266 3029 2267
rect 3174 2266 3181 2267
rect 3326 2266 3333 2267
rect 3478 2266 3485 2267
rect 3639 2266 3648 2267
rect 3775 2266 3781 2267
rect 3790 2267 3791 2268
rect 3795 2267 3796 2271
rect 3798 2269 3799 2273
rect 3803 2269 3804 2273
rect 3798 2268 3804 2269
rect 3790 2266 3796 2267
rect 110 2265 116 2266
rect 1934 2265 1940 2266
rect 110 2261 111 2265
rect 115 2261 116 2265
rect 110 2260 116 2261
rect 158 2264 164 2265
rect 422 2264 428 2265
rect 710 2264 716 2265
rect 998 2264 1004 2265
rect 1294 2264 1300 2265
rect 158 2260 159 2264
rect 163 2260 164 2264
rect 158 2259 164 2260
rect 255 2263 261 2264
rect 255 2259 256 2263
rect 260 2262 261 2263
rect 295 2263 301 2264
rect 295 2262 296 2263
rect 260 2260 296 2262
rect 260 2259 261 2260
rect 255 2258 261 2259
rect 295 2259 296 2260
rect 300 2259 301 2263
rect 422 2260 423 2264
rect 427 2260 428 2264
rect 422 2259 428 2260
rect 518 2263 525 2264
rect 518 2259 519 2263
rect 524 2259 525 2263
rect 710 2260 711 2264
rect 715 2260 716 2264
rect 710 2259 716 2260
rect 807 2263 816 2264
rect 807 2259 808 2263
rect 815 2259 816 2263
rect 998 2260 999 2264
rect 1003 2260 1004 2264
rect 998 2259 1004 2260
rect 1094 2263 1101 2264
rect 1094 2259 1095 2263
rect 1100 2259 1101 2263
rect 1294 2260 1295 2264
rect 1299 2260 1300 2264
rect 1294 2259 1300 2260
rect 1386 2263 1397 2264
rect 1386 2259 1387 2263
rect 1391 2259 1392 2263
rect 1396 2259 1397 2263
rect 1934 2261 1935 2265
rect 1939 2261 1940 2265
rect 1934 2260 1940 2261
rect 295 2258 301 2259
rect 518 2258 525 2259
rect 807 2258 816 2259
rect 1094 2258 1101 2259
rect 1386 2258 1397 2259
rect 1994 2257 2000 2258
rect 1974 2256 1980 2257
rect 1974 2252 1975 2256
rect 1979 2252 1980 2256
rect 1994 2253 1995 2257
rect 1999 2253 2000 2257
rect 1994 2252 2000 2253
rect 2130 2257 2136 2258
rect 2130 2253 2131 2257
rect 2135 2253 2136 2257
rect 2130 2252 2136 2253
rect 2266 2257 2272 2258
rect 2266 2253 2267 2257
rect 2271 2253 2272 2257
rect 2266 2252 2272 2253
rect 2418 2257 2424 2258
rect 2418 2253 2419 2257
rect 2423 2253 2424 2257
rect 2418 2252 2424 2253
rect 2578 2257 2584 2258
rect 2578 2253 2579 2257
rect 2583 2253 2584 2257
rect 2578 2252 2584 2253
rect 2738 2257 2744 2258
rect 2738 2253 2739 2257
rect 2743 2253 2744 2257
rect 2738 2252 2744 2253
rect 2898 2257 2904 2258
rect 2898 2253 2899 2257
rect 2903 2253 2904 2257
rect 2898 2252 2904 2253
rect 3050 2257 3056 2258
rect 3050 2253 3051 2257
rect 3055 2253 3056 2257
rect 3050 2252 3056 2253
rect 3202 2257 3208 2258
rect 3202 2253 3203 2257
rect 3207 2253 3208 2257
rect 3202 2252 3208 2253
rect 3354 2257 3360 2258
rect 3354 2253 3355 2257
rect 3359 2253 3360 2257
rect 3354 2252 3360 2253
rect 3514 2257 3520 2258
rect 3514 2253 3515 2257
rect 3519 2253 3520 2257
rect 3514 2252 3520 2253
rect 3650 2257 3656 2258
rect 3650 2253 3651 2257
rect 3655 2253 3656 2257
rect 3650 2252 3656 2253
rect 3798 2256 3804 2257
rect 3798 2252 3799 2256
rect 3803 2252 3804 2256
rect 1974 2251 1980 2252
rect 3798 2251 3804 2252
rect 130 2249 136 2250
rect 110 2248 116 2249
rect 110 2244 111 2248
rect 115 2244 116 2248
rect 130 2245 131 2249
rect 135 2245 136 2249
rect 130 2244 136 2245
rect 394 2249 400 2250
rect 394 2245 395 2249
rect 399 2245 400 2249
rect 394 2244 400 2245
rect 682 2249 688 2250
rect 682 2245 683 2249
rect 687 2245 688 2249
rect 682 2244 688 2245
rect 970 2249 976 2250
rect 970 2245 971 2249
rect 975 2245 976 2249
rect 970 2244 976 2245
rect 1266 2249 1272 2250
rect 1266 2245 1267 2249
rect 1271 2245 1272 2249
rect 1266 2244 1272 2245
rect 1934 2248 1940 2249
rect 1934 2244 1935 2248
rect 1939 2244 1940 2248
rect 110 2243 116 2244
rect 1934 2243 1940 2244
rect 3146 2239 3152 2240
rect 3146 2235 3147 2239
rect 3151 2238 3152 2239
rect 3326 2239 3332 2240
rect 3326 2238 3327 2239
rect 3151 2236 3327 2238
rect 3151 2235 3152 2236
rect 3146 2234 3152 2235
rect 3326 2235 3327 2236
rect 3331 2235 3332 2239
rect 3326 2234 3332 2235
rect 3838 2229 3844 2230
rect 5662 2229 5668 2230
rect 3838 2225 3839 2229
rect 3843 2225 3844 2229
rect 3838 2224 3844 2225
rect 4590 2228 4596 2229
rect 4726 2228 4732 2229
rect 4862 2228 4868 2229
rect 4998 2228 5004 2229
rect 5134 2228 5140 2229
rect 5270 2228 5276 2229
rect 5406 2228 5412 2229
rect 5542 2228 5548 2229
rect 4590 2224 4591 2228
rect 4595 2224 4596 2228
rect 4590 2223 4596 2224
rect 4687 2227 4696 2228
rect 4687 2223 4688 2227
rect 4695 2223 4696 2227
rect 4726 2224 4727 2228
rect 4731 2224 4732 2228
rect 4726 2223 4732 2224
rect 4823 2227 4832 2228
rect 4823 2223 4824 2227
rect 4831 2223 4832 2227
rect 4862 2224 4863 2228
rect 4867 2224 4868 2228
rect 4862 2223 4868 2224
rect 4959 2227 4968 2228
rect 4959 2223 4960 2227
rect 4967 2223 4968 2227
rect 4998 2224 4999 2228
rect 5003 2224 5004 2228
rect 4998 2223 5004 2224
rect 5095 2227 5104 2228
rect 5095 2223 5096 2227
rect 5103 2223 5104 2227
rect 5134 2224 5135 2228
rect 5139 2224 5140 2228
rect 5134 2223 5140 2224
rect 5231 2227 5240 2228
rect 5231 2223 5232 2227
rect 5239 2223 5240 2227
rect 5270 2224 5271 2228
rect 5275 2224 5276 2228
rect 5270 2223 5276 2224
rect 5367 2227 5376 2228
rect 5367 2223 5368 2227
rect 5375 2223 5376 2227
rect 5406 2224 5407 2228
rect 5411 2224 5412 2228
rect 5406 2223 5412 2224
rect 5498 2227 5509 2228
rect 5498 2223 5499 2227
rect 5503 2223 5504 2227
rect 5508 2223 5509 2227
rect 5542 2224 5543 2228
rect 5547 2224 5548 2228
rect 5542 2223 5548 2224
rect 5639 2227 5648 2228
rect 5639 2223 5640 2227
rect 5647 2223 5648 2227
rect 5662 2225 5663 2229
rect 5667 2225 5668 2229
rect 5662 2224 5668 2225
rect 4687 2222 4696 2223
rect 4823 2222 4832 2223
rect 4959 2222 4968 2223
rect 5095 2222 5104 2223
rect 5231 2222 5240 2223
rect 5367 2222 5376 2223
rect 5498 2222 5509 2223
rect 5639 2222 5648 2223
rect 4562 2213 4568 2214
rect 3838 2212 3844 2213
rect 3838 2208 3839 2212
rect 3843 2208 3844 2212
rect 4562 2209 4563 2213
rect 4567 2209 4568 2213
rect 4562 2208 4568 2209
rect 4698 2213 4704 2214
rect 4698 2209 4699 2213
rect 4703 2209 4704 2213
rect 4698 2208 4704 2209
rect 4834 2213 4840 2214
rect 4834 2209 4835 2213
rect 4839 2209 4840 2213
rect 4834 2208 4840 2209
rect 4970 2213 4976 2214
rect 4970 2209 4971 2213
rect 4975 2209 4976 2213
rect 4970 2208 4976 2209
rect 5106 2213 5112 2214
rect 5106 2209 5107 2213
rect 5111 2209 5112 2213
rect 5106 2208 5112 2209
rect 5242 2213 5248 2214
rect 5242 2209 5243 2213
rect 5247 2209 5248 2213
rect 5242 2208 5248 2209
rect 5378 2213 5384 2214
rect 5378 2209 5379 2213
rect 5383 2209 5384 2213
rect 5378 2208 5384 2209
rect 5514 2213 5520 2214
rect 5514 2209 5515 2213
rect 5519 2209 5520 2213
rect 5514 2208 5520 2209
rect 5662 2212 5668 2213
rect 5662 2208 5663 2212
rect 5667 2208 5668 2212
rect 2114 2207 2120 2208
rect 2114 2206 2115 2207
rect 2093 2204 2115 2206
rect 2114 2203 2115 2204
rect 2119 2203 2120 2207
rect 2114 2202 2120 2203
rect 2122 2207 2128 2208
rect 2122 2203 2123 2207
rect 2127 2206 2128 2207
rect 2258 2207 2264 2208
rect 2127 2204 2137 2206
rect 2127 2203 2128 2204
rect 2122 2202 2128 2203
rect 2258 2203 2259 2207
rect 2263 2206 2264 2207
rect 2407 2207 2413 2208
rect 2263 2204 2273 2206
rect 2263 2203 2264 2204
rect 2258 2202 2264 2203
rect 2407 2203 2408 2207
rect 2412 2206 2413 2207
rect 2850 2207 2856 2208
rect 2850 2206 2851 2207
rect 2412 2204 2425 2206
rect 2412 2203 2413 2204
rect 2407 2202 2413 2203
rect 250 2199 256 2200
rect 250 2198 251 2199
rect 229 2196 251 2198
rect 250 2195 251 2196
rect 255 2195 256 2199
rect 250 2194 256 2195
rect 295 2199 301 2200
rect 295 2195 296 2199
rect 300 2198 301 2199
rect 810 2199 816 2200
rect 300 2196 401 2198
rect 300 2195 301 2196
rect 295 2194 301 2195
rect 780 2190 782 2197
rect 810 2195 811 2199
rect 815 2198 816 2199
rect 1374 2199 1380 2200
rect 1374 2198 1375 2199
rect 815 2196 977 2198
rect 1365 2196 1375 2198
rect 815 2195 816 2196
rect 810 2194 816 2195
rect 1374 2195 1375 2196
rect 1379 2195 1380 2199
rect 2676 2198 2678 2205
rect 2837 2204 2851 2206
rect 2850 2203 2851 2204
rect 2855 2203 2856 2207
rect 3146 2207 3152 2208
rect 2850 2202 2856 2203
rect 2858 2199 2864 2200
rect 2858 2198 2859 2199
rect 2676 2196 2859 2198
rect 1374 2194 1380 2195
rect 2858 2195 2859 2196
rect 2863 2195 2864 2199
rect 2996 2198 2998 2205
rect 3146 2203 3147 2207
rect 3151 2203 3152 2207
rect 3422 2207 3428 2208
rect 3146 2202 3152 2203
rect 3174 2199 3180 2200
rect 3174 2198 3175 2199
rect 2996 2196 3175 2198
rect 2858 2194 2864 2195
rect 3174 2195 3175 2196
rect 3179 2195 3180 2199
rect 3300 2198 3302 2205
rect 3422 2203 3423 2207
rect 3427 2203 3428 2207
rect 3422 2202 3428 2203
rect 3558 2207 3564 2208
rect 3558 2203 3559 2207
rect 3563 2203 3564 2207
rect 3558 2202 3564 2203
rect 3642 2207 3648 2208
rect 3838 2207 3844 2208
rect 5662 2207 5668 2208
rect 3642 2203 3643 2207
rect 3647 2206 3648 2207
rect 3647 2204 3657 2206
rect 3647 2203 3648 2204
rect 3642 2202 3648 2203
rect 3478 2199 3484 2200
rect 3478 2198 3479 2199
rect 3300 2196 3479 2198
rect 3174 2194 3180 2195
rect 3478 2195 3479 2196
rect 3483 2195 3484 2199
rect 3478 2194 3484 2195
rect 1386 2191 1392 2192
rect 1386 2190 1387 2191
rect 780 2188 1387 2190
rect 1386 2187 1387 2188
rect 1391 2187 1392 2191
rect 1386 2186 1392 2187
rect 2538 2175 2544 2176
rect 2538 2174 2539 2175
rect 2340 2172 2539 2174
rect 2340 2170 2342 2172
rect 2538 2171 2539 2172
rect 2543 2171 2544 2175
rect 3774 2175 3780 2176
rect 3774 2174 3775 2175
rect 2538 2170 2544 2171
rect 3468 2172 3775 2174
rect 2332 2168 2342 2170
rect 2332 2166 2334 2168
rect 2229 2164 2334 2166
rect 3018 2167 3024 2168
rect 2338 2163 2344 2164
rect 526 2159 532 2160
rect 526 2158 527 2159
rect 259 2156 527 2158
rect 259 2154 261 2156
rect 526 2155 527 2156
rect 531 2155 532 2159
rect 2338 2159 2339 2163
rect 2343 2159 2344 2163
rect 2338 2158 2344 2159
rect 2538 2163 2544 2164
rect 2538 2159 2539 2163
rect 2543 2159 2544 2163
rect 2538 2158 2544 2159
rect 2738 2163 2744 2164
rect 2738 2159 2739 2163
rect 2743 2159 2744 2163
rect 3018 2163 3019 2167
rect 3023 2163 3024 2167
rect 3468 2166 3470 2172
rect 3774 2171 3775 2172
rect 3779 2171 3780 2175
rect 3774 2170 3780 2171
rect 3397 2164 3470 2166
rect 3018 2162 3024 2163
rect 3122 2163 3128 2164
rect 2738 2158 2744 2159
rect 3122 2159 3123 2163
rect 3127 2159 3128 2163
rect 3122 2158 3128 2159
rect 3578 2163 3584 2164
rect 3578 2159 3579 2163
rect 3583 2159 3584 2163
rect 3578 2158 3584 2159
rect 3658 2163 3664 2164
rect 3658 2159 3659 2163
rect 3663 2159 3664 2163
rect 4690 2163 4696 2164
rect 3658 2158 3664 2159
rect 526 2154 532 2155
rect 1094 2155 1100 2156
rect 229 2152 261 2154
rect 498 2151 504 2152
rect 498 2147 499 2151
rect 503 2147 504 2151
rect 498 2146 504 2147
rect 738 2151 744 2152
rect 738 2147 739 2151
rect 743 2147 744 2151
rect 1094 2151 1095 2155
rect 1099 2151 1100 2155
rect 2118 2155 2124 2156
rect 2118 2154 2119 2155
rect 1885 2152 2119 2154
rect 1094 2150 1100 2151
rect 1450 2151 1456 2152
rect 738 2146 744 2147
rect 1450 2147 1451 2151
rect 1455 2147 1456 2151
rect 2118 2151 2119 2152
rect 2123 2151 2124 2155
rect 4660 2154 4662 2161
rect 4690 2159 4691 2163
rect 4695 2162 4696 2163
rect 4826 2163 4832 2164
rect 4695 2160 4705 2162
rect 4695 2159 4696 2160
rect 4690 2158 4696 2159
rect 4826 2159 4827 2163
rect 4831 2162 4832 2163
rect 4962 2163 4968 2164
rect 4831 2160 4841 2162
rect 4831 2159 4832 2160
rect 4826 2158 4832 2159
rect 4962 2159 4963 2163
rect 4967 2162 4968 2163
rect 5098 2163 5104 2164
rect 4967 2160 4977 2162
rect 4967 2159 4968 2160
rect 4962 2158 4968 2159
rect 5098 2159 5099 2163
rect 5103 2162 5104 2163
rect 5234 2163 5240 2164
rect 5103 2160 5113 2162
rect 5103 2159 5104 2160
rect 5098 2158 5104 2159
rect 5234 2159 5235 2163
rect 5239 2162 5240 2163
rect 5370 2163 5376 2164
rect 5239 2160 5249 2162
rect 5239 2159 5240 2160
rect 5234 2158 5240 2159
rect 5370 2159 5371 2163
rect 5375 2162 5376 2163
rect 5634 2163 5640 2164
rect 5634 2162 5635 2163
rect 5375 2160 5385 2162
rect 5613 2160 5635 2162
rect 5375 2159 5376 2160
rect 5370 2158 5376 2159
rect 5634 2159 5635 2160
rect 5639 2159 5640 2163
rect 5634 2158 5640 2159
rect 5166 2155 5172 2156
rect 5166 2154 5167 2155
rect 4660 2152 5167 2154
rect 2118 2150 2124 2151
rect 5166 2151 5167 2152
rect 5171 2151 5172 2155
rect 5166 2150 5172 2151
rect 1450 2146 1456 2147
rect 5350 2123 5356 2124
rect 5350 2122 5351 2123
rect 5299 2120 5351 2122
rect 5299 2118 5301 2120
rect 5350 2119 5351 2120
rect 5355 2119 5356 2123
rect 5350 2118 5356 2119
rect 1974 2116 1980 2117
rect 3798 2116 3804 2117
rect 5196 2116 5301 2118
rect 498 2115 504 2116
rect 498 2111 499 2115
rect 503 2114 504 2115
rect 854 2115 860 2116
rect 854 2114 855 2115
rect 503 2112 855 2114
rect 503 2111 504 2112
rect 498 2110 504 2111
rect 854 2111 855 2112
rect 859 2111 860 2115
rect 1974 2112 1975 2116
rect 1979 2112 1980 2116
rect 1974 2111 1980 2112
rect 2130 2115 2136 2116
rect 2130 2111 2131 2115
rect 2135 2111 2136 2115
rect 854 2110 860 2111
rect 2130 2110 2136 2111
rect 2330 2115 2336 2116
rect 2330 2111 2331 2115
rect 2335 2111 2336 2115
rect 2330 2110 2336 2111
rect 2530 2115 2536 2116
rect 2530 2111 2531 2115
rect 2535 2111 2536 2115
rect 2530 2110 2536 2111
rect 2730 2115 2736 2116
rect 2730 2111 2731 2115
rect 2735 2111 2736 2115
rect 2730 2110 2736 2111
rect 2922 2115 2928 2116
rect 2922 2111 2923 2115
rect 2927 2111 2928 2115
rect 2922 2110 2928 2111
rect 3114 2115 3120 2116
rect 3114 2111 3115 2115
rect 3119 2111 3120 2115
rect 3114 2110 3120 2111
rect 3298 2115 3304 2116
rect 3298 2111 3299 2115
rect 3303 2111 3304 2115
rect 3298 2110 3304 2111
rect 3482 2115 3488 2116
rect 3482 2111 3483 2115
rect 3487 2111 3488 2115
rect 3482 2110 3488 2111
rect 3650 2115 3656 2116
rect 3650 2111 3651 2115
rect 3655 2111 3656 2115
rect 3798 2112 3799 2116
rect 3803 2112 3804 2116
rect 5082 2115 5088 2116
rect 5082 2114 5083 2115
rect 5053 2112 5083 2114
rect 3798 2111 3804 2112
rect 5082 2111 5083 2112
rect 5087 2111 5088 2115
rect 5196 2114 5198 2116
rect 5410 2115 5416 2116
rect 5410 2114 5411 2115
rect 5189 2112 5198 2114
rect 5325 2112 5411 2114
rect 3650 2110 3656 2111
rect 5082 2110 5088 2111
rect 5410 2111 5411 2112
rect 5415 2111 5416 2115
rect 5410 2110 5416 2111
rect 110 2104 116 2105
rect 1934 2104 1940 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 130 2103 136 2104
rect 130 2099 131 2103
rect 135 2099 136 2103
rect 130 2098 136 2099
rect 402 2103 408 2104
rect 402 2099 403 2103
rect 407 2099 408 2103
rect 402 2098 408 2099
rect 730 2103 736 2104
rect 730 2099 731 2103
rect 735 2099 736 2103
rect 730 2098 736 2099
rect 1082 2103 1088 2104
rect 1082 2099 1083 2103
rect 1087 2099 1088 2103
rect 1082 2098 1088 2099
rect 1442 2103 1448 2104
rect 1442 2099 1443 2103
rect 1447 2099 1448 2103
rect 1442 2098 1448 2099
rect 1786 2103 1792 2104
rect 1786 2099 1787 2103
rect 1791 2099 1792 2103
rect 1934 2100 1935 2104
rect 1939 2100 1940 2104
rect 2158 2100 2164 2101
rect 2358 2100 2364 2101
rect 2558 2100 2564 2101
rect 2758 2100 2764 2101
rect 2950 2100 2956 2101
rect 3142 2100 3148 2101
rect 3326 2100 3332 2101
rect 3510 2100 3516 2101
rect 3678 2100 3684 2101
rect 1934 2099 1940 2100
rect 1974 2099 1980 2100
rect 1786 2098 1792 2099
rect 1974 2095 1975 2099
rect 1979 2095 1980 2099
rect 2158 2096 2159 2100
rect 2163 2096 2164 2100
rect 2158 2095 2164 2096
rect 2255 2099 2261 2100
rect 2255 2095 2256 2099
rect 2260 2098 2261 2099
rect 2338 2099 2344 2100
rect 2338 2098 2339 2099
rect 2260 2096 2339 2098
rect 2260 2095 2261 2096
rect 1974 2094 1980 2095
rect 2255 2094 2261 2095
rect 2338 2095 2339 2096
rect 2343 2095 2344 2099
rect 2358 2096 2359 2100
rect 2363 2096 2364 2100
rect 2358 2095 2364 2096
rect 2455 2099 2461 2100
rect 2455 2095 2456 2099
rect 2460 2098 2461 2099
rect 2538 2099 2544 2100
rect 2538 2098 2539 2099
rect 2460 2096 2539 2098
rect 2460 2095 2461 2096
rect 2338 2094 2344 2095
rect 2455 2094 2461 2095
rect 2538 2095 2539 2096
rect 2543 2095 2544 2099
rect 2558 2096 2559 2100
rect 2563 2096 2564 2100
rect 2558 2095 2564 2096
rect 2655 2099 2661 2100
rect 2655 2095 2656 2099
rect 2660 2098 2661 2099
rect 2738 2099 2744 2100
rect 2738 2098 2739 2099
rect 2660 2096 2739 2098
rect 2660 2095 2661 2096
rect 2538 2094 2544 2095
rect 2655 2094 2661 2095
rect 2738 2095 2739 2096
rect 2743 2095 2744 2099
rect 2758 2096 2759 2100
rect 2763 2096 2764 2100
rect 2758 2095 2764 2096
rect 2850 2099 2861 2100
rect 2850 2095 2851 2099
rect 2855 2095 2856 2099
rect 2860 2095 2861 2099
rect 2950 2096 2951 2100
rect 2955 2096 2956 2100
rect 2950 2095 2956 2096
rect 3047 2099 3053 2100
rect 3047 2095 3048 2099
rect 3052 2098 3053 2099
rect 3122 2099 3128 2100
rect 3122 2098 3123 2099
rect 3052 2096 3123 2098
rect 3052 2095 3053 2096
rect 2738 2094 2744 2095
rect 2850 2094 2861 2095
rect 3047 2094 3053 2095
rect 3122 2095 3123 2096
rect 3127 2095 3128 2099
rect 3142 2096 3143 2100
rect 3147 2096 3148 2100
rect 3142 2095 3148 2096
rect 3238 2099 3245 2100
rect 3238 2095 3239 2099
rect 3244 2095 3245 2099
rect 3326 2096 3327 2100
rect 3331 2096 3332 2100
rect 3326 2095 3332 2096
rect 3422 2099 3429 2100
rect 3422 2095 3423 2099
rect 3428 2095 3429 2099
rect 3510 2096 3511 2100
rect 3515 2096 3516 2100
rect 3510 2095 3516 2096
rect 3607 2099 3613 2100
rect 3607 2095 3608 2099
rect 3612 2098 3613 2099
rect 3658 2099 3664 2100
rect 3658 2098 3659 2099
rect 3612 2096 3659 2098
rect 3612 2095 3613 2096
rect 3122 2094 3128 2095
rect 3238 2094 3245 2095
rect 3422 2094 3429 2095
rect 3607 2094 3613 2095
rect 3658 2095 3659 2096
rect 3663 2095 3664 2099
rect 3678 2096 3679 2100
rect 3683 2096 3684 2100
rect 3678 2095 3684 2096
rect 3774 2099 3781 2100
rect 3774 2095 3775 2099
rect 3780 2095 3781 2099
rect 3658 2094 3664 2095
rect 3774 2094 3781 2095
rect 3798 2099 3804 2100
rect 3798 2095 3799 2099
rect 3803 2095 3804 2099
rect 3798 2094 3804 2095
rect 158 2088 164 2089
rect 430 2088 436 2089
rect 758 2088 764 2089
rect 1110 2088 1116 2089
rect 1470 2088 1476 2089
rect 1814 2088 1820 2089
rect 110 2087 116 2088
rect 110 2083 111 2087
rect 115 2083 116 2087
rect 158 2084 159 2088
rect 163 2084 164 2088
rect 158 2083 164 2084
rect 250 2087 261 2088
rect 250 2083 251 2087
rect 255 2083 256 2087
rect 260 2083 261 2087
rect 430 2084 431 2088
rect 435 2084 436 2088
rect 430 2083 436 2084
rect 526 2087 533 2088
rect 526 2083 527 2087
rect 532 2083 533 2087
rect 758 2084 759 2088
rect 763 2084 764 2088
rect 758 2083 764 2084
rect 854 2087 861 2088
rect 854 2083 855 2087
rect 860 2083 861 2087
rect 1110 2084 1111 2088
rect 1115 2084 1116 2088
rect 1110 2083 1116 2084
rect 1207 2087 1213 2088
rect 1207 2083 1208 2087
rect 1212 2086 1213 2087
rect 1450 2087 1456 2088
rect 1450 2086 1451 2087
rect 1212 2084 1451 2086
rect 1212 2083 1213 2084
rect 110 2082 116 2083
rect 250 2082 261 2083
rect 526 2082 533 2083
rect 854 2082 861 2083
rect 1207 2082 1213 2083
rect 1450 2083 1451 2084
rect 1455 2083 1456 2087
rect 1470 2084 1471 2088
rect 1475 2084 1476 2088
rect 1470 2083 1476 2084
rect 1566 2087 1573 2088
rect 1566 2083 1567 2087
rect 1572 2083 1573 2087
rect 1814 2084 1815 2088
rect 1819 2084 1820 2088
rect 1814 2083 1820 2084
rect 1910 2087 1917 2088
rect 1910 2083 1911 2087
rect 1916 2083 1917 2087
rect 1450 2082 1456 2083
rect 1566 2082 1573 2083
rect 1910 2082 1917 2083
rect 1934 2087 1940 2088
rect 1934 2083 1935 2087
rect 1939 2083 1940 2087
rect 1934 2082 1940 2083
rect 3838 2064 3844 2065
rect 5662 2064 5668 2065
rect 3838 2060 3839 2064
rect 3843 2060 3844 2064
rect 3838 2059 3844 2060
rect 4954 2063 4960 2064
rect 4954 2059 4955 2063
rect 4959 2059 4960 2063
rect 4954 2058 4960 2059
rect 5090 2063 5096 2064
rect 5090 2059 5091 2063
rect 5095 2059 5096 2063
rect 5090 2058 5096 2059
rect 5226 2063 5232 2064
rect 5226 2059 5227 2063
rect 5231 2059 5232 2063
rect 5662 2060 5663 2064
rect 5667 2060 5668 2064
rect 5662 2059 5668 2060
rect 5226 2058 5232 2059
rect 5082 2055 5088 2056
rect 5082 2051 5083 2055
rect 5087 2054 5088 2055
rect 5087 2052 5218 2054
rect 5087 2051 5088 2052
rect 5082 2050 5088 2051
rect 4982 2048 4988 2049
rect 5118 2048 5124 2049
rect 5216 2048 5218 2052
rect 5254 2048 5260 2049
rect 3838 2047 3844 2048
rect 3838 2043 3839 2047
rect 3843 2043 3844 2047
rect 4982 2044 4983 2048
rect 4987 2044 4988 2048
rect 4982 2043 4988 2044
rect 5074 2047 5085 2048
rect 5074 2043 5075 2047
rect 5079 2043 5080 2047
rect 5084 2043 5085 2047
rect 5118 2044 5119 2048
rect 5123 2044 5124 2048
rect 5118 2043 5124 2044
rect 5215 2047 5221 2048
rect 5215 2043 5216 2047
rect 5220 2043 5221 2047
rect 5254 2044 5255 2048
rect 5259 2044 5260 2048
rect 5254 2043 5260 2044
rect 5350 2047 5357 2048
rect 5350 2043 5351 2047
rect 5356 2043 5357 2047
rect 3838 2042 3844 2043
rect 5074 2042 5085 2043
rect 5215 2042 5221 2043
rect 5350 2042 5357 2043
rect 5662 2047 5668 2048
rect 5662 2043 5663 2047
rect 5667 2043 5668 2047
rect 5662 2042 5668 2043
rect 1974 2033 1980 2034
rect 3798 2033 3804 2034
rect 1974 2029 1975 2033
rect 1979 2029 1980 2033
rect 1974 2028 1980 2029
rect 2022 2032 2028 2033
rect 2278 2032 2284 2033
rect 2550 2032 2556 2033
rect 2798 2032 2804 2033
rect 3030 2032 3036 2033
rect 3254 2032 3260 2033
rect 3478 2032 3484 2033
rect 3678 2032 3684 2033
rect 2022 2028 2023 2032
rect 2027 2028 2028 2032
rect 2022 2027 2028 2028
rect 2118 2031 2125 2032
rect 2118 2027 2119 2031
rect 2124 2027 2125 2031
rect 2278 2028 2279 2032
rect 2283 2028 2284 2032
rect 2278 2027 2284 2028
rect 2374 2031 2381 2032
rect 2374 2027 2375 2031
rect 2380 2027 2381 2031
rect 2550 2028 2551 2032
rect 2555 2028 2556 2032
rect 2550 2027 2556 2028
rect 2646 2031 2653 2032
rect 2646 2027 2647 2031
rect 2652 2027 2653 2031
rect 2798 2028 2799 2032
rect 2803 2028 2804 2032
rect 2798 2027 2804 2028
rect 2890 2031 2901 2032
rect 2890 2027 2891 2031
rect 2895 2027 2896 2031
rect 2900 2027 2901 2031
rect 3030 2028 3031 2032
rect 3035 2028 3036 2032
rect 3030 2027 3036 2028
rect 3122 2031 3133 2032
rect 3122 2027 3123 2031
rect 3127 2027 3128 2031
rect 3132 2027 3133 2031
rect 3254 2028 3255 2032
rect 3259 2028 3260 2032
rect 3254 2027 3260 2028
rect 3350 2031 3357 2032
rect 3350 2027 3351 2031
rect 3356 2027 3357 2031
rect 3478 2028 3479 2032
rect 3483 2028 3484 2032
rect 3478 2027 3484 2028
rect 3575 2031 3584 2032
rect 3575 2027 3576 2031
rect 3583 2027 3584 2031
rect 3678 2028 3679 2032
rect 3683 2028 3684 2032
rect 3678 2027 3684 2028
rect 3770 2031 3781 2032
rect 3770 2027 3771 2031
rect 3775 2027 3776 2031
rect 3780 2027 3781 2031
rect 3798 2029 3799 2033
rect 3803 2029 3804 2033
rect 3798 2028 3804 2029
rect 2118 2026 2125 2027
rect 2374 2026 2381 2027
rect 2646 2026 2653 2027
rect 2890 2026 2901 2027
rect 3122 2026 3133 2027
rect 3350 2026 3357 2027
rect 3575 2026 3584 2027
rect 3770 2026 3781 2027
rect 110 2025 116 2026
rect 1934 2025 1940 2026
rect 110 2021 111 2025
rect 115 2021 116 2025
rect 110 2020 116 2021
rect 222 2024 228 2025
rect 382 2024 388 2025
rect 558 2024 564 2025
rect 750 2024 756 2025
rect 958 2024 964 2025
rect 1166 2024 1172 2025
rect 1382 2024 1388 2025
rect 1606 2024 1612 2025
rect 1814 2024 1820 2025
rect 222 2020 223 2024
rect 227 2020 228 2024
rect 222 2019 228 2020
rect 319 2023 328 2024
rect 319 2019 320 2023
rect 327 2019 328 2023
rect 382 2020 383 2024
rect 387 2020 388 2024
rect 382 2019 388 2020
rect 479 2023 485 2024
rect 479 2019 480 2023
rect 484 2022 485 2023
rect 495 2023 501 2024
rect 495 2022 496 2023
rect 484 2020 496 2022
rect 484 2019 485 2020
rect 319 2018 328 2019
rect 479 2018 485 2019
rect 495 2019 496 2020
rect 500 2019 501 2023
rect 558 2020 559 2024
rect 563 2020 564 2024
rect 558 2019 564 2020
rect 655 2023 661 2024
rect 655 2019 656 2023
rect 660 2022 661 2023
rect 738 2023 744 2024
rect 738 2022 739 2023
rect 660 2020 739 2022
rect 660 2019 661 2020
rect 495 2018 501 2019
rect 655 2018 661 2019
rect 738 2019 739 2020
rect 743 2019 744 2023
rect 750 2020 751 2024
rect 755 2020 756 2024
rect 750 2019 756 2020
rect 842 2023 853 2024
rect 842 2019 843 2023
rect 847 2019 848 2023
rect 852 2019 853 2023
rect 958 2020 959 2024
rect 963 2020 964 2024
rect 958 2019 964 2020
rect 1054 2023 1061 2024
rect 1054 2019 1055 2023
rect 1060 2019 1061 2023
rect 1166 2020 1167 2024
rect 1171 2020 1172 2024
rect 1166 2019 1172 2020
rect 1258 2023 1269 2024
rect 1258 2019 1259 2023
rect 1263 2019 1264 2023
rect 1268 2019 1269 2023
rect 1382 2020 1383 2024
rect 1387 2020 1388 2024
rect 1382 2019 1388 2020
rect 1479 2023 1488 2024
rect 1479 2019 1480 2023
rect 1487 2019 1488 2023
rect 1606 2020 1607 2024
rect 1611 2020 1612 2024
rect 1606 2019 1612 2020
rect 1702 2023 1709 2024
rect 1702 2019 1703 2023
rect 1708 2019 1709 2023
rect 1814 2020 1815 2024
rect 1819 2020 1820 2024
rect 1814 2019 1820 2020
rect 1911 2023 1917 2024
rect 1911 2019 1912 2023
rect 1916 2019 1917 2023
rect 1934 2021 1935 2025
rect 1939 2021 1940 2025
rect 1934 2020 1940 2021
rect 738 2018 744 2019
rect 842 2018 853 2019
rect 1054 2018 1061 2019
rect 1258 2018 1269 2019
rect 1479 2018 1488 2019
rect 1702 2018 1709 2019
rect 1911 2018 1917 2019
rect 194 2009 200 2010
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 194 2005 195 2009
rect 199 2005 200 2009
rect 194 2004 200 2005
rect 354 2009 360 2010
rect 354 2005 355 2009
rect 359 2005 360 2009
rect 354 2004 360 2005
rect 530 2009 536 2010
rect 530 2005 531 2009
rect 535 2005 536 2009
rect 530 2004 536 2005
rect 722 2009 728 2010
rect 722 2005 723 2009
rect 727 2005 728 2009
rect 722 2004 728 2005
rect 930 2009 936 2010
rect 930 2005 931 2009
rect 935 2005 936 2009
rect 930 2004 936 2005
rect 1138 2009 1144 2010
rect 1138 2005 1139 2009
rect 1143 2005 1144 2009
rect 1138 2004 1144 2005
rect 1354 2009 1360 2010
rect 1354 2005 1355 2009
rect 1359 2005 1360 2009
rect 1354 2004 1360 2005
rect 1578 2009 1584 2010
rect 1578 2005 1579 2009
rect 1583 2005 1584 2009
rect 1578 2004 1584 2005
rect 1786 2009 1792 2010
rect 1786 2005 1787 2009
rect 1791 2005 1792 2009
rect 1786 2004 1792 2005
rect 110 2003 116 2004
rect 1234 2003 1240 2004
rect 1234 1999 1235 2003
rect 1239 2002 1240 2003
rect 1566 2003 1572 2004
rect 1566 2002 1567 2003
rect 1239 2000 1567 2002
rect 1239 1999 1240 2000
rect 1234 1998 1240 1999
rect 1566 1999 1567 2000
rect 1571 1999 1572 2003
rect 1566 1998 1572 1999
rect 1674 2003 1680 2004
rect 1674 1999 1675 2003
rect 1679 2002 1680 2003
rect 1912 2002 1914 2018
rect 1994 2017 2000 2018
rect 1974 2016 1980 2017
rect 1974 2012 1975 2016
rect 1979 2012 1980 2016
rect 1994 2013 1995 2017
rect 1999 2013 2000 2017
rect 1994 2012 2000 2013
rect 2250 2017 2256 2018
rect 2250 2013 2251 2017
rect 2255 2013 2256 2017
rect 2250 2012 2256 2013
rect 2522 2017 2528 2018
rect 2522 2013 2523 2017
rect 2527 2013 2528 2017
rect 2522 2012 2528 2013
rect 2770 2017 2776 2018
rect 2770 2013 2771 2017
rect 2775 2013 2776 2017
rect 2770 2012 2776 2013
rect 3002 2017 3008 2018
rect 3002 2013 3003 2017
rect 3007 2013 3008 2017
rect 3002 2012 3008 2013
rect 3226 2017 3232 2018
rect 3226 2013 3227 2017
rect 3231 2013 3232 2017
rect 3226 2012 3232 2013
rect 3450 2017 3456 2018
rect 3450 2013 3451 2017
rect 3455 2013 3456 2017
rect 3450 2012 3456 2013
rect 3650 2017 3656 2018
rect 3650 2013 3651 2017
rect 3655 2013 3656 2017
rect 3650 2012 3656 2013
rect 3798 2016 3804 2017
rect 3798 2012 3799 2016
rect 3803 2012 3804 2016
rect 1974 2011 1980 2012
rect 3798 2011 3804 2012
rect 1934 2008 1940 2009
rect 1934 2004 1935 2008
rect 1939 2004 1940 2008
rect 1934 2003 1940 2004
rect 2866 2003 2872 2004
rect 1679 2000 1914 2002
rect 1679 1999 1680 2000
rect 1674 1998 1680 1999
rect 2866 1999 2867 2003
rect 2871 2002 2872 2003
rect 3122 2003 3128 2004
rect 3122 2002 3123 2003
rect 2871 2000 3123 2002
rect 2871 1999 2872 2000
rect 2866 1998 2872 1999
rect 3122 1999 3123 2000
rect 3127 1999 3128 2003
rect 3122 1998 3128 1999
rect 3546 1999 3552 2000
rect 3546 1995 3547 1999
rect 3551 1998 3552 1999
rect 3770 1999 3776 2000
rect 3770 1998 3771 1999
rect 3551 1996 3771 1998
rect 3551 1995 3552 1996
rect 3546 1994 3552 1995
rect 3770 1995 3771 1996
rect 3775 1995 3776 1999
rect 3770 1994 3776 1995
rect 3838 1989 3844 1990
rect 5662 1989 5668 1990
rect 1026 1987 1032 1988
rect 1026 1983 1027 1987
rect 1031 1986 1032 1987
rect 1258 1987 1264 1988
rect 1258 1986 1259 1987
rect 1031 1984 1259 1986
rect 1031 1983 1032 1984
rect 1026 1982 1032 1983
rect 1258 1983 1259 1984
rect 1263 1983 1264 1987
rect 3838 1985 3839 1989
rect 3843 1985 3844 1989
rect 3838 1984 3844 1985
rect 4726 1988 4732 1989
rect 4862 1988 4868 1989
rect 5006 1988 5012 1989
rect 5158 1988 5164 1989
rect 5318 1988 5324 1989
rect 5486 1988 5492 1989
rect 4726 1984 4727 1988
rect 4731 1984 4732 1988
rect 4726 1983 4732 1984
rect 4823 1987 4832 1988
rect 4823 1983 4824 1987
rect 4831 1983 4832 1987
rect 4862 1984 4863 1988
rect 4867 1984 4868 1988
rect 4862 1983 4868 1984
rect 4959 1987 4965 1988
rect 4959 1983 4960 1987
rect 4964 1986 4965 1987
rect 4970 1987 4976 1988
rect 4970 1986 4971 1987
rect 4964 1984 4971 1986
rect 4964 1983 4965 1984
rect 1258 1982 1264 1983
rect 4823 1982 4832 1983
rect 4959 1982 4965 1983
rect 4970 1983 4971 1984
rect 4975 1983 4976 1987
rect 5006 1984 5007 1988
rect 5011 1984 5012 1988
rect 5006 1983 5012 1984
rect 5103 1987 5109 1988
rect 5103 1983 5104 1987
rect 5108 1986 5109 1987
rect 5119 1987 5125 1988
rect 5119 1986 5120 1987
rect 5108 1984 5120 1986
rect 5108 1983 5109 1984
rect 4970 1982 4976 1983
rect 5103 1982 5109 1983
rect 5119 1983 5120 1984
rect 5124 1983 5125 1987
rect 5158 1984 5159 1988
rect 5163 1984 5164 1988
rect 5158 1983 5164 1984
rect 5250 1987 5261 1988
rect 5250 1983 5251 1987
rect 5255 1983 5256 1987
rect 5260 1983 5261 1987
rect 5318 1984 5319 1988
rect 5323 1984 5324 1988
rect 5318 1983 5324 1984
rect 5410 1987 5421 1988
rect 5410 1983 5411 1987
rect 5415 1983 5416 1987
rect 5420 1983 5421 1987
rect 5486 1984 5487 1988
rect 5491 1984 5492 1988
rect 5486 1983 5492 1984
rect 5582 1987 5589 1988
rect 5582 1983 5583 1987
rect 5588 1983 5589 1987
rect 5662 1985 5663 1989
rect 5667 1985 5668 1989
rect 5662 1984 5668 1985
rect 5119 1982 5125 1983
rect 5250 1982 5261 1983
rect 5410 1982 5421 1983
rect 5582 1982 5589 1983
rect 4698 1973 4704 1974
rect 3838 1972 3844 1973
rect 3838 1968 3839 1972
rect 3843 1968 3844 1972
rect 4698 1969 4699 1973
rect 4703 1969 4704 1973
rect 4698 1968 4704 1969
rect 4834 1973 4840 1974
rect 4834 1969 4835 1973
rect 4839 1969 4840 1973
rect 4834 1968 4840 1969
rect 4978 1973 4984 1974
rect 4978 1969 4979 1973
rect 4983 1969 4984 1973
rect 4978 1968 4984 1969
rect 5130 1973 5136 1974
rect 5130 1969 5131 1973
rect 5135 1969 5136 1973
rect 5130 1968 5136 1969
rect 5290 1973 5296 1974
rect 5290 1969 5291 1973
rect 5295 1969 5296 1973
rect 5290 1968 5296 1969
rect 5458 1973 5464 1974
rect 5458 1969 5459 1973
rect 5463 1969 5464 1973
rect 5458 1968 5464 1969
rect 5662 1972 5668 1973
rect 5662 1968 5663 1972
rect 5667 1968 5668 1972
rect 2442 1967 2448 1968
rect 314 1959 320 1960
rect 314 1958 315 1959
rect 293 1956 315 1958
rect 314 1955 315 1956
rect 319 1955 320 1959
rect 314 1954 320 1955
rect 322 1959 328 1960
rect 322 1955 323 1959
rect 327 1958 328 1959
rect 495 1959 501 1960
rect 327 1956 361 1958
rect 327 1955 328 1956
rect 322 1954 328 1955
rect 495 1955 496 1959
rect 500 1958 501 1959
rect 1026 1959 1032 1960
rect 500 1956 537 1958
rect 500 1955 501 1956
rect 495 1954 501 1955
rect 820 1950 822 1957
rect 1026 1955 1027 1959
rect 1031 1955 1032 1959
rect 1026 1954 1032 1955
rect 1234 1959 1240 1960
rect 1234 1955 1235 1959
rect 1239 1955 1240 1959
rect 1674 1959 1680 1960
rect 1234 1954 1240 1955
rect 1054 1951 1060 1952
rect 1054 1950 1055 1951
rect 820 1948 1055 1950
rect 1054 1947 1055 1948
rect 1059 1947 1060 1951
rect 1452 1950 1454 1957
rect 1674 1955 1675 1959
rect 1679 1955 1680 1959
rect 1910 1959 1916 1960
rect 1910 1958 1911 1959
rect 1885 1956 1911 1958
rect 1674 1954 1680 1955
rect 1910 1955 1911 1956
rect 1915 1955 1916 1959
rect 2092 1958 2094 1965
rect 2349 1964 2438 1966
rect 2374 1959 2380 1960
rect 2374 1958 2375 1959
rect 2092 1956 2375 1958
rect 1910 1954 1916 1955
rect 2374 1955 2375 1956
rect 2379 1955 2380 1959
rect 2436 1958 2438 1964
rect 2442 1963 2443 1967
rect 2447 1966 2448 1967
rect 2866 1967 2872 1968
rect 2447 1964 2529 1966
rect 2447 1963 2448 1964
rect 2442 1962 2448 1963
rect 2866 1963 2867 1967
rect 2871 1963 2872 1967
rect 3238 1967 3244 1968
rect 2866 1962 2872 1963
rect 2646 1959 2652 1960
rect 2646 1958 2647 1959
rect 2436 1956 2647 1958
rect 2374 1954 2380 1955
rect 2646 1955 2647 1956
rect 2651 1955 2652 1959
rect 3100 1958 3102 1965
rect 3238 1963 3239 1967
rect 3243 1963 3244 1967
rect 3238 1962 3244 1963
rect 3546 1967 3552 1968
rect 3546 1963 3547 1967
rect 3551 1963 3552 1967
rect 3770 1967 3776 1968
rect 3838 1967 3844 1968
rect 5662 1967 5668 1968
rect 3770 1966 3771 1967
rect 3749 1964 3771 1966
rect 3546 1962 3552 1963
rect 3770 1963 3771 1964
rect 3775 1963 3776 1967
rect 3770 1962 3776 1963
rect 3350 1959 3356 1960
rect 3350 1958 3351 1959
rect 3100 1956 3351 1958
rect 2646 1954 2652 1955
rect 3350 1955 3351 1956
rect 3355 1955 3356 1959
rect 3350 1954 3356 1955
rect 1702 1951 1708 1952
rect 1702 1950 1703 1951
rect 1452 1948 1703 1950
rect 1054 1946 1060 1947
rect 1702 1947 1703 1948
rect 1707 1947 1708 1951
rect 1702 1946 1708 1947
rect 842 1927 848 1928
rect 842 1926 843 1927
rect 816 1924 843 1926
rect 506 1923 512 1924
rect 506 1922 507 1923
rect 384 1920 507 1922
rect 384 1918 386 1920
rect 506 1919 507 1920
rect 511 1919 512 1923
rect 506 1918 512 1919
rect 816 1918 818 1924
rect 842 1923 843 1924
rect 847 1923 848 1927
rect 842 1922 848 1923
rect 2206 1923 2212 1924
rect 2206 1922 2207 1923
rect 2093 1920 2207 1922
rect 1474 1919 1480 1920
rect 1474 1918 1475 1919
rect 293 1916 386 1918
rect 693 1916 818 1918
rect 1381 1916 1475 1918
rect 826 1915 832 1916
rect 480 1910 482 1913
rect 574 1911 580 1912
rect 574 1910 575 1911
rect 480 1908 575 1910
rect 574 1907 575 1908
rect 579 1907 580 1911
rect 826 1911 827 1915
rect 831 1911 832 1915
rect 826 1910 832 1911
rect 1058 1915 1064 1916
rect 1058 1911 1059 1915
rect 1063 1911 1064 1915
rect 1474 1915 1475 1916
rect 1479 1915 1480 1919
rect 1474 1914 1480 1915
rect 1482 1919 1488 1920
rect 1482 1915 1483 1919
rect 1487 1918 1488 1919
rect 2206 1919 2207 1920
rect 2211 1919 2212 1923
rect 2890 1923 2896 1924
rect 2890 1922 2891 1923
rect 2717 1920 2891 1922
rect 2206 1918 2212 1919
rect 2322 1919 2328 1920
rect 1487 1916 1529 1918
rect 1487 1915 1488 1916
rect 1482 1914 1488 1915
rect 1778 1915 1784 1916
rect 1058 1910 1064 1911
rect 1778 1911 1779 1915
rect 1783 1911 1784 1915
rect 2322 1915 2323 1919
rect 2327 1915 2328 1919
rect 2890 1919 2891 1920
rect 2895 1919 2896 1923
rect 3534 1923 3540 1924
rect 3534 1922 3535 1923
rect 3517 1920 3535 1922
rect 2890 1918 2896 1919
rect 2906 1919 2912 1920
rect 2322 1914 2328 1915
rect 2906 1915 2907 1919
rect 2911 1915 2912 1919
rect 2906 1914 2912 1915
rect 3170 1919 3176 1920
rect 3170 1915 3171 1919
rect 3175 1915 3176 1919
rect 3534 1919 3535 1920
rect 3539 1919 3540 1923
rect 4826 1923 4832 1924
rect 3534 1918 3540 1919
rect 3658 1919 3664 1920
rect 3170 1914 3176 1915
rect 3658 1915 3659 1919
rect 3663 1915 3664 1919
rect 3658 1914 3664 1915
rect 4796 1914 4798 1921
rect 4826 1919 4827 1923
rect 4831 1922 4832 1923
rect 5074 1923 5080 1924
rect 4831 1920 4841 1922
rect 4831 1919 4832 1920
rect 4826 1918 4832 1919
rect 5074 1919 5075 1923
rect 5079 1919 5080 1923
rect 5074 1918 5080 1919
rect 5119 1923 5125 1924
rect 5119 1919 5120 1923
rect 5124 1922 5125 1923
rect 5358 1923 5364 1924
rect 5124 1920 5137 1922
rect 5124 1919 5125 1920
rect 5119 1918 5125 1919
rect 5358 1919 5359 1923
rect 5363 1919 5364 1923
rect 5646 1923 5652 1924
rect 5646 1922 5647 1923
rect 5557 1920 5647 1922
rect 5358 1918 5364 1919
rect 5646 1919 5647 1920
rect 5651 1919 5652 1923
rect 5646 1918 5652 1919
rect 5250 1915 5256 1916
rect 5250 1914 5251 1915
rect 4796 1912 5251 1914
rect 1778 1910 1784 1911
rect 5250 1911 5251 1912
rect 5255 1911 5256 1915
rect 5250 1910 5256 1911
rect 574 1906 580 1907
rect 4490 1891 4496 1892
rect 4490 1890 4491 1891
rect 4373 1888 4491 1890
rect 4490 1887 4491 1888
rect 4495 1887 4496 1891
rect 4970 1891 4976 1892
rect 4490 1886 4496 1887
rect 4506 1887 4512 1888
rect 4506 1883 4507 1887
rect 4511 1883 4512 1887
rect 4506 1882 4512 1883
rect 4738 1887 4744 1888
rect 4738 1883 4739 1887
rect 4743 1883 4744 1887
rect 4970 1887 4971 1891
rect 4975 1890 4976 1891
rect 5338 1891 5344 1892
rect 5338 1890 5339 1891
rect 4975 1888 4985 1890
rect 5333 1888 5339 1890
rect 4975 1887 4976 1888
rect 4970 1886 4976 1887
rect 5338 1887 5339 1888
rect 5343 1887 5344 1891
rect 5338 1886 5344 1887
rect 5582 1891 5588 1892
rect 5582 1887 5583 1891
rect 5587 1887 5588 1891
rect 5582 1886 5588 1887
rect 4738 1882 4744 1883
rect 1974 1872 1980 1873
rect 3798 1872 3804 1873
rect 110 1868 116 1869
rect 1934 1868 1940 1869
rect 110 1864 111 1868
rect 115 1864 116 1868
rect 110 1863 116 1864
rect 194 1867 200 1868
rect 194 1863 195 1867
rect 199 1863 200 1867
rect 194 1862 200 1863
rect 386 1867 392 1868
rect 386 1863 387 1867
rect 391 1863 392 1867
rect 386 1862 392 1863
rect 594 1867 600 1868
rect 594 1863 595 1867
rect 599 1863 600 1867
rect 594 1862 600 1863
rect 818 1867 824 1868
rect 818 1863 819 1867
rect 823 1863 824 1867
rect 818 1862 824 1863
rect 1050 1867 1056 1868
rect 1050 1863 1051 1867
rect 1055 1863 1056 1867
rect 1050 1862 1056 1863
rect 1282 1867 1288 1868
rect 1282 1863 1283 1867
rect 1287 1863 1288 1867
rect 1282 1862 1288 1863
rect 1522 1867 1528 1868
rect 1522 1863 1523 1867
rect 1527 1863 1528 1867
rect 1522 1862 1528 1863
rect 1770 1867 1776 1868
rect 1770 1863 1771 1867
rect 1775 1863 1776 1867
rect 1934 1864 1935 1868
rect 1939 1864 1940 1868
rect 1974 1868 1975 1872
rect 1979 1868 1980 1872
rect 1974 1867 1980 1868
rect 1994 1871 2000 1872
rect 1994 1867 1995 1871
rect 1999 1867 2000 1871
rect 1994 1866 2000 1867
rect 2314 1871 2320 1872
rect 2314 1867 2315 1871
rect 2319 1867 2320 1871
rect 2314 1866 2320 1867
rect 2618 1871 2624 1872
rect 2618 1867 2619 1871
rect 2623 1867 2624 1871
rect 2618 1866 2624 1867
rect 2898 1871 2904 1872
rect 2898 1867 2899 1871
rect 2903 1867 2904 1871
rect 2898 1866 2904 1867
rect 3162 1871 3168 1872
rect 3162 1867 3163 1871
rect 3167 1867 3168 1871
rect 3162 1866 3168 1867
rect 3418 1871 3424 1872
rect 3418 1867 3419 1871
rect 3423 1867 3424 1871
rect 3418 1866 3424 1867
rect 3650 1871 3656 1872
rect 3650 1867 3651 1871
rect 3655 1867 3656 1871
rect 3798 1868 3799 1872
rect 3803 1868 3804 1872
rect 3798 1867 3804 1868
rect 3650 1866 3656 1867
rect 1934 1863 1940 1864
rect 1770 1862 1776 1863
rect 1474 1859 1480 1860
rect 1474 1855 1475 1859
rect 1479 1858 1480 1859
rect 1479 1856 1898 1858
rect 2022 1856 2028 1857
rect 2342 1856 2348 1857
rect 2646 1856 2652 1857
rect 2926 1856 2932 1857
rect 3190 1856 3196 1857
rect 3446 1856 3452 1857
rect 3678 1856 3684 1857
rect 1479 1855 1480 1856
rect 1474 1854 1480 1855
rect 1896 1854 1898 1856
rect 1974 1855 1980 1856
rect 1895 1853 1901 1854
rect 222 1852 228 1853
rect 414 1852 420 1853
rect 622 1852 628 1853
rect 846 1852 852 1853
rect 1078 1852 1084 1853
rect 1310 1852 1316 1853
rect 1550 1852 1556 1853
rect 1798 1852 1804 1853
rect 110 1851 116 1852
rect 110 1847 111 1851
rect 115 1847 116 1851
rect 222 1848 223 1852
rect 227 1848 228 1852
rect 222 1847 228 1848
rect 314 1851 325 1852
rect 314 1847 315 1851
rect 319 1847 320 1851
rect 324 1847 325 1851
rect 414 1848 415 1852
rect 419 1848 420 1852
rect 414 1847 420 1848
rect 506 1851 517 1852
rect 506 1847 507 1851
rect 511 1847 512 1851
rect 516 1847 517 1851
rect 622 1848 623 1852
rect 627 1848 628 1852
rect 622 1847 628 1848
rect 719 1851 725 1852
rect 719 1847 720 1851
rect 724 1850 725 1851
rect 826 1851 832 1852
rect 826 1850 827 1851
rect 724 1848 827 1850
rect 724 1847 725 1848
rect 110 1846 116 1847
rect 314 1846 325 1847
rect 506 1846 517 1847
rect 719 1846 725 1847
rect 826 1847 827 1848
rect 831 1847 832 1851
rect 846 1848 847 1852
rect 851 1848 852 1852
rect 846 1847 852 1848
rect 943 1851 949 1852
rect 943 1847 944 1851
rect 948 1850 949 1851
rect 1058 1851 1064 1852
rect 1058 1850 1059 1851
rect 948 1848 1059 1850
rect 948 1847 949 1848
rect 826 1846 832 1847
rect 943 1846 949 1847
rect 1058 1847 1059 1848
rect 1063 1847 1064 1851
rect 1078 1848 1079 1852
rect 1083 1848 1084 1852
rect 1078 1847 1084 1848
rect 1170 1851 1181 1852
rect 1170 1847 1171 1851
rect 1175 1847 1176 1851
rect 1180 1847 1181 1851
rect 1310 1848 1311 1852
rect 1315 1848 1316 1852
rect 1310 1847 1316 1848
rect 1406 1851 1413 1852
rect 1406 1847 1407 1851
rect 1412 1847 1413 1851
rect 1550 1848 1551 1852
rect 1555 1848 1556 1852
rect 1550 1847 1556 1848
rect 1647 1851 1653 1852
rect 1647 1847 1648 1851
rect 1652 1850 1653 1851
rect 1778 1851 1784 1852
rect 1778 1850 1779 1851
rect 1652 1848 1779 1850
rect 1652 1847 1653 1848
rect 1058 1846 1064 1847
rect 1170 1846 1181 1847
rect 1406 1846 1413 1847
rect 1647 1846 1653 1847
rect 1778 1847 1779 1848
rect 1783 1847 1784 1851
rect 1798 1848 1799 1852
rect 1803 1848 1804 1852
rect 1895 1849 1896 1853
rect 1900 1849 1901 1853
rect 1895 1848 1901 1849
rect 1934 1851 1940 1852
rect 1798 1847 1804 1848
rect 1934 1847 1935 1851
rect 1939 1847 1940 1851
rect 1974 1851 1975 1855
rect 1979 1851 1980 1855
rect 2022 1852 2023 1856
rect 2027 1852 2028 1856
rect 2022 1851 2028 1852
rect 2119 1855 2125 1856
rect 2119 1851 2120 1855
rect 2124 1854 2125 1855
rect 2322 1855 2328 1856
rect 2322 1854 2323 1855
rect 2124 1852 2323 1854
rect 2124 1851 2125 1852
rect 1974 1850 1980 1851
rect 2119 1850 2125 1851
rect 2322 1851 2323 1852
rect 2327 1851 2328 1855
rect 2342 1852 2343 1856
rect 2347 1852 2348 1856
rect 2342 1851 2348 1852
rect 2439 1855 2448 1856
rect 2439 1851 2440 1855
rect 2447 1851 2448 1855
rect 2646 1852 2647 1856
rect 2651 1852 2652 1856
rect 2646 1851 2652 1852
rect 2743 1855 2749 1856
rect 2743 1851 2744 1855
rect 2748 1854 2749 1855
rect 2906 1855 2912 1856
rect 2906 1854 2907 1855
rect 2748 1852 2907 1854
rect 2748 1851 2749 1852
rect 2322 1850 2328 1851
rect 2439 1850 2448 1851
rect 2743 1850 2749 1851
rect 2906 1851 2907 1852
rect 2911 1851 2912 1855
rect 2926 1852 2927 1856
rect 2931 1852 2932 1856
rect 2926 1851 2932 1852
rect 3023 1855 3029 1856
rect 3023 1851 3024 1855
rect 3028 1854 3029 1855
rect 3170 1855 3176 1856
rect 3170 1854 3171 1855
rect 3028 1852 3171 1854
rect 3028 1851 3029 1852
rect 2906 1850 2912 1851
rect 3023 1850 3029 1851
rect 3170 1851 3171 1852
rect 3175 1851 3176 1855
rect 3190 1852 3191 1856
rect 3195 1852 3196 1856
rect 3190 1851 3196 1852
rect 3286 1855 3293 1856
rect 3286 1851 3287 1855
rect 3292 1851 3293 1855
rect 3446 1852 3447 1856
rect 3451 1852 3452 1856
rect 3446 1851 3452 1852
rect 3543 1855 3549 1856
rect 3543 1851 3544 1855
rect 3548 1854 3549 1855
rect 3658 1855 3664 1856
rect 3658 1854 3659 1855
rect 3548 1852 3659 1854
rect 3548 1851 3549 1852
rect 3170 1850 3176 1851
rect 3286 1850 3293 1851
rect 3543 1850 3549 1851
rect 3658 1851 3659 1852
rect 3663 1851 3664 1855
rect 3678 1852 3679 1856
rect 3683 1852 3684 1856
rect 3678 1851 3684 1852
rect 3770 1855 3781 1856
rect 3770 1851 3771 1855
rect 3775 1851 3776 1855
rect 3780 1851 3781 1855
rect 3658 1850 3664 1851
rect 3770 1850 3781 1851
rect 3798 1855 3804 1856
rect 3798 1851 3799 1855
rect 3803 1851 3804 1855
rect 3798 1850 3804 1851
rect 1778 1846 1784 1847
rect 1934 1846 1940 1847
rect 3838 1840 3844 1841
rect 5662 1840 5668 1841
rect 3838 1836 3839 1840
rect 3843 1836 3844 1840
rect 3838 1835 3844 1836
rect 4274 1839 4280 1840
rect 4274 1835 4275 1839
rect 4279 1835 4280 1839
rect 4274 1834 4280 1835
rect 4498 1839 4504 1840
rect 4498 1835 4499 1839
rect 4503 1835 4504 1839
rect 4498 1834 4504 1835
rect 4730 1839 4736 1840
rect 4730 1835 4731 1839
rect 4735 1835 4736 1839
rect 4730 1834 4736 1835
rect 4978 1839 4984 1840
rect 4978 1835 4979 1839
rect 4983 1835 4984 1839
rect 4978 1834 4984 1835
rect 5234 1839 5240 1840
rect 5234 1835 5235 1839
rect 5239 1835 5240 1839
rect 5234 1834 5240 1835
rect 5498 1839 5504 1840
rect 5498 1835 5499 1839
rect 5503 1835 5504 1839
rect 5662 1836 5663 1840
rect 5667 1836 5668 1840
rect 5662 1835 5668 1836
rect 5498 1834 5504 1835
rect 4490 1831 4496 1832
rect 4490 1827 4491 1831
rect 4495 1830 4496 1831
rect 4495 1828 5106 1830
rect 4495 1827 4496 1828
rect 4490 1826 4496 1827
rect 5104 1826 5106 1828
rect 5103 1825 5109 1826
rect 4302 1824 4308 1825
rect 4526 1824 4532 1825
rect 4758 1824 4764 1825
rect 5006 1824 5012 1825
rect 3838 1823 3844 1824
rect 3838 1819 3839 1823
rect 3843 1819 3844 1823
rect 4302 1820 4303 1824
rect 4307 1820 4308 1824
rect 4302 1819 4308 1820
rect 4399 1823 4405 1824
rect 4399 1819 4400 1823
rect 4404 1822 4405 1823
rect 4506 1823 4512 1824
rect 4506 1822 4507 1823
rect 4404 1820 4507 1822
rect 4404 1819 4405 1820
rect 3838 1818 3844 1819
rect 4399 1818 4405 1819
rect 4506 1819 4507 1820
rect 4511 1819 4512 1823
rect 4526 1820 4527 1824
rect 4531 1820 4532 1824
rect 4526 1819 4532 1820
rect 4623 1823 4629 1824
rect 4623 1819 4624 1823
rect 4628 1822 4629 1823
rect 4738 1823 4744 1824
rect 4738 1822 4739 1823
rect 4628 1820 4739 1822
rect 4628 1819 4629 1820
rect 4506 1818 4512 1819
rect 4623 1818 4629 1819
rect 4738 1819 4739 1820
rect 4743 1819 4744 1823
rect 4758 1820 4759 1824
rect 4763 1820 4764 1824
rect 4758 1819 4764 1820
rect 4855 1823 4864 1824
rect 4855 1819 4856 1823
rect 4863 1819 4864 1823
rect 5006 1820 5007 1824
rect 5011 1820 5012 1824
rect 5103 1821 5104 1825
rect 5108 1821 5109 1825
rect 5103 1820 5109 1821
rect 5262 1824 5268 1825
rect 5526 1824 5532 1825
rect 5262 1820 5263 1824
rect 5267 1820 5268 1824
rect 5006 1819 5012 1820
rect 5262 1819 5268 1820
rect 5358 1823 5365 1824
rect 5358 1819 5359 1823
rect 5364 1819 5365 1823
rect 5526 1820 5527 1824
rect 5531 1820 5532 1824
rect 5526 1819 5532 1820
rect 5622 1823 5629 1824
rect 5622 1819 5623 1823
rect 5628 1819 5629 1823
rect 4738 1818 4744 1819
rect 4855 1818 4864 1819
rect 5358 1818 5365 1819
rect 5622 1818 5629 1819
rect 5662 1823 5668 1824
rect 5662 1819 5663 1823
rect 5667 1819 5668 1823
rect 5662 1818 5668 1819
rect 1974 1793 1980 1794
rect 3798 1793 3804 1794
rect 1974 1789 1975 1793
rect 1979 1789 1980 1793
rect 1974 1788 1980 1789
rect 2110 1792 2116 1793
rect 2390 1792 2396 1793
rect 2662 1792 2668 1793
rect 2926 1792 2932 1793
rect 3182 1792 3188 1793
rect 3438 1792 3444 1793
rect 3678 1792 3684 1793
rect 2110 1788 2111 1792
rect 2115 1788 2116 1792
rect 2110 1787 2116 1788
rect 2206 1791 2213 1792
rect 2206 1787 2207 1791
rect 2212 1787 2213 1791
rect 2390 1788 2391 1792
rect 2395 1788 2396 1792
rect 2390 1787 2396 1788
rect 2486 1791 2493 1792
rect 2486 1787 2487 1791
rect 2492 1787 2493 1791
rect 2662 1788 2663 1792
rect 2667 1788 2668 1792
rect 2662 1787 2668 1788
rect 2754 1791 2765 1792
rect 2754 1787 2755 1791
rect 2759 1787 2760 1791
rect 2764 1787 2765 1791
rect 2926 1788 2927 1792
rect 2931 1788 2932 1792
rect 2926 1787 2932 1788
rect 3018 1791 3029 1792
rect 3018 1787 3019 1791
rect 3023 1787 3024 1791
rect 3028 1787 3029 1791
rect 3182 1788 3183 1792
rect 3187 1788 3188 1792
rect 3182 1787 3188 1788
rect 3278 1791 3285 1792
rect 3278 1787 3279 1791
rect 3284 1787 3285 1791
rect 3438 1788 3439 1792
rect 3443 1788 3444 1792
rect 3438 1787 3444 1788
rect 3534 1791 3541 1792
rect 3534 1787 3535 1791
rect 3540 1787 3541 1791
rect 3678 1788 3679 1792
rect 3683 1788 3684 1792
rect 3678 1787 3684 1788
rect 3770 1791 3781 1792
rect 3770 1787 3771 1791
rect 3775 1787 3776 1791
rect 3780 1787 3781 1791
rect 3798 1789 3799 1793
rect 3803 1789 3804 1793
rect 3798 1788 3804 1789
rect 2206 1786 2213 1787
rect 2486 1786 2493 1787
rect 2754 1786 2765 1787
rect 3018 1786 3029 1787
rect 3278 1786 3285 1787
rect 3534 1786 3541 1787
rect 3770 1786 3781 1787
rect 110 1777 116 1778
rect 1934 1777 1940 1778
rect 2082 1777 2088 1778
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 110 1772 116 1773
rect 158 1776 164 1777
rect 302 1776 308 1777
rect 478 1776 484 1777
rect 654 1776 660 1777
rect 830 1776 836 1777
rect 1006 1776 1012 1777
rect 1182 1776 1188 1777
rect 1358 1776 1364 1777
rect 1534 1776 1540 1777
rect 1710 1776 1716 1777
rect 158 1772 159 1776
rect 163 1772 164 1776
rect 158 1771 164 1772
rect 255 1775 261 1776
rect 255 1771 256 1775
rect 260 1774 261 1775
rect 266 1775 272 1776
rect 266 1774 267 1775
rect 260 1772 267 1774
rect 260 1771 261 1772
rect 255 1770 261 1771
rect 266 1771 267 1772
rect 271 1771 272 1775
rect 302 1772 303 1776
rect 307 1772 308 1776
rect 302 1771 308 1772
rect 399 1775 405 1776
rect 399 1771 400 1775
rect 404 1774 405 1775
rect 418 1775 424 1776
rect 418 1774 419 1775
rect 404 1772 419 1774
rect 404 1771 405 1772
rect 266 1770 272 1771
rect 399 1770 405 1771
rect 418 1771 419 1772
rect 423 1771 424 1775
rect 478 1772 479 1776
rect 483 1772 484 1776
rect 478 1771 484 1772
rect 574 1775 581 1776
rect 574 1771 575 1775
rect 580 1771 581 1775
rect 654 1772 655 1776
rect 659 1772 660 1776
rect 654 1771 660 1772
rect 751 1775 757 1776
rect 751 1771 752 1775
rect 756 1774 757 1775
rect 770 1775 776 1776
rect 770 1774 771 1775
rect 756 1772 771 1774
rect 756 1771 757 1772
rect 418 1770 424 1771
rect 574 1770 581 1771
rect 751 1770 757 1771
rect 770 1771 771 1772
rect 775 1771 776 1775
rect 830 1772 831 1776
rect 835 1772 836 1776
rect 830 1771 836 1772
rect 926 1775 933 1776
rect 926 1771 927 1775
rect 932 1771 933 1775
rect 1006 1772 1007 1776
rect 1011 1772 1012 1776
rect 1006 1771 1012 1772
rect 1098 1775 1109 1776
rect 1098 1771 1099 1775
rect 1103 1771 1104 1775
rect 1108 1771 1109 1775
rect 1182 1772 1183 1776
rect 1187 1772 1188 1776
rect 1182 1771 1188 1772
rect 1279 1775 1285 1776
rect 1279 1771 1280 1775
rect 1284 1774 1285 1775
rect 1290 1775 1296 1776
rect 1290 1774 1291 1775
rect 1284 1772 1291 1774
rect 1284 1771 1285 1772
rect 770 1770 776 1771
rect 926 1770 933 1771
rect 1098 1770 1109 1771
rect 1279 1770 1285 1771
rect 1290 1771 1291 1772
rect 1295 1771 1296 1775
rect 1358 1772 1359 1776
rect 1363 1772 1364 1776
rect 1358 1771 1364 1772
rect 1455 1775 1461 1776
rect 1455 1771 1456 1775
rect 1460 1774 1461 1775
rect 1470 1775 1476 1776
rect 1470 1774 1471 1775
rect 1460 1772 1471 1774
rect 1460 1771 1461 1772
rect 1290 1770 1296 1771
rect 1455 1770 1461 1771
rect 1470 1771 1471 1772
rect 1475 1771 1476 1775
rect 1534 1772 1535 1776
rect 1539 1772 1540 1776
rect 1534 1771 1540 1772
rect 1631 1775 1637 1776
rect 1631 1771 1632 1775
rect 1636 1774 1637 1775
rect 1646 1775 1652 1776
rect 1646 1774 1647 1775
rect 1636 1772 1647 1774
rect 1636 1771 1637 1772
rect 1470 1770 1476 1771
rect 1631 1770 1637 1771
rect 1646 1771 1647 1772
rect 1651 1771 1652 1775
rect 1710 1772 1711 1776
rect 1715 1772 1716 1776
rect 1710 1771 1716 1772
rect 1806 1775 1813 1776
rect 1806 1771 1807 1775
rect 1812 1771 1813 1775
rect 1934 1773 1935 1777
rect 1939 1773 1940 1777
rect 1934 1772 1940 1773
rect 1974 1776 1980 1777
rect 1974 1772 1975 1776
rect 1979 1772 1980 1776
rect 2082 1773 2083 1777
rect 2087 1773 2088 1777
rect 2082 1772 2088 1773
rect 2362 1777 2368 1778
rect 2362 1773 2363 1777
rect 2367 1773 2368 1777
rect 2362 1772 2368 1773
rect 2634 1777 2640 1778
rect 2634 1773 2635 1777
rect 2639 1773 2640 1777
rect 2634 1772 2640 1773
rect 2898 1777 2904 1778
rect 2898 1773 2899 1777
rect 2903 1773 2904 1777
rect 2898 1772 2904 1773
rect 3154 1777 3160 1778
rect 3154 1773 3155 1777
rect 3159 1773 3160 1777
rect 3154 1772 3160 1773
rect 3410 1777 3416 1778
rect 3410 1773 3411 1777
rect 3415 1773 3416 1777
rect 3410 1772 3416 1773
rect 3650 1777 3656 1778
rect 3650 1773 3651 1777
rect 3655 1773 3656 1777
rect 3650 1772 3656 1773
rect 3798 1776 3804 1777
rect 3798 1772 3799 1776
rect 3803 1772 3804 1776
rect 1974 1771 1980 1772
rect 3798 1771 3804 1772
rect 1646 1770 1652 1771
rect 1806 1770 1813 1771
rect 130 1761 136 1762
rect 110 1760 116 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 130 1757 131 1761
rect 135 1757 136 1761
rect 130 1756 136 1757
rect 274 1761 280 1762
rect 274 1757 275 1761
rect 279 1757 280 1761
rect 274 1756 280 1757
rect 450 1761 456 1762
rect 450 1757 451 1761
rect 455 1757 456 1761
rect 450 1756 456 1757
rect 626 1761 632 1762
rect 626 1757 627 1761
rect 631 1757 632 1761
rect 626 1756 632 1757
rect 802 1761 808 1762
rect 802 1757 803 1761
rect 807 1757 808 1761
rect 802 1756 808 1757
rect 978 1761 984 1762
rect 978 1757 979 1761
rect 983 1757 984 1761
rect 978 1756 984 1757
rect 1154 1761 1160 1762
rect 1154 1757 1155 1761
rect 1159 1757 1160 1761
rect 1154 1756 1160 1757
rect 1330 1761 1336 1762
rect 1330 1757 1331 1761
rect 1335 1757 1336 1761
rect 1330 1756 1336 1757
rect 1506 1761 1512 1762
rect 1506 1757 1507 1761
rect 1511 1757 1512 1761
rect 1506 1756 1512 1757
rect 1682 1761 1688 1762
rect 1682 1757 1683 1761
rect 1687 1757 1688 1761
rect 1682 1756 1688 1757
rect 1934 1760 1940 1761
rect 1934 1756 1935 1760
rect 1939 1756 1940 1760
rect 110 1755 116 1756
rect 1934 1755 1940 1756
rect 3838 1757 3844 1758
rect 5662 1757 5668 1758
rect 3838 1753 3839 1757
rect 3843 1753 3844 1757
rect 3838 1752 3844 1753
rect 3886 1756 3892 1757
rect 4086 1756 4092 1757
rect 4342 1756 4348 1757
rect 4622 1756 4628 1757
rect 4926 1756 4932 1757
rect 5246 1756 5252 1757
rect 5542 1756 5548 1757
rect 3886 1752 3887 1756
rect 3891 1752 3892 1756
rect 3886 1751 3892 1752
rect 3982 1755 3989 1756
rect 3982 1751 3983 1755
rect 3988 1751 3989 1755
rect 4086 1752 4087 1756
rect 4091 1752 4092 1756
rect 4086 1751 4092 1752
rect 4183 1755 4189 1756
rect 4183 1751 4184 1755
rect 4188 1754 4189 1755
rect 4222 1755 4228 1756
rect 4222 1754 4223 1755
rect 4188 1752 4223 1754
rect 4188 1751 4189 1752
rect 3982 1750 3989 1751
rect 4183 1750 4189 1751
rect 4222 1751 4223 1752
rect 4227 1751 4228 1755
rect 4342 1752 4343 1756
rect 4347 1752 4348 1756
rect 4342 1751 4348 1752
rect 4434 1755 4445 1756
rect 4434 1751 4435 1755
rect 4439 1751 4440 1755
rect 4444 1751 4445 1755
rect 4622 1752 4623 1756
rect 4627 1752 4628 1756
rect 4622 1751 4628 1752
rect 4714 1755 4725 1756
rect 4714 1751 4715 1755
rect 4719 1751 4720 1755
rect 4724 1751 4725 1755
rect 4926 1752 4927 1756
rect 4931 1752 4932 1756
rect 4926 1751 4932 1752
rect 5022 1755 5029 1756
rect 5022 1751 5023 1755
rect 5028 1751 5029 1755
rect 5246 1752 5247 1756
rect 5251 1752 5252 1756
rect 5246 1751 5252 1752
rect 5338 1755 5349 1756
rect 5338 1751 5339 1755
rect 5343 1751 5344 1755
rect 5348 1751 5349 1755
rect 5542 1752 5543 1756
rect 5547 1752 5548 1756
rect 5542 1751 5548 1752
rect 5634 1755 5645 1756
rect 5634 1751 5635 1755
rect 5639 1751 5640 1755
rect 5644 1751 5645 1755
rect 5662 1753 5663 1757
rect 5667 1753 5668 1757
rect 5662 1752 5668 1753
rect 4222 1750 4228 1751
rect 4434 1750 4445 1751
rect 4714 1750 4725 1751
rect 5022 1750 5029 1751
rect 5338 1750 5349 1751
rect 5634 1750 5645 1751
rect 3858 1741 3864 1742
rect 3838 1740 3844 1741
rect 722 1739 728 1740
rect 722 1735 723 1739
rect 727 1738 728 1739
rect 1098 1739 1104 1740
rect 1098 1738 1099 1739
rect 727 1736 1099 1738
rect 727 1735 728 1736
rect 722 1734 728 1735
rect 1098 1735 1099 1736
rect 1103 1735 1104 1739
rect 3838 1736 3839 1740
rect 3843 1736 3844 1740
rect 3858 1737 3859 1741
rect 3863 1737 3864 1741
rect 3858 1736 3864 1737
rect 4058 1741 4064 1742
rect 4058 1737 4059 1741
rect 4063 1737 4064 1741
rect 4058 1736 4064 1737
rect 4314 1741 4320 1742
rect 4314 1737 4315 1741
rect 4319 1737 4320 1741
rect 4314 1736 4320 1737
rect 4594 1741 4600 1742
rect 4594 1737 4595 1741
rect 4599 1737 4600 1741
rect 4594 1736 4600 1737
rect 4898 1741 4904 1742
rect 4898 1737 4899 1741
rect 4903 1737 4904 1741
rect 4898 1736 4904 1737
rect 5218 1741 5224 1742
rect 5218 1737 5219 1741
rect 5223 1737 5224 1741
rect 5218 1736 5224 1737
rect 5514 1741 5520 1742
rect 5514 1737 5515 1741
rect 5519 1737 5520 1741
rect 5514 1736 5520 1737
rect 5662 1740 5668 1741
rect 5662 1736 5663 1740
rect 5667 1736 5668 1740
rect 3838 1735 3844 1736
rect 5662 1735 5668 1736
rect 1098 1734 1104 1735
rect 2610 1727 2616 1728
rect 2610 1726 2611 1727
rect 2180 1718 2182 1725
rect 2461 1724 2611 1726
rect 2610 1723 2611 1724
rect 2615 1723 2616 1727
rect 3286 1727 3292 1728
rect 3286 1726 3287 1727
rect 2733 1724 2781 1726
rect 2997 1724 3158 1726
rect 3253 1724 3287 1726
rect 2610 1722 2616 1723
rect 2486 1719 2492 1720
rect 2486 1718 2487 1719
rect 2180 1716 2487 1718
rect 2486 1715 2487 1716
rect 2491 1715 2492 1719
rect 2779 1718 2781 1724
rect 3018 1719 3024 1720
rect 3018 1718 3019 1719
rect 2779 1716 3019 1718
rect 2486 1714 2492 1715
rect 3018 1715 3019 1716
rect 3023 1715 3024 1719
rect 3156 1718 3158 1724
rect 3286 1723 3287 1724
rect 3291 1723 3292 1727
rect 3982 1727 3988 1728
rect 3982 1726 3983 1727
rect 3509 1724 3621 1726
rect 3749 1724 3983 1726
rect 3286 1722 3292 1723
rect 3278 1719 3284 1720
rect 3278 1718 3279 1719
rect 3156 1716 3279 1718
rect 3018 1714 3024 1715
rect 3278 1715 3279 1716
rect 3283 1715 3284 1719
rect 3619 1718 3621 1724
rect 3982 1723 3983 1724
rect 3987 1723 3988 1727
rect 3982 1722 3988 1723
rect 3770 1719 3776 1720
rect 3770 1718 3771 1719
rect 3619 1716 3771 1718
rect 3278 1714 3284 1715
rect 3770 1715 3771 1716
rect 3775 1715 3776 1719
rect 3770 1714 3776 1715
rect 250 1711 256 1712
rect 250 1710 251 1711
rect 229 1708 251 1710
rect 250 1707 251 1708
rect 255 1707 256 1711
rect 250 1706 256 1707
rect 266 1711 272 1712
rect 266 1707 267 1711
rect 271 1710 272 1711
rect 418 1711 424 1712
rect 271 1708 281 1710
rect 271 1707 272 1708
rect 266 1706 272 1707
rect 418 1707 419 1711
rect 423 1710 424 1711
rect 722 1711 728 1712
rect 423 1708 457 1710
rect 423 1707 424 1708
rect 418 1706 424 1707
rect 722 1707 723 1711
rect 727 1707 728 1711
rect 722 1706 728 1707
rect 770 1711 776 1712
rect 770 1707 771 1711
rect 775 1710 776 1711
rect 1406 1711 1412 1712
rect 775 1708 809 1710
rect 1077 1708 1101 1710
rect 775 1707 776 1708
rect 770 1706 776 1707
rect 1099 1702 1101 1708
rect 1170 1703 1176 1704
rect 1170 1702 1171 1703
rect 1099 1700 1171 1702
rect 1170 1699 1171 1700
rect 1175 1699 1176 1703
rect 1252 1702 1254 1709
rect 1406 1707 1407 1711
rect 1411 1707 1412 1711
rect 1406 1706 1412 1707
rect 1470 1711 1476 1712
rect 1470 1707 1471 1711
rect 1475 1710 1476 1711
rect 1646 1711 1652 1712
rect 1475 1708 1513 1710
rect 1475 1707 1476 1708
rect 1470 1706 1476 1707
rect 1646 1707 1647 1711
rect 1651 1710 1652 1711
rect 1651 1708 1689 1710
rect 1651 1707 1652 1708
rect 1646 1706 1652 1707
rect 1806 1703 1812 1704
rect 1806 1702 1807 1703
rect 1252 1700 1807 1702
rect 1170 1698 1176 1699
rect 1806 1699 1807 1700
rect 1811 1699 1812 1703
rect 1806 1698 1812 1699
rect 3978 1691 3984 1692
rect 3978 1690 3979 1691
rect 3957 1688 3979 1690
rect 3978 1687 3979 1688
rect 3983 1687 3984 1691
rect 4222 1691 4228 1692
rect 3978 1686 3984 1687
rect 4156 1682 4158 1689
rect 4222 1687 4223 1691
rect 4227 1690 4228 1691
rect 4858 1691 4864 1692
rect 4227 1688 4321 1690
rect 4693 1688 4854 1690
rect 4227 1687 4228 1688
rect 4222 1686 4228 1687
rect 4714 1683 4720 1684
rect 4714 1682 4715 1683
rect 4156 1680 4715 1682
rect 1266 1679 1272 1680
rect 1266 1678 1267 1679
rect 1144 1676 1267 1678
rect 926 1675 932 1676
rect 926 1671 927 1675
rect 931 1671 932 1675
rect 1144 1674 1146 1676
rect 1266 1675 1267 1676
rect 1271 1675 1272 1679
rect 4714 1679 4715 1680
rect 4719 1679 4720 1683
rect 4852 1682 4854 1688
rect 4858 1687 4859 1691
rect 4863 1690 4864 1691
rect 5394 1691 5400 1692
rect 5394 1690 5395 1691
rect 4863 1688 4905 1690
rect 5317 1688 5395 1690
rect 4863 1687 4864 1688
rect 4858 1686 4864 1687
rect 5394 1687 5395 1688
rect 5399 1687 5400 1691
rect 5622 1691 5628 1692
rect 5622 1690 5623 1691
rect 5613 1688 5623 1690
rect 5394 1686 5400 1687
rect 5622 1687 5623 1688
rect 5627 1687 5628 1691
rect 5622 1686 5628 1687
rect 5022 1683 5028 1684
rect 5022 1682 5023 1683
rect 4852 1680 5023 1682
rect 4714 1678 4720 1679
rect 5022 1679 5023 1680
rect 5027 1679 5028 1683
rect 5022 1678 5028 1679
rect 1266 1674 1272 1675
rect 1290 1675 1296 1676
rect 1109 1672 1146 1674
rect 926 1670 932 1671
rect 1242 1671 1248 1672
rect 1242 1667 1243 1671
rect 1247 1667 1248 1671
rect 1290 1671 1291 1675
rect 1295 1671 1296 1675
rect 1290 1670 1296 1671
rect 1426 1671 1432 1672
rect 1242 1666 1248 1667
rect 1426 1667 1427 1671
rect 1431 1667 1432 1671
rect 1426 1666 1432 1667
rect 1562 1671 1568 1672
rect 1562 1667 1563 1671
rect 1567 1667 1568 1671
rect 1562 1666 1568 1667
rect 2754 1663 2760 1664
rect 2754 1662 2755 1663
rect 2725 1660 2755 1662
rect 2178 1659 2184 1660
rect 2178 1655 2179 1659
rect 2183 1655 2184 1659
rect 2178 1654 2184 1655
rect 2226 1659 2232 1660
rect 2226 1655 2227 1659
rect 2231 1655 2232 1659
rect 2226 1654 2232 1655
rect 2362 1659 2368 1660
rect 2362 1655 2363 1659
rect 2367 1655 2368 1659
rect 2362 1654 2368 1655
rect 2498 1659 2504 1660
rect 2498 1655 2499 1659
rect 2503 1655 2504 1659
rect 2754 1659 2755 1660
rect 2759 1659 2760 1663
rect 2754 1658 2760 1659
rect 2778 1659 2784 1660
rect 2498 1654 2504 1655
rect 2778 1655 2779 1659
rect 2783 1655 2784 1659
rect 2778 1654 2784 1655
rect 2922 1659 2928 1660
rect 2922 1655 2923 1659
rect 2927 1655 2928 1659
rect 4262 1659 4268 1660
rect 4262 1658 4263 1659
rect 2922 1654 2928 1655
rect 3996 1656 4263 1658
rect 3996 1654 3998 1656
rect 4262 1655 4263 1656
rect 4267 1655 4268 1659
rect 4262 1654 4268 1655
rect 4434 1655 4440 1656
rect 4434 1654 4435 1655
rect 3957 1652 3998 1654
rect 4421 1652 4435 1654
rect 4002 1651 4008 1652
rect 4002 1647 4003 1651
rect 4007 1647 4008 1651
rect 4002 1646 4008 1647
rect 4146 1651 4152 1652
rect 4146 1647 4147 1651
rect 4151 1647 4152 1651
rect 4434 1651 4435 1652
rect 4439 1651 4440 1655
rect 5402 1655 5408 1656
rect 5402 1654 5403 1655
rect 5373 1652 5403 1654
rect 4434 1650 4440 1651
rect 4538 1651 4544 1652
rect 4146 1646 4152 1647
rect 4538 1647 4539 1651
rect 4543 1647 4544 1651
rect 4538 1646 4544 1647
rect 4770 1651 4776 1652
rect 4770 1647 4771 1651
rect 4775 1647 4776 1651
rect 4770 1646 4776 1647
rect 5018 1651 5024 1652
rect 5018 1647 5019 1651
rect 5023 1647 5024 1651
rect 5402 1651 5403 1652
rect 5407 1651 5408 1655
rect 5634 1655 5640 1656
rect 5634 1654 5635 1655
rect 5613 1652 5635 1654
rect 5402 1650 5408 1651
rect 5634 1651 5635 1652
rect 5639 1651 5640 1655
rect 5634 1650 5640 1651
rect 5018 1646 5024 1647
rect 1242 1643 1248 1644
rect 1242 1639 1243 1643
rect 1247 1642 1248 1643
rect 1678 1643 1684 1644
rect 1678 1642 1679 1643
rect 1247 1640 1679 1642
rect 1247 1639 1248 1640
rect 1242 1638 1248 1639
rect 1678 1639 1679 1640
rect 1683 1639 1684 1643
rect 1678 1638 1684 1639
rect 110 1624 116 1625
rect 1934 1624 1940 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 110 1619 116 1620
rect 874 1623 880 1624
rect 874 1619 875 1623
rect 879 1619 880 1623
rect 874 1618 880 1619
rect 1010 1623 1016 1624
rect 1010 1619 1011 1623
rect 1015 1619 1016 1623
rect 1010 1618 1016 1619
rect 1146 1623 1152 1624
rect 1146 1619 1147 1623
rect 1151 1619 1152 1623
rect 1146 1618 1152 1619
rect 1282 1623 1288 1624
rect 1282 1619 1283 1623
rect 1287 1619 1288 1623
rect 1282 1618 1288 1619
rect 1418 1623 1424 1624
rect 1418 1619 1419 1623
rect 1423 1619 1424 1623
rect 1418 1618 1424 1619
rect 1554 1623 1560 1624
rect 1554 1619 1555 1623
rect 1559 1619 1560 1623
rect 1934 1620 1935 1624
rect 1939 1620 1940 1624
rect 1934 1619 1940 1620
rect 1554 1618 1560 1619
rect 1974 1612 1980 1613
rect 3798 1612 3804 1613
rect 902 1608 908 1609
rect 1038 1608 1044 1609
rect 1174 1608 1180 1609
rect 1310 1608 1316 1609
rect 1446 1608 1452 1609
rect 1582 1608 1588 1609
rect 1974 1608 1975 1612
rect 1979 1608 1980 1612
rect 110 1607 116 1608
rect 110 1603 111 1607
rect 115 1603 116 1607
rect 902 1604 903 1608
rect 907 1604 908 1608
rect 902 1603 908 1604
rect 998 1607 1005 1608
rect 998 1603 999 1607
rect 1004 1603 1005 1607
rect 1038 1604 1039 1608
rect 1043 1604 1044 1608
rect 1038 1603 1044 1604
rect 1134 1607 1141 1608
rect 1134 1603 1135 1607
rect 1140 1603 1141 1607
rect 1174 1604 1175 1608
rect 1179 1604 1180 1608
rect 1174 1603 1180 1604
rect 1266 1607 1277 1608
rect 1266 1603 1267 1607
rect 1271 1603 1272 1607
rect 1276 1603 1277 1607
rect 1310 1604 1311 1608
rect 1315 1604 1316 1608
rect 1310 1603 1316 1604
rect 1407 1607 1413 1608
rect 1407 1603 1408 1607
rect 1412 1606 1413 1607
rect 1426 1607 1432 1608
rect 1426 1606 1427 1607
rect 1412 1604 1427 1606
rect 1412 1603 1413 1604
rect 110 1602 116 1603
rect 998 1602 1005 1603
rect 1134 1602 1141 1603
rect 1266 1602 1277 1603
rect 1407 1602 1413 1603
rect 1426 1603 1427 1604
rect 1431 1603 1432 1607
rect 1446 1604 1447 1608
rect 1451 1604 1452 1608
rect 1446 1603 1452 1604
rect 1543 1607 1549 1608
rect 1543 1603 1544 1607
rect 1548 1606 1549 1607
rect 1562 1607 1568 1608
rect 1562 1606 1563 1607
rect 1548 1604 1563 1606
rect 1548 1603 1549 1604
rect 1426 1602 1432 1603
rect 1543 1602 1549 1603
rect 1562 1603 1563 1604
rect 1567 1603 1568 1607
rect 1582 1604 1583 1608
rect 1587 1604 1588 1608
rect 1582 1603 1588 1604
rect 1678 1607 1685 1608
rect 1678 1603 1679 1607
rect 1684 1603 1685 1607
rect 1562 1602 1568 1603
rect 1678 1602 1685 1603
rect 1934 1607 1940 1608
rect 1974 1607 1980 1608
rect 2082 1611 2088 1612
rect 2082 1607 2083 1611
rect 2087 1607 2088 1611
rect 1934 1603 1935 1607
rect 1939 1603 1940 1607
rect 2082 1606 2088 1607
rect 2218 1611 2224 1612
rect 2218 1607 2219 1611
rect 2223 1607 2224 1611
rect 2218 1606 2224 1607
rect 2354 1611 2360 1612
rect 2354 1607 2355 1611
rect 2359 1607 2360 1611
rect 2354 1606 2360 1607
rect 2490 1611 2496 1612
rect 2490 1607 2491 1611
rect 2495 1607 2496 1611
rect 2490 1606 2496 1607
rect 2626 1611 2632 1612
rect 2626 1607 2627 1611
rect 2631 1607 2632 1611
rect 2626 1606 2632 1607
rect 2770 1611 2776 1612
rect 2770 1607 2771 1611
rect 2775 1607 2776 1611
rect 2770 1606 2776 1607
rect 2914 1611 2920 1612
rect 2914 1607 2915 1611
rect 2919 1607 2920 1611
rect 3798 1608 3799 1612
rect 3803 1608 3804 1612
rect 3798 1607 3804 1608
rect 2914 1606 2920 1607
rect 1934 1602 1940 1603
rect 3838 1604 3844 1605
rect 5662 1604 5668 1605
rect 3838 1600 3839 1604
rect 3843 1600 3844 1604
rect 3838 1599 3844 1600
rect 3858 1603 3864 1604
rect 3858 1599 3859 1603
rect 3863 1599 3864 1603
rect 3858 1598 3864 1599
rect 3994 1603 4000 1604
rect 3994 1599 3995 1603
rect 3999 1599 4000 1603
rect 3994 1598 4000 1599
rect 4138 1603 4144 1604
rect 4138 1599 4139 1603
rect 4143 1599 4144 1603
rect 4138 1598 4144 1599
rect 4322 1603 4328 1604
rect 4322 1599 4323 1603
rect 4327 1599 4328 1603
rect 4322 1598 4328 1599
rect 4530 1603 4536 1604
rect 4530 1599 4531 1603
rect 4535 1599 4536 1603
rect 4530 1598 4536 1599
rect 4762 1603 4768 1604
rect 4762 1599 4763 1603
rect 4767 1599 4768 1603
rect 4762 1598 4768 1599
rect 5010 1603 5016 1604
rect 5010 1599 5011 1603
rect 5015 1599 5016 1603
rect 5010 1598 5016 1599
rect 5274 1603 5280 1604
rect 5274 1599 5275 1603
rect 5279 1599 5280 1603
rect 5274 1598 5280 1599
rect 5514 1603 5520 1604
rect 5514 1599 5515 1603
rect 5519 1599 5520 1603
rect 5662 1600 5663 1604
rect 5667 1600 5668 1604
rect 5662 1599 5668 1600
rect 5514 1598 5520 1599
rect 2110 1596 2116 1597
rect 2246 1596 2252 1597
rect 2382 1596 2388 1597
rect 2518 1596 2524 1597
rect 2654 1596 2660 1597
rect 2798 1596 2804 1597
rect 2942 1596 2948 1597
rect 1974 1595 1980 1596
rect 1974 1591 1975 1595
rect 1979 1591 1980 1595
rect 2110 1592 2111 1596
rect 2115 1592 2116 1596
rect 2110 1591 2116 1592
rect 2207 1595 2213 1596
rect 2207 1591 2208 1595
rect 2212 1594 2213 1595
rect 2226 1595 2232 1596
rect 2226 1594 2227 1595
rect 2212 1592 2227 1594
rect 2212 1591 2213 1592
rect 1974 1590 1980 1591
rect 2207 1590 2213 1591
rect 2226 1591 2227 1592
rect 2231 1591 2232 1595
rect 2246 1592 2247 1596
rect 2251 1592 2252 1596
rect 2246 1591 2252 1592
rect 2343 1595 2349 1596
rect 2343 1591 2344 1595
rect 2348 1594 2349 1595
rect 2362 1595 2368 1596
rect 2362 1594 2363 1595
rect 2348 1592 2363 1594
rect 2348 1591 2349 1592
rect 2226 1590 2232 1591
rect 2343 1590 2349 1591
rect 2362 1591 2363 1592
rect 2367 1591 2368 1595
rect 2382 1592 2383 1596
rect 2387 1592 2388 1596
rect 2382 1591 2388 1592
rect 2479 1595 2485 1596
rect 2479 1591 2480 1595
rect 2484 1594 2485 1595
rect 2498 1595 2504 1596
rect 2498 1594 2499 1595
rect 2484 1592 2499 1594
rect 2484 1591 2485 1592
rect 2362 1590 2368 1591
rect 2479 1590 2485 1591
rect 2498 1591 2499 1592
rect 2503 1591 2504 1595
rect 2518 1592 2519 1596
rect 2523 1592 2524 1596
rect 2518 1591 2524 1592
rect 2610 1595 2621 1596
rect 2610 1591 2611 1595
rect 2615 1591 2616 1595
rect 2620 1591 2621 1595
rect 2654 1592 2655 1596
rect 2659 1592 2660 1596
rect 2654 1591 2660 1592
rect 2751 1595 2757 1596
rect 2751 1591 2752 1595
rect 2756 1594 2757 1595
rect 2778 1595 2784 1596
rect 2778 1594 2779 1595
rect 2756 1592 2779 1594
rect 2756 1591 2757 1592
rect 2498 1590 2504 1591
rect 2610 1590 2621 1591
rect 2751 1590 2757 1591
rect 2778 1591 2779 1592
rect 2783 1591 2784 1595
rect 2798 1592 2799 1596
rect 2803 1592 2804 1596
rect 2798 1591 2804 1592
rect 2895 1595 2901 1596
rect 2895 1591 2896 1595
rect 2900 1594 2901 1595
rect 2922 1595 2928 1596
rect 2922 1594 2923 1595
rect 2900 1592 2923 1594
rect 2900 1591 2901 1592
rect 2778 1590 2784 1591
rect 2895 1590 2901 1591
rect 2922 1591 2923 1592
rect 2927 1591 2928 1595
rect 2942 1592 2943 1596
rect 2947 1592 2948 1596
rect 2942 1591 2948 1592
rect 3038 1595 3045 1596
rect 3038 1591 3039 1595
rect 3044 1591 3045 1595
rect 2922 1590 2928 1591
rect 3038 1590 3045 1591
rect 3798 1595 3804 1596
rect 3798 1591 3799 1595
rect 3803 1591 3804 1595
rect 3798 1590 3804 1591
rect 3886 1588 3892 1589
rect 4022 1588 4028 1589
rect 4166 1588 4172 1589
rect 4350 1588 4356 1589
rect 4558 1588 4564 1589
rect 4790 1588 4796 1589
rect 5038 1588 5044 1589
rect 5302 1588 5308 1589
rect 5542 1588 5548 1589
rect 3838 1587 3844 1588
rect 3838 1583 3839 1587
rect 3843 1583 3844 1587
rect 3886 1584 3887 1588
rect 3891 1584 3892 1588
rect 3886 1583 3892 1584
rect 3978 1587 3989 1588
rect 3978 1583 3979 1587
rect 3983 1583 3984 1587
rect 3988 1583 3989 1587
rect 4022 1584 4023 1588
rect 4027 1584 4028 1588
rect 4022 1583 4028 1584
rect 4119 1587 4125 1588
rect 4119 1583 4120 1587
rect 4124 1586 4125 1587
rect 4146 1587 4152 1588
rect 4146 1586 4147 1587
rect 4124 1584 4147 1586
rect 4124 1583 4125 1584
rect 3838 1582 3844 1583
rect 3978 1582 3989 1583
rect 4119 1582 4125 1583
rect 4146 1583 4147 1584
rect 4151 1583 4152 1587
rect 4166 1584 4167 1588
rect 4171 1584 4172 1588
rect 4166 1583 4172 1584
rect 4262 1587 4269 1588
rect 4262 1583 4263 1587
rect 4268 1583 4269 1587
rect 4350 1584 4351 1588
rect 4355 1584 4356 1588
rect 4350 1583 4356 1584
rect 4447 1587 4453 1588
rect 4447 1583 4448 1587
rect 4452 1586 4453 1587
rect 4538 1587 4544 1588
rect 4538 1586 4539 1587
rect 4452 1584 4539 1586
rect 4452 1583 4453 1584
rect 4146 1582 4152 1583
rect 4262 1582 4269 1583
rect 4447 1582 4453 1583
rect 4538 1583 4539 1584
rect 4543 1583 4544 1587
rect 4558 1584 4559 1588
rect 4563 1584 4564 1588
rect 4558 1583 4564 1584
rect 4655 1587 4661 1588
rect 4655 1583 4656 1587
rect 4660 1586 4661 1587
rect 4770 1587 4776 1588
rect 4770 1586 4771 1587
rect 4660 1584 4771 1586
rect 4660 1583 4661 1584
rect 4538 1582 4544 1583
rect 4655 1582 4661 1583
rect 4770 1583 4771 1584
rect 4775 1583 4776 1587
rect 4790 1584 4791 1588
rect 4795 1584 4796 1588
rect 4790 1583 4796 1584
rect 4887 1587 4893 1588
rect 4887 1583 4888 1587
rect 4892 1586 4893 1587
rect 5018 1587 5024 1588
rect 5018 1586 5019 1587
rect 4892 1584 5019 1586
rect 4892 1583 4893 1584
rect 4770 1582 4776 1583
rect 4887 1582 4893 1583
rect 5018 1583 5019 1584
rect 5023 1583 5024 1587
rect 5038 1584 5039 1588
rect 5043 1584 5044 1588
rect 5038 1583 5044 1584
rect 5130 1587 5141 1588
rect 5130 1583 5131 1587
rect 5135 1583 5136 1587
rect 5140 1583 5141 1587
rect 5302 1584 5303 1588
rect 5307 1584 5308 1588
rect 5302 1583 5308 1584
rect 5394 1587 5405 1588
rect 5394 1583 5395 1587
rect 5399 1583 5400 1587
rect 5404 1583 5405 1587
rect 5542 1584 5543 1588
rect 5547 1584 5548 1588
rect 5542 1583 5548 1584
rect 5638 1587 5645 1588
rect 5638 1583 5639 1587
rect 5644 1583 5645 1587
rect 5018 1582 5024 1583
rect 5130 1582 5141 1583
rect 5394 1582 5405 1583
rect 5638 1582 5645 1583
rect 5662 1587 5668 1588
rect 5662 1583 5663 1587
rect 5667 1583 5668 1587
rect 5662 1582 5668 1583
rect 2178 1547 2184 1548
rect 2178 1543 2179 1547
rect 2183 1546 2184 1547
rect 2183 1544 2242 1546
rect 2183 1543 2184 1544
rect 2178 1542 2184 1543
rect 1974 1533 1980 1534
rect 110 1529 116 1530
rect 1934 1529 1940 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 158 1528 164 1529
rect 390 1528 396 1529
rect 630 1528 636 1529
rect 870 1528 876 1529
rect 1110 1528 1116 1529
rect 1350 1528 1356 1529
rect 158 1524 159 1528
rect 163 1524 164 1528
rect 158 1523 164 1524
rect 250 1527 261 1528
rect 250 1523 251 1527
rect 255 1523 256 1527
rect 260 1523 261 1527
rect 390 1524 391 1528
rect 395 1524 396 1528
rect 390 1523 396 1524
rect 487 1527 493 1528
rect 487 1523 488 1527
rect 492 1526 493 1527
rect 518 1527 524 1528
rect 518 1526 519 1527
rect 492 1524 519 1526
rect 492 1523 493 1524
rect 250 1522 261 1523
rect 487 1522 493 1523
rect 518 1523 519 1524
rect 523 1523 524 1527
rect 630 1524 631 1528
rect 635 1524 636 1528
rect 630 1523 636 1524
rect 727 1527 736 1528
rect 727 1523 728 1527
rect 735 1523 736 1527
rect 870 1524 871 1528
rect 875 1524 876 1528
rect 870 1523 876 1524
rect 967 1527 973 1528
rect 967 1523 968 1527
rect 972 1526 973 1527
rect 990 1527 996 1528
rect 990 1526 991 1527
rect 972 1524 991 1526
rect 972 1523 973 1524
rect 518 1522 524 1523
rect 727 1522 736 1523
rect 967 1522 973 1523
rect 990 1523 991 1524
rect 995 1523 996 1527
rect 1110 1524 1111 1528
rect 1115 1524 1116 1528
rect 1110 1523 1116 1524
rect 1207 1527 1213 1528
rect 1207 1523 1208 1527
rect 1212 1526 1213 1527
rect 1231 1527 1237 1528
rect 1231 1526 1232 1527
rect 1212 1524 1232 1526
rect 1212 1523 1213 1524
rect 990 1522 996 1523
rect 1207 1522 1213 1523
rect 1231 1523 1232 1524
rect 1236 1523 1237 1527
rect 1350 1524 1351 1528
rect 1355 1524 1356 1528
rect 1350 1523 1356 1524
rect 1442 1527 1453 1528
rect 1442 1523 1443 1527
rect 1447 1523 1448 1527
rect 1452 1523 1453 1527
rect 1934 1525 1935 1529
rect 1939 1525 1940 1529
rect 1974 1529 1975 1533
rect 1979 1529 1980 1533
rect 1974 1528 1980 1529
rect 2142 1532 2148 1533
rect 2240 1532 2242 1544
rect 3798 1533 3804 1534
rect 2278 1532 2284 1533
rect 2414 1532 2420 1533
rect 2550 1532 2556 1533
rect 2686 1532 2692 1533
rect 2822 1532 2828 1533
rect 2958 1532 2964 1533
rect 3094 1532 3100 1533
rect 3230 1532 3236 1533
rect 2142 1528 2143 1532
rect 2147 1528 2148 1532
rect 2142 1527 2148 1528
rect 2239 1531 2245 1532
rect 2239 1527 2240 1531
rect 2244 1527 2245 1531
rect 2278 1528 2279 1532
rect 2283 1528 2284 1532
rect 2278 1527 2284 1528
rect 2374 1531 2381 1532
rect 2374 1527 2375 1531
rect 2380 1527 2381 1531
rect 2414 1528 2415 1532
rect 2419 1528 2420 1532
rect 2414 1527 2420 1528
rect 2511 1531 2520 1532
rect 2511 1527 2512 1531
rect 2519 1527 2520 1531
rect 2550 1528 2551 1532
rect 2555 1528 2556 1532
rect 2550 1527 2556 1528
rect 2647 1531 2656 1532
rect 2647 1527 2648 1531
rect 2655 1527 2656 1531
rect 2686 1528 2687 1532
rect 2691 1528 2692 1532
rect 2686 1527 2692 1528
rect 2783 1531 2792 1532
rect 2783 1527 2784 1531
rect 2791 1527 2792 1531
rect 2822 1528 2823 1532
rect 2827 1528 2828 1532
rect 2822 1527 2828 1528
rect 2914 1531 2925 1532
rect 2914 1527 2915 1531
rect 2919 1527 2920 1531
rect 2924 1527 2925 1531
rect 2958 1528 2959 1532
rect 2963 1528 2964 1532
rect 2958 1527 2964 1528
rect 3055 1531 3064 1532
rect 3055 1527 3056 1531
rect 3063 1527 3064 1531
rect 3094 1528 3095 1532
rect 3099 1528 3100 1532
rect 3094 1527 3100 1528
rect 3191 1531 3200 1532
rect 3191 1527 3192 1531
rect 3199 1527 3200 1531
rect 3230 1528 3231 1532
rect 3235 1528 3236 1532
rect 3230 1527 3236 1528
rect 3322 1531 3333 1532
rect 3322 1527 3323 1531
rect 3327 1527 3328 1531
rect 3332 1527 3333 1531
rect 3798 1529 3799 1533
rect 3803 1529 3804 1533
rect 3798 1528 3804 1529
rect 2239 1526 2245 1527
rect 2374 1526 2381 1527
rect 2511 1526 2520 1527
rect 2647 1526 2656 1527
rect 2783 1526 2792 1527
rect 2914 1526 2925 1527
rect 3055 1526 3064 1527
rect 3191 1526 3200 1527
rect 3322 1526 3333 1527
rect 1934 1524 1940 1525
rect 3838 1525 3844 1526
rect 5662 1525 5668 1526
rect 1231 1522 1237 1523
rect 1442 1522 1453 1523
rect 3838 1521 3839 1525
rect 3843 1521 3844 1525
rect 3838 1520 3844 1521
rect 3886 1524 3892 1525
rect 4110 1524 4116 1525
rect 4342 1524 4348 1525
rect 4574 1524 4580 1525
rect 4814 1524 4820 1525
rect 5062 1524 5068 1525
rect 5310 1524 5316 1525
rect 5542 1524 5548 1525
rect 3886 1520 3887 1524
rect 3891 1520 3892 1524
rect 3886 1519 3892 1520
rect 3983 1523 3989 1524
rect 3983 1519 3984 1523
rect 3988 1522 3989 1523
rect 4002 1523 4008 1524
rect 4002 1522 4003 1523
rect 3988 1520 4003 1522
rect 3988 1519 3989 1520
rect 3983 1518 3989 1519
rect 4002 1519 4003 1520
rect 4007 1519 4008 1523
rect 4110 1520 4111 1524
rect 4115 1520 4116 1524
rect 4110 1519 4116 1520
rect 4206 1523 4213 1524
rect 4206 1519 4207 1523
rect 4212 1519 4213 1523
rect 4342 1520 4343 1524
rect 4347 1520 4348 1524
rect 4342 1519 4348 1520
rect 4439 1523 4445 1524
rect 4439 1519 4440 1523
rect 4444 1522 4445 1523
rect 4447 1523 4453 1524
rect 4447 1522 4448 1523
rect 4444 1520 4448 1522
rect 4444 1519 4445 1520
rect 4002 1518 4008 1519
rect 4206 1518 4213 1519
rect 4439 1518 4445 1519
rect 4447 1519 4448 1520
rect 4452 1519 4453 1523
rect 4574 1520 4575 1524
rect 4579 1520 4580 1524
rect 4574 1519 4580 1520
rect 4671 1523 4677 1524
rect 4671 1519 4672 1523
rect 4676 1522 4677 1523
rect 4702 1523 4708 1524
rect 4702 1522 4703 1523
rect 4676 1520 4703 1522
rect 4676 1519 4677 1520
rect 4447 1518 4453 1519
rect 4671 1518 4677 1519
rect 4702 1519 4703 1520
rect 4707 1519 4708 1523
rect 4814 1520 4815 1524
rect 4819 1520 4820 1524
rect 4814 1519 4820 1520
rect 4911 1523 4917 1524
rect 4911 1519 4912 1523
rect 4916 1522 4917 1523
rect 4950 1523 4956 1524
rect 4950 1522 4951 1523
rect 4916 1520 4951 1522
rect 4916 1519 4917 1520
rect 4702 1518 4708 1519
rect 4911 1518 4917 1519
rect 4950 1519 4951 1520
rect 4955 1519 4956 1523
rect 5062 1520 5063 1524
rect 5067 1520 5068 1524
rect 5062 1519 5068 1520
rect 5154 1523 5165 1524
rect 5154 1519 5155 1523
rect 5159 1519 5160 1523
rect 5164 1519 5165 1523
rect 5310 1520 5311 1524
rect 5315 1520 5316 1524
rect 5310 1519 5316 1520
rect 5402 1523 5413 1524
rect 5402 1519 5403 1523
rect 5407 1519 5408 1523
rect 5412 1519 5413 1523
rect 5542 1520 5543 1524
rect 5547 1520 5548 1524
rect 5542 1519 5548 1520
rect 5639 1524 5645 1525
rect 5639 1520 5640 1524
rect 5644 1523 5645 1524
rect 5647 1523 5653 1524
rect 5644 1521 5648 1523
rect 5644 1520 5645 1521
rect 5639 1519 5645 1520
rect 5647 1519 5648 1521
rect 5652 1519 5653 1523
rect 5662 1521 5663 1525
rect 5667 1521 5668 1525
rect 5662 1520 5668 1521
rect 4950 1518 4956 1519
rect 5154 1518 5165 1519
rect 5402 1518 5413 1519
rect 5647 1518 5653 1519
rect 2114 1517 2120 1518
rect 1974 1516 1980 1517
rect 130 1513 136 1514
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 130 1509 131 1513
rect 135 1509 136 1513
rect 130 1508 136 1509
rect 362 1513 368 1514
rect 362 1509 363 1513
rect 367 1509 368 1513
rect 362 1508 368 1509
rect 602 1513 608 1514
rect 602 1509 603 1513
rect 607 1509 608 1513
rect 602 1508 608 1509
rect 842 1513 848 1514
rect 842 1509 843 1513
rect 847 1509 848 1513
rect 842 1508 848 1509
rect 1082 1513 1088 1514
rect 1082 1509 1083 1513
rect 1087 1509 1088 1513
rect 1082 1508 1088 1509
rect 1322 1513 1328 1514
rect 1322 1509 1323 1513
rect 1327 1509 1328 1513
rect 1322 1508 1328 1509
rect 1934 1512 1940 1513
rect 1934 1508 1935 1512
rect 1939 1508 1940 1512
rect 1974 1512 1975 1516
rect 1979 1512 1980 1516
rect 2114 1513 2115 1517
rect 2119 1513 2120 1517
rect 2114 1512 2120 1513
rect 2250 1517 2256 1518
rect 2250 1513 2251 1517
rect 2255 1513 2256 1517
rect 2250 1512 2256 1513
rect 2386 1517 2392 1518
rect 2386 1513 2387 1517
rect 2391 1513 2392 1517
rect 2386 1512 2392 1513
rect 2522 1517 2528 1518
rect 2522 1513 2523 1517
rect 2527 1513 2528 1517
rect 2522 1512 2528 1513
rect 2658 1517 2664 1518
rect 2658 1513 2659 1517
rect 2663 1513 2664 1517
rect 2658 1512 2664 1513
rect 2794 1517 2800 1518
rect 2794 1513 2795 1517
rect 2799 1513 2800 1517
rect 2794 1512 2800 1513
rect 2930 1517 2936 1518
rect 2930 1513 2931 1517
rect 2935 1513 2936 1517
rect 2930 1512 2936 1513
rect 3066 1517 3072 1518
rect 3066 1513 3067 1517
rect 3071 1513 3072 1517
rect 3066 1512 3072 1513
rect 3202 1517 3208 1518
rect 3202 1513 3203 1517
rect 3207 1513 3208 1517
rect 3202 1512 3208 1513
rect 3798 1516 3804 1517
rect 3798 1512 3799 1516
rect 3803 1512 3804 1516
rect 1974 1511 1980 1512
rect 3798 1511 3804 1512
rect 3858 1509 3864 1510
rect 110 1507 116 1508
rect 458 1507 464 1508
rect 458 1503 459 1507
rect 463 1506 464 1507
rect 998 1507 1004 1508
rect 1934 1507 1940 1508
rect 3838 1508 3844 1509
rect 998 1506 999 1507
rect 463 1504 999 1506
rect 463 1503 464 1504
rect 458 1502 464 1503
rect 998 1503 999 1504
rect 1003 1503 1004 1507
rect 3838 1504 3839 1508
rect 3843 1504 3844 1508
rect 3858 1505 3859 1509
rect 3863 1505 3864 1509
rect 3858 1504 3864 1505
rect 4082 1509 4088 1510
rect 4082 1505 4083 1509
rect 4087 1505 4088 1509
rect 4082 1504 4088 1505
rect 4314 1509 4320 1510
rect 4314 1505 4315 1509
rect 4319 1505 4320 1509
rect 4314 1504 4320 1505
rect 4546 1509 4552 1510
rect 4546 1505 4547 1509
rect 4551 1505 4552 1509
rect 4546 1504 4552 1505
rect 4786 1509 4792 1510
rect 4786 1505 4787 1509
rect 4791 1505 4792 1509
rect 4786 1504 4792 1505
rect 5034 1509 5040 1510
rect 5034 1505 5035 1509
rect 5039 1505 5040 1509
rect 5034 1504 5040 1505
rect 5282 1509 5288 1510
rect 5282 1505 5283 1509
rect 5287 1505 5288 1509
rect 5282 1504 5288 1505
rect 5514 1509 5520 1510
rect 5514 1505 5515 1509
rect 5519 1505 5520 1509
rect 5514 1504 5520 1505
rect 5662 1508 5668 1509
rect 5662 1504 5663 1508
rect 5667 1504 5668 1508
rect 3838 1503 3844 1504
rect 3954 1503 3960 1504
rect 998 1502 1004 1503
rect 3954 1499 3955 1503
rect 3959 1502 3960 1503
rect 4206 1503 4212 1504
rect 4206 1502 4207 1503
rect 3959 1500 4207 1502
rect 3959 1499 3960 1500
rect 3954 1498 3960 1499
rect 4206 1499 4207 1500
rect 4211 1499 4212 1503
rect 4206 1498 4212 1499
rect 4418 1503 4424 1504
rect 4418 1499 4419 1503
rect 4423 1502 4424 1503
rect 5154 1503 5160 1504
rect 5662 1503 5668 1504
rect 5154 1502 5155 1503
rect 4423 1500 5155 1502
rect 4423 1499 4424 1500
rect 4418 1498 4424 1499
rect 5154 1499 5155 1500
rect 5159 1499 5160 1503
rect 5154 1498 5160 1499
rect 4410 1495 4416 1496
rect 2346 1491 2352 1492
rect 2346 1487 2347 1491
rect 2351 1490 2352 1491
rect 2914 1491 2920 1492
rect 2914 1490 2915 1491
rect 2351 1488 2915 1490
rect 2351 1487 2352 1488
rect 2346 1486 2352 1487
rect 2914 1487 2915 1488
rect 2919 1487 2920 1491
rect 4410 1491 4411 1495
rect 4415 1494 4416 1495
rect 5130 1495 5136 1496
rect 5130 1494 5131 1495
rect 4415 1492 5131 1494
rect 4415 1491 4416 1492
rect 4410 1490 4416 1491
rect 5130 1491 5131 1492
rect 5135 1491 5136 1495
rect 5130 1490 5136 1491
rect 2914 1486 2920 1487
rect 2346 1467 2352 1468
rect 458 1463 464 1464
rect 229 1460 261 1462
rect 259 1454 261 1460
rect 458 1459 459 1463
rect 463 1459 464 1463
rect 458 1458 464 1459
rect 518 1463 524 1464
rect 518 1459 519 1463
rect 523 1462 524 1463
rect 1134 1463 1140 1464
rect 523 1460 609 1462
rect 523 1459 524 1460
rect 518 1458 524 1459
rect 454 1455 460 1456
rect 454 1454 455 1455
rect 259 1452 455 1454
rect 454 1451 455 1452
rect 459 1451 460 1455
rect 940 1454 942 1461
rect 1134 1459 1135 1463
rect 1139 1459 1140 1463
rect 1134 1458 1140 1459
rect 1231 1463 1237 1464
rect 1231 1459 1232 1463
rect 1236 1462 1237 1463
rect 1236 1460 1329 1462
rect 1236 1459 1237 1460
rect 1231 1458 1237 1459
rect 2212 1458 2214 1465
rect 2346 1463 2347 1467
rect 2351 1463 2352 1467
rect 2514 1467 2520 1468
rect 2346 1462 2352 1463
rect 2374 1459 2380 1460
rect 2374 1458 2375 1459
rect 2212 1456 2375 1458
rect 1442 1455 1448 1456
rect 1442 1454 1443 1455
rect 940 1452 1443 1454
rect 454 1450 460 1451
rect 1442 1451 1443 1452
rect 1447 1451 1448 1455
rect 2374 1455 2375 1456
rect 2379 1455 2380 1459
rect 2484 1458 2486 1465
rect 2514 1463 2515 1467
rect 2519 1466 2520 1467
rect 2650 1467 2656 1468
rect 2519 1464 2529 1466
rect 2519 1463 2520 1464
rect 2514 1462 2520 1463
rect 2650 1463 2651 1467
rect 2655 1466 2656 1467
rect 2786 1467 2792 1468
rect 2655 1464 2665 1466
rect 2655 1463 2656 1464
rect 2650 1462 2656 1463
rect 2786 1463 2787 1467
rect 2791 1466 2792 1467
rect 3038 1467 3044 1468
rect 3038 1466 3039 1467
rect 2791 1464 2801 1466
rect 3029 1464 3039 1466
rect 2791 1463 2792 1464
rect 2786 1462 2792 1463
rect 3038 1463 3039 1464
rect 3043 1463 3044 1467
rect 3038 1462 3044 1463
rect 3058 1467 3064 1468
rect 3058 1463 3059 1467
rect 3063 1466 3064 1467
rect 3194 1467 3200 1468
rect 3063 1464 3073 1466
rect 3063 1463 3064 1464
rect 3058 1462 3064 1463
rect 3194 1463 3195 1467
rect 3199 1466 3200 1467
rect 3199 1464 3209 1466
rect 3199 1463 3200 1464
rect 3194 1462 3200 1463
rect 2814 1459 2820 1460
rect 2814 1458 2815 1459
rect 2484 1456 2815 1458
rect 2374 1454 2380 1455
rect 2814 1455 2815 1456
rect 2819 1455 2820 1459
rect 2814 1454 2820 1455
rect 3954 1459 3960 1460
rect 3954 1455 3955 1459
rect 3959 1455 3960 1459
rect 4202 1459 4208 1460
rect 4202 1458 4203 1459
rect 4181 1456 4203 1458
rect 3954 1454 3960 1455
rect 4202 1455 4203 1456
rect 4207 1455 4208 1459
rect 4202 1454 4208 1455
rect 4410 1459 4416 1460
rect 4410 1455 4411 1459
rect 4415 1455 4416 1459
rect 4410 1454 4416 1455
rect 4447 1459 4453 1460
rect 4447 1455 4448 1459
rect 4452 1458 4453 1459
rect 4702 1459 4708 1460
rect 4452 1456 4553 1458
rect 4452 1455 4453 1456
rect 4447 1454 4453 1455
rect 4702 1455 4703 1459
rect 4707 1458 4708 1459
rect 4950 1459 4956 1460
rect 4707 1456 4793 1458
rect 4707 1455 4708 1456
rect 4702 1454 4708 1455
rect 4950 1455 4951 1459
rect 4955 1458 4956 1459
rect 5638 1459 5644 1460
rect 5638 1458 5639 1459
rect 4955 1456 5041 1458
rect 4955 1455 4956 1456
rect 4950 1454 4956 1455
rect 1442 1450 1448 1451
rect 5380 1450 5382 1457
rect 5613 1456 5639 1458
rect 5638 1455 5639 1456
rect 5643 1455 5644 1459
rect 5638 1454 5644 1455
rect 5542 1451 5548 1452
rect 5542 1450 5543 1451
rect 5380 1448 5543 1450
rect 5542 1447 5543 1448
rect 5547 1447 5548 1451
rect 5542 1446 5548 1447
rect 3982 1427 3988 1428
rect 3982 1426 3983 1427
rect 3957 1424 3983 1426
rect 3982 1423 3983 1424
rect 3987 1423 3988 1427
rect 4418 1427 4424 1428
rect 3982 1422 3988 1423
rect 4090 1423 4096 1424
rect 254 1419 260 1420
rect 254 1418 255 1419
rect 229 1416 255 1418
rect 254 1415 255 1416
rect 259 1415 260 1419
rect 730 1419 736 1420
rect 254 1414 260 1415
rect 338 1415 344 1416
rect 338 1411 339 1415
rect 343 1411 344 1415
rect 338 1410 344 1411
rect 650 1415 656 1416
rect 650 1411 651 1415
rect 655 1411 656 1415
rect 730 1415 731 1419
rect 735 1418 736 1419
rect 990 1419 996 1420
rect 735 1416 785 1418
rect 735 1415 736 1416
rect 730 1414 736 1415
rect 990 1415 991 1419
rect 995 1418 996 1419
rect 2991 1419 2997 1420
rect 2991 1418 2992 1419
rect 995 1416 1009 1418
rect 2949 1416 2992 1418
rect 995 1415 996 1416
rect 990 1414 996 1415
rect 2194 1415 2200 1416
rect 650 1410 656 1411
rect 2194 1411 2195 1415
rect 2199 1411 2200 1415
rect 2194 1410 2200 1411
rect 2250 1415 2256 1416
rect 2250 1411 2251 1415
rect 2255 1411 2256 1415
rect 2250 1410 2256 1411
rect 2394 1415 2400 1416
rect 2394 1411 2395 1415
rect 2399 1411 2400 1415
rect 2394 1410 2400 1411
rect 2546 1415 2552 1416
rect 2546 1411 2547 1415
rect 2551 1411 2552 1415
rect 2546 1410 2552 1411
rect 2698 1415 2704 1416
rect 2698 1411 2699 1415
rect 2703 1411 2704 1415
rect 2991 1415 2992 1416
rect 2996 1415 2997 1419
rect 3151 1419 3157 1420
rect 3151 1418 3152 1419
rect 3109 1416 3152 1418
rect 2991 1414 2997 1415
rect 3151 1415 3152 1416
rect 3156 1415 3157 1419
rect 3322 1419 3328 1420
rect 3322 1418 3323 1419
rect 3269 1416 3323 1418
rect 3151 1414 3157 1415
rect 3322 1415 3323 1416
rect 3327 1415 3328 1419
rect 4090 1419 4091 1423
rect 4095 1419 4096 1423
rect 4418 1423 4419 1427
rect 4423 1423 4424 1427
rect 5534 1427 5540 1428
rect 5534 1426 5535 1427
rect 5517 1424 5535 1426
rect 4418 1422 4424 1423
rect 4554 1423 4560 1424
rect 4090 1418 4096 1419
rect 4554 1419 4555 1423
rect 4559 1419 4560 1423
rect 4554 1418 4560 1419
rect 4778 1423 4784 1424
rect 4778 1419 4779 1423
rect 4783 1419 4784 1423
rect 4778 1418 4784 1419
rect 4994 1423 5000 1424
rect 4994 1419 4995 1423
rect 4999 1419 5000 1423
rect 4994 1418 5000 1419
rect 5210 1423 5216 1424
rect 5210 1419 5211 1423
rect 5215 1419 5216 1423
rect 5534 1423 5535 1424
rect 5539 1423 5540 1427
rect 5534 1422 5540 1423
rect 5210 1418 5216 1419
rect 3322 1414 3328 1415
rect 2698 1410 2704 1411
rect 650 1395 656 1396
rect 650 1391 651 1395
rect 655 1394 656 1395
rect 1126 1395 1132 1396
rect 1126 1394 1127 1395
rect 655 1392 1127 1394
rect 655 1391 656 1392
rect 650 1390 656 1391
rect 1126 1391 1127 1392
rect 1131 1391 1132 1395
rect 1126 1390 1132 1391
rect 3838 1376 3844 1377
rect 5662 1376 5668 1377
rect 3838 1372 3839 1376
rect 3843 1372 3844 1376
rect 3838 1371 3844 1372
rect 3858 1375 3864 1376
rect 3858 1371 3859 1375
rect 3863 1371 3864 1375
rect 3858 1370 3864 1371
rect 4082 1375 4088 1376
rect 4082 1371 4083 1375
rect 4087 1371 4088 1375
rect 4082 1370 4088 1371
rect 4322 1375 4328 1376
rect 4322 1371 4323 1375
rect 4327 1371 4328 1375
rect 4322 1370 4328 1371
rect 4546 1375 4552 1376
rect 4546 1371 4547 1375
rect 4551 1371 4552 1375
rect 4546 1370 4552 1371
rect 4770 1375 4776 1376
rect 4770 1371 4771 1375
rect 4775 1371 4776 1375
rect 4770 1370 4776 1371
rect 4986 1375 4992 1376
rect 4986 1371 4987 1375
rect 4991 1371 4992 1375
rect 4986 1370 4992 1371
rect 5202 1375 5208 1376
rect 5202 1371 5203 1375
rect 5207 1371 5208 1375
rect 5202 1370 5208 1371
rect 5418 1375 5424 1376
rect 5418 1371 5419 1375
rect 5423 1371 5424 1375
rect 5662 1372 5663 1376
rect 5667 1372 5668 1376
rect 5662 1371 5668 1372
rect 5418 1370 5424 1371
rect 110 1368 116 1369
rect 1934 1368 1940 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 130 1367 136 1368
rect 130 1363 131 1367
rect 135 1363 136 1367
rect 130 1362 136 1363
rect 330 1367 336 1368
rect 330 1363 331 1367
rect 335 1363 336 1367
rect 330 1362 336 1363
rect 554 1367 560 1368
rect 554 1363 555 1367
rect 559 1363 560 1367
rect 554 1362 560 1363
rect 778 1367 784 1368
rect 778 1363 779 1367
rect 783 1363 784 1367
rect 778 1362 784 1363
rect 1002 1367 1008 1368
rect 1002 1363 1003 1367
rect 1007 1363 1008 1367
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 1934 1363 1940 1364
rect 1974 1368 1980 1369
rect 3798 1368 3804 1369
rect 1974 1364 1975 1368
rect 1979 1364 1980 1368
rect 1974 1363 1980 1364
rect 2098 1367 2104 1368
rect 2098 1363 2099 1367
rect 2103 1363 2104 1367
rect 1002 1362 1008 1363
rect 2098 1362 2104 1363
rect 2242 1367 2248 1368
rect 2242 1363 2243 1367
rect 2247 1363 2248 1367
rect 2242 1362 2248 1363
rect 2386 1367 2392 1368
rect 2386 1363 2387 1367
rect 2391 1363 2392 1367
rect 2386 1362 2392 1363
rect 2538 1367 2544 1368
rect 2538 1363 2539 1367
rect 2543 1363 2544 1367
rect 2538 1362 2544 1363
rect 2690 1367 2696 1368
rect 2690 1363 2691 1367
rect 2695 1363 2696 1367
rect 2690 1362 2696 1363
rect 2850 1367 2856 1368
rect 2850 1363 2851 1367
rect 2855 1363 2856 1367
rect 2850 1362 2856 1363
rect 3010 1367 3016 1368
rect 3010 1363 3011 1367
rect 3015 1363 3016 1367
rect 3010 1362 3016 1363
rect 3170 1367 3176 1368
rect 3170 1363 3171 1367
rect 3175 1363 3176 1367
rect 3798 1364 3799 1368
rect 3803 1364 3804 1368
rect 3798 1363 3804 1364
rect 3170 1362 3176 1363
rect 3886 1360 3892 1361
rect 4110 1360 4116 1361
rect 4350 1360 4356 1361
rect 4574 1360 4580 1361
rect 4798 1360 4804 1361
rect 5014 1360 5020 1361
rect 5230 1360 5236 1361
rect 5446 1360 5452 1361
rect 2991 1359 2997 1360
rect 2991 1355 2992 1359
rect 2996 1358 2997 1359
rect 3151 1359 3157 1360
rect 2996 1356 3138 1358
rect 2996 1355 2997 1356
rect 2991 1354 2997 1355
rect 158 1352 164 1353
rect 358 1352 364 1353
rect 582 1352 588 1353
rect 806 1352 812 1353
rect 1030 1352 1036 1353
rect 2126 1352 2132 1353
rect 2270 1352 2276 1353
rect 2414 1352 2420 1353
rect 2566 1352 2572 1353
rect 2718 1352 2724 1353
rect 2878 1352 2884 1353
rect 3038 1352 3044 1353
rect 3136 1352 3138 1356
rect 3151 1355 3152 1359
rect 3156 1358 3157 1359
rect 3838 1359 3844 1360
rect 3156 1356 3298 1358
rect 3156 1355 3157 1356
rect 3151 1354 3157 1355
rect 3198 1352 3204 1353
rect 3296 1352 3298 1356
rect 3838 1355 3839 1359
rect 3843 1355 3844 1359
rect 3886 1356 3887 1360
rect 3891 1356 3892 1360
rect 3886 1355 3892 1356
rect 3983 1359 3989 1360
rect 3983 1355 3984 1359
rect 3988 1358 3989 1359
rect 4090 1359 4096 1360
rect 4090 1358 4091 1359
rect 3988 1356 4091 1358
rect 3988 1355 3989 1356
rect 3838 1354 3844 1355
rect 3983 1354 3989 1355
rect 4090 1355 4091 1356
rect 4095 1355 4096 1359
rect 4110 1356 4111 1360
rect 4115 1356 4116 1360
rect 4110 1355 4116 1356
rect 4202 1359 4213 1360
rect 4202 1355 4203 1359
rect 4207 1355 4208 1359
rect 4212 1355 4213 1359
rect 4350 1356 4351 1360
rect 4355 1356 4356 1360
rect 4350 1355 4356 1356
rect 4447 1359 4453 1360
rect 4447 1355 4448 1359
rect 4452 1358 4453 1359
rect 4554 1359 4560 1360
rect 4554 1358 4555 1359
rect 4452 1356 4555 1358
rect 4452 1355 4453 1356
rect 4090 1354 4096 1355
rect 4202 1354 4213 1355
rect 4447 1354 4453 1355
rect 4554 1355 4555 1356
rect 4559 1355 4560 1359
rect 4574 1356 4575 1360
rect 4579 1356 4580 1360
rect 4574 1355 4580 1356
rect 4671 1359 4677 1360
rect 4671 1355 4672 1359
rect 4676 1358 4677 1359
rect 4778 1359 4784 1360
rect 4778 1358 4779 1359
rect 4676 1356 4779 1358
rect 4676 1355 4677 1356
rect 4554 1354 4560 1355
rect 4671 1354 4677 1355
rect 4778 1355 4779 1356
rect 4783 1355 4784 1359
rect 4798 1356 4799 1360
rect 4803 1356 4804 1360
rect 4798 1355 4804 1356
rect 4895 1359 4901 1360
rect 4895 1355 4896 1359
rect 4900 1358 4901 1359
rect 4994 1359 5000 1360
rect 4994 1358 4995 1359
rect 4900 1356 4995 1358
rect 4900 1355 4901 1356
rect 4778 1354 4784 1355
rect 4895 1354 4901 1355
rect 4994 1355 4995 1356
rect 4999 1355 5000 1359
rect 5014 1356 5015 1360
rect 5019 1356 5020 1360
rect 5014 1355 5020 1356
rect 5111 1359 5117 1360
rect 5111 1355 5112 1359
rect 5116 1358 5117 1359
rect 5210 1359 5216 1360
rect 5210 1358 5211 1359
rect 5116 1356 5211 1358
rect 5116 1355 5117 1356
rect 4994 1354 5000 1355
rect 5111 1354 5117 1355
rect 5210 1355 5211 1356
rect 5215 1355 5216 1359
rect 5230 1356 5231 1360
rect 5235 1356 5236 1360
rect 5230 1355 5236 1356
rect 5322 1359 5333 1360
rect 5322 1355 5323 1359
rect 5327 1355 5328 1359
rect 5332 1355 5333 1359
rect 5446 1356 5447 1360
rect 5451 1356 5452 1360
rect 5446 1355 5452 1356
rect 5542 1359 5549 1360
rect 5542 1355 5543 1359
rect 5548 1355 5549 1359
rect 5210 1354 5216 1355
rect 5322 1354 5333 1355
rect 5542 1354 5549 1355
rect 5662 1359 5668 1360
rect 5662 1355 5663 1359
rect 5667 1355 5668 1359
rect 5662 1354 5668 1355
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 158 1348 159 1352
rect 163 1348 164 1352
rect 158 1347 164 1348
rect 255 1351 261 1352
rect 255 1347 256 1351
rect 260 1350 261 1351
rect 338 1351 344 1352
rect 338 1350 339 1351
rect 260 1348 339 1350
rect 260 1347 261 1348
rect 110 1346 116 1347
rect 255 1346 261 1347
rect 338 1347 339 1348
rect 343 1347 344 1351
rect 358 1348 359 1352
rect 363 1348 364 1352
rect 358 1347 364 1348
rect 454 1351 461 1352
rect 454 1347 455 1351
rect 460 1347 461 1351
rect 582 1348 583 1352
rect 587 1348 588 1352
rect 582 1347 588 1348
rect 674 1351 685 1352
rect 674 1347 675 1351
rect 679 1347 680 1351
rect 684 1347 685 1351
rect 806 1348 807 1352
rect 811 1348 812 1352
rect 806 1347 812 1348
rect 902 1351 909 1352
rect 902 1347 903 1351
rect 908 1347 909 1351
rect 1030 1348 1031 1352
rect 1035 1348 1036 1352
rect 1030 1347 1036 1348
rect 1126 1351 1133 1352
rect 1126 1347 1127 1351
rect 1132 1347 1133 1351
rect 338 1346 344 1347
rect 454 1346 461 1347
rect 674 1346 685 1347
rect 902 1346 909 1347
rect 1126 1346 1133 1347
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 1934 1346 1940 1347
rect 1974 1351 1980 1352
rect 1974 1347 1975 1351
rect 1979 1347 1980 1351
rect 2126 1348 2127 1352
rect 2131 1348 2132 1352
rect 2126 1347 2132 1348
rect 2223 1351 2229 1352
rect 2223 1347 2224 1351
rect 2228 1350 2229 1351
rect 2250 1351 2256 1352
rect 2250 1350 2251 1351
rect 2228 1348 2251 1350
rect 2228 1347 2229 1348
rect 1974 1346 1980 1347
rect 2223 1346 2229 1347
rect 2250 1347 2251 1348
rect 2255 1347 2256 1351
rect 2270 1348 2271 1352
rect 2275 1348 2276 1352
rect 2270 1347 2276 1348
rect 2367 1351 2373 1352
rect 2367 1347 2368 1351
rect 2372 1350 2373 1351
rect 2394 1351 2400 1352
rect 2394 1350 2395 1351
rect 2372 1348 2395 1350
rect 2372 1347 2373 1348
rect 2250 1346 2256 1347
rect 2367 1346 2373 1347
rect 2394 1347 2395 1348
rect 2399 1347 2400 1351
rect 2414 1348 2415 1352
rect 2419 1348 2420 1352
rect 2414 1347 2420 1348
rect 2511 1351 2517 1352
rect 2511 1347 2512 1351
rect 2516 1350 2517 1351
rect 2546 1351 2552 1352
rect 2546 1350 2547 1351
rect 2516 1348 2547 1350
rect 2516 1347 2517 1348
rect 2394 1346 2400 1347
rect 2511 1346 2517 1347
rect 2546 1347 2547 1348
rect 2551 1347 2552 1351
rect 2566 1348 2567 1352
rect 2571 1348 2572 1352
rect 2566 1347 2572 1348
rect 2663 1351 2669 1352
rect 2663 1347 2664 1351
rect 2668 1350 2669 1351
rect 2698 1351 2704 1352
rect 2698 1350 2699 1351
rect 2668 1348 2699 1350
rect 2668 1347 2669 1348
rect 2546 1346 2552 1347
rect 2663 1346 2669 1347
rect 2698 1347 2699 1348
rect 2703 1347 2704 1351
rect 2718 1348 2719 1352
rect 2723 1348 2724 1352
rect 2718 1347 2724 1348
rect 2814 1351 2821 1352
rect 2814 1347 2815 1351
rect 2820 1347 2821 1351
rect 2878 1348 2879 1352
rect 2883 1348 2884 1352
rect 2878 1347 2884 1348
rect 2975 1351 2981 1352
rect 2975 1347 2976 1351
rect 2980 1350 2981 1351
rect 2983 1351 2989 1352
rect 2983 1350 2984 1351
rect 2980 1348 2984 1350
rect 2980 1347 2981 1348
rect 2698 1346 2704 1347
rect 2814 1346 2821 1347
rect 2975 1346 2981 1347
rect 2983 1347 2984 1348
rect 2988 1347 2989 1351
rect 3038 1348 3039 1352
rect 3043 1348 3044 1352
rect 3038 1347 3044 1348
rect 3135 1351 3141 1352
rect 3135 1347 3136 1351
rect 3140 1347 3141 1351
rect 3198 1348 3199 1352
rect 3203 1348 3204 1352
rect 3198 1347 3204 1348
rect 3295 1351 3301 1352
rect 3295 1347 3296 1351
rect 3300 1347 3301 1351
rect 2983 1346 2989 1347
rect 3135 1346 3141 1347
rect 3295 1346 3301 1347
rect 3798 1351 3804 1352
rect 3798 1347 3799 1351
rect 3803 1347 3804 1351
rect 3798 1346 3804 1347
rect 2194 1319 2200 1320
rect 2194 1315 2195 1319
rect 2199 1318 2200 1319
rect 2886 1319 2892 1320
rect 2886 1318 2887 1319
rect 2199 1316 2887 1318
rect 2199 1315 2200 1316
rect 2194 1314 2200 1315
rect 2886 1315 2887 1316
rect 2891 1315 2892 1319
rect 2886 1314 2892 1315
rect 3838 1301 3844 1302
rect 5662 1301 5668 1302
rect 3838 1297 3839 1301
rect 3843 1297 3844 1301
rect 3838 1296 3844 1297
rect 3886 1300 3892 1301
rect 4118 1300 4124 1301
rect 4390 1300 4396 1301
rect 4670 1300 4676 1301
rect 4966 1300 4972 1301
rect 5262 1300 5268 1301
rect 5542 1300 5548 1301
rect 3886 1296 3887 1300
rect 3891 1296 3892 1300
rect 3886 1295 3892 1296
rect 3982 1299 3989 1300
rect 3982 1295 3983 1299
rect 3988 1295 3989 1299
rect 4118 1296 4119 1300
rect 4123 1296 4124 1300
rect 4118 1295 4124 1296
rect 4215 1299 4224 1300
rect 4215 1295 4216 1299
rect 4223 1295 4224 1299
rect 4390 1296 4391 1300
rect 4395 1296 4396 1300
rect 4390 1295 4396 1296
rect 4487 1299 4496 1300
rect 4487 1295 4488 1299
rect 4495 1295 4496 1299
rect 4670 1296 4671 1300
rect 4675 1296 4676 1300
rect 4670 1295 4676 1296
rect 4766 1299 4773 1300
rect 4766 1295 4767 1299
rect 4772 1295 4773 1299
rect 4966 1296 4967 1300
rect 4971 1296 4972 1300
rect 4966 1295 4972 1296
rect 5063 1299 5072 1300
rect 5063 1295 5064 1299
rect 5071 1295 5072 1299
rect 5262 1296 5263 1300
rect 5267 1296 5268 1300
rect 5262 1295 5268 1296
rect 5354 1299 5365 1300
rect 5354 1295 5355 1299
rect 5359 1295 5360 1299
rect 5364 1295 5365 1299
rect 5542 1296 5543 1300
rect 5547 1296 5548 1300
rect 5542 1295 5548 1296
rect 5634 1299 5645 1300
rect 5634 1295 5635 1299
rect 5639 1295 5640 1299
rect 5644 1295 5645 1299
rect 5662 1297 5663 1301
rect 5667 1297 5668 1301
rect 5662 1296 5668 1297
rect 3982 1294 3989 1295
rect 4215 1294 4224 1295
rect 4487 1294 4496 1295
rect 4766 1294 4773 1295
rect 5063 1294 5072 1295
rect 5354 1294 5365 1295
rect 5634 1294 5645 1295
rect 110 1293 116 1294
rect 1934 1293 1940 1294
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 158 1292 164 1293
rect 366 1292 372 1293
rect 606 1292 612 1293
rect 846 1292 852 1293
rect 1086 1292 1092 1293
rect 158 1288 159 1292
rect 163 1288 164 1292
rect 158 1287 164 1288
rect 254 1291 261 1292
rect 254 1287 255 1291
rect 260 1287 261 1291
rect 366 1288 367 1292
rect 371 1288 372 1292
rect 366 1287 372 1288
rect 462 1291 469 1292
rect 462 1287 463 1291
rect 468 1287 469 1291
rect 606 1288 607 1292
rect 611 1288 612 1292
rect 606 1287 612 1288
rect 702 1291 709 1292
rect 702 1287 703 1291
rect 708 1287 709 1291
rect 846 1288 847 1292
rect 851 1288 852 1292
rect 846 1287 852 1288
rect 943 1291 949 1292
rect 943 1287 944 1291
rect 948 1290 949 1291
rect 970 1291 976 1292
rect 970 1290 971 1291
rect 948 1288 971 1290
rect 948 1287 949 1288
rect 254 1286 261 1287
rect 462 1286 469 1287
rect 702 1286 709 1287
rect 943 1286 949 1287
rect 970 1287 971 1288
rect 975 1287 976 1291
rect 1086 1288 1087 1292
rect 1091 1288 1092 1292
rect 1086 1287 1092 1288
rect 1178 1291 1189 1292
rect 1178 1287 1179 1291
rect 1183 1287 1184 1291
rect 1188 1287 1189 1291
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 1934 1288 1940 1289
rect 1974 1289 1980 1290
rect 3798 1289 3804 1290
rect 970 1286 976 1287
rect 1178 1286 1189 1287
rect 1974 1285 1975 1289
rect 1979 1285 1980 1289
rect 1974 1284 1980 1285
rect 2022 1288 2028 1289
rect 2174 1288 2180 1289
rect 2366 1288 2372 1289
rect 2574 1288 2580 1289
rect 2790 1288 2796 1289
rect 3014 1288 3020 1289
rect 3238 1288 3244 1289
rect 3470 1288 3476 1289
rect 3678 1288 3684 1289
rect 2022 1284 2023 1288
rect 2027 1284 2028 1288
rect 2022 1283 2028 1284
rect 2119 1287 2125 1288
rect 2119 1283 2120 1287
rect 2124 1286 2125 1287
rect 2135 1287 2141 1288
rect 2135 1286 2136 1287
rect 2124 1284 2136 1286
rect 2124 1283 2125 1284
rect 2119 1282 2125 1283
rect 2135 1283 2136 1284
rect 2140 1283 2141 1287
rect 2174 1284 2175 1288
rect 2179 1284 2180 1288
rect 2174 1283 2180 1284
rect 2271 1287 2277 1288
rect 2271 1283 2272 1287
rect 2276 1286 2277 1287
rect 2310 1287 2316 1288
rect 2310 1286 2311 1287
rect 2276 1284 2311 1286
rect 2276 1283 2277 1284
rect 2135 1282 2141 1283
rect 2271 1282 2277 1283
rect 2310 1283 2311 1284
rect 2315 1283 2316 1287
rect 2366 1284 2367 1288
rect 2371 1284 2372 1288
rect 2366 1283 2372 1284
rect 2463 1287 2472 1288
rect 2463 1283 2464 1287
rect 2471 1283 2472 1287
rect 2574 1284 2575 1288
rect 2579 1284 2580 1288
rect 2574 1283 2580 1284
rect 2671 1287 2680 1288
rect 2671 1283 2672 1287
rect 2679 1283 2680 1287
rect 2790 1284 2791 1288
rect 2795 1284 2796 1288
rect 2790 1283 2796 1284
rect 2886 1287 2893 1288
rect 2886 1283 2887 1287
rect 2892 1283 2893 1287
rect 3014 1284 3015 1288
rect 3019 1284 3020 1288
rect 3014 1283 3020 1284
rect 3111 1287 3120 1288
rect 3111 1283 3112 1287
rect 3119 1283 3120 1287
rect 3238 1284 3239 1288
rect 3243 1284 3244 1288
rect 3238 1283 3244 1284
rect 3334 1287 3341 1288
rect 3334 1283 3335 1287
rect 3340 1283 3341 1287
rect 3470 1284 3471 1288
rect 3475 1284 3476 1288
rect 3470 1283 3476 1284
rect 3567 1287 3573 1288
rect 3567 1283 3568 1287
rect 3572 1286 3573 1287
rect 3591 1287 3597 1288
rect 3591 1286 3592 1287
rect 3572 1284 3592 1286
rect 3572 1283 3573 1284
rect 2310 1282 2316 1283
rect 2463 1282 2472 1283
rect 2671 1282 2680 1283
rect 2886 1282 2893 1283
rect 3111 1282 3120 1283
rect 3334 1282 3341 1283
rect 3567 1282 3573 1283
rect 3591 1283 3592 1284
rect 3596 1283 3597 1287
rect 3678 1284 3679 1288
rect 3683 1284 3684 1288
rect 3678 1283 3684 1284
rect 3775 1287 3781 1288
rect 3775 1283 3776 1287
rect 3780 1286 3781 1287
rect 3790 1287 3796 1288
rect 3790 1286 3791 1287
rect 3780 1284 3791 1286
rect 3780 1283 3781 1284
rect 3591 1282 3597 1283
rect 3775 1282 3781 1283
rect 3790 1283 3791 1284
rect 3795 1283 3796 1287
rect 3798 1285 3799 1289
rect 3803 1285 3804 1289
rect 3858 1285 3864 1286
rect 3798 1284 3804 1285
rect 3838 1284 3844 1285
rect 3790 1282 3796 1283
rect 3838 1280 3839 1284
rect 3843 1280 3844 1284
rect 3858 1281 3859 1285
rect 3863 1281 3864 1285
rect 3858 1280 3864 1281
rect 4090 1285 4096 1286
rect 4090 1281 4091 1285
rect 4095 1281 4096 1285
rect 4090 1280 4096 1281
rect 4362 1285 4368 1286
rect 4362 1281 4363 1285
rect 4367 1281 4368 1285
rect 4362 1280 4368 1281
rect 4642 1285 4648 1286
rect 4642 1281 4643 1285
rect 4647 1281 4648 1285
rect 4642 1280 4648 1281
rect 4938 1285 4944 1286
rect 4938 1281 4939 1285
rect 4943 1281 4944 1285
rect 4938 1280 4944 1281
rect 5234 1285 5240 1286
rect 5234 1281 5235 1285
rect 5239 1281 5240 1285
rect 5234 1280 5240 1281
rect 5514 1285 5520 1286
rect 5514 1281 5515 1285
rect 5519 1281 5520 1285
rect 5514 1280 5520 1281
rect 5662 1284 5668 1285
rect 5662 1280 5663 1284
rect 5667 1280 5668 1284
rect 3838 1279 3844 1280
rect 5662 1279 5668 1280
rect 130 1277 136 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 130 1273 131 1277
rect 135 1273 136 1277
rect 130 1272 136 1273
rect 338 1277 344 1278
rect 338 1273 339 1277
rect 343 1273 344 1277
rect 338 1272 344 1273
rect 578 1277 584 1278
rect 578 1273 579 1277
rect 583 1273 584 1277
rect 578 1272 584 1273
rect 818 1277 824 1278
rect 818 1273 819 1277
rect 823 1273 824 1277
rect 818 1272 824 1273
rect 1058 1277 1064 1278
rect 1058 1273 1059 1277
rect 1063 1273 1064 1277
rect 1058 1272 1064 1273
rect 1934 1276 1940 1277
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 1994 1273 2000 1274
rect 110 1271 116 1272
rect 1934 1271 1940 1272
rect 1974 1272 1980 1273
rect 1974 1268 1975 1272
rect 1979 1268 1980 1272
rect 1994 1269 1995 1273
rect 1999 1269 2000 1273
rect 1994 1268 2000 1269
rect 2146 1273 2152 1274
rect 2146 1269 2147 1273
rect 2151 1269 2152 1273
rect 2146 1268 2152 1269
rect 2338 1273 2344 1274
rect 2338 1269 2339 1273
rect 2343 1269 2344 1273
rect 2338 1268 2344 1269
rect 2546 1273 2552 1274
rect 2546 1269 2547 1273
rect 2551 1269 2552 1273
rect 2546 1268 2552 1269
rect 2762 1273 2768 1274
rect 2762 1269 2763 1273
rect 2767 1269 2768 1273
rect 2762 1268 2768 1269
rect 2986 1273 2992 1274
rect 2986 1269 2987 1273
rect 2991 1269 2992 1273
rect 2986 1268 2992 1269
rect 3210 1273 3216 1274
rect 3210 1269 3211 1273
rect 3215 1269 3216 1273
rect 3210 1268 3216 1269
rect 3442 1273 3448 1274
rect 3442 1269 3443 1273
rect 3447 1269 3448 1273
rect 3442 1268 3448 1269
rect 3650 1273 3656 1274
rect 3650 1269 3651 1273
rect 3655 1269 3656 1273
rect 3650 1268 3656 1269
rect 3798 1272 3804 1273
rect 3798 1268 3799 1272
rect 3803 1268 3804 1272
rect 1974 1267 1980 1268
rect 3798 1267 3804 1268
rect 3790 1235 3796 1236
rect 3790 1231 3791 1235
rect 3795 1234 3796 1235
rect 4134 1235 4140 1236
rect 3795 1232 3865 1234
rect 3795 1231 3796 1232
rect 3790 1230 3796 1231
rect 4134 1231 4135 1235
rect 4139 1231 4140 1235
rect 4134 1230 4140 1231
rect 4218 1235 4224 1236
rect 4218 1231 4219 1235
rect 4223 1234 4224 1235
rect 4490 1235 4496 1236
rect 4223 1232 4369 1234
rect 4223 1231 4224 1232
rect 4218 1230 4224 1231
rect 4490 1231 4491 1235
rect 4495 1234 4496 1235
rect 5066 1235 5072 1236
rect 4495 1232 4649 1234
rect 4495 1231 4496 1232
rect 4490 1230 4496 1231
rect 250 1227 256 1228
rect 250 1226 251 1227
rect 229 1224 251 1226
rect 250 1223 251 1224
rect 255 1223 256 1227
rect 674 1227 680 1228
rect 250 1222 256 1223
rect 436 1218 438 1225
rect 674 1223 675 1227
rect 679 1223 680 1227
rect 674 1222 680 1223
rect 902 1227 908 1228
rect 902 1223 903 1227
rect 907 1223 908 1227
rect 902 1222 908 1223
rect 970 1227 976 1228
rect 970 1223 971 1227
rect 975 1226 976 1227
rect 5036 1226 5038 1233
rect 5066 1231 5067 1235
rect 5071 1234 5072 1235
rect 5647 1235 5653 1236
rect 5647 1234 5648 1235
rect 5071 1232 5241 1234
rect 5613 1232 5648 1234
rect 5071 1231 5072 1232
rect 5066 1230 5072 1231
rect 5647 1231 5648 1232
rect 5652 1231 5653 1235
rect 5647 1230 5653 1231
rect 5322 1227 5328 1228
rect 5322 1226 5323 1227
rect 975 1224 1065 1226
rect 5036 1224 5323 1226
rect 975 1223 976 1224
rect 970 1222 976 1223
rect 1914 1223 1920 1224
rect 702 1219 708 1220
rect 702 1218 703 1219
rect 436 1216 703 1218
rect 702 1215 703 1216
rect 707 1215 708 1219
rect 1914 1219 1915 1223
rect 1919 1222 1920 1223
rect 2135 1223 2141 1224
rect 1919 1220 2001 1222
rect 1919 1219 1920 1220
rect 1914 1218 1920 1219
rect 2135 1219 2136 1223
rect 2140 1222 2141 1223
rect 2310 1223 2316 1224
rect 2140 1220 2153 1222
rect 2140 1219 2141 1220
rect 2135 1218 2141 1219
rect 2310 1219 2311 1223
rect 2315 1222 2316 1223
rect 2466 1223 2472 1224
rect 2315 1220 2345 1222
rect 2315 1219 2316 1220
rect 2310 1218 2316 1219
rect 2466 1219 2467 1223
rect 2471 1222 2472 1223
rect 2674 1223 2680 1224
rect 2471 1220 2553 1222
rect 2471 1219 2472 1220
rect 2466 1218 2472 1219
rect 2674 1219 2675 1223
rect 2679 1222 2680 1223
rect 2983 1223 2989 1224
rect 2679 1220 2769 1222
rect 2679 1219 2680 1220
rect 2674 1218 2680 1219
rect 2983 1219 2984 1223
rect 2988 1222 2989 1223
rect 3114 1223 3120 1224
rect 2988 1220 2993 1222
rect 2988 1219 2989 1220
rect 2983 1218 2989 1219
rect 3114 1219 3115 1223
rect 3119 1222 3120 1223
rect 3582 1223 3588 1224
rect 3582 1222 3583 1223
rect 3119 1220 3217 1222
rect 3541 1220 3583 1222
rect 3119 1219 3120 1220
rect 3114 1218 3120 1219
rect 3582 1219 3583 1220
rect 3587 1219 3588 1223
rect 3582 1218 3588 1219
rect 3591 1223 3597 1224
rect 3591 1219 3592 1223
rect 3596 1222 3597 1223
rect 5322 1223 5323 1224
rect 5327 1223 5328 1227
rect 5322 1222 5328 1223
rect 3596 1220 3657 1222
rect 3596 1219 3597 1220
rect 3591 1218 3597 1219
rect 702 1214 708 1215
rect 1178 1191 1184 1192
rect 1178 1190 1179 1191
rect 1024 1188 1179 1190
rect 266 1183 272 1184
rect 266 1182 267 1183
rect 229 1180 267 1182
rect 266 1179 267 1180
rect 271 1179 272 1183
rect 462 1183 468 1184
rect 266 1178 272 1179
rect 370 1179 376 1180
rect 370 1175 371 1179
rect 375 1175 376 1179
rect 462 1179 463 1183
rect 467 1179 468 1183
rect 914 1183 920 1184
rect 914 1182 915 1183
rect 861 1180 915 1182
rect 462 1178 468 1179
rect 610 1179 616 1180
rect 370 1174 376 1175
rect 610 1175 611 1179
rect 615 1175 616 1179
rect 914 1179 915 1180
rect 919 1179 920 1183
rect 1024 1182 1026 1188
rect 1178 1187 1179 1188
rect 1183 1187 1184 1191
rect 1178 1186 1184 1187
rect 1334 1187 1340 1188
rect 1334 1186 1335 1187
rect 1216 1184 1335 1186
rect 1216 1182 1218 1184
rect 1334 1183 1335 1184
rect 1339 1183 1340 1187
rect 4334 1187 4340 1188
rect 4334 1186 4335 1187
rect 4172 1184 4335 1186
rect 1334 1182 1340 1183
rect 3239 1183 3245 1184
rect 3239 1182 3240 1183
rect 1021 1180 1026 1182
rect 1173 1180 1218 1182
rect 3181 1180 3240 1182
rect 914 1178 920 1179
rect 1226 1179 1232 1180
rect 610 1174 616 1175
rect 1226 1175 1227 1179
rect 1231 1175 1232 1179
rect 1226 1174 1232 1175
rect 1370 1179 1376 1180
rect 1370 1175 1371 1179
rect 1375 1175 1376 1179
rect 1370 1174 1376 1175
rect 1514 1179 1520 1180
rect 1514 1175 1515 1179
rect 1519 1175 1520 1179
rect 1514 1174 1520 1175
rect 1658 1179 1664 1180
rect 1658 1175 1659 1179
rect 1663 1175 1664 1179
rect 1658 1174 1664 1175
rect 1794 1179 1800 1180
rect 1794 1175 1795 1179
rect 1799 1175 1800 1179
rect 1794 1174 1800 1175
rect 2818 1179 2824 1180
rect 2818 1175 2819 1179
rect 2823 1175 2824 1179
rect 2818 1174 2824 1175
rect 2906 1179 2912 1180
rect 2906 1175 2907 1179
rect 2911 1175 2912 1179
rect 3239 1179 3240 1180
rect 3244 1179 3245 1183
rect 3239 1178 3245 1179
rect 3334 1183 3340 1184
rect 3334 1179 3335 1183
rect 3339 1179 3340 1183
rect 3642 1183 3648 1184
rect 3642 1182 3643 1183
rect 3565 1180 3643 1182
rect 3334 1178 3340 1179
rect 3642 1179 3643 1180
rect 3647 1179 3648 1183
rect 3642 1178 3648 1179
rect 3670 1183 3676 1184
rect 3670 1179 3671 1183
rect 3675 1179 3676 1183
rect 4172 1182 4174 1184
rect 4334 1183 4335 1184
rect 4339 1183 4340 1187
rect 4334 1182 4340 1183
rect 4682 1183 4688 1184
rect 4682 1182 4683 1183
rect 4109 1180 4174 1182
rect 4533 1180 4683 1182
rect 3670 1178 3676 1179
rect 4218 1179 4224 1180
rect 2906 1174 2912 1175
rect 4218 1175 4219 1179
rect 4223 1175 4224 1179
rect 4682 1179 4683 1180
rect 4687 1179 4688 1183
rect 4682 1178 4688 1179
rect 4766 1183 4772 1184
rect 4766 1179 4767 1183
rect 4771 1179 4772 1183
rect 5354 1183 5360 1184
rect 5354 1182 5355 1183
rect 5349 1180 5355 1182
rect 4766 1178 4772 1179
rect 4970 1179 4976 1180
rect 4218 1174 4224 1175
rect 4970 1175 4971 1179
rect 4975 1175 4976 1179
rect 5354 1179 5355 1180
rect 5359 1179 5360 1183
rect 5634 1183 5640 1184
rect 5634 1182 5635 1183
rect 5613 1180 5635 1182
rect 5354 1178 5360 1179
rect 5634 1179 5635 1180
rect 5639 1179 5640 1183
rect 5634 1178 5640 1179
rect 4970 1174 4976 1175
rect 2818 1159 2824 1160
rect 370 1155 376 1156
rect 370 1151 371 1155
rect 375 1154 376 1155
rect 726 1155 732 1156
rect 726 1154 727 1155
rect 375 1152 727 1154
rect 375 1151 376 1152
rect 370 1150 376 1151
rect 726 1151 727 1152
rect 731 1151 732 1155
rect 2818 1155 2819 1159
rect 2823 1158 2824 1159
rect 3202 1159 3208 1160
rect 3202 1158 3203 1159
rect 2823 1156 3203 1158
rect 2823 1155 2824 1156
rect 2818 1154 2824 1155
rect 3202 1155 3203 1156
rect 3207 1155 3208 1159
rect 3202 1154 3208 1155
rect 726 1150 732 1151
rect 110 1132 116 1133
rect 1934 1132 1940 1133
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 130 1131 136 1132
rect 130 1127 131 1131
rect 135 1127 136 1131
rect 130 1126 136 1127
rect 274 1131 280 1132
rect 274 1127 275 1131
rect 279 1127 280 1131
rect 274 1126 280 1127
rect 442 1131 448 1132
rect 442 1127 443 1131
rect 447 1127 448 1131
rect 442 1126 448 1127
rect 602 1131 608 1132
rect 602 1127 603 1131
rect 607 1127 608 1131
rect 602 1126 608 1127
rect 762 1131 768 1132
rect 762 1127 763 1131
rect 767 1127 768 1131
rect 762 1126 768 1127
rect 922 1131 928 1132
rect 922 1127 923 1131
rect 927 1127 928 1131
rect 922 1126 928 1127
rect 1074 1131 1080 1132
rect 1074 1127 1075 1131
rect 1079 1127 1080 1131
rect 1074 1126 1080 1127
rect 1218 1131 1224 1132
rect 1218 1127 1219 1131
rect 1223 1127 1224 1131
rect 1218 1126 1224 1127
rect 1362 1131 1368 1132
rect 1362 1127 1363 1131
rect 1367 1127 1368 1131
rect 1362 1126 1368 1127
rect 1506 1131 1512 1132
rect 1506 1127 1507 1131
rect 1511 1127 1512 1131
rect 1506 1126 1512 1127
rect 1650 1131 1656 1132
rect 1650 1127 1651 1131
rect 1655 1127 1656 1131
rect 1650 1126 1656 1127
rect 1786 1131 1792 1132
rect 1786 1127 1787 1131
rect 1791 1127 1792 1131
rect 1934 1128 1935 1132
rect 1939 1128 1940 1132
rect 1934 1127 1940 1128
rect 1974 1132 1980 1133
rect 3798 1132 3804 1133
rect 1974 1128 1975 1132
rect 1979 1128 1980 1132
rect 1974 1127 1980 1128
rect 2722 1131 2728 1132
rect 2722 1127 2723 1131
rect 2727 1127 2728 1131
rect 1786 1126 1792 1127
rect 2722 1126 2728 1127
rect 2898 1131 2904 1132
rect 2898 1127 2899 1131
rect 2903 1127 2904 1131
rect 2898 1126 2904 1127
rect 3082 1131 3088 1132
rect 3082 1127 3083 1131
rect 3087 1127 3088 1131
rect 3082 1126 3088 1127
rect 3274 1131 3280 1132
rect 3274 1127 3275 1131
rect 3279 1127 3280 1131
rect 3274 1126 3280 1127
rect 3466 1131 3472 1132
rect 3466 1127 3467 1131
rect 3471 1127 3472 1131
rect 3466 1126 3472 1127
rect 3650 1131 3656 1132
rect 3650 1127 3651 1131
rect 3655 1127 3656 1131
rect 3798 1128 3799 1132
rect 3803 1128 3804 1132
rect 3798 1127 3804 1128
rect 3838 1132 3844 1133
rect 5662 1132 5668 1133
rect 3838 1128 3839 1132
rect 3843 1128 3844 1132
rect 3838 1127 3844 1128
rect 4010 1131 4016 1132
rect 4010 1127 4011 1131
rect 4015 1127 4016 1131
rect 3650 1126 3656 1127
rect 4010 1126 4016 1127
rect 4210 1131 4216 1132
rect 4210 1127 4211 1131
rect 4215 1127 4216 1131
rect 4210 1126 4216 1127
rect 4434 1131 4440 1132
rect 4434 1127 4435 1131
rect 4439 1127 4440 1131
rect 4434 1126 4440 1127
rect 4690 1131 4696 1132
rect 4690 1127 4691 1131
rect 4695 1127 4696 1131
rect 4690 1126 4696 1127
rect 4962 1131 4968 1132
rect 4962 1127 4963 1131
rect 4967 1127 4968 1131
rect 4962 1126 4968 1127
rect 5250 1131 5256 1132
rect 5250 1127 5251 1131
rect 5255 1127 5256 1131
rect 5250 1126 5256 1127
rect 5514 1131 5520 1132
rect 5514 1127 5515 1131
rect 5519 1127 5520 1131
rect 5662 1128 5663 1132
rect 5667 1128 5668 1132
rect 5662 1127 5668 1128
rect 5514 1126 5520 1127
rect 914 1123 920 1124
rect 914 1119 915 1123
rect 919 1122 920 1123
rect 3239 1123 3245 1124
rect 919 1120 1050 1122
rect 919 1119 920 1120
rect 914 1118 920 1119
rect 1048 1118 1050 1120
rect 3239 1119 3240 1123
rect 3244 1122 3245 1123
rect 3642 1123 3648 1124
rect 3244 1120 3402 1122
rect 3244 1119 3245 1120
rect 3239 1118 3245 1119
rect 1047 1117 1053 1118
rect 158 1116 164 1117
rect 302 1116 308 1117
rect 470 1116 476 1117
rect 630 1116 636 1117
rect 790 1116 796 1117
rect 950 1116 956 1117
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 158 1112 159 1116
rect 163 1112 164 1116
rect 158 1111 164 1112
rect 250 1115 261 1116
rect 250 1111 251 1115
rect 255 1111 256 1115
rect 260 1111 261 1115
rect 302 1112 303 1116
rect 307 1112 308 1116
rect 302 1111 308 1112
rect 398 1115 405 1116
rect 398 1111 399 1115
rect 404 1111 405 1115
rect 470 1112 471 1116
rect 475 1112 476 1116
rect 470 1111 476 1112
rect 567 1115 573 1116
rect 567 1111 568 1115
rect 572 1114 573 1115
rect 610 1115 616 1116
rect 610 1114 611 1115
rect 572 1112 611 1114
rect 572 1111 573 1112
rect 110 1110 116 1111
rect 250 1110 261 1111
rect 398 1110 405 1111
rect 567 1110 573 1111
rect 610 1111 611 1112
rect 615 1111 616 1115
rect 630 1112 631 1116
rect 635 1112 636 1116
rect 630 1111 636 1112
rect 726 1115 733 1116
rect 726 1111 727 1115
rect 732 1111 733 1115
rect 790 1112 791 1116
rect 795 1112 796 1116
rect 790 1111 796 1112
rect 886 1115 893 1116
rect 886 1111 887 1115
rect 892 1111 893 1115
rect 950 1112 951 1116
rect 955 1112 956 1116
rect 1047 1113 1048 1117
rect 1052 1113 1053 1117
rect 1047 1112 1053 1113
rect 1102 1116 1108 1117
rect 1246 1116 1252 1117
rect 1390 1116 1396 1117
rect 1534 1116 1540 1117
rect 1678 1116 1684 1117
rect 1814 1116 1820 1117
rect 2750 1116 2756 1117
rect 2926 1116 2932 1117
rect 3110 1116 3116 1117
rect 3302 1116 3308 1117
rect 3400 1116 3402 1120
rect 3642 1119 3643 1123
rect 3647 1122 3648 1123
rect 4682 1123 4688 1124
rect 3647 1120 3778 1122
rect 3647 1119 3648 1120
rect 3642 1118 3648 1119
rect 3494 1116 3500 1117
rect 3678 1116 3684 1117
rect 3776 1116 3778 1120
rect 4682 1119 4683 1123
rect 4687 1122 4688 1123
rect 4687 1120 5090 1122
rect 4687 1119 4688 1120
rect 4682 1118 4688 1119
rect 4038 1116 4044 1117
rect 4238 1116 4244 1117
rect 4462 1116 4468 1117
rect 4718 1116 4724 1117
rect 4990 1116 4996 1117
rect 5088 1116 5090 1120
rect 5278 1116 5284 1117
rect 5542 1116 5548 1117
rect 1102 1112 1103 1116
rect 1107 1112 1108 1116
rect 950 1111 956 1112
rect 1102 1111 1108 1112
rect 1199 1115 1205 1116
rect 1199 1111 1200 1115
rect 1204 1114 1205 1115
rect 1226 1115 1232 1116
rect 1226 1114 1227 1115
rect 1204 1112 1227 1114
rect 1204 1111 1205 1112
rect 610 1110 616 1111
rect 726 1110 733 1111
rect 886 1110 893 1111
rect 1199 1110 1205 1111
rect 1226 1111 1227 1112
rect 1231 1111 1232 1115
rect 1246 1112 1247 1116
rect 1251 1112 1252 1116
rect 1246 1111 1252 1112
rect 1343 1115 1349 1116
rect 1343 1111 1344 1115
rect 1348 1114 1349 1115
rect 1370 1115 1376 1116
rect 1370 1114 1371 1115
rect 1348 1112 1371 1114
rect 1348 1111 1349 1112
rect 1226 1110 1232 1111
rect 1343 1110 1349 1111
rect 1370 1111 1371 1112
rect 1375 1111 1376 1115
rect 1390 1112 1391 1116
rect 1395 1112 1396 1116
rect 1390 1111 1396 1112
rect 1487 1115 1493 1116
rect 1487 1111 1488 1115
rect 1492 1114 1493 1115
rect 1514 1115 1520 1116
rect 1514 1114 1515 1115
rect 1492 1112 1515 1114
rect 1492 1111 1493 1112
rect 1370 1110 1376 1111
rect 1487 1110 1493 1111
rect 1514 1111 1515 1112
rect 1519 1111 1520 1115
rect 1534 1112 1535 1116
rect 1539 1112 1540 1116
rect 1534 1111 1540 1112
rect 1631 1115 1637 1116
rect 1631 1111 1632 1115
rect 1636 1114 1637 1115
rect 1658 1115 1664 1116
rect 1658 1114 1659 1115
rect 1636 1112 1659 1114
rect 1636 1111 1637 1112
rect 1514 1110 1520 1111
rect 1631 1110 1637 1111
rect 1658 1111 1659 1112
rect 1663 1111 1664 1115
rect 1678 1112 1679 1116
rect 1683 1112 1684 1116
rect 1678 1111 1684 1112
rect 1775 1115 1781 1116
rect 1775 1111 1776 1115
rect 1780 1114 1781 1115
rect 1794 1115 1800 1116
rect 1794 1114 1795 1115
rect 1780 1112 1795 1114
rect 1780 1111 1781 1112
rect 1658 1110 1664 1111
rect 1775 1110 1781 1111
rect 1794 1111 1795 1112
rect 1799 1111 1800 1115
rect 1814 1112 1815 1116
rect 1819 1112 1820 1116
rect 1814 1111 1820 1112
rect 1911 1115 1920 1116
rect 1911 1111 1912 1115
rect 1919 1111 1920 1115
rect 1794 1110 1800 1111
rect 1911 1110 1920 1111
rect 1934 1115 1940 1116
rect 1934 1111 1935 1115
rect 1939 1111 1940 1115
rect 1934 1110 1940 1111
rect 1974 1115 1980 1116
rect 1974 1111 1975 1115
rect 1979 1111 1980 1115
rect 2750 1112 2751 1116
rect 2755 1112 2756 1116
rect 2750 1111 2756 1112
rect 2847 1115 2853 1116
rect 2847 1111 2848 1115
rect 2852 1114 2853 1115
rect 2906 1115 2912 1116
rect 2906 1114 2907 1115
rect 2852 1112 2907 1114
rect 2852 1111 2853 1112
rect 1974 1110 1980 1111
rect 2847 1110 2853 1111
rect 2906 1111 2907 1112
rect 2911 1111 2912 1115
rect 2926 1112 2927 1116
rect 2931 1112 2932 1116
rect 2926 1111 2932 1112
rect 3018 1115 3029 1116
rect 3018 1111 3019 1115
rect 3023 1111 3024 1115
rect 3028 1111 3029 1115
rect 3110 1112 3111 1116
rect 3115 1112 3116 1116
rect 3110 1111 3116 1112
rect 3202 1115 3213 1116
rect 3202 1111 3203 1115
rect 3207 1111 3208 1115
rect 3212 1111 3213 1115
rect 3302 1112 3303 1116
rect 3307 1112 3308 1116
rect 3302 1111 3308 1112
rect 3399 1115 3405 1116
rect 3399 1111 3400 1115
rect 3404 1111 3405 1115
rect 3494 1112 3495 1116
rect 3499 1112 3500 1116
rect 3494 1111 3500 1112
rect 3586 1115 3597 1116
rect 3586 1111 3587 1115
rect 3591 1111 3592 1115
rect 3596 1111 3597 1115
rect 3678 1112 3679 1116
rect 3683 1112 3684 1116
rect 3678 1111 3684 1112
rect 3775 1115 3781 1116
rect 3775 1111 3776 1115
rect 3780 1111 3781 1115
rect 2906 1110 2912 1111
rect 3018 1110 3029 1111
rect 3202 1110 3213 1111
rect 3399 1110 3405 1111
rect 3586 1110 3597 1111
rect 3775 1110 3781 1111
rect 3798 1115 3804 1116
rect 3798 1111 3799 1115
rect 3803 1111 3804 1115
rect 3798 1110 3804 1111
rect 3838 1115 3844 1116
rect 3838 1111 3839 1115
rect 3843 1111 3844 1115
rect 4038 1112 4039 1116
rect 4043 1112 4044 1116
rect 4038 1111 4044 1112
rect 4134 1115 4141 1116
rect 4134 1111 4135 1115
rect 4140 1111 4141 1115
rect 4238 1112 4239 1116
rect 4243 1112 4244 1116
rect 4238 1111 4244 1112
rect 4334 1115 4341 1116
rect 4334 1111 4335 1115
rect 4340 1111 4341 1115
rect 4462 1112 4463 1116
rect 4467 1112 4468 1116
rect 4462 1111 4468 1112
rect 4559 1115 4565 1116
rect 4559 1111 4560 1115
rect 4564 1114 4565 1115
rect 4578 1115 4584 1116
rect 4578 1114 4579 1115
rect 4564 1112 4579 1114
rect 4564 1111 4565 1112
rect 3838 1110 3844 1111
rect 4134 1110 4141 1111
rect 4334 1110 4341 1111
rect 4559 1110 4565 1111
rect 4578 1111 4579 1112
rect 4583 1111 4584 1115
rect 4718 1112 4719 1116
rect 4723 1112 4724 1116
rect 4718 1111 4724 1112
rect 4815 1115 4821 1116
rect 4815 1111 4816 1115
rect 4820 1114 4821 1115
rect 4970 1115 4976 1116
rect 4970 1114 4971 1115
rect 4820 1112 4971 1114
rect 4820 1111 4821 1112
rect 4578 1110 4584 1111
rect 4815 1110 4821 1111
rect 4970 1111 4971 1112
rect 4975 1111 4976 1115
rect 4990 1112 4991 1116
rect 4995 1112 4996 1116
rect 4990 1111 4996 1112
rect 5087 1115 5093 1116
rect 5087 1111 5088 1115
rect 5092 1111 5093 1115
rect 5278 1112 5279 1116
rect 5283 1112 5284 1116
rect 5278 1111 5284 1112
rect 5374 1115 5381 1116
rect 5374 1111 5375 1115
rect 5380 1111 5381 1115
rect 5542 1112 5543 1116
rect 5547 1112 5548 1116
rect 5542 1111 5548 1112
rect 5638 1115 5645 1116
rect 5638 1111 5639 1115
rect 5644 1111 5645 1115
rect 4970 1110 4976 1111
rect 5087 1110 5093 1111
rect 5374 1110 5381 1111
rect 5638 1110 5645 1111
rect 5662 1115 5668 1116
rect 5662 1111 5663 1115
rect 5667 1111 5668 1115
rect 5662 1110 5668 1111
rect 110 1049 116 1050
rect 1934 1049 1940 1050
rect 110 1045 111 1049
rect 115 1045 116 1049
rect 110 1044 116 1045
rect 174 1048 180 1049
rect 414 1048 420 1049
rect 638 1048 644 1049
rect 854 1048 860 1049
rect 1054 1048 1060 1049
rect 1238 1048 1244 1049
rect 1422 1048 1428 1049
rect 1606 1048 1612 1049
rect 1790 1048 1796 1049
rect 174 1044 175 1048
rect 179 1044 180 1048
rect 174 1043 180 1044
rect 266 1047 277 1048
rect 266 1043 267 1047
rect 271 1043 272 1047
rect 276 1043 277 1047
rect 414 1044 415 1048
rect 419 1044 420 1048
rect 414 1043 420 1044
rect 511 1047 520 1048
rect 511 1043 512 1047
rect 519 1043 520 1047
rect 638 1044 639 1048
rect 643 1044 644 1048
rect 638 1043 644 1044
rect 734 1047 741 1048
rect 734 1043 735 1047
rect 740 1043 741 1047
rect 854 1044 855 1048
rect 859 1044 860 1048
rect 854 1043 860 1044
rect 951 1047 960 1048
rect 951 1043 952 1047
rect 959 1043 960 1047
rect 1054 1044 1055 1048
rect 1059 1044 1060 1048
rect 1054 1043 1060 1044
rect 1151 1047 1160 1048
rect 1151 1043 1152 1047
rect 1159 1043 1160 1047
rect 1238 1044 1239 1048
rect 1243 1044 1244 1048
rect 1238 1043 1244 1044
rect 1334 1047 1341 1048
rect 1334 1043 1335 1047
rect 1340 1043 1341 1047
rect 1422 1044 1423 1048
rect 1427 1044 1428 1048
rect 1422 1043 1428 1044
rect 1518 1047 1525 1048
rect 1518 1043 1519 1047
rect 1524 1043 1525 1047
rect 1606 1044 1607 1048
rect 1611 1044 1612 1048
rect 1606 1043 1612 1044
rect 1702 1047 1709 1048
rect 1702 1043 1703 1047
rect 1708 1043 1709 1047
rect 1790 1044 1791 1048
rect 1795 1044 1796 1048
rect 1790 1043 1796 1044
rect 1886 1047 1893 1048
rect 1886 1043 1887 1047
rect 1892 1043 1893 1047
rect 1934 1045 1935 1049
rect 1939 1045 1940 1049
rect 1934 1044 1940 1045
rect 1974 1045 1980 1046
rect 3798 1045 3804 1046
rect 266 1042 277 1043
rect 511 1042 520 1043
rect 734 1042 741 1043
rect 951 1042 960 1043
rect 1151 1042 1160 1043
rect 1334 1042 1341 1043
rect 1518 1042 1525 1043
rect 1702 1042 1709 1043
rect 1886 1042 1893 1043
rect 1974 1041 1975 1045
rect 1979 1041 1980 1045
rect 1974 1040 1980 1041
rect 2558 1044 2564 1045
rect 2750 1044 2756 1045
rect 2950 1044 2956 1045
rect 3150 1044 3156 1045
rect 3358 1044 3364 1045
rect 3574 1044 3580 1045
rect 2558 1040 2559 1044
rect 2563 1040 2564 1044
rect 2558 1039 2564 1040
rect 2650 1043 2661 1044
rect 2650 1039 2651 1043
rect 2655 1039 2656 1043
rect 2660 1039 2661 1043
rect 2750 1040 2751 1044
rect 2755 1040 2756 1044
rect 2750 1039 2756 1040
rect 2842 1043 2853 1044
rect 2842 1039 2843 1043
rect 2847 1039 2848 1043
rect 2852 1039 2853 1043
rect 2950 1040 2951 1044
rect 2955 1040 2956 1044
rect 2950 1039 2956 1040
rect 3047 1043 3056 1044
rect 3047 1039 3048 1043
rect 3055 1039 3056 1043
rect 3150 1040 3151 1044
rect 3155 1040 3156 1044
rect 3150 1039 3156 1040
rect 3242 1043 3253 1044
rect 3242 1039 3243 1043
rect 3247 1039 3248 1043
rect 3252 1039 3253 1043
rect 3358 1040 3359 1044
rect 3363 1040 3364 1044
rect 3358 1039 3364 1040
rect 3455 1043 3464 1044
rect 3455 1039 3456 1043
rect 3463 1039 3464 1043
rect 3574 1040 3575 1044
rect 3579 1040 3580 1044
rect 3574 1039 3580 1040
rect 3670 1043 3677 1044
rect 3670 1039 3671 1043
rect 3676 1039 3677 1043
rect 3798 1041 3799 1045
rect 3803 1041 3804 1045
rect 3798 1040 3804 1041
rect 3838 1045 3844 1046
rect 5639 1045 5645 1046
rect 3838 1041 3839 1045
rect 3843 1041 3844 1045
rect 3838 1040 3844 1041
rect 4094 1044 4100 1045
rect 4390 1044 4396 1045
rect 4686 1044 4692 1045
rect 4974 1044 4980 1045
rect 5262 1044 5268 1045
rect 5542 1044 5548 1045
rect 4094 1040 4095 1044
rect 4099 1040 4100 1044
rect 4094 1039 4100 1040
rect 4191 1043 4197 1044
rect 4191 1039 4192 1043
rect 4196 1042 4197 1043
rect 4218 1043 4224 1044
rect 4218 1042 4219 1043
rect 4196 1040 4219 1042
rect 4196 1039 4197 1040
rect 2650 1038 2661 1039
rect 2842 1038 2853 1039
rect 3047 1038 3056 1039
rect 3242 1038 3253 1039
rect 3455 1038 3464 1039
rect 3670 1038 3677 1039
rect 4191 1038 4197 1039
rect 4218 1039 4219 1040
rect 4223 1039 4224 1043
rect 4390 1040 4391 1044
rect 4395 1040 4396 1044
rect 4390 1039 4396 1040
rect 4482 1043 4493 1044
rect 4482 1039 4483 1043
rect 4487 1039 4488 1043
rect 4492 1039 4493 1043
rect 4686 1040 4687 1044
rect 4691 1040 4692 1044
rect 4686 1039 4692 1040
rect 4778 1043 4789 1044
rect 4778 1039 4779 1043
rect 4783 1039 4784 1043
rect 4788 1039 4789 1043
rect 4974 1040 4975 1044
rect 4979 1040 4980 1044
rect 4974 1039 4980 1040
rect 5071 1043 5080 1044
rect 5071 1039 5072 1043
rect 5079 1039 5080 1043
rect 5262 1040 5263 1044
rect 5267 1040 5268 1044
rect 5262 1039 5268 1040
rect 5354 1043 5365 1044
rect 5354 1039 5355 1043
rect 5359 1039 5360 1043
rect 5364 1039 5365 1043
rect 5542 1040 5543 1044
rect 5547 1040 5548 1044
rect 5639 1041 5640 1045
rect 5644 1041 5645 1045
rect 5639 1040 5645 1041
rect 5662 1045 5668 1046
rect 5662 1041 5663 1045
rect 5667 1041 5668 1045
rect 5662 1040 5668 1041
rect 5542 1039 5548 1040
rect 4218 1038 4224 1039
rect 4482 1038 4493 1039
rect 4778 1038 4789 1039
rect 5071 1038 5080 1039
rect 5354 1038 5365 1039
rect 5640 1034 5642 1040
rect 5646 1035 5652 1036
rect 5646 1034 5647 1035
rect 146 1033 152 1034
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 146 1029 147 1033
rect 151 1029 152 1033
rect 146 1028 152 1029
rect 386 1033 392 1034
rect 386 1029 387 1033
rect 391 1029 392 1033
rect 386 1028 392 1029
rect 610 1033 616 1034
rect 610 1029 611 1033
rect 615 1029 616 1033
rect 610 1028 616 1029
rect 826 1033 832 1034
rect 826 1029 827 1033
rect 831 1029 832 1033
rect 826 1028 832 1029
rect 1026 1033 1032 1034
rect 1026 1029 1027 1033
rect 1031 1029 1032 1033
rect 1026 1028 1032 1029
rect 1210 1033 1216 1034
rect 1210 1029 1211 1033
rect 1215 1029 1216 1033
rect 1210 1028 1216 1029
rect 1394 1033 1400 1034
rect 1394 1029 1395 1033
rect 1399 1029 1400 1033
rect 1394 1028 1400 1029
rect 1578 1033 1584 1034
rect 1578 1029 1579 1033
rect 1583 1029 1584 1033
rect 1578 1028 1584 1029
rect 1762 1033 1768 1034
rect 1762 1029 1763 1033
rect 1767 1029 1768 1033
rect 1762 1028 1768 1029
rect 1934 1032 1940 1033
rect 5640 1032 5647 1034
rect 1934 1028 1935 1032
rect 1939 1028 1940 1032
rect 5646 1031 5647 1032
rect 5651 1031 5652 1035
rect 5646 1030 5652 1031
rect 2530 1029 2536 1030
rect 110 1027 116 1028
rect 1934 1027 1940 1028
rect 1974 1028 1980 1029
rect 1974 1024 1975 1028
rect 1979 1024 1980 1028
rect 2530 1025 2531 1029
rect 2535 1025 2536 1029
rect 2530 1024 2536 1025
rect 2722 1029 2728 1030
rect 2722 1025 2723 1029
rect 2727 1025 2728 1029
rect 2722 1024 2728 1025
rect 2922 1029 2928 1030
rect 2922 1025 2923 1029
rect 2927 1025 2928 1029
rect 2922 1024 2928 1025
rect 3122 1029 3128 1030
rect 3122 1025 3123 1029
rect 3127 1025 3128 1029
rect 3122 1024 3128 1025
rect 3330 1029 3336 1030
rect 3330 1025 3331 1029
rect 3335 1025 3336 1029
rect 3330 1024 3336 1025
rect 3546 1029 3552 1030
rect 4066 1029 4072 1030
rect 3546 1025 3547 1029
rect 3551 1025 3552 1029
rect 3546 1024 3552 1025
rect 3798 1028 3804 1029
rect 3798 1024 3799 1028
rect 3803 1024 3804 1028
rect 1974 1023 1980 1024
rect 3798 1023 3804 1024
rect 3838 1028 3844 1029
rect 3838 1024 3839 1028
rect 3843 1024 3844 1028
rect 4066 1025 4067 1029
rect 4071 1025 4072 1029
rect 4066 1024 4072 1025
rect 4362 1029 4368 1030
rect 4362 1025 4363 1029
rect 4367 1025 4368 1029
rect 4362 1024 4368 1025
rect 4658 1029 4664 1030
rect 4658 1025 4659 1029
rect 4663 1025 4664 1029
rect 4658 1024 4664 1025
rect 4946 1029 4952 1030
rect 4946 1025 4947 1029
rect 4951 1025 4952 1029
rect 4946 1024 4952 1025
rect 5234 1029 5240 1030
rect 5234 1025 5235 1029
rect 5239 1025 5240 1029
rect 5234 1024 5240 1025
rect 5514 1029 5520 1030
rect 5514 1025 5515 1029
rect 5519 1025 5520 1029
rect 5514 1024 5520 1025
rect 5662 1028 5668 1029
rect 5662 1024 5663 1028
rect 5667 1024 5668 1028
rect 3838 1023 3844 1024
rect 5662 1023 5668 1024
rect 1490 1011 1496 1012
rect 1490 1007 1491 1011
rect 1495 1010 1496 1011
rect 1702 1011 1708 1012
rect 1702 1010 1703 1011
rect 1495 1008 1703 1010
rect 1495 1007 1496 1008
rect 1490 1006 1496 1007
rect 1702 1007 1703 1008
rect 1707 1007 1708 1011
rect 1702 1006 1708 1007
rect 2626 1011 2632 1012
rect 2626 1007 2627 1011
rect 2631 1010 2632 1011
rect 2842 1011 2848 1012
rect 2842 1010 2843 1011
rect 2631 1008 2843 1010
rect 2631 1007 2632 1008
rect 2626 1006 2632 1007
rect 2842 1007 2843 1008
rect 2847 1007 2848 1011
rect 2842 1006 2848 1007
rect 318 983 324 984
rect 318 982 319 983
rect 245 980 319 982
rect 318 979 319 980
rect 323 979 324 983
rect 318 978 324 979
rect 398 983 404 984
rect 398 979 399 983
rect 403 979 404 983
rect 398 978 404 979
rect 514 983 520 984
rect 514 979 515 983
rect 519 982 520 983
rect 886 983 892 984
rect 519 980 617 982
rect 519 979 520 980
rect 514 978 520 979
rect 886 979 887 983
rect 891 979 892 983
rect 886 978 892 979
rect 954 983 960 984
rect 954 979 955 983
rect 959 982 960 983
rect 1490 983 1496 984
rect 959 980 1033 982
rect 959 979 960 980
rect 954 978 960 979
rect 1308 974 1310 981
rect 1490 979 1491 983
rect 1495 979 1496 983
rect 1906 983 1912 984
rect 1906 982 1907 983
rect 1490 978 1496 979
rect 1518 975 1524 976
rect 1518 974 1519 975
rect 1308 972 1519 974
rect 1518 971 1519 972
rect 1523 971 1524 975
rect 1676 974 1678 981
rect 1861 980 1907 982
rect 1906 979 1907 980
rect 1911 979 1912 983
rect 1906 978 1912 979
rect 2626 979 2632 980
rect 1886 975 1892 976
rect 1886 974 1887 975
rect 1676 972 1887 974
rect 1518 970 1524 971
rect 1886 971 1887 972
rect 1891 971 1892 975
rect 2626 975 2627 979
rect 2631 975 2632 979
rect 3018 979 3024 980
rect 2626 974 2632 975
rect 1886 970 1892 971
rect 2820 970 2822 977
rect 3018 975 3019 979
rect 3023 975 3024 979
rect 3018 974 3024 975
rect 3050 979 3056 980
rect 3050 975 3051 979
rect 3055 978 3056 979
rect 3458 979 3464 980
rect 3055 976 3129 978
rect 3055 975 3056 976
rect 3050 974 3056 975
rect 3242 971 3248 972
rect 3242 970 3243 971
rect 2820 968 3243 970
rect 3242 967 3243 968
rect 3247 967 3248 971
rect 3428 970 3430 977
rect 3458 975 3459 979
rect 3463 978 3464 979
rect 4274 979 4280 980
rect 4274 978 4275 979
rect 3463 976 3553 978
rect 4165 976 4275 978
rect 3463 975 3464 976
rect 3458 974 3464 975
rect 4274 975 4275 976
rect 4279 975 4280 979
rect 4578 979 4584 980
rect 4274 974 4280 975
rect 3530 971 3536 972
rect 3530 970 3531 971
rect 3428 968 3531 970
rect 3242 966 3248 967
rect 3530 967 3531 968
rect 3535 967 3536 971
rect 4460 970 4462 977
rect 4578 975 4579 979
rect 4583 978 4584 979
rect 5074 979 5080 980
rect 4583 976 4665 978
rect 4583 975 4584 976
rect 4578 974 4584 975
rect 4778 971 4784 972
rect 4778 970 4779 971
rect 4460 968 4779 970
rect 3530 966 3536 967
rect 4778 967 4779 968
rect 4783 967 4784 971
rect 5044 970 5046 977
rect 5074 975 5075 979
rect 5079 978 5080 979
rect 5638 979 5644 980
rect 5638 978 5639 979
rect 5079 976 5241 978
rect 5613 976 5639 978
rect 5079 975 5080 976
rect 5074 974 5080 975
rect 5638 975 5639 976
rect 5643 975 5644 979
rect 5638 974 5644 975
rect 5374 971 5380 972
rect 5374 970 5375 971
rect 5044 968 5375 970
rect 4778 966 4784 967
rect 5374 967 5375 968
rect 5379 967 5380 971
rect 5374 966 5380 967
rect 2342 951 2348 952
rect 2342 950 2343 951
rect 2200 948 2343 950
rect 538 947 544 948
rect 538 946 539 947
rect 401 944 539 946
rect 401 942 403 944
rect 538 943 539 944
rect 543 943 544 947
rect 2200 946 2202 948
rect 2342 947 2343 948
rect 2347 947 2348 951
rect 2342 946 2348 947
rect 2650 947 2656 948
rect 2650 946 2651 947
rect 2093 944 2202 946
rect 2565 944 2651 946
rect 538 942 544 943
rect 734 943 740 944
rect 293 940 403 942
rect 426 939 432 940
rect 426 935 427 939
rect 431 935 432 939
rect 734 939 735 943
rect 739 939 740 943
rect 1154 943 1160 944
rect 734 938 740 939
rect 938 939 944 940
rect 426 934 432 935
rect 938 935 939 939
rect 943 935 944 939
rect 1154 939 1155 943
rect 1159 942 1160 943
rect 1986 943 1992 944
rect 1986 942 1987 943
rect 1159 940 1225 942
rect 1885 940 1987 942
rect 1159 939 1160 940
rect 1154 938 1160 939
rect 1522 939 1528 940
rect 938 934 944 935
rect 1522 935 1523 939
rect 1527 935 1528 939
rect 1986 939 1987 940
rect 1991 939 1992 943
rect 1986 938 1992 939
rect 2314 943 2320 944
rect 2314 939 2315 943
rect 2319 939 2320 943
rect 2650 943 2651 944
rect 2655 943 2656 947
rect 2650 942 2656 943
rect 2714 943 2720 944
rect 2314 938 2320 939
rect 2714 939 2715 943
rect 2719 939 2720 943
rect 2714 938 2720 939
rect 3034 943 3040 944
rect 3034 939 3035 943
rect 3039 939 3040 943
rect 3034 938 3040 939
rect 3178 943 3184 944
rect 3178 939 3179 943
rect 3183 939 3184 943
rect 3178 938 3184 939
rect 3418 943 3424 944
rect 3418 939 3419 943
rect 3423 939 3424 943
rect 3418 938 3424 939
rect 3982 943 3988 944
rect 3982 939 3983 943
rect 3987 939 3988 943
rect 4482 943 4488 944
rect 4482 942 4483 943
rect 4477 940 4483 942
rect 3982 938 3988 939
rect 4162 939 4168 940
rect 1522 934 1528 935
rect 4162 935 4163 939
rect 4167 935 4168 939
rect 4482 939 4483 940
rect 4487 939 4488 943
rect 5175 943 5181 944
rect 5175 942 5176 943
rect 5125 940 5176 942
rect 4482 938 4488 939
rect 4602 939 4608 940
rect 4162 934 4168 935
rect 4602 935 4603 939
rect 4607 935 4608 939
rect 4602 934 4608 935
rect 4818 939 4824 940
rect 4818 935 4819 939
rect 4823 935 4824 939
rect 5175 939 5176 940
rect 5180 939 5181 943
rect 5354 943 5360 944
rect 5354 942 5355 943
rect 5341 940 5355 942
rect 5175 938 5181 939
rect 5354 939 5355 940
rect 5359 939 5360 943
rect 5598 943 5604 944
rect 5598 942 5599 943
rect 5565 940 5599 942
rect 5354 938 5360 939
rect 5598 939 5599 940
rect 5603 939 5604 943
rect 5598 938 5604 939
rect 4818 934 4824 935
rect 5534 915 5540 916
rect 5534 911 5535 915
rect 5539 914 5540 915
rect 5590 915 5596 916
rect 5590 914 5591 915
rect 5539 912 5591 914
rect 5539 911 5540 912
rect 5534 910 5540 911
rect 5590 911 5591 912
rect 5595 911 5596 915
rect 5590 910 5596 911
rect 3034 903 3040 904
rect 3034 899 3035 903
rect 3039 902 3040 903
rect 3206 903 3212 904
rect 3206 902 3207 903
rect 3039 900 3207 902
rect 3039 899 3040 900
rect 3034 898 3040 899
rect 3206 899 3207 900
rect 3211 899 3212 903
rect 3206 898 3212 899
rect 1974 896 1980 897
rect 3798 896 3804 897
rect 110 892 116 893
rect 1934 892 1940 893
rect 110 888 111 892
rect 115 888 116 892
rect 110 887 116 888
rect 194 891 200 892
rect 194 887 195 891
rect 199 887 200 891
rect 194 886 200 887
rect 418 891 424 892
rect 418 887 419 891
rect 423 887 424 891
rect 418 886 424 887
rect 666 891 672 892
rect 666 887 667 891
rect 671 887 672 891
rect 666 886 672 887
rect 930 891 936 892
rect 930 887 931 891
rect 935 887 936 891
rect 930 886 936 887
rect 1218 891 1224 892
rect 1218 887 1219 891
rect 1223 887 1224 891
rect 1218 886 1224 887
rect 1514 891 1520 892
rect 1514 887 1515 891
rect 1519 887 1520 891
rect 1514 886 1520 887
rect 1786 891 1792 892
rect 1786 887 1787 891
rect 1791 887 1792 891
rect 1934 888 1935 892
rect 1939 888 1940 892
rect 1974 892 1975 896
rect 1979 892 1980 896
rect 1974 891 1980 892
rect 1994 895 2000 896
rect 1994 891 1995 895
rect 1999 891 2000 895
rect 1994 890 2000 891
rect 2218 895 2224 896
rect 2218 891 2219 895
rect 2223 891 2224 895
rect 2218 890 2224 891
rect 2466 895 2472 896
rect 2466 891 2467 895
rect 2471 891 2472 895
rect 2466 890 2472 891
rect 2706 895 2712 896
rect 2706 891 2707 895
rect 2711 891 2712 895
rect 2706 890 2712 891
rect 2938 895 2944 896
rect 2938 891 2939 895
rect 2943 891 2944 895
rect 2938 890 2944 891
rect 3170 895 3176 896
rect 3170 891 3171 895
rect 3175 891 3176 895
rect 3170 890 3176 891
rect 3410 895 3416 896
rect 3410 891 3411 895
rect 3415 891 3416 895
rect 3798 892 3799 896
rect 3803 892 3804 896
rect 3798 891 3804 892
rect 3838 892 3844 893
rect 5662 892 5668 893
rect 3410 890 3416 891
rect 3838 888 3839 892
rect 3843 888 3844 892
rect 1934 887 1940 888
rect 1986 887 1992 888
rect 3838 887 3844 888
rect 3930 891 3936 892
rect 3930 887 3931 891
rect 3935 887 3936 891
rect 1786 886 1792 887
rect 1986 883 1987 887
rect 1991 886 1992 887
rect 3930 886 3936 887
rect 4154 891 4160 892
rect 4154 887 4155 891
rect 4159 887 4160 891
rect 4154 886 4160 887
rect 4378 891 4384 892
rect 4378 887 4379 891
rect 4383 887 4384 891
rect 4378 886 4384 887
rect 4594 891 4600 892
rect 4594 887 4595 891
rect 4599 887 4600 891
rect 4594 886 4600 887
rect 4810 891 4816 892
rect 4810 887 4811 891
rect 4815 887 4816 891
rect 4810 886 4816 887
rect 5026 891 5032 892
rect 5026 887 5027 891
rect 5031 887 5032 891
rect 5026 886 5032 887
rect 5242 891 5248 892
rect 5242 887 5243 891
rect 5247 887 5248 891
rect 5242 886 5248 887
rect 5466 891 5472 892
rect 5466 887 5467 891
rect 5471 887 5472 891
rect 5662 888 5663 892
rect 5667 888 5668 892
rect 5662 887 5668 888
rect 5466 886 5472 887
rect 1991 884 2122 886
rect 1991 883 1992 884
rect 1986 882 1992 883
rect 2022 880 2028 881
rect 2120 880 2122 884
rect 5175 883 5181 884
rect 2246 880 2252 881
rect 2494 880 2500 881
rect 2734 880 2740 881
rect 2966 880 2972 881
rect 3198 880 3204 881
rect 3438 880 3444 881
rect 1974 879 1980 880
rect 222 876 228 877
rect 446 876 452 877
rect 694 876 700 877
rect 958 876 964 877
rect 1055 876 1061 877
rect 110 875 116 876
rect 110 871 111 875
rect 115 871 116 875
rect 222 872 223 876
rect 227 872 228 876
rect 222 871 228 872
rect 318 875 325 876
rect 318 871 319 875
rect 324 871 325 875
rect 446 872 447 876
rect 451 872 452 876
rect 446 871 452 872
rect 538 875 549 876
rect 538 871 539 875
rect 543 871 544 875
rect 548 871 549 875
rect 694 872 695 876
rect 699 872 700 876
rect 694 871 700 872
rect 791 875 797 876
rect 791 871 792 875
rect 796 874 797 875
rect 938 875 944 876
rect 938 874 939 875
rect 796 872 939 874
rect 796 871 797 872
rect 110 870 116 871
rect 318 870 325 871
rect 538 870 549 871
rect 791 870 797 871
rect 938 871 939 872
rect 943 871 944 875
rect 958 872 959 876
rect 963 872 964 876
rect 958 871 964 872
rect 1054 875 1056 876
rect 1054 871 1055 875
rect 1060 872 1061 876
rect 1059 871 1061 872
rect 1246 876 1252 877
rect 1542 876 1548 877
rect 1814 876 1820 877
rect 1246 872 1247 876
rect 1251 872 1252 876
rect 1246 871 1252 872
rect 1343 875 1349 876
rect 1343 871 1344 875
rect 1348 874 1349 875
rect 1522 875 1528 876
rect 1522 874 1523 875
rect 1348 872 1523 874
rect 1348 871 1349 872
rect 938 870 944 871
rect 1054 870 1060 871
rect 1343 870 1349 871
rect 1522 871 1523 872
rect 1527 871 1528 875
rect 1542 872 1543 876
rect 1547 872 1548 876
rect 1542 871 1548 872
rect 1638 875 1645 876
rect 1638 871 1639 875
rect 1644 871 1645 875
rect 1814 872 1815 876
rect 1819 872 1820 876
rect 1814 871 1820 872
rect 1906 875 1917 876
rect 1906 871 1907 875
rect 1911 871 1912 875
rect 1916 871 1917 875
rect 1522 870 1528 871
rect 1638 870 1645 871
rect 1906 870 1917 871
rect 1934 875 1940 876
rect 1934 871 1935 875
rect 1939 871 1940 875
rect 1974 875 1975 879
rect 1979 875 1980 879
rect 2022 876 2023 880
rect 2027 876 2028 880
rect 2022 875 2028 876
rect 2119 879 2125 880
rect 2119 875 2120 879
rect 2124 875 2125 879
rect 2246 876 2247 880
rect 2251 876 2252 880
rect 2246 875 2252 876
rect 2342 879 2349 880
rect 2342 875 2343 879
rect 2348 875 2349 879
rect 2494 876 2495 880
rect 2499 876 2500 880
rect 2494 875 2500 876
rect 2591 879 2597 880
rect 2591 875 2592 879
rect 2596 878 2597 879
rect 2714 879 2720 880
rect 2714 878 2715 879
rect 2596 876 2715 878
rect 2596 875 2597 876
rect 1974 874 1980 875
rect 2119 874 2125 875
rect 2342 874 2349 875
rect 2591 874 2597 875
rect 2714 875 2715 876
rect 2719 875 2720 879
rect 2734 876 2735 880
rect 2739 876 2740 880
rect 2734 875 2740 876
rect 2830 879 2837 880
rect 2830 875 2831 879
rect 2836 875 2837 879
rect 2966 876 2967 880
rect 2971 876 2972 880
rect 2966 875 2972 876
rect 3063 879 3069 880
rect 3063 875 3064 879
rect 3068 878 3069 879
rect 3178 879 3184 880
rect 3178 878 3179 879
rect 3068 876 3179 878
rect 3068 875 3069 876
rect 2714 874 2720 875
rect 2830 874 2837 875
rect 3063 874 3069 875
rect 3178 875 3179 876
rect 3183 875 3184 879
rect 3198 876 3199 880
rect 3203 876 3204 880
rect 3198 875 3204 876
rect 3295 879 3301 880
rect 3295 875 3296 879
rect 3300 878 3301 879
rect 3418 879 3424 880
rect 3418 878 3419 879
rect 3300 876 3419 878
rect 3300 875 3301 876
rect 3178 874 3184 875
rect 3295 874 3301 875
rect 3418 875 3419 876
rect 3423 875 3424 879
rect 3438 876 3439 880
rect 3443 876 3444 880
rect 3438 875 3444 876
rect 3530 879 3541 880
rect 3530 875 3531 879
rect 3535 875 3536 879
rect 3540 875 3541 879
rect 3418 874 3424 875
rect 3530 874 3541 875
rect 3798 879 3804 880
rect 3798 875 3799 879
rect 3803 875 3804 879
rect 5175 879 5176 883
rect 5180 882 5181 883
rect 5180 880 5370 882
rect 5180 879 5181 880
rect 5175 878 5181 879
rect 5368 878 5370 880
rect 5367 877 5373 878
rect 3958 876 3964 877
rect 4182 876 4188 877
rect 4406 876 4412 877
rect 4622 876 4628 877
rect 4838 876 4844 877
rect 5054 876 5060 877
rect 5270 876 5276 877
rect 3798 874 3804 875
rect 3838 875 3844 876
rect 1934 870 1940 871
rect 3838 871 3839 875
rect 3843 871 3844 875
rect 3958 872 3959 876
rect 3963 872 3964 876
rect 3958 871 3964 872
rect 4055 875 4061 876
rect 4055 871 4056 875
rect 4060 874 4061 875
rect 4162 875 4168 876
rect 4162 874 4163 875
rect 4060 872 4163 874
rect 4060 871 4061 872
rect 3838 870 3844 871
rect 4055 870 4061 871
rect 4162 871 4163 872
rect 4167 871 4168 875
rect 4182 872 4183 876
rect 4187 872 4188 876
rect 4182 871 4188 872
rect 4274 875 4285 876
rect 4274 871 4275 875
rect 4279 871 4280 875
rect 4284 871 4285 875
rect 4406 872 4407 876
rect 4411 872 4412 876
rect 4406 871 4412 872
rect 4503 875 4509 876
rect 4503 871 4504 875
rect 4508 874 4509 875
rect 4602 875 4608 876
rect 4602 874 4603 875
rect 4508 872 4603 874
rect 4508 871 4509 872
rect 4162 870 4168 871
rect 4274 870 4285 871
rect 4503 870 4509 871
rect 4602 871 4603 872
rect 4607 871 4608 875
rect 4622 872 4623 876
rect 4627 872 4628 876
rect 4622 871 4628 872
rect 4719 875 4725 876
rect 4719 871 4720 875
rect 4724 874 4725 875
rect 4818 875 4824 876
rect 4818 874 4819 875
rect 4724 872 4819 874
rect 4724 871 4725 872
rect 4602 870 4608 871
rect 4719 870 4725 871
rect 4818 871 4819 872
rect 4823 871 4824 875
rect 4838 872 4839 876
rect 4843 872 4844 876
rect 4838 871 4844 872
rect 4930 875 4941 876
rect 4930 871 4931 875
rect 4935 871 4936 875
rect 4940 871 4941 875
rect 5054 872 5055 876
rect 5059 872 5060 876
rect 5054 871 5060 872
rect 5151 875 5160 876
rect 5151 871 5152 875
rect 5159 871 5160 875
rect 5270 872 5271 876
rect 5275 872 5276 876
rect 5367 873 5368 877
rect 5372 873 5373 877
rect 5367 872 5373 873
rect 5494 876 5500 877
rect 5494 872 5495 876
rect 5499 872 5500 876
rect 5270 871 5276 872
rect 5494 871 5500 872
rect 5590 875 5597 876
rect 5590 871 5591 875
rect 5596 871 5597 875
rect 4818 870 4824 871
rect 4930 870 4941 871
rect 5151 870 5160 871
rect 5590 870 5597 871
rect 5662 875 5668 876
rect 5662 871 5663 875
rect 5667 871 5668 875
rect 5662 870 5668 871
rect 538 859 544 860
rect 538 855 539 859
rect 543 858 544 859
rect 1054 859 1060 860
rect 1054 858 1055 859
rect 543 856 1055 858
rect 543 855 544 856
rect 538 854 544 855
rect 1054 855 1055 856
rect 1059 855 1060 859
rect 1054 854 1060 855
rect 1974 821 1980 822
rect 3798 821 3804 822
rect 1974 817 1975 821
rect 1979 817 1980 821
rect 1974 816 1980 817
rect 2222 820 2228 821
rect 2438 820 2444 821
rect 2662 820 2668 821
rect 2886 820 2892 821
rect 3110 820 3116 821
rect 3334 820 3340 821
rect 3558 820 3564 821
rect 2222 816 2223 820
rect 2227 816 2228 820
rect 2222 815 2228 816
rect 2314 819 2325 820
rect 2314 815 2315 819
rect 2319 815 2320 819
rect 2324 815 2325 819
rect 2438 816 2439 820
rect 2443 816 2444 820
rect 2438 815 2444 816
rect 2534 819 2541 820
rect 2534 815 2535 819
rect 2540 815 2541 819
rect 2662 816 2663 820
rect 2667 816 2668 820
rect 2662 815 2668 816
rect 2758 819 2765 820
rect 2758 815 2759 819
rect 2764 815 2765 819
rect 2886 816 2887 820
rect 2891 816 2892 820
rect 2886 815 2892 816
rect 2978 819 2989 820
rect 2978 815 2979 819
rect 2983 815 2984 819
rect 2988 815 2989 819
rect 3110 816 3111 820
rect 3115 816 3116 820
rect 3110 815 3116 816
rect 3206 819 3213 820
rect 3206 815 3207 819
rect 3212 815 3213 819
rect 3334 816 3335 820
rect 3339 816 3340 820
rect 3334 815 3340 816
rect 3430 819 3437 820
rect 3430 815 3431 819
rect 3436 815 3437 819
rect 3558 816 3559 820
rect 3563 816 3564 820
rect 3558 815 3564 816
rect 3650 819 3661 820
rect 3650 815 3651 819
rect 3655 815 3656 819
rect 3660 815 3661 819
rect 3798 817 3799 821
rect 3803 817 3804 821
rect 3798 816 3804 817
rect 3838 817 3844 818
rect 5662 817 5668 818
rect 2314 814 2325 815
rect 2534 814 2541 815
rect 2758 814 2765 815
rect 2978 814 2989 815
rect 3206 814 3213 815
rect 3430 814 3437 815
rect 3650 814 3661 815
rect 3838 813 3839 817
rect 3843 813 3844 817
rect 3838 812 3844 813
rect 3886 816 3892 817
rect 4110 816 4116 817
rect 4342 816 4348 817
rect 4574 816 4580 817
rect 4798 816 4804 817
rect 5030 816 5036 817
rect 5262 816 5268 817
rect 5494 816 5500 817
rect 3886 812 3887 816
rect 3891 812 3892 816
rect 3886 811 3892 812
rect 3982 815 3989 816
rect 3982 811 3983 815
rect 3988 811 3989 815
rect 4110 812 4111 816
rect 4115 812 4116 816
rect 4110 811 4116 812
rect 4206 815 4213 816
rect 4206 811 4207 815
rect 4212 811 4213 815
rect 4342 812 4343 816
rect 4347 812 4348 816
rect 4342 811 4348 812
rect 4439 815 4445 816
rect 4439 811 4440 815
rect 4444 814 4445 815
rect 4495 815 4501 816
rect 4495 814 4496 815
rect 4444 812 4496 814
rect 4444 811 4445 812
rect 3982 810 3989 811
rect 4206 810 4213 811
rect 4439 810 4445 811
rect 4495 811 4496 812
rect 4500 811 4501 815
rect 4574 812 4575 816
rect 4579 812 4580 816
rect 4574 811 4580 812
rect 4671 815 4680 816
rect 4671 811 4672 815
rect 4679 811 4680 815
rect 4798 812 4799 816
rect 4803 812 4804 816
rect 4798 811 4804 812
rect 4890 815 4901 816
rect 4890 811 4891 815
rect 4895 811 4896 815
rect 4900 811 4901 815
rect 5030 812 5031 816
rect 5035 812 5036 816
rect 5030 811 5036 812
rect 5122 815 5133 816
rect 5122 811 5123 815
rect 5127 811 5128 815
rect 5132 811 5133 815
rect 5262 812 5263 816
rect 5267 812 5268 816
rect 5262 811 5268 812
rect 5354 815 5365 816
rect 5354 811 5355 815
rect 5359 811 5360 815
rect 5364 811 5365 815
rect 5494 812 5495 816
rect 5499 812 5500 816
rect 5494 811 5500 812
rect 5591 815 5597 816
rect 5591 811 5592 815
rect 5596 811 5597 815
rect 5662 813 5663 817
rect 5667 813 5668 817
rect 5662 812 5668 813
rect 4495 810 4501 811
rect 4671 810 4680 811
rect 4890 810 4901 811
rect 5122 810 5133 811
rect 5354 810 5365 811
rect 5591 810 5597 811
rect 2194 805 2200 806
rect 1974 804 1980 805
rect 1974 800 1975 804
rect 1979 800 1980 804
rect 2194 801 2195 805
rect 2199 801 2200 805
rect 2194 800 2200 801
rect 2410 805 2416 806
rect 2410 801 2411 805
rect 2415 801 2416 805
rect 2410 800 2416 801
rect 2634 805 2640 806
rect 2634 801 2635 805
rect 2639 801 2640 805
rect 2634 800 2640 801
rect 2858 805 2864 806
rect 2858 801 2859 805
rect 2863 801 2864 805
rect 2858 800 2864 801
rect 3082 805 3088 806
rect 3082 801 3083 805
rect 3087 801 3088 805
rect 3082 800 3088 801
rect 3306 805 3312 806
rect 3306 801 3307 805
rect 3311 801 3312 805
rect 3306 800 3312 801
rect 3530 805 3536 806
rect 3530 801 3531 805
rect 3535 801 3536 805
rect 3530 800 3536 801
rect 3798 804 3804 805
rect 3798 800 3799 804
rect 3803 800 3804 804
rect 3858 801 3864 802
rect 1974 799 1980 800
rect 3798 799 3804 800
rect 3838 800 3844 801
rect 3838 796 3839 800
rect 3843 796 3844 800
rect 3858 797 3859 801
rect 3863 797 3864 801
rect 3858 796 3864 797
rect 4082 801 4088 802
rect 4082 797 4083 801
rect 4087 797 4088 801
rect 4082 796 4088 797
rect 4314 801 4320 802
rect 4314 797 4315 801
rect 4319 797 4320 801
rect 4314 796 4320 797
rect 4546 801 4552 802
rect 4546 797 4547 801
rect 4551 797 4552 801
rect 4546 796 4552 797
rect 4770 801 4776 802
rect 4770 797 4771 801
rect 4775 797 4776 801
rect 4770 796 4776 797
rect 5002 801 5008 802
rect 5002 797 5003 801
rect 5007 797 5008 801
rect 5002 796 5008 797
rect 5234 801 5240 802
rect 5234 797 5235 801
rect 5239 797 5240 801
rect 5234 796 5240 797
rect 5466 801 5472 802
rect 5466 797 5467 801
rect 5471 797 5472 801
rect 5466 796 5472 797
rect 5662 800 5668 801
rect 5662 796 5663 800
rect 5667 796 5668 800
rect 3838 795 3844 796
rect 5662 795 5668 796
rect 110 793 116 794
rect 1934 793 1940 794
rect 110 789 111 793
rect 115 789 116 793
rect 110 788 116 789
rect 222 792 228 793
rect 446 792 452 793
rect 662 792 668 793
rect 878 792 884 793
rect 1086 792 1092 793
rect 1294 792 1300 793
rect 1510 792 1516 793
rect 222 788 223 792
rect 227 788 228 792
rect 222 787 228 788
rect 319 791 325 792
rect 319 787 320 791
rect 324 790 325 791
rect 426 791 432 792
rect 426 790 427 791
rect 324 788 427 790
rect 324 787 325 788
rect 319 786 325 787
rect 426 787 427 788
rect 431 787 432 791
rect 446 788 447 792
rect 451 788 452 792
rect 446 787 452 788
rect 543 791 552 792
rect 543 787 544 791
rect 551 787 552 791
rect 662 788 663 792
rect 667 788 668 792
rect 662 787 668 788
rect 759 791 768 792
rect 759 787 760 791
rect 767 787 768 791
rect 878 788 879 792
rect 883 788 884 792
rect 878 787 884 788
rect 974 791 981 792
rect 974 787 975 791
rect 980 787 981 791
rect 1086 788 1087 792
rect 1091 788 1092 792
rect 1086 787 1092 788
rect 1178 791 1189 792
rect 1178 787 1179 791
rect 1183 787 1184 791
rect 1188 787 1189 791
rect 1294 788 1295 792
rect 1299 788 1300 792
rect 1294 787 1300 788
rect 1386 791 1397 792
rect 1386 787 1387 791
rect 1391 787 1392 791
rect 1396 787 1397 791
rect 1510 788 1511 792
rect 1515 788 1516 792
rect 1510 787 1516 788
rect 1606 791 1613 792
rect 1606 787 1607 791
rect 1612 787 1613 791
rect 1934 789 1935 793
rect 1939 789 1940 793
rect 1934 788 1940 789
rect 426 786 432 787
rect 543 786 552 787
rect 759 786 768 787
rect 974 786 981 787
rect 1178 786 1189 787
rect 1386 786 1397 787
rect 1606 786 1613 787
rect 3178 783 3184 784
rect 3178 779 3179 783
rect 3183 782 3184 783
rect 3430 783 3436 784
rect 3430 782 3431 783
rect 3183 780 3431 782
rect 3183 779 3184 780
rect 3178 778 3184 779
rect 3430 779 3431 780
rect 3435 779 3436 783
rect 3430 778 3436 779
rect 3954 783 3960 784
rect 3954 779 3955 783
rect 3959 782 3960 783
rect 4206 783 4212 784
rect 4206 782 4207 783
rect 3959 780 4207 782
rect 3959 779 3960 780
rect 3954 778 3960 779
rect 4206 779 4207 780
rect 4211 779 4212 783
rect 4206 778 4212 779
rect 194 777 200 778
rect 110 776 116 777
rect 110 772 111 776
rect 115 772 116 776
rect 194 773 195 777
rect 199 773 200 777
rect 194 772 200 773
rect 418 777 424 778
rect 418 773 419 777
rect 423 773 424 777
rect 418 772 424 773
rect 634 777 640 778
rect 634 773 635 777
rect 639 773 640 777
rect 634 772 640 773
rect 850 777 856 778
rect 850 773 851 777
rect 855 773 856 777
rect 850 772 856 773
rect 1058 777 1064 778
rect 1058 773 1059 777
rect 1063 773 1064 777
rect 1058 772 1064 773
rect 1266 777 1272 778
rect 1266 773 1267 777
rect 1271 773 1272 777
rect 1266 772 1272 773
rect 1482 777 1488 778
rect 1482 773 1483 777
rect 1487 773 1488 777
rect 1482 772 1488 773
rect 1934 776 1940 777
rect 1934 772 1935 776
rect 1939 772 1940 776
rect 110 771 116 772
rect 1934 771 1940 772
rect 2830 755 2836 756
rect 2292 746 2294 753
rect 2509 752 2638 754
rect 2733 752 2781 754
rect 2534 747 2540 748
rect 2534 746 2535 747
rect 2292 744 2535 746
rect 2534 743 2535 744
rect 2539 743 2540 747
rect 2636 746 2638 752
rect 2758 747 2764 748
rect 2758 746 2759 747
rect 2636 744 2759 746
rect 2534 742 2540 743
rect 2758 743 2759 744
rect 2763 743 2764 747
rect 2779 746 2781 752
rect 2830 751 2831 755
rect 2835 754 2836 755
rect 3178 755 3184 756
rect 2835 752 2865 754
rect 2835 751 2836 752
rect 2830 750 2836 751
rect 3178 751 3179 755
rect 3183 751 3184 755
rect 3506 755 3512 756
rect 3178 750 3184 751
rect 2978 747 2984 748
rect 2978 746 2979 747
rect 2779 744 2979 746
rect 2758 742 2764 743
rect 2978 743 2979 744
rect 2983 743 2984 747
rect 3404 746 3406 753
rect 3506 751 3507 755
rect 3511 754 3512 755
rect 3511 752 3537 754
rect 3511 751 3512 752
rect 3506 750 3512 751
rect 3954 751 3960 752
rect 3650 747 3656 748
rect 3650 746 3651 747
rect 3404 744 3651 746
rect 2978 742 2984 743
rect 3650 743 3651 744
rect 3655 743 3656 747
rect 3954 747 3955 751
rect 3959 747 3960 751
rect 4202 751 4208 752
rect 4202 750 4203 751
rect 4181 748 4203 750
rect 3954 746 3960 747
rect 4202 747 4203 748
rect 4207 747 4208 751
rect 4495 751 4501 752
rect 4413 748 4461 750
rect 4202 746 4208 747
rect 3650 742 3656 743
rect 4459 742 4461 748
rect 4495 747 4496 751
rect 4500 750 4501 751
rect 4674 751 4680 752
rect 4500 748 4553 750
rect 4500 747 4501 748
rect 4495 746 4501 747
rect 4674 747 4675 751
rect 4679 750 4680 751
rect 5154 751 5160 752
rect 4679 748 4777 750
rect 4679 747 4680 748
rect 4674 746 4680 747
rect 4930 743 4936 744
rect 4930 742 4931 743
rect 4459 740 4931 742
rect 4930 739 4931 740
rect 4935 739 4936 743
rect 5100 742 5102 749
rect 5154 747 5155 751
rect 5159 750 5160 751
rect 5646 751 5652 752
rect 5646 750 5647 751
rect 5159 748 5241 750
rect 5565 748 5647 750
rect 5159 747 5160 748
rect 5154 746 5160 747
rect 5646 747 5647 748
rect 5651 747 5652 751
rect 5646 746 5652 747
rect 5354 743 5360 744
rect 5354 742 5355 743
rect 5100 740 5355 742
rect 4930 738 4936 739
rect 5354 739 5355 740
rect 5359 739 5360 743
rect 5354 738 5360 739
rect 4650 735 4656 736
rect 4650 731 4651 735
rect 4655 734 4656 735
rect 5122 735 5128 736
rect 5122 734 5123 735
rect 4655 732 5123 734
rect 4655 731 4656 732
rect 4650 730 4656 731
rect 5122 731 5123 732
rect 5127 731 5128 735
rect 5122 730 5128 731
rect 538 727 544 728
rect 538 726 539 727
rect 292 718 294 725
rect 517 724 539 726
rect 538 723 539 724
rect 543 723 544 727
rect 538 722 544 723
rect 546 727 552 728
rect 546 723 547 727
rect 551 726 552 727
rect 762 727 768 728
rect 551 724 641 726
rect 551 723 552 724
rect 546 722 552 723
rect 762 723 763 727
rect 767 726 768 727
rect 1638 727 1644 728
rect 1638 726 1639 727
rect 767 724 857 726
rect 767 723 768 724
rect 762 722 768 723
rect 562 719 568 720
rect 562 718 563 719
rect 292 716 563 718
rect 562 715 563 716
rect 567 715 568 719
rect 1156 718 1158 725
rect 1365 724 1470 726
rect 1581 724 1639 726
rect 1386 719 1392 720
rect 1386 718 1387 719
rect 1156 716 1387 718
rect 562 714 568 715
rect 1386 715 1387 716
rect 1391 715 1392 719
rect 1468 718 1470 724
rect 1638 723 1639 724
rect 1643 723 1644 727
rect 1638 722 1644 723
rect 4678 723 4684 724
rect 4678 722 4679 723
rect 4459 720 4679 722
rect 1606 719 1612 720
rect 1606 718 1607 719
rect 1468 716 1607 718
rect 1386 714 1392 715
rect 1606 715 1607 716
rect 1611 715 1612 719
rect 3982 719 3988 720
rect 3982 718 3983 719
rect 3957 716 3983 718
rect 1606 714 1612 715
rect 3982 715 3983 716
rect 3987 715 3988 719
rect 4459 718 4461 720
rect 4678 719 4679 720
rect 4683 719 4684 723
rect 4678 718 4684 719
rect 4890 719 4896 720
rect 4890 718 4891 719
rect 4421 716 4461 718
rect 4877 716 4891 718
rect 3982 714 3988 715
rect 4090 715 4096 716
rect 4090 711 4091 715
rect 4095 711 4096 715
rect 4090 710 4096 711
rect 4650 715 4656 716
rect 4650 711 4651 715
rect 4655 711 4656 715
rect 4890 715 4891 716
rect 4895 715 4896 719
rect 5638 719 5644 720
rect 5638 718 5639 719
rect 5557 716 5639 718
rect 4890 714 4896 715
rect 5010 715 5016 716
rect 4650 710 4656 711
rect 5010 711 5011 715
rect 5015 711 5016 715
rect 5010 710 5016 711
rect 5234 715 5240 716
rect 5234 711 5235 715
rect 5239 711 5240 715
rect 5638 715 5639 716
rect 5643 715 5644 719
rect 5638 714 5644 715
rect 5234 710 5240 711
rect 3647 707 3653 708
rect 3647 706 3648 707
rect 3613 704 3648 706
rect 3474 703 3480 704
rect 3474 699 3475 703
rect 3479 699 3480 703
rect 3647 703 3648 704
rect 3652 703 3653 707
rect 3774 707 3780 708
rect 3774 706 3775 707
rect 3749 704 3775 706
rect 3647 702 3653 703
rect 3774 703 3775 704
rect 3779 703 3780 707
rect 3774 702 3780 703
rect 3474 698 3480 699
rect 254 687 260 688
rect 254 686 255 687
rect 229 684 255 686
rect 254 683 255 684
rect 259 683 260 687
rect 762 687 768 688
rect 762 686 763 687
rect 709 684 763 686
rect 254 682 260 683
rect 282 683 288 684
rect 282 679 283 683
rect 287 679 288 683
rect 282 678 288 679
rect 450 683 456 684
rect 450 679 451 683
rect 455 679 456 683
rect 762 683 763 684
rect 767 683 768 687
rect 910 687 916 688
rect 910 686 911 687
rect 869 684 911 686
rect 762 682 768 683
rect 910 683 911 684
rect 915 683 916 687
rect 910 682 916 683
rect 974 687 980 688
rect 974 683 975 687
rect 979 683 980 687
rect 1178 687 1184 688
rect 1178 686 1179 687
rect 1173 684 1179 686
rect 974 682 980 683
rect 1178 683 1179 684
rect 1183 683 1184 687
rect 1178 682 1184 683
rect 1226 683 1232 684
rect 450 678 456 679
rect 1226 679 1227 683
rect 1231 679 1232 683
rect 1226 678 1232 679
rect 1370 683 1376 684
rect 1370 679 1371 683
rect 1375 679 1376 683
rect 1370 678 1376 679
rect 1514 683 1520 684
rect 1514 679 1515 683
rect 1519 679 1520 683
rect 1514 678 1520 679
rect 1658 683 1664 684
rect 1658 679 1659 683
rect 1663 679 1664 683
rect 1658 678 1664 679
rect 1794 683 1800 684
rect 1794 679 1795 683
rect 1799 679 1800 683
rect 1794 678 1800 679
rect 3838 668 3844 669
rect 5662 668 5668 669
rect 3838 664 3839 668
rect 3843 664 3844 668
rect 3474 663 3480 664
rect 3474 659 3475 663
rect 3479 662 3480 663
rect 3638 663 3644 664
rect 3838 663 3844 664
rect 3858 667 3864 668
rect 3858 663 3859 667
rect 3863 663 3864 667
rect 3638 662 3639 663
rect 3479 660 3639 662
rect 3479 659 3480 660
rect 3474 658 3480 659
rect 3638 659 3639 660
rect 3643 659 3644 663
rect 3858 662 3864 663
rect 4082 667 4088 668
rect 4082 663 4083 667
rect 4087 663 4088 667
rect 4082 662 4088 663
rect 4322 667 4328 668
rect 4322 663 4323 667
rect 4327 663 4328 667
rect 4322 662 4328 663
rect 4554 667 4560 668
rect 4554 663 4555 667
rect 4559 663 4560 667
rect 4554 662 4560 663
rect 4778 667 4784 668
rect 4778 663 4779 667
rect 4783 663 4784 667
rect 4778 662 4784 663
rect 5002 667 5008 668
rect 5002 663 5003 667
rect 5007 663 5008 667
rect 5002 662 5008 663
rect 5226 667 5232 668
rect 5226 663 5227 667
rect 5231 663 5232 667
rect 5226 662 5232 663
rect 5458 667 5464 668
rect 5458 663 5459 667
rect 5463 663 5464 667
rect 5662 664 5663 668
rect 5667 664 5668 668
rect 5662 663 5668 664
rect 5458 662 5464 663
rect 3638 658 3644 659
rect 1974 656 1980 657
rect 3798 656 3804 657
rect 1974 652 1975 656
rect 1979 652 1980 656
rect 1974 651 1980 652
rect 3378 655 3384 656
rect 3378 651 3379 655
rect 3383 651 3384 655
rect 3378 650 3384 651
rect 3514 655 3520 656
rect 3514 651 3515 655
rect 3519 651 3520 655
rect 3514 650 3520 651
rect 3650 655 3656 656
rect 3650 651 3651 655
rect 3655 651 3656 655
rect 3798 652 3799 656
rect 3803 652 3804 656
rect 3886 652 3892 653
rect 4110 652 4116 653
rect 4350 652 4356 653
rect 4582 652 4588 653
rect 4806 652 4812 653
rect 5030 652 5036 653
rect 5254 652 5260 653
rect 5486 652 5492 653
rect 3798 651 3804 652
rect 3838 651 3844 652
rect 3650 650 3656 651
rect 3838 647 3839 651
rect 3843 647 3844 651
rect 3886 648 3887 652
rect 3891 648 3892 652
rect 3886 647 3892 648
rect 3983 651 3989 652
rect 3983 647 3984 651
rect 3988 650 3989 651
rect 4090 651 4096 652
rect 4090 650 4091 651
rect 3988 648 4091 650
rect 3988 647 3989 648
rect 3838 646 3844 647
rect 3983 646 3989 647
rect 4090 647 4091 648
rect 4095 647 4096 651
rect 4110 648 4111 652
rect 4115 648 4116 652
rect 4110 647 4116 648
rect 4202 651 4213 652
rect 4202 647 4203 651
rect 4207 647 4208 651
rect 4212 647 4213 651
rect 4350 648 4351 652
rect 4355 648 4356 652
rect 4350 647 4356 648
rect 4446 651 4453 652
rect 4446 647 4447 651
rect 4452 647 4453 651
rect 4582 648 4583 652
rect 4587 648 4588 652
rect 4582 647 4588 648
rect 4678 651 4685 652
rect 4678 647 4679 651
rect 4684 647 4685 651
rect 4806 648 4807 652
rect 4811 648 4812 652
rect 4806 647 4812 648
rect 4903 651 4909 652
rect 4903 647 4904 651
rect 4908 650 4909 651
rect 5010 651 5016 652
rect 5010 650 5011 651
rect 4908 648 5011 650
rect 4908 647 4909 648
rect 4090 646 4096 647
rect 4202 646 4213 647
rect 4446 646 4453 647
rect 4678 646 4685 647
rect 4903 646 4909 647
rect 5010 647 5011 648
rect 5015 647 5016 651
rect 5030 648 5031 652
rect 5035 648 5036 652
rect 5030 647 5036 648
rect 5127 651 5133 652
rect 5127 647 5128 651
rect 5132 650 5133 651
rect 5234 651 5240 652
rect 5234 650 5235 651
rect 5132 648 5235 650
rect 5132 647 5133 648
rect 5010 646 5016 647
rect 5127 646 5133 647
rect 5234 647 5235 648
rect 5239 647 5240 651
rect 5254 648 5255 652
rect 5259 648 5260 652
rect 5254 647 5260 648
rect 5346 651 5357 652
rect 5346 647 5347 651
rect 5351 647 5352 651
rect 5356 647 5357 651
rect 5486 648 5487 652
rect 5491 648 5492 652
rect 5486 647 5492 648
rect 5582 651 5589 652
rect 5582 647 5583 651
rect 5588 647 5589 651
rect 5234 646 5240 647
rect 5346 646 5357 647
rect 5582 646 5589 647
rect 5662 651 5668 652
rect 5662 647 5663 651
rect 5667 647 5668 651
rect 5662 646 5668 647
rect 3672 644 3779 646
rect 3647 643 3653 644
rect 3406 640 3412 641
rect 3542 640 3548 641
rect 1974 639 1980 640
rect 110 636 116 637
rect 1934 636 1940 637
rect 110 632 111 636
rect 115 632 116 636
rect 110 631 116 632
rect 130 635 136 636
rect 130 631 131 635
rect 135 631 136 635
rect 130 630 136 631
rect 274 635 280 636
rect 274 631 275 635
rect 279 631 280 635
rect 274 630 280 631
rect 442 635 448 636
rect 442 631 443 635
rect 447 631 448 635
rect 442 630 448 631
rect 610 635 616 636
rect 610 631 611 635
rect 615 631 616 635
rect 610 630 616 631
rect 770 635 776 636
rect 770 631 771 635
rect 775 631 776 635
rect 770 630 776 631
rect 922 635 928 636
rect 922 631 923 635
rect 927 631 928 635
rect 922 630 928 631
rect 1074 635 1080 636
rect 1074 631 1075 635
rect 1079 631 1080 635
rect 1074 630 1080 631
rect 1218 635 1224 636
rect 1218 631 1219 635
rect 1223 631 1224 635
rect 1218 630 1224 631
rect 1362 635 1368 636
rect 1362 631 1363 635
rect 1367 631 1368 635
rect 1362 630 1368 631
rect 1506 635 1512 636
rect 1506 631 1507 635
rect 1511 631 1512 635
rect 1506 630 1512 631
rect 1650 635 1656 636
rect 1650 631 1651 635
rect 1655 631 1656 635
rect 1650 630 1656 631
rect 1786 635 1792 636
rect 1786 631 1787 635
rect 1791 631 1792 635
rect 1934 632 1935 636
rect 1939 632 1940 636
rect 1974 635 1975 639
rect 1979 635 1980 639
rect 3406 636 3407 640
rect 3411 636 3412 640
rect 3406 635 3412 636
rect 3503 639 3512 640
rect 3503 635 3504 639
rect 3511 635 3512 639
rect 3542 636 3543 640
rect 3547 636 3548 640
rect 3542 635 3548 636
rect 3638 639 3645 640
rect 3638 635 3639 639
rect 3644 635 3645 639
rect 3647 639 3648 643
rect 3652 642 3653 643
rect 3672 642 3674 644
rect 3652 640 3674 642
rect 3678 640 3684 641
rect 3777 640 3779 644
rect 3652 639 3653 640
rect 3647 638 3653 639
rect 3678 636 3679 640
rect 3683 636 3684 640
rect 3678 635 3684 636
rect 3775 639 3781 640
rect 3775 635 3776 639
rect 3780 635 3781 639
rect 1974 634 1980 635
rect 3503 634 3512 635
rect 3638 634 3645 635
rect 3775 634 3781 635
rect 3798 639 3804 640
rect 3798 635 3799 639
rect 3803 635 3804 639
rect 3798 634 3804 635
rect 1934 631 1940 632
rect 1786 630 1792 631
rect 762 627 768 628
rect 762 623 763 627
rect 767 626 768 627
rect 910 627 916 628
rect 767 624 891 626
rect 767 623 768 624
rect 762 622 768 623
rect 158 620 164 621
rect 302 620 308 621
rect 470 620 476 621
rect 638 620 644 621
rect 798 620 804 621
rect 110 619 116 620
rect 110 615 111 619
rect 115 615 116 619
rect 158 616 159 620
rect 163 616 164 620
rect 158 615 164 616
rect 255 619 261 620
rect 255 615 256 619
rect 260 618 261 619
rect 282 619 288 620
rect 282 618 283 619
rect 260 616 283 618
rect 260 615 261 616
rect 110 614 116 615
rect 255 614 261 615
rect 282 615 283 616
rect 287 615 288 619
rect 302 616 303 620
rect 307 616 308 620
rect 302 615 308 616
rect 399 619 405 620
rect 399 615 400 619
rect 404 618 405 619
rect 450 619 456 620
rect 450 618 451 619
rect 404 616 451 618
rect 404 615 405 616
rect 282 614 288 615
rect 399 614 405 615
rect 450 615 451 616
rect 455 615 456 619
rect 470 616 471 620
rect 475 616 476 620
rect 470 615 476 616
rect 562 619 573 620
rect 562 615 563 619
rect 567 615 568 619
rect 572 615 573 619
rect 638 616 639 620
rect 643 616 644 620
rect 638 615 644 616
rect 734 619 741 620
rect 734 615 735 619
rect 740 615 741 619
rect 798 616 799 620
rect 803 616 804 620
rect 889 618 891 624
rect 910 623 911 627
rect 915 626 916 627
rect 915 624 1051 626
rect 915 623 916 624
rect 910 622 916 623
rect 950 620 956 621
rect 1049 620 1051 624
rect 1102 620 1108 621
rect 1246 620 1252 621
rect 1390 620 1396 621
rect 1534 620 1540 621
rect 1678 620 1684 621
rect 1814 620 1820 621
rect 895 619 901 620
rect 895 618 896 619
rect 889 616 896 618
rect 798 615 804 616
rect 895 615 896 616
rect 900 615 901 619
rect 950 616 951 620
rect 955 616 956 620
rect 950 615 956 616
rect 1047 619 1053 620
rect 1047 615 1048 619
rect 1052 615 1053 619
rect 1102 616 1103 620
rect 1107 616 1108 620
rect 1102 615 1108 616
rect 1199 619 1205 620
rect 1199 615 1200 619
rect 1204 618 1205 619
rect 1226 619 1232 620
rect 1226 618 1227 619
rect 1204 616 1227 618
rect 1204 615 1205 616
rect 450 614 456 615
rect 562 614 573 615
rect 734 614 741 615
rect 895 614 901 615
rect 1047 614 1053 615
rect 1199 614 1205 615
rect 1226 615 1227 616
rect 1231 615 1232 619
rect 1246 616 1247 620
rect 1251 616 1252 620
rect 1246 615 1252 616
rect 1343 619 1349 620
rect 1343 615 1344 619
rect 1348 618 1349 619
rect 1370 619 1376 620
rect 1370 618 1371 619
rect 1348 616 1371 618
rect 1348 615 1349 616
rect 1226 614 1232 615
rect 1343 614 1349 615
rect 1370 615 1371 616
rect 1375 615 1376 619
rect 1390 616 1391 620
rect 1395 616 1396 620
rect 1390 615 1396 616
rect 1487 619 1493 620
rect 1487 615 1488 619
rect 1492 618 1493 619
rect 1514 619 1520 620
rect 1514 618 1515 619
rect 1492 616 1515 618
rect 1492 615 1493 616
rect 1370 614 1376 615
rect 1487 614 1493 615
rect 1514 615 1515 616
rect 1519 615 1520 619
rect 1534 616 1535 620
rect 1539 616 1540 620
rect 1534 615 1540 616
rect 1631 619 1637 620
rect 1631 615 1632 619
rect 1636 618 1637 619
rect 1658 619 1664 620
rect 1658 618 1659 619
rect 1636 616 1659 618
rect 1636 615 1637 616
rect 1514 614 1520 615
rect 1631 614 1637 615
rect 1658 615 1659 616
rect 1663 615 1664 619
rect 1678 616 1679 620
rect 1683 616 1684 620
rect 1678 615 1684 616
rect 1775 619 1781 620
rect 1775 615 1776 619
rect 1780 618 1781 619
rect 1794 619 1800 620
rect 1794 618 1795 619
rect 1780 616 1795 618
rect 1780 615 1781 616
rect 1658 614 1664 615
rect 1775 614 1781 615
rect 1794 615 1795 616
rect 1799 615 1800 619
rect 1814 616 1815 620
rect 1819 616 1820 620
rect 1814 615 1820 616
rect 1910 619 1917 620
rect 1910 615 1911 619
rect 1916 615 1917 619
rect 1794 614 1800 615
rect 1910 614 1917 615
rect 1934 619 1940 620
rect 1934 615 1935 619
rect 1939 615 1940 619
rect 1934 614 1940 615
rect 3838 585 3844 586
rect 5662 585 5668 586
rect 3838 581 3839 585
rect 3843 581 3844 585
rect 3838 580 3844 581
rect 3886 584 3892 585
rect 4142 584 4148 585
rect 4406 584 4412 585
rect 4646 584 4652 585
rect 4878 584 4884 585
rect 5094 584 5100 585
rect 5310 584 5316 585
rect 5526 584 5532 585
rect 3886 580 3887 584
rect 3891 580 3892 584
rect 3886 579 3892 580
rect 3982 583 3989 584
rect 3982 579 3983 583
rect 3988 579 3989 583
rect 4142 580 4143 584
rect 4147 580 4148 584
rect 4142 579 4148 580
rect 4238 583 4245 584
rect 4238 579 4239 583
rect 4244 579 4245 583
rect 4406 580 4407 584
rect 4411 580 4412 584
rect 4406 579 4412 580
rect 4502 583 4509 584
rect 4502 579 4503 583
rect 4508 579 4509 583
rect 4646 580 4647 584
rect 4651 580 4652 584
rect 4646 579 4652 580
rect 4743 583 4749 584
rect 4743 579 4744 583
rect 4748 582 4749 583
rect 4766 583 4772 584
rect 4766 582 4767 583
rect 4748 580 4767 582
rect 4748 579 4749 580
rect 3982 578 3989 579
rect 4238 578 4245 579
rect 4502 578 4509 579
rect 4743 578 4749 579
rect 4766 579 4767 580
rect 4771 579 4772 583
rect 4878 580 4879 584
rect 4883 580 4884 584
rect 4878 579 4884 580
rect 4975 583 4984 584
rect 4975 579 4976 583
rect 4983 579 4984 583
rect 5094 580 5095 584
rect 5099 580 5100 584
rect 5094 579 5100 580
rect 5191 583 5200 584
rect 5191 579 5192 583
rect 5199 579 5200 583
rect 5310 580 5311 584
rect 5315 580 5316 584
rect 5310 579 5316 580
rect 5402 583 5413 584
rect 5402 579 5403 583
rect 5407 579 5408 583
rect 5412 579 5413 583
rect 5526 580 5527 584
rect 5531 580 5532 584
rect 5526 579 5532 580
rect 5622 583 5629 584
rect 5622 579 5623 583
rect 5628 579 5629 583
rect 5662 581 5663 585
rect 5667 581 5668 585
rect 5662 580 5668 581
rect 4766 578 4772 579
rect 4975 578 4984 579
rect 5191 578 5200 579
rect 5402 578 5413 579
rect 5622 578 5629 579
rect 1974 573 1980 574
rect 3798 573 3804 574
rect 1974 569 1975 573
rect 1979 569 1980 573
rect 1974 568 1980 569
rect 3270 572 3276 573
rect 3406 572 3412 573
rect 3542 572 3548 573
rect 3678 572 3684 573
rect 3270 568 3271 572
rect 3275 568 3276 572
rect 3270 567 3276 568
rect 3367 571 3376 572
rect 3367 567 3368 571
rect 3375 567 3376 571
rect 3406 568 3407 572
rect 3411 568 3412 572
rect 3406 567 3412 568
rect 3503 571 3512 572
rect 3503 567 3504 571
rect 3511 567 3512 571
rect 3542 568 3543 572
rect 3547 568 3548 572
rect 3542 567 3548 568
rect 3639 571 3648 572
rect 3639 567 3640 571
rect 3647 567 3648 571
rect 3678 568 3679 572
rect 3683 568 3684 572
rect 3678 567 3684 568
rect 3774 571 3781 572
rect 3774 567 3775 571
rect 3780 567 3781 571
rect 3798 569 3799 573
rect 3803 569 3804 573
rect 3858 569 3864 570
rect 3798 568 3804 569
rect 3838 568 3844 569
rect 3367 566 3376 567
rect 3503 566 3512 567
rect 3639 566 3648 567
rect 3774 566 3781 567
rect 3838 564 3839 568
rect 3843 564 3844 568
rect 3858 565 3859 569
rect 3863 565 3864 569
rect 3858 564 3864 565
rect 4114 569 4120 570
rect 4114 565 4115 569
rect 4119 565 4120 569
rect 4114 564 4120 565
rect 4378 569 4384 570
rect 4378 565 4379 569
rect 4383 565 4384 569
rect 4378 564 4384 565
rect 4618 569 4624 570
rect 4618 565 4619 569
rect 4623 565 4624 569
rect 4618 564 4624 565
rect 4850 569 4856 570
rect 4850 565 4851 569
rect 4855 565 4856 569
rect 4850 564 4856 565
rect 5066 569 5072 570
rect 5066 565 5067 569
rect 5071 565 5072 569
rect 5066 564 5072 565
rect 5282 569 5288 570
rect 5282 565 5283 569
rect 5287 565 5288 569
rect 5282 564 5288 565
rect 5498 569 5504 570
rect 5498 565 5499 569
rect 5503 565 5504 569
rect 5498 564 5504 565
rect 5662 568 5668 569
rect 5662 564 5663 568
rect 5667 564 5668 568
rect 3838 563 3844 564
rect 5662 563 5668 564
rect 3242 557 3248 558
rect 1974 556 1980 557
rect 1974 552 1975 556
rect 1979 552 1980 556
rect 3242 553 3243 557
rect 3247 553 3248 557
rect 3242 552 3248 553
rect 3378 557 3384 558
rect 3378 553 3379 557
rect 3383 553 3384 557
rect 3378 552 3384 553
rect 3514 557 3520 558
rect 3514 553 3515 557
rect 3519 553 3520 557
rect 3514 552 3520 553
rect 3650 557 3656 558
rect 3650 553 3651 557
rect 3655 553 3656 557
rect 3650 552 3656 553
rect 3798 556 3804 557
rect 3798 552 3799 556
rect 3803 552 3804 556
rect 1974 551 1980 552
rect 3798 551 3804 552
rect 4714 555 4720 556
rect 4714 551 4715 555
rect 4719 554 4720 555
rect 5346 555 5352 556
rect 5346 554 5347 555
rect 4719 552 5347 554
rect 4719 551 4720 552
rect 4714 550 4720 551
rect 5346 551 5347 552
rect 5351 551 5352 555
rect 5346 550 5352 551
rect 110 549 116 550
rect 1934 549 1940 550
rect 110 545 111 549
rect 115 545 116 549
rect 110 544 116 545
rect 158 548 164 549
rect 374 548 380 549
rect 598 548 604 549
rect 806 548 812 549
rect 998 548 1004 549
rect 1174 548 1180 549
rect 1342 548 1348 549
rect 1510 548 1516 549
rect 1670 548 1676 549
rect 1814 548 1820 549
rect 158 544 159 548
rect 163 544 164 548
rect 158 543 164 544
rect 254 547 261 548
rect 254 543 255 547
rect 260 543 261 547
rect 374 544 375 548
rect 379 544 380 548
rect 374 543 380 544
rect 466 547 477 548
rect 466 543 467 547
rect 471 543 472 547
rect 476 543 477 547
rect 598 544 599 548
rect 603 544 604 548
rect 598 543 604 544
rect 695 547 704 548
rect 695 543 696 547
rect 703 543 704 547
rect 806 544 807 548
rect 811 544 812 548
rect 806 543 812 544
rect 903 547 909 548
rect 903 543 904 547
rect 908 546 909 547
rect 934 547 940 548
rect 934 546 935 547
rect 908 544 935 546
rect 908 543 909 544
rect 254 542 261 543
rect 466 542 477 543
rect 695 542 704 543
rect 903 542 909 543
rect 934 543 935 544
rect 939 543 940 547
rect 998 544 999 548
rect 1003 544 1004 548
rect 998 543 1004 544
rect 1094 547 1101 548
rect 1094 543 1095 547
rect 1100 543 1101 547
rect 1174 544 1175 548
rect 1179 544 1180 548
rect 1174 543 1180 544
rect 1271 547 1280 548
rect 1271 543 1272 547
rect 1279 543 1280 547
rect 1342 544 1343 548
rect 1347 544 1348 548
rect 1342 543 1348 544
rect 1439 547 1448 548
rect 1439 543 1440 547
rect 1447 543 1448 547
rect 1510 544 1511 548
rect 1515 544 1516 548
rect 1510 543 1516 544
rect 1607 547 1616 548
rect 1607 543 1608 547
rect 1615 543 1616 547
rect 1670 544 1671 548
rect 1675 544 1676 548
rect 1670 543 1676 544
rect 1767 547 1776 548
rect 1767 543 1768 547
rect 1775 543 1776 547
rect 1814 544 1815 548
rect 1819 544 1820 548
rect 1814 543 1820 544
rect 1911 547 1917 548
rect 1911 543 1912 547
rect 1916 546 1917 547
rect 1926 547 1932 548
rect 1926 546 1927 547
rect 1916 544 1927 546
rect 1916 543 1917 544
rect 934 542 940 543
rect 1094 542 1101 543
rect 1271 542 1280 543
rect 1439 542 1448 543
rect 1607 542 1616 543
rect 1767 542 1776 543
rect 1911 542 1917 543
rect 1926 543 1927 544
rect 1931 543 1932 547
rect 1934 545 1935 549
rect 1939 545 1940 549
rect 1934 544 1940 545
rect 4778 547 4784 548
rect 1926 542 1932 543
rect 4778 543 4779 547
rect 4783 546 4784 547
rect 5402 547 5408 548
rect 5402 546 5403 547
rect 4783 544 5403 546
rect 4783 543 4784 544
rect 4778 542 4784 543
rect 5402 543 5403 544
rect 5407 543 5408 547
rect 5402 542 5408 543
rect 130 533 136 534
rect 110 532 116 533
rect 110 528 111 532
rect 115 528 116 532
rect 130 529 131 533
rect 135 529 136 533
rect 130 528 136 529
rect 346 533 352 534
rect 346 529 347 533
rect 351 529 352 533
rect 346 528 352 529
rect 570 533 576 534
rect 570 529 571 533
rect 575 529 576 533
rect 570 528 576 529
rect 778 533 784 534
rect 778 529 779 533
rect 783 529 784 533
rect 778 528 784 529
rect 970 533 976 534
rect 970 529 971 533
rect 975 529 976 533
rect 970 528 976 529
rect 1146 533 1152 534
rect 1146 529 1147 533
rect 1151 529 1152 533
rect 1146 528 1152 529
rect 1314 533 1320 534
rect 1314 529 1315 533
rect 1319 529 1320 533
rect 1314 528 1320 529
rect 1482 533 1488 534
rect 1482 529 1483 533
rect 1487 529 1488 533
rect 1482 528 1488 529
rect 1642 533 1648 534
rect 1642 529 1643 533
rect 1647 529 1648 533
rect 1642 528 1648 529
rect 1786 533 1792 534
rect 1786 529 1787 533
rect 1791 529 1792 533
rect 1786 528 1792 529
rect 1934 532 1940 533
rect 1934 528 1935 532
rect 1939 528 1940 532
rect 110 527 116 528
rect 1934 527 1940 528
rect 4014 519 4020 520
rect 3956 510 3958 517
rect 4014 515 4015 519
rect 4019 518 4020 519
rect 4446 519 4452 520
rect 4019 516 4121 518
rect 4019 515 4020 516
rect 4014 514 4020 515
rect 4446 515 4447 519
rect 4451 515 4452 519
rect 4446 514 4452 515
rect 4714 519 4720 520
rect 4714 515 4715 519
rect 4719 515 4720 519
rect 4714 514 4720 515
rect 4766 519 4772 520
rect 4766 515 4767 519
rect 4771 518 4772 519
rect 4978 519 4984 520
rect 4771 516 4857 518
rect 4771 515 4772 516
rect 4766 514 4772 515
rect 4978 515 4979 519
rect 4983 518 4984 519
rect 5194 519 5200 520
rect 4983 516 5073 518
rect 4983 515 4984 516
rect 4978 514 4984 515
rect 5194 515 5195 519
rect 5199 518 5200 519
rect 5582 519 5588 520
rect 5199 516 5289 518
rect 5199 515 5200 516
rect 5194 514 5200 515
rect 5582 515 5583 519
rect 5587 515 5588 519
rect 5582 514 5588 515
rect 4238 511 4244 512
rect 4238 510 4239 511
rect 3956 508 4239 510
rect 3370 507 3376 508
rect 3340 498 3342 505
rect 3370 503 3371 507
rect 3375 506 3376 507
rect 3506 507 3512 508
rect 3375 504 3385 506
rect 3375 503 3376 504
rect 3370 502 3376 503
rect 3506 503 3507 507
rect 3511 506 3512 507
rect 3642 507 3648 508
rect 3511 504 3521 506
rect 3511 503 3512 504
rect 3506 502 3512 503
rect 3642 503 3643 507
rect 3647 506 3648 507
rect 4238 507 4239 508
rect 4243 507 4244 511
rect 4238 506 4244 507
rect 3647 504 3657 506
rect 3647 503 3648 504
rect 3642 502 3648 503
rect 3658 499 3664 500
rect 3658 498 3659 499
rect 3340 496 3659 498
rect 3658 495 3659 496
rect 3663 495 3664 499
rect 3658 494 3664 495
rect 734 491 740 492
rect 734 490 735 491
rect 668 488 735 490
rect 335 483 341 484
rect 229 480 261 482
rect 259 474 261 480
rect 335 479 336 483
rect 340 482 341 483
rect 340 480 353 482
rect 668 481 670 488
rect 734 487 735 488
rect 739 487 740 491
rect 734 486 740 487
rect 698 483 704 484
rect 340 479 341 480
rect 335 478 341 479
rect 698 479 699 483
rect 703 482 704 483
rect 934 483 940 484
rect 703 480 785 482
rect 703 479 704 480
rect 698 478 704 479
rect 934 479 935 483
rect 939 482 940 483
rect 1274 483 1280 484
rect 939 480 977 482
rect 939 479 940 480
rect 934 478 940 479
rect 466 475 472 476
rect 466 474 467 475
rect 259 472 467 474
rect 466 471 467 472
rect 471 471 472 475
rect 1244 474 1246 481
rect 1274 479 1275 483
rect 1279 482 1280 483
rect 1442 483 1448 484
rect 1279 480 1321 482
rect 1279 479 1280 480
rect 1274 478 1280 479
rect 1442 479 1443 483
rect 1447 482 1448 483
rect 1610 483 1616 484
rect 1447 480 1489 482
rect 1447 479 1448 480
rect 1442 478 1448 479
rect 1610 479 1611 483
rect 1615 482 1616 483
rect 1770 483 1776 484
rect 1615 480 1649 482
rect 1615 479 1616 480
rect 1610 478 1616 479
rect 1770 479 1771 483
rect 1775 482 1776 483
rect 1775 480 1793 482
rect 1775 479 1776 480
rect 1770 478 1776 479
rect 1910 475 1916 476
rect 1910 474 1911 475
rect 1244 472 1911 474
rect 466 470 472 471
rect 1910 471 1911 472
rect 1915 471 1916 475
rect 1910 470 1916 471
rect 4162 471 4168 472
rect 4162 470 4163 471
rect 3989 468 4163 470
rect 4162 467 4163 468
rect 4167 467 4168 471
rect 4294 471 4300 472
rect 4294 470 4295 471
rect 4269 468 4295 470
rect 4162 466 4168 467
rect 4294 467 4295 468
rect 4299 467 4300 471
rect 4294 466 4300 467
rect 4502 471 4508 472
rect 4502 467 4503 471
rect 4507 467 4508 471
rect 4502 466 4508 467
rect 4778 471 4784 472
rect 4778 467 4779 471
rect 4783 467 4784 471
rect 4778 466 4784 467
rect 4914 467 4920 468
rect 4914 463 4915 467
rect 4919 463 4920 467
rect 4914 462 4920 463
rect 5130 467 5136 468
rect 5130 463 5131 467
rect 5135 463 5136 467
rect 5130 462 5136 463
rect 5338 467 5344 468
rect 5338 463 5339 467
rect 5343 463 5344 467
rect 5338 462 5344 463
rect 5522 467 5528 468
rect 5522 463 5523 467
rect 5527 463 5528 467
rect 5522 462 5528 463
rect 607 459 613 460
rect 607 458 608 459
rect 432 456 608 458
rect 432 450 434 456
rect 607 455 608 456
rect 612 455 613 459
rect 607 454 613 455
rect 1926 455 1932 456
rect 598 451 604 452
rect 598 450 599 451
rect 293 448 434 450
rect 573 448 599 450
rect 598 447 599 448
rect 603 447 604 451
rect 943 451 949 452
rect 943 450 944 451
rect 853 448 944 450
rect 598 446 604 447
rect 943 447 944 448
rect 948 447 949 451
rect 943 446 949 447
rect 1094 451 1100 452
rect 1094 447 1095 451
rect 1099 447 1100 451
rect 1926 451 1927 455
rect 1931 454 1932 455
rect 3014 455 3020 456
rect 1931 452 2001 454
rect 1931 451 1932 452
rect 1926 450 1932 451
rect 2162 451 2168 452
rect 1094 446 1100 447
rect 1338 447 1344 448
rect 1338 443 1339 447
rect 1343 443 1344 447
rect 2162 447 2163 451
rect 2167 447 2168 451
rect 2162 446 2168 447
rect 2354 451 2360 452
rect 2354 447 2355 451
rect 2359 447 2360 451
rect 2354 446 2360 447
rect 2546 451 2552 452
rect 2546 447 2547 451
rect 2551 447 2552 451
rect 2546 446 2552 447
rect 2746 451 2752 452
rect 2746 447 2747 451
rect 2751 447 2752 451
rect 3014 451 3015 455
rect 3019 451 3020 455
rect 3014 450 3020 451
rect 3138 451 3144 452
rect 2746 446 2752 447
rect 3138 447 3139 451
rect 3143 447 3144 451
rect 3138 446 3144 447
rect 3338 451 3344 452
rect 3338 447 3339 451
rect 3343 447 3344 451
rect 3338 446 3344 447
rect 3538 451 3544 452
rect 3538 447 3539 451
rect 3543 447 3544 451
rect 3538 446 3544 447
rect 1338 442 1344 443
rect 3838 420 3844 421
rect 5662 420 5668 421
rect 3838 416 3839 420
rect 3843 416 3844 420
rect 3838 415 3844 416
rect 3890 419 3896 420
rect 3890 415 3891 419
rect 3895 415 3896 419
rect 3890 414 3896 415
rect 4170 419 4176 420
rect 4170 415 4171 419
rect 4175 415 4176 419
rect 4170 414 4176 415
rect 4434 419 4440 420
rect 4434 415 4435 419
rect 4439 415 4440 419
rect 4434 414 4440 415
rect 4682 419 4688 420
rect 4682 415 4683 419
rect 4687 415 4688 419
rect 4682 414 4688 415
rect 4906 419 4912 420
rect 4906 415 4907 419
rect 4911 415 4912 419
rect 4906 414 4912 415
rect 5122 419 5128 420
rect 5122 415 5123 419
rect 5127 415 5128 419
rect 5122 414 5128 415
rect 5330 419 5336 420
rect 5330 415 5331 419
rect 5335 415 5336 419
rect 5330 414 5336 415
rect 5514 419 5520 420
rect 5514 415 5515 419
rect 5519 415 5520 419
rect 5662 416 5663 420
rect 5667 416 5668 420
rect 5662 415 5668 416
rect 5514 414 5520 415
rect 4162 411 4168 412
rect 4162 407 4163 411
rect 4167 410 4168 411
rect 4167 408 4298 410
rect 4167 407 4168 408
rect 4162 406 4168 407
rect 1974 404 1980 405
rect 3798 404 3804 405
rect 3918 404 3924 405
rect 4198 404 4204 405
rect 4296 404 4298 408
rect 4462 404 4468 405
rect 4710 404 4716 405
rect 4934 404 4940 405
rect 5150 404 5156 405
rect 5358 404 5364 405
rect 5542 404 5548 405
rect 110 400 116 401
rect 1934 400 1940 401
rect 110 396 111 400
rect 115 396 116 400
rect 110 395 116 396
rect 194 399 200 400
rect 194 395 195 399
rect 199 395 200 399
rect 194 394 200 395
rect 474 399 480 400
rect 474 395 475 399
rect 479 395 480 399
rect 474 394 480 395
rect 754 399 760 400
rect 754 395 755 399
rect 759 395 760 399
rect 754 394 760 395
rect 1042 399 1048 400
rect 1042 395 1043 399
rect 1047 395 1048 399
rect 1042 394 1048 395
rect 1330 399 1336 400
rect 1330 395 1331 399
rect 1335 395 1336 399
rect 1934 396 1935 400
rect 1939 396 1940 400
rect 1974 400 1975 404
rect 1979 400 1980 404
rect 1974 399 1980 400
rect 1994 403 2000 404
rect 1994 399 1995 403
rect 1999 399 2000 403
rect 1994 398 2000 399
rect 2154 403 2160 404
rect 2154 399 2155 403
rect 2159 399 2160 403
rect 2154 398 2160 399
rect 2346 403 2352 404
rect 2346 399 2347 403
rect 2351 399 2352 403
rect 2346 398 2352 399
rect 2538 403 2544 404
rect 2538 399 2539 403
rect 2543 399 2544 403
rect 2538 398 2544 399
rect 2738 403 2744 404
rect 2738 399 2739 403
rect 2743 399 2744 403
rect 2738 398 2744 399
rect 2930 403 2936 404
rect 2930 399 2931 403
rect 2935 399 2936 403
rect 2930 398 2936 399
rect 3130 403 3136 404
rect 3130 399 3131 403
rect 3135 399 3136 403
rect 3130 398 3136 399
rect 3330 403 3336 404
rect 3330 399 3331 403
rect 3335 399 3336 403
rect 3330 398 3336 399
rect 3530 403 3536 404
rect 3530 399 3531 403
rect 3535 399 3536 403
rect 3798 400 3799 404
rect 3803 400 3804 404
rect 3798 399 3804 400
rect 3838 403 3844 404
rect 3838 399 3839 403
rect 3843 399 3844 403
rect 3918 400 3919 404
rect 3923 400 3924 404
rect 3918 399 3924 400
rect 4014 403 4021 404
rect 4014 399 4015 403
rect 4020 399 4021 403
rect 4198 400 4199 404
rect 4203 400 4204 404
rect 4198 399 4204 400
rect 4295 403 4301 404
rect 4295 399 4296 403
rect 4300 399 4301 403
rect 4462 400 4463 404
rect 4467 400 4468 404
rect 4462 399 4468 400
rect 4554 403 4565 404
rect 4554 399 4555 403
rect 4559 399 4560 403
rect 4564 399 4565 403
rect 4710 400 4711 404
rect 4715 400 4716 404
rect 4710 399 4716 400
rect 4807 403 4813 404
rect 4807 399 4808 403
rect 4812 402 4813 403
rect 4914 403 4920 404
rect 4914 402 4915 403
rect 4812 400 4915 402
rect 4812 399 4813 400
rect 3530 398 3536 399
rect 3838 398 3844 399
rect 4014 398 4021 399
rect 4295 398 4301 399
rect 4554 398 4565 399
rect 4807 398 4813 399
rect 4914 399 4915 400
rect 4919 399 4920 403
rect 4934 400 4935 404
rect 4939 400 4940 404
rect 4934 399 4940 400
rect 5031 403 5037 404
rect 5031 399 5032 403
rect 5036 402 5037 403
rect 5130 403 5136 404
rect 5130 402 5131 403
rect 5036 400 5131 402
rect 5036 399 5037 400
rect 4914 398 4920 399
rect 5031 398 5037 399
rect 5130 399 5131 400
rect 5135 399 5136 403
rect 5150 400 5151 404
rect 5155 400 5156 404
rect 5150 399 5156 400
rect 5247 403 5253 404
rect 5247 399 5248 403
rect 5252 402 5253 403
rect 5338 403 5344 404
rect 5338 402 5339 403
rect 5252 400 5339 402
rect 5252 399 5253 400
rect 5130 398 5136 399
rect 5247 398 5253 399
rect 5338 399 5339 400
rect 5343 399 5344 403
rect 5358 400 5359 404
rect 5363 400 5364 404
rect 5358 399 5364 400
rect 5455 403 5461 404
rect 5455 399 5456 403
rect 5460 402 5461 403
rect 5522 403 5528 404
rect 5522 402 5523 403
rect 5460 400 5523 402
rect 5460 399 5461 400
rect 5338 398 5344 399
rect 5455 398 5461 399
rect 5522 399 5523 400
rect 5527 399 5528 403
rect 5542 400 5543 404
rect 5547 400 5548 404
rect 5542 399 5548 400
rect 5638 403 5645 404
rect 5638 399 5639 403
rect 5644 399 5645 403
rect 5522 398 5528 399
rect 5638 398 5645 399
rect 5662 403 5668 404
rect 5662 399 5663 403
rect 5667 399 5668 403
rect 5662 398 5668 399
rect 1934 395 1940 396
rect 1330 394 1336 395
rect 943 391 949 392
rect 943 387 944 391
rect 948 390 949 391
rect 948 388 1458 390
rect 2022 388 2028 389
rect 2182 388 2188 389
rect 2374 388 2380 389
rect 2566 388 2572 389
rect 2766 388 2772 389
rect 2958 388 2964 389
rect 3158 388 3164 389
rect 3358 388 3364 389
rect 3558 388 3564 389
rect 948 387 949 388
rect 943 386 949 387
rect 1456 386 1458 388
rect 1974 387 1980 388
rect 1455 385 1461 386
rect 222 384 228 385
rect 502 384 508 385
rect 782 384 788 385
rect 1070 384 1076 385
rect 1358 384 1364 385
rect 110 383 116 384
rect 110 379 111 383
rect 115 379 116 383
rect 222 380 223 384
rect 227 380 228 384
rect 222 379 228 380
rect 319 383 325 384
rect 319 379 320 383
rect 324 382 325 383
rect 335 383 341 384
rect 335 382 336 383
rect 324 380 336 382
rect 324 379 325 380
rect 110 378 116 379
rect 319 378 325 379
rect 335 379 336 380
rect 340 379 341 383
rect 502 380 503 384
rect 507 380 508 384
rect 502 379 508 380
rect 599 383 605 384
rect 599 379 600 383
rect 604 382 605 383
rect 607 383 613 384
rect 607 382 608 383
rect 604 380 608 382
rect 604 379 605 380
rect 335 378 341 379
rect 599 378 605 379
rect 607 379 608 380
rect 612 379 613 383
rect 782 380 783 384
rect 787 380 788 384
rect 782 379 788 380
rect 878 383 885 384
rect 878 379 879 383
rect 884 379 885 383
rect 1070 380 1071 384
rect 1075 380 1076 384
rect 1070 379 1076 380
rect 1167 383 1173 384
rect 1167 379 1168 383
rect 1172 382 1173 383
rect 1338 383 1344 384
rect 1338 382 1339 383
rect 1172 380 1339 382
rect 1172 379 1173 380
rect 607 378 613 379
rect 878 378 885 379
rect 1167 378 1173 379
rect 1338 379 1339 380
rect 1343 379 1344 383
rect 1358 380 1359 384
rect 1363 380 1364 384
rect 1455 381 1456 385
rect 1460 381 1461 385
rect 1455 380 1461 381
rect 1934 383 1940 384
rect 1358 379 1364 380
rect 1934 379 1935 383
rect 1939 379 1940 383
rect 1974 383 1975 387
rect 1979 383 1980 387
rect 2022 384 2023 388
rect 2027 384 2028 388
rect 2022 383 2028 384
rect 2119 387 2125 388
rect 2119 383 2120 387
rect 2124 386 2125 387
rect 2162 387 2168 388
rect 2162 386 2163 387
rect 2124 384 2163 386
rect 2124 383 2125 384
rect 1974 382 1980 383
rect 2119 382 2125 383
rect 2162 383 2163 384
rect 2167 383 2168 387
rect 2182 384 2183 388
rect 2187 384 2188 388
rect 2182 383 2188 384
rect 2279 387 2285 388
rect 2279 383 2280 387
rect 2284 386 2285 387
rect 2354 387 2360 388
rect 2354 386 2355 387
rect 2284 384 2355 386
rect 2284 383 2285 384
rect 2162 382 2168 383
rect 2279 382 2285 383
rect 2354 383 2355 384
rect 2359 383 2360 387
rect 2374 384 2375 388
rect 2379 384 2380 388
rect 2374 383 2380 384
rect 2471 387 2477 388
rect 2471 383 2472 387
rect 2476 386 2477 387
rect 2546 387 2552 388
rect 2546 386 2547 387
rect 2476 384 2547 386
rect 2476 383 2477 384
rect 2354 382 2360 383
rect 2471 382 2477 383
rect 2546 383 2547 384
rect 2551 383 2552 387
rect 2566 384 2567 388
rect 2571 384 2572 388
rect 2566 383 2572 384
rect 2663 387 2669 388
rect 2663 383 2664 387
rect 2668 386 2669 387
rect 2746 387 2752 388
rect 2746 386 2747 387
rect 2668 384 2747 386
rect 2668 383 2669 384
rect 2546 382 2552 383
rect 2663 382 2669 383
rect 2746 383 2747 384
rect 2751 383 2752 387
rect 2766 384 2767 388
rect 2771 384 2772 388
rect 2766 383 2772 384
rect 2858 387 2869 388
rect 2858 383 2859 387
rect 2863 383 2864 387
rect 2868 383 2869 387
rect 2958 384 2959 388
rect 2963 384 2964 388
rect 2958 383 2964 384
rect 3055 387 3061 388
rect 3055 383 3056 387
rect 3060 386 3061 387
rect 3138 387 3144 388
rect 3138 386 3139 387
rect 3060 384 3139 386
rect 3060 383 3061 384
rect 2746 382 2752 383
rect 2858 382 2869 383
rect 3055 382 3061 383
rect 3138 383 3139 384
rect 3143 383 3144 387
rect 3158 384 3159 388
rect 3163 384 3164 388
rect 3158 383 3164 384
rect 3255 387 3261 388
rect 3255 383 3256 387
rect 3260 386 3261 387
rect 3338 387 3344 388
rect 3338 386 3339 387
rect 3260 384 3339 386
rect 3260 383 3261 384
rect 3138 382 3144 383
rect 3255 382 3261 383
rect 3338 383 3339 384
rect 3343 383 3344 387
rect 3358 384 3359 388
rect 3363 384 3364 388
rect 3358 383 3364 384
rect 3455 387 3461 388
rect 3455 383 3456 387
rect 3460 386 3461 387
rect 3538 387 3544 388
rect 3538 386 3539 387
rect 3460 384 3539 386
rect 3460 383 3461 384
rect 3338 382 3344 383
rect 3455 382 3461 383
rect 3538 383 3539 384
rect 3543 383 3544 387
rect 3558 384 3559 388
rect 3563 384 3564 388
rect 3558 383 3564 384
rect 3655 387 3664 388
rect 3655 383 3656 387
rect 3663 383 3664 387
rect 3538 382 3544 383
rect 3655 382 3664 383
rect 3798 387 3804 388
rect 3798 383 3799 387
rect 3803 383 3804 387
rect 3798 382 3804 383
rect 1338 378 1344 379
rect 1934 378 1940 379
rect 3838 341 3844 342
rect 5662 341 5668 342
rect 3838 337 3839 341
rect 3843 337 3844 341
rect 3838 336 3844 337
rect 4006 340 4012 341
rect 4198 340 4204 341
rect 4422 340 4428 341
rect 4678 340 4684 341
rect 4966 340 4972 341
rect 5262 340 5268 341
rect 5542 340 5548 341
rect 4006 336 4007 340
rect 4011 336 4012 340
rect 4006 335 4012 336
rect 4103 339 4109 340
rect 4103 335 4104 339
rect 4108 338 4109 339
rect 4134 339 4140 340
rect 4134 338 4135 339
rect 4108 336 4135 338
rect 4108 335 4109 336
rect 4103 334 4109 335
rect 4134 335 4135 336
rect 4139 335 4140 339
rect 4198 336 4199 340
rect 4203 336 4204 340
rect 4198 335 4204 336
rect 4294 339 4301 340
rect 4294 335 4295 339
rect 4300 335 4301 339
rect 4422 336 4423 340
rect 4427 336 4428 340
rect 4422 335 4428 336
rect 4519 339 4525 340
rect 4519 335 4520 339
rect 4524 338 4525 339
rect 4558 339 4564 340
rect 4558 338 4559 339
rect 4524 336 4559 338
rect 4524 335 4525 336
rect 4134 334 4140 335
rect 4294 334 4301 335
rect 4519 334 4525 335
rect 4558 335 4559 336
rect 4563 335 4564 339
rect 4678 336 4679 340
rect 4683 336 4684 340
rect 4678 335 4684 336
rect 4775 339 4784 340
rect 4775 335 4776 339
rect 4783 335 4784 339
rect 4966 336 4967 340
rect 4971 336 4972 340
rect 4966 335 4972 336
rect 5063 339 5072 340
rect 5063 335 5064 339
rect 5071 335 5072 339
rect 5262 336 5263 340
rect 5267 336 5268 340
rect 5262 335 5268 336
rect 5354 339 5365 340
rect 5354 335 5355 339
rect 5359 335 5360 339
rect 5364 335 5365 339
rect 5542 336 5543 340
rect 5547 336 5548 340
rect 5542 335 5548 336
rect 5634 339 5645 340
rect 5634 335 5635 339
rect 5639 335 5640 339
rect 5644 335 5645 339
rect 5662 337 5663 341
rect 5667 337 5668 341
rect 5662 336 5668 337
rect 4558 334 4564 335
rect 4775 334 4784 335
rect 5063 334 5072 335
rect 5354 334 5365 335
rect 5634 334 5645 335
rect 110 325 116 326
rect 1934 325 1940 326
rect 3978 325 3984 326
rect 110 321 111 325
rect 115 321 116 325
rect 110 320 116 321
rect 310 324 316 325
rect 502 324 508 325
rect 694 324 700 325
rect 886 324 892 325
rect 1078 324 1084 325
rect 310 320 311 324
rect 315 320 316 324
rect 310 319 316 320
rect 407 323 413 324
rect 407 319 408 323
rect 412 322 413 323
rect 430 323 436 324
rect 430 322 431 323
rect 412 320 431 322
rect 412 319 413 320
rect 407 318 413 319
rect 430 319 431 320
rect 435 319 436 323
rect 502 320 503 324
rect 507 320 508 324
rect 502 319 508 320
rect 598 323 605 324
rect 598 319 599 323
rect 604 319 605 323
rect 694 320 695 324
rect 699 320 700 324
rect 694 319 700 320
rect 791 323 797 324
rect 791 319 792 323
rect 796 322 797 323
rect 799 323 805 324
rect 799 322 800 323
rect 796 320 800 322
rect 796 319 797 320
rect 430 318 436 319
rect 598 318 605 319
rect 791 318 797 319
rect 799 319 800 320
rect 804 319 805 323
rect 886 320 887 324
rect 891 320 892 324
rect 886 319 892 320
rect 983 323 989 324
rect 983 319 984 323
rect 988 322 989 323
rect 991 323 997 324
rect 991 322 992 323
rect 988 320 992 322
rect 988 319 989 320
rect 799 318 805 319
rect 983 318 989 319
rect 991 319 992 320
rect 996 319 997 323
rect 1078 320 1079 324
rect 1083 320 1084 324
rect 1078 319 1084 320
rect 1174 323 1181 324
rect 1174 319 1175 323
rect 1180 319 1181 323
rect 1934 321 1935 325
rect 1939 321 1940 325
rect 1934 320 1940 321
rect 3838 324 3844 325
rect 3838 320 3839 324
rect 3843 320 3844 324
rect 3978 321 3979 325
rect 3983 321 3984 325
rect 3978 320 3984 321
rect 4170 325 4176 326
rect 4170 321 4171 325
rect 4175 321 4176 325
rect 4170 320 4176 321
rect 4394 325 4400 326
rect 4394 321 4395 325
rect 4399 321 4400 325
rect 4394 320 4400 321
rect 4650 325 4656 326
rect 4650 321 4651 325
rect 4655 321 4656 325
rect 4650 320 4656 321
rect 4938 325 4944 326
rect 4938 321 4939 325
rect 4943 321 4944 325
rect 4938 320 4944 321
rect 5234 325 5240 326
rect 5234 321 5235 325
rect 5239 321 5240 325
rect 5234 320 5240 321
rect 5514 325 5520 326
rect 5514 321 5515 325
rect 5519 321 5520 325
rect 5514 320 5520 321
rect 5662 324 5668 325
rect 5662 320 5663 324
rect 5667 320 5668 324
rect 991 318 997 319
rect 1174 318 1181 319
rect 3014 319 3020 320
rect 3838 319 3844 320
rect 5662 319 5668 320
rect 3014 315 3015 319
rect 3019 318 3020 319
rect 3019 316 3618 318
rect 3019 315 3020 316
rect 3014 314 3020 315
rect 282 309 288 310
rect 110 308 116 309
rect 110 304 111 308
rect 115 304 116 308
rect 282 305 283 309
rect 287 305 288 309
rect 282 304 288 305
rect 474 309 480 310
rect 474 305 475 309
rect 479 305 480 309
rect 474 304 480 305
rect 666 309 672 310
rect 666 305 667 309
rect 671 305 672 309
rect 666 304 672 305
rect 858 309 864 310
rect 858 305 859 309
rect 863 305 864 309
rect 858 304 864 305
rect 1050 309 1056 310
rect 1050 305 1051 309
rect 1055 305 1056 309
rect 1050 304 1056 305
rect 1934 308 1940 309
rect 1934 304 1935 308
rect 1939 304 1940 308
rect 110 303 116 304
rect 1934 303 1940 304
rect 1974 305 1980 306
rect 1974 301 1975 305
rect 1979 301 1980 305
rect 1974 300 1980 301
rect 2022 304 2028 305
rect 2158 304 2164 305
rect 2294 304 2300 305
rect 2430 304 2436 305
rect 2566 304 2572 305
rect 2702 304 2708 305
rect 2838 304 2844 305
rect 2974 304 2980 305
rect 3110 304 3116 305
rect 3246 304 3252 305
rect 3382 304 3388 305
rect 3518 304 3524 305
rect 3616 304 3618 316
rect 3798 305 3804 306
rect 2022 300 2023 304
rect 2027 300 2028 304
rect 2022 299 2028 300
rect 2119 303 2128 304
rect 2119 299 2120 303
rect 2127 299 2128 303
rect 2158 300 2159 304
rect 2163 300 2164 304
rect 2158 299 2164 300
rect 2255 303 2264 304
rect 2255 299 2256 303
rect 2263 299 2264 303
rect 2294 300 2295 304
rect 2299 300 2300 304
rect 2294 299 2300 300
rect 2391 303 2400 304
rect 2391 299 2392 303
rect 2399 299 2400 303
rect 2430 300 2431 304
rect 2435 300 2436 304
rect 2430 299 2436 300
rect 2527 303 2536 304
rect 2527 299 2528 303
rect 2535 299 2536 303
rect 2566 300 2567 304
rect 2571 300 2572 304
rect 2566 299 2572 300
rect 2663 303 2672 304
rect 2663 299 2664 303
rect 2671 299 2672 303
rect 2702 300 2703 304
rect 2707 300 2708 304
rect 2702 299 2708 300
rect 2794 303 2805 304
rect 2794 299 2795 303
rect 2799 299 2800 303
rect 2804 299 2805 303
rect 2838 300 2839 304
rect 2843 300 2844 304
rect 2838 299 2844 300
rect 2935 303 2944 304
rect 2935 299 2936 303
rect 2943 299 2944 303
rect 2974 300 2975 304
rect 2979 300 2980 304
rect 2974 299 2980 300
rect 3071 303 3080 304
rect 3071 299 3072 303
rect 3079 299 3080 303
rect 3110 300 3111 304
rect 3115 300 3116 304
rect 3110 299 3116 300
rect 3207 303 3216 304
rect 3207 299 3208 303
rect 3215 299 3216 303
rect 3246 300 3247 304
rect 3251 300 3252 304
rect 3246 299 3252 300
rect 3343 303 3352 304
rect 3343 299 3344 303
rect 3351 299 3352 303
rect 3382 300 3383 304
rect 3387 300 3388 304
rect 3382 299 3388 300
rect 3479 303 3488 304
rect 3479 299 3480 303
rect 3487 299 3488 303
rect 3518 300 3519 304
rect 3523 300 3524 304
rect 3518 299 3524 300
rect 3615 303 3621 304
rect 3615 299 3616 303
rect 3620 299 3621 303
rect 3798 301 3799 305
rect 3803 301 3804 305
rect 3798 300 3804 301
rect 2119 298 2128 299
rect 2255 298 2264 299
rect 2391 298 2400 299
rect 2527 298 2536 299
rect 2663 298 2672 299
rect 2794 298 2805 299
rect 2935 298 2944 299
rect 3071 298 3080 299
rect 3207 298 3216 299
rect 3343 298 3352 299
rect 3479 298 3488 299
rect 3615 298 3621 299
rect 1994 289 2000 290
rect 1974 288 1980 289
rect 1974 284 1975 288
rect 1979 284 1980 288
rect 1994 285 1995 289
rect 1999 285 2000 289
rect 1994 284 2000 285
rect 2130 289 2136 290
rect 2130 285 2131 289
rect 2135 285 2136 289
rect 2130 284 2136 285
rect 2266 289 2272 290
rect 2266 285 2267 289
rect 2271 285 2272 289
rect 2266 284 2272 285
rect 2402 289 2408 290
rect 2402 285 2403 289
rect 2407 285 2408 289
rect 2402 284 2408 285
rect 2538 289 2544 290
rect 2538 285 2539 289
rect 2543 285 2544 289
rect 2538 284 2544 285
rect 2674 289 2680 290
rect 2674 285 2675 289
rect 2679 285 2680 289
rect 2674 284 2680 285
rect 2810 289 2816 290
rect 2810 285 2811 289
rect 2815 285 2816 289
rect 2810 284 2816 285
rect 2946 289 2952 290
rect 2946 285 2947 289
rect 2951 285 2952 289
rect 2946 284 2952 285
rect 3082 289 3088 290
rect 3082 285 3083 289
rect 3087 285 3088 289
rect 3082 284 3088 285
rect 3218 289 3224 290
rect 3218 285 3219 289
rect 3223 285 3224 289
rect 3218 284 3224 285
rect 3354 289 3360 290
rect 3354 285 3355 289
rect 3359 285 3360 289
rect 3354 284 3360 285
rect 3490 289 3496 290
rect 3490 285 3491 289
rect 3495 285 3496 289
rect 3490 284 3496 285
rect 3798 288 3804 289
rect 3798 284 3799 288
rect 3803 284 3804 288
rect 1974 283 1980 284
rect 2090 283 2096 284
rect 2090 279 2091 283
rect 2095 282 2096 283
rect 2858 283 2864 284
rect 3798 283 3804 284
rect 2858 282 2859 283
rect 2095 280 2859 282
rect 2095 279 2096 280
rect 2090 278 2096 279
rect 2858 279 2859 280
rect 2863 279 2864 283
rect 2858 278 2864 279
rect 4114 275 4120 276
rect 4114 274 4115 275
rect 4077 272 4115 274
rect 4114 271 4115 272
rect 4119 271 4120 275
rect 4114 270 4120 271
rect 4134 275 4140 276
rect 4134 271 4135 275
rect 4139 274 4140 275
rect 4550 275 4556 276
rect 4550 274 4551 275
rect 4139 272 4177 274
rect 4493 272 4551 274
rect 4139 271 4140 272
rect 4134 270 4140 271
rect 4550 271 4551 272
rect 4555 271 4556 275
rect 4550 270 4556 271
rect 4558 275 4564 276
rect 4558 271 4559 275
rect 4563 274 4564 275
rect 4778 275 4784 276
rect 4563 272 4657 274
rect 4563 271 4564 272
rect 4558 270 4564 271
rect 4778 271 4779 275
rect 4783 274 4784 275
rect 5066 275 5072 276
rect 4783 272 4945 274
rect 4783 271 4784 272
rect 4778 270 4784 271
rect 5066 271 5067 275
rect 5071 274 5072 275
rect 5622 275 5628 276
rect 5622 274 5623 275
rect 5071 272 5241 274
rect 5613 272 5623 274
rect 5071 271 5072 272
rect 5066 270 5072 271
rect 5622 271 5623 272
rect 5627 271 5628 275
rect 5622 270 5628 271
rect 386 259 392 260
rect 386 258 387 259
rect 381 256 387 258
rect 386 255 387 256
rect 391 255 392 259
rect 386 254 392 255
rect 430 259 436 260
rect 430 255 431 259
rect 435 258 436 259
rect 878 259 884 260
rect 435 256 481 258
rect 435 255 436 256
rect 430 254 436 255
rect 764 250 766 257
rect 878 255 879 259
rect 883 255 884 259
rect 878 254 884 255
rect 991 259 997 260
rect 991 255 992 259
rect 996 258 997 259
rect 996 256 1057 258
rect 996 255 997 256
rect 991 254 997 255
rect 4722 255 4728 256
rect 1174 251 1180 252
rect 1174 250 1175 251
rect 764 248 1175 250
rect 1174 247 1175 248
rect 1179 247 1180 251
rect 4722 251 4723 255
rect 4727 254 4728 255
rect 5354 255 5360 256
rect 5354 254 5355 255
rect 4727 252 5355 254
rect 4727 251 4728 252
rect 4722 250 4728 251
rect 5354 251 5355 252
rect 5359 251 5360 255
rect 5354 250 5360 251
rect 1174 246 1180 247
rect 2090 239 2096 240
rect 2090 235 2091 239
rect 2095 235 2096 239
rect 2090 234 2096 235
rect 2122 239 2128 240
rect 2122 235 2123 239
rect 2127 238 2128 239
rect 2258 239 2264 240
rect 2127 236 2137 238
rect 2127 235 2128 236
rect 2122 234 2128 235
rect 2258 235 2259 239
rect 2263 238 2264 239
rect 2394 239 2400 240
rect 2263 236 2273 238
rect 2263 235 2264 236
rect 2258 234 2264 235
rect 2394 235 2395 239
rect 2399 238 2400 239
rect 2530 239 2536 240
rect 2399 236 2409 238
rect 2399 235 2400 236
rect 2394 234 2400 235
rect 2530 235 2531 239
rect 2535 238 2536 239
rect 2666 239 2672 240
rect 2535 236 2545 238
rect 2535 235 2536 236
rect 2530 234 2536 235
rect 2666 235 2667 239
rect 2671 238 2672 239
rect 2906 239 2912 240
rect 2671 236 2681 238
rect 2671 235 2672 236
rect 2666 234 2672 235
rect 2906 235 2907 239
rect 2911 235 2912 239
rect 2906 234 2912 235
rect 2938 239 2944 240
rect 2938 235 2939 239
rect 2943 238 2944 239
rect 3074 239 3080 240
rect 2943 236 2953 238
rect 2943 235 2944 236
rect 2938 234 2944 235
rect 3074 235 3075 239
rect 3079 238 3080 239
rect 3210 239 3216 240
rect 3079 236 3089 238
rect 3079 235 3080 236
rect 3074 234 3080 235
rect 3210 235 3211 239
rect 3215 238 3216 239
rect 3346 239 3352 240
rect 3215 236 3225 238
rect 3215 235 3216 236
rect 3210 234 3216 235
rect 3346 235 3347 239
rect 3351 238 3352 239
rect 3482 239 3488 240
rect 3351 236 3361 238
rect 3351 235 3352 236
rect 3346 234 3352 235
rect 3482 235 3483 239
rect 3487 238 3488 239
rect 3487 236 3497 238
rect 3487 235 3488 236
rect 3482 234 3488 235
rect 522 199 528 200
rect 522 198 523 199
rect 259 196 523 198
rect 259 190 261 196
rect 522 195 523 196
rect 527 195 528 199
rect 1206 199 1212 200
rect 1206 198 1207 199
rect 522 194 528 195
rect 792 196 1207 198
rect 666 191 672 192
rect 666 190 667 191
rect 229 188 261 190
rect 637 188 667 190
rect 274 187 280 188
rect 274 183 275 187
rect 279 183 280 187
rect 274 182 280 183
rect 498 187 504 188
rect 498 183 499 187
rect 503 183 504 187
rect 666 187 667 188
rect 671 187 672 191
rect 792 190 794 196
rect 1206 195 1207 196
rect 1211 195 1212 199
rect 4250 199 4256 200
rect 4250 198 4251 199
rect 1206 194 1212 195
rect 3996 196 4251 198
rect 773 188 794 190
rect 799 191 805 192
rect 666 186 672 187
rect 799 187 800 191
rect 804 190 805 191
rect 3996 190 3998 196
rect 4250 195 4251 196
rect 4255 195 4256 199
rect 4250 194 4256 195
rect 4394 191 4400 192
rect 4394 190 4395 191
rect 804 188 817 190
rect 3957 188 3998 190
rect 4365 188 4395 190
rect 804 187 805 188
rect 799 186 805 187
rect 954 187 960 188
rect 498 182 504 183
rect 954 183 955 187
rect 959 183 960 187
rect 954 182 960 183
rect 1090 187 1096 188
rect 1090 183 1091 187
rect 1095 183 1096 187
rect 1090 182 1096 183
rect 4002 187 4008 188
rect 4002 183 4003 187
rect 4007 183 4008 187
rect 4002 182 4008 183
rect 4226 187 4232 188
rect 4226 183 4227 187
rect 4231 183 4232 187
rect 4394 187 4395 188
rect 4399 187 4400 191
rect 4722 191 4728 192
rect 4394 186 4400 187
rect 4530 187 4536 188
rect 4226 182 4232 183
rect 4530 183 4531 187
rect 4535 183 4536 187
rect 4722 187 4723 191
rect 4727 187 4728 191
rect 5502 191 5508 192
rect 5502 190 5503 191
rect 5397 188 5503 190
rect 4722 186 4728 187
rect 4850 187 4856 188
rect 4530 182 4536 183
rect 4850 183 4851 187
rect 4855 183 4856 187
rect 4850 182 4856 183
rect 5074 187 5080 188
rect 5074 183 5075 187
rect 5079 183 5080 187
rect 5502 187 5503 188
rect 5507 187 5508 191
rect 5634 191 5640 192
rect 5634 190 5635 191
rect 5613 188 5635 190
rect 5502 186 5508 187
rect 5634 187 5635 188
rect 5639 187 5640 191
rect 5634 186 5640 187
rect 5074 182 5080 183
rect 2114 175 2120 176
rect 2114 174 2115 175
rect 2093 172 2115 174
rect 2114 171 2115 172
rect 2119 171 2120 175
rect 2114 170 2120 171
rect 2138 171 2144 172
rect 2138 167 2139 171
rect 2143 167 2144 171
rect 2138 166 2144 167
rect 2274 171 2280 172
rect 2274 167 2275 171
rect 2279 167 2280 171
rect 2274 166 2280 167
rect 2410 171 2416 172
rect 2410 167 2411 171
rect 2415 167 2416 171
rect 2410 166 2416 167
rect 2546 171 2552 172
rect 2546 167 2547 171
rect 2551 167 2552 171
rect 2546 166 2552 167
rect 2682 171 2688 172
rect 2682 167 2683 171
rect 2687 167 2688 171
rect 2682 166 2688 167
rect 2818 171 2824 172
rect 2818 167 2819 171
rect 2823 167 2824 171
rect 2818 166 2824 167
rect 2954 171 2960 172
rect 2954 167 2955 171
rect 2959 167 2960 171
rect 2954 166 2960 167
rect 3090 171 3096 172
rect 3090 167 3091 171
rect 3095 167 3096 171
rect 3090 166 3096 167
rect 3226 171 3232 172
rect 3226 167 3227 171
rect 3231 167 3232 171
rect 3226 166 3232 167
rect 3362 171 3368 172
rect 3362 167 3363 171
rect 3367 167 3368 171
rect 3362 166 3368 167
rect 3498 171 3504 172
rect 3498 167 3499 171
rect 3503 167 3504 171
rect 3498 166 3504 167
rect 3634 171 3640 172
rect 3634 167 3635 171
rect 3639 167 3640 171
rect 3634 166 3640 167
rect 498 159 504 160
rect 498 155 499 159
rect 503 158 504 159
rect 658 159 664 160
rect 658 158 659 159
rect 503 156 659 158
rect 503 155 504 156
rect 498 154 504 155
rect 658 155 659 156
rect 663 155 664 159
rect 658 154 664 155
rect 4226 159 4232 160
rect 4226 155 4227 159
rect 4231 158 4232 159
rect 4386 159 4392 160
rect 4386 158 4387 159
rect 4231 156 4387 158
rect 4231 155 4232 156
rect 4226 154 4232 155
rect 4386 155 4387 156
rect 4391 155 4392 159
rect 4386 154 4392 155
rect 4530 155 4536 156
rect 4530 151 4531 155
rect 4535 154 4536 155
rect 5186 155 5192 156
rect 5186 154 5187 155
rect 4535 152 5187 154
rect 4535 151 4536 152
rect 4530 150 4536 151
rect 5186 151 5187 152
rect 5191 151 5192 155
rect 5186 150 5192 151
rect 110 140 116 141
rect 1934 140 1940 141
rect 110 136 111 140
rect 115 136 116 140
rect 110 135 116 136
rect 130 139 136 140
rect 130 135 131 139
rect 135 135 136 139
rect 130 134 136 135
rect 266 139 272 140
rect 266 135 267 139
rect 271 135 272 139
rect 266 134 272 135
rect 402 139 408 140
rect 402 135 403 139
rect 407 135 408 139
rect 402 134 408 135
rect 538 139 544 140
rect 538 135 539 139
rect 543 135 544 139
rect 538 134 544 135
rect 674 139 680 140
rect 674 135 675 139
rect 679 135 680 139
rect 674 134 680 135
rect 810 139 816 140
rect 810 135 811 139
rect 815 135 816 139
rect 810 134 816 135
rect 946 139 952 140
rect 946 135 947 139
rect 951 135 952 139
rect 946 134 952 135
rect 1082 139 1088 140
rect 1082 135 1083 139
rect 1087 135 1088 139
rect 1934 136 1935 140
rect 1939 136 1940 140
rect 1934 135 1940 136
rect 3838 140 3844 141
rect 5662 140 5668 141
rect 3838 136 3839 140
rect 3843 136 3844 140
rect 3838 135 3844 136
rect 3858 139 3864 140
rect 3858 135 3859 139
rect 3863 135 3864 139
rect 1082 134 1088 135
rect 3858 134 3864 135
rect 3994 139 4000 140
rect 3994 135 3995 139
rect 3999 135 4000 139
rect 3994 134 4000 135
rect 4130 139 4136 140
rect 4130 135 4131 139
rect 4135 135 4136 139
rect 4130 134 4136 135
rect 4266 139 4272 140
rect 4266 135 4267 139
rect 4271 135 4272 139
rect 4266 134 4272 135
rect 4434 139 4440 140
rect 4434 135 4435 139
rect 4439 135 4440 139
rect 4434 134 4440 135
rect 4626 139 4632 140
rect 4626 135 4627 139
rect 4631 135 4632 139
rect 4626 134 4632 135
rect 4842 139 4848 140
rect 4842 135 4843 139
rect 4847 135 4848 139
rect 4842 134 4848 135
rect 5066 139 5072 140
rect 5066 135 5067 139
rect 5071 135 5072 139
rect 5066 134 5072 135
rect 5298 139 5304 140
rect 5298 135 5299 139
rect 5303 135 5304 139
rect 5298 134 5304 135
rect 5514 139 5520 140
rect 5514 135 5515 139
rect 5519 135 5520 139
rect 5662 136 5663 140
rect 5667 136 5668 140
rect 5662 135 5668 136
rect 5514 134 5520 135
rect 666 131 672 132
rect 666 127 667 131
rect 671 130 672 131
rect 4394 131 4400 132
rect 671 128 802 130
rect 671 127 672 128
rect 666 126 672 127
rect 800 126 802 128
rect 4394 127 4395 131
rect 4399 130 4400 131
rect 5502 131 5508 132
rect 4399 128 4562 130
rect 4399 127 4400 128
rect 4394 126 4400 127
rect 799 125 805 126
rect 158 124 164 125
rect 294 124 300 125
rect 430 124 436 125
rect 566 124 572 125
rect 702 124 708 125
rect 110 123 116 124
rect 110 119 111 123
rect 115 119 116 123
rect 158 120 159 124
rect 163 120 164 124
rect 158 119 164 120
rect 255 123 261 124
rect 255 119 256 123
rect 260 122 261 123
rect 274 123 280 124
rect 274 122 275 123
rect 260 120 275 122
rect 260 119 261 120
rect 110 118 116 119
rect 255 118 261 119
rect 274 119 275 120
rect 279 119 280 123
rect 294 120 295 124
rect 299 120 300 124
rect 294 119 300 120
rect 386 123 397 124
rect 386 119 387 123
rect 391 119 392 123
rect 396 119 397 123
rect 430 120 431 124
rect 435 120 436 124
rect 430 119 436 120
rect 522 123 533 124
rect 522 119 523 123
rect 527 119 528 123
rect 532 119 533 123
rect 566 120 567 124
rect 571 120 572 124
rect 566 119 572 120
rect 662 123 669 124
rect 662 119 663 123
rect 668 119 669 123
rect 702 120 703 124
rect 707 120 708 124
rect 799 121 800 125
rect 804 121 805 125
rect 799 120 805 121
rect 838 124 844 125
rect 974 124 980 125
rect 1110 124 1116 125
rect 1974 124 1980 125
rect 3798 124 3804 125
rect 3886 124 3892 125
rect 4022 124 4028 125
rect 4158 124 4164 125
rect 4294 124 4300 125
rect 4462 124 4468 125
rect 4560 124 4562 128
rect 5502 127 5503 131
rect 5507 130 5508 131
rect 5507 128 5642 130
rect 5507 127 5508 128
rect 5502 126 5508 127
rect 5640 126 5642 128
rect 5639 125 5645 126
rect 4654 124 4660 125
rect 4870 124 4876 125
rect 5094 124 5100 125
rect 5326 124 5332 125
rect 838 120 839 124
rect 843 120 844 124
rect 702 119 708 120
rect 838 119 844 120
rect 935 123 941 124
rect 935 119 936 123
rect 940 122 941 123
rect 954 123 960 124
rect 954 122 955 123
rect 940 120 955 122
rect 940 119 941 120
rect 274 118 280 119
rect 386 118 397 119
rect 522 118 533 119
rect 662 118 669 119
rect 935 118 941 119
rect 954 119 955 120
rect 959 119 960 123
rect 974 120 975 124
rect 979 120 980 124
rect 974 119 980 120
rect 1071 123 1077 124
rect 1071 119 1072 123
rect 1076 122 1077 123
rect 1090 123 1096 124
rect 1090 122 1091 123
rect 1076 120 1091 122
rect 1076 119 1077 120
rect 954 118 960 119
rect 1071 118 1077 119
rect 1090 119 1091 120
rect 1095 119 1096 123
rect 1110 120 1111 124
rect 1115 120 1116 124
rect 1110 119 1116 120
rect 1206 123 1213 124
rect 1206 119 1207 123
rect 1212 119 1213 123
rect 1090 118 1096 119
rect 1206 118 1213 119
rect 1934 123 1940 124
rect 1934 119 1935 123
rect 1939 119 1940 123
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 1994 123 2000 124
rect 1994 119 1995 123
rect 1999 119 2000 123
rect 1934 118 1940 119
rect 1994 118 2000 119
rect 2130 123 2136 124
rect 2130 119 2131 123
rect 2135 119 2136 123
rect 2130 118 2136 119
rect 2266 123 2272 124
rect 2266 119 2267 123
rect 2271 119 2272 123
rect 2266 118 2272 119
rect 2402 123 2408 124
rect 2402 119 2403 123
rect 2407 119 2408 123
rect 2402 118 2408 119
rect 2538 123 2544 124
rect 2538 119 2539 123
rect 2543 119 2544 123
rect 2538 118 2544 119
rect 2674 123 2680 124
rect 2674 119 2675 123
rect 2679 119 2680 123
rect 2674 118 2680 119
rect 2810 123 2816 124
rect 2810 119 2811 123
rect 2815 119 2816 123
rect 2810 118 2816 119
rect 2946 123 2952 124
rect 2946 119 2947 123
rect 2951 119 2952 123
rect 2946 118 2952 119
rect 3082 123 3088 124
rect 3082 119 3083 123
rect 3087 119 3088 123
rect 3082 118 3088 119
rect 3218 123 3224 124
rect 3218 119 3219 123
rect 3223 119 3224 123
rect 3218 118 3224 119
rect 3354 123 3360 124
rect 3354 119 3355 123
rect 3359 119 3360 123
rect 3354 118 3360 119
rect 3490 123 3496 124
rect 3490 119 3491 123
rect 3495 119 3496 123
rect 3490 118 3496 119
rect 3626 123 3632 124
rect 3626 119 3627 123
rect 3631 119 3632 123
rect 3798 120 3799 124
rect 3803 120 3804 124
rect 3798 119 3804 120
rect 3838 123 3844 124
rect 3838 119 3839 123
rect 3843 119 3844 123
rect 3886 120 3887 124
rect 3891 120 3892 124
rect 3886 119 3892 120
rect 3983 123 3989 124
rect 3983 119 3984 123
rect 3988 122 3989 123
rect 4002 123 4008 124
rect 4002 122 4003 123
rect 3988 120 4003 122
rect 3988 119 3989 120
rect 3626 118 3632 119
rect 3838 118 3844 119
rect 3983 118 3989 119
rect 4002 119 4003 120
rect 4007 119 4008 123
rect 4022 120 4023 124
rect 4027 120 4028 124
rect 4022 119 4028 120
rect 4114 123 4125 124
rect 4114 119 4115 123
rect 4119 119 4120 123
rect 4124 119 4125 123
rect 4158 120 4159 124
rect 4163 120 4164 124
rect 4158 119 4164 120
rect 4250 123 4261 124
rect 4250 119 4251 123
rect 4255 119 4256 123
rect 4260 119 4261 123
rect 4294 120 4295 124
rect 4299 120 4300 124
rect 4294 119 4300 120
rect 4390 123 4397 124
rect 4390 119 4391 123
rect 4396 119 4397 123
rect 4462 120 4463 124
rect 4467 120 4468 124
rect 4462 119 4468 120
rect 4559 123 4565 124
rect 4559 119 4560 123
rect 4564 119 4565 123
rect 4654 120 4655 124
rect 4659 120 4660 124
rect 4654 119 4660 120
rect 4751 123 4757 124
rect 4751 119 4752 123
rect 4756 122 4757 123
rect 4850 123 4856 124
rect 4850 122 4851 123
rect 4756 120 4851 122
rect 4756 119 4757 120
rect 4002 118 4008 119
rect 4114 118 4125 119
rect 4250 118 4261 119
rect 4390 118 4397 119
rect 4559 118 4565 119
rect 4751 118 4757 119
rect 4850 119 4851 120
rect 4855 119 4856 123
rect 4870 120 4871 124
rect 4875 120 4876 124
rect 4870 119 4876 120
rect 4967 123 4973 124
rect 4967 119 4968 123
rect 4972 122 4973 123
rect 5074 123 5080 124
rect 5074 122 5075 123
rect 4972 120 5075 122
rect 4972 119 4973 120
rect 4850 118 4856 119
rect 4967 118 4973 119
rect 5074 119 5075 120
rect 5079 119 5080 123
rect 5094 120 5095 124
rect 5099 120 5100 124
rect 5094 119 5100 120
rect 5186 123 5197 124
rect 5186 119 5187 123
rect 5191 119 5192 123
rect 5196 119 5197 123
rect 5326 120 5327 124
rect 5331 120 5332 124
rect 5326 119 5332 120
rect 5542 124 5548 125
rect 5542 120 5543 124
rect 5547 120 5548 124
rect 5639 121 5640 125
rect 5644 121 5645 125
rect 5639 120 5645 121
rect 5662 123 5668 124
rect 5542 119 5548 120
rect 5662 119 5663 123
rect 5667 119 5668 123
rect 5074 118 5080 119
rect 5186 118 5197 119
rect 5662 118 5668 119
rect 2022 108 2028 109
rect 2158 108 2164 109
rect 2294 108 2300 109
rect 2430 108 2436 109
rect 2566 108 2572 109
rect 2702 108 2708 109
rect 2838 108 2844 109
rect 2974 108 2980 109
rect 3110 108 3116 109
rect 3246 108 3252 109
rect 3382 108 3388 109
rect 3518 108 3524 109
rect 3654 108 3660 109
rect 1974 107 1980 108
rect 1974 103 1975 107
rect 1979 103 1980 107
rect 2022 104 2023 108
rect 2027 104 2028 108
rect 2022 103 2028 104
rect 2119 107 2125 108
rect 2119 103 2120 107
rect 2124 106 2125 107
rect 2138 107 2144 108
rect 2138 106 2139 107
rect 2124 104 2139 106
rect 2124 103 2125 104
rect 1974 102 1980 103
rect 2119 102 2125 103
rect 2138 103 2139 104
rect 2143 103 2144 107
rect 2158 104 2159 108
rect 2163 104 2164 108
rect 2158 103 2164 104
rect 2255 107 2261 108
rect 2255 103 2256 107
rect 2260 106 2261 107
rect 2274 107 2280 108
rect 2274 106 2275 107
rect 2260 104 2275 106
rect 2260 103 2261 104
rect 2138 102 2144 103
rect 2255 102 2261 103
rect 2274 103 2275 104
rect 2279 103 2280 107
rect 2294 104 2295 108
rect 2299 104 2300 108
rect 2294 103 2300 104
rect 2391 107 2397 108
rect 2391 103 2392 107
rect 2396 106 2397 107
rect 2410 107 2416 108
rect 2410 106 2411 107
rect 2396 104 2411 106
rect 2396 103 2397 104
rect 2274 102 2280 103
rect 2391 102 2397 103
rect 2410 103 2411 104
rect 2415 103 2416 107
rect 2430 104 2431 108
rect 2435 104 2436 108
rect 2430 103 2436 104
rect 2527 107 2533 108
rect 2527 103 2528 107
rect 2532 106 2533 107
rect 2546 107 2552 108
rect 2546 106 2547 107
rect 2532 104 2547 106
rect 2532 103 2533 104
rect 2410 102 2416 103
rect 2527 102 2533 103
rect 2546 103 2547 104
rect 2551 103 2552 107
rect 2566 104 2567 108
rect 2571 104 2572 108
rect 2566 103 2572 104
rect 2663 107 2669 108
rect 2663 103 2664 107
rect 2668 106 2669 107
rect 2682 107 2688 108
rect 2682 106 2683 107
rect 2668 104 2683 106
rect 2668 103 2669 104
rect 2546 102 2552 103
rect 2663 102 2669 103
rect 2682 103 2683 104
rect 2687 103 2688 107
rect 2702 104 2703 108
rect 2707 104 2708 108
rect 2702 103 2708 104
rect 2799 107 2805 108
rect 2799 103 2800 107
rect 2804 106 2805 107
rect 2818 107 2824 108
rect 2818 106 2819 107
rect 2804 104 2819 106
rect 2804 103 2805 104
rect 2682 102 2688 103
rect 2799 102 2805 103
rect 2818 103 2819 104
rect 2823 103 2824 107
rect 2838 104 2839 108
rect 2843 104 2844 108
rect 2838 103 2844 104
rect 2935 107 2941 108
rect 2935 103 2936 107
rect 2940 106 2941 107
rect 2954 107 2960 108
rect 2954 106 2955 107
rect 2940 104 2955 106
rect 2940 103 2941 104
rect 2818 102 2824 103
rect 2935 102 2941 103
rect 2954 103 2955 104
rect 2959 103 2960 107
rect 2974 104 2975 108
rect 2979 104 2980 108
rect 2974 103 2980 104
rect 3071 107 3077 108
rect 3071 103 3072 107
rect 3076 106 3077 107
rect 3090 107 3096 108
rect 3090 106 3091 107
rect 3076 104 3091 106
rect 3076 103 3077 104
rect 2954 102 2960 103
rect 3071 102 3077 103
rect 3090 103 3091 104
rect 3095 103 3096 107
rect 3110 104 3111 108
rect 3115 104 3116 108
rect 3110 103 3116 104
rect 3207 107 3213 108
rect 3207 103 3208 107
rect 3212 106 3213 107
rect 3226 107 3232 108
rect 3226 106 3227 107
rect 3212 104 3227 106
rect 3212 103 3213 104
rect 3090 102 3096 103
rect 3207 102 3213 103
rect 3226 103 3227 104
rect 3231 103 3232 107
rect 3246 104 3247 108
rect 3251 104 3252 108
rect 3246 103 3252 104
rect 3343 107 3349 108
rect 3343 103 3344 107
rect 3348 106 3349 107
rect 3362 107 3368 108
rect 3362 106 3363 107
rect 3348 104 3363 106
rect 3348 103 3349 104
rect 3226 102 3232 103
rect 3343 102 3349 103
rect 3362 103 3363 104
rect 3367 103 3368 107
rect 3382 104 3383 108
rect 3387 104 3388 108
rect 3382 103 3388 104
rect 3479 107 3485 108
rect 3479 103 3480 107
rect 3484 106 3485 107
rect 3498 107 3504 108
rect 3498 106 3499 107
rect 3484 104 3499 106
rect 3484 103 3485 104
rect 3362 102 3368 103
rect 3479 102 3485 103
rect 3498 103 3499 104
rect 3503 103 3504 107
rect 3518 104 3519 108
rect 3523 104 3524 108
rect 3518 103 3524 104
rect 3615 107 3621 108
rect 3615 103 3616 107
rect 3620 106 3621 107
rect 3634 107 3640 108
rect 3634 106 3635 107
rect 3620 104 3635 106
rect 3620 103 3621 104
rect 3498 102 3504 103
rect 3615 102 3621 103
rect 3634 103 3635 104
rect 3639 103 3640 107
rect 3654 104 3655 108
rect 3659 104 3660 108
rect 3654 103 3660 104
rect 3750 107 3757 108
rect 3750 103 3751 107
rect 3756 103 3757 107
rect 3634 102 3640 103
rect 3750 102 3757 103
rect 3798 107 3804 108
rect 3798 103 3799 107
rect 3803 103 3804 107
rect 3798 102 3804 103
<< m3c >>
rect 1679 5743 1683 5747
rect 379 5735 383 5739
rect 643 5735 647 5739
rect 915 5735 919 5739
rect 1459 5735 1463 5739
rect 1731 5735 1735 5739
rect 111 5688 115 5692
rect 131 5687 135 5691
rect 371 5687 375 5691
rect 635 5687 639 5691
rect 907 5687 911 5691
rect 1179 5687 1183 5691
rect 1451 5687 1455 5691
rect 1723 5687 1727 5691
rect 1935 5688 1939 5692
rect 1975 5689 1979 5693
rect 2511 5688 2515 5692
rect 2663 5688 2667 5692
rect 2755 5687 2759 5691
rect 2815 5688 2819 5692
rect 2907 5687 2911 5691
rect 2975 5688 2979 5692
rect 3071 5687 3072 5691
rect 3072 5687 3075 5691
rect 3143 5688 3147 5692
rect 3239 5687 3240 5691
rect 3240 5687 3243 5691
rect 3319 5688 3323 5692
rect 3415 5687 3416 5691
rect 3416 5687 3419 5691
rect 3495 5688 3499 5692
rect 3591 5687 3592 5691
rect 3592 5687 3595 5691
rect 3799 5689 3803 5693
rect 111 5671 115 5675
rect 159 5672 163 5676
rect 379 5671 383 5675
rect 399 5672 403 5676
rect 643 5671 647 5675
rect 663 5672 667 5676
rect 915 5671 919 5675
rect 935 5672 939 5676
rect 1031 5671 1032 5675
rect 1032 5671 1035 5675
rect 1207 5672 1211 5676
rect 1459 5671 1463 5675
rect 1479 5672 1483 5676
rect 1731 5671 1735 5675
rect 1751 5672 1755 5676
rect 1847 5671 1848 5675
rect 1848 5671 1851 5675
rect 1935 5671 1939 5675
rect 1975 5672 1979 5676
rect 2483 5673 2487 5677
rect 2635 5673 2639 5677
rect 2787 5673 2791 5677
rect 2947 5673 2951 5677
rect 3115 5673 3119 5677
rect 3291 5673 3295 5677
rect 3467 5673 3471 5677
rect 3799 5672 3803 5676
rect 3211 5667 3215 5671
rect 3415 5667 3419 5671
rect 4203 5651 4207 5655
rect 4251 5651 4255 5655
rect 4387 5651 4391 5655
rect 4523 5651 4527 5655
rect 4659 5651 4663 5655
rect 4795 5651 4799 5655
rect 4931 5651 4935 5655
rect 5067 5651 5071 5655
rect 5203 5651 5207 5655
rect 111 5613 115 5617
rect 455 5612 459 5616
rect 647 5612 651 5616
rect 747 5611 748 5615
rect 748 5611 751 5615
rect 855 5612 859 5616
rect 967 5611 971 5615
rect 1087 5612 1091 5616
rect 1179 5611 1183 5615
rect 1327 5612 1331 5616
rect 1583 5612 1587 5616
rect 1679 5611 1680 5615
rect 1680 5611 1683 5615
rect 1815 5612 1819 5616
rect 1927 5611 1931 5615
rect 1935 5613 1939 5617
rect 2907 5615 2911 5619
rect 3071 5615 3075 5619
rect 3211 5623 3215 5627
rect 3239 5615 3243 5619
rect 3775 5623 3779 5627
rect 3591 5615 3595 5619
rect 3839 5604 3843 5608
rect 4107 5603 4111 5607
rect 4243 5603 4247 5607
rect 4379 5603 4383 5607
rect 4515 5603 4519 5607
rect 4651 5603 4655 5607
rect 4787 5603 4791 5607
rect 4923 5603 4927 5607
rect 5059 5603 5063 5607
rect 5195 5603 5199 5607
rect 5663 5604 5667 5608
rect 111 5596 115 5600
rect 427 5597 431 5601
rect 619 5597 623 5601
rect 827 5597 831 5601
rect 1059 5597 1063 5601
rect 1299 5597 1303 5601
rect 1555 5597 1559 5601
rect 1787 5597 1791 5601
rect 1935 5596 1939 5600
rect 1927 5583 1931 5587
rect 2779 5591 2783 5595
rect 2443 5579 2447 5583
rect 2755 5583 2759 5587
rect 3839 5587 3843 5591
rect 4135 5588 4139 5592
rect 4251 5587 4255 5591
rect 4271 5588 4275 5592
rect 4387 5587 4391 5591
rect 4407 5588 4411 5592
rect 4523 5587 4527 5591
rect 4543 5588 4547 5592
rect 4659 5587 4663 5591
rect 4679 5588 4683 5592
rect 4795 5587 4799 5591
rect 4815 5588 4819 5592
rect 4931 5587 4935 5591
rect 4951 5588 4955 5592
rect 5067 5587 5071 5591
rect 5087 5588 5091 5592
rect 5203 5587 5207 5591
rect 5223 5588 5227 5592
rect 5315 5587 5319 5591
rect 5663 5587 5667 5591
rect 3083 5579 3087 5583
rect 3283 5579 3287 5583
rect 3483 5579 3487 5583
rect 3659 5579 3663 5583
rect 4203 5555 4207 5559
rect 4399 5555 4403 5559
rect 747 5547 751 5551
rect 967 5547 971 5551
rect 1319 5547 1323 5551
rect 1847 5547 1851 5551
rect 1031 5539 1035 5543
rect 1975 5532 1979 5536
rect 1995 5531 1999 5535
rect 2203 5531 2207 5535
rect 2435 5531 2439 5535
rect 2659 5531 2663 5535
rect 2867 5531 2871 5535
rect 3075 5531 3079 5535
rect 3275 5531 3279 5535
rect 3475 5531 3479 5535
rect 3651 5531 3655 5535
rect 3799 5532 3803 5536
rect 883 5515 887 5519
rect 931 5511 935 5515
rect 1067 5511 1071 5515
rect 1203 5511 1207 5515
rect 1427 5511 1431 5515
rect 1975 5515 1979 5519
rect 2023 5516 2027 5520
rect 2123 5515 2124 5519
rect 2124 5515 2127 5519
rect 2231 5516 2235 5520
rect 2443 5515 2447 5519
rect 2463 5516 2467 5520
rect 2559 5515 2560 5519
rect 2560 5515 2563 5519
rect 2687 5516 2691 5520
rect 2779 5515 2783 5519
rect 2895 5516 2899 5520
rect 3083 5515 3087 5519
rect 3103 5516 3107 5520
rect 3283 5515 3287 5519
rect 3303 5516 3307 5520
rect 3483 5515 3487 5519
rect 3503 5516 3507 5520
rect 3659 5515 3663 5519
rect 3679 5516 3683 5520
rect 3775 5515 3776 5519
rect 3776 5515 3779 5519
rect 3799 5515 3803 5519
rect 3839 5497 3843 5501
rect 4303 5496 4307 5500
rect 4399 5495 4400 5499
rect 4400 5495 4403 5499
rect 4511 5496 4515 5500
rect 4603 5495 4607 5499
rect 4719 5496 4723 5500
rect 4819 5495 4820 5499
rect 4820 5495 4823 5499
rect 4927 5496 4931 5500
rect 5023 5495 5024 5499
rect 5024 5495 5027 5499
rect 5135 5496 5139 5500
rect 5231 5495 5232 5499
rect 5232 5495 5235 5499
rect 5663 5497 5667 5501
rect 3839 5480 3843 5484
rect 4275 5481 4279 5485
rect 4483 5481 4487 5485
rect 4691 5481 4695 5485
rect 4899 5481 4903 5485
rect 5107 5481 5111 5485
rect 5663 5480 5667 5484
rect 111 5464 115 5468
rect 787 5463 791 5467
rect 923 5463 927 5467
rect 1059 5463 1063 5467
rect 1195 5463 1199 5467
rect 1331 5463 1335 5467
rect 1935 5464 1939 5468
rect 1975 5457 1979 5461
rect 2023 5456 2027 5460
rect 2115 5455 2119 5459
rect 2167 5456 2171 5460
rect 2279 5455 2283 5459
rect 2343 5456 2347 5460
rect 2443 5455 2444 5459
rect 2444 5455 2447 5459
rect 2527 5456 2531 5460
rect 2719 5456 2723 5460
rect 2911 5456 2915 5460
rect 3011 5455 3012 5459
rect 3012 5455 3015 5459
rect 3111 5456 3115 5460
rect 3211 5455 3212 5459
rect 3212 5455 3215 5459
rect 3311 5456 3315 5460
rect 3799 5457 3803 5461
rect 111 5447 115 5451
rect 815 5448 819 5452
rect 931 5447 935 5451
rect 951 5448 955 5452
rect 1067 5447 1071 5451
rect 1087 5448 1091 5452
rect 1203 5447 1207 5451
rect 1223 5448 1227 5452
rect 1319 5447 1320 5451
rect 1320 5447 1323 5451
rect 1359 5448 1363 5452
rect 1455 5448 1456 5451
rect 1456 5448 1459 5451
rect 1455 5447 1459 5448
rect 1935 5447 1939 5451
rect 1975 5440 1979 5444
rect 1995 5441 1999 5445
rect 2139 5441 2143 5445
rect 2315 5441 2319 5445
rect 2499 5441 2503 5445
rect 2691 5441 2695 5445
rect 2883 5441 2887 5445
rect 3083 5441 3087 5445
rect 3283 5441 3287 5445
rect 3799 5440 3803 5444
rect 4559 5431 4563 5435
rect 4603 5423 4607 5427
rect 4819 5431 4823 5435
rect 5315 5431 5319 5435
rect 5231 5423 5235 5427
rect 1251 5415 1255 5419
rect 1455 5415 1459 5419
rect 2123 5391 2127 5395
rect 2279 5391 2283 5395
rect 2559 5391 2563 5395
rect 2979 5391 2983 5395
rect 3011 5391 3015 5395
rect 3211 5391 3215 5395
rect 3787 5375 3791 5379
rect 4723 5379 4727 5383
rect 111 5369 115 5373
rect 903 5368 907 5372
rect 1003 5367 1004 5371
rect 1004 5367 1007 5371
rect 1039 5368 1043 5372
rect 1135 5367 1136 5371
rect 1136 5367 1139 5371
rect 1183 5368 1187 5372
rect 1275 5367 1279 5371
rect 1335 5368 1339 5372
rect 1427 5367 1431 5371
rect 1495 5368 1499 5372
rect 1595 5367 1596 5371
rect 1596 5367 1599 5371
rect 1663 5368 1667 5372
rect 1759 5367 1760 5371
rect 1760 5367 1763 5371
rect 1815 5368 1819 5372
rect 1907 5367 1911 5371
rect 1935 5369 1939 5373
rect 4003 5371 4007 5375
rect 4139 5371 4143 5375
rect 4283 5371 4287 5375
rect 4699 5371 4703 5375
rect 4931 5375 4935 5379
rect 5023 5375 5027 5379
rect 111 5352 115 5356
rect 875 5353 879 5357
rect 1011 5353 1015 5357
rect 1155 5353 1159 5357
rect 1307 5353 1311 5357
rect 1467 5353 1471 5357
rect 1635 5353 1639 5357
rect 1787 5353 1791 5357
rect 1935 5352 1939 5356
rect 2147 5331 2151 5335
rect 2443 5335 2447 5339
rect 3759 5339 3763 5343
rect 2867 5331 2871 5335
rect 3659 5331 3663 5335
rect 3839 5324 3843 5328
rect 3859 5323 3863 5327
rect 3995 5323 3999 5327
rect 4131 5323 4135 5327
rect 4275 5323 4279 5327
rect 4435 5323 4439 5327
rect 4603 5323 4607 5327
rect 4779 5323 4783 5327
rect 4963 5323 4967 5327
rect 5663 5324 5667 5328
rect 2147 5311 2151 5315
rect 2583 5311 2587 5315
rect 4931 5315 4935 5319
rect 1003 5303 1007 5307
rect 1251 5303 1255 5307
rect 1275 5295 1279 5299
rect 1551 5303 1555 5307
rect 1595 5303 1599 5307
rect 2115 5303 2119 5307
rect 3839 5307 3843 5311
rect 3887 5308 3891 5312
rect 4003 5307 4007 5311
rect 4023 5308 4027 5312
rect 4139 5307 4143 5311
rect 4159 5308 4163 5312
rect 4283 5307 4287 5311
rect 4303 5308 4307 5312
rect 4395 5307 4399 5311
rect 4463 5308 4467 5312
rect 4559 5307 4560 5311
rect 4560 5307 4563 5311
rect 4631 5308 4635 5312
rect 4723 5307 4727 5311
rect 4807 5308 4811 5312
rect 4899 5307 4903 5311
rect 4991 5308 4995 5312
rect 5663 5307 5667 5311
rect 1759 5295 1763 5299
rect 1975 5284 1979 5288
rect 2051 5283 2055 5287
rect 2459 5283 2463 5287
rect 2859 5283 2863 5287
rect 3267 5283 3271 5287
rect 3651 5283 3655 5287
rect 3799 5284 3803 5288
rect 863 5271 867 5275
rect 4067 5275 4071 5279
rect 4391 5275 4395 5279
rect 995 5263 999 5267
rect 1135 5267 1139 5271
rect 1251 5263 1255 5267
rect 1543 5267 1547 5271
rect 1779 5267 1783 5271
rect 1907 5267 1911 5271
rect 1975 5267 1979 5271
rect 2079 5268 2083 5272
rect 2199 5267 2203 5271
rect 2487 5268 2491 5272
rect 2583 5267 2584 5271
rect 2584 5267 2587 5271
rect 2887 5268 2891 5272
rect 2979 5267 2983 5271
rect 3295 5268 3299 5272
rect 3659 5267 3663 5271
rect 3679 5268 3683 5272
rect 3787 5267 3791 5271
rect 3799 5267 3803 5271
rect 3839 5245 3843 5249
rect 3999 5244 4003 5248
rect 4099 5243 4100 5247
rect 4100 5243 4103 5247
rect 4199 5244 4203 5248
rect 4299 5243 4300 5247
rect 4300 5243 4303 5247
rect 4399 5244 4403 5248
rect 4491 5243 4495 5247
rect 4607 5244 4611 5248
rect 4699 5243 4703 5247
rect 4823 5244 4827 5248
rect 4923 5243 4924 5247
rect 4924 5243 4927 5247
rect 5039 5244 5043 5248
rect 5135 5243 5136 5247
rect 5136 5243 5139 5247
rect 5663 5245 5667 5249
rect 995 5235 999 5239
rect 1367 5235 1371 5239
rect 3839 5228 3843 5232
rect 3971 5229 3975 5233
rect 4171 5229 4175 5233
rect 4371 5229 4375 5233
rect 4579 5229 4583 5233
rect 4795 5229 4799 5233
rect 5011 5229 5015 5233
rect 5663 5228 5667 5232
rect 111 5216 115 5220
rect 587 5215 591 5219
rect 739 5215 743 5219
rect 899 5215 903 5219
rect 1067 5215 1071 5219
rect 1243 5215 1247 5219
rect 1427 5215 1431 5219
rect 1619 5215 1623 5219
rect 1787 5215 1791 5219
rect 1935 5216 1939 5220
rect 1779 5207 1783 5211
rect 1975 5209 1979 5213
rect 2239 5208 2243 5212
rect 2335 5207 2336 5211
rect 2336 5207 2339 5211
rect 2591 5208 2595 5212
rect 2867 5207 2871 5211
rect 2943 5208 2947 5212
rect 3039 5207 3040 5211
rect 3040 5207 3043 5211
rect 3303 5208 3307 5212
rect 3595 5207 3599 5211
rect 3663 5208 3667 5212
rect 3759 5207 3760 5211
rect 3760 5207 3763 5211
rect 3799 5209 3803 5213
rect 111 5199 115 5203
rect 615 5200 619 5204
rect 711 5199 712 5203
rect 712 5199 715 5203
rect 767 5200 771 5204
rect 863 5199 864 5203
rect 864 5199 867 5203
rect 927 5200 931 5204
rect 1095 5200 1099 5204
rect 1251 5199 1255 5203
rect 1271 5200 1275 5204
rect 1367 5199 1368 5203
rect 1368 5199 1371 5203
rect 1455 5200 1459 5204
rect 1551 5199 1552 5203
rect 1552 5199 1555 5203
rect 1647 5200 1651 5204
rect 1747 5199 1748 5203
rect 1748 5199 1751 5203
rect 1815 5200 1819 5204
rect 1935 5199 1939 5203
rect 1975 5192 1979 5196
rect 2211 5193 2215 5197
rect 2563 5193 2567 5197
rect 2915 5193 2919 5197
rect 3275 5193 3279 5197
rect 3635 5193 3639 5197
rect 3799 5192 3803 5196
rect 4067 5179 4071 5183
rect 4099 5179 4103 5183
rect 4299 5179 4303 5183
rect 4715 5179 4719 5183
rect 4899 5179 4903 5183
rect 4923 5179 4927 5183
rect 2199 5143 2203 5147
rect 2639 5143 2643 5147
rect 3039 5143 3043 5147
rect 3595 5143 3599 5147
rect 3115 5135 3119 5139
rect 111 5129 115 5133
rect 367 5128 371 5132
rect 467 5127 468 5131
rect 468 5127 471 5131
rect 535 5128 539 5132
rect 631 5127 632 5131
rect 632 5127 635 5131
rect 711 5128 715 5132
rect 895 5128 899 5132
rect 1015 5127 1019 5131
rect 1079 5128 1083 5132
rect 1171 5127 1175 5131
rect 1263 5128 1267 5132
rect 1447 5128 1451 5132
rect 1543 5127 1544 5131
rect 1544 5127 1547 5131
rect 1631 5128 1635 5132
rect 1727 5127 1728 5131
rect 1728 5127 1731 5131
rect 1815 5128 1819 5132
rect 1911 5127 1912 5131
rect 1912 5127 1915 5131
rect 1935 5129 1939 5133
rect 4491 5127 4495 5131
rect 4603 5123 4607 5127
rect 5135 5127 5139 5131
rect 111 5112 115 5116
rect 339 5113 343 5117
rect 507 5113 511 5117
rect 683 5113 687 5117
rect 867 5113 871 5117
rect 1051 5113 1055 5117
rect 1235 5113 1239 5117
rect 1419 5113 1423 5117
rect 1603 5113 1607 5117
rect 1787 5113 1791 5117
rect 1935 5112 1939 5116
rect 435 5107 439 5111
rect 2335 5111 2339 5115
rect 1171 5107 1175 5111
rect 2839 5111 2843 5115
rect 3227 5111 3231 5115
rect 3599 5115 3603 5119
rect 3483 5107 3487 5111
rect 3839 5076 3843 5080
rect 4099 5075 4103 5079
rect 4347 5075 4351 5079
rect 4595 5075 4599 5079
rect 4843 5075 4847 5079
rect 5099 5075 5103 5079
rect 5663 5076 5667 5080
rect 435 5063 439 5067
rect 467 5063 471 5067
rect 703 5063 707 5067
rect 1015 5063 1019 5067
rect 1331 5063 1335 5067
rect 1747 5063 1751 5067
rect 1975 5060 1979 5064
rect 2267 5059 2271 5063
rect 1911 5055 1915 5059
rect 2515 5059 2519 5063
rect 2755 5059 2759 5063
rect 2995 5059 2999 5063
rect 3235 5059 3239 5063
rect 3475 5059 3479 5063
rect 3799 5060 3803 5064
rect 3839 5059 3843 5063
rect 4127 5060 4131 5064
rect 4223 5059 4224 5063
rect 4224 5059 4227 5063
rect 4375 5060 4379 5064
rect 4623 5060 4627 5064
rect 4715 5059 4719 5063
rect 4871 5060 4875 5064
rect 4967 5059 4968 5063
rect 4968 5059 4971 5063
rect 5127 5060 5131 5064
rect 5663 5059 5667 5063
rect 3227 5051 3231 5055
rect 1975 5043 1979 5047
rect 2295 5044 2299 5048
rect 2391 5043 2392 5047
rect 2392 5043 2395 5047
rect 2543 5044 2547 5048
rect 2639 5043 2640 5047
rect 2640 5043 2643 5047
rect 2783 5044 2787 5048
rect 3023 5044 3027 5048
rect 3115 5043 3119 5047
rect 3263 5044 3267 5048
rect 3503 5044 3507 5048
rect 3599 5043 3600 5047
rect 3600 5043 3603 5047
rect 3799 5043 3803 5047
rect 227 5023 231 5027
rect 331 5023 335 5027
rect 631 5027 635 5031
rect 819 5023 823 5027
rect 1091 5023 1095 5027
rect 1467 5023 1471 5027
rect 1727 5027 1731 5031
rect 227 4987 231 4991
rect 1207 4987 1211 4991
rect 1467 4991 1471 4995
rect 1783 4991 1787 4995
rect 3839 4985 3843 4989
rect 3983 4984 3987 4988
rect 4083 4983 4084 4987
rect 4084 4983 4087 4987
rect 4223 4984 4227 4988
rect 4319 4983 4320 4987
rect 4320 4983 4323 4987
rect 4447 4984 4451 4988
rect 4603 4983 4607 4987
rect 4655 4984 4659 4988
rect 4751 4983 4752 4987
rect 4752 4983 4755 4987
rect 4855 4984 4859 4988
rect 4951 4983 4952 4987
rect 4952 4983 4955 4987
rect 5039 4984 5043 4988
rect 5151 4983 5155 4987
rect 5215 4984 5219 4988
rect 5315 4983 5316 4987
rect 5316 4983 5319 4987
rect 5391 4984 5395 4988
rect 5543 4984 5547 4988
rect 5635 4983 5639 4987
rect 5663 4985 5667 4989
rect 111 4976 115 4980
rect 131 4975 135 4979
rect 323 4975 327 4979
rect 555 4975 559 4979
rect 811 4975 815 4979
rect 1083 4975 1087 4979
rect 1371 4975 1375 4979
rect 1659 4975 1663 4979
rect 1935 4976 1939 4980
rect 1331 4967 1335 4971
rect 3839 4968 3843 4972
rect 3955 4969 3959 4973
rect 4195 4969 4199 4973
rect 4419 4969 4423 4973
rect 4627 4969 4631 4973
rect 4827 4969 4831 4973
rect 5011 4969 5015 4973
rect 5187 4969 5191 4973
rect 5363 4969 5367 4973
rect 5515 4969 5519 4973
rect 5663 4968 5667 4972
rect 111 4959 115 4963
rect 159 4960 163 4964
rect 331 4959 335 4963
rect 351 4960 355 4964
rect 447 4959 448 4963
rect 448 4959 451 4963
rect 583 4960 587 4964
rect 819 4959 823 4963
rect 839 4960 843 4964
rect 1091 4959 1095 4963
rect 1111 4960 1115 4964
rect 1207 4959 1208 4963
rect 1208 4959 1211 4963
rect 1399 4960 1403 4964
rect 1687 4960 1691 4964
rect 1783 4959 1784 4963
rect 1784 4959 1787 4963
rect 1935 4959 1939 4963
rect 1975 4953 1979 4957
rect 2183 4952 2187 4956
rect 2283 4951 2284 4955
rect 2284 4951 2287 4955
rect 2319 4952 2323 4956
rect 2419 4951 2420 4955
rect 2420 4951 2423 4955
rect 2455 4952 2459 4956
rect 2555 4951 2556 4955
rect 2556 4951 2559 4955
rect 2599 4952 2603 4956
rect 2691 4951 2695 4955
rect 2743 4952 2747 4956
rect 2839 4951 2840 4955
rect 2840 4951 2843 4955
rect 2895 4952 2899 4956
rect 2987 4951 2991 4955
rect 3047 4952 3051 4956
rect 3143 4951 3144 4955
rect 3144 4951 3147 4955
rect 3199 4952 3203 4956
rect 3295 4951 3296 4955
rect 3296 4951 3299 4955
rect 3351 4952 3355 4956
rect 3483 4951 3487 4955
rect 3799 4953 3803 4957
rect 1975 4936 1979 4940
rect 2155 4937 2159 4941
rect 2291 4937 2295 4941
rect 2427 4937 2431 4941
rect 2571 4937 2575 4941
rect 2715 4937 2719 4941
rect 2867 4937 2871 4941
rect 3019 4937 3023 4941
rect 3171 4937 3175 4941
rect 3323 4937 3327 4941
rect 3799 4936 3803 4940
rect 4215 4919 4219 4923
rect 4427 4919 4431 4923
rect 4319 4911 4323 4915
rect 4967 4919 4971 4923
rect 4951 4911 4955 4915
rect 5151 4919 5155 4923
rect 5315 4919 5319 4923
rect 5495 4911 5499 4915
rect 2283 4887 2287 4891
rect 2419 4887 2423 4891
rect 2555 4887 2559 4891
rect 111 4877 115 4881
rect 159 4876 163 4880
rect 251 4875 255 4879
rect 295 4876 299 4880
rect 387 4875 391 4879
rect 431 4876 435 4880
rect 531 4875 532 4879
rect 532 4875 535 4879
rect 567 4876 571 4880
rect 667 4875 668 4879
rect 668 4875 671 4879
rect 703 4876 707 4880
rect 799 4875 800 4879
rect 800 4875 803 4879
rect 1935 4877 1939 4881
rect 2391 4879 2395 4883
rect 2851 4887 2855 4891
rect 3003 4887 3007 4891
rect 3143 4887 3147 4891
rect 3295 4887 3299 4891
rect 2987 4879 2991 4883
rect 111 4860 115 4864
rect 131 4861 135 4865
rect 267 4861 271 4865
rect 403 4861 407 4865
rect 539 4861 543 4865
rect 675 4861 679 4865
rect 1935 4860 1939 4864
rect 4083 4863 4087 4867
rect 4631 4867 4635 4871
rect 4603 4859 4607 4863
rect 4751 4863 4755 4867
rect 4883 4859 4887 4863
rect 5051 4859 5055 4863
rect 5331 4863 5335 4867
rect 5379 4859 5383 4863
rect 5635 4863 5639 4867
rect 2691 4851 2695 4855
rect 2579 4843 2583 4847
rect 2731 4843 2735 4847
rect 3019 4847 3023 4851
rect 3303 4851 3307 4855
rect 3343 4839 3347 4843
rect 387 4803 391 4807
rect 447 4811 451 4815
rect 531 4811 535 4815
rect 667 4811 671 4815
rect 3839 4812 3843 4816
rect 3859 4811 3863 4815
rect 4075 4811 4079 4815
rect 4299 4811 4303 4815
rect 4507 4811 4511 4815
rect 4699 4811 4703 4815
rect 4875 4811 4879 4815
rect 5043 4811 5047 4815
rect 5211 4811 5215 4815
rect 5371 4811 5375 4815
rect 5515 4811 5519 4815
rect 5663 4812 5667 4816
rect 799 4803 803 4807
rect 1975 4796 1979 4800
rect 2427 4795 2431 4799
rect 2571 4795 2575 4799
rect 2723 4795 2727 4799
rect 2875 4795 2879 4799
rect 3027 4795 3031 4799
rect 3179 4795 3183 4799
rect 3799 4796 3803 4800
rect 3839 4795 3843 4799
rect 3887 4796 3891 4800
rect 3983 4795 3984 4799
rect 3984 4795 3987 4799
rect 4103 4796 4107 4800
rect 4327 4796 4331 4800
rect 4427 4795 4428 4799
rect 4428 4795 4431 4799
rect 4535 4796 4539 4800
rect 4631 4795 4632 4799
rect 4632 4795 4635 4799
rect 4727 4796 4731 4800
rect 4883 4795 4887 4799
rect 4903 4796 4907 4800
rect 5051 4795 5055 4799
rect 5071 4796 5075 4800
rect 5167 4795 5168 4799
rect 5168 4795 5171 4799
rect 5239 4796 5243 4800
rect 5379 4795 5383 4799
rect 5399 4796 5403 4800
rect 5495 4795 5496 4799
rect 5496 4795 5499 4799
rect 5543 4796 5547 4800
rect 5639 4795 5640 4799
rect 5640 4795 5643 4799
rect 5663 4795 5667 4799
rect 3019 4787 3023 4791
rect 1975 4779 1979 4783
rect 2455 4780 2459 4784
rect 2579 4779 2583 4783
rect 2599 4780 2603 4784
rect 2731 4779 2735 4783
rect 2751 4780 2755 4784
rect 2851 4779 2852 4783
rect 2852 4779 2855 4783
rect 2903 4780 2907 4784
rect 3003 4779 3004 4783
rect 3004 4779 3007 4783
rect 3055 4780 3059 4784
rect 3207 4780 3211 4784
rect 3303 4779 3304 4783
rect 3304 4779 3307 4783
rect 3799 4779 3803 4783
rect 251 4767 255 4771
rect 275 4763 279 4767
rect 411 4763 415 4767
rect 547 4763 551 4767
rect 683 4763 687 4767
rect 4603 4751 4607 4755
rect 3839 4737 3843 4741
rect 4943 4736 4947 4740
rect 5087 4736 5091 4740
rect 5239 4736 5243 4740
rect 5331 4735 5335 4739
rect 5399 4736 5403 4740
rect 5491 4735 5495 4739
rect 5543 4736 5547 4740
rect 5663 4737 5667 4741
rect 111 4716 115 4720
rect 131 4715 135 4719
rect 267 4715 271 4719
rect 403 4715 407 4719
rect 539 4715 543 4719
rect 675 4715 679 4719
rect 1935 4716 1939 4720
rect 1975 4717 1979 4721
rect 2023 4716 2027 4720
rect 2123 4715 2124 4719
rect 2124 4715 2127 4719
rect 2159 4716 2163 4720
rect 2259 4715 2260 4719
rect 2260 4715 2263 4719
rect 2295 4716 2299 4720
rect 2395 4715 2396 4719
rect 2396 4715 2399 4719
rect 2431 4716 2435 4720
rect 2531 4715 2532 4719
rect 2532 4715 2535 4719
rect 2567 4716 2571 4720
rect 2667 4715 2668 4719
rect 2668 4715 2671 4719
rect 2703 4716 2707 4720
rect 2803 4715 2804 4719
rect 2804 4715 2807 4719
rect 2839 4716 2843 4720
rect 2939 4715 2940 4719
rect 2940 4715 2943 4719
rect 2975 4716 2979 4720
rect 3075 4715 3076 4719
rect 3076 4715 3079 4719
rect 3111 4716 3115 4720
rect 3211 4715 3212 4719
rect 3212 4715 3215 4719
rect 3247 4716 3251 4720
rect 3343 4715 3344 4719
rect 3344 4715 3347 4719
rect 3399 4716 3403 4720
rect 3543 4716 3547 4720
rect 3639 4715 3640 4719
rect 3640 4715 3643 4719
rect 3679 4716 3683 4720
rect 3771 4715 3775 4719
rect 3799 4717 3803 4721
rect 3839 4720 3843 4724
rect 4915 4721 4919 4725
rect 5059 4721 5063 4725
rect 5211 4721 5215 4725
rect 5371 4721 5375 4725
rect 5515 4721 5519 4725
rect 5663 4720 5667 4724
rect 111 4699 115 4703
rect 159 4700 163 4704
rect 275 4699 279 4703
rect 295 4700 299 4704
rect 411 4699 415 4703
rect 431 4700 435 4704
rect 547 4699 551 4703
rect 567 4700 571 4704
rect 683 4699 687 4703
rect 703 4700 707 4704
rect 803 4699 804 4703
rect 804 4699 807 4703
rect 1935 4699 1939 4703
rect 1975 4700 1979 4704
rect 1995 4701 1999 4705
rect 2131 4701 2135 4705
rect 2267 4701 2271 4705
rect 2403 4701 2407 4705
rect 2539 4701 2543 4705
rect 2675 4701 2679 4705
rect 2811 4701 2815 4705
rect 2947 4701 2951 4705
rect 3083 4701 3087 4705
rect 3219 4701 3223 4705
rect 3371 4701 3375 4705
rect 3515 4701 3519 4705
rect 3651 4701 3655 4705
rect 3799 4700 3803 4704
rect 5167 4671 5171 4675
rect 5463 4671 5467 4675
rect 5639 4671 5643 4675
rect 5491 4663 5495 4667
rect 2123 4651 2127 4655
rect 2259 4651 2263 4655
rect 2395 4651 2399 4655
rect 2531 4651 2535 4655
rect 2667 4651 2671 4655
rect 2803 4651 2807 4655
rect 2939 4651 2943 4655
rect 3075 4651 3079 4655
rect 3211 4651 3215 4655
rect 2443 4643 2447 4647
rect 3983 4651 3987 4655
rect 3771 4643 3775 4647
rect 111 4633 115 4637
rect 159 4632 163 4636
rect 295 4632 299 4636
rect 395 4631 396 4635
rect 396 4631 399 4635
rect 431 4632 435 4636
rect 531 4631 532 4635
rect 532 4631 535 4635
rect 567 4632 571 4636
rect 667 4631 668 4635
rect 668 4631 671 4635
rect 703 4632 707 4636
rect 795 4631 799 4635
rect 1935 4633 1939 4637
rect 111 4616 115 4620
rect 131 4617 135 4621
rect 267 4617 271 4621
rect 403 4617 407 4621
rect 539 4617 543 4621
rect 675 4617 679 4621
rect 1935 4616 1939 4620
rect 4867 4611 4871 4615
rect 4963 4611 4967 4615
rect 5155 4611 5159 4615
rect 5347 4611 5351 4615
rect 2567 4587 2571 4591
rect 2639 4587 2643 4591
rect 3067 4587 3071 4591
rect 3467 4587 3471 4591
rect 3639 4587 3643 4591
rect 395 4567 399 4571
rect 531 4567 535 4571
rect 667 4567 671 4571
rect 3839 4564 3843 4568
rect 4771 4563 4775 4567
rect 803 4559 807 4563
rect 4955 4563 4959 4567
rect 5147 4563 5151 4567
rect 5339 4563 5343 4567
rect 5515 4563 5519 4567
rect 5663 4564 5667 4568
rect 3839 4547 3843 4551
rect 4799 4548 4803 4552
rect 4963 4547 4967 4551
rect 4983 4548 4987 4552
rect 5155 4547 5159 4551
rect 5175 4548 5179 4552
rect 5347 4547 5351 4551
rect 5367 4548 5371 4552
rect 5463 4547 5464 4551
rect 5464 4547 5467 4551
rect 5543 4548 5547 4552
rect 5643 4547 5644 4551
rect 5644 4547 5647 4551
rect 5663 4547 5667 4551
rect 1975 4536 1979 4540
rect 2323 4535 2327 4539
rect 795 4531 799 4535
rect 2579 4535 2583 4539
rect 2827 4535 2831 4539
rect 3075 4535 3079 4539
rect 3315 4535 3319 4539
rect 3563 4535 3567 4539
rect 3799 4536 3803 4540
rect 523 4523 527 4527
rect 699 4523 703 4527
rect 883 4523 887 4527
rect 1067 4523 1071 4527
rect 1419 4527 1423 4531
rect 1435 4523 1439 4527
rect 1627 4523 1631 4527
rect 1795 4523 1799 4527
rect 2567 4527 2571 4531
rect 3067 4527 3071 4531
rect 3467 4527 3471 4531
rect 1975 4519 1979 4523
rect 2351 4520 2355 4524
rect 2443 4519 2447 4523
rect 2607 4520 2611 4524
rect 2855 4520 2859 4524
rect 2951 4519 2952 4523
rect 2952 4519 2955 4523
rect 3103 4520 3107 4524
rect 3343 4520 3347 4524
rect 3591 4520 3595 4524
rect 3799 4519 3803 4523
rect 111 4476 115 4480
rect 339 4475 343 4479
rect 515 4475 519 4479
rect 691 4475 695 4479
rect 875 4475 879 4479
rect 1059 4475 1063 4479
rect 1243 4475 1247 4479
rect 1427 4475 1431 4479
rect 1619 4475 1623 4479
rect 1787 4475 1791 4479
rect 1935 4476 1939 4480
rect 3839 4477 3843 4481
rect 4487 4476 4491 4480
rect 4671 4476 4675 4480
rect 4879 4476 4883 4480
rect 4979 4475 4980 4479
rect 4980 4475 4983 4479
rect 5095 4476 5099 4480
rect 5327 4476 5331 4480
rect 5423 4475 5424 4479
rect 5424 4475 5427 4479
rect 5543 4476 5547 4480
rect 5635 4475 5639 4479
rect 5663 4477 5667 4481
rect 111 4459 115 4463
rect 367 4460 371 4464
rect 523 4459 527 4463
rect 543 4460 547 4464
rect 699 4459 703 4463
rect 719 4460 723 4464
rect 883 4459 887 4463
rect 903 4460 907 4464
rect 1067 4459 1071 4463
rect 1087 4460 1091 4464
rect 1179 4459 1183 4463
rect 1271 4460 1275 4464
rect 1435 4459 1439 4463
rect 1455 4460 1459 4464
rect 1627 4459 1631 4463
rect 1647 4460 1651 4464
rect 1795 4459 1799 4463
rect 1815 4460 1819 4464
rect 1911 4459 1912 4463
rect 1912 4459 1915 4463
rect 1935 4459 1939 4463
rect 3839 4460 3843 4464
rect 4459 4461 4463 4465
rect 4643 4461 4647 4465
rect 4851 4461 4855 4465
rect 5067 4461 5071 4465
rect 5299 4461 5303 4465
rect 5515 4461 5519 4465
rect 5663 4460 5667 4464
rect 1975 4453 1979 4457
rect 2543 4452 2547 4456
rect 2639 4451 2640 4455
rect 2640 4451 2643 4455
rect 2783 4452 2787 4456
rect 3015 4452 3019 4456
rect 3127 4451 3131 4455
rect 3247 4452 3251 4456
rect 3347 4451 3348 4455
rect 3348 4451 3351 4455
rect 3471 4452 3475 4456
rect 3571 4451 3572 4455
rect 3572 4451 3575 4455
rect 3679 4452 3683 4456
rect 3771 4451 3775 4455
rect 3799 4453 3803 4457
rect 1975 4436 1979 4440
rect 2515 4437 2519 4441
rect 2755 4437 2759 4441
rect 2987 4437 2991 4441
rect 3219 4437 3223 4441
rect 3443 4437 3447 4441
rect 3651 4437 3655 4441
rect 3799 4436 3803 4440
rect 4551 4411 4555 4415
rect 4979 4411 4983 4415
rect 5643 4411 5647 4415
rect 111 4401 115 4405
rect 567 4400 571 4404
rect 667 4399 668 4403
rect 668 4399 671 4403
rect 711 4400 715 4404
rect 863 4400 867 4404
rect 963 4399 964 4403
rect 964 4399 967 4403
rect 1023 4400 1027 4404
rect 1123 4399 1124 4403
rect 1124 4399 1127 4403
rect 1183 4400 1187 4404
rect 1279 4399 1280 4403
rect 1280 4399 1283 4403
rect 1343 4400 1347 4404
rect 1435 4399 1439 4403
rect 1503 4400 1507 4404
rect 1595 4399 1599 4403
rect 1671 4400 1675 4404
rect 1771 4399 1772 4403
rect 1772 4399 1775 4403
rect 1815 4400 1819 4404
rect 1927 4399 1931 4403
rect 1935 4401 1939 4405
rect 111 4384 115 4388
rect 539 4385 543 4389
rect 683 4385 687 4389
rect 835 4385 839 4389
rect 995 4385 999 4389
rect 1155 4385 1159 4389
rect 1315 4385 1319 4389
rect 1475 4385 1479 4389
rect 1643 4385 1647 4389
rect 2951 4395 2955 4399
rect 1787 4385 1791 4389
rect 1935 4384 1939 4388
rect 3127 4387 3131 4391
rect 3347 4387 3351 4391
rect 3571 4387 3575 4391
rect 2927 4379 2931 4383
rect 3779 4355 3783 4359
rect 1927 4343 1931 4347
rect 3359 4347 3363 4351
rect 4003 4351 4007 4355
rect 4139 4351 4143 4355
rect 4379 4351 4383 4355
rect 4491 4351 4495 4355
rect 4723 4351 4727 4355
rect 4987 4351 4991 4355
rect 5259 4351 5263 4355
rect 5635 4355 5639 4359
rect 667 4335 671 4339
rect 963 4335 967 4339
rect 1123 4335 1127 4339
rect 1175 4327 1179 4331
rect 1543 4335 1547 4339
rect 1595 4327 1599 4331
rect 1771 4335 1775 4339
rect 2387 4339 2391 4343
rect 3243 4339 3247 4343
rect 3771 4343 3775 4347
rect 1911 4327 1915 4331
rect 3839 4304 3843 4308
rect 3859 4303 3863 4307
rect 3995 4303 3999 4307
rect 4131 4303 4135 4307
rect 4283 4303 4287 4307
rect 4483 4303 4487 4307
rect 4715 4303 4719 4307
rect 4979 4303 4983 4307
rect 5251 4303 5255 4307
rect 5515 4303 5519 4307
rect 5663 4304 5667 4308
rect 1047 4295 1051 4299
rect 1975 4292 1979 4296
rect 1207 4287 1211 4291
rect 1995 4291 1999 4295
rect 779 4279 783 4283
rect 1279 4283 1283 4287
rect 1715 4287 1719 4291
rect 2379 4291 2383 4295
rect 2803 4291 2807 4295
rect 3235 4291 3239 4295
rect 3651 4291 3655 4295
rect 3799 4292 3803 4296
rect 3839 4287 3843 4291
rect 3887 4288 3891 4292
rect 4003 4287 4007 4291
rect 4023 4288 4027 4292
rect 4139 4287 4143 4291
rect 4159 4288 4163 4292
rect 4255 4287 4256 4291
rect 4256 4287 4259 4291
rect 4311 4288 4315 4292
rect 4491 4287 4495 4291
rect 4511 4288 4515 4292
rect 4723 4287 4727 4291
rect 4743 4288 4747 4292
rect 4987 4287 4991 4291
rect 5007 4288 5011 4292
rect 5259 4287 5263 4291
rect 5279 4288 5283 4292
rect 5543 4288 5547 4292
rect 5639 4287 5640 4291
rect 5640 4287 5643 4291
rect 5663 4287 5667 4291
rect 1879 4275 1883 4279
rect 1975 4275 1979 4279
rect 2023 4276 2027 4280
rect 2387 4275 2391 4279
rect 2407 4276 2411 4280
rect 2503 4275 2504 4279
rect 2504 4275 2507 4279
rect 2831 4276 2835 4280
rect 2927 4275 2928 4279
rect 2928 4275 2931 4279
rect 3263 4276 3267 4280
rect 3359 4275 3360 4279
rect 3360 4275 3363 4279
rect 3679 4276 3683 4280
rect 3779 4275 3780 4279
rect 3780 4275 3783 4279
rect 3799 4275 3803 4279
rect 4551 4275 4555 4279
rect 111 4232 115 4236
rect 627 4231 631 4235
rect 771 4231 775 4235
rect 923 4231 927 4235
rect 1083 4231 1087 4235
rect 1251 4231 1255 4235
rect 1419 4231 1423 4235
rect 1595 4231 1599 4235
rect 1935 4232 1939 4236
rect 3839 4229 3843 4233
rect 3887 4228 3891 4232
rect 3987 4227 3988 4231
rect 3988 4227 3991 4231
rect 4023 4228 4027 4232
rect 4123 4227 4124 4231
rect 4124 4227 4127 4231
rect 4159 4228 4163 4232
rect 4303 4228 4307 4232
rect 4447 4227 4451 4231
rect 4503 4228 4507 4232
rect 4735 4228 4739 4232
rect 4999 4228 5003 4232
rect 5099 4227 5100 4231
rect 5100 4227 5103 4231
rect 5271 4228 5275 4232
rect 5367 4227 5368 4231
rect 5368 4227 5371 4231
rect 5543 4228 5547 4232
rect 5663 4229 5667 4233
rect 111 4215 115 4219
rect 655 4216 659 4220
rect 779 4215 783 4219
rect 799 4216 803 4220
rect 895 4215 896 4219
rect 896 4215 899 4219
rect 951 4216 955 4220
rect 1047 4215 1048 4219
rect 1048 4215 1051 4219
rect 1111 4216 1115 4220
rect 1207 4215 1208 4219
rect 1208 4215 1211 4219
rect 1279 4216 1283 4220
rect 1447 4216 1451 4220
rect 1543 4215 1544 4219
rect 1544 4215 1547 4219
rect 1623 4216 1627 4220
rect 1715 4215 1719 4219
rect 1935 4215 1939 4219
rect 3839 4212 3843 4216
rect 3859 4213 3863 4217
rect 3995 4213 3999 4217
rect 4131 4213 4135 4217
rect 4275 4213 4279 4217
rect 4475 4213 4479 4217
rect 4707 4213 4711 4217
rect 4971 4213 4975 4217
rect 5243 4213 5247 4217
rect 5515 4213 5519 4217
rect 5663 4212 5667 4216
rect 1975 4189 1979 4193
rect 2023 4188 2027 4192
rect 2123 4187 2124 4191
rect 2124 4187 2127 4191
rect 2191 4188 2195 4192
rect 2287 4187 2288 4191
rect 2288 4187 2291 4191
rect 2383 4188 2387 4192
rect 2479 4187 2480 4191
rect 2480 4187 2483 4191
rect 2583 4188 2587 4192
rect 2683 4187 2684 4191
rect 2684 4187 2687 4191
rect 2783 4188 2787 4192
rect 2883 4187 2884 4191
rect 2884 4187 2887 4191
rect 2983 4188 2987 4192
rect 3243 4187 3247 4191
rect 3799 4189 3803 4193
rect 1975 4172 1979 4176
rect 1995 4173 1999 4177
rect 2163 4173 2167 4177
rect 2355 4173 2359 4177
rect 2555 4173 2559 4177
rect 2755 4173 2759 4177
rect 2955 4173 2959 4177
rect 3799 4172 3803 4176
rect 3987 4163 3991 4167
rect 4123 4163 4127 4167
rect 4447 4163 4451 4167
rect 5099 4163 5103 4167
rect 5639 4163 5643 4167
rect 111 4153 115 4157
rect 519 4152 523 4156
rect 703 4152 707 4156
rect 803 4151 804 4155
rect 804 4151 807 4155
rect 895 4152 899 4156
rect 995 4151 996 4155
rect 996 4151 999 4155
rect 1103 4152 1107 4156
rect 1203 4151 1204 4155
rect 1204 4151 1207 4155
rect 1327 4152 1331 4156
rect 1419 4151 1423 4155
rect 1551 4152 1555 4156
rect 1651 4151 1652 4155
rect 1652 4151 1655 4155
rect 1783 4152 1787 4156
rect 1879 4151 1880 4155
rect 1880 4151 1883 4155
rect 1935 4153 1939 4157
rect 4255 4155 4259 4159
rect 111 4136 115 4140
rect 491 4137 495 4141
rect 675 4137 679 4141
rect 867 4137 871 4141
rect 1075 4137 1079 4141
rect 1299 4137 1303 4141
rect 1523 4137 1527 4141
rect 1755 4137 1759 4141
rect 1935 4136 1939 4140
rect 587 4123 591 4127
rect 1419 4123 1423 4127
rect 2123 4123 2127 4127
rect 2503 4123 2507 4127
rect 2567 4123 2571 4127
rect 2683 4123 2687 4127
rect 2883 4123 2887 4127
rect 2479 4115 2483 4119
rect 587 4087 591 4091
rect 887 4087 891 4091
rect 995 4087 999 4091
rect 1203 4087 1207 4091
rect 1615 4087 1619 4091
rect 1651 4087 1655 4091
rect 2287 4091 2291 4095
rect 2539 4087 2543 4091
rect 2747 4091 2751 4095
rect 3079 4095 3083 4099
rect 5091 4099 5095 4103
rect 5231 4095 5235 4099
rect 3139 4087 3143 4091
rect 4707 4087 4711 4091
rect 4843 4087 4847 4091
rect 5203 4087 5207 4091
rect 5339 4087 5343 4091
rect 5423 4091 5427 4095
rect 463 4059 467 4063
rect 795 4055 799 4059
rect 803 4055 807 4059
rect 1187 4051 1191 4055
rect 1587 4051 1591 4055
rect 1907 4055 1911 4059
rect 2539 4059 2543 4063
rect 2739 4059 2743 4063
rect 5203 4059 5207 4063
rect 5367 4059 5371 4063
rect 5339 4051 5343 4055
rect 5499 4051 5503 4055
rect 1975 4040 1979 4044
rect 2075 4039 2079 4043
rect 2259 4039 2263 4043
rect 2443 4039 2447 4043
rect 2619 4039 2623 4043
rect 2787 4039 2791 4043
rect 2955 4039 2959 4043
rect 3131 4039 3135 4043
rect 3799 4040 3803 4044
rect 3839 4040 3843 4044
rect 4563 4039 4567 4043
rect 4699 4039 4703 4043
rect 4835 4039 4839 4043
rect 4971 4039 4975 4043
rect 5107 4039 5111 4043
rect 5243 4039 5247 4043
rect 5379 4039 5383 4043
rect 5515 4039 5519 4043
rect 5663 4040 5667 4044
rect 1587 4031 1591 4035
rect 1915 4031 1919 4035
rect 2747 4031 2751 4035
rect 1975 4023 1979 4027
rect 2103 4024 2107 4028
rect 2195 4023 2199 4027
rect 2287 4024 2291 4028
rect 2471 4024 2475 4028
rect 2567 4023 2568 4027
rect 2568 4023 2571 4027
rect 2647 4024 2651 4028
rect 2743 4023 2744 4027
rect 2744 4023 2747 4027
rect 2815 4024 2819 4028
rect 2983 4024 2987 4028
rect 3079 4023 3080 4027
rect 3080 4023 3083 4027
rect 3159 4024 3163 4028
rect 3799 4023 3803 4027
rect 3839 4023 3843 4027
rect 4591 4024 4595 4028
rect 4707 4023 4711 4027
rect 4727 4024 4731 4028
rect 4843 4023 4847 4027
rect 4863 4024 4867 4028
rect 4959 4023 4960 4027
rect 4960 4023 4963 4027
rect 4999 4024 5003 4028
rect 5091 4023 5095 4027
rect 5135 4024 5139 4028
rect 5231 4023 5232 4027
rect 5232 4023 5235 4027
rect 5271 4024 5275 4028
rect 5367 4023 5368 4027
rect 5368 4023 5371 4027
rect 5407 4024 5411 4028
rect 5499 4023 5503 4027
rect 5543 4024 5547 4028
rect 5639 4023 5640 4027
rect 5640 4023 5643 4027
rect 5663 4023 5667 4027
rect 111 4004 115 4008
rect 131 4003 135 4007
rect 339 4003 343 4007
rect 595 4003 599 4007
rect 875 4003 879 4007
rect 1179 4003 1183 4007
rect 1491 4003 1495 4007
rect 1787 4003 1791 4007
rect 1935 4004 1939 4008
rect 795 3995 799 3999
rect 111 3987 115 3991
rect 159 3988 163 3992
rect 255 3987 256 3991
rect 256 3987 259 3991
rect 367 3988 371 3992
rect 463 3987 464 3991
rect 464 3987 467 3991
rect 623 3988 627 3992
rect 903 3988 907 3992
rect 1187 3987 1191 3991
rect 1207 3988 1211 3992
rect 1519 3988 1523 3992
rect 1615 3987 1616 3991
rect 1616 3987 1619 3991
rect 1815 3988 1819 3992
rect 1915 3987 1916 3991
rect 1916 3987 1919 3991
rect 1935 3987 1939 3991
rect 1975 3957 1979 3961
rect 2127 3956 2131 3960
rect 2311 3956 2315 3960
rect 2487 3956 2491 3960
rect 2579 3955 2583 3959
rect 2663 3956 2667 3960
rect 2831 3956 2835 3960
rect 2927 3955 2928 3959
rect 2928 3955 2931 3959
rect 2999 3956 3003 3960
rect 3139 3955 3143 3959
rect 3175 3956 3179 3960
rect 3267 3955 3271 3959
rect 3351 3956 3355 3960
rect 3447 3955 3448 3959
rect 3448 3955 3451 3959
rect 3799 3957 3803 3961
rect 363 3939 367 3943
rect 1975 3940 1979 3944
rect 2099 3941 2103 3945
rect 2283 3941 2287 3945
rect 2459 3941 2463 3945
rect 2635 3941 2639 3945
rect 2803 3941 2807 3945
rect 2971 3941 2975 3945
rect 3147 3941 3151 3945
rect 3839 3945 3843 3949
rect 3323 3941 3327 3945
rect 4359 3944 4363 3948
rect 3799 3940 3803 3944
rect 4471 3943 4475 3947
rect 4543 3944 4547 3948
rect 4643 3943 4644 3947
rect 4644 3943 4647 3947
rect 4735 3944 4739 3948
rect 4827 3943 4831 3947
rect 4927 3944 4931 3948
rect 5023 3943 5024 3947
rect 5024 3943 5027 3947
rect 5127 3944 5131 3948
rect 5327 3944 5331 3948
rect 5423 3943 5424 3947
rect 5424 3943 5427 3947
rect 5527 3944 5531 3948
rect 5619 3943 5623 3947
rect 5663 3945 5667 3949
rect 111 3925 115 3929
rect 159 3924 163 3928
rect 275 3923 279 3927
rect 343 3924 347 3928
rect 439 3923 440 3927
rect 440 3923 443 3927
rect 567 3924 571 3928
rect 695 3923 699 3927
rect 807 3924 811 3928
rect 943 3923 947 3927
rect 1055 3924 1059 3928
rect 1311 3924 1315 3928
rect 1575 3924 1579 3928
rect 1815 3924 1819 3928
rect 1907 3923 1911 3927
rect 1935 3925 1939 3929
rect 3839 3928 3843 3932
rect 4331 3929 4335 3933
rect 4515 3929 4519 3933
rect 4707 3929 4711 3933
rect 4899 3929 4903 3933
rect 5099 3929 5103 3933
rect 5299 3929 5303 3933
rect 5499 3929 5503 3933
rect 5663 3928 5667 3932
rect 2731 3919 2735 3923
rect 3267 3919 3271 3923
rect 111 3908 115 3912
rect 131 3909 135 3913
rect 315 3909 319 3913
rect 539 3909 543 3913
rect 779 3909 783 3913
rect 1027 3909 1031 3913
rect 1283 3909 1287 3913
rect 1547 3909 1551 3913
rect 1787 3909 1791 3913
rect 1935 3908 1939 3912
rect 4427 3911 4431 3915
rect 4827 3911 4831 3915
rect 2195 3891 2199 3895
rect 2731 3891 2735 3895
rect 2927 3891 2931 3895
rect 3283 3891 3287 3895
rect 3447 3883 3451 3887
rect 4427 3879 4431 3883
rect 4471 3879 4475 3883
rect 4959 3879 4963 3883
rect 5035 3879 5039 3883
rect 5639 3879 5643 3883
rect 5023 3871 5027 3875
rect 255 3859 259 3863
rect 275 3859 279 3863
rect 439 3859 443 3863
rect 695 3859 699 3863
rect 943 3859 947 3863
rect 1379 3859 1383 3863
rect 2579 3859 2583 3863
rect 2531 3847 2535 3851
rect 2939 3851 2943 3855
rect 2955 3847 2959 3851
rect 3163 3847 3167 3851
rect 3391 3851 3395 3855
rect 3571 3847 3575 3851
rect 4475 3839 4479 3843
rect 4635 3839 4639 3843
rect 4643 3839 4647 3843
rect 5099 3839 5103 3843
rect 5447 3843 5451 3847
rect 5619 3839 5623 3843
rect 363 3819 367 3823
rect 483 3815 487 3819
rect 715 3815 719 3819
rect 971 3815 975 3819
rect 1243 3815 1247 3819
rect 1611 3815 1615 3819
rect 1855 3819 1859 3823
rect 1975 3800 1979 3804
rect 2291 3799 2295 3803
rect 2523 3799 2527 3803
rect 2739 3799 2743 3803
rect 2947 3799 2951 3803
rect 3155 3799 3159 3803
rect 3355 3799 3359 3803
rect 3563 3799 3567 3803
rect 3799 3800 3803 3804
rect 1611 3791 1615 3795
rect 1911 3791 1915 3795
rect 2939 3791 2943 3795
rect 1975 3783 1979 3787
rect 2319 3784 2323 3788
rect 2531 3783 2535 3787
rect 2551 3784 2555 3788
rect 2647 3783 2648 3787
rect 2648 3783 2651 3787
rect 2767 3784 2771 3788
rect 2955 3783 2959 3787
rect 2975 3784 2979 3788
rect 3163 3783 3167 3787
rect 3183 3784 3187 3788
rect 3283 3783 3284 3787
rect 3284 3783 3287 3787
rect 3383 3784 3387 3788
rect 3571 3783 3575 3787
rect 3591 3784 3595 3788
rect 3839 3788 3843 3792
rect 4051 3787 4055 3791
rect 3799 3783 3803 3787
rect 4267 3787 4271 3791
rect 4483 3787 4487 3791
rect 4699 3787 4703 3791
rect 4907 3787 4911 3791
rect 5115 3787 5119 3791
rect 5323 3787 5327 3791
rect 5515 3787 5519 3791
rect 5663 3788 5667 3792
rect 4475 3779 4479 3783
rect 4635 3779 4639 3783
rect 5099 3779 5103 3783
rect 111 3768 115 3772
rect 267 3767 271 3771
rect 475 3767 479 3771
rect 707 3767 711 3771
rect 963 3767 967 3771
rect 1235 3767 1239 3771
rect 1515 3767 1519 3771
rect 1787 3767 1791 3771
rect 1935 3768 1939 3772
rect 3839 3771 3843 3775
rect 4079 3772 4083 3776
rect 4171 3771 4175 3775
rect 4295 3772 4299 3776
rect 4511 3772 4515 3776
rect 4727 3772 4731 3776
rect 4935 3772 4939 3776
rect 5035 3771 5036 3775
rect 5036 3771 5039 3775
rect 5143 3772 5147 3776
rect 5351 3772 5355 3776
rect 5447 3771 5448 3775
rect 5448 3771 5451 3775
rect 5543 3772 5547 3776
rect 5663 3771 5667 3775
rect 1379 3759 1383 3763
rect 111 3751 115 3755
rect 295 3752 299 3756
rect 483 3751 487 3755
rect 503 3752 507 3756
rect 715 3751 719 3755
rect 735 3752 739 3756
rect 971 3751 975 3755
rect 991 3752 995 3756
rect 1243 3751 1247 3755
rect 1263 3752 1267 3756
rect 1543 3752 1547 3756
rect 1815 3752 1819 3756
rect 1911 3751 1912 3755
rect 1912 3751 1915 3755
rect 1935 3751 1939 3755
rect 699 3735 703 3739
rect 1975 3721 1979 3725
rect 2407 3720 2411 3724
rect 2503 3719 2504 3723
rect 2504 3719 2507 3723
rect 2647 3720 2651 3724
rect 2743 3719 2744 3723
rect 2744 3719 2747 3723
rect 2871 3720 2875 3724
rect 2971 3719 2972 3723
rect 2972 3719 2975 3723
rect 3087 3720 3091 3724
rect 3187 3719 3188 3723
rect 3188 3719 3191 3723
rect 3295 3720 3299 3724
rect 3391 3719 3392 3723
rect 3392 3719 3395 3723
rect 3495 3720 3499 3724
rect 3591 3719 3592 3723
rect 3592 3719 3595 3723
rect 3679 3720 3683 3724
rect 3771 3719 3775 3723
rect 3799 3721 3803 3725
rect 1975 3704 1979 3708
rect 2379 3705 2383 3709
rect 2619 3705 2623 3709
rect 2843 3705 2847 3709
rect 3059 3705 3063 3709
rect 3267 3705 3271 3709
rect 3467 3705 3471 3709
rect 3651 3705 3655 3709
rect 3799 3704 3803 3708
rect 111 3689 115 3693
rect 631 3688 635 3692
rect 731 3687 732 3691
rect 732 3687 735 3691
rect 775 3688 779 3692
rect 927 3688 931 3692
rect 1027 3687 1028 3691
rect 1028 3687 1031 3691
rect 1087 3688 1091 3692
rect 1187 3687 1188 3691
rect 1188 3687 1191 3691
rect 1255 3688 1259 3692
rect 1347 3687 1351 3691
rect 1423 3688 1427 3692
rect 1523 3687 1524 3691
rect 1524 3687 1527 3691
rect 1591 3688 1595 3692
rect 1691 3687 1692 3691
rect 1692 3687 1695 3691
rect 1759 3688 1763 3692
rect 1855 3687 1856 3691
rect 1856 3687 1859 3691
rect 1935 3689 1939 3693
rect 2939 3683 2943 3687
rect 3591 3683 3595 3687
rect 3839 3685 3843 3689
rect 3887 3684 3891 3688
rect 3983 3683 3984 3687
rect 3984 3683 3987 3687
rect 4055 3684 4059 3688
rect 4183 3683 4187 3687
rect 4247 3684 4251 3688
rect 4439 3684 4443 3688
rect 4567 3683 4571 3687
rect 4631 3684 4635 3688
rect 4723 3683 4727 3687
rect 5663 3685 5667 3689
rect 111 3672 115 3676
rect 603 3673 607 3677
rect 747 3673 751 3677
rect 899 3673 903 3677
rect 1059 3673 1063 3677
rect 1227 3673 1231 3677
rect 1395 3673 1399 3677
rect 1563 3673 1567 3677
rect 1731 3673 1735 3677
rect 1935 3672 1939 3676
rect 3839 3668 3843 3672
rect 3859 3669 3863 3673
rect 4027 3669 4031 3673
rect 4219 3669 4223 3673
rect 4411 3669 4415 3673
rect 4603 3669 4607 3673
rect 5663 3668 5667 3672
rect 2639 3655 2643 3659
rect 2939 3655 2943 3659
rect 2971 3655 2975 3659
rect 3187 3655 3191 3659
rect 2743 3647 2747 3651
rect 3983 3655 3987 3659
rect 3771 3647 3775 3651
rect 699 3623 703 3627
rect 731 3623 735 3627
rect 1027 3623 1031 3627
rect 1187 3623 1191 3627
rect 1523 3623 1527 3627
rect 1691 3623 1695 3627
rect 1851 3615 1855 3619
rect 2503 3615 2507 3619
rect 3955 3619 3959 3623
rect 4171 3619 4175 3623
rect 4183 3619 4187 3623
rect 4567 3619 4571 3623
rect 2555 3611 2559 3615
rect 2691 3611 2695 3615
rect 1347 3587 1351 3591
rect 1371 3587 1375 3591
rect 3779 3587 3783 3591
rect 4723 3595 4727 3599
rect 4003 3583 4007 3587
rect 4139 3583 4143 3587
rect 4275 3583 4279 3587
rect 4411 3583 4415 3587
rect 4683 3583 4687 3587
rect 4819 3583 4823 3587
rect 4955 3583 4959 3587
rect 5091 3583 5095 3587
rect 923 3575 927 3579
rect 1059 3575 1063 3579
rect 1195 3575 1199 3579
rect 1331 3575 1335 3579
rect 1603 3575 1607 3579
rect 1739 3575 1743 3579
rect 1975 3564 1979 3568
rect 2411 3563 2415 3567
rect 2547 3563 2551 3567
rect 2683 3563 2687 3567
rect 3799 3564 3803 3568
rect 1975 3547 1979 3551
rect 2439 3548 2443 3552
rect 2555 3547 2559 3551
rect 2575 3548 2579 3552
rect 2691 3547 2695 3551
rect 2711 3548 2715 3552
rect 2807 3547 2808 3551
rect 2808 3547 2811 3551
rect 3799 3547 3803 3551
rect 3839 3536 3843 3540
rect 3859 3535 3863 3539
rect 3995 3535 3999 3539
rect 4131 3535 4135 3539
rect 4267 3535 4271 3539
rect 4403 3535 4407 3539
rect 4539 3535 4543 3539
rect 4675 3535 4679 3539
rect 4811 3535 4815 3539
rect 4947 3535 4951 3539
rect 5083 3535 5087 3539
rect 5663 3536 5667 3540
rect 111 3528 115 3532
rect 779 3527 783 3531
rect 915 3527 919 3531
rect 1051 3527 1055 3531
rect 1187 3527 1191 3531
rect 1323 3527 1327 3531
rect 1459 3527 1463 3531
rect 1595 3527 1599 3531
rect 1731 3527 1735 3531
rect 1935 3528 1939 3532
rect 3839 3519 3843 3523
rect 3887 3520 3891 3524
rect 4003 3519 4007 3523
rect 4023 3520 4027 3524
rect 4139 3519 4143 3523
rect 4159 3520 4163 3524
rect 4275 3519 4279 3523
rect 4295 3520 4299 3524
rect 4411 3519 4415 3523
rect 4431 3520 4435 3524
rect 4527 3519 4528 3523
rect 4528 3519 4531 3523
rect 4567 3520 4571 3524
rect 4683 3519 4687 3523
rect 4703 3520 4707 3524
rect 4819 3519 4823 3523
rect 4839 3520 4843 3524
rect 4955 3519 4959 3523
rect 4975 3520 4979 3524
rect 5091 3519 5095 3523
rect 5111 3520 5115 3524
rect 5207 3519 5208 3523
rect 5208 3519 5211 3523
rect 5663 3519 5667 3523
rect 111 3511 115 3515
rect 807 3512 811 3516
rect 923 3511 927 3515
rect 943 3512 947 3516
rect 1059 3511 1063 3515
rect 1079 3512 1083 3516
rect 1195 3511 1199 3515
rect 1215 3512 1219 3516
rect 1331 3511 1335 3515
rect 1351 3512 1355 3516
rect 1447 3511 1448 3515
rect 1448 3511 1451 3515
rect 1487 3512 1491 3516
rect 1603 3511 1607 3515
rect 1623 3512 1627 3516
rect 1739 3511 1743 3515
rect 1759 3512 1763 3516
rect 1851 3511 1855 3515
rect 1935 3511 1939 3515
rect 4899 3483 4903 3487
rect 5207 3483 5211 3487
rect 1975 3449 1979 3453
rect 2599 3448 2603 3452
rect 2699 3447 2700 3451
rect 2700 3447 2703 3451
rect 2823 3448 2827 3452
rect 2915 3447 2919 3451
rect 3047 3448 3051 3452
rect 3147 3447 3148 3451
rect 3148 3447 3151 3451
rect 3263 3448 3267 3452
rect 3363 3447 3364 3451
rect 3364 3447 3367 3451
rect 3479 3448 3483 3452
rect 3599 3447 3603 3451
rect 3679 3448 3683 3452
rect 3779 3447 3780 3451
rect 3780 3447 3783 3451
rect 3799 3449 3803 3453
rect 3839 3453 3843 3457
rect 4831 3452 4835 3456
rect 4931 3451 4932 3455
rect 4932 3451 4935 3455
rect 4967 3452 4971 3456
rect 5067 3451 5068 3455
rect 5068 3451 5071 3455
rect 5103 3452 5107 3456
rect 5203 3451 5204 3455
rect 5204 3451 5207 3455
rect 5239 3452 5243 3456
rect 5339 3451 5340 3455
rect 5340 3451 5343 3455
rect 5375 3452 5379 3456
rect 5471 3451 5472 3455
rect 5472 3451 5475 3455
rect 5663 3453 5667 3457
rect 111 3429 115 3433
rect 727 3428 731 3432
rect 827 3427 828 3431
rect 828 3427 831 3431
rect 863 3428 867 3432
rect 963 3427 964 3431
rect 964 3427 967 3431
rect 999 3428 1003 3432
rect 1135 3428 1139 3432
rect 1235 3427 1236 3431
rect 1236 3427 1239 3431
rect 1271 3428 1275 3432
rect 1371 3427 1372 3431
rect 1372 3427 1375 3431
rect 1407 3428 1411 3432
rect 1507 3427 1508 3431
rect 1508 3427 1511 3431
rect 1543 3428 1547 3432
rect 1643 3427 1644 3431
rect 1644 3427 1647 3431
rect 1679 3428 1683 3432
rect 1779 3427 1780 3431
rect 1780 3427 1783 3431
rect 1815 3428 1819 3432
rect 1907 3427 1911 3431
rect 1935 3429 1939 3433
rect 1975 3432 1979 3436
rect 2571 3433 2575 3437
rect 2795 3433 2799 3437
rect 3019 3433 3023 3437
rect 3235 3433 3239 3437
rect 3451 3433 3455 3437
rect 3651 3433 3655 3437
rect 3799 3432 3803 3436
rect 3839 3436 3843 3440
rect 4803 3437 4807 3441
rect 4939 3437 4943 3441
rect 5075 3437 5079 3441
rect 5211 3437 5215 3441
rect 5347 3437 5351 3441
rect 5663 3436 5667 3440
rect 111 3412 115 3416
rect 699 3413 703 3417
rect 835 3413 839 3417
rect 971 3413 975 3417
rect 1107 3413 1111 3417
rect 1243 3413 1247 3417
rect 1379 3413 1383 3417
rect 1515 3413 1519 3417
rect 1651 3413 1655 3417
rect 1787 3413 1791 3417
rect 1935 3412 1939 3416
rect 2807 3383 2811 3387
rect 3115 3383 3119 3387
rect 3147 3383 3151 3387
rect 3363 3383 3367 3387
rect 3599 3383 3603 3387
rect 4899 3387 4903 3391
rect 4931 3387 4935 3391
rect 5067 3387 5071 3391
rect 5203 3387 5207 3391
rect 5339 3387 5343 3391
rect 2915 3375 2919 3379
rect 827 3363 831 3367
rect 963 3363 967 3367
rect 1235 3363 1239 3367
rect 1447 3363 1451 3367
rect 1507 3363 1511 3367
rect 1643 3363 1647 3367
rect 1779 3363 1783 3367
rect 875 3355 879 3359
rect 4263 3359 4267 3363
rect 5303 3359 5307 3363
rect 4147 3351 4151 3355
rect 4523 3351 4527 3355
rect 4699 3351 4703 3355
rect 5471 3355 5475 3359
rect 2699 3343 2703 3347
rect 3071 3343 3075 3347
rect 5419 3347 5423 3351
rect 1159 3335 1163 3339
rect 3091 3339 3095 3343
rect 3275 3339 3279 3343
rect 1019 3327 1023 3331
rect 1463 3331 1467 3335
rect 1907 3331 1911 3335
rect 1131 3323 1135 3327
rect 1435 3323 1439 3327
rect 1659 3323 1663 3327
rect 1795 3323 1799 3327
rect 3839 3304 3843 3308
rect 3859 3303 3863 3307
rect 3115 3299 3119 3303
rect 4139 3303 4143 3307
rect 4427 3303 4431 3307
rect 4691 3303 4695 3307
rect 4939 3303 4943 3307
rect 5179 3303 5183 3307
rect 5427 3303 5431 3307
rect 5663 3304 5667 3308
rect 1975 3292 1979 3296
rect 2531 3291 2535 3295
rect 2715 3291 2719 3295
rect 2899 3291 2903 3295
rect 3083 3291 3087 3295
rect 3267 3291 3271 3295
rect 3799 3292 3803 3296
rect 5419 3295 5423 3299
rect 3839 3287 3843 3291
rect 3887 3288 3891 3292
rect 4167 3288 4171 3292
rect 4263 3287 4264 3291
rect 4264 3287 4267 3291
rect 4455 3288 4459 3292
rect 4699 3287 4703 3291
rect 4719 3288 4723 3292
rect 4819 3287 4820 3291
rect 4820 3287 4823 3291
rect 4967 3288 4971 3292
rect 5059 3287 5063 3291
rect 5207 3288 5211 3292
rect 5303 3287 5304 3291
rect 5304 3287 5307 3291
rect 5455 3288 5459 3292
rect 5663 3287 5667 3291
rect 111 3276 115 3280
rect 755 3275 759 3279
rect 891 3275 895 3279
rect 1035 3275 1039 3279
rect 1187 3275 1191 3279
rect 1339 3275 1343 3279
rect 1491 3275 1495 3279
rect 1651 3275 1655 3279
rect 1787 3275 1791 3279
rect 1935 3276 1939 3280
rect 1975 3275 1979 3279
rect 2559 3276 2563 3280
rect 2655 3275 2656 3279
rect 2656 3275 2659 3279
rect 2743 3276 2747 3280
rect 2927 3276 2931 3280
rect 3091 3275 3095 3279
rect 3111 3276 3115 3280
rect 3275 3275 3279 3279
rect 3295 3276 3299 3280
rect 3403 3275 3407 3279
rect 3799 3275 3803 3279
rect 1019 3267 1023 3271
rect 111 3259 115 3263
rect 783 3260 787 3264
rect 875 3259 879 3263
rect 919 3260 923 3264
rect 1011 3259 1015 3263
rect 1063 3260 1067 3264
rect 1159 3259 1160 3263
rect 1160 3259 1163 3263
rect 1215 3260 1219 3264
rect 1367 3260 1371 3264
rect 1463 3259 1464 3263
rect 1464 3259 1467 3263
rect 1519 3260 1523 3264
rect 1659 3259 1663 3263
rect 1679 3260 1683 3264
rect 1795 3259 1799 3263
rect 1815 3260 1819 3264
rect 1911 3259 1912 3263
rect 1912 3259 1915 3263
rect 1935 3259 1939 3263
rect 1131 3215 1135 3219
rect 111 3201 115 3205
rect 1435 3215 1439 3219
rect 1975 3217 1979 3221
rect 2023 3216 2027 3220
rect 2143 3215 2147 3219
rect 2255 3216 2259 3220
rect 2347 3215 2351 3219
rect 2503 3216 2507 3220
rect 2595 3215 2599 3219
rect 2743 3216 2747 3220
rect 2855 3215 2859 3219
rect 2975 3216 2979 3220
rect 3071 3215 3072 3219
rect 3072 3215 3075 3219
rect 3207 3216 3211 3220
rect 3299 3215 3303 3219
rect 3447 3216 3451 3220
rect 3543 3215 3544 3219
rect 3544 3215 3547 3219
rect 3799 3217 3803 3221
rect 391 3200 395 3204
rect 491 3199 492 3203
rect 492 3199 495 3203
rect 647 3200 651 3204
rect 743 3199 744 3203
rect 744 3199 747 3203
rect 927 3200 931 3204
rect 1019 3199 1023 3203
rect 1223 3200 1227 3204
rect 1527 3200 1531 3204
rect 1815 3200 1819 3204
rect 1927 3199 1931 3203
rect 1935 3201 1939 3205
rect 1975 3200 1979 3204
rect 1995 3201 1999 3205
rect 2227 3201 2231 3205
rect 2475 3201 2479 3205
rect 2715 3201 2719 3205
rect 2947 3201 2951 3205
rect 3179 3201 3183 3205
rect 3839 3205 3843 3209
rect 3419 3201 3423 3205
rect 3911 3204 3915 3208
rect 3799 3200 3803 3204
rect 4147 3203 4151 3207
rect 4183 3204 4187 3208
rect 4439 3204 4443 3208
rect 4535 3203 4536 3207
rect 4536 3203 4539 3207
rect 4687 3204 4691 3208
rect 4779 3203 4783 3207
rect 4935 3204 4939 3208
rect 5031 3203 5032 3207
rect 5032 3203 5035 3207
rect 5191 3204 5195 3208
rect 5287 3203 5288 3207
rect 5288 3203 5291 3207
rect 5663 3205 5667 3209
rect 111 3184 115 3188
rect 363 3185 367 3189
rect 619 3185 623 3189
rect 899 3185 903 3189
rect 1195 3185 1199 3189
rect 1499 3185 1503 3189
rect 1787 3185 1791 3189
rect 1935 3184 1939 3188
rect 3839 3188 3843 3192
rect 3883 3189 3887 3193
rect 4155 3189 4159 3193
rect 4411 3189 4415 3193
rect 4659 3189 4663 3193
rect 4907 3189 4911 3193
rect 5163 3189 5167 3193
rect 5663 3188 5667 3192
rect 1927 3151 1931 3155
rect 2143 3151 2147 3155
rect 2655 3151 2659 3155
rect 2855 3151 2859 3155
rect 2899 3143 2903 3147
rect 3403 3151 3407 3155
rect 3543 3143 3547 3147
rect 743 3127 747 3131
rect 1011 3135 1015 3139
rect 1027 3135 1031 3139
rect 1575 3135 1579 3139
rect 1911 3135 1915 3139
rect 4051 3139 4055 3143
rect 1019 3127 1023 3131
rect 4779 3131 4783 3135
rect 4819 3139 4823 3143
rect 5031 3139 5035 3143
rect 5287 3131 5291 3135
rect 2595 3119 2599 3123
rect 2875 3115 2879 3119
rect 3299 3119 3303 3123
rect 3379 3115 3383 3119
rect 3659 3115 3663 3119
rect 4095 3103 4099 3107
rect 431 3095 435 3099
rect 4227 3099 4231 3103
rect 4339 3099 4343 3103
rect 4535 3103 4539 3107
rect 4723 3099 4727 3103
rect 4923 3099 4927 3103
rect 491 3091 495 3095
rect 499 3083 503 3087
rect 803 3087 807 3091
rect 907 3087 911 3091
rect 1267 3091 1271 3095
rect 1283 3087 1287 3091
rect 1459 3087 1463 3091
rect 2347 3091 2351 3095
rect 2875 3075 2879 3079
rect 3215 3075 3219 3079
rect 1975 3068 1979 3072
rect 2483 3067 2487 3071
rect 2779 3067 2783 3071
rect 3075 3067 3079 3071
rect 3371 3067 3375 3071
rect 3651 3067 3655 3071
rect 3799 3068 3803 3072
rect 1975 3051 1979 3055
rect 2511 3052 2515 3056
rect 2607 3051 2608 3055
rect 2608 3051 2611 3055
rect 2807 3052 2811 3056
rect 2899 3051 2903 3055
rect 3103 3052 3107 3056
rect 3379 3051 3383 3055
rect 3399 3052 3403 3056
rect 3659 3051 3663 3055
rect 3679 3052 3683 3056
rect 3771 3051 3775 3055
rect 3799 3051 3803 3055
rect 3839 3052 3843 3056
rect 3931 3051 3935 3055
rect 4131 3051 4135 3055
rect 4331 3051 4335 3055
rect 4523 3051 4527 3055
rect 4715 3051 4719 3055
rect 4915 3051 4919 3055
rect 5663 3052 5667 3056
rect 111 3040 115 3044
rect 131 3039 135 3043
rect 307 3039 311 3043
rect 507 3039 511 3043
rect 707 3039 711 3043
rect 899 3039 903 3043
rect 1091 3039 1095 3043
rect 1275 3039 1279 3043
rect 1451 3039 1455 3043
rect 1627 3039 1631 3043
rect 1787 3039 1791 3043
rect 1935 3040 1939 3044
rect 499 3031 503 3035
rect 1267 3031 1271 3035
rect 3839 3035 3843 3039
rect 3959 3036 3963 3040
rect 4051 3035 4055 3039
rect 4159 3036 4163 3040
rect 4339 3035 4343 3039
rect 4359 3036 4363 3040
rect 4467 3035 4471 3039
rect 4551 3036 4555 3040
rect 4723 3035 4727 3039
rect 4743 3036 4747 3040
rect 4923 3035 4927 3039
rect 4943 3036 4947 3040
rect 5039 3035 5040 3039
rect 5040 3035 5043 3039
rect 5663 3035 5667 3039
rect 111 3023 115 3027
rect 159 3024 163 3028
rect 251 3023 255 3027
rect 335 3024 339 3028
rect 431 3023 432 3027
rect 432 3023 435 3027
rect 535 3024 539 3028
rect 735 3024 739 3028
rect 907 3023 911 3027
rect 927 3024 931 3028
rect 1027 3023 1028 3027
rect 1028 3023 1031 3027
rect 1119 3024 1123 3028
rect 1283 3023 1287 3027
rect 1303 3024 1307 3028
rect 1459 3023 1463 3027
rect 1479 3024 1483 3028
rect 1575 3023 1576 3027
rect 1576 3023 1579 3027
rect 1655 3024 1659 3028
rect 1815 3024 1819 3028
rect 1935 3023 1939 3027
rect 1975 2985 1979 2989
rect 2191 2984 2195 2988
rect 2287 2983 2288 2987
rect 2288 2983 2291 2987
rect 2351 2984 2355 2988
rect 2447 2983 2448 2987
rect 2448 2983 2451 2987
rect 2519 2984 2523 2988
rect 2639 2983 2643 2987
rect 2703 2984 2707 2988
rect 2795 2983 2799 2987
rect 2903 2984 2907 2988
rect 3003 2983 3004 2987
rect 3004 2983 3007 2987
rect 3119 2984 3123 2988
rect 3215 2983 3216 2987
rect 3216 2983 3219 2987
rect 3335 2984 3339 2988
rect 3427 2983 3431 2987
rect 3559 2984 3563 2988
rect 3651 2983 3655 2987
rect 3799 2985 3803 2989
rect 1975 2968 1979 2972
rect 2163 2969 2167 2973
rect 2323 2969 2327 2973
rect 2491 2969 2495 2973
rect 2675 2969 2679 2973
rect 2875 2969 2879 2973
rect 3091 2969 3095 2973
rect 3307 2969 3311 2973
rect 3531 2969 3535 2973
rect 3799 2968 3803 2972
rect 111 2961 115 2965
rect 159 2960 163 2964
rect 295 2960 299 2964
rect 395 2959 396 2963
rect 396 2959 399 2963
rect 431 2960 435 2964
rect 531 2959 532 2963
rect 532 2959 535 2963
rect 567 2960 571 2964
rect 659 2959 663 2963
rect 703 2960 707 2964
rect 803 2959 804 2963
rect 804 2959 807 2963
rect 1935 2961 1939 2965
rect 3839 2953 3843 2957
rect 3999 2952 4003 2956
rect 111 2944 115 2948
rect 131 2945 135 2949
rect 267 2945 271 2949
rect 403 2945 407 2949
rect 539 2945 543 2949
rect 675 2945 679 2949
rect 1935 2944 1939 2948
rect 2259 2947 2263 2951
rect 4095 2951 4096 2955
rect 4096 2951 4099 2955
rect 4159 2952 4163 2956
rect 2447 2947 2451 2951
rect 4335 2952 4339 2956
rect 4443 2951 4447 2955
rect 4519 2952 4523 2956
rect 4619 2951 4620 2955
rect 4620 2951 4623 2955
rect 4719 2952 4723 2956
rect 4819 2951 4820 2955
rect 4820 2951 4823 2955
rect 4927 2952 4931 2956
rect 5019 2951 5023 2955
rect 5135 2952 5139 2956
rect 5287 2951 5291 2955
rect 5351 2952 5355 2956
rect 5483 2951 5487 2955
rect 5543 2952 5547 2956
rect 5635 2951 5639 2955
rect 5663 2953 5667 2957
rect 3839 2936 3843 2940
rect 3971 2937 3975 2941
rect 4131 2937 4135 2941
rect 4307 2937 4311 2941
rect 4491 2937 4495 2941
rect 4691 2937 4695 2941
rect 4899 2937 4903 2941
rect 5107 2937 5111 2941
rect 5323 2937 5327 2941
rect 5515 2937 5519 2941
rect 5663 2936 5667 2940
rect 2259 2919 2263 2923
rect 2607 2919 2611 2923
rect 2639 2919 2643 2923
rect 2959 2919 2963 2923
rect 3003 2919 3007 2923
rect 2795 2911 2799 2915
rect 3771 2919 3775 2923
rect 3651 2911 3655 2915
rect 251 2895 255 2899
rect 395 2895 399 2899
rect 531 2895 535 2899
rect 759 2895 763 2899
rect 2091 2879 2095 2883
rect 2139 2879 2143 2883
rect 2287 2883 2291 2887
rect 2411 2879 2415 2883
rect 2547 2879 2551 2883
rect 2719 2883 2723 2887
rect 2843 2879 2847 2883
rect 3147 2883 3151 2887
rect 3307 2883 3311 2887
rect 3427 2883 3431 2887
rect 3983 2887 3987 2891
rect 4467 2887 4471 2891
rect 4619 2887 4623 2891
rect 4819 2887 4823 2891
rect 5019 2879 5023 2883
rect 5287 2887 5291 2891
rect 5483 2887 5487 2891
rect 5375 2879 5379 2883
rect 659 2867 663 2871
rect 371 2855 375 2859
rect 507 2855 511 2859
rect 895 2859 899 2863
rect 2091 2851 2095 2855
rect 2663 2851 2667 2855
rect 1975 2832 1979 2836
rect 1995 2831 1999 2835
rect 2131 2831 2135 2835
rect 2267 2831 2271 2835
rect 2403 2831 2407 2835
rect 2539 2831 2543 2835
rect 2683 2831 2687 2835
rect 2835 2831 2839 2835
rect 2995 2831 2999 2835
rect 3155 2831 3159 2835
rect 3315 2831 3319 2835
rect 3799 2832 3803 2836
rect 3955 2835 3959 2839
rect 4203 2839 4207 2843
rect 4443 2839 4447 2843
rect 4699 2835 4703 2839
rect 4971 2835 4975 2839
rect 5391 2839 5395 2843
rect 5635 2839 5639 2843
rect 3147 2823 3151 2827
rect 3307 2823 3311 2827
rect 1975 2815 1979 2819
rect 2023 2816 2027 2820
rect 2139 2815 2143 2819
rect 2159 2816 2163 2820
rect 2251 2815 2255 2819
rect 2295 2816 2299 2820
rect 2411 2815 2415 2819
rect 2431 2816 2435 2820
rect 2547 2815 2551 2819
rect 2567 2816 2571 2820
rect 2663 2815 2664 2819
rect 2664 2815 2667 2819
rect 2711 2816 2715 2820
rect 2843 2815 2847 2819
rect 2863 2816 2867 2820
rect 2959 2815 2960 2819
rect 2960 2815 2963 2819
rect 3023 2816 3027 2820
rect 3119 2815 3120 2819
rect 3120 2815 3123 2819
rect 3183 2816 3187 2820
rect 3343 2816 3347 2820
rect 3799 2815 3803 2819
rect 111 2808 115 2812
rect 227 2807 231 2811
rect 363 2807 367 2811
rect 499 2807 503 2811
rect 635 2807 639 2811
rect 771 2807 775 2811
rect 1935 2808 1939 2812
rect 111 2791 115 2795
rect 255 2792 259 2796
rect 371 2791 375 2795
rect 391 2792 395 2796
rect 507 2791 511 2795
rect 527 2792 531 2796
rect 663 2792 667 2796
rect 759 2791 760 2795
rect 760 2791 763 2795
rect 799 2792 803 2796
rect 1935 2791 1939 2795
rect 3839 2788 3843 2792
rect 3859 2787 3863 2791
rect 4011 2787 4015 2791
rect 4211 2787 4215 2791
rect 4435 2787 4439 2791
rect 4691 2787 4695 2791
rect 4963 2787 4967 2791
rect 5251 2787 5255 2791
rect 5515 2787 5519 2791
rect 5663 2788 5667 2792
rect 919 2775 923 2779
rect 4203 2779 4207 2783
rect 3839 2771 3843 2775
rect 3887 2772 3891 2776
rect 3983 2771 3984 2775
rect 3984 2771 3987 2775
rect 4039 2772 4043 2776
rect 4239 2772 4243 2776
rect 4463 2772 4467 2776
rect 4699 2771 4703 2775
rect 4719 2772 4723 2776
rect 4971 2771 4975 2775
rect 4991 2772 4995 2776
rect 5279 2772 5283 2776
rect 5375 2771 5376 2775
rect 5376 2771 5379 2775
rect 5543 2772 5547 2776
rect 5643 2771 5644 2775
rect 5644 2771 5647 2775
rect 5663 2771 5667 2775
rect 1975 2753 1979 2757
rect 2023 2752 2027 2756
rect 2115 2751 2119 2755
rect 2159 2752 2163 2756
rect 2259 2751 2260 2755
rect 2260 2751 2263 2755
rect 2303 2752 2307 2756
rect 2403 2751 2404 2755
rect 2404 2751 2407 2755
rect 2463 2752 2467 2756
rect 2559 2751 2560 2755
rect 2560 2751 2563 2755
rect 2623 2752 2627 2756
rect 2719 2751 2720 2755
rect 2720 2751 2723 2755
rect 2783 2752 2787 2756
rect 2875 2751 2879 2755
rect 2943 2752 2947 2756
rect 3035 2751 3039 2755
rect 3103 2752 3107 2756
rect 3199 2751 3200 2755
rect 3200 2751 3203 2755
rect 3799 2753 3803 2757
rect 1975 2736 1979 2740
rect 1995 2737 1999 2741
rect 2131 2737 2135 2741
rect 2275 2737 2279 2741
rect 2435 2737 2439 2741
rect 2595 2737 2599 2741
rect 2755 2737 2759 2741
rect 2915 2737 2919 2741
rect 3075 2737 3079 2741
rect 3799 2736 3803 2740
rect 3955 2739 3959 2743
rect 4063 2739 4067 2743
rect 111 2729 115 2733
rect 375 2728 379 2732
rect 475 2727 476 2731
rect 476 2727 479 2731
rect 575 2728 579 2732
rect 675 2727 676 2731
rect 676 2727 679 2731
rect 799 2728 803 2732
rect 895 2727 896 2731
rect 896 2727 899 2731
rect 1039 2728 1043 2732
rect 1295 2728 1299 2732
rect 1387 2727 1391 2731
rect 1567 2728 1571 2732
rect 1659 2727 1663 2731
rect 1815 2728 1819 2732
rect 1911 2727 1912 2731
rect 1912 2727 1915 2731
rect 1935 2729 1939 2733
rect 111 2712 115 2716
rect 347 2713 351 2717
rect 547 2713 551 2717
rect 771 2713 775 2717
rect 1011 2713 1015 2717
rect 1267 2713 1271 2717
rect 1539 2713 1543 2717
rect 1787 2713 1791 2717
rect 1935 2712 1939 2716
rect 4363 2715 4367 2719
rect 3839 2701 3843 2705
rect 3967 2700 3971 2704
rect 4063 2699 4064 2703
rect 4064 2699 4067 2703
rect 4223 2700 4227 2704
rect 4423 2699 4427 2703
rect 4527 2700 4531 2704
rect 4627 2699 4628 2703
rect 4628 2699 4631 2703
rect 4863 2700 4867 2704
rect 4983 2699 4987 2703
rect 5215 2700 5219 2704
rect 5543 2700 5547 2704
rect 5635 2699 5639 2703
rect 5663 2701 5667 2705
rect 2251 2687 2255 2691
rect 2259 2687 2263 2691
rect 2403 2687 2407 2691
rect 2559 2679 2563 2683
rect 2823 2687 2827 2691
rect 2875 2679 2879 2683
rect 3119 2687 3123 2691
rect 3839 2684 3843 2688
rect 3939 2685 3943 2689
rect 4195 2685 4199 2689
rect 4499 2685 4503 2689
rect 4835 2685 4839 2689
rect 5187 2685 5191 2689
rect 5515 2685 5519 2689
rect 5663 2684 5667 2688
rect 3199 2679 3203 2683
rect 475 2663 479 2667
rect 675 2663 679 2667
rect 919 2663 923 2667
rect 507 2655 511 2659
rect 2115 2663 2119 2667
rect 1911 2655 1915 2659
rect 3035 2655 3039 2659
rect 663 2635 667 2639
rect 635 2627 639 2631
rect 855 2631 859 2635
rect 1159 2639 1163 2643
rect 1387 2643 1391 2647
rect 2795 2643 2799 2647
rect 2979 2643 2983 2647
rect 1495 2635 1499 2639
rect 1467 2627 1471 2631
rect 1659 2631 1663 2635
rect 1723 2627 1727 2631
rect 4423 2635 4427 2639
rect 4627 2635 4631 2639
rect 4983 2635 4987 2639
rect 5643 2635 5647 2639
rect 4187 2627 4191 2631
rect 1467 2599 1471 2603
rect 1839 2599 1843 2603
rect 1975 2596 1979 2600
rect 2699 2595 2703 2599
rect 2835 2595 2839 2599
rect 2971 2595 2975 2599
rect 3799 2596 3803 2600
rect 3987 2599 3991 2603
rect 4075 2599 4079 2603
rect 4363 2603 4367 2607
rect 4499 2599 4503 2603
rect 4739 2599 4743 2603
rect 5003 2599 5007 2603
rect 5443 2603 5447 2607
rect 5635 2603 5639 2607
rect 111 2580 115 2584
rect 387 2579 391 2583
rect 539 2579 543 2583
rect 699 2579 703 2583
rect 867 2579 871 2583
rect 1035 2579 1039 2583
rect 1203 2579 1207 2583
rect 1371 2579 1375 2583
rect 1539 2579 1543 2583
rect 1715 2579 1719 2583
rect 1935 2580 1939 2584
rect 1975 2579 1979 2583
rect 2727 2580 2731 2584
rect 2823 2579 2824 2583
rect 2824 2579 2827 2583
rect 2863 2580 2867 2584
rect 2979 2579 2983 2583
rect 2999 2580 3003 2584
rect 3095 2579 3096 2583
rect 3096 2579 3099 2583
rect 3799 2579 3803 2583
rect 855 2571 859 2575
rect 111 2563 115 2567
rect 415 2564 419 2568
rect 507 2563 511 2567
rect 567 2564 571 2568
rect 663 2563 664 2567
rect 664 2563 667 2567
rect 727 2564 731 2568
rect 823 2563 824 2567
rect 824 2563 827 2567
rect 895 2564 899 2568
rect 1063 2564 1067 2568
rect 1159 2563 1160 2567
rect 1160 2563 1163 2567
rect 1231 2564 1235 2568
rect 1327 2563 1328 2567
rect 1328 2563 1331 2567
rect 1399 2564 1403 2568
rect 1495 2563 1496 2567
rect 1496 2563 1499 2567
rect 1567 2564 1571 2568
rect 1723 2563 1727 2567
rect 1743 2564 1747 2568
rect 1839 2563 1840 2567
rect 1840 2563 1843 2567
rect 1935 2563 1939 2567
rect 3839 2552 3843 2556
rect 3891 2551 3895 2555
rect 4067 2551 4071 2555
rect 4267 2551 4271 2555
rect 4491 2551 4495 2555
rect 4731 2551 4735 2555
rect 4995 2551 4999 2555
rect 5267 2551 5271 2555
rect 5515 2551 5519 2555
rect 5663 2552 5667 2556
rect 2795 2535 2799 2539
rect 1975 2521 1979 2525
rect 3839 2535 3843 2539
rect 3919 2536 3923 2540
rect 4075 2535 4079 2539
rect 4095 2536 4099 2540
rect 4187 2535 4191 2539
rect 4295 2536 4299 2540
rect 4499 2535 4503 2539
rect 4519 2536 4523 2540
rect 4739 2535 4743 2539
rect 4759 2536 4763 2540
rect 5003 2535 5007 2539
rect 5023 2536 5027 2540
rect 5115 2535 5119 2539
rect 5295 2536 5299 2540
rect 5391 2535 5392 2539
rect 5392 2535 5395 2539
rect 5543 2536 5547 2540
rect 5635 2535 5639 2539
rect 5663 2535 5667 2539
rect 2607 2520 2611 2524
rect 2703 2519 2704 2523
rect 2704 2519 2707 2523
rect 2759 2520 2763 2524
rect 2911 2520 2915 2524
rect 3003 2519 3007 2523
rect 3063 2520 3067 2524
rect 3163 2519 3164 2523
rect 3164 2519 3167 2523
rect 3223 2520 3227 2524
rect 3319 2519 3320 2523
rect 3320 2519 3323 2523
rect 3799 2521 3803 2525
rect 111 2505 115 2509
rect 327 2504 331 2508
rect 427 2503 428 2507
rect 428 2503 431 2507
rect 535 2504 539 2508
rect 635 2503 636 2507
rect 636 2503 639 2507
rect 735 2504 739 2508
rect 919 2504 923 2508
rect 1031 2503 1035 2507
rect 1095 2504 1099 2508
rect 1187 2503 1191 2507
rect 1271 2504 1275 2508
rect 1371 2503 1372 2507
rect 1372 2503 1375 2507
rect 1439 2504 1443 2508
rect 1539 2503 1540 2507
rect 1540 2503 1543 2507
rect 1607 2504 1611 2508
rect 1707 2503 1708 2507
rect 1708 2503 1711 2507
rect 1775 2504 1779 2508
rect 1867 2503 1871 2507
rect 1935 2505 1939 2509
rect 1975 2504 1979 2508
rect 2579 2505 2583 2509
rect 2731 2505 2735 2509
rect 2883 2505 2887 2509
rect 3035 2505 3039 2509
rect 3195 2505 3199 2509
rect 3799 2504 3803 2508
rect 111 2488 115 2492
rect 299 2489 303 2493
rect 507 2489 511 2493
rect 707 2489 711 2493
rect 891 2489 895 2493
rect 1067 2489 1071 2493
rect 1243 2489 1247 2493
rect 1411 2489 1415 2493
rect 1579 2489 1583 2493
rect 1747 2489 1751 2493
rect 1935 2488 1939 2492
rect 3839 2473 3843 2477
rect 3887 2472 3891 2476
rect 3987 2471 3988 2475
rect 3988 2471 3991 2475
rect 4087 2472 4091 2476
rect 4183 2471 4184 2475
rect 4184 2471 4187 2475
rect 4319 2472 4323 2476
rect 4439 2471 4443 2475
rect 4567 2472 4571 2476
rect 4711 2471 4715 2475
rect 4823 2472 4827 2476
rect 4975 2471 4979 2475
rect 5087 2472 5091 2476
rect 5351 2472 5355 2476
rect 5443 2471 5447 2475
rect 5663 2473 5667 2477
rect 2691 2455 2695 2459
rect 2703 2455 2707 2459
rect 3095 2455 3099 2459
rect 3163 2455 3167 2459
rect 3839 2456 3843 2460
rect 3859 2457 3863 2461
rect 4059 2457 4063 2461
rect 4291 2457 4295 2461
rect 4539 2457 4543 2461
rect 4795 2457 4799 2461
rect 5059 2457 5063 2461
rect 5323 2457 5327 2461
rect 5663 2456 5667 2460
rect 3319 2447 3323 2451
rect 427 2439 431 2443
rect 823 2439 827 2443
rect 1031 2439 1035 2443
rect 1327 2439 1331 2443
rect 1371 2439 1375 2443
rect 1539 2439 1543 2443
rect 1707 2439 1711 2443
rect 227 2399 231 2403
rect 519 2403 523 2407
rect 699 2399 703 2403
rect 1187 2403 1191 2407
rect 1867 2411 1871 2415
rect 1915 2407 1919 2411
rect 2703 2411 2707 2415
rect 1259 2399 1263 2403
rect 1795 2399 1799 2403
rect 2579 2403 2583 2407
rect 3003 2407 3007 2411
rect 3155 2403 3159 2407
rect 3443 2403 3447 2407
rect 4211 2407 4215 2411
rect 4387 2407 4391 2411
rect 4439 2407 4443 2411
rect 4711 2407 4715 2411
rect 4975 2407 4979 2411
rect 5407 2407 5411 2411
rect 4183 2399 4187 2403
rect 227 2371 231 2375
rect 815 2371 819 2375
rect 3791 2375 3795 2379
rect 4099 2371 4103 2375
rect 4587 2371 4591 2375
rect 4819 2371 4823 2375
rect 5051 2371 5055 2375
rect 5499 2375 5503 2379
rect 5635 2375 5639 2379
rect 111 2352 115 2356
rect 131 2351 135 2355
rect 403 2351 407 2355
rect 691 2351 695 2355
rect 971 2351 975 2355
rect 1251 2351 1255 2355
rect 1531 2351 1535 2355
rect 1787 2351 1791 2355
rect 1935 2352 1939 2356
rect 1975 2356 1979 2360
rect 1995 2355 1999 2359
rect 2275 2355 2279 2359
rect 2571 2355 2575 2359
rect 2859 2355 2863 2359
rect 3147 2355 3151 2359
rect 3435 2355 3439 2359
rect 3799 2356 3803 2360
rect 111 2335 115 2339
rect 159 2336 163 2340
rect 431 2336 435 2340
rect 699 2335 703 2339
rect 719 2336 723 2340
rect 815 2335 816 2339
rect 816 2335 819 2339
rect 999 2336 1003 2340
rect 1259 2335 1263 2339
rect 1279 2336 1283 2340
rect 1375 2335 1376 2339
rect 1376 2335 1379 2339
rect 1559 2336 1563 2340
rect 1795 2335 1799 2339
rect 1815 2336 1819 2340
rect 1915 2335 1916 2339
rect 1916 2335 1919 2339
rect 1935 2335 1939 2339
rect 1975 2339 1979 2343
rect 2023 2340 2027 2344
rect 2115 2339 2119 2343
rect 2303 2340 2307 2344
rect 2579 2339 2583 2343
rect 2599 2340 2603 2344
rect 2691 2339 2695 2343
rect 2887 2340 2891 2344
rect 3155 2339 3159 2343
rect 3175 2340 3179 2344
rect 3443 2339 3447 2343
rect 3463 2340 3467 2344
rect 3559 2339 3560 2343
rect 3560 2339 3563 2343
rect 3799 2339 3803 2343
rect 3839 2324 3843 2328
rect 3859 2323 3863 2327
rect 4091 2323 4095 2327
rect 4339 2323 4343 2327
rect 4579 2323 4583 2327
rect 4811 2323 4815 2327
rect 5043 2323 5047 2327
rect 5283 2323 5287 2327
rect 5515 2323 5519 2327
rect 5663 2324 5667 2328
rect 3839 2307 3843 2311
rect 3887 2308 3891 2312
rect 4099 2307 4103 2311
rect 4119 2308 4123 2312
rect 4211 2307 4215 2311
rect 4367 2308 4371 2312
rect 4587 2307 4591 2311
rect 4607 2308 4611 2312
rect 4819 2307 4823 2311
rect 4839 2308 4843 2312
rect 5051 2307 5055 2311
rect 5071 2308 5075 2312
rect 5167 2307 5168 2311
rect 5168 2307 5171 2311
rect 5311 2308 5315 2312
rect 5407 2307 5408 2311
rect 5408 2307 5411 2311
rect 5543 2308 5547 2312
rect 5635 2307 5639 2311
rect 5663 2307 5667 2311
rect 1975 2269 1979 2273
rect 2023 2268 2027 2272
rect 2123 2267 2124 2271
rect 2124 2267 2127 2271
rect 2159 2268 2163 2272
rect 2259 2267 2260 2271
rect 2260 2267 2263 2271
rect 2295 2268 2299 2272
rect 2447 2268 2451 2272
rect 2539 2267 2543 2271
rect 2607 2268 2611 2272
rect 2703 2267 2704 2271
rect 2704 2267 2707 2271
rect 2767 2268 2771 2272
rect 2859 2267 2863 2271
rect 2927 2268 2931 2272
rect 3019 2267 3023 2271
rect 3079 2268 3083 2272
rect 3175 2267 3176 2271
rect 3176 2267 3179 2271
rect 3231 2268 3235 2272
rect 3327 2267 3328 2271
rect 3328 2267 3331 2271
rect 3383 2268 3387 2272
rect 3479 2267 3480 2271
rect 3480 2267 3483 2271
rect 3543 2268 3547 2272
rect 3643 2267 3644 2271
rect 3644 2267 3647 2271
rect 3679 2268 3683 2272
rect 3791 2267 3795 2271
rect 3799 2269 3803 2273
rect 111 2261 115 2265
rect 159 2260 163 2264
rect 423 2260 427 2264
rect 519 2259 520 2263
rect 520 2259 523 2263
rect 711 2260 715 2264
rect 811 2259 812 2263
rect 812 2259 815 2263
rect 999 2260 1003 2264
rect 1095 2259 1096 2263
rect 1096 2259 1099 2263
rect 1295 2260 1299 2264
rect 1387 2259 1391 2263
rect 1935 2261 1939 2265
rect 1975 2252 1979 2256
rect 1995 2253 1999 2257
rect 2131 2253 2135 2257
rect 2267 2253 2271 2257
rect 2419 2253 2423 2257
rect 2579 2253 2583 2257
rect 2739 2253 2743 2257
rect 2899 2253 2903 2257
rect 3051 2253 3055 2257
rect 3203 2253 3207 2257
rect 3355 2253 3359 2257
rect 3515 2253 3519 2257
rect 3651 2253 3655 2257
rect 3799 2252 3803 2256
rect 111 2244 115 2248
rect 131 2245 135 2249
rect 395 2245 399 2249
rect 683 2245 687 2249
rect 971 2245 975 2249
rect 1267 2245 1271 2249
rect 1935 2244 1939 2248
rect 3147 2235 3151 2239
rect 3327 2235 3331 2239
rect 3839 2225 3843 2229
rect 4591 2224 4595 2228
rect 4691 2223 4692 2227
rect 4692 2223 4695 2227
rect 4727 2224 4731 2228
rect 4827 2223 4828 2227
rect 4828 2223 4831 2227
rect 4863 2224 4867 2228
rect 4963 2223 4964 2227
rect 4964 2223 4967 2227
rect 4999 2224 5003 2228
rect 5099 2223 5100 2227
rect 5100 2223 5103 2227
rect 5135 2224 5139 2228
rect 5235 2223 5236 2227
rect 5236 2223 5239 2227
rect 5271 2224 5275 2228
rect 5371 2223 5372 2227
rect 5372 2223 5375 2227
rect 5407 2224 5411 2228
rect 5499 2223 5503 2227
rect 5543 2224 5547 2228
rect 5643 2223 5644 2227
rect 5644 2223 5647 2227
rect 5663 2225 5667 2229
rect 3839 2208 3843 2212
rect 4563 2209 4567 2213
rect 4699 2209 4703 2213
rect 4835 2209 4839 2213
rect 4971 2209 4975 2213
rect 5107 2209 5111 2213
rect 5243 2209 5247 2213
rect 5379 2209 5383 2213
rect 5515 2209 5519 2213
rect 5663 2208 5667 2212
rect 2115 2203 2119 2207
rect 2123 2203 2127 2207
rect 2259 2203 2263 2207
rect 251 2195 255 2199
rect 811 2195 815 2199
rect 1375 2195 1379 2199
rect 2851 2203 2855 2207
rect 2859 2195 2863 2199
rect 3147 2203 3151 2207
rect 3175 2195 3179 2199
rect 3423 2203 3427 2207
rect 3559 2203 3563 2207
rect 3643 2203 3647 2207
rect 3479 2195 3483 2199
rect 1387 2187 1391 2191
rect 2539 2171 2543 2175
rect 527 2155 531 2159
rect 2339 2159 2343 2163
rect 2539 2159 2543 2163
rect 2739 2159 2743 2163
rect 3019 2163 3023 2167
rect 3775 2171 3779 2175
rect 3123 2159 3127 2163
rect 3579 2159 3583 2163
rect 3659 2159 3663 2163
rect 499 2147 503 2151
rect 739 2147 743 2151
rect 1095 2151 1099 2155
rect 1451 2147 1455 2151
rect 2119 2151 2123 2155
rect 4691 2159 4695 2163
rect 4827 2159 4831 2163
rect 4963 2159 4967 2163
rect 5099 2159 5103 2163
rect 5235 2159 5239 2163
rect 5371 2159 5375 2163
rect 5635 2159 5639 2163
rect 5167 2151 5171 2155
rect 5351 2119 5355 2123
rect 499 2111 503 2115
rect 855 2111 859 2115
rect 1975 2112 1979 2116
rect 2131 2111 2135 2115
rect 2331 2111 2335 2115
rect 2531 2111 2535 2115
rect 2731 2111 2735 2115
rect 2923 2111 2927 2115
rect 3115 2111 3119 2115
rect 3299 2111 3303 2115
rect 3483 2111 3487 2115
rect 3651 2111 3655 2115
rect 3799 2112 3803 2116
rect 5083 2111 5087 2115
rect 5411 2111 5415 2115
rect 111 2100 115 2104
rect 131 2099 135 2103
rect 403 2099 407 2103
rect 731 2099 735 2103
rect 1083 2099 1087 2103
rect 1443 2099 1447 2103
rect 1787 2099 1791 2103
rect 1935 2100 1939 2104
rect 1975 2095 1979 2099
rect 2159 2096 2163 2100
rect 2339 2095 2343 2099
rect 2359 2096 2363 2100
rect 2539 2095 2543 2099
rect 2559 2096 2563 2100
rect 2739 2095 2743 2099
rect 2759 2096 2763 2100
rect 2851 2095 2855 2099
rect 2951 2096 2955 2100
rect 3123 2095 3127 2099
rect 3143 2096 3147 2100
rect 3239 2095 3240 2099
rect 3240 2095 3243 2099
rect 3327 2096 3331 2100
rect 3423 2095 3424 2099
rect 3424 2095 3427 2099
rect 3511 2096 3515 2100
rect 3659 2095 3663 2099
rect 3679 2096 3683 2100
rect 3775 2095 3776 2099
rect 3776 2095 3779 2099
rect 3799 2095 3803 2099
rect 111 2083 115 2087
rect 159 2084 163 2088
rect 251 2083 255 2087
rect 431 2084 435 2088
rect 527 2083 528 2087
rect 528 2083 531 2087
rect 759 2084 763 2088
rect 855 2083 856 2087
rect 856 2083 859 2087
rect 1111 2084 1115 2088
rect 1451 2083 1455 2087
rect 1471 2084 1475 2088
rect 1567 2083 1568 2087
rect 1568 2083 1571 2087
rect 1815 2084 1819 2088
rect 1911 2083 1912 2087
rect 1912 2083 1915 2087
rect 1935 2083 1939 2087
rect 3839 2060 3843 2064
rect 4955 2059 4959 2063
rect 5091 2059 5095 2063
rect 5227 2059 5231 2063
rect 5663 2060 5667 2064
rect 5083 2051 5087 2055
rect 3839 2043 3843 2047
rect 4983 2044 4987 2048
rect 5075 2043 5079 2047
rect 5119 2044 5123 2048
rect 5255 2044 5259 2048
rect 5351 2043 5352 2047
rect 5352 2043 5355 2047
rect 5663 2043 5667 2047
rect 1975 2029 1979 2033
rect 2023 2028 2027 2032
rect 2119 2027 2120 2031
rect 2120 2027 2123 2031
rect 2279 2028 2283 2032
rect 2375 2027 2376 2031
rect 2376 2027 2379 2031
rect 2551 2028 2555 2032
rect 2647 2027 2648 2031
rect 2648 2027 2651 2031
rect 2799 2028 2803 2032
rect 2891 2027 2895 2031
rect 3031 2028 3035 2032
rect 3123 2027 3127 2031
rect 3255 2028 3259 2032
rect 3351 2027 3352 2031
rect 3352 2027 3355 2031
rect 3479 2028 3483 2032
rect 3579 2027 3580 2031
rect 3580 2027 3583 2031
rect 3679 2028 3683 2032
rect 3771 2027 3775 2031
rect 3799 2029 3803 2033
rect 111 2021 115 2025
rect 223 2020 227 2024
rect 323 2019 324 2023
rect 324 2019 327 2023
rect 383 2020 387 2024
rect 559 2020 563 2024
rect 739 2019 743 2023
rect 751 2020 755 2024
rect 843 2019 847 2023
rect 959 2020 963 2024
rect 1055 2019 1056 2023
rect 1056 2019 1059 2023
rect 1167 2020 1171 2024
rect 1259 2019 1263 2023
rect 1383 2020 1387 2024
rect 1483 2019 1484 2023
rect 1484 2019 1487 2023
rect 1607 2020 1611 2024
rect 1703 2019 1704 2023
rect 1704 2019 1707 2023
rect 1815 2020 1819 2024
rect 1935 2021 1939 2025
rect 111 2004 115 2008
rect 195 2005 199 2009
rect 355 2005 359 2009
rect 531 2005 535 2009
rect 723 2005 727 2009
rect 931 2005 935 2009
rect 1139 2005 1143 2009
rect 1355 2005 1359 2009
rect 1579 2005 1583 2009
rect 1787 2005 1791 2009
rect 1235 1999 1239 2003
rect 1567 1999 1571 2003
rect 1675 1999 1679 2003
rect 1975 2012 1979 2016
rect 1995 2013 1999 2017
rect 2251 2013 2255 2017
rect 2523 2013 2527 2017
rect 2771 2013 2775 2017
rect 3003 2013 3007 2017
rect 3227 2013 3231 2017
rect 3451 2013 3455 2017
rect 3651 2013 3655 2017
rect 3799 2012 3803 2016
rect 1935 2004 1939 2008
rect 2867 1999 2871 2003
rect 3123 1999 3127 2003
rect 3547 1995 3551 1999
rect 3771 1995 3775 1999
rect 1027 1983 1031 1987
rect 1259 1983 1263 1987
rect 3839 1985 3843 1989
rect 4727 1984 4731 1988
rect 4827 1983 4828 1987
rect 4828 1983 4831 1987
rect 4863 1984 4867 1988
rect 4971 1983 4975 1987
rect 5007 1984 5011 1988
rect 5159 1984 5163 1988
rect 5251 1983 5255 1987
rect 5319 1984 5323 1988
rect 5411 1983 5415 1987
rect 5487 1984 5491 1988
rect 5583 1983 5584 1987
rect 5584 1983 5587 1987
rect 5663 1985 5667 1989
rect 3839 1968 3843 1972
rect 4699 1969 4703 1973
rect 4835 1969 4839 1973
rect 4979 1969 4983 1973
rect 5131 1969 5135 1973
rect 5291 1969 5295 1973
rect 5459 1969 5463 1973
rect 5663 1968 5667 1972
rect 315 1955 319 1959
rect 323 1955 327 1959
rect 1027 1955 1031 1959
rect 1235 1955 1239 1959
rect 1055 1947 1059 1951
rect 1675 1955 1679 1959
rect 1911 1955 1915 1959
rect 2375 1955 2379 1959
rect 2443 1963 2447 1967
rect 2867 1963 2871 1967
rect 2647 1955 2651 1959
rect 3239 1963 3243 1967
rect 3547 1963 3551 1967
rect 3771 1963 3775 1967
rect 3351 1955 3355 1959
rect 1703 1947 1707 1951
rect 507 1919 511 1923
rect 843 1923 847 1927
rect 575 1907 579 1911
rect 827 1911 831 1915
rect 1059 1911 1063 1915
rect 1475 1915 1479 1919
rect 1483 1915 1487 1919
rect 2207 1919 2211 1923
rect 1779 1911 1783 1915
rect 2323 1915 2327 1919
rect 2891 1919 2895 1923
rect 2907 1915 2911 1919
rect 3171 1915 3175 1919
rect 3535 1919 3539 1923
rect 3659 1915 3663 1919
rect 4827 1919 4831 1923
rect 5075 1919 5079 1923
rect 5359 1919 5363 1923
rect 5647 1919 5651 1923
rect 5251 1911 5255 1915
rect 4491 1887 4495 1891
rect 4507 1883 4511 1887
rect 4739 1883 4743 1887
rect 4971 1887 4975 1891
rect 5339 1887 5343 1891
rect 5583 1887 5587 1891
rect 111 1864 115 1868
rect 195 1863 199 1867
rect 387 1863 391 1867
rect 595 1863 599 1867
rect 819 1863 823 1867
rect 1051 1863 1055 1867
rect 1283 1863 1287 1867
rect 1523 1863 1527 1867
rect 1771 1863 1775 1867
rect 1935 1864 1939 1868
rect 1975 1868 1979 1872
rect 1995 1867 1999 1871
rect 2315 1867 2319 1871
rect 2619 1867 2623 1871
rect 2899 1867 2903 1871
rect 3163 1867 3167 1871
rect 3419 1867 3423 1871
rect 3651 1867 3655 1871
rect 3799 1868 3803 1872
rect 1475 1855 1479 1859
rect 111 1847 115 1851
rect 223 1848 227 1852
rect 315 1847 319 1851
rect 415 1848 419 1852
rect 507 1847 511 1851
rect 623 1848 627 1852
rect 827 1847 831 1851
rect 847 1848 851 1852
rect 1059 1847 1063 1851
rect 1079 1848 1083 1852
rect 1171 1847 1175 1851
rect 1311 1848 1315 1852
rect 1407 1847 1408 1851
rect 1408 1847 1411 1851
rect 1551 1848 1555 1852
rect 1779 1847 1783 1851
rect 1799 1848 1803 1852
rect 1935 1847 1939 1851
rect 1975 1851 1979 1855
rect 2023 1852 2027 1856
rect 2323 1851 2327 1855
rect 2343 1852 2347 1856
rect 2443 1851 2444 1855
rect 2444 1851 2447 1855
rect 2647 1852 2651 1856
rect 2907 1851 2911 1855
rect 2927 1852 2931 1856
rect 3171 1851 3175 1855
rect 3191 1852 3195 1856
rect 3287 1851 3288 1855
rect 3288 1851 3291 1855
rect 3447 1852 3451 1856
rect 3659 1851 3663 1855
rect 3679 1852 3683 1856
rect 3771 1851 3775 1855
rect 3799 1851 3803 1855
rect 3839 1836 3843 1840
rect 4275 1835 4279 1839
rect 4499 1835 4503 1839
rect 4731 1835 4735 1839
rect 4979 1835 4983 1839
rect 5235 1835 5239 1839
rect 5499 1835 5503 1839
rect 5663 1836 5667 1840
rect 4491 1827 4495 1831
rect 3839 1819 3843 1823
rect 4303 1820 4307 1824
rect 4507 1819 4511 1823
rect 4527 1820 4531 1824
rect 4739 1819 4743 1823
rect 4759 1820 4763 1824
rect 4859 1819 4860 1823
rect 4860 1819 4863 1823
rect 5007 1820 5011 1824
rect 5263 1820 5267 1824
rect 5359 1819 5360 1823
rect 5360 1819 5363 1823
rect 5527 1820 5531 1824
rect 5623 1819 5624 1823
rect 5624 1819 5627 1823
rect 5663 1819 5667 1823
rect 1975 1789 1979 1793
rect 2111 1788 2115 1792
rect 2207 1787 2208 1791
rect 2208 1787 2211 1791
rect 2391 1788 2395 1792
rect 2487 1787 2488 1791
rect 2488 1787 2491 1791
rect 2663 1788 2667 1792
rect 2755 1787 2759 1791
rect 2927 1788 2931 1792
rect 3019 1787 3023 1791
rect 3183 1788 3187 1792
rect 3279 1787 3280 1791
rect 3280 1787 3283 1791
rect 3439 1788 3443 1792
rect 3535 1787 3536 1791
rect 3536 1787 3539 1791
rect 3679 1788 3683 1792
rect 3771 1787 3775 1791
rect 3799 1789 3803 1793
rect 111 1773 115 1777
rect 159 1772 163 1776
rect 267 1771 271 1775
rect 303 1772 307 1776
rect 419 1771 423 1775
rect 479 1772 483 1776
rect 575 1771 576 1775
rect 576 1771 579 1775
rect 655 1772 659 1776
rect 771 1771 775 1775
rect 831 1772 835 1776
rect 927 1771 928 1775
rect 928 1771 931 1775
rect 1007 1772 1011 1776
rect 1099 1771 1103 1775
rect 1183 1772 1187 1776
rect 1291 1771 1295 1775
rect 1359 1772 1363 1776
rect 1471 1771 1475 1775
rect 1535 1772 1539 1776
rect 1647 1771 1651 1775
rect 1711 1772 1715 1776
rect 1807 1771 1808 1775
rect 1808 1771 1811 1775
rect 1935 1773 1939 1777
rect 1975 1772 1979 1776
rect 2083 1773 2087 1777
rect 2363 1773 2367 1777
rect 2635 1773 2639 1777
rect 2899 1773 2903 1777
rect 3155 1773 3159 1777
rect 3411 1773 3415 1777
rect 3651 1773 3655 1777
rect 3799 1772 3803 1776
rect 111 1756 115 1760
rect 131 1757 135 1761
rect 275 1757 279 1761
rect 451 1757 455 1761
rect 627 1757 631 1761
rect 803 1757 807 1761
rect 979 1757 983 1761
rect 1155 1757 1159 1761
rect 1331 1757 1335 1761
rect 1507 1757 1511 1761
rect 1683 1757 1687 1761
rect 1935 1756 1939 1760
rect 3839 1753 3843 1757
rect 3887 1752 3891 1756
rect 3983 1751 3984 1755
rect 3984 1751 3987 1755
rect 4087 1752 4091 1756
rect 4223 1751 4227 1755
rect 4343 1752 4347 1756
rect 4435 1751 4439 1755
rect 4623 1752 4627 1756
rect 4715 1751 4719 1755
rect 4927 1752 4931 1756
rect 5023 1751 5024 1755
rect 5024 1751 5027 1755
rect 5247 1752 5251 1756
rect 5339 1751 5343 1755
rect 5543 1752 5547 1756
rect 5635 1751 5639 1755
rect 5663 1753 5667 1757
rect 723 1735 727 1739
rect 1099 1735 1103 1739
rect 3839 1736 3843 1740
rect 3859 1737 3863 1741
rect 4059 1737 4063 1741
rect 4315 1737 4319 1741
rect 4595 1737 4599 1741
rect 4899 1737 4903 1741
rect 5219 1737 5223 1741
rect 5515 1737 5519 1741
rect 5663 1736 5667 1740
rect 2611 1723 2615 1727
rect 2487 1715 2491 1719
rect 3019 1715 3023 1719
rect 3287 1723 3291 1727
rect 3279 1715 3283 1719
rect 3983 1723 3987 1727
rect 3771 1715 3775 1719
rect 251 1707 255 1711
rect 267 1707 271 1711
rect 419 1707 423 1711
rect 723 1707 727 1711
rect 771 1707 775 1711
rect 1171 1699 1175 1703
rect 1407 1707 1411 1711
rect 1471 1707 1475 1711
rect 1647 1707 1651 1711
rect 1807 1699 1811 1703
rect 3979 1687 3983 1691
rect 4223 1687 4227 1691
rect 927 1671 931 1675
rect 1267 1675 1271 1679
rect 4715 1679 4719 1683
rect 4859 1687 4863 1691
rect 5395 1687 5399 1691
rect 5623 1687 5627 1691
rect 5023 1679 5027 1683
rect 1243 1667 1247 1671
rect 1291 1671 1295 1675
rect 1427 1667 1431 1671
rect 1563 1667 1567 1671
rect 2179 1655 2183 1659
rect 2227 1655 2231 1659
rect 2363 1655 2367 1659
rect 2499 1655 2503 1659
rect 2755 1659 2759 1663
rect 2779 1655 2783 1659
rect 2923 1655 2927 1659
rect 4263 1655 4267 1659
rect 4003 1647 4007 1651
rect 4147 1647 4151 1651
rect 4435 1651 4439 1655
rect 4539 1647 4543 1651
rect 4771 1647 4775 1651
rect 5019 1647 5023 1651
rect 5403 1651 5407 1655
rect 5635 1651 5639 1655
rect 1243 1639 1247 1643
rect 1679 1639 1683 1643
rect 111 1620 115 1624
rect 875 1619 879 1623
rect 1011 1619 1015 1623
rect 1147 1619 1151 1623
rect 1283 1619 1287 1623
rect 1419 1619 1423 1623
rect 1555 1619 1559 1623
rect 1935 1620 1939 1624
rect 1975 1608 1979 1612
rect 111 1603 115 1607
rect 903 1604 907 1608
rect 999 1603 1000 1607
rect 1000 1603 1003 1607
rect 1039 1604 1043 1608
rect 1135 1603 1136 1607
rect 1136 1603 1139 1607
rect 1175 1604 1179 1608
rect 1267 1603 1271 1607
rect 1311 1604 1315 1608
rect 1427 1603 1431 1607
rect 1447 1604 1451 1608
rect 1563 1603 1567 1607
rect 1583 1604 1587 1608
rect 1679 1603 1680 1607
rect 1680 1603 1683 1607
rect 2083 1607 2087 1611
rect 1935 1603 1939 1607
rect 2219 1607 2223 1611
rect 2355 1607 2359 1611
rect 2491 1607 2495 1611
rect 2627 1607 2631 1611
rect 2771 1607 2775 1611
rect 2915 1607 2919 1611
rect 3799 1608 3803 1612
rect 3839 1600 3843 1604
rect 3859 1599 3863 1603
rect 3995 1599 3999 1603
rect 4139 1599 4143 1603
rect 4323 1599 4327 1603
rect 4531 1599 4535 1603
rect 4763 1599 4767 1603
rect 5011 1599 5015 1603
rect 5275 1599 5279 1603
rect 5515 1599 5519 1603
rect 5663 1600 5667 1604
rect 1975 1591 1979 1595
rect 2111 1592 2115 1596
rect 2227 1591 2231 1595
rect 2247 1592 2251 1596
rect 2363 1591 2367 1595
rect 2383 1592 2387 1596
rect 2499 1591 2503 1595
rect 2519 1592 2523 1596
rect 2611 1591 2615 1595
rect 2655 1592 2659 1596
rect 2779 1591 2783 1595
rect 2799 1592 2803 1596
rect 2923 1591 2927 1595
rect 2943 1592 2947 1596
rect 3039 1591 3040 1595
rect 3040 1591 3043 1595
rect 3799 1591 3803 1595
rect 3839 1583 3843 1587
rect 3887 1584 3891 1588
rect 3979 1583 3983 1587
rect 4023 1584 4027 1588
rect 4147 1583 4151 1587
rect 4167 1584 4171 1588
rect 4263 1583 4264 1587
rect 4264 1583 4267 1587
rect 4351 1584 4355 1588
rect 4539 1583 4543 1587
rect 4559 1584 4563 1588
rect 4771 1583 4775 1587
rect 4791 1584 4795 1588
rect 5019 1583 5023 1587
rect 5039 1584 5043 1588
rect 5131 1583 5135 1587
rect 5303 1584 5307 1588
rect 5395 1583 5399 1587
rect 5543 1584 5547 1588
rect 5639 1583 5640 1587
rect 5640 1583 5643 1587
rect 5663 1583 5667 1587
rect 2179 1543 2183 1547
rect 111 1525 115 1529
rect 159 1524 163 1528
rect 251 1523 255 1527
rect 391 1524 395 1528
rect 519 1523 523 1527
rect 631 1524 635 1528
rect 731 1523 732 1527
rect 732 1523 735 1527
rect 871 1524 875 1528
rect 991 1523 995 1527
rect 1111 1524 1115 1528
rect 1351 1524 1355 1528
rect 1443 1523 1447 1527
rect 1935 1525 1939 1529
rect 1975 1529 1979 1533
rect 2143 1528 2147 1532
rect 2279 1528 2283 1532
rect 2375 1527 2376 1531
rect 2376 1527 2379 1531
rect 2415 1528 2419 1532
rect 2515 1527 2516 1531
rect 2516 1527 2519 1531
rect 2551 1528 2555 1532
rect 2651 1527 2652 1531
rect 2652 1527 2655 1531
rect 2687 1528 2691 1532
rect 2787 1527 2788 1531
rect 2788 1527 2791 1531
rect 2823 1528 2827 1532
rect 2915 1527 2919 1531
rect 2959 1528 2963 1532
rect 3059 1527 3060 1531
rect 3060 1527 3063 1531
rect 3095 1528 3099 1532
rect 3195 1527 3196 1531
rect 3196 1527 3199 1531
rect 3231 1528 3235 1532
rect 3323 1527 3327 1531
rect 3799 1529 3803 1533
rect 3839 1521 3843 1525
rect 3887 1520 3891 1524
rect 4003 1519 4007 1523
rect 4111 1520 4115 1524
rect 4207 1519 4208 1523
rect 4208 1519 4211 1523
rect 4343 1520 4347 1524
rect 4575 1520 4579 1524
rect 4703 1519 4707 1523
rect 4815 1520 4819 1524
rect 4951 1519 4955 1523
rect 5063 1520 5067 1524
rect 5155 1519 5159 1523
rect 5311 1520 5315 1524
rect 5403 1519 5407 1523
rect 5543 1520 5547 1524
rect 5663 1521 5667 1525
rect 111 1508 115 1512
rect 131 1509 135 1513
rect 363 1509 367 1513
rect 603 1509 607 1513
rect 843 1509 847 1513
rect 1083 1509 1087 1513
rect 1323 1509 1327 1513
rect 1935 1508 1939 1512
rect 1975 1512 1979 1516
rect 2115 1513 2119 1517
rect 2251 1513 2255 1517
rect 2387 1513 2391 1517
rect 2523 1513 2527 1517
rect 2659 1513 2663 1517
rect 2795 1513 2799 1517
rect 2931 1513 2935 1517
rect 3067 1513 3071 1517
rect 3203 1513 3207 1517
rect 3799 1512 3803 1516
rect 459 1503 463 1507
rect 999 1503 1003 1507
rect 3839 1504 3843 1508
rect 3859 1505 3863 1509
rect 4083 1505 4087 1509
rect 4315 1505 4319 1509
rect 4547 1505 4551 1509
rect 4787 1505 4791 1509
rect 5035 1505 5039 1509
rect 5283 1505 5287 1509
rect 5515 1505 5519 1509
rect 5663 1504 5667 1508
rect 3955 1499 3959 1503
rect 4207 1499 4211 1503
rect 4419 1499 4423 1503
rect 5155 1499 5159 1503
rect 2347 1487 2351 1491
rect 2915 1487 2919 1491
rect 4411 1491 4415 1495
rect 5131 1491 5135 1495
rect 459 1459 463 1463
rect 519 1459 523 1463
rect 455 1451 459 1455
rect 1135 1459 1139 1463
rect 2347 1463 2351 1467
rect 1443 1451 1447 1455
rect 2375 1455 2379 1459
rect 2515 1463 2519 1467
rect 2651 1463 2655 1467
rect 2787 1463 2791 1467
rect 3039 1463 3043 1467
rect 3059 1463 3063 1467
rect 3195 1463 3199 1467
rect 2815 1455 2819 1459
rect 3955 1455 3959 1459
rect 4203 1455 4207 1459
rect 4411 1455 4415 1459
rect 4703 1455 4707 1459
rect 4951 1455 4955 1459
rect 5639 1455 5643 1459
rect 5543 1447 5547 1451
rect 3983 1423 3987 1427
rect 255 1415 259 1419
rect 339 1411 343 1415
rect 651 1411 655 1415
rect 731 1415 735 1419
rect 991 1415 995 1419
rect 2195 1411 2199 1415
rect 2251 1411 2255 1415
rect 2395 1411 2399 1415
rect 2547 1411 2551 1415
rect 2699 1411 2703 1415
rect 3323 1415 3327 1419
rect 4091 1419 4095 1423
rect 4419 1423 4423 1427
rect 4555 1419 4559 1423
rect 4779 1419 4783 1423
rect 4995 1419 4999 1423
rect 5211 1419 5215 1423
rect 5535 1423 5539 1427
rect 651 1391 655 1395
rect 1127 1391 1131 1395
rect 3839 1372 3843 1376
rect 3859 1371 3863 1375
rect 4083 1371 4087 1375
rect 4323 1371 4327 1375
rect 4547 1371 4551 1375
rect 4771 1371 4775 1375
rect 4987 1371 4991 1375
rect 5203 1371 5207 1375
rect 5419 1371 5423 1375
rect 5663 1372 5667 1376
rect 111 1364 115 1368
rect 131 1363 135 1367
rect 331 1363 335 1367
rect 555 1363 559 1367
rect 779 1363 783 1367
rect 1003 1363 1007 1367
rect 1935 1364 1939 1368
rect 1975 1364 1979 1368
rect 2099 1363 2103 1367
rect 2243 1363 2247 1367
rect 2387 1363 2391 1367
rect 2539 1363 2543 1367
rect 2691 1363 2695 1367
rect 2851 1363 2855 1367
rect 3011 1363 3015 1367
rect 3171 1363 3175 1367
rect 3799 1364 3803 1368
rect 3839 1355 3843 1359
rect 3887 1356 3891 1360
rect 4091 1355 4095 1359
rect 4111 1356 4115 1360
rect 4203 1355 4207 1359
rect 4351 1356 4355 1360
rect 4555 1355 4559 1359
rect 4575 1356 4579 1360
rect 4779 1355 4783 1359
rect 4799 1356 4803 1360
rect 4995 1355 4999 1359
rect 5015 1356 5019 1360
rect 5211 1355 5215 1359
rect 5231 1356 5235 1360
rect 5323 1355 5327 1359
rect 5447 1356 5451 1360
rect 5543 1355 5544 1359
rect 5544 1355 5547 1359
rect 5663 1355 5667 1359
rect 111 1347 115 1351
rect 159 1348 163 1352
rect 339 1347 343 1351
rect 359 1348 363 1352
rect 455 1347 456 1351
rect 456 1347 459 1351
rect 583 1348 587 1352
rect 675 1347 679 1351
rect 807 1348 811 1352
rect 903 1347 904 1351
rect 904 1347 907 1351
rect 1031 1348 1035 1352
rect 1127 1347 1128 1351
rect 1128 1347 1131 1351
rect 1935 1347 1939 1351
rect 1975 1347 1979 1351
rect 2127 1348 2131 1352
rect 2251 1347 2255 1351
rect 2271 1348 2275 1352
rect 2395 1347 2399 1351
rect 2415 1348 2419 1352
rect 2547 1347 2551 1351
rect 2567 1348 2571 1352
rect 2699 1347 2703 1351
rect 2719 1348 2723 1352
rect 2815 1347 2816 1351
rect 2816 1347 2819 1351
rect 2879 1348 2883 1352
rect 3039 1348 3043 1352
rect 3199 1348 3203 1352
rect 3799 1347 3803 1351
rect 2195 1315 2199 1319
rect 2887 1315 2891 1319
rect 3839 1297 3843 1301
rect 3887 1296 3891 1300
rect 3983 1295 3984 1299
rect 3984 1295 3987 1299
rect 4119 1296 4123 1300
rect 4219 1295 4220 1299
rect 4220 1295 4223 1299
rect 4391 1296 4395 1300
rect 4491 1295 4492 1299
rect 4492 1295 4495 1299
rect 4671 1296 4675 1300
rect 4767 1295 4768 1299
rect 4768 1295 4771 1299
rect 4967 1296 4971 1300
rect 5067 1295 5068 1299
rect 5068 1295 5071 1299
rect 5263 1296 5267 1300
rect 5355 1295 5359 1299
rect 5543 1296 5547 1300
rect 5635 1295 5639 1299
rect 5663 1297 5667 1301
rect 111 1289 115 1293
rect 159 1288 163 1292
rect 255 1287 256 1291
rect 256 1287 259 1291
rect 367 1288 371 1292
rect 463 1287 464 1291
rect 464 1287 467 1291
rect 607 1288 611 1292
rect 703 1287 704 1291
rect 704 1287 707 1291
rect 847 1288 851 1292
rect 971 1287 975 1291
rect 1087 1288 1091 1292
rect 1179 1287 1183 1291
rect 1935 1289 1939 1293
rect 1975 1285 1979 1289
rect 2023 1284 2027 1288
rect 2175 1284 2179 1288
rect 2311 1283 2315 1287
rect 2367 1284 2371 1288
rect 2467 1283 2468 1287
rect 2468 1283 2471 1287
rect 2575 1284 2579 1288
rect 2675 1283 2676 1287
rect 2676 1283 2679 1287
rect 2791 1284 2795 1288
rect 2887 1283 2888 1287
rect 2888 1283 2891 1287
rect 3015 1284 3019 1288
rect 3115 1283 3116 1287
rect 3116 1283 3119 1287
rect 3239 1284 3243 1288
rect 3335 1283 3336 1287
rect 3336 1283 3339 1287
rect 3471 1284 3475 1288
rect 3679 1284 3683 1288
rect 3791 1283 3795 1287
rect 3799 1285 3803 1289
rect 3839 1280 3843 1284
rect 3859 1281 3863 1285
rect 4091 1281 4095 1285
rect 4363 1281 4367 1285
rect 4643 1281 4647 1285
rect 4939 1281 4943 1285
rect 5235 1281 5239 1285
rect 5515 1281 5519 1285
rect 5663 1280 5667 1284
rect 111 1272 115 1276
rect 131 1273 135 1277
rect 339 1273 343 1277
rect 579 1273 583 1277
rect 819 1273 823 1277
rect 1059 1273 1063 1277
rect 1935 1272 1939 1276
rect 1975 1268 1979 1272
rect 1995 1269 1999 1273
rect 2147 1269 2151 1273
rect 2339 1269 2343 1273
rect 2547 1269 2551 1273
rect 2763 1269 2767 1273
rect 2987 1269 2991 1273
rect 3211 1269 3215 1273
rect 3443 1269 3447 1273
rect 3651 1269 3655 1273
rect 3799 1268 3803 1272
rect 3791 1231 3795 1235
rect 4135 1231 4139 1235
rect 4219 1231 4223 1235
rect 4491 1231 4495 1235
rect 251 1223 255 1227
rect 675 1223 679 1227
rect 903 1223 907 1227
rect 971 1223 975 1227
rect 5067 1231 5071 1235
rect 703 1215 707 1219
rect 1915 1219 1919 1223
rect 2311 1219 2315 1223
rect 2467 1219 2471 1223
rect 2675 1219 2679 1223
rect 3115 1219 3119 1223
rect 3583 1219 3587 1223
rect 5323 1223 5327 1227
rect 267 1179 271 1183
rect 371 1175 375 1179
rect 463 1179 467 1183
rect 611 1175 615 1179
rect 915 1179 919 1183
rect 1179 1187 1183 1191
rect 1335 1183 1339 1187
rect 1227 1175 1231 1179
rect 1371 1175 1375 1179
rect 1515 1175 1519 1179
rect 1659 1175 1663 1179
rect 1795 1175 1799 1179
rect 2819 1175 2823 1179
rect 2907 1175 2911 1179
rect 3335 1179 3339 1183
rect 3643 1179 3647 1183
rect 3671 1179 3675 1183
rect 4335 1183 4339 1187
rect 4219 1175 4223 1179
rect 4683 1179 4687 1183
rect 4767 1179 4771 1183
rect 4971 1175 4975 1179
rect 5355 1179 5359 1183
rect 5635 1179 5639 1183
rect 371 1151 375 1155
rect 727 1151 731 1155
rect 2819 1155 2823 1159
rect 3203 1155 3207 1159
rect 111 1128 115 1132
rect 131 1127 135 1131
rect 275 1127 279 1131
rect 443 1127 447 1131
rect 603 1127 607 1131
rect 763 1127 767 1131
rect 923 1127 927 1131
rect 1075 1127 1079 1131
rect 1219 1127 1223 1131
rect 1363 1127 1367 1131
rect 1507 1127 1511 1131
rect 1651 1127 1655 1131
rect 1787 1127 1791 1131
rect 1935 1128 1939 1132
rect 1975 1128 1979 1132
rect 2723 1127 2727 1131
rect 2899 1127 2903 1131
rect 3083 1127 3087 1131
rect 3275 1127 3279 1131
rect 3467 1127 3471 1131
rect 3651 1127 3655 1131
rect 3799 1128 3803 1132
rect 3839 1128 3843 1132
rect 4011 1127 4015 1131
rect 4211 1127 4215 1131
rect 4435 1127 4439 1131
rect 4691 1127 4695 1131
rect 4963 1127 4967 1131
rect 5251 1127 5255 1131
rect 5515 1127 5519 1131
rect 5663 1128 5667 1132
rect 915 1119 919 1123
rect 111 1111 115 1115
rect 159 1112 163 1116
rect 251 1111 255 1115
rect 303 1112 307 1116
rect 399 1111 400 1115
rect 400 1111 403 1115
rect 471 1112 475 1116
rect 611 1111 615 1115
rect 631 1112 635 1116
rect 727 1111 728 1115
rect 728 1111 731 1115
rect 791 1112 795 1116
rect 887 1111 888 1115
rect 888 1111 891 1115
rect 951 1112 955 1116
rect 3643 1119 3647 1123
rect 4683 1119 4687 1123
rect 1103 1112 1107 1116
rect 1227 1111 1231 1115
rect 1247 1112 1251 1116
rect 1371 1111 1375 1115
rect 1391 1112 1395 1116
rect 1515 1111 1519 1115
rect 1535 1112 1539 1116
rect 1659 1111 1663 1115
rect 1679 1112 1683 1116
rect 1795 1111 1799 1115
rect 1815 1112 1819 1116
rect 1915 1111 1916 1115
rect 1916 1111 1919 1115
rect 1935 1111 1939 1115
rect 1975 1111 1979 1115
rect 2751 1112 2755 1116
rect 2907 1111 2911 1115
rect 2927 1112 2931 1116
rect 3019 1111 3023 1115
rect 3111 1112 3115 1116
rect 3203 1111 3207 1115
rect 3303 1112 3307 1116
rect 3495 1112 3499 1116
rect 3587 1111 3591 1115
rect 3679 1112 3683 1116
rect 3799 1111 3803 1115
rect 3839 1111 3843 1115
rect 4039 1112 4043 1116
rect 4135 1111 4136 1115
rect 4136 1111 4139 1115
rect 4239 1112 4243 1116
rect 4335 1111 4336 1115
rect 4336 1111 4339 1115
rect 4463 1112 4467 1116
rect 4579 1111 4583 1115
rect 4719 1112 4723 1116
rect 4971 1111 4975 1115
rect 4991 1112 4995 1116
rect 5279 1112 5283 1116
rect 5375 1111 5376 1115
rect 5376 1111 5379 1115
rect 5543 1112 5547 1116
rect 5639 1111 5640 1115
rect 5640 1111 5643 1115
rect 5663 1111 5667 1115
rect 111 1045 115 1049
rect 175 1044 179 1048
rect 267 1043 271 1047
rect 415 1044 419 1048
rect 515 1043 516 1047
rect 516 1043 519 1047
rect 639 1044 643 1048
rect 735 1043 736 1047
rect 736 1043 739 1047
rect 855 1044 859 1048
rect 955 1043 956 1047
rect 956 1043 959 1047
rect 1055 1044 1059 1048
rect 1155 1043 1156 1047
rect 1156 1043 1159 1047
rect 1239 1044 1243 1048
rect 1335 1043 1336 1047
rect 1336 1043 1339 1047
rect 1423 1044 1427 1048
rect 1519 1043 1520 1047
rect 1520 1043 1523 1047
rect 1607 1044 1611 1048
rect 1703 1043 1704 1047
rect 1704 1043 1707 1047
rect 1791 1044 1795 1048
rect 1887 1043 1888 1047
rect 1888 1043 1891 1047
rect 1935 1045 1939 1049
rect 1975 1041 1979 1045
rect 2559 1040 2563 1044
rect 2651 1039 2655 1043
rect 2751 1040 2755 1044
rect 2843 1039 2847 1043
rect 2951 1040 2955 1044
rect 3051 1039 3052 1043
rect 3052 1039 3055 1043
rect 3151 1040 3155 1044
rect 3243 1039 3247 1043
rect 3359 1040 3363 1044
rect 3459 1039 3460 1043
rect 3460 1039 3463 1043
rect 3575 1040 3579 1044
rect 3671 1039 3672 1043
rect 3672 1039 3675 1043
rect 3799 1041 3803 1045
rect 3839 1041 3843 1045
rect 4095 1040 4099 1044
rect 4219 1039 4223 1043
rect 4391 1040 4395 1044
rect 4483 1039 4487 1043
rect 4687 1040 4691 1044
rect 4779 1039 4783 1043
rect 4975 1040 4979 1044
rect 5075 1039 5076 1043
rect 5076 1039 5079 1043
rect 5263 1040 5267 1044
rect 5355 1039 5359 1043
rect 5543 1040 5547 1044
rect 5663 1041 5667 1045
rect 111 1028 115 1032
rect 147 1029 151 1033
rect 387 1029 391 1033
rect 611 1029 615 1033
rect 827 1029 831 1033
rect 1027 1029 1031 1033
rect 1211 1029 1215 1033
rect 1395 1029 1399 1033
rect 1579 1029 1583 1033
rect 1763 1029 1767 1033
rect 1935 1028 1939 1032
rect 5647 1031 5651 1035
rect 1975 1024 1979 1028
rect 2531 1025 2535 1029
rect 2723 1025 2727 1029
rect 2923 1025 2927 1029
rect 3123 1025 3127 1029
rect 3331 1025 3335 1029
rect 3547 1025 3551 1029
rect 3799 1024 3803 1028
rect 3839 1024 3843 1028
rect 4067 1025 4071 1029
rect 4363 1025 4367 1029
rect 4659 1025 4663 1029
rect 4947 1025 4951 1029
rect 5235 1025 5239 1029
rect 5515 1025 5519 1029
rect 5663 1024 5667 1028
rect 1491 1007 1495 1011
rect 1703 1007 1707 1011
rect 2627 1007 2631 1011
rect 2843 1007 2847 1011
rect 319 979 323 983
rect 399 979 403 983
rect 515 979 519 983
rect 887 979 891 983
rect 955 979 959 983
rect 1491 979 1495 983
rect 1519 971 1523 975
rect 1907 979 1911 983
rect 1887 971 1891 975
rect 2627 975 2631 979
rect 3019 975 3023 979
rect 3051 975 3055 979
rect 3243 967 3247 971
rect 3459 975 3463 979
rect 4275 975 4279 979
rect 3531 967 3535 971
rect 4579 975 4583 979
rect 4779 967 4783 971
rect 5075 975 5079 979
rect 5639 975 5643 979
rect 5375 967 5379 971
rect 539 943 543 947
rect 2343 947 2347 951
rect 427 935 431 939
rect 735 939 739 943
rect 939 935 943 939
rect 1155 939 1159 943
rect 1523 935 1527 939
rect 1987 939 1991 943
rect 2315 939 2319 943
rect 2651 943 2655 947
rect 2715 939 2719 943
rect 3035 939 3039 943
rect 3179 939 3183 943
rect 3419 939 3423 943
rect 3983 939 3987 943
rect 4163 935 4167 939
rect 4483 939 4487 943
rect 4603 935 4607 939
rect 4819 935 4823 939
rect 5355 939 5359 943
rect 5599 939 5603 943
rect 5535 911 5539 915
rect 5591 911 5595 915
rect 3035 899 3039 903
rect 3207 899 3211 903
rect 111 888 115 892
rect 195 887 199 891
rect 419 887 423 891
rect 667 887 671 891
rect 931 887 935 891
rect 1219 887 1223 891
rect 1515 887 1519 891
rect 1787 887 1791 891
rect 1935 888 1939 892
rect 1975 892 1979 896
rect 1995 891 1999 895
rect 2219 891 2223 895
rect 2467 891 2471 895
rect 2707 891 2711 895
rect 2939 891 2943 895
rect 3171 891 3175 895
rect 3411 891 3415 895
rect 3799 892 3803 896
rect 3839 888 3843 892
rect 3931 887 3935 891
rect 1987 883 1991 887
rect 4155 887 4159 891
rect 4379 887 4383 891
rect 4595 887 4599 891
rect 4811 887 4815 891
rect 5027 887 5031 891
rect 5243 887 5247 891
rect 5467 887 5471 891
rect 5663 888 5667 892
rect 111 871 115 875
rect 223 872 227 876
rect 319 871 320 875
rect 320 871 323 875
rect 447 872 451 876
rect 539 871 543 875
rect 695 872 699 876
rect 939 871 943 875
rect 959 872 963 876
rect 1055 872 1056 875
rect 1056 872 1059 875
rect 1055 871 1059 872
rect 1247 872 1251 876
rect 1523 871 1527 875
rect 1543 872 1547 876
rect 1639 871 1640 875
rect 1640 871 1643 875
rect 1815 872 1819 876
rect 1907 871 1911 875
rect 1935 871 1939 875
rect 1975 875 1979 879
rect 2023 876 2027 880
rect 2247 876 2251 880
rect 2343 875 2344 879
rect 2344 875 2347 879
rect 2495 876 2499 880
rect 2715 875 2719 879
rect 2735 876 2739 880
rect 2831 875 2832 879
rect 2832 875 2835 879
rect 2967 876 2971 880
rect 3179 875 3183 879
rect 3199 876 3203 880
rect 3419 875 3423 879
rect 3439 876 3443 880
rect 3531 875 3535 879
rect 3799 875 3803 879
rect 3839 871 3843 875
rect 3959 872 3963 876
rect 4163 871 4167 875
rect 4183 872 4187 876
rect 4275 871 4279 875
rect 4407 872 4411 876
rect 4603 871 4607 875
rect 4623 872 4627 876
rect 4819 871 4823 875
rect 4839 872 4843 876
rect 4931 871 4935 875
rect 5055 872 5059 876
rect 5155 871 5156 875
rect 5156 871 5159 875
rect 5271 872 5275 876
rect 5495 872 5499 876
rect 5591 871 5592 875
rect 5592 871 5595 875
rect 5663 871 5667 875
rect 539 855 543 859
rect 1055 855 1059 859
rect 1975 817 1979 821
rect 2223 816 2227 820
rect 2315 815 2319 819
rect 2439 816 2443 820
rect 2535 815 2536 819
rect 2536 815 2539 819
rect 2663 816 2667 820
rect 2759 815 2760 819
rect 2760 815 2763 819
rect 2887 816 2891 820
rect 2979 815 2983 819
rect 3111 816 3115 820
rect 3207 815 3208 819
rect 3208 815 3211 819
rect 3335 816 3339 820
rect 3431 815 3432 819
rect 3432 815 3435 819
rect 3559 816 3563 820
rect 3651 815 3655 819
rect 3799 817 3803 821
rect 3839 813 3843 817
rect 3887 812 3891 816
rect 3983 811 3984 815
rect 3984 811 3987 815
rect 4111 812 4115 816
rect 4207 811 4208 815
rect 4208 811 4211 815
rect 4343 812 4347 816
rect 4575 812 4579 816
rect 4675 811 4676 815
rect 4676 811 4679 815
rect 4799 812 4803 816
rect 4891 811 4895 815
rect 5031 812 5035 816
rect 5123 811 5127 815
rect 5263 812 5267 816
rect 5355 811 5359 815
rect 5495 812 5499 816
rect 5592 811 5596 815
rect 5663 813 5667 817
rect 1975 800 1979 804
rect 2195 801 2199 805
rect 2411 801 2415 805
rect 2635 801 2639 805
rect 2859 801 2863 805
rect 3083 801 3087 805
rect 3307 801 3311 805
rect 3531 801 3535 805
rect 3799 800 3803 804
rect 3839 796 3843 800
rect 3859 797 3863 801
rect 4083 797 4087 801
rect 4315 797 4319 801
rect 4547 797 4551 801
rect 4771 797 4775 801
rect 5003 797 5007 801
rect 5235 797 5239 801
rect 5467 797 5471 801
rect 5663 796 5667 800
rect 111 789 115 793
rect 223 788 227 792
rect 427 787 431 791
rect 447 788 451 792
rect 547 787 548 791
rect 548 787 551 791
rect 663 788 667 792
rect 763 787 764 791
rect 764 787 767 791
rect 879 788 883 792
rect 975 787 976 791
rect 976 787 979 791
rect 1087 788 1091 792
rect 1179 787 1183 791
rect 1295 788 1299 792
rect 1387 787 1391 791
rect 1511 788 1515 792
rect 1607 787 1608 791
rect 1608 787 1611 791
rect 1935 789 1939 793
rect 3179 779 3183 783
rect 3431 779 3435 783
rect 3955 779 3959 783
rect 4207 779 4211 783
rect 111 772 115 776
rect 195 773 199 777
rect 419 773 423 777
rect 635 773 639 777
rect 851 773 855 777
rect 1059 773 1063 777
rect 1267 773 1271 777
rect 1483 773 1487 777
rect 1935 772 1939 776
rect 2535 743 2539 747
rect 2759 743 2763 747
rect 2831 751 2835 755
rect 3179 751 3183 755
rect 2979 743 2983 747
rect 3507 751 3511 755
rect 3651 743 3655 747
rect 3955 747 3959 751
rect 4203 747 4207 751
rect 4675 747 4679 751
rect 4931 739 4935 743
rect 5155 747 5159 751
rect 5647 747 5651 751
rect 5355 739 5359 743
rect 4651 731 4655 735
rect 5123 731 5127 735
rect 539 723 543 727
rect 547 723 551 727
rect 763 723 767 727
rect 563 715 567 719
rect 1387 715 1391 719
rect 1639 723 1643 727
rect 1607 715 1611 719
rect 3983 715 3987 719
rect 4679 719 4683 723
rect 4091 711 4095 715
rect 4651 711 4655 715
rect 4891 715 4895 719
rect 5011 711 5015 715
rect 5235 711 5239 715
rect 5639 715 5643 719
rect 3475 699 3479 703
rect 3775 703 3779 707
rect 255 683 259 687
rect 283 679 287 683
rect 451 679 455 683
rect 763 683 767 687
rect 911 683 915 687
rect 975 683 979 687
rect 1179 683 1183 687
rect 1227 679 1231 683
rect 1371 679 1375 683
rect 1515 679 1519 683
rect 1659 679 1663 683
rect 1795 679 1799 683
rect 3839 664 3843 668
rect 3475 659 3479 663
rect 3859 663 3863 667
rect 3639 659 3643 663
rect 4083 663 4087 667
rect 4323 663 4327 667
rect 4555 663 4559 667
rect 4779 663 4783 667
rect 5003 663 5007 667
rect 5227 663 5231 667
rect 5459 663 5463 667
rect 5663 664 5667 668
rect 1975 652 1979 656
rect 3379 651 3383 655
rect 3515 651 3519 655
rect 3651 651 3655 655
rect 3799 652 3803 656
rect 3839 647 3843 651
rect 3887 648 3891 652
rect 4091 647 4095 651
rect 4111 648 4115 652
rect 4203 647 4207 651
rect 4351 648 4355 652
rect 4447 647 4448 651
rect 4448 647 4451 651
rect 4583 648 4587 652
rect 4679 647 4680 651
rect 4680 647 4683 651
rect 4807 648 4811 652
rect 5011 647 5015 651
rect 5031 648 5035 652
rect 5235 647 5239 651
rect 5255 648 5259 652
rect 5347 647 5351 651
rect 5487 648 5491 652
rect 5583 647 5584 651
rect 5584 647 5587 651
rect 5663 647 5667 651
rect 111 632 115 636
rect 131 631 135 635
rect 275 631 279 635
rect 443 631 447 635
rect 611 631 615 635
rect 771 631 775 635
rect 923 631 927 635
rect 1075 631 1079 635
rect 1219 631 1223 635
rect 1363 631 1367 635
rect 1507 631 1511 635
rect 1651 631 1655 635
rect 1787 631 1791 635
rect 1935 632 1939 636
rect 1975 635 1979 639
rect 3407 636 3411 640
rect 3507 635 3508 639
rect 3508 635 3511 639
rect 3543 636 3547 640
rect 3639 635 3640 639
rect 3640 635 3643 639
rect 3679 636 3683 640
rect 3799 635 3803 639
rect 763 623 767 627
rect 111 615 115 619
rect 159 616 163 620
rect 283 615 287 619
rect 303 616 307 620
rect 451 615 455 619
rect 471 616 475 620
rect 563 615 567 619
rect 639 616 643 620
rect 735 615 736 619
rect 736 615 739 619
rect 799 616 803 620
rect 911 623 915 627
rect 951 616 955 620
rect 1103 616 1107 620
rect 1227 615 1231 619
rect 1247 616 1251 620
rect 1371 615 1375 619
rect 1391 616 1395 620
rect 1515 615 1519 619
rect 1535 616 1539 620
rect 1659 615 1663 619
rect 1679 616 1683 620
rect 1795 615 1799 619
rect 1815 616 1819 620
rect 1911 615 1912 619
rect 1912 615 1915 619
rect 1935 615 1939 619
rect 3839 581 3843 585
rect 3887 580 3891 584
rect 3983 579 3984 583
rect 3984 579 3987 583
rect 4143 580 4147 584
rect 4239 579 4240 583
rect 4240 579 4243 583
rect 4407 580 4411 584
rect 4503 579 4504 583
rect 4504 579 4507 583
rect 4647 580 4651 584
rect 4767 579 4771 583
rect 4879 580 4883 584
rect 4979 579 4980 583
rect 4980 579 4983 583
rect 5095 580 5099 584
rect 5195 579 5196 583
rect 5196 579 5199 583
rect 5311 580 5315 584
rect 5403 579 5407 583
rect 5527 580 5531 584
rect 5623 579 5624 583
rect 5624 579 5627 583
rect 5663 581 5667 585
rect 1975 569 1979 573
rect 3271 568 3275 572
rect 3371 567 3372 571
rect 3372 567 3375 571
rect 3407 568 3411 572
rect 3507 567 3508 571
rect 3508 567 3511 571
rect 3543 568 3547 572
rect 3643 567 3644 571
rect 3644 567 3647 571
rect 3679 568 3683 572
rect 3775 567 3776 571
rect 3776 567 3779 571
rect 3799 569 3803 573
rect 3839 564 3843 568
rect 3859 565 3863 569
rect 4115 565 4119 569
rect 4379 565 4383 569
rect 4619 565 4623 569
rect 4851 565 4855 569
rect 5067 565 5071 569
rect 5283 565 5287 569
rect 5499 565 5503 569
rect 5663 564 5667 568
rect 1975 552 1979 556
rect 3243 553 3247 557
rect 3379 553 3383 557
rect 3515 553 3519 557
rect 3651 553 3655 557
rect 3799 552 3803 556
rect 4715 551 4719 555
rect 5347 551 5351 555
rect 111 545 115 549
rect 159 544 163 548
rect 255 543 256 547
rect 256 543 259 547
rect 375 544 379 548
rect 467 543 471 547
rect 599 544 603 548
rect 699 543 700 547
rect 700 543 703 547
rect 807 544 811 548
rect 935 543 939 547
rect 999 544 1003 548
rect 1095 543 1096 547
rect 1096 543 1099 547
rect 1175 544 1179 548
rect 1275 543 1276 547
rect 1276 543 1279 547
rect 1343 544 1347 548
rect 1443 543 1444 547
rect 1444 543 1447 547
rect 1511 544 1515 548
rect 1611 543 1612 547
rect 1612 543 1615 547
rect 1671 544 1675 548
rect 1771 543 1772 547
rect 1772 543 1775 547
rect 1815 544 1819 548
rect 1927 543 1931 547
rect 1935 545 1939 549
rect 4779 543 4783 547
rect 5403 543 5407 547
rect 111 528 115 532
rect 131 529 135 533
rect 347 529 351 533
rect 571 529 575 533
rect 779 529 783 533
rect 971 529 975 533
rect 1147 529 1151 533
rect 1315 529 1319 533
rect 1483 529 1487 533
rect 1643 529 1647 533
rect 1787 529 1791 533
rect 1935 528 1939 532
rect 4015 515 4019 519
rect 4447 515 4451 519
rect 4715 515 4719 519
rect 4767 515 4771 519
rect 4979 515 4983 519
rect 5195 515 5199 519
rect 5583 515 5587 519
rect 3371 503 3375 507
rect 3507 503 3511 507
rect 3643 503 3647 507
rect 4239 507 4243 511
rect 3659 495 3663 499
rect 735 487 739 491
rect 699 479 703 483
rect 935 479 939 483
rect 467 471 471 475
rect 1275 479 1279 483
rect 1443 479 1447 483
rect 1611 479 1615 483
rect 1771 479 1775 483
rect 1911 471 1915 475
rect 4163 467 4167 471
rect 4295 467 4299 471
rect 4503 467 4507 471
rect 4779 467 4783 471
rect 4915 463 4919 467
rect 5131 463 5135 467
rect 5339 463 5343 467
rect 5523 463 5527 467
rect 599 447 603 451
rect 1095 447 1099 451
rect 1927 451 1931 455
rect 1339 443 1343 447
rect 2163 447 2167 451
rect 2355 447 2359 451
rect 2547 447 2551 451
rect 2747 447 2751 451
rect 3015 451 3019 455
rect 3139 447 3143 451
rect 3339 447 3343 451
rect 3539 447 3543 451
rect 3839 416 3843 420
rect 3891 415 3895 419
rect 4171 415 4175 419
rect 4435 415 4439 419
rect 4683 415 4687 419
rect 4907 415 4911 419
rect 5123 415 5127 419
rect 5331 415 5335 419
rect 5515 415 5519 419
rect 5663 416 5667 420
rect 4163 407 4167 411
rect 111 396 115 400
rect 195 395 199 399
rect 475 395 479 399
rect 755 395 759 399
rect 1043 395 1047 399
rect 1331 395 1335 399
rect 1935 396 1939 400
rect 1975 400 1979 404
rect 1995 399 1999 403
rect 2155 399 2159 403
rect 2347 399 2351 403
rect 2539 399 2543 403
rect 2739 399 2743 403
rect 2931 399 2935 403
rect 3131 399 3135 403
rect 3331 399 3335 403
rect 3531 399 3535 403
rect 3799 400 3803 404
rect 3839 399 3843 403
rect 3919 400 3923 404
rect 4015 399 4016 403
rect 4016 399 4019 403
rect 4199 400 4203 404
rect 4463 400 4467 404
rect 4555 399 4559 403
rect 4711 400 4715 404
rect 4915 399 4919 403
rect 4935 400 4939 404
rect 5131 399 5135 403
rect 5151 400 5155 404
rect 5339 399 5343 403
rect 5359 400 5363 404
rect 5523 399 5527 403
rect 5543 400 5547 404
rect 5639 399 5640 403
rect 5640 399 5643 403
rect 5663 399 5667 403
rect 111 379 115 383
rect 223 380 227 384
rect 503 380 507 384
rect 783 380 787 384
rect 879 379 880 383
rect 880 379 883 383
rect 1071 380 1075 384
rect 1339 379 1343 383
rect 1359 380 1363 384
rect 1935 379 1939 383
rect 1975 383 1979 387
rect 2023 384 2027 388
rect 2163 383 2167 387
rect 2183 384 2187 388
rect 2355 383 2359 387
rect 2375 384 2379 388
rect 2547 383 2551 387
rect 2567 384 2571 388
rect 2747 383 2751 387
rect 2767 384 2771 388
rect 2859 383 2863 387
rect 2959 384 2963 388
rect 3139 383 3143 387
rect 3159 384 3163 388
rect 3339 383 3343 387
rect 3359 384 3363 388
rect 3539 383 3543 387
rect 3559 384 3563 388
rect 3659 383 3660 387
rect 3660 383 3663 387
rect 3799 383 3803 387
rect 3839 337 3843 341
rect 4007 336 4011 340
rect 4135 335 4139 339
rect 4199 336 4203 340
rect 4295 335 4296 339
rect 4296 335 4299 339
rect 4423 336 4427 340
rect 4559 335 4563 339
rect 4679 336 4683 340
rect 4779 335 4780 339
rect 4780 335 4783 339
rect 4967 336 4971 340
rect 5067 335 5068 339
rect 5068 335 5071 339
rect 5263 336 5267 340
rect 5355 335 5359 339
rect 5543 336 5547 340
rect 5635 335 5639 339
rect 5663 337 5667 341
rect 111 321 115 325
rect 311 320 315 324
rect 431 319 435 323
rect 503 320 507 324
rect 599 319 600 323
rect 600 319 603 323
rect 695 320 699 324
rect 887 320 891 324
rect 1079 320 1083 324
rect 1175 319 1176 323
rect 1176 319 1179 323
rect 1935 321 1939 325
rect 3839 320 3843 324
rect 3979 321 3983 325
rect 4171 321 4175 325
rect 4395 321 4399 325
rect 4651 321 4655 325
rect 4939 321 4943 325
rect 5235 321 5239 325
rect 5515 321 5519 325
rect 5663 320 5667 324
rect 3015 315 3019 319
rect 111 304 115 308
rect 283 305 287 309
rect 475 305 479 309
rect 667 305 671 309
rect 859 305 863 309
rect 1051 305 1055 309
rect 1935 304 1939 308
rect 1975 301 1979 305
rect 2023 300 2027 304
rect 2123 299 2124 303
rect 2124 299 2127 303
rect 2159 300 2163 304
rect 2259 299 2260 303
rect 2260 299 2263 303
rect 2295 300 2299 304
rect 2395 299 2396 303
rect 2396 299 2399 303
rect 2431 300 2435 304
rect 2531 299 2532 303
rect 2532 299 2535 303
rect 2567 300 2571 304
rect 2667 299 2668 303
rect 2668 299 2671 303
rect 2703 300 2707 304
rect 2795 299 2799 303
rect 2839 300 2843 304
rect 2939 299 2940 303
rect 2940 299 2943 303
rect 2975 300 2979 304
rect 3075 299 3076 303
rect 3076 299 3079 303
rect 3111 300 3115 304
rect 3211 299 3212 303
rect 3212 299 3215 303
rect 3247 300 3251 304
rect 3347 299 3348 303
rect 3348 299 3351 303
rect 3383 300 3387 304
rect 3483 299 3484 303
rect 3484 299 3487 303
rect 3519 300 3523 304
rect 3799 301 3803 305
rect 1975 284 1979 288
rect 1995 285 1999 289
rect 2131 285 2135 289
rect 2267 285 2271 289
rect 2403 285 2407 289
rect 2539 285 2543 289
rect 2675 285 2679 289
rect 2811 285 2815 289
rect 2947 285 2951 289
rect 3083 285 3087 289
rect 3219 285 3223 289
rect 3355 285 3359 289
rect 3491 285 3495 289
rect 3799 284 3803 288
rect 2091 279 2095 283
rect 2859 279 2863 283
rect 4115 271 4119 275
rect 4135 271 4139 275
rect 4551 271 4555 275
rect 4559 271 4563 275
rect 4779 271 4783 275
rect 5067 271 5071 275
rect 5623 271 5627 275
rect 387 255 391 259
rect 431 255 435 259
rect 879 255 883 259
rect 1175 247 1179 251
rect 4723 251 4727 255
rect 5355 251 5359 255
rect 2091 235 2095 239
rect 2123 235 2127 239
rect 2259 235 2263 239
rect 2395 235 2399 239
rect 2531 235 2535 239
rect 2667 235 2671 239
rect 2907 235 2911 239
rect 2939 235 2943 239
rect 3075 235 3079 239
rect 3211 235 3215 239
rect 3347 235 3351 239
rect 3483 235 3487 239
rect 523 195 527 199
rect 275 183 279 187
rect 499 183 503 187
rect 667 187 671 191
rect 1207 195 1211 199
rect 4251 195 4255 199
rect 955 183 959 187
rect 1091 183 1095 187
rect 4003 183 4007 187
rect 4227 183 4231 187
rect 4395 187 4399 191
rect 4531 183 4535 187
rect 4723 187 4727 191
rect 4851 183 4855 187
rect 5075 183 5079 187
rect 5503 187 5507 191
rect 5635 187 5639 191
rect 2115 171 2119 175
rect 2139 167 2143 171
rect 2275 167 2279 171
rect 2411 167 2415 171
rect 2547 167 2551 171
rect 2683 167 2687 171
rect 2819 167 2823 171
rect 2955 167 2959 171
rect 3091 167 3095 171
rect 3227 167 3231 171
rect 3363 167 3367 171
rect 3499 167 3503 171
rect 3635 167 3639 171
rect 499 155 503 159
rect 659 155 663 159
rect 4227 155 4231 159
rect 4387 155 4391 159
rect 4531 151 4535 155
rect 5187 151 5191 155
rect 111 136 115 140
rect 131 135 135 139
rect 267 135 271 139
rect 403 135 407 139
rect 539 135 543 139
rect 675 135 679 139
rect 811 135 815 139
rect 947 135 951 139
rect 1083 135 1087 139
rect 1935 136 1939 140
rect 3839 136 3843 140
rect 3859 135 3863 139
rect 3995 135 3999 139
rect 4131 135 4135 139
rect 4267 135 4271 139
rect 4435 135 4439 139
rect 4627 135 4631 139
rect 4843 135 4847 139
rect 5067 135 5071 139
rect 5299 135 5303 139
rect 5515 135 5519 139
rect 5663 136 5667 140
rect 667 127 671 131
rect 4395 127 4399 131
rect 111 119 115 123
rect 159 120 163 124
rect 275 119 279 123
rect 295 120 299 124
rect 387 119 391 123
rect 431 120 435 124
rect 523 119 527 123
rect 567 120 571 124
rect 663 119 664 123
rect 664 119 667 123
rect 703 120 707 124
rect 5503 127 5507 131
rect 839 120 843 124
rect 955 119 959 123
rect 975 120 979 124
rect 1091 119 1095 123
rect 1111 120 1115 124
rect 1207 119 1208 123
rect 1208 119 1211 123
rect 1935 119 1939 123
rect 1975 120 1979 124
rect 1995 119 1999 123
rect 2131 119 2135 123
rect 2267 119 2271 123
rect 2403 119 2407 123
rect 2539 119 2543 123
rect 2675 119 2679 123
rect 2811 119 2815 123
rect 2947 119 2951 123
rect 3083 119 3087 123
rect 3219 119 3223 123
rect 3355 119 3359 123
rect 3491 119 3495 123
rect 3627 119 3631 123
rect 3799 120 3803 124
rect 3839 119 3843 123
rect 3887 120 3891 124
rect 4003 119 4007 123
rect 4023 120 4027 124
rect 4115 119 4119 123
rect 4159 120 4163 124
rect 4251 119 4255 123
rect 4295 120 4299 124
rect 4391 119 4392 123
rect 4392 119 4395 123
rect 4463 120 4467 124
rect 4655 120 4659 124
rect 4851 119 4855 123
rect 4871 120 4875 124
rect 5075 119 5079 123
rect 5095 120 5099 124
rect 5187 119 5191 123
rect 5327 120 5331 124
rect 5543 120 5547 124
rect 5663 119 5667 123
rect 1975 103 1979 107
rect 2023 104 2027 108
rect 2139 103 2143 107
rect 2159 104 2163 108
rect 2275 103 2279 107
rect 2295 104 2299 108
rect 2411 103 2415 107
rect 2431 104 2435 108
rect 2547 103 2551 107
rect 2567 104 2571 108
rect 2683 103 2687 107
rect 2703 104 2707 108
rect 2819 103 2823 107
rect 2839 104 2843 108
rect 2955 103 2959 107
rect 2975 104 2979 108
rect 3091 103 3095 107
rect 3111 104 3115 108
rect 3227 103 3231 107
rect 3247 104 3251 108
rect 3363 103 3367 107
rect 3383 104 3387 108
rect 3499 103 3503 107
rect 3519 104 3523 108
rect 3635 103 3639 107
rect 3655 104 3659 108
rect 3751 103 3752 107
rect 3752 103 3755 107
rect 3799 103 3803 107
<< m3 >>
rect 111 5758 115 5759
rect 111 5753 115 5754
rect 131 5758 135 5759
rect 131 5753 135 5754
rect 371 5758 375 5759
rect 371 5753 375 5754
rect 635 5758 639 5759
rect 635 5753 639 5754
rect 907 5758 911 5759
rect 907 5753 911 5754
rect 1179 5758 1183 5759
rect 1179 5753 1183 5754
rect 1451 5758 1455 5759
rect 1451 5753 1455 5754
rect 1723 5758 1727 5759
rect 1723 5753 1727 5754
rect 1935 5758 1939 5759
rect 1935 5753 1939 5754
rect 112 5693 114 5753
rect 110 5692 116 5693
rect 132 5692 134 5753
rect 372 5692 374 5753
rect 378 5739 384 5740
rect 378 5735 379 5739
rect 383 5735 384 5739
rect 378 5734 384 5735
rect 110 5688 111 5692
rect 115 5688 116 5692
rect 110 5687 116 5688
rect 130 5691 136 5692
rect 130 5687 131 5691
rect 135 5687 136 5691
rect 130 5686 136 5687
rect 370 5691 376 5692
rect 370 5687 371 5691
rect 375 5687 376 5691
rect 370 5686 376 5687
rect 158 5676 164 5677
rect 380 5676 382 5734
rect 636 5692 638 5753
rect 642 5739 648 5740
rect 642 5735 643 5739
rect 647 5735 648 5739
rect 642 5734 648 5735
rect 634 5691 640 5692
rect 634 5687 635 5691
rect 639 5687 640 5691
rect 634 5686 640 5687
rect 398 5676 404 5677
rect 644 5676 646 5734
rect 908 5692 910 5753
rect 914 5739 920 5740
rect 914 5735 915 5739
rect 919 5735 920 5739
rect 914 5734 920 5735
rect 906 5691 912 5692
rect 906 5687 907 5691
rect 911 5687 912 5691
rect 906 5686 912 5687
rect 662 5676 668 5677
rect 916 5676 918 5734
rect 1180 5692 1182 5753
rect 1452 5692 1454 5753
rect 1678 5747 1684 5748
rect 1678 5743 1679 5747
rect 1683 5743 1684 5747
rect 1678 5742 1684 5743
rect 1458 5739 1464 5740
rect 1458 5735 1459 5739
rect 1463 5735 1464 5739
rect 1458 5734 1464 5735
rect 1178 5691 1184 5692
rect 1178 5687 1179 5691
rect 1183 5687 1184 5691
rect 1178 5686 1184 5687
rect 1450 5691 1456 5692
rect 1450 5687 1451 5691
rect 1455 5687 1456 5691
rect 1450 5686 1456 5687
rect 934 5676 940 5677
rect 1206 5676 1212 5677
rect 1460 5676 1462 5734
rect 1478 5676 1484 5677
rect 110 5675 116 5676
rect 110 5671 111 5675
rect 115 5671 116 5675
rect 158 5672 159 5676
rect 163 5672 164 5676
rect 158 5671 164 5672
rect 378 5675 384 5676
rect 378 5671 379 5675
rect 383 5671 384 5675
rect 398 5672 399 5676
rect 403 5672 404 5676
rect 398 5671 404 5672
rect 642 5675 648 5676
rect 642 5671 643 5675
rect 647 5671 648 5675
rect 662 5672 663 5676
rect 667 5672 668 5676
rect 662 5671 668 5672
rect 914 5675 920 5676
rect 914 5671 915 5675
rect 919 5671 920 5675
rect 934 5672 935 5676
rect 939 5672 940 5676
rect 934 5671 940 5672
rect 1030 5675 1036 5676
rect 1030 5671 1031 5675
rect 1035 5671 1036 5675
rect 1206 5672 1207 5676
rect 1211 5672 1212 5676
rect 1206 5671 1212 5672
rect 1458 5675 1464 5676
rect 1458 5671 1459 5675
rect 1463 5671 1464 5675
rect 1478 5672 1479 5676
rect 1483 5672 1484 5676
rect 1478 5671 1484 5672
rect 110 5670 116 5671
rect 112 5647 114 5670
rect 160 5647 162 5671
rect 378 5670 384 5671
rect 400 5647 402 5671
rect 642 5670 648 5671
rect 664 5647 666 5671
rect 914 5670 920 5671
rect 936 5647 938 5671
rect 1030 5670 1036 5671
rect 111 5646 115 5647
rect 111 5641 115 5642
rect 159 5646 163 5647
rect 159 5641 163 5642
rect 399 5646 403 5647
rect 399 5641 403 5642
rect 455 5646 459 5647
rect 455 5641 459 5642
rect 647 5646 651 5647
rect 647 5641 651 5642
rect 663 5646 667 5647
rect 663 5641 667 5642
rect 855 5646 859 5647
rect 855 5641 859 5642
rect 935 5646 939 5647
rect 935 5641 939 5642
rect 112 5618 114 5641
rect 110 5617 116 5618
rect 456 5617 458 5641
rect 648 5617 650 5641
rect 856 5617 858 5641
rect 110 5613 111 5617
rect 115 5613 116 5617
rect 110 5612 116 5613
rect 454 5616 460 5617
rect 454 5612 455 5616
rect 459 5612 460 5616
rect 454 5611 460 5612
rect 646 5616 652 5617
rect 854 5616 860 5617
rect 646 5612 647 5616
rect 651 5612 652 5616
rect 646 5611 652 5612
rect 746 5615 752 5616
rect 746 5611 747 5615
rect 751 5611 752 5615
rect 854 5612 855 5616
rect 859 5612 860 5616
rect 854 5611 860 5612
rect 966 5615 972 5616
rect 966 5611 967 5615
rect 971 5611 972 5615
rect 746 5610 752 5611
rect 966 5610 972 5611
rect 426 5601 432 5602
rect 110 5600 116 5601
rect 110 5596 111 5600
rect 115 5596 116 5600
rect 426 5597 427 5601
rect 431 5597 432 5601
rect 426 5596 432 5597
rect 618 5601 624 5602
rect 618 5597 619 5601
rect 623 5597 624 5601
rect 618 5596 624 5597
rect 110 5595 116 5596
rect 112 5535 114 5595
rect 428 5535 430 5596
rect 620 5535 622 5596
rect 748 5552 750 5610
rect 826 5601 832 5602
rect 826 5597 827 5601
rect 831 5597 832 5601
rect 826 5596 832 5597
rect 746 5551 752 5552
rect 746 5547 747 5551
rect 751 5547 752 5551
rect 746 5546 752 5547
rect 828 5535 830 5596
rect 883 5564 887 5565
rect 883 5559 887 5560
rect 111 5534 115 5535
rect 111 5529 115 5530
rect 427 5534 431 5535
rect 427 5529 431 5530
rect 619 5534 623 5535
rect 619 5529 623 5530
rect 787 5534 791 5535
rect 787 5529 791 5530
rect 827 5534 831 5535
rect 827 5529 831 5530
rect 112 5469 114 5529
rect 110 5468 116 5469
rect 788 5468 790 5529
rect 884 5520 886 5559
rect 968 5552 970 5610
rect 966 5551 972 5552
rect 966 5547 967 5551
rect 971 5547 972 5551
rect 966 5546 972 5547
rect 1032 5544 1034 5670
rect 1208 5647 1210 5671
rect 1458 5670 1464 5671
rect 1480 5647 1482 5671
rect 1087 5646 1091 5647
rect 1087 5641 1091 5642
rect 1207 5646 1211 5647
rect 1207 5641 1211 5642
rect 1327 5646 1331 5647
rect 1327 5641 1331 5642
rect 1479 5646 1483 5647
rect 1479 5641 1483 5642
rect 1583 5646 1587 5647
rect 1583 5641 1587 5642
rect 1088 5617 1090 5641
rect 1328 5617 1330 5641
rect 1584 5617 1586 5641
rect 1086 5616 1092 5617
rect 1326 5616 1332 5617
rect 1086 5612 1087 5616
rect 1091 5612 1092 5616
rect 1086 5611 1092 5612
rect 1178 5615 1184 5616
rect 1178 5611 1179 5615
rect 1183 5611 1184 5615
rect 1326 5612 1327 5616
rect 1331 5612 1332 5616
rect 1326 5611 1332 5612
rect 1582 5616 1588 5617
rect 1680 5616 1682 5742
rect 1724 5692 1726 5753
rect 1730 5739 1736 5740
rect 1730 5735 1731 5739
rect 1735 5735 1736 5739
rect 1730 5734 1736 5735
rect 1722 5691 1728 5692
rect 1722 5687 1723 5691
rect 1727 5687 1728 5691
rect 1722 5686 1728 5687
rect 1732 5676 1734 5734
rect 1936 5693 1938 5753
rect 1975 5722 1979 5723
rect 1975 5717 1979 5718
rect 2511 5722 2515 5723
rect 2511 5717 2515 5718
rect 2663 5722 2667 5723
rect 2663 5717 2667 5718
rect 2815 5722 2819 5723
rect 2815 5717 2819 5718
rect 2975 5722 2979 5723
rect 2975 5717 2979 5718
rect 3143 5722 3147 5723
rect 3143 5717 3147 5718
rect 3319 5722 3323 5723
rect 3319 5717 3323 5718
rect 3495 5722 3499 5723
rect 3495 5717 3499 5718
rect 3799 5722 3803 5723
rect 3799 5717 3803 5718
rect 1976 5694 1978 5717
rect 1974 5693 1980 5694
rect 2512 5693 2514 5717
rect 2664 5693 2666 5717
rect 2816 5693 2818 5717
rect 2976 5693 2978 5717
rect 3144 5693 3146 5717
rect 3320 5693 3322 5717
rect 3496 5693 3498 5717
rect 3800 5694 3802 5717
rect 3798 5693 3804 5694
rect 1934 5692 1940 5693
rect 1934 5688 1935 5692
rect 1939 5688 1940 5692
rect 1974 5689 1975 5693
rect 1979 5689 1980 5693
rect 1974 5688 1980 5689
rect 2510 5692 2516 5693
rect 2510 5688 2511 5692
rect 2515 5688 2516 5692
rect 1934 5687 1940 5688
rect 2510 5687 2516 5688
rect 2662 5692 2668 5693
rect 2814 5692 2820 5693
rect 2974 5692 2980 5693
rect 3142 5692 3148 5693
rect 3318 5692 3324 5693
rect 3494 5692 3500 5693
rect 2662 5688 2663 5692
rect 2667 5688 2668 5692
rect 2662 5687 2668 5688
rect 2754 5691 2760 5692
rect 2754 5687 2755 5691
rect 2759 5687 2760 5691
rect 2814 5688 2815 5692
rect 2819 5688 2820 5692
rect 2814 5687 2820 5688
rect 2906 5691 2912 5692
rect 2906 5687 2907 5691
rect 2911 5687 2912 5691
rect 2974 5688 2975 5692
rect 2979 5688 2980 5692
rect 2974 5687 2980 5688
rect 3070 5691 3076 5692
rect 3070 5687 3071 5691
rect 3075 5687 3076 5691
rect 3142 5688 3143 5692
rect 3147 5688 3148 5692
rect 3142 5687 3148 5688
rect 3238 5691 3244 5692
rect 3238 5687 3239 5691
rect 3243 5687 3244 5691
rect 3318 5688 3319 5692
rect 3323 5688 3324 5692
rect 3318 5687 3324 5688
rect 3414 5691 3420 5692
rect 3414 5687 3415 5691
rect 3419 5687 3420 5691
rect 3494 5688 3495 5692
rect 3499 5688 3500 5692
rect 3494 5687 3500 5688
rect 3590 5691 3596 5692
rect 3590 5687 3591 5691
rect 3595 5687 3596 5691
rect 3798 5689 3799 5693
rect 3803 5689 3804 5693
rect 3798 5688 3804 5689
rect 2754 5686 2760 5687
rect 2906 5686 2912 5687
rect 3070 5686 3076 5687
rect 3238 5686 3244 5687
rect 3414 5686 3420 5687
rect 3590 5686 3596 5687
rect 2482 5677 2488 5678
rect 1750 5676 1756 5677
rect 1974 5676 1980 5677
rect 1730 5675 1736 5676
rect 1730 5671 1731 5675
rect 1735 5671 1736 5675
rect 1750 5672 1751 5676
rect 1755 5672 1756 5676
rect 1750 5671 1756 5672
rect 1846 5675 1852 5676
rect 1846 5671 1847 5675
rect 1851 5671 1852 5675
rect 1730 5670 1736 5671
rect 1752 5647 1754 5671
rect 1846 5670 1852 5671
rect 1934 5675 1940 5676
rect 1934 5671 1935 5675
rect 1939 5671 1940 5675
rect 1974 5672 1975 5676
rect 1979 5672 1980 5676
rect 2482 5673 2483 5677
rect 2487 5673 2488 5677
rect 2482 5672 2488 5673
rect 2634 5677 2640 5678
rect 2634 5673 2635 5677
rect 2639 5673 2640 5677
rect 2634 5672 2640 5673
rect 1974 5671 1980 5672
rect 1934 5670 1940 5671
rect 1751 5646 1755 5647
rect 1751 5641 1755 5642
rect 1815 5646 1819 5647
rect 1815 5641 1819 5642
rect 1816 5617 1818 5641
rect 1814 5616 1820 5617
rect 1582 5612 1583 5616
rect 1587 5612 1588 5616
rect 1582 5611 1588 5612
rect 1678 5615 1684 5616
rect 1678 5611 1679 5615
rect 1683 5611 1684 5615
rect 1814 5612 1815 5616
rect 1819 5612 1820 5616
rect 1814 5611 1820 5612
rect 1178 5610 1184 5611
rect 1678 5610 1684 5611
rect 1058 5601 1064 5602
rect 1058 5597 1059 5601
rect 1063 5597 1064 5601
rect 1058 5596 1064 5597
rect 1030 5543 1036 5544
rect 1030 5539 1031 5543
rect 1035 5539 1036 5543
rect 1030 5538 1036 5539
rect 1060 5535 1062 5596
rect 1180 5565 1182 5610
rect 1298 5601 1304 5602
rect 1298 5597 1299 5601
rect 1303 5597 1304 5601
rect 1298 5596 1304 5597
rect 1554 5601 1560 5602
rect 1554 5597 1555 5601
rect 1559 5597 1560 5601
rect 1554 5596 1560 5597
rect 1786 5601 1792 5602
rect 1786 5597 1787 5601
rect 1791 5597 1792 5601
rect 1786 5596 1792 5597
rect 1179 5564 1183 5565
rect 1179 5559 1183 5560
rect 1300 5535 1302 5596
rect 1318 5551 1324 5552
rect 1318 5547 1319 5551
rect 1323 5547 1324 5551
rect 1318 5546 1324 5547
rect 923 5534 927 5535
rect 923 5529 927 5530
rect 1059 5534 1063 5535
rect 1059 5529 1063 5530
rect 1195 5534 1199 5535
rect 1195 5529 1199 5530
rect 1299 5534 1303 5535
rect 1299 5529 1303 5530
rect 882 5519 888 5520
rect 882 5515 883 5519
rect 887 5515 888 5519
rect 882 5514 888 5515
rect 924 5468 926 5529
rect 930 5515 936 5516
rect 930 5511 931 5515
rect 935 5511 936 5515
rect 930 5510 936 5511
rect 110 5464 111 5468
rect 115 5464 116 5468
rect 110 5463 116 5464
rect 786 5467 792 5468
rect 786 5463 787 5467
rect 791 5463 792 5467
rect 786 5462 792 5463
rect 922 5467 928 5468
rect 922 5463 923 5467
rect 927 5463 928 5467
rect 922 5462 928 5463
rect 814 5452 820 5453
rect 932 5452 934 5510
rect 1060 5468 1062 5529
rect 1066 5515 1072 5516
rect 1066 5511 1067 5515
rect 1071 5511 1072 5515
rect 1066 5510 1072 5511
rect 1058 5467 1064 5468
rect 1058 5463 1059 5467
rect 1063 5463 1064 5467
rect 1058 5462 1064 5463
rect 950 5452 956 5453
rect 1068 5452 1070 5510
rect 1196 5468 1198 5529
rect 1202 5515 1208 5516
rect 1202 5511 1203 5515
rect 1207 5511 1208 5515
rect 1202 5510 1208 5511
rect 1194 5467 1200 5468
rect 1194 5463 1195 5467
rect 1199 5463 1200 5467
rect 1194 5462 1200 5463
rect 1086 5452 1092 5453
rect 1204 5452 1206 5510
rect 1222 5452 1228 5453
rect 1320 5452 1322 5546
rect 1556 5535 1558 5596
rect 1788 5535 1790 5596
rect 1848 5552 1850 5670
rect 1936 5647 1938 5670
rect 1935 5646 1939 5647
rect 1935 5641 1939 5642
rect 1936 5618 1938 5641
rect 1934 5617 1940 5618
rect 1926 5615 1932 5616
rect 1926 5611 1927 5615
rect 1931 5611 1932 5615
rect 1934 5613 1935 5617
rect 1939 5613 1940 5617
rect 1934 5612 1940 5613
rect 1926 5610 1932 5611
rect 1928 5588 1930 5610
rect 1976 5603 1978 5671
rect 2484 5603 2486 5672
rect 2636 5603 2638 5672
rect 1975 5602 1979 5603
rect 1934 5600 1940 5601
rect 1934 5596 1935 5600
rect 1939 5596 1940 5600
rect 1975 5597 1979 5598
rect 1995 5602 1999 5603
rect 1995 5597 1999 5598
rect 2203 5602 2207 5603
rect 2203 5597 2207 5598
rect 2435 5602 2439 5603
rect 2435 5597 2439 5598
rect 2483 5602 2487 5603
rect 2483 5597 2487 5598
rect 2635 5602 2639 5603
rect 2635 5597 2639 5598
rect 2659 5602 2663 5603
rect 2659 5597 2663 5598
rect 1934 5595 1940 5596
rect 1926 5587 1932 5588
rect 1926 5583 1927 5587
rect 1931 5583 1932 5587
rect 1926 5582 1932 5583
rect 1846 5551 1852 5552
rect 1846 5547 1847 5551
rect 1851 5547 1852 5551
rect 1846 5546 1852 5547
rect 1936 5535 1938 5595
rect 1976 5537 1978 5597
rect 1974 5536 1980 5537
rect 1996 5536 1998 5597
rect 2204 5536 2206 5597
rect 2436 5536 2438 5597
rect 2442 5583 2448 5584
rect 2442 5579 2443 5583
rect 2447 5579 2448 5583
rect 2442 5578 2448 5579
rect 1331 5534 1335 5535
rect 1331 5529 1335 5530
rect 1555 5534 1559 5535
rect 1555 5529 1559 5530
rect 1787 5534 1791 5535
rect 1787 5529 1791 5530
rect 1935 5534 1939 5535
rect 1974 5532 1975 5536
rect 1979 5532 1980 5536
rect 1974 5531 1980 5532
rect 1994 5535 2000 5536
rect 1994 5531 1995 5535
rect 1999 5531 2000 5535
rect 1994 5530 2000 5531
rect 2202 5535 2208 5536
rect 2202 5531 2203 5535
rect 2207 5531 2208 5535
rect 2202 5530 2208 5531
rect 2434 5535 2440 5536
rect 2434 5531 2435 5535
rect 2439 5531 2440 5535
rect 2434 5530 2440 5531
rect 1935 5529 1939 5530
rect 1332 5468 1334 5529
rect 1426 5515 1432 5516
rect 1426 5511 1427 5515
rect 1431 5511 1432 5515
rect 1426 5510 1432 5511
rect 1330 5467 1336 5468
rect 1330 5463 1331 5467
rect 1335 5463 1336 5467
rect 1330 5462 1336 5463
rect 1358 5452 1364 5453
rect 110 5451 116 5452
rect 110 5447 111 5451
rect 115 5447 116 5451
rect 814 5448 815 5452
rect 819 5448 820 5452
rect 814 5447 820 5448
rect 930 5451 936 5452
rect 930 5447 931 5451
rect 935 5447 936 5451
rect 950 5448 951 5452
rect 955 5448 956 5452
rect 950 5447 956 5448
rect 1066 5451 1072 5452
rect 1066 5447 1067 5451
rect 1071 5447 1072 5451
rect 1086 5448 1087 5452
rect 1091 5448 1092 5452
rect 1086 5447 1092 5448
rect 1202 5451 1208 5452
rect 1202 5447 1203 5451
rect 1207 5447 1208 5451
rect 1222 5448 1223 5452
rect 1227 5448 1228 5452
rect 1222 5447 1228 5448
rect 1318 5451 1324 5452
rect 1318 5447 1319 5451
rect 1323 5447 1324 5451
rect 1358 5448 1359 5452
rect 1363 5448 1364 5452
rect 1358 5447 1364 5448
rect 110 5446 116 5447
rect 112 5403 114 5446
rect 816 5403 818 5447
rect 930 5446 936 5447
rect 952 5403 954 5447
rect 1066 5446 1072 5447
rect 1088 5403 1090 5447
rect 1202 5446 1208 5447
rect 1224 5403 1226 5447
rect 1318 5446 1324 5447
rect 1250 5419 1256 5420
rect 1250 5415 1251 5419
rect 1255 5415 1256 5419
rect 1250 5414 1256 5415
rect 111 5402 115 5403
rect 111 5397 115 5398
rect 815 5402 819 5403
rect 815 5397 819 5398
rect 903 5402 907 5403
rect 903 5397 907 5398
rect 951 5402 955 5403
rect 951 5397 955 5398
rect 1039 5402 1043 5403
rect 1039 5397 1043 5398
rect 1087 5402 1091 5403
rect 1087 5397 1091 5398
rect 1183 5402 1187 5403
rect 1183 5397 1187 5398
rect 1223 5402 1227 5403
rect 1223 5397 1227 5398
rect 112 5374 114 5397
rect 110 5373 116 5374
rect 904 5373 906 5397
rect 1040 5373 1042 5397
rect 1184 5373 1186 5397
rect 110 5369 111 5373
rect 115 5369 116 5373
rect 110 5368 116 5369
rect 902 5372 908 5373
rect 1038 5372 1044 5373
rect 1182 5372 1188 5373
rect 902 5368 903 5372
rect 907 5368 908 5372
rect 902 5367 908 5368
rect 1002 5371 1008 5372
rect 1002 5367 1003 5371
rect 1007 5367 1008 5371
rect 1038 5368 1039 5372
rect 1043 5368 1044 5372
rect 1038 5367 1044 5368
rect 1134 5371 1140 5372
rect 1134 5367 1135 5371
rect 1139 5367 1140 5371
rect 1182 5368 1183 5372
rect 1187 5368 1188 5372
rect 1182 5367 1188 5368
rect 1002 5366 1008 5367
rect 1134 5366 1140 5367
rect 874 5357 880 5358
rect 110 5356 116 5357
rect 110 5352 111 5356
rect 115 5352 116 5356
rect 874 5353 875 5357
rect 879 5353 880 5357
rect 874 5352 880 5353
rect 110 5351 116 5352
rect 112 5287 114 5351
rect 876 5287 878 5352
rect 1004 5308 1006 5366
rect 1010 5357 1016 5358
rect 1010 5353 1011 5357
rect 1015 5353 1016 5357
rect 1010 5352 1016 5353
rect 1002 5307 1008 5308
rect 1002 5303 1003 5307
rect 1007 5303 1008 5307
rect 1002 5302 1008 5303
rect 1012 5287 1014 5352
rect 111 5286 115 5287
rect 111 5281 115 5282
rect 587 5286 591 5287
rect 587 5281 591 5282
rect 739 5286 743 5287
rect 739 5281 743 5282
rect 875 5286 879 5287
rect 875 5281 879 5282
rect 899 5286 903 5287
rect 899 5281 903 5282
rect 1011 5286 1015 5287
rect 1011 5281 1015 5282
rect 1067 5286 1071 5287
rect 1067 5281 1071 5282
rect 112 5221 114 5281
rect 110 5220 116 5221
rect 588 5220 590 5281
rect 740 5220 742 5281
rect 862 5275 868 5276
rect 862 5271 863 5275
rect 867 5271 868 5275
rect 862 5270 868 5271
rect 110 5216 111 5220
rect 115 5216 116 5220
rect 110 5215 116 5216
rect 586 5219 592 5220
rect 586 5215 587 5219
rect 591 5215 592 5219
rect 586 5214 592 5215
rect 738 5219 744 5220
rect 738 5215 739 5219
rect 743 5215 744 5219
rect 738 5214 744 5215
rect 614 5204 620 5205
rect 766 5204 772 5205
rect 864 5204 866 5270
rect 900 5220 902 5281
rect 994 5267 1000 5268
rect 994 5263 995 5267
rect 999 5263 1000 5267
rect 994 5262 1000 5263
rect 996 5240 998 5262
rect 994 5239 1000 5240
rect 994 5235 995 5239
rect 999 5235 1000 5239
rect 994 5234 1000 5235
rect 1068 5220 1070 5281
rect 1136 5272 1138 5366
rect 1154 5357 1160 5358
rect 1154 5353 1155 5357
rect 1159 5353 1160 5357
rect 1154 5352 1160 5353
rect 1156 5287 1158 5352
rect 1252 5308 1254 5414
rect 1360 5403 1362 5447
rect 1335 5402 1339 5403
rect 1335 5397 1339 5398
rect 1359 5402 1363 5403
rect 1359 5397 1363 5398
rect 1336 5373 1338 5397
rect 1334 5372 1340 5373
rect 1428 5372 1430 5510
rect 1936 5469 1938 5529
rect 2022 5520 2028 5521
rect 2230 5520 2236 5521
rect 2444 5520 2446 5578
rect 2660 5536 2662 5597
rect 2756 5588 2758 5686
rect 2786 5677 2792 5678
rect 2786 5673 2787 5677
rect 2791 5673 2792 5677
rect 2786 5672 2792 5673
rect 2788 5603 2790 5672
rect 2908 5620 2910 5686
rect 2946 5677 2952 5678
rect 2946 5673 2947 5677
rect 2951 5673 2952 5677
rect 2946 5672 2952 5673
rect 2906 5619 2912 5620
rect 2906 5615 2907 5619
rect 2911 5615 2912 5619
rect 2906 5614 2912 5615
rect 2948 5603 2950 5672
rect 3072 5620 3074 5686
rect 3114 5677 3120 5678
rect 3114 5673 3115 5677
rect 3119 5673 3120 5677
rect 3114 5672 3120 5673
rect 3070 5619 3076 5620
rect 3070 5615 3071 5619
rect 3075 5615 3076 5619
rect 3070 5614 3076 5615
rect 3116 5603 3118 5672
rect 3210 5671 3216 5672
rect 3210 5667 3211 5671
rect 3215 5667 3216 5671
rect 3210 5666 3216 5667
rect 3212 5628 3214 5666
rect 3210 5627 3216 5628
rect 3210 5623 3211 5627
rect 3215 5623 3216 5627
rect 3210 5622 3216 5623
rect 3240 5620 3242 5686
rect 3290 5677 3296 5678
rect 3290 5673 3291 5677
rect 3295 5673 3296 5677
rect 3290 5672 3296 5673
rect 3416 5672 3418 5686
rect 3466 5677 3472 5678
rect 3466 5673 3467 5677
rect 3471 5673 3472 5677
rect 3466 5672 3472 5673
rect 3238 5619 3244 5620
rect 3238 5615 3239 5619
rect 3243 5615 3244 5619
rect 3238 5614 3244 5615
rect 3292 5603 3294 5672
rect 3414 5671 3420 5672
rect 3414 5667 3415 5671
rect 3419 5667 3420 5671
rect 3414 5666 3420 5667
rect 3468 5603 3470 5672
rect 3592 5620 3594 5686
rect 3798 5676 3804 5677
rect 3798 5672 3799 5676
rect 3803 5672 3804 5676
rect 3798 5671 3804 5672
rect 3839 5674 3843 5675
rect 3774 5627 3780 5628
rect 3774 5623 3775 5627
rect 3779 5623 3780 5627
rect 3774 5622 3780 5623
rect 3590 5619 3596 5620
rect 3590 5615 3591 5619
rect 3595 5615 3596 5619
rect 3590 5614 3596 5615
rect 2787 5602 2791 5603
rect 2787 5597 2791 5598
rect 2867 5602 2871 5603
rect 2867 5597 2871 5598
rect 2947 5602 2951 5603
rect 2947 5597 2951 5598
rect 3075 5602 3079 5603
rect 3075 5597 3079 5598
rect 3115 5602 3119 5603
rect 3115 5597 3119 5598
rect 3275 5602 3279 5603
rect 3275 5597 3279 5598
rect 3291 5602 3295 5603
rect 3291 5597 3295 5598
rect 3467 5602 3471 5603
rect 3467 5597 3471 5598
rect 3475 5602 3479 5603
rect 3475 5597 3479 5598
rect 3651 5602 3655 5603
rect 3651 5597 3655 5598
rect 2778 5595 2784 5596
rect 2778 5591 2779 5595
rect 2783 5591 2784 5595
rect 2778 5590 2784 5591
rect 2754 5587 2760 5588
rect 2754 5583 2755 5587
rect 2759 5583 2760 5587
rect 2754 5582 2760 5583
rect 2658 5535 2664 5536
rect 2658 5531 2659 5535
rect 2663 5531 2664 5535
rect 2658 5530 2664 5531
rect 2462 5520 2468 5521
rect 2686 5520 2692 5521
rect 2780 5520 2782 5590
rect 2868 5536 2870 5597
rect 3076 5536 3078 5597
rect 3082 5583 3088 5584
rect 3082 5579 3083 5583
rect 3087 5579 3088 5583
rect 3082 5578 3088 5579
rect 2866 5535 2872 5536
rect 2866 5531 2867 5535
rect 2871 5531 2872 5535
rect 2866 5530 2872 5531
rect 3074 5535 3080 5536
rect 3074 5531 3075 5535
rect 3079 5531 3080 5535
rect 3074 5530 3080 5531
rect 2894 5520 2900 5521
rect 3084 5520 3086 5578
rect 3276 5536 3278 5597
rect 3282 5583 3288 5584
rect 3282 5579 3283 5583
rect 3287 5579 3288 5583
rect 3282 5578 3288 5579
rect 3274 5535 3280 5536
rect 3274 5531 3275 5535
rect 3279 5531 3280 5535
rect 3274 5530 3280 5531
rect 3102 5520 3108 5521
rect 3284 5520 3286 5578
rect 3476 5536 3478 5597
rect 3482 5583 3488 5584
rect 3482 5579 3483 5583
rect 3487 5579 3488 5583
rect 3482 5578 3488 5579
rect 3474 5535 3480 5536
rect 3474 5531 3475 5535
rect 3479 5531 3480 5535
rect 3474 5530 3480 5531
rect 3302 5520 3308 5521
rect 3484 5520 3486 5578
rect 3652 5536 3654 5597
rect 3658 5583 3664 5584
rect 3658 5579 3659 5583
rect 3663 5579 3664 5583
rect 3658 5578 3664 5579
rect 3650 5535 3656 5536
rect 3650 5531 3651 5535
rect 3655 5531 3656 5535
rect 3650 5530 3656 5531
rect 3502 5520 3508 5521
rect 3660 5520 3662 5578
rect 3678 5520 3684 5521
rect 3776 5520 3778 5622
rect 3800 5603 3802 5671
rect 3839 5669 3843 5670
rect 4107 5674 4111 5675
rect 4107 5669 4111 5670
rect 4243 5674 4247 5675
rect 4243 5669 4247 5670
rect 4379 5674 4383 5675
rect 4379 5669 4383 5670
rect 4515 5674 4519 5675
rect 4515 5669 4519 5670
rect 4651 5674 4655 5675
rect 4651 5669 4655 5670
rect 4787 5674 4791 5675
rect 4787 5669 4791 5670
rect 4923 5674 4927 5675
rect 4923 5669 4927 5670
rect 5059 5674 5063 5675
rect 5059 5669 5063 5670
rect 5195 5674 5199 5675
rect 5195 5669 5199 5670
rect 5663 5674 5667 5675
rect 5663 5669 5667 5670
rect 3840 5609 3842 5669
rect 3838 5608 3844 5609
rect 4108 5608 4110 5669
rect 4202 5655 4208 5656
rect 4202 5651 4203 5655
rect 4207 5651 4208 5655
rect 4202 5650 4208 5651
rect 3838 5604 3839 5608
rect 3843 5604 3844 5608
rect 3838 5603 3844 5604
rect 4106 5607 4112 5608
rect 4106 5603 4107 5607
rect 4111 5603 4112 5607
rect 3799 5602 3803 5603
rect 4106 5602 4112 5603
rect 3799 5597 3803 5598
rect 3800 5537 3802 5597
rect 4134 5592 4140 5593
rect 3838 5591 3844 5592
rect 3838 5587 3839 5591
rect 3843 5587 3844 5591
rect 4134 5588 4135 5592
rect 4139 5588 4140 5592
rect 4134 5587 4140 5588
rect 3838 5586 3844 5587
rect 3798 5536 3804 5537
rect 3798 5532 3799 5536
rect 3803 5532 3804 5536
rect 3798 5531 3804 5532
rect 3840 5531 3842 5586
rect 4136 5531 4138 5587
rect 4204 5560 4206 5650
rect 4244 5608 4246 5669
rect 4250 5655 4256 5656
rect 4250 5651 4251 5655
rect 4255 5651 4256 5655
rect 4250 5650 4256 5651
rect 4242 5607 4248 5608
rect 4242 5603 4243 5607
rect 4247 5603 4248 5607
rect 4242 5602 4248 5603
rect 4252 5592 4254 5650
rect 4380 5608 4382 5669
rect 4386 5655 4392 5656
rect 4386 5651 4387 5655
rect 4391 5651 4392 5655
rect 4386 5650 4392 5651
rect 4378 5607 4384 5608
rect 4378 5603 4379 5607
rect 4383 5603 4384 5607
rect 4378 5602 4384 5603
rect 4270 5592 4276 5593
rect 4388 5592 4390 5650
rect 4516 5608 4518 5669
rect 4522 5655 4528 5656
rect 4522 5651 4523 5655
rect 4527 5651 4528 5655
rect 4522 5650 4528 5651
rect 4514 5607 4520 5608
rect 4514 5603 4515 5607
rect 4519 5603 4520 5607
rect 4514 5602 4520 5603
rect 4406 5592 4412 5593
rect 4524 5592 4526 5650
rect 4652 5608 4654 5669
rect 4658 5655 4664 5656
rect 4658 5651 4659 5655
rect 4663 5651 4664 5655
rect 4658 5650 4664 5651
rect 4650 5607 4656 5608
rect 4650 5603 4651 5607
rect 4655 5603 4656 5607
rect 4650 5602 4656 5603
rect 4542 5592 4548 5593
rect 4660 5592 4662 5650
rect 4788 5608 4790 5669
rect 4794 5655 4800 5656
rect 4794 5651 4795 5655
rect 4799 5651 4800 5655
rect 4794 5650 4800 5651
rect 4786 5607 4792 5608
rect 4786 5603 4787 5607
rect 4791 5603 4792 5607
rect 4786 5602 4792 5603
rect 4678 5592 4684 5593
rect 4796 5592 4798 5650
rect 4924 5608 4926 5669
rect 4930 5655 4936 5656
rect 4930 5651 4931 5655
rect 4935 5651 4936 5655
rect 4930 5650 4936 5651
rect 4922 5607 4928 5608
rect 4922 5603 4923 5607
rect 4927 5603 4928 5607
rect 4922 5602 4928 5603
rect 4814 5592 4820 5593
rect 4932 5592 4934 5650
rect 5060 5608 5062 5669
rect 5066 5655 5072 5656
rect 5066 5651 5067 5655
rect 5071 5651 5072 5655
rect 5066 5650 5072 5651
rect 5058 5607 5064 5608
rect 5058 5603 5059 5607
rect 5063 5603 5064 5607
rect 5058 5602 5064 5603
rect 4950 5592 4956 5593
rect 5068 5592 5070 5650
rect 5196 5608 5198 5669
rect 5202 5655 5208 5656
rect 5202 5651 5203 5655
rect 5207 5651 5208 5655
rect 5202 5650 5208 5651
rect 5194 5607 5200 5608
rect 5194 5603 5195 5607
rect 5199 5603 5200 5607
rect 5194 5602 5200 5603
rect 5086 5592 5092 5593
rect 5204 5592 5206 5650
rect 5664 5609 5666 5669
rect 5662 5608 5668 5609
rect 5662 5604 5663 5608
rect 5667 5604 5668 5608
rect 5662 5603 5668 5604
rect 5222 5592 5228 5593
rect 4250 5591 4256 5592
rect 4250 5587 4251 5591
rect 4255 5587 4256 5591
rect 4270 5588 4271 5592
rect 4275 5588 4276 5592
rect 4270 5587 4276 5588
rect 4386 5591 4392 5592
rect 4386 5587 4387 5591
rect 4391 5587 4392 5591
rect 4406 5588 4407 5592
rect 4411 5588 4412 5592
rect 4406 5587 4412 5588
rect 4522 5591 4528 5592
rect 4522 5587 4523 5591
rect 4527 5587 4528 5591
rect 4542 5588 4543 5592
rect 4547 5588 4548 5592
rect 4542 5587 4548 5588
rect 4658 5591 4664 5592
rect 4658 5587 4659 5591
rect 4663 5587 4664 5591
rect 4678 5588 4679 5592
rect 4683 5588 4684 5592
rect 4678 5587 4684 5588
rect 4794 5591 4800 5592
rect 4794 5587 4795 5591
rect 4799 5587 4800 5591
rect 4814 5588 4815 5592
rect 4819 5588 4820 5592
rect 4814 5587 4820 5588
rect 4930 5591 4936 5592
rect 4930 5587 4931 5591
rect 4935 5587 4936 5591
rect 4950 5588 4951 5592
rect 4955 5588 4956 5592
rect 4950 5587 4956 5588
rect 5066 5591 5072 5592
rect 5066 5587 5067 5591
rect 5071 5587 5072 5591
rect 5086 5588 5087 5592
rect 5091 5588 5092 5592
rect 5086 5587 5092 5588
rect 5202 5591 5208 5592
rect 5202 5587 5203 5591
rect 5207 5587 5208 5591
rect 5222 5588 5223 5592
rect 5227 5588 5228 5592
rect 5222 5587 5228 5588
rect 5314 5591 5320 5592
rect 5314 5587 5315 5591
rect 5319 5587 5320 5591
rect 4250 5586 4256 5587
rect 4202 5559 4208 5560
rect 4202 5555 4203 5559
rect 4207 5555 4208 5559
rect 4202 5554 4208 5555
rect 4272 5531 4274 5587
rect 4386 5586 4392 5587
rect 4398 5559 4404 5560
rect 4398 5555 4399 5559
rect 4403 5555 4404 5559
rect 4398 5554 4404 5555
rect 3839 5530 3843 5531
rect 3839 5525 3843 5526
rect 4135 5530 4139 5531
rect 4135 5525 4139 5526
rect 4271 5530 4275 5531
rect 4271 5525 4275 5526
rect 4303 5530 4307 5531
rect 4303 5525 4307 5526
rect 1974 5519 1980 5520
rect 1974 5515 1975 5519
rect 1979 5515 1980 5519
rect 2022 5516 2023 5520
rect 2027 5516 2028 5520
rect 2022 5515 2028 5516
rect 2122 5519 2128 5520
rect 2122 5515 2123 5519
rect 2127 5515 2128 5519
rect 2230 5516 2231 5520
rect 2235 5516 2236 5520
rect 2230 5515 2236 5516
rect 2442 5519 2448 5520
rect 2442 5515 2443 5519
rect 2447 5515 2448 5519
rect 2462 5516 2463 5520
rect 2467 5516 2468 5520
rect 2462 5515 2468 5516
rect 2558 5519 2564 5520
rect 2558 5515 2559 5519
rect 2563 5515 2564 5519
rect 2686 5516 2687 5520
rect 2691 5516 2692 5520
rect 2686 5515 2692 5516
rect 2778 5519 2784 5520
rect 2778 5515 2779 5519
rect 2783 5515 2784 5519
rect 2894 5516 2895 5520
rect 2899 5516 2900 5520
rect 2894 5515 2900 5516
rect 3082 5519 3088 5520
rect 3082 5515 3083 5519
rect 3087 5515 3088 5519
rect 3102 5516 3103 5520
rect 3107 5516 3108 5520
rect 3102 5515 3108 5516
rect 3282 5519 3288 5520
rect 3282 5515 3283 5519
rect 3287 5515 3288 5519
rect 3302 5516 3303 5520
rect 3307 5516 3308 5520
rect 3302 5515 3308 5516
rect 3482 5519 3488 5520
rect 3482 5515 3483 5519
rect 3487 5515 3488 5519
rect 3502 5516 3503 5520
rect 3507 5516 3508 5520
rect 3502 5515 3508 5516
rect 3658 5519 3664 5520
rect 3658 5515 3659 5519
rect 3663 5515 3664 5519
rect 3678 5516 3679 5520
rect 3683 5516 3684 5520
rect 3678 5515 3684 5516
rect 3774 5519 3780 5520
rect 3774 5515 3775 5519
rect 3779 5515 3780 5519
rect 1974 5514 1980 5515
rect 1976 5491 1978 5514
rect 2024 5491 2026 5515
rect 2122 5514 2128 5515
rect 1975 5490 1979 5491
rect 1975 5485 1979 5486
rect 2023 5490 2027 5491
rect 2023 5485 2027 5486
rect 1934 5468 1940 5469
rect 1934 5464 1935 5468
rect 1939 5464 1940 5468
rect 1934 5463 1940 5464
rect 1976 5462 1978 5485
rect 1974 5461 1980 5462
rect 2024 5461 2026 5485
rect 1974 5457 1975 5461
rect 1979 5457 1980 5461
rect 1974 5456 1980 5457
rect 2022 5460 2028 5461
rect 2022 5456 2023 5460
rect 2027 5456 2028 5460
rect 2022 5455 2028 5456
rect 2114 5459 2120 5460
rect 2114 5455 2115 5459
rect 2119 5455 2120 5459
rect 2114 5454 2120 5455
rect 1454 5451 1460 5452
rect 1454 5447 1455 5451
rect 1459 5447 1460 5451
rect 1454 5446 1460 5447
rect 1934 5451 1940 5452
rect 1934 5447 1935 5451
rect 1939 5447 1940 5451
rect 1934 5446 1940 5447
rect 1456 5420 1458 5446
rect 1454 5419 1460 5420
rect 1454 5415 1455 5419
rect 1459 5415 1460 5419
rect 1454 5414 1460 5415
rect 1936 5403 1938 5446
rect 1994 5445 2000 5446
rect 1974 5444 1980 5445
rect 1974 5440 1975 5444
rect 1979 5440 1980 5444
rect 1994 5441 1995 5445
rect 1999 5441 2000 5445
rect 1994 5440 2000 5441
rect 1974 5439 1980 5440
rect 1495 5402 1499 5403
rect 1495 5397 1499 5398
rect 1663 5402 1667 5403
rect 1663 5397 1667 5398
rect 1815 5402 1819 5403
rect 1815 5397 1819 5398
rect 1935 5402 1939 5403
rect 1935 5397 1939 5398
rect 1496 5373 1498 5397
rect 1664 5373 1666 5397
rect 1816 5373 1818 5397
rect 1936 5374 1938 5397
rect 1934 5373 1940 5374
rect 1494 5372 1500 5373
rect 1662 5372 1668 5373
rect 1814 5372 1820 5373
rect 1274 5371 1280 5372
rect 1274 5367 1275 5371
rect 1279 5367 1280 5371
rect 1334 5368 1335 5372
rect 1339 5368 1340 5372
rect 1334 5367 1340 5368
rect 1426 5371 1432 5372
rect 1426 5367 1427 5371
rect 1431 5367 1432 5371
rect 1494 5368 1495 5372
rect 1499 5368 1500 5372
rect 1494 5367 1500 5368
rect 1594 5371 1600 5372
rect 1594 5367 1595 5371
rect 1599 5367 1600 5371
rect 1662 5368 1663 5372
rect 1667 5368 1668 5372
rect 1662 5367 1668 5368
rect 1758 5371 1764 5372
rect 1758 5367 1759 5371
rect 1763 5367 1764 5371
rect 1814 5368 1815 5372
rect 1819 5368 1820 5372
rect 1814 5367 1820 5368
rect 1906 5371 1912 5372
rect 1906 5367 1907 5371
rect 1911 5367 1912 5371
rect 1934 5369 1935 5373
rect 1939 5369 1940 5373
rect 1934 5368 1940 5369
rect 1274 5366 1280 5367
rect 1426 5366 1432 5367
rect 1594 5366 1600 5367
rect 1758 5366 1764 5367
rect 1906 5366 1912 5367
rect 1250 5307 1256 5308
rect 1250 5303 1251 5307
rect 1255 5303 1256 5307
rect 1250 5302 1256 5303
rect 1276 5300 1278 5366
rect 1306 5357 1312 5358
rect 1306 5353 1307 5357
rect 1311 5353 1312 5357
rect 1306 5352 1312 5353
rect 1466 5357 1472 5358
rect 1466 5353 1467 5357
rect 1471 5353 1472 5357
rect 1466 5352 1472 5353
rect 1274 5299 1280 5300
rect 1274 5295 1275 5299
rect 1279 5295 1280 5299
rect 1274 5294 1280 5295
rect 1308 5287 1310 5352
rect 1468 5287 1470 5352
rect 1596 5308 1598 5366
rect 1634 5357 1640 5358
rect 1634 5353 1635 5357
rect 1639 5353 1640 5357
rect 1634 5352 1640 5353
rect 1550 5307 1556 5308
rect 1550 5303 1551 5307
rect 1555 5303 1556 5307
rect 1550 5302 1556 5303
rect 1594 5307 1600 5308
rect 1594 5303 1595 5307
rect 1599 5303 1600 5307
rect 1594 5302 1600 5303
rect 1155 5286 1159 5287
rect 1155 5281 1159 5282
rect 1243 5286 1247 5287
rect 1243 5281 1247 5282
rect 1307 5286 1311 5287
rect 1307 5281 1311 5282
rect 1427 5286 1431 5287
rect 1427 5281 1431 5282
rect 1467 5286 1471 5287
rect 1467 5281 1471 5282
rect 1134 5271 1140 5272
rect 1134 5267 1135 5271
rect 1139 5267 1140 5271
rect 1134 5266 1140 5267
rect 1244 5220 1246 5281
rect 1250 5267 1256 5268
rect 1250 5263 1251 5267
rect 1255 5263 1256 5267
rect 1250 5262 1256 5263
rect 898 5219 904 5220
rect 898 5215 899 5219
rect 903 5215 904 5219
rect 898 5214 904 5215
rect 1066 5219 1072 5220
rect 1066 5215 1067 5219
rect 1071 5215 1072 5219
rect 1066 5214 1072 5215
rect 1242 5219 1248 5220
rect 1242 5215 1243 5219
rect 1247 5215 1248 5219
rect 1242 5214 1248 5215
rect 926 5204 932 5205
rect 110 5203 116 5204
rect 110 5199 111 5203
rect 115 5199 116 5203
rect 614 5200 615 5204
rect 619 5200 620 5204
rect 614 5199 620 5200
rect 710 5203 716 5204
rect 710 5199 711 5203
rect 715 5199 716 5203
rect 766 5200 767 5204
rect 771 5200 772 5204
rect 766 5199 772 5200
rect 862 5203 868 5204
rect 862 5199 863 5203
rect 867 5199 868 5203
rect 926 5200 927 5204
rect 931 5200 932 5204
rect 926 5199 932 5200
rect 1094 5204 1100 5205
rect 1252 5204 1254 5262
rect 1366 5239 1372 5240
rect 1366 5235 1367 5239
rect 1371 5235 1372 5239
rect 1366 5234 1372 5235
rect 1270 5204 1276 5205
rect 1368 5204 1370 5234
rect 1428 5220 1430 5281
rect 1542 5271 1548 5272
rect 1542 5267 1543 5271
rect 1547 5267 1548 5271
rect 1542 5266 1548 5267
rect 1426 5219 1432 5220
rect 1426 5215 1427 5219
rect 1431 5215 1432 5219
rect 1426 5214 1432 5215
rect 1454 5204 1460 5205
rect 1094 5200 1095 5204
rect 1099 5200 1100 5204
rect 1094 5199 1100 5200
rect 1250 5203 1256 5204
rect 1250 5199 1251 5203
rect 1255 5199 1256 5203
rect 1270 5200 1271 5204
rect 1275 5200 1276 5204
rect 1270 5199 1276 5200
rect 1366 5203 1372 5204
rect 1366 5199 1367 5203
rect 1371 5199 1372 5203
rect 1454 5200 1455 5204
rect 1459 5200 1460 5204
rect 1454 5199 1460 5200
rect 110 5198 116 5199
rect 112 5163 114 5198
rect 616 5163 618 5199
rect 710 5198 716 5199
rect 712 5195 714 5198
rect 704 5193 714 5195
rect 111 5162 115 5163
rect 111 5157 115 5158
rect 367 5162 371 5163
rect 367 5157 371 5158
rect 535 5162 539 5163
rect 535 5157 539 5158
rect 615 5162 619 5163
rect 615 5157 619 5158
rect 112 5134 114 5157
rect 110 5133 116 5134
rect 368 5133 370 5157
rect 536 5133 538 5157
rect 110 5129 111 5133
rect 115 5129 116 5133
rect 110 5128 116 5129
rect 366 5132 372 5133
rect 534 5132 540 5133
rect 366 5128 367 5132
rect 371 5128 372 5132
rect 366 5127 372 5128
rect 466 5131 472 5132
rect 466 5127 467 5131
rect 471 5127 472 5131
rect 534 5128 535 5132
rect 539 5128 540 5132
rect 534 5127 540 5128
rect 630 5131 636 5132
rect 630 5127 631 5131
rect 635 5127 636 5131
rect 466 5126 472 5127
rect 630 5126 636 5127
rect 338 5117 344 5118
rect 110 5116 116 5117
rect 110 5112 111 5116
rect 115 5112 116 5116
rect 338 5113 339 5117
rect 343 5113 344 5117
rect 338 5112 344 5113
rect 110 5111 116 5112
rect 112 5047 114 5111
rect 340 5047 342 5112
rect 434 5111 440 5112
rect 434 5107 435 5111
rect 439 5107 440 5111
rect 434 5106 440 5107
rect 436 5068 438 5106
rect 468 5068 470 5126
rect 506 5117 512 5118
rect 506 5113 507 5117
rect 511 5113 512 5117
rect 506 5112 512 5113
rect 434 5067 440 5068
rect 434 5063 435 5067
rect 439 5063 440 5067
rect 434 5062 440 5063
rect 466 5067 472 5068
rect 466 5063 467 5067
rect 471 5063 472 5067
rect 466 5062 472 5063
rect 508 5047 510 5112
rect 111 5046 115 5047
rect 111 5041 115 5042
rect 131 5046 135 5047
rect 131 5041 135 5042
rect 323 5046 327 5047
rect 323 5041 327 5042
rect 339 5046 343 5047
rect 339 5041 343 5042
rect 507 5046 511 5047
rect 507 5041 511 5042
rect 555 5046 559 5047
rect 555 5041 559 5042
rect 112 4981 114 5041
rect 110 4980 116 4981
rect 132 4980 134 5041
rect 226 5027 232 5028
rect 226 5023 227 5027
rect 231 5023 232 5027
rect 226 5022 232 5023
rect 228 4992 230 5022
rect 226 4991 232 4992
rect 226 4987 227 4991
rect 231 4987 232 4991
rect 226 4986 232 4987
rect 324 4980 326 5041
rect 330 5027 336 5028
rect 330 5023 331 5027
rect 335 5023 336 5027
rect 330 5022 336 5023
rect 110 4976 111 4980
rect 115 4976 116 4980
rect 110 4975 116 4976
rect 130 4979 136 4980
rect 130 4975 131 4979
rect 135 4975 136 4979
rect 130 4974 136 4975
rect 322 4979 328 4980
rect 322 4975 323 4979
rect 327 4975 328 4979
rect 322 4974 328 4975
rect 158 4964 164 4965
rect 332 4964 334 5022
rect 556 4980 558 5041
rect 632 5032 634 5126
rect 682 5117 688 5118
rect 682 5113 683 5117
rect 687 5113 688 5117
rect 682 5112 688 5113
rect 684 5047 686 5112
rect 704 5068 706 5193
rect 768 5163 770 5199
rect 862 5198 868 5199
rect 928 5163 930 5199
rect 1096 5163 1098 5199
rect 1250 5198 1256 5199
rect 1272 5163 1274 5199
rect 1366 5198 1372 5199
rect 1456 5163 1458 5199
rect 711 5162 715 5163
rect 711 5157 715 5158
rect 767 5162 771 5163
rect 767 5157 771 5158
rect 895 5162 899 5163
rect 895 5157 899 5158
rect 927 5162 931 5163
rect 927 5157 931 5158
rect 1079 5162 1083 5163
rect 1079 5157 1083 5158
rect 1095 5162 1099 5163
rect 1095 5157 1099 5158
rect 1263 5162 1267 5163
rect 1263 5157 1267 5158
rect 1271 5162 1275 5163
rect 1271 5157 1275 5158
rect 1447 5162 1451 5163
rect 1447 5157 1451 5158
rect 1455 5162 1459 5163
rect 1455 5157 1459 5158
rect 712 5133 714 5157
rect 896 5133 898 5157
rect 1080 5133 1082 5157
rect 1264 5133 1266 5157
rect 1448 5133 1450 5157
rect 710 5132 716 5133
rect 710 5128 711 5132
rect 715 5128 716 5132
rect 710 5127 716 5128
rect 894 5132 900 5133
rect 1078 5132 1084 5133
rect 1262 5132 1268 5133
rect 894 5128 895 5132
rect 899 5128 900 5132
rect 894 5127 900 5128
rect 1014 5131 1020 5132
rect 1014 5127 1015 5131
rect 1019 5127 1020 5131
rect 1078 5128 1079 5132
rect 1083 5128 1084 5132
rect 1078 5127 1084 5128
rect 1170 5131 1176 5132
rect 1170 5127 1171 5131
rect 1175 5127 1176 5131
rect 1262 5128 1263 5132
rect 1267 5128 1268 5132
rect 1262 5127 1268 5128
rect 1446 5132 1452 5133
rect 1544 5132 1546 5266
rect 1552 5204 1554 5302
rect 1636 5287 1638 5352
rect 1760 5300 1762 5366
rect 1786 5357 1792 5358
rect 1786 5353 1787 5357
rect 1791 5353 1792 5357
rect 1786 5352 1792 5353
rect 1758 5299 1764 5300
rect 1758 5295 1759 5299
rect 1763 5295 1764 5299
rect 1758 5294 1764 5295
rect 1788 5287 1790 5352
rect 1619 5286 1623 5287
rect 1619 5281 1623 5282
rect 1635 5286 1639 5287
rect 1635 5281 1639 5282
rect 1787 5286 1791 5287
rect 1787 5281 1791 5282
rect 1620 5220 1622 5281
rect 1778 5271 1784 5272
rect 1778 5267 1779 5271
rect 1783 5267 1784 5271
rect 1778 5266 1784 5267
rect 1618 5219 1624 5220
rect 1618 5215 1619 5219
rect 1623 5215 1624 5219
rect 1618 5214 1624 5215
rect 1780 5212 1782 5266
rect 1788 5220 1790 5281
rect 1908 5272 1910 5366
rect 1934 5356 1940 5357
rect 1934 5352 1935 5356
rect 1939 5352 1940 5356
rect 1976 5355 1978 5439
rect 1996 5355 1998 5440
rect 1934 5351 1940 5352
rect 1975 5354 1979 5355
rect 1936 5287 1938 5351
rect 1975 5349 1979 5350
rect 1995 5354 1999 5355
rect 1995 5349 1999 5350
rect 2051 5354 2055 5355
rect 2051 5349 2055 5350
rect 1976 5289 1978 5349
rect 1974 5288 1980 5289
rect 2052 5288 2054 5349
rect 2116 5308 2118 5454
rect 2124 5396 2126 5514
rect 2232 5491 2234 5515
rect 2442 5514 2448 5515
rect 2464 5491 2466 5515
rect 2558 5514 2564 5515
rect 2167 5490 2171 5491
rect 2167 5485 2171 5486
rect 2231 5490 2235 5491
rect 2231 5485 2235 5486
rect 2343 5490 2347 5491
rect 2343 5485 2347 5486
rect 2463 5490 2467 5491
rect 2463 5485 2467 5486
rect 2527 5490 2531 5491
rect 2527 5485 2531 5486
rect 2168 5461 2170 5485
rect 2344 5461 2346 5485
rect 2528 5461 2530 5485
rect 2166 5460 2172 5461
rect 2342 5460 2348 5461
rect 2526 5460 2532 5461
rect 2166 5456 2167 5460
rect 2171 5456 2172 5460
rect 2166 5455 2172 5456
rect 2278 5459 2284 5460
rect 2278 5455 2279 5459
rect 2283 5455 2284 5459
rect 2342 5456 2343 5460
rect 2347 5456 2348 5460
rect 2342 5455 2348 5456
rect 2442 5459 2448 5460
rect 2442 5455 2443 5459
rect 2447 5455 2448 5459
rect 2526 5456 2527 5460
rect 2531 5456 2532 5460
rect 2526 5455 2532 5456
rect 2278 5454 2284 5455
rect 2442 5454 2448 5455
rect 2138 5445 2144 5446
rect 2138 5441 2139 5445
rect 2143 5441 2144 5445
rect 2138 5440 2144 5441
rect 2122 5395 2128 5396
rect 2122 5391 2123 5395
rect 2127 5391 2128 5395
rect 2122 5390 2128 5391
rect 2140 5355 2142 5440
rect 2280 5396 2282 5454
rect 2314 5445 2320 5446
rect 2314 5441 2315 5445
rect 2319 5441 2320 5445
rect 2314 5440 2320 5441
rect 2278 5395 2284 5396
rect 2278 5391 2279 5395
rect 2283 5391 2284 5395
rect 2278 5390 2284 5391
rect 2316 5355 2318 5440
rect 2139 5354 2143 5355
rect 2139 5349 2143 5350
rect 2315 5354 2319 5355
rect 2315 5349 2319 5350
rect 2444 5340 2446 5454
rect 2498 5445 2504 5446
rect 2498 5441 2499 5445
rect 2503 5441 2504 5445
rect 2498 5440 2504 5441
rect 2500 5355 2502 5440
rect 2560 5396 2562 5514
rect 2688 5491 2690 5515
rect 2778 5514 2784 5515
rect 2896 5491 2898 5515
rect 3082 5514 3088 5515
rect 3104 5491 3106 5515
rect 3282 5514 3288 5515
rect 3304 5491 3306 5515
rect 3482 5514 3488 5515
rect 3504 5491 3506 5515
rect 3658 5514 3664 5515
rect 3680 5491 3682 5515
rect 3774 5514 3780 5515
rect 3798 5519 3804 5520
rect 3798 5515 3799 5519
rect 3803 5515 3804 5519
rect 3798 5514 3804 5515
rect 3800 5491 3802 5514
rect 3840 5502 3842 5525
rect 3838 5501 3844 5502
rect 4304 5501 4306 5525
rect 3838 5497 3839 5501
rect 3843 5497 3844 5501
rect 3838 5496 3844 5497
rect 4302 5500 4308 5501
rect 4400 5500 4402 5554
rect 4408 5531 4410 5587
rect 4522 5586 4528 5587
rect 4544 5531 4546 5587
rect 4658 5586 4664 5587
rect 4680 5531 4682 5587
rect 4794 5586 4800 5587
rect 4816 5531 4818 5587
rect 4930 5586 4936 5587
rect 4952 5531 4954 5587
rect 5066 5586 5072 5587
rect 5088 5531 5090 5587
rect 5202 5586 5208 5587
rect 5224 5531 5226 5587
rect 5314 5586 5320 5587
rect 5662 5591 5668 5592
rect 5662 5587 5663 5591
rect 5667 5587 5668 5591
rect 5662 5586 5668 5587
rect 4407 5530 4411 5531
rect 4407 5525 4411 5526
rect 4511 5530 4515 5531
rect 4511 5525 4515 5526
rect 4543 5530 4547 5531
rect 4543 5525 4547 5526
rect 4679 5530 4683 5531
rect 4679 5525 4683 5526
rect 4719 5530 4723 5531
rect 4719 5525 4723 5526
rect 4815 5530 4819 5531
rect 4815 5525 4819 5526
rect 4927 5530 4931 5531
rect 4927 5525 4931 5526
rect 4951 5530 4955 5531
rect 4951 5525 4955 5526
rect 5087 5530 5091 5531
rect 5087 5525 5091 5526
rect 5135 5530 5139 5531
rect 5135 5525 5139 5526
rect 5223 5530 5227 5531
rect 5223 5525 5227 5526
rect 4512 5501 4514 5525
rect 4720 5501 4722 5525
rect 4928 5501 4930 5525
rect 5136 5501 5138 5525
rect 4510 5500 4516 5501
rect 4718 5500 4724 5501
rect 4926 5500 4932 5501
rect 5134 5500 5140 5501
rect 4302 5496 4303 5500
rect 4307 5496 4308 5500
rect 4302 5495 4308 5496
rect 4398 5499 4404 5500
rect 4398 5495 4399 5499
rect 4403 5495 4404 5499
rect 4510 5496 4511 5500
rect 4515 5496 4516 5500
rect 4510 5495 4516 5496
rect 4602 5499 4608 5500
rect 4602 5495 4603 5499
rect 4607 5495 4608 5499
rect 4718 5496 4719 5500
rect 4723 5496 4724 5500
rect 4718 5495 4724 5496
rect 4818 5499 4824 5500
rect 4818 5495 4819 5499
rect 4823 5495 4824 5499
rect 4926 5496 4927 5500
rect 4931 5496 4932 5500
rect 4926 5495 4932 5496
rect 5022 5499 5028 5500
rect 5022 5495 5023 5499
rect 5027 5495 5028 5499
rect 5134 5496 5135 5500
rect 5139 5496 5140 5500
rect 5134 5495 5140 5496
rect 5230 5499 5236 5500
rect 5230 5495 5231 5499
rect 5235 5495 5236 5499
rect 4398 5494 4404 5495
rect 4602 5494 4608 5495
rect 4818 5494 4824 5495
rect 5022 5494 5028 5495
rect 5230 5494 5236 5495
rect 2687 5490 2691 5491
rect 2687 5485 2691 5486
rect 2719 5490 2723 5491
rect 2719 5485 2723 5486
rect 2895 5490 2899 5491
rect 2895 5485 2899 5486
rect 2911 5490 2915 5491
rect 2911 5485 2915 5486
rect 3103 5490 3107 5491
rect 3103 5485 3107 5486
rect 3111 5490 3115 5491
rect 3111 5485 3115 5486
rect 3303 5490 3307 5491
rect 3303 5485 3307 5486
rect 3311 5490 3315 5491
rect 3311 5485 3315 5486
rect 3503 5490 3507 5491
rect 3503 5485 3507 5486
rect 3679 5490 3683 5491
rect 3679 5485 3683 5486
rect 3799 5490 3803 5491
rect 3799 5485 3803 5486
rect 4274 5485 4280 5486
rect 2720 5461 2722 5485
rect 2912 5461 2914 5485
rect 3112 5461 3114 5485
rect 3312 5461 3314 5485
rect 3800 5462 3802 5485
rect 3838 5484 3844 5485
rect 3838 5480 3839 5484
rect 3843 5480 3844 5484
rect 4274 5481 4275 5485
rect 4279 5481 4280 5485
rect 4274 5480 4280 5481
rect 4482 5485 4488 5486
rect 4482 5481 4483 5485
rect 4487 5481 4488 5485
rect 4482 5480 4488 5481
rect 3838 5479 3844 5480
rect 3798 5461 3804 5462
rect 2718 5460 2724 5461
rect 2718 5456 2719 5460
rect 2723 5456 2724 5460
rect 2718 5455 2724 5456
rect 2910 5460 2916 5461
rect 3110 5460 3116 5461
rect 3310 5460 3316 5461
rect 2910 5456 2911 5460
rect 2915 5456 2916 5460
rect 2910 5455 2916 5456
rect 3010 5459 3016 5460
rect 3010 5455 3011 5459
rect 3015 5455 3016 5459
rect 3110 5456 3111 5460
rect 3115 5456 3116 5460
rect 3110 5455 3116 5456
rect 3210 5459 3216 5460
rect 3210 5455 3211 5459
rect 3215 5455 3216 5459
rect 3310 5456 3311 5460
rect 3315 5456 3316 5460
rect 3798 5457 3799 5461
rect 3803 5457 3804 5461
rect 3798 5456 3804 5457
rect 3310 5455 3316 5456
rect 3010 5454 3016 5455
rect 3210 5454 3216 5455
rect 2690 5445 2696 5446
rect 2690 5441 2691 5445
rect 2695 5441 2696 5445
rect 2690 5440 2696 5441
rect 2882 5445 2888 5446
rect 2882 5441 2883 5445
rect 2887 5441 2888 5445
rect 2882 5440 2888 5441
rect 2558 5395 2564 5396
rect 2558 5391 2559 5395
rect 2563 5391 2564 5395
rect 2558 5390 2564 5391
rect 2692 5355 2694 5440
rect 2884 5355 2886 5440
rect 3012 5396 3014 5454
rect 3082 5445 3088 5446
rect 3082 5441 3083 5445
rect 3087 5441 3088 5445
rect 3082 5440 3088 5441
rect 2978 5395 2984 5396
rect 2978 5391 2979 5395
rect 2983 5391 2984 5395
rect 2978 5390 2984 5391
rect 3010 5395 3016 5396
rect 3010 5391 3011 5395
rect 3015 5391 3016 5395
rect 3010 5390 3016 5391
rect 2459 5354 2463 5355
rect 2459 5349 2463 5350
rect 2499 5354 2503 5355
rect 2499 5349 2503 5350
rect 2691 5354 2695 5355
rect 2691 5349 2695 5350
rect 2859 5354 2863 5355
rect 2859 5349 2863 5350
rect 2883 5354 2887 5355
rect 2883 5349 2887 5350
rect 2442 5339 2448 5340
rect 2146 5335 2152 5336
rect 2146 5331 2147 5335
rect 2151 5331 2152 5335
rect 2442 5335 2443 5339
rect 2447 5335 2448 5339
rect 2442 5334 2448 5335
rect 2146 5330 2152 5331
rect 2148 5316 2150 5330
rect 2146 5315 2152 5316
rect 2146 5311 2147 5315
rect 2151 5311 2152 5315
rect 2146 5310 2152 5311
rect 2114 5307 2120 5308
rect 2114 5303 2115 5307
rect 2119 5303 2120 5307
rect 2114 5302 2120 5303
rect 2460 5288 2462 5349
rect 2582 5315 2588 5316
rect 2582 5311 2583 5315
rect 2587 5311 2588 5315
rect 2582 5310 2588 5311
rect 1935 5286 1939 5287
rect 1974 5284 1975 5288
rect 1979 5284 1980 5288
rect 1974 5283 1980 5284
rect 2050 5287 2056 5288
rect 2050 5283 2051 5287
rect 2055 5283 2056 5287
rect 2050 5282 2056 5283
rect 2458 5287 2464 5288
rect 2458 5283 2459 5287
rect 2463 5283 2464 5287
rect 2458 5282 2464 5283
rect 1935 5281 1939 5282
rect 1906 5271 1912 5272
rect 1906 5267 1907 5271
rect 1911 5267 1912 5271
rect 1906 5266 1912 5267
rect 1936 5221 1938 5281
rect 2078 5272 2084 5273
rect 2486 5272 2492 5273
rect 2584 5272 2586 5310
rect 2860 5288 2862 5349
rect 2866 5335 2872 5336
rect 2866 5331 2867 5335
rect 2871 5331 2872 5335
rect 2866 5330 2872 5331
rect 2858 5287 2864 5288
rect 2858 5283 2859 5287
rect 2863 5283 2864 5287
rect 2858 5282 2864 5283
rect 1974 5271 1980 5272
rect 1974 5267 1975 5271
rect 1979 5267 1980 5271
rect 2078 5268 2079 5272
rect 2083 5268 2084 5272
rect 2078 5267 2084 5268
rect 2198 5271 2204 5272
rect 2198 5267 2199 5271
rect 2203 5267 2204 5271
rect 2486 5268 2487 5272
rect 2491 5268 2492 5272
rect 2486 5267 2492 5268
rect 2582 5271 2588 5272
rect 2582 5267 2583 5271
rect 2587 5267 2588 5271
rect 1974 5266 1980 5267
rect 1976 5243 1978 5266
rect 2080 5243 2082 5267
rect 2198 5266 2204 5267
rect 1975 5242 1979 5243
rect 1975 5237 1979 5238
rect 2079 5242 2083 5243
rect 2079 5237 2083 5238
rect 1934 5220 1940 5221
rect 1786 5219 1792 5220
rect 1786 5215 1787 5219
rect 1791 5215 1792 5219
rect 1934 5216 1935 5220
rect 1939 5216 1940 5220
rect 1934 5215 1940 5216
rect 1786 5214 1792 5215
rect 1976 5214 1978 5237
rect 1974 5213 1980 5214
rect 1778 5211 1784 5212
rect 1778 5207 1779 5211
rect 1783 5207 1784 5211
rect 1974 5209 1975 5213
rect 1979 5209 1980 5213
rect 1974 5208 1980 5209
rect 1778 5206 1784 5207
rect 1646 5204 1652 5205
rect 1814 5204 1820 5205
rect 1550 5203 1556 5204
rect 1550 5199 1551 5203
rect 1555 5199 1556 5203
rect 1646 5200 1647 5204
rect 1651 5200 1652 5204
rect 1646 5199 1652 5200
rect 1746 5203 1752 5204
rect 1746 5199 1747 5203
rect 1751 5199 1752 5203
rect 1814 5200 1815 5204
rect 1819 5200 1820 5204
rect 1814 5199 1820 5200
rect 1934 5203 1940 5204
rect 1934 5199 1935 5203
rect 1939 5199 1940 5203
rect 1550 5198 1556 5199
rect 1648 5163 1650 5199
rect 1746 5198 1752 5199
rect 1631 5162 1635 5163
rect 1631 5157 1635 5158
rect 1647 5162 1651 5163
rect 1647 5157 1651 5158
rect 1632 5133 1634 5157
rect 1630 5132 1636 5133
rect 1446 5128 1447 5132
rect 1451 5128 1452 5132
rect 1446 5127 1452 5128
rect 1542 5131 1548 5132
rect 1542 5127 1543 5131
rect 1547 5127 1548 5131
rect 1630 5128 1631 5132
rect 1635 5128 1636 5132
rect 1630 5127 1636 5128
rect 1726 5131 1732 5132
rect 1726 5127 1727 5131
rect 1731 5127 1732 5131
rect 1014 5126 1020 5127
rect 1170 5126 1176 5127
rect 1542 5126 1548 5127
rect 1726 5126 1732 5127
rect 866 5117 872 5118
rect 866 5113 867 5117
rect 871 5113 872 5117
rect 866 5112 872 5113
rect 702 5067 708 5068
rect 702 5063 703 5067
rect 707 5063 708 5067
rect 702 5062 708 5063
rect 868 5047 870 5112
rect 1016 5068 1018 5126
rect 1050 5117 1056 5118
rect 1050 5113 1051 5117
rect 1055 5113 1056 5117
rect 1050 5112 1056 5113
rect 1172 5112 1174 5126
rect 1234 5117 1240 5118
rect 1234 5113 1235 5117
rect 1239 5113 1240 5117
rect 1234 5112 1240 5113
rect 1418 5117 1424 5118
rect 1418 5113 1419 5117
rect 1423 5113 1424 5117
rect 1418 5112 1424 5113
rect 1602 5117 1608 5118
rect 1602 5113 1603 5117
rect 1607 5113 1608 5117
rect 1602 5112 1608 5113
rect 1014 5067 1020 5068
rect 1014 5063 1015 5067
rect 1019 5063 1020 5067
rect 1014 5062 1020 5063
rect 1052 5047 1054 5112
rect 1170 5111 1176 5112
rect 1170 5107 1171 5111
rect 1175 5107 1176 5111
rect 1170 5106 1176 5107
rect 1236 5047 1238 5112
rect 1330 5067 1336 5068
rect 1330 5063 1331 5067
rect 1335 5063 1336 5067
rect 1330 5062 1336 5063
rect 683 5046 687 5047
rect 683 5041 687 5042
rect 811 5046 815 5047
rect 811 5041 815 5042
rect 867 5046 871 5047
rect 867 5041 871 5042
rect 1051 5046 1055 5047
rect 1051 5041 1055 5042
rect 1083 5046 1087 5047
rect 1083 5041 1087 5042
rect 1235 5046 1239 5047
rect 1235 5041 1239 5042
rect 630 5031 636 5032
rect 630 5027 631 5031
rect 635 5027 636 5031
rect 630 5026 636 5027
rect 812 4980 814 5041
rect 818 5027 824 5028
rect 818 5023 819 5027
rect 823 5023 824 5027
rect 818 5022 824 5023
rect 554 4979 560 4980
rect 554 4975 555 4979
rect 559 4975 560 4979
rect 554 4974 560 4975
rect 810 4979 816 4980
rect 810 4975 811 4979
rect 815 4975 816 4979
rect 810 4974 816 4975
rect 350 4964 356 4965
rect 582 4964 588 4965
rect 820 4964 822 5022
rect 1084 4980 1086 5041
rect 1090 5027 1096 5028
rect 1090 5023 1091 5027
rect 1095 5023 1096 5027
rect 1090 5022 1096 5023
rect 1082 4979 1088 4980
rect 1082 4975 1083 4979
rect 1087 4975 1088 4979
rect 1082 4974 1088 4975
rect 838 4964 844 4965
rect 1092 4964 1094 5022
rect 1206 4991 1212 4992
rect 1206 4987 1207 4991
rect 1211 4987 1212 4991
rect 1206 4986 1212 4987
rect 1110 4964 1116 4965
rect 1208 4964 1210 4986
rect 1332 4972 1334 5062
rect 1420 5047 1422 5112
rect 1604 5047 1606 5112
rect 1371 5046 1375 5047
rect 1371 5041 1375 5042
rect 1419 5046 1423 5047
rect 1419 5041 1423 5042
rect 1603 5046 1607 5047
rect 1603 5041 1607 5042
rect 1659 5046 1663 5047
rect 1659 5041 1663 5042
rect 1372 4980 1374 5041
rect 1466 5027 1472 5028
rect 1466 5023 1467 5027
rect 1471 5023 1472 5027
rect 1466 5022 1472 5023
rect 1468 4996 1470 5022
rect 1466 4995 1472 4996
rect 1466 4991 1467 4995
rect 1471 4991 1472 4995
rect 1466 4990 1472 4991
rect 1660 4980 1662 5041
rect 1728 5032 1730 5126
rect 1748 5068 1750 5198
rect 1816 5163 1818 5199
rect 1934 5198 1940 5199
rect 1936 5163 1938 5198
rect 1974 5196 1980 5197
rect 1974 5192 1975 5196
rect 1979 5192 1980 5196
rect 1974 5191 1980 5192
rect 1815 5162 1819 5163
rect 1815 5157 1819 5158
rect 1935 5162 1939 5163
rect 1935 5157 1939 5158
rect 1816 5133 1818 5157
rect 1936 5134 1938 5157
rect 1934 5133 1940 5134
rect 1814 5132 1820 5133
rect 1814 5128 1815 5132
rect 1819 5128 1820 5132
rect 1814 5127 1820 5128
rect 1910 5131 1916 5132
rect 1910 5127 1911 5131
rect 1915 5127 1916 5131
rect 1934 5129 1935 5133
rect 1939 5129 1940 5133
rect 1976 5131 1978 5191
rect 2200 5148 2202 5266
rect 2488 5243 2490 5267
rect 2582 5266 2588 5267
rect 2239 5242 2243 5243
rect 2239 5237 2243 5238
rect 2487 5242 2491 5243
rect 2487 5237 2491 5238
rect 2591 5242 2595 5243
rect 2591 5237 2595 5238
rect 2240 5213 2242 5237
rect 2592 5213 2594 5237
rect 2238 5212 2244 5213
rect 2590 5212 2596 5213
rect 2868 5212 2870 5330
rect 2886 5272 2892 5273
rect 2980 5272 2982 5390
rect 3084 5355 3086 5440
rect 3212 5396 3214 5454
rect 3282 5445 3288 5446
rect 3282 5441 3283 5445
rect 3287 5441 3288 5445
rect 3282 5440 3288 5441
rect 3798 5444 3804 5445
rect 3798 5440 3799 5444
rect 3803 5440 3804 5444
rect 3210 5395 3216 5396
rect 3210 5391 3211 5395
rect 3215 5391 3216 5395
rect 3210 5390 3216 5391
rect 3284 5355 3286 5440
rect 3798 5439 3804 5440
rect 3786 5379 3792 5380
rect 3786 5375 3787 5379
rect 3791 5375 3792 5379
rect 3786 5374 3792 5375
rect 3083 5354 3087 5355
rect 3083 5349 3087 5350
rect 3267 5354 3271 5355
rect 3267 5349 3271 5350
rect 3283 5354 3287 5355
rect 3283 5349 3287 5350
rect 3651 5354 3655 5355
rect 3651 5349 3655 5350
rect 3268 5288 3270 5349
rect 3652 5288 3654 5349
rect 3758 5343 3764 5344
rect 3758 5339 3759 5343
rect 3763 5339 3764 5343
rect 3758 5338 3764 5339
rect 3658 5335 3664 5336
rect 3658 5331 3659 5335
rect 3663 5331 3664 5335
rect 3658 5330 3664 5331
rect 3266 5287 3272 5288
rect 3266 5283 3267 5287
rect 3271 5283 3272 5287
rect 3266 5282 3272 5283
rect 3650 5287 3656 5288
rect 3650 5283 3651 5287
rect 3655 5283 3656 5287
rect 3650 5282 3656 5283
rect 3294 5272 3300 5273
rect 3660 5272 3662 5330
rect 3678 5272 3684 5273
rect 2886 5268 2887 5272
rect 2891 5268 2892 5272
rect 2886 5267 2892 5268
rect 2978 5271 2984 5272
rect 2978 5267 2979 5271
rect 2983 5267 2984 5271
rect 3294 5268 3295 5272
rect 3299 5268 3300 5272
rect 3294 5267 3300 5268
rect 3658 5271 3664 5272
rect 3658 5267 3659 5271
rect 3663 5267 3664 5271
rect 3678 5268 3679 5272
rect 3683 5268 3684 5272
rect 3678 5267 3684 5268
rect 2888 5243 2890 5267
rect 2978 5266 2984 5267
rect 3296 5243 3298 5267
rect 3658 5266 3664 5267
rect 3680 5243 3682 5267
rect 2887 5242 2891 5243
rect 2887 5237 2891 5238
rect 2943 5242 2947 5243
rect 2943 5237 2947 5238
rect 3295 5242 3299 5243
rect 3295 5237 3299 5238
rect 3303 5242 3307 5243
rect 3303 5237 3307 5238
rect 3663 5242 3667 5243
rect 3663 5237 3667 5238
rect 3679 5242 3683 5243
rect 3679 5237 3683 5238
rect 2944 5213 2946 5237
rect 3304 5213 3306 5237
rect 3664 5213 3666 5237
rect 2942 5212 2948 5213
rect 3302 5212 3308 5213
rect 3662 5212 3668 5213
rect 3760 5212 3762 5338
rect 3788 5272 3790 5374
rect 3800 5355 3802 5439
rect 3840 5395 3842 5479
rect 4276 5395 4278 5480
rect 4484 5395 4486 5480
rect 4558 5435 4564 5436
rect 4558 5431 4559 5435
rect 4563 5431 4564 5435
rect 4558 5430 4564 5431
rect 3839 5394 3843 5395
rect 3839 5389 3843 5390
rect 3859 5394 3863 5395
rect 3859 5389 3863 5390
rect 3995 5394 3999 5395
rect 3995 5389 3999 5390
rect 4131 5394 4135 5395
rect 4131 5389 4135 5390
rect 4275 5394 4279 5395
rect 4275 5389 4279 5390
rect 4435 5394 4439 5395
rect 4435 5389 4439 5390
rect 4483 5394 4487 5395
rect 4483 5389 4487 5390
rect 3799 5354 3803 5355
rect 3799 5349 3803 5350
rect 3800 5289 3802 5349
rect 3840 5329 3842 5389
rect 3838 5328 3844 5329
rect 3860 5328 3862 5389
rect 3996 5328 3998 5389
rect 4002 5375 4008 5376
rect 4002 5371 4003 5375
rect 4007 5371 4008 5375
rect 4002 5370 4008 5371
rect 3838 5324 3839 5328
rect 3843 5324 3844 5328
rect 3838 5323 3844 5324
rect 3858 5327 3864 5328
rect 3858 5323 3859 5327
rect 3863 5323 3864 5327
rect 3858 5322 3864 5323
rect 3994 5327 4000 5328
rect 3994 5323 3995 5327
rect 3999 5323 4000 5327
rect 3994 5322 4000 5323
rect 3886 5312 3892 5313
rect 4004 5312 4006 5370
rect 4132 5328 4134 5389
rect 4138 5375 4144 5376
rect 4138 5371 4139 5375
rect 4143 5371 4144 5375
rect 4138 5370 4144 5371
rect 4130 5327 4136 5328
rect 4130 5323 4131 5327
rect 4135 5323 4136 5327
rect 4130 5322 4136 5323
rect 4022 5312 4028 5313
rect 4140 5312 4142 5370
rect 4276 5328 4278 5389
rect 4282 5375 4288 5376
rect 4282 5371 4283 5375
rect 4287 5371 4288 5375
rect 4282 5370 4288 5371
rect 4274 5327 4280 5328
rect 4274 5323 4275 5327
rect 4279 5323 4280 5327
rect 4274 5322 4280 5323
rect 4158 5312 4164 5313
rect 4284 5312 4286 5370
rect 4436 5328 4438 5389
rect 4434 5327 4440 5328
rect 4434 5323 4435 5327
rect 4439 5323 4440 5327
rect 4434 5322 4440 5323
rect 4302 5312 4308 5313
rect 4462 5312 4468 5313
rect 4560 5312 4562 5430
rect 4604 5428 4606 5494
rect 4690 5485 4696 5486
rect 4690 5481 4691 5485
rect 4695 5481 4696 5485
rect 4690 5480 4696 5481
rect 4602 5427 4608 5428
rect 4602 5423 4603 5427
rect 4607 5423 4608 5427
rect 4602 5422 4608 5423
rect 4692 5395 4694 5480
rect 4820 5436 4822 5494
rect 4898 5485 4904 5486
rect 4898 5481 4899 5485
rect 4903 5481 4904 5485
rect 4898 5480 4904 5481
rect 4818 5435 4824 5436
rect 4818 5431 4819 5435
rect 4823 5431 4824 5435
rect 4818 5430 4824 5431
rect 4900 5395 4902 5480
rect 4603 5394 4607 5395
rect 4603 5389 4607 5390
rect 4691 5394 4695 5395
rect 4691 5389 4695 5390
rect 4779 5394 4783 5395
rect 4779 5389 4783 5390
rect 4899 5394 4903 5395
rect 4899 5389 4903 5390
rect 4963 5394 4967 5395
rect 4963 5389 4967 5390
rect 4604 5328 4606 5389
rect 4722 5383 4728 5384
rect 4722 5379 4723 5383
rect 4727 5379 4728 5383
rect 4722 5378 4728 5379
rect 4698 5375 4704 5376
rect 4698 5371 4699 5375
rect 4703 5371 4704 5375
rect 4698 5370 4704 5371
rect 4602 5327 4608 5328
rect 4602 5323 4603 5327
rect 4607 5323 4608 5327
rect 4602 5322 4608 5323
rect 4630 5312 4636 5313
rect 3838 5311 3844 5312
rect 3838 5307 3839 5311
rect 3843 5307 3844 5311
rect 3886 5308 3887 5312
rect 3891 5308 3892 5312
rect 3886 5307 3892 5308
rect 4002 5311 4008 5312
rect 4002 5307 4003 5311
rect 4007 5307 4008 5311
rect 4022 5308 4023 5312
rect 4027 5308 4028 5312
rect 4022 5307 4028 5308
rect 4138 5311 4144 5312
rect 4138 5307 4139 5311
rect 4143 5307 4144 5311
rect 4158 5308 4159 5312
rect 4163 5308 4164 5312
rect 4158 5307 4164 5308
rect 4282 5311 4288 5312
rect 4282 5307 4283 5311
rect 4287 5307 4288 5311
rect 4302 5308 4303 5312
rect 4307 5308 4308 5312
rect 4302 5307 4308 5308
rect 4394 5311 4400 5312
rect 4394 5307 4395 5311
rect 4399 5307 4400 5311
rect 4462 5308 4463 5312
rect 4467 5308 4468 5312
rect 4462 5307 4468 5308
rect 4558 5311 4564 5312
rect 4558 5307 4559 5311
rect 4563 5307 4564 5311
rect 4630 5308 4631 5312
rect 4635 5308 4636 5312
rect 4630 5307 4636 5308
rect 3838 5306 3844 5307
rect 3798 5288 3804 5289
rect 3798 5284 3799 5288
rect 3803 5284 3804 5288
rect 3798 5283 3804 5284
rect 3840 5279 3842 5306
rect 3888 5279 3890 5307
rect 4002 5306 4008 5307
rect 4024 5279 4026 5307
rect 4138 5306 4144 5307
rect 4066 5279 4072 5280
rect 4160 5279 4162 5307
rect 4282 5306 4288 5307
rect 4304 5279 4306 5307
rect 4394 5306 4400 5307
rect 4396 5293 4398 5306
rect 4392 5291 4398 5293
rect 4392 5280 4394 5291
rect 4390 5279 4396 5280
rect 4464 5279 4466 5307
rect 4558 5306 4564 5307
rect 4632 5279 4634 5307
rect 3839 5278 3843 5279
rect 3839 5273 3843 5274
rect 3887 5278 3891 5279
rect 3887 5273 3891 5274
rect 3999 5278 4003 5279
rect 3999 5273 4003 5274
rect 4023 5278 4027 5279
rect 4066 5275 4067 5279
rect 4071 5275 4072 5279
rect 4066 5274 4072 5275
rect 4159 5278 4163 5279
rect 4023 5273 4027 5274
rect 3786 5271 3792 5272
rect 3786 5267 3787 5271
rect 3791 5267 3792 5271
rect 3786 5266 3792 5267
rect 3798 5271 3804 5272
rect 3798 5267 3799 5271
rect 3803 5267 3804 5271
rect 3798 5266 3804 5267
rect 3800 5243 3802 5266
rect 3840 5250 3842 5273
rect 3838 5249 3844 5250
rect 4000 5249 4002 5273
rect 3838 5245 3839 5249
rect 3843 5245 3844 5249
rect 3838 5244 3844 5245
rect 3998 5248 4004 5249
rect 3998 5244 3999 5248
rect 4003 5244 4004 5248
rect 3998 5243 4004 5244
rect 3799 5242 3803 5243
rect 3799 5237 3803 5238
rect 3800 5214 3802 5237
rect 3970 5233 3976 5234
rect 3838 5232 3844 5233
rect 3838 5228 3839 5232
rect 3843 5228 3844 5232
rect 3970 5229 3971 5233
rect 3975 5229 3976 5233
rect 3970 5228 3976 5229
rect 3838 5227 3844 5228
rect 3798 5213 3804 5214
rect 2238 5208 2239 5212
rect 2243 5208 2244 5212
rect 2238 5207 2244 5208
rect 2334 5211 2340 5212
rect 2334 5207 2335 5211
rect 2339 5207 2340 5211
rect 2590 5208 2591 5212
rect 2595 5208 2596 5212
rect 2590 5207 2596 5208
rect 2866 5211 2872 5212
rect 2866 5207 2867 5211
rect 2871 5207 2872 5211
rect 2942 5208 2943 5212
rect 2947 5208 2948 5212
rect 2942 5207 2948 5208
rect 3038 5211 3044 5212
rect 3038 5207 3039 5211
rect 3043 5207 3044 5211
rect 3302 5208 3303 5212
rect 3307 5208 3308 5212
rect 3302 5207 3308 5208
rect 3594 5211 3600 5212
rect 3594 5207 3595 5211
rect 3599 5207 3600 5211
rect 3662 5208 3663 5212
rect 3667 5208 3668 5212
rect 3662 5207 3668 5208
rect 3758 5211 3764 5212
rect 3758 5207 3759 5211
rect 3763 5207 3764 5211
rect 3798 5209 3799 5213
rect 3803 5209 3804 5213
rect 3798 5208 3804 5209
rect 2334 5206 2340 5207
rect 2866 5206 2872 5207
rect 3038 5206 3044 5207
rect 3594 5206 3600 5207
rect 3758 5206 3764 5207
rect 2210 5197 2216 5198
rect 2210 5193 2211 5197
rect 2215 5193 2216 5197
rect 2210 5192 2216 5193
rect 2198 5147 2204 5148
rect 2198 5143 2199 5147
rect 2203 5143 2204 5147
rect 2198 5142 2204 5143
rect 2212 5131 2214 5192
rect 1934 5128 1940 5129
rect 1975 5130 1979 5131
rect 1910 5126 1916 5127
rect 1786 5117 1792 5118
rect 1786 5113 1787 5117
rect 1791 5113 1792 5117
rect 1786 5112 1792 5113
rect 1746 5067 1752 5068
rect 1746 5063 1747 5067
rect 1751 5063 1752 5067
rect 1746 5062 1752 5063
rect 1788 5047 1790 5112
rect 1912 5060 1914 5126
rect 1975 5125 1979 5126
rect 2211 5130 2215 5131
rect 2211 5125 2215 5126
rect 2267 5130 2271 5131
rect 2267 5125 2271 5126
rect 1934 5116 1940 5117
rect 1934 5112 1935 5116
rect 1939 5112 1940 5116
rect 1934 5111 1940 5112
rect 1910 5059 1916 5060
rect 1910 5055 1911 5059
rect 1915 5055 1916 5059
rect 1910 5054 1916 5055
rect 1936 5047 1938 5111
rect 1976 5065 1978 5125
rect 1974 5064 1980 5065
rect 2268 5064 2270 5125
rect 2336 5116 2338 5206
rect 2562 5197 2568 5198
rect 2562 5193 2563 5197
rect 2567 5193 2568 5197
rect 2562 5192 2568 5193
rect 2914 5197 2920 5198
rect 2914 5193 2915 5197
rect 2919 5193 2920 5197
rect 2914 5192 2920 5193
rect 2564 5131 2566 5192
rect 2638 5147 2644 5148
rect 2638 5143 2639 5147
rect 2643 5143 2644 5147
rect 2638 5142 2644 5143
rect 2515 5130 2519 5131
rect 2515 5125 2519 5126
rect 2563 5130 2567 5131
rect 2563 5125 2567 5126
rect 2334 5115 2340 5116
rect 2334 5111 2335 5115
rect 2339 5111 2340 5115
rect 2334 5110 2340 5111
rect 2516 5064 2518 5125
rect 1974 5060 1975 5064
rect 1979 5060 1980 5064
rect 1974 5059 1980 5060
rect 2266 5063 2272 5064
rect 2266 5059 2267 5063
rect 2271 5059 2272 5063
rect 2266 5058 2272 5059
rect 2514 5063 2520 5064
rect 2514 5059 2515 5063
rect 2519 5059 2520 5063
rect 2514 5058 2520 5059
rect 2294 5048 2300 5049
rect 2542 5048 2548 5049
rect 2640 5048 2642 5142
rect 2916 5131 2918 5192
rect 3040 5148 3042 5206
rect 3274 5197 3280 5198
rect 3274 5193 3275 5197
rect 3279 5193 3280 5197
rect 3274 5192 3280 5193
rect 3038 5147 3044 5148
rect 3038 5143 3039 5147
rect 3043 5143 3044 5147
rect 3038 5142 3044 5143
rect 3114 5139 3120 5140
rect 3114 5135 3115 5139
rect 3119 5135 3120 5139
rect 3114 5134 3120 5135
rect 2755 5130 2759 5131
rect 2755 5125 2759 5126
rect 2915 5130 2919 5131
rect 2915 5125 2919 5126
rect 2995 5130 2999 5131
rect 2995 5125 2999 5126
rect 2756 5064 2758 5125
rect 2838 5115 2844 5116
rect 2838 5111 2839 5115
rect 2843 5111 2844 5115
rect 2838 5110 2844 5111
rect 2754 5063 2760 5064
rect 2754 5059 2755 5063
rect 2759 5059 2760 5063
rect 2754 5058 2760 5059
rect 2782 5048 2788 5049
rect 1974 5047 1980 5048
rect 1787 5046 1791 5047
rect 1787 5041 1791 5042
rect 1935 5046 1939 5047
rect 1974 5043 1975 5047
rect 1979 5043 1980 5047
rect 2294 5044 2295 5048
rect 2299 5044 2300 5048
rect 2294 5043 2300 5044
rect 2390 5047 2396 5048
rect 2390 5043 2391 5047
rect 2395 5043 2396 5047
rect 2542 5044 2543 5048
rect 2547 5044 2548 5048
rect 2542 5043 2548 5044
rect 2638 5047 2644 5048
rect 2638 5043 2639 5047
rect 2643 5043 2644 5047
rect 2782 5044 2783 5048
rect 2787 5044 2788 5048
rect 2782 5043 2788 5044
rect 1974 5042 1980 5043
rect 1935 5041 1939 5042
rect 1726 5031 1732 5032
rect 1726 5027 1727 5031
rect 1731 5027 1732 5031
rect 1726 5026 1732 5027
rect 1782 4995 1788 4996
rect 1782 4991 1783 4995
rect 1787 4991 1788 4995
rect 1782 4990 1788 4991
rect 1370 4979 1376 4980
rect 1370 4975 1371 4979
rect 1375 4975 1376 4979
rect 1370 4974 1376 4975
rect 1658 4979 1664 4980
rect 1658 4975 1659 4979
rect 1663 4975 1664 4979
rect 1658 4974 1664 4975
rect 1330 4971 1336 4972
rect 1330 4967 1331 4971
rect 1335 4967 1336 4971
rect 1330 4966 1336 4967
rect 1398 4964 1404 4965
rect 110 4963 116 4964
rect 110 4959 111 4963
rect 115 4959 116 4963
rect 158 4960 159 4964
rect 163 4960 164 4964
rect 158 4959 164 4960
rect 330 4963 336 4964
rect 330 4959 331 4963
rect 335 4959 336 4963
rect 350 4960 351 4964
rect 355 4960 356 4964
rect 350 4959 356 4960
rect 446 4963 452 4964
rect 446 4959 447 4963
rect 451 4959 452 4963
rect 582 4960 583 4964
rect 587 4960 588 4964
rect 582 4959 588 4960
rect 818 4963 824 4964
rect 818 4959 819 4963
rect 823 4959 824 4963
rect 838 4960 839 4964
rect 843 4960 844 4964
rect 838 4959 844 4960
rect 1090 4963 1096 4964
rect 1090 4959 1091 4963
rect 1095 4959 1096 4963
rect 1110 4960 1111 4964
rect 1115 4960 1116 4964
rect 1110 4959 1116 4960
rect 1206 4963 1212 4964
rect 1206 4959 1207 4963
rect 1211 4959 1212 4963
rect 1398 4960 1399 4964
rect 1403 4960 1404 4964
rect 1398 4959 1404 4960
rect 1686 4964 1692 4965
rect 1784 4964 1786 4990
rect 1936 4981 1938 5041
rect 1976 4987 1978 5042
rect 2296 4987 2298 5043
rect 2390 5042 2396 5043
rect 1975 4986 1979 4987
rect 1975 4981 1979 4982
rect 2183 4986 2187 4987
rect 2183 4981 2187 4982
rect 2295 4986 2299 4987
rect 2295 4981 2299 4982
rect 2319 4986 2323 4987
rect 2319 4981 2323 4982
rect 1934 4980 1940 4981
rect 1934 4976 1935 4980
rect 1939 4976 1940 4980
rect 1934 4975 1940 4976
rect 1686 4960 1687 4964
rect 1691 4960 1692 4964
rect 1686 4959 1692 4960
rect 1782 4963 1788 4964
rect 1782 4959 1783 4963
rect 1787 4959 1788 4963
rect 110 4958 116 4959
rect 112 4911 114 4958
rect 160 4911 162 4959
rect 330 4958 336 4959
rect 352 4911 354 4959
rect 446 4958 452 4959
rect 111 4910 115 4911
rect 111 4905 115 4906
rect 159 4910 163 4911
rect 159 4905 163 4906
rect 295 4910 299 4911
rect 295 4905 299 4906
rect 351 4910 355 4911
rect 351 4905 355 4906
rect 431 4910 435 4911
rect 431 4905 435 4906
rect 112 4882 114 4905
rect 110 4881 116 4882
rect 160 4881 162 4905
rect 296 4881 298 4905
rect 432 4881 434 4905
rect 110 4877 111 4881
rect 115 4877 116 4881
rect 110 4876 116 4877
rect 158 4880 164 4881
rect 294 4880 300 4881
rect 430 4880 436 4881
rect 158 4876 159 4880
rect 163 4876 164 4880
rect 158 4875 164 4876
rect 250 4879 256 4880
rect 250 4875 251 4879
rect 255 4875 256 4879
rect 294 4876 295 4880
rect 299 4876 300 4880
rect 294 4875 300 4876
rect 386 4879 392 4880
rect 386 4875 387 4879
rect 391 4875 392 4879
rect 430 4876 431 4880
rect 435 4876 436 4880
rect 430 4875 436 4876
rect 250 4874 256 4875
rect 386 4874 392 4875
rect 130 4865 136 4866
rect 110 4864 116 4865
rect 110 4860 111 4864
rect 115 4860 116 4864
rect 130 4861 131 4865
rect 135 4861 136 4865
rect 130 4860 136 4861
rect 110 4859 116 4860
rect 112 4787 114 4859
rect 132 4787 134 4860
rect 111 4786 115 4787
rect 111 4781 115 4782
rect 131 4786 135 4787
rect 131 4781 135 4782
rect 112 4721 114 4781
rect 110 4720 116 4721
rect 132 4720 134 4781
rect 252 4772 254 4874
rect 266 4865 272 4866
rect 266 4861 267 4865
rect 271 4861 272 4865
rect 266 4860 272 4861
rect 268 4787 270 4860
rect 388 4808 390 4874
rect 402 4865 408 4866
rect 402 4861 403 4865
rect 407 4861 408 4865
rect 402 4860 408 4861
rect 386 4807 392 4808
rect 386 4803 387 4807
rect 391 4803 392 4807
rect 386 4802 392 4803
rect 404 4787 406 4860
rect 448 4816 450 4958
rect 584 4911 586 4959
rect 818 4958 824 4959
rect 840 4911 842 4959
rect 1090 4958 1096 4959
rect 1112 4911 1114 4959
rect 1206 4958 1212 4959
rect 1400 4911 1402 4959
rect 1688 4911 1690 4959
rect 1782 4958 1788 4959
rect 1934 4963 1940 4964
rect 1934 4959 1935 4963
rect 1939 4959 1940 4963
rect 1934 4958 1940 4959
rect 1976 4958 1978 4981
rect 1936 4911 1938 4958
rect 1974 4957 1980 4958
rect 2184 4957 2186 4981
rect 2320 4957 2322 4981
rect 1974 4953 1975 4957
rect 1979 4953 1980 4957
rect 1974 4952 1980 4953
rect 2182 4956 2188 4957
rect 2318 4956 2324 4957
rect 2182 4952 2183 4956
rect 2187 4952 2188 4956
rect 2182 4951 2188 4952
rect 2282 4955 2288 4956
rect 2282 4951 2283 4955
rect 2287 4951 2288 4955
rect 2318 4952 2319 4956
rect 2323 4952 2324 4956
rect 2318 4951 2324 4952
rect 2282 4950 2288 4951
rect 2154 4941 2160 4942
rect 1974 4940 1980 4941
rect 1974 4936 1975 4940
rect 1979 4936 1980 4940
rect 2154 4937 2155 4941
rect 2159 4937 2160 4941
rect 2154 4936 2160 4937
rect 1974 4935 1980 4936
rect 567 4910 571 4911
rect 567 4905 571 4906
rect 583 4910 587 4911
rect 583 4905 587 4906
rect 703 4910 707 4911
rect 703 4905 707 4906
rect 839 4910 843 4911
rect 839 4905 843 4906
rect 1111 4910 1115 4911
rect 1111 4905 1115 4906
rect 1399 4910 1403 4911
rect 1399 4905 1403 4906
rect 1687 4910 1691 4911
rect 1687 4905 1691 4906
rect 1935 4910 1939 4911
rect 1935 4905 1939 4906
rect 568 4881 570 4905
rect 704 4881 706 4905
rect 1936 4882 1938 4905
rect 1934 4881 1940 4882
rect 566 4880 572 4881
rect 702 4880 708 4881
rect 530 4879 536 4880
rect 530 4875 531 4879
rect 535 4875 536 4879
rect 566 4876 567 4880
rect 571 4876 572 4880
rect 566 4875 572 4876
rect 666 4879 672 4880
rect 666 4875 667 4879
rect 671 4875 672 4879
rect 702 4876 703 4880
rect 707 4876 708 4880
rect 702 4875 708 4876
rect 798 4879 804 4880
rect 798 4875 799 4879
rect 803 4875 804 4879
rect 1934 4877 1935 4881
rect 1939 4877 1940 4881
rect 1934 4876 1940 4877
rect 530 4874 536 4875
rect 666 4874 672 4875
rect 798 4874 804 4875
rect 532 4816 534 4874
rect 538 4865 544 4866
rect 538 4861 539 4865
rect 543 4861 544 4865
rect 538 4860 544 4861
rect 446 4815 452 4816
rect 446 4811 447 4815
rect 451 4811 452 4815
rect 446 4810 452 4811
rect 530 4815 536 4816
rect 530 4811 531 4815
rect 535 4811 536 4815
rect 530 4810 536 4811
rect 540 4787 542 4860
rect 668 4816 670 4874
rect 674 4865 680 4866
rect 674 4861 675 4865
rect 679 4861 680 4865
rect 674 4860 680 4861
rect 666 4815 672 4816
rect 666 4811 667 4815
rect 671 4811 672 4815
rect 666 4810 672 4811
rect 676 4787 678 4860
rect 800 4808 802 4874
rect 1976 4867 1978 4935
rect 2156 4867 2158 4936
rect 2284 4892 2286 4950
rect 2290 4941 2296 4942
rect 2290 4937 2291 4941
rect 2295 4937 2296 4941
rect 2290 4936 2296 4937
rect 2282 4891 2288 4892
rect 2282 4887 2283 4891
rect 2287 4887 2288 4891
rect 2282 4886 2288 4887
rect 2292 4867 2294 4936
rect 2392 4884 2394 5042
rect 2544 4987 2546 5043
rect 2638 5042 2644 5043
rect 2784 4987 2786 5043
rect 2455 4986 2459 4987
rect 2455 4981 2459 4982
rect 2543 4986 2547 4987
rect 2543 4981 2547 4982
rect 2599 4986 2603 4987
rect 2599 4981 2603 4982
rect 2743 4986 2747 4987
rect 2743 4981 2747 4982
rect 2783 4986 2787 4987
rect 2783 4981 2787 4982
rect 2456 4957 2458 4981
rect 2600 4957 2602 4981
rect 2744 4957 2746 4981
rect 2454 4956 2460 4957
rect 2598 4956 2604 4957
rect 2742 4956 2748 4957
rect 2840 4956 2842 5110
rect 2996 5064 2998 5125
rect 2994 5063 3000 5064
rect 2994 5059 2995 5063
rect 2999 5059 3000 5063
rect 2994 5058 3000 5059
rect 3022 5048 3028 5049
rect 3116 5048 3118 5134
rect 3276 5131 3278 5192
rect 3596 5148 3598 5206
rect 3634 5197 3640 5198
rect 3634 5193 3635 5197
rect 3639 5193 3640 5197
rect 3634 5192 3640 5193
rect 3798 5196 3804 5197
rect 3798 5192 3799 5196
rect 3803 5192 3804 5196
rect 3594 5147 3600 5148
rect 3594 5143 3595 5147
rect 3599 5143 3600 5147
rect 3594 5142 3600 5143
rect 3636 5131 3638 5192
rect 3798 5191 3804 5192
rect 3800 5131 3802 5191
rect 3840 5147 3842 5227
rect 3972 5147 3974 5228
rect 4068 5184 4070 5274
rect 4159 5273 4163 5274
rect 4199 5278 4203 5279
rect 4199 5273 4203 5274
rect 4303 5278 4307 5279
rect 4390 5275 4391 5279
rect 4395 5275 4396 5279
rect 4390 5274 4396 5275
rect 4399 5278 4403 5279
rect 4303 5273 4307 5274
rect 4399 5273 4403 5274
rect 4463 5278 4467 5279
rect 4463 5273 4467 5274
rect 4607 5278 4611 5279
rect 4607 5273 4611 5274
rect 4631 5278 4635 5279
rect 4631 5273 4635 5274
rect 4200 5249 4202 5273
rect 4400 5249 4402 5273
rect 4608 5249 4610 5273
rect 4198 5248 4204 5249
rect 4398 5248 4404 5249
rect 4606 5248 4612 5249
rect 4700 5248 4702 5370
rect 4724 5312 4726 5378
rect 4780 5328 4782 5389
rect 4930 5379 4936 5380
rect 4930 5375 4931 5379
rect 4935 5375 4936 5379
rect 4930 5374 4936 5375
rect 4778 5327 4784 5328
rect 4778 5323 4779 5327
rect 4783 5323 4784 5327
rect 4778 5322 4784 5323
rect 4932 5320 4934 5374
rect 4964 5328 4966 5389
rect 5024 5380 5026 5494
rect 5106 5485 5112 5486
rect 5106 5481 5107 5485
rect 5111 5481 5112 5485
rect 5106 5480 5112 5481
rect 5108 5395 5110 5480
rect 5232 5428 5234 5494
rect 5316 5436 5318 5586
rect 5664 5531 5666 5586
rect 5663 5530 5667 5531
rect 5663 5525 5667 5526
rect 5664 5502 5666 5525
rect 5662 5501 5668 5502
rect 5662 5497 5663 5501
rect 5667 5497 5668 5501
rect 5662 5496 5668 5497
rect 5662 5484 5668 5485
rect 5662 5480 5663 5484
rect 5667 5480 5668 5484
rect 5662 5479 5668 5480
rect 5314 5435 5320 5436
rect 5314 5431 5315 5435
rect 5319 5431 5320 5435
rect 5314 5430 5320 5431
rect 5230 5427 5236 5428
rect 5230 5423 5231 5427
rect 5235 5423 5236 5427
rect 5230 5422 5236 5423
rect 5664 5395 5666 5479
rect 5107 5394 5111 5395
rect 5107 5389 5111 5390
rect 5663 5394 5667 5395
rect 5663 5389 5667 5390
rect 5022 5379 5028 5380
rect 5022 5375 5023 5379
rect 5027 5375 5028 5379
rect 5022 5374 5028 5375
rect 5664 5329 5666 5389
rect 5662 5328 5668 5329
rect 4962 5327 4968 5328
rect 4962 5323 4963 5327
rect 4967 5323 4968 5327
rect 5662 5324 5663 5328
rect 5667 5324 5668 5328
rect 5662 5323 5668 5324
rect 4962 5322 4968 5323
rect 4930 5319 4936 5320
rect 4930 5315 4931 5319
rect 4935 5315 4936 5319
rect 4930 5314 4936 5315
rect 4806 5312 4812 5313
rect 4990 5312 4996 5313
rect 4722 5311 4728 5312
rect 4722 5307 4723 5311
rect 4727 5307 4728 5311
rect 4806 5308 4807 5312
rect 4811 5308 4812 5312
rect 4806 5307 4812 5308
rect 4898 5311 4904 5312
rect 4898 5307 4899 5311
rect 4903 5307 4904 5311
rect 4990 5308 4991 5312
rect 4995 5308 4996 5312
rect 4990 5307 4996 5308
rect 5662 5311 5668 5312
rect 5662 5307 5663 5311
rect 5667 5307 5668 5311
rect 4722 5306 4728 5307
rect 4808 5279 4810 5307
rect 4898 5306 4904 5307
rect 4807 5278 4811 5279
rect 4807 5273 4811 5274
rect 4823 5278 4827 5279
rect 4823 5273 4827 5274
rect 4824 5249 4826 5273
rect 4822 5248 4828 5249
rect 4098 5247 4104 5248
rect 4098 5243 4099 5247
rect 4103 5243 4104 5247
rect 4198 5244 4199 5248
rect 4203 5244 4204 5248
rect 4198 5243 4204 5244
rect 4298 5247 4304 5248
rect 4298 5243 4299 5247
rect 4303 5243 4304 5247
rect 4398 5244 4399 5248
rect 4403 5244 4404 5248
rect 4398 5243 4404 5244
rect 4490 5247 4496 5248
rect 4490 5243 4491 5247
rect 4495 5243 4496 5247
rect 4606 5244 4607 5248
rect 4611 5244 4612 5248
rect 4606 5243 4612 5244
rect 4698 5247 4704 5248
rect 4698 5243 4699 5247
rect 4703 5243 4704 5247
rect 4822 5244 4823 5248
rect 4827 5244 4828 5248
rect 4822 5243 4828 5244
rect 4098 5242 4104 5243
rect 4298 5242 4304 5243
rect 4490 5242 4496 5243
rect 4698 5242 4704 5243
rect 4100 5184 4102 5242
rect 4170 5233 4176 5234
rect 4170 5229 4171 5233
rect 4175 5229 4176 5233
rect 4170 5228 4176 5229
rect 4066 5183 4072 5184
rect 4066 5179 4067 5183
rect 4071 5179 4072 5183
rect 4066 5178 4072 5179
rect 4098 5183 4104 5184
rect 4098 5179 4099 5183
rect 4103 5179 4104 5183
rect 4098 5178 4104 5179
rect 4172 5147 4174 5228
rect 4300 5184 4302 5242
rect 4370 5233 4376 5234
rect 4370 5229 4371 5233
rect 4375 5229 4376 5233
rect 4370 5228 4376 5229
rect 4298 5183 4304 5184
rect 4298 5179 4299 5183
rect 4303 5179 4304 5183
rect 4298 5178 4304 5179
rect 4372 5147 4374 5228
rect 3839 5146 3843 5147
rect 3839 5141 3843 5142
rect 3971 5146 3975 5147
rect 3971 5141 3975 5142
rect 4099 5146 4103 5147
rect 4099 5141 4103 5142
rect 4171 5146 4175 5147
rect 4171 5141 4175 5142
rect 4347 5146 4351 5147
rect 4347 5141 4351 5142
rect 4371 5146 4375 5147
rect 4371 5141 4375 5142
rect 3235 5130 3239 5131
rect 3235 5125 3239 5126
rect 3275 5130 3279 5131
rect 3275 5125 3279 5126
rect 3475 5130 3479 5131
rect 3475 5125 3479 5126
rect 3635 5130 3639 5131
rect 3635 5125 3639 5126
rect 3799 5130 3803 5131
rect 3799 5125 3803 5126
rect 3226 5115 3232 5116
rect 3226 5111 3227 5115
rect 3231 5111 3232 5115
rect 3226 5110 3232 5111
rect 3228 5056 3230 5110
rect 3236 5064 3238 5125
rect 3476 5064 3478 5125
rect 3598 5119 3604 5120
rect 3598 5115 3599 5119
rect 3603 5115 3604 5119
rect 3598 5114 3604 5115
rect 3482 5111 3488 5112
rect 3482 5107 3483 5111
rect 3487 5107 3488 5111
rect 3482 5106 3488 5107
rect 3234 5063 3240 5064
rect 3234 5059 3235 5063
rect 3239 5059 3240 5063
rect 3234 5058 3240 5059
rect 3474 5063 3480 5064
rect 3474 5059 3475 5063
rect 3479 5059 3480 5063
rect 3474 5058 3480 5059
rect 3226 5055 3232 5056
rect 3226 5051 3227 5055
rect 3231 5051 3232 5055
rect 3226 5050 3232 5051
rect 3262 5048 3268 5049
rect 3022 5044 3023 5048
rect 3027 5044 3028 5048
rect 3022 5043 3028 5044
rect 3114 5047 3120 5048
rect 3114 5043 3115 5047
rect 3119 5043 3120 5047
rect 3262 5044 3263 5048
rect 3267 5044 3268 5048
rect 3262 5043 3268 5044
rect 3024 4987 3026 5043
rect 3114 5042 3120 5043
rect 3264 4987 3266 5043
rect 2895 4986 2899 4987
rect 2895 4981 2899 4982
rect 3023 4986 3027 4987
rect 3023 4981 3027 4982
rect 3047 4986 3051 4987
rect 3047 4981 3051 4982
rect 3199 4986 3203 4987
rect 3199 4981 3203 4982
rect 3263 4986 3267 4987
rect 3263 4981 3267 4982
rect 3351 4986 3355 4987
rect 3351 4981 3355 4982
rect 2896 4957 2898 4981
rect 3048 4957 3050 4981
rect 3200 4957 3202 4981
rect 3352 4957 3354 4981
rect 2894 4956 2900 4957
rect 3046 4956 3052 4957
rect 3198 4956 3204 4957
rect 3350 4956 3356 4957
rect 3484 4956 3486 5106
rect 3502 5048 3508 5049
rect 3600 5048 3602 5114
rect 3800 5065 3802 5125
rect 3840 5081 3842 5141
rect 3838 5080 3844 5081
rect 4100 5080 4102 5141
rect 4348 5080 4350 5141
rect 4492 5132 4494 5242
rect 4578 5233 4584 5234
rect 4578 5229 4579 5233
rect 4583 5229 4584 5233
rect 4578 5228 4584 5229
rect 4794 5233 4800 5234
rect 4794 5229 4795 5233
rect 4799 5229 4800 5233
rect 4794 5228 4800 5229
rect 4580 5147 4582 5228
rect 4714 5183 4720 5184
rect 4714 5179 4715 5183
rect 4719 5179 4720 5183
rect 4714 5178 4720 5179
rect 4579 5146 4583 5147
rect 4579 5141 4583 5142
rect 4595 5146 4599 5147
rect 4595 5141 4599 5142
rect 4490 5131 4496 5132
rect 4490 5127 4491 5131
rect 4495 5127 4496 5131
rect 4490 5126 4496 5127
rect 4596 5080 4598 5141
rect 4602 5127 4608 5128
rect 4602 5123 4603 5127
rect 4607 5123 4608 5127
rect 4602 5122 4608 5123
rect 3838 5076 3839 5080
rect 3843 5076 3844 5080
rect 3838 5075 3844 5076
rect 4098 5079 4104 5080
rect 4098 5075 4099 5079
rect 4103 5075 4104 5079
rect 4098 5074 4104 5075
rect 4346 5079 4352 5080
rect 4346 5075 4347 5079
rect 4351 5075 4352 5079
rect 4346 5074 4352 5075
rect 4594 5079 4600 5080
rect 4594 5075 4595 5079
rect 4599 5075 4600 5079
rect 4594 5074 4600 5075
rect 3798 5064 3804 5065
rect 4126 5064 4132 5065
rect 4374 5064 4380 5065
rect 3798 5060 3799 5064
rect 3803 5060 3804 5064
rect 3798 5059 3804 5060
rect 3838 5063 3844 5064
rect 3838 5059 3839 5063
rect 3843 5059 3844 5063
rect 4126 5060 4127 5064
rect 4131 5060 4132 5064
rect 4126 5059 4132 5060
rect 4222 5063 4228 5064
rect 4222 5059 4223 5063
rect 4227 5059 4228 5063
rect 4374 5060 4375 5064
rect 4379 5060 4380 5064
rect 4374 5059 4380 5060
rect 3838 5058 3844 5059
rect 3502 5044 3503 5048
rect 3507 5044 3508 5048
rect 3502 5043 3508 5044
rect 3598 5047 3604 5048
rect 3598 5043 3599 5047
rect 3603 5043 3604 5047
rect 3504 4987 3506 5043
rect 3598 5042 3604 5043
rect 3798 5047 3804 5048
rect 3798 5043 3799 5047
rect 3803 5043 3804 5047
rect 3798 5042 3804 5043
rect 3800 4987 3802 5042
rect 3840 5019 3842 5058
rect 4128 5019 4130 5059
rect 4216 5058 4228 5059
rect 4216 5057 4226 5058
rect 3839 5018 3843 5019
rect 3839 5013 3843 5014
rect 3983 5018 3987 5019
rect 3983 5013 3987 5014
rect 4127 5018 4131 5019
rect 4127 5013 4131 5014
rect 3840 4990 3842 5013
rect 3838 4989 3844 4990
rect 3984 4989 3986 5013
rect 3503 4986 3507 4987
rect 3503 4981 3507 4982
rect 3799 4986 3803 4987
rect 3838 4985 3839 4989
rect 3843 4985 3844 4989
rect 3838 4984 3844 4985
rect 3982 4988 3988 4989
rect 3982 4984 3983 4988
rect 3987 4984 3988 4988
rect 3982 4983 3988 4984
rect 4082 4987 4088 4988
rect 4082 4983 4083 4987
rect 4087 4983 4088 4987
rect 4082 4982 4088 4983
rect 3799 4981 3803 4982
rect 3800 4958 3802 4981
rect 3954 4973 3960 4974
rect 3838 4972 3844 4973
rect 3838 4968 3839 4972
rect 3843 4968 3844 4972
rect 3954 4969 3955 4973
rect 3959 4969 3960 4973
rect 3954 4968 3960 4969
rect 3838 4967 3844 4968
rect 3798 4957 3804 4958
rect 2418 4955 2424 4956
rect 2418 4951 2419 4955
rect 2423 4951 2424 4955
rect 2454 4952 2455 4956
rect 2459 4952 2460 4956
rect 2454 4951 2460 4952
rect 2554 4955 2560 4956
rect 2554 4951 2555 4955
rect 2559 4951 2560 4955
rect 2598 4952 2599 4956
rect 2603 4952 2604 4956
rect 2598 4951 2604 4952
rect 2690 4955 2696 4956
rect 2690 4951 2691 4955
rect 2695 4951 2696 4955
rect 2742 4952 2743 4956
rect 2747 4952 2748 4956
rect 2742 4951 2748 4952
rect 2838 4955 2844 4956
rect 2838 4951 2839 4955
rect 2843 4951 2844 4955
rect 2894 4952 2895 4956
rect 2899 4952 2900 4956
rect 2894 4951 2900 4952
rect 2986 4955 2992 4956
rect 2986 4951 2987 4955
rect 2991 4951 2992 4955
rect 3046 4952 3047 4956
rect 3051 4952 3052 4956
rect 3046 4951 3052 4952
rect 3142 4955 3148 4956
rect 3142 4951 3143 4955
rect 3147 4951 3148 4955
rect 3198 4952 3199 4956
rect 3203 4952 3204 4956
rect 3198 4951 3204 4952
rect 3294 4955 3300 4956
rect 3294 4951 3295 4955
rect 3299 4951 3300 4955
rect 3350 4952 3351 4956
rect 3355 4952 3356 4956
rect 3350 4951 3356 4952
rect 3482 4955 3488 4956
rect 3482 4951 3483 4955
rect 3487 4951 3488 4955
rect 3798 4953 3799 4957
rect 3803 4953 3804 4957
rect 3798 4952 3804 4953
rect 2418 4950 2424 4951
rect 2554 4950 2560 4951
rect 2690 4950 2696 4951
rect 2838 4950 2844 4951
rect 2986 4950 2992 4951
rect 3142 4950 3148 4951
rect 3294 4950 3300 4951
rect 3482 4950 3488 4951
rect 2420 4892 2422 4950
rect 2426 4941 2432 4942
rect 2426 4937 2427 4941
rect 2431 4937 2432 4941
rect 2426 4936 2432 4937
rect 2418 4891 2424 4892
rect 2418 4887 2419 4891
rect 2423 4887 2424 4891
rect 2418 4886 2424 4887
rect 2390 4883 2396 4884
rect 2390 4879 2391 4883
rect 2395 4879 2396 4883
rect 2390 4878 2396 4879
rect 2428 4867 2430 4936
rect 2556 4892 2558 4950
rect 2570 4941 2576 4942
rect 2570 4937 2571 4941
rect 2575 4937 2576 4941
rect 2570 4936 2576 4937
rect 2554 4891 2560 4892
rect 2554 4887 2555 4891
rect 2559 4887 2560 4891
rect 2554 4886 2560 4887
rect 2572 4867 2574 4936
rect 1975 4866 1979 4867
rect 1934 4864 1940 4865
rect 1934 4860 1935 4864
rect 1939 4860 1940 4864
rect 1975 4861 1979 4862
rect 2155 4866 2159 4867
rect 2155 4861 2159 4862
rect 2291 4866 2295 4867
rect 2291 4861 2295 4862
rect 2427 4866 2431 4867
rect 2427 4861 2431 4862
rect 2571 4866 2575 4867
rect 2571 4861 2575 4862
rect 1934 4859 1940 4860
rect 798 4807 804 4808
rect 798 4803 799 4807
rect 803 4803 804 4807
rect 798 4802 804 4803
rect 1936 4787 1938 4859
rect 1976 4801 1978 4861
rect 1974 4800 1980 4801
rect 2428 4800 2430 4861
rect 2572 4800 2574 4861
rect 2692 4856 2694 4950
rect 2714 4941 2720 4942
rect 2714 4937 2715 4941
rect 2719 4937 2720 4941
rect 2714 4936 2720 4937
rect 2866 4941 2872 4942
rect 2866 4937 2867 4941
rect 2871 4937 2872 4941
rect 2866 4936 2872 4937
rect 2716 4867 2718 4936
rect 2850 4891 2856 4892
rect 2850 4887 2851 4891
rect 2855 4887 2856 4891
rect 2850 4886 2856 4887
rect 2715 4866 2719 4867
rect 2715 4861 2719 4862
rect 2723 4866 2727 4867
rect 2723 4861 2727 4862
rect 2690 4855 2696 4856
rect 2690 4851 2691 4855
rect 2695 4851 2696 4855
rect 2690 4850 2696 4851
rect 2578 4847 2584 4848
rect 2578 4843 2579 4847
rect 2583 4843 2584 4847
rect 2578 4842 2584 4843
rect 1974 4796 1975 4800
rect 1979 4796 1980 4800
rect 1974 4795 1980 4796
rect 2426 4799 2432 4800
rect 2426 4795 2427 4799
rect 2431 4795 2432 4799
rect 2426 4794 2432 4795
rect 2570 4799 2576 4800
rect 2570 4795 2571 4799
rect 2575 4795 2576 4799
rect 2570 4794 2576 4795
rect 267 4786 271 4787
rect 267 4781 271 4782
rect 403 4786 407 4787
rect 403 4781 407 4782
rect 539 4786 543 4787
rect 539 4781 543 4782
rect 675 4786 679 4787
rect 675 4781 679 4782
rect 1935 4786 1939 4787
rect 2454 4784 2460 4785
rect 2580 4784 2582 4842
rect 2724 4800 2726 4861
rect 2730 4847 2736 4848
rect 2730 4843 2731 4847
rect 2735 4843 2736 4847
rect 2730 4842 2736 4843
rect 2722 4799 2728 4800
rect 2722 4795 2723 4799
rect 2727 4795 2728 4799
rect 2722 4794 2728 4795
rect 2598 4784 2604 4785
rect 2732 4784 2734 4842
rect 2750 4784 2756 4785
rect 2852 4784 2854 4886
rect 2868 4867 2870 4936
rect 2988 4884 2990 4950
rect 3018 4941 3024 4942
rect 3018 4937 3019 4941
rect 3023 4937 3024 4941
rect 3018 4936 3024 4937
rect 3002 4891 3008 4892
rect 3002 4887 3003 4891
rect 3007 4887 3008 4891
rect 3002 4886 3008 4887
rect 2986 4883 2992 4884
rect 2986 4879 2987 4883
rect 2991 4879 2992 4883
rect 2986 4878 2992 4879
rect 2867 4866 2871 4867
rect 2867 4861 2871 4862
rect 2875 4866 2879 4867
rect 2875 4861 2879 4862
rect 2876 4800 2878 4861
rect 2874 4799 2880 4800
rect 2874 4795 2875 4799
rect 2879 4795 2880 4799
rect 2874 4794 2880 4795
rect 2902 4784 2908 4785
rect 3004 4784 3006 4886
rect 3020 4867 3022 4936
rect 3144 4892 3146 4950
rect 3170 4941 3176 4942
rect 3170 4937 3171 4941
rect 3175 4937 3176 4941
rect 3170 4936 3176 4937
rect 3142 4891 3148 4892
rect 3142 4887 3143 4891
rect 3147 4887 3148 4891
rect 3142 4886 3148 4887
rect 3172 4867 3174 4936
rect 3296 4892 3298 4950
rect 3322 4941 3328 4942
rect 3322 4937 3323 4941
rect 3327 4937 3328 4941
rect 3322 4936 3328 4937
rect 3798 4940 3804 4941
rect 3798 4936 3799 4940
rect 3803 4936 3804 4940
rect 3294 4891 3300 4892
rect 3294 4887 3295 4891
rect 3299 4887 3300 4891
rect 3294 4886 3300 4887
rect 3324 4867 3326 4936
rect 3798 4935 3804 4936
rect 3800 4867 3802 4935
rect 3840 4883 3842 4967
rect 3956 4883 3958 4968
rect 3839 4882 3843 4883
rect 3839 4877 3843 4878
rect 3859 4882 3863 4883
rect 3859 4877 3863 4878
rect 3955 4882 3959 4883
rect 3955 4877 3959 4878
rect 4075 4882 4079 4883
rect 4075 4877 4079 4878
rect 3019 4866 3023 4867
rect 3019 4861 3023 4862
rect 3027 4866 3031 4867
rect 3027 4861 3031 4862
rect 3171 4866 3175 4867
rect 3171 4861 3175 4862
rect 3179 4866 3183 4867
rect 3179 4861 3183 4862
rect 3323 4866 3327 4867
rect 3323 4861 3327 4862
rect 3799 4866 3803 4867
rect 3799 4861 3803 4862
rect 3018 4851 3024 4852
rect 3018 4847 3019 4851
rect 3023 4847 3024 4851
rect 3018 4846 3024 4847
rect 3020 4792 3022 4846
rect 3028 4800 3030 4861
rect 3180 4800 3182 4861
rect 3302 4855 3308 4856
rect 3302 4851 3303 4855
rect 3307 4851 3308 4855
rect 3302 4850 3308 4851
rect 3026 4799 3032 4800
rect 3026 4795 3027 4799
rect 3031 4795 3032 4799
rect 3026 4794 3032 4795
rect 3178 4799 3184 4800
rect 3178 4795 3179 4799
rect 3183 4795 3184 4799
rect 3178 4794 3184 4795
rect 3018 4791 3024 4792
rect 3018 4787 3019 4791
rect 3023 4787 3024 4791
rect 3018 4786 3024 4787
rect 3054 4784 3060 4785
rect 1935 4781 1939 4782
rect 1974 4783 1980 4784
rect 250 4771 256 4772
rect 250 4767 251 4771
rect 255 4767 256 4771
rect 250 4766 256 4767
rect 268 4720 270 4781
rect 274 4767 280 4768
rect 274 4763 275 4767
rect 279 4763 280 4767
rect 274 4762 280 4763
rect 110 4716 111 4720
rect 115 4716 116 4720
rect 110 4715 116 4716
rect 130 4719 136 4720
rect 130 4715 131 4719
rect 135 4715 136 4719
rect 130 4714 136 4715
rect 266 4719 272 4720
rect 266 4715 267 4719
rect 271 4715 272 4719
rect 266 4714 272 4715
rect 158 4704 164 4705
rect 276 4704 278 4762
rect 404 4720 406 4781
rect 410 4767 416 4768
rect 410 4763 411 4767
rect 415 4763 416 4767
rect 410 4762 416 4763
rect 402 4719 408 4720
rect 402 4715 403 4719
rect 407 4715 408 4719
rect 402 4714 408 4715
rect 294 4704 300 4705
rect 412 4704 414 4762
rect 540 4720 542 4781
rect 546 4767 552 4768
rect 546 4763 547 4767
rect 551 4763 552 4767
rect 546 4762 552 4763
rect 538 4719 544 4720
rect 538 4715 539 4719
rect 543 4715 544 4719
rect 538 4714 544 4715
rect 430 4704 436 4705
rect 548 4704 550 4762
rect 676 4720 678 4781
rect 682 4767 688 4768
rect 682 4763 683 4767
rect 687 4763 688 4767
rect 682 4762 688 4763
rect 674 4719 680 4720
rect 674 4715 675 4719
rect 679 4715 680 4719
rect 674 4714 680 4715
rect 566 4704 572 4705
rect 684 4704 686 4762
rect 1936 4721 1938 4781
rect 1974 4779 1975 4783
rect 1979 4779 1980 4783
rect 2454 4780 2455 4784
rect 2459 4780 2460 4784
rect 2454 4779 2460 4780
rect 2578 4783 2584 4784
rect 2578 4779 2579 4783
rect 2583 4779 2584 4783
rect 2598 4780 2599 4784
rect 2603 4780 2604 4784
rect 2598 4779 2604 4780
rect 2730 4783 2736 4784
rect 2730 4779 2731 4783
rect 2735 4779 2736 4783
rect 2750 4780 2751 4784
rect 2755 4780 2756 4784
rect 2750 4779 2756 4780
rect 2850 4783 2856 4784
rect 2850 4779 2851 4783
rect 2855 4779 2856 4783
rect 2902 4780 2903 4784
rect 2907 4780 2908 4784
rect 2902 4779 2908 4780
rect 3002 4783 3008 4784
rect 3002 4779 3003 4783
rect 3007 4779 3008 4783
rect 3054 4780 3055 4784
rect 3059 4780 3060 4784
rect 3054 4779 3060 4780
rect 3206 4784 3212 4785
rect 3304 4784 3306 4850
rect 3342 4843 3348 4844
rect 3342 4839 3343 4843
rect 3347 4839 3348 4843
rect 3342 4838 3348 4839
rect 3206 4780 3207 4784
rect 3211 4780 3212 4784
rect 3206 4779 3212 4780
rect 3302 4783 3308 4784
rect 3302 4779 3303 4783
rect 3307 4779 3308 4783
rect 1974 4778 1980 4779
rect 1976 4751 1978 4778
rect 2456 4751 2458 4779
rect 2578 4778 2584 4779
rect 2600 4751 2602 4779
rect 2730 4778 2736 4779
rect 2752 4751 2754 4779
rect 2850 4778 2856 4779
rect 2904 4751 2906 4779
rect 3002 4778 3008 4779
rect 3056 4751 3058 4779
rect 3208 4751 3210 4779
rect 3302 4778 3308 4779
rect 1975 4750 1979 4751
rect 1975 4745 1979 4746
rect 2023 4750 2027 4751
rect 2023 4745 2027 4746
rect 2159 4750 2163 4751
rect 2159 4745 2163 4746
rect 2295 4750 2299 4751
rect 2295 4745 2299 4746
rect 2431 4750 2435 4751
rect 2431 4745 2435 4746
rect 2455 4750 2459 4751
rect 2455 4745 2459 4746
rect 2567 4750 2571 4751
rect 2567 4745 2571 4746
rect 2599 4750 2603 4751
rect 2599 4745 2603 4746
rect 2703 4750 2707 4751
rect 2703 4745 2707 4746
rect 2751 4750 2755 4751
rect 2751 4745 2755 4746
rect 2839 4750 2843 4751
rect 2839 4745 2843 4746
rect 2903 4750 2907 4751
rect 2903 4745 2907 4746
rect 2975 4750 2979 4751
rect 2975 4745 2979 4746
rect 3055 4750 3059 4751
rect 3055 4745 3059 4746
rect 3111 4750 3115 4751
rect 3111 4745 3115 4746
rect 3207 4750 3211 4751
rect 3207 4745 3211 4746
rect 3247 4750 3251 4751
rect 3247 4745 3251 4746
rect 1976 4722 1978 4745
rect 1974 4721 1980 4722
rect 2024 4721 2026 4745
rect 2160 4721 2162 4745
rect 2296 4721 2298 4745
rect 2432 4721 2434 4745
rect 2568 4721 2570 4745
rect 2704 4721 2706 4745
rect 2840 4721 2842 4745
rect 2976 4721 2978 4745
rect 3112 4721 3114 4745
rect 3248 4721 3250 4745
rect 1934 4720 1940 4721
rect 1934 4716 1935 4720
rect 1939 4716 1940 4720
rect 1974 4717 1975 4721
rect 1979 4717 1980 4721
rect 1974 4716 1980 4717
rect 2022 4720 2028 4721
rect 2158 4720 2164 4721
rect 2294 4720 2300 4721
rect 2430 4720 2436 4721
rect 2566 4720 2572 4721
rect 2702 4720 2708 4721
rect 2838 4720 2844 4721
rect 2974 4720 2980 4721
rect 3110 4720 3116 4721
rect 3246 4720 3252 4721
rect 3344 4720 3346 4838
rect 3800 4801 3802 4861
rect 3840 4817 3842 4877
rect 3838 4816 3844 4817
rect 3860 4816 3862 4877
rect 4076 4816 4078 4877
rect 4084 4868 4086 4982
rect 4194 4973 4200 4974
rect 4194 4969 4195 4973
rect 4199 4969 4200 4973
rect 4194 4968 4200 4969
rect 4196 4883 4198 4968
rect 4216 4924 4218 5057
rect 4376 5019 4378 5059
rect 4223 5018 4227 5019
rect 4223 5013 4227 5014
rect 4375 5018 4379 5019
rect 4375 5013 4379 5014
rect 4447 5018 4451 5019
rect 4447 5013 4451 5014
rect 4224 4989 4226 5013
rect 4448 4989 4450 5013
rect 4222 4988 4228 4989
rect 4446 4988 4452 4989
rect 4604 4988 4606 5122
rect 4622 5064 4628 5065
rect 4716 5064 4718 5178
rect 4796 5147 4798 5228
rect 4900 5184 4902 5306
rect 4992 5279 4994 5307
rect 5662 5306 5668 5307
rect 5664 5279 5666 5306
rect 4991 5278 4995 5279
rect 4991 5273 4995 5274
rect 5039 5278 5043 5279
rect 5039 5273 5043 5274
rect 5663 5278 5667 5279
rect 5663 5273 5667 5274
rect 5040 5249 5042 5273
rect 5664 5250 5666 5273
rect 5662 5249 5668 5250
rect 5038 5248 5044 5249
rect 4922 5247 4928 5248
rect 4922 5243 4923 5247
rect 4927 5243 4928 5247
rect 5038 5244 5039 5248
rect 5043 5244 5044 5248
rect 5038 5243 5044 5244
rect 5134 5247 5140 5248
rect 5134 5243 5135 5247
rect 5139 5243 5140 5247
rect 5662 5245 5663 5249
rect 5667 5245 5668 5249
rect 5662 5244 5668 5245
rect 4922 5242 4928 5243
rect 5134 5242 5140 5243
rect 4924 5184 4926 5242
rect 5010 5233 5016 5234
rect 5010 5229 5011 5233
rect 5015 5229 5016 5233
rect 5010 5228 5016 5229
rect 4898 5183 4904 5184
rect 4898 5179 4899 5183
rect 4903 5179 4904 5183
rect 4898 5178 4904 5179
rect 4922 5183 4928 5184
rect 4922 5179 4923 5183
rect 4927 5179 4928 5183
rect 4922 5178 4928 5179
rect 5012 5147 5014 5228
rect 4795 5146 4799 5147
rect 4795 5141 4799 5142
rect 4843 5146 4847 5147
rect 4843 5141 4847 5142
rect 5011 5146 5015 5147
rect 5011 5141 5015 5142
rect 5099 5146 5103 5147
rect 5099 5141 5103 5142
rect 4844 5080 4846 5141
rect 5100 5080 5102 5141
rect 5136 5132 5138 5242
rect 5662 5232 5668 5233
rect 5662 5228 5663 5232
rect 5667 5228 5668 5232
rect 5662 5227 5668 5228
rect 5664 5147 5666 5227
rect 5663 5146 5667 5147
rect 5663 5141 5667 5142
rect 5134 5131 5140 5132
rect 5134 5127 5135 5131
rect 5139 5127 5140 5131
rect 5134 5126 5140 5127
rect 5664 5081 5666 5141
rect 5662 5080 5668 5081
rect 4842 5079 4848 5080
rect 4842 5075 4843 5079
rect 4847 5075 4848 5079
rect 4842 5074 4848 5075
rect 5098 5079 5104 5080
rect 5098 5075 5099 5079
rect 5103 5075 5104 5079
rect 5662 5076 5663 5080
rect 5667 5076 5668 5080
rect 5662 5075 5668 5076
rect 5098 5074 5104 5075
rect 4870 5064 4876 5065
rect 5126 5064 5132 5065
rect 4622 5060 4623 5064
rect 4627 5060 4628 5064
rect 4622 5059 4628 5060
rect 4714 5063 4720 5064
rect 4714 5059 4715 5063
rect 4719 5059 4720 5063
rect 4870 5060 4871 5064
rect 4875 5060 4876 5064
rect 4870 5059 4876 5060
rect 4966 5063 4972 5064
rect 4966 5059 4967 5063
rect 4971 5059 4972 5063
rect 5126 5060 5127 5064
rect 5131 5060 5132 5064
rect 5126 5059 5132 5060
rect 5662 5063 5668 5064
rect 5662 5059 5663 5063
rect 5667 5059 5668 5063
rect 4624 5019 4626 5059
rect 4714 5058 4720 5059
rect 4872 5019 4874 5059
rect 4966 5058 4972 5059
rect 4623 5018 4627 5019
rect 4623 5013 4627 5014
rect 4655 5018 4659 5019
rect 4655 5013 4659 5014
rect 4855 5018 4859 5019
rect 4855 5013 4859 5014
rect 4871 5018 4875 5019
rect 4871 5013 4875 5014
rect 4656 4989 4658 5013
rect 4856 4989 4858 5013
rect 4654 4988 4660 4989
rect 4854 4988 4860 4989
rect 4222 4984 4223 4988
rect 4227 4984 4228 4988
rect 4222 4983 4228 4984
rect 4318 4987 4324 4988
rect 4318 4983 4319 4987
rect 4323 4983 4324 4987
rect 4446 4984 4447 4988
rect 4451 4984 4452 4988
rect 4446 4983 4452 4984
rect 4602 4987 4608 4988
rect 4602 4983 4603 4987
rect 4607 4983 4608 4987
rect 4654 4984 4655 4988
rect 4659 4984 4660 4988
rect 4654 4983 4660 4984
rect 4750 4987 4756 4988
rect 4750 4983 4751 4987
rect 4755 4983 4756 4987
rect 4854 4984 4855 4988
rect 4859 4984 4860 4988
rect 4854 4983 4860 4984
rect 4950 4987 4956 4988
rect 4950 4983 4951 4987
rect 4955 4983 4956 4987
rect 4318 4982 4324 4983
rect 4602 4982 4608 4983
rect 4750 4982 4756 4983
rect 4950 4982 4956 4983
rect 4214 4923 4220 4924
rect 4214 4919 4215 4923
rect 4219 4919 4220 4923
rect 4214 4918 4220 4919
rect 4320 4916 4322 4982
rect 4418 4973 4424 4974
rect 4418 4969 4419 4973
rect 4423 4969 4424 4973
rect 4418 4968 4424 4969
rect 4626 4973 4632 4974
rect 4626 4969 4627 4973
rect 4631 4969 4632 4973
rect 4626 4968 4632 4969
rect 4318 4915 4324 4916
rect 4318 4911 4319 4915
rect 4323 4911 4324 4915
rect 4318 4910 4324 4911
rect 4420 4883 4422 4968
rect 4426 4923 4432 4924
rect 4426 4919 4427 4923
rect 4431 4919 4432 4923
rect 4426 4918 4432 4919
rect 4195 4882 4199 4883
rect 4195 4877 4199 4878
rect 4299 4882 4303 4883
rect 4299 4877 4303 4878
rect 4419 4882 4423 4883
rect 4419 4877 4423 4878
rect 4082 4867 4088 4868
rect 4082 4863 4083 4867
rect 4087 4863 4088 4867
rect 4082 4862 4088 4863
rect 4300 4816 4302 4877
rect 3838 4812 3839 4816
rect 3843 4812 3844 4816
rect 3838 4811 3844 4812
rect 3858 4815 3864 4816
rect 3858 4811 3859 4815
rect 3863 4811 3864 4815
rect 3858 4810 3864 4811
rect 4074 4815 4080 4816
rect 4074 4811 4075 4815
rect 4079 4811 4080 4815
rect 4074 4810 4080 4811
rect 4298 4815 4304 4816
rect 4298 4811 4299 4815
rect 4303 4811 4304 4815
rect 4298 4810 4304 4811
rect 3798 4800 3804 4801
rect 3886 4800 3892 4801
rect 4102 4800 4108 4801
rect 3798 4796 3799 4800
rect 3803 4796 3804 4800
rect 3798 4795 3804 4796
rect 3838 4799 3844 4800
rect 3838 4795 3839 4799
rect 3843 4795 3844 4799
rect 3886 4796 3887 4800
rect 3891 4796 3892 4800
rect 3886 4795 3892 4796
rect 3982 4799 3988 4800
rect 3982 4795 3983 4799
rect 3987 4795 3988 4799
rect 4102 4796 4103 4800
rect 4107 4796 4108 4800
rect 4102 4795 4108 4796
rect 4326 4800 4332 4801
rect 4428 4800 4430 4918
rect 4628 4883 4630 4968
rect 4507 4882 4511 4883
rect 4507 4877 4511 4878
rect 4627 4882 4631 4883
rect 4627 4877 4631 4878
rect 4699 4882 4703 4883
rect 4699 4877 4703 4878
rect 4508 4816 4510 4877
rect 4630 4871 4636 4872
rect 4630 4867 4631 4871
rect 4635 4867 4636 4871
rect 4630 4866 4636 4867
rect 4602 4863 4608 4864
rect 4602 4859 4603 4863
rect 4607 4859 4608 4863
rect 4602 4858 4608 4859
rect 4506 4815 4512 4816
rect 4506 4811 4507 4815
rect 4511 4811 4512 4815
rect 4506 4810 4512 4811
rect 4534 4800 4540 4801
rect 4326 4796 4327 4800
rect 4331 4796 4332 4800
rect 4326 4795 4332 4796
rect 4426 4799 4432 4800
rect 4426 4795 4427 4799
rect 4431 4795 4432 4799
rect 4534 4796 4535 4800
rect 4539 4796 4540 4800
rect 4534 4795 4540 4796
rect 3838 4794 3844 4795
rect 3798 4783 3804 4784
rect 3798 4779 3799 4783
rect 3803 4779 3804 4783
rect 3798 4778 3804 4779
rect 3800 4751 3802 4778
rect 3840 4771 3842 4794
rect 3888 4771 3890 4795
rect 3982 4794 3988 4795
rect 3839 4770 3843 4771
rect 3839 4765 3843 4766
rect 3887 4770 3891 4771
rect 3887 4765 3891 4766
rect 3399 4750 3403 4751
rect 3399 4745 3403 4746
rect 3543 4750 3547 4751
rect 3543 4745 3547 4746
rect 3679 4750 3683 4751
rect 3679 4745 3683 4746
rect 3799 4750 3803 4751
rect 3799 4745 3803 4746
rect 3400 4721 3402 4745
rect 3544 4721 3546 4745
rect 3680 4721 3682 4745
rect 3800 4722 3802 4745
rect 3840 4742 3842 4765
rect 3838 4741 3844 4742
rect 3838 4737 3839 4741
rect 3843 4737 3844 4741
rect 3838 4736 3844 4737
rect 3838 4724 3844 4725
rect 3798 4721 3804 4722
rect 3398 4720 3404 4721
rect 2022 4716 2023 4720
rect 2027 4716 2028 4720
rect 1934 4715 1940 4716
rect 2022 4715 2028 4716
rect 2122 4719 2128 4720
rect 2122 4715 2123 4719
rect 2127 4715 2128 4719
rect 2158 4716 2159 4720
rect 2163 4716 2164 4720
rect 2158 4715 2164 4716
rect 2258 4719 2264 4720
rect 2258 4715 2259 4719
rect 2263 4715 2264 4719
rect 2294 4716 2295 4720
rect 2299 4716 2300 4720
rect 2294 4715 2300 4716
rect 2394 4719 2400 4720
rect 2394 4715 2395 4719
rect 2399 4715 2400 4719
rect 2430 4716 2431 4720
rect 2435 4716 2436 4720
rect 2430 4715 2436 4716
rect 2530 4719 2536 4720
rect 2530 4715 2531 4719
rect 2535 4715 2536 4719
rect 2566 4716 2567 4720
rect 2571 4716 2572 4720
rect 2566 4715 2572 4716
rect 2666 4719 2672 4720
rect 2666 4715 2667 4719
rect 2671 4715 2672 4719
rect 2702 4716 2703 4720
rect 2707 4716 2708 4720
rect 2702 4715 2708 4716
rect 2802 4719 2808 4720
rect 2802 4715 2803 4719
rect 2807 4715 2808 4719
rect 2838 4716 2839 4720
rect 2843 4716 2844 4720
rect 2838 4715 2844 4716
rect 2938 4719 2944 4720
rect 2938 4715 2939 4719
rect 2943 4715 2944 4719
rect 2974 4716 2975 4720
rect 2979 4716 2980 4720
rect 2974 4715 2980 4716
rect 3074 4719 3080 4720
rect 3074 4715 3075 4719
rect 3079 4715 3080 4719
rect 3110 4716 3111 4720
rect 3115 4716 3116 4720
rect 3110 4715 3116 4716
rect 3210 4719 3216 4720
rect 3210 4715 3211 4719
rect 3215 4715 3216 4719
rect 3246 4716 3247 4720
rect 3251 4716 3252 4720
rect 3246 4715 3252 4716
rect 3342 4719 3348 4720
rect 3342 4715 3343 4719
rect 3347 4715 3348 4719
rect 3398 4716 3399 4720
rect 3403 4716 3404 4720
rect 3398 4715 3404 4716
rect 3542 4720 3548 4721
rect 3678 4720 3684 4721
rect 3542 4716 3543 4720
rect 3547 4716 3548 4720
rect 3542 4715 3548 4716
rect 3638 4719 3644 4720
rect 3638 4715 3639 4719
rect 3643 4715 3644 4719
rect 3678 4716 3679 4720
rect 3683 4716 3684 4720
rect 3678 4715 3684 4716
rect 3770 4719 3776 4720
rect 3770 4715 3771 4719
rect 3775 4715 3776 4719
rect 3798 4717 3799 4721
rect 3803 4717 3804 4721
rect 3838 4720 3839 4724
rect 3843 4720 3844 4724
rect 3838 4719 3844 4720
rect 3798 4716 3804 4717
rect 2122 4714 2128 4715
rect 2258 4714 2264 4715
rect 2394 4714 2400 4715
rect 2530 4714 2536 4715
rect 2666 4714 2672 4715
rect 2802 4714 2808 4715
rect 2938 4714 2944 4715
rect 3074 4714 3080 4715
rect 3210 4714 3216 4715
rect 3342 4714 3348 4715
rect 3638 4714 3644 4715
rect 3770 4714 3776 4715
rect 1994 4705 2000 4706
rect 702 4704 708 4705
rect 1974 4704 1980 4705
rect 110 4703 116 4704
rect 110 4699 111 4703
rect 115 4699 116 4703
rect 158 4700 159 4704
rect 163 4700 164 4704
rect 158 4699 164 4700
rect 274 4703 280 4704
rect 274 4699 275 4703
rect 279 4699 280 4703
rect 294 4700 295 4704
rect 299 4700 300 4704
rect 294 4699 300 4700
rect 410 4703 416 4704
rect 410 4699 411 4703
rect 415 4699 416 4703
rect 430 4700 431 4704
rect 435 4700 436 4704
rect 430 4699 436 4700
rect 546 4703 552 4704
rect 546 4699 547 4703
rect 551 4699 552 4703
rect 566 4700 567 4704
rect 571 4700 572 4704
rect 566 4699 572 4700
rect 682 4703 688 4704
rect 682 4699 683 4703
rect 687 4699 688 4703
rect 702 4700 703 4704
rect 707 4700 708 4704
rect 702 4699 708 4700
rect 802 4703 808 4704
rect 802 4699 803 4703
rect 807 4699 808 4703
rect 110 4698 116 4699
rect 112 4667 114 4698
rect 160 4667 162 4699
rect 274 4698 280 4699
rect 296 4667 298 4699
rect 410 4698 416 4699
rect 432 4667 434 4699
rect 546 4698 552 4699
rect 568 4667 570 4699
rect 682 4698 688 4699
rect 704 4667 706 4699
rect 802 4698 808 4699
rect 1934 4703 1940 4704
rect 1934 4699 1935 4703
rect 1939 4699 1940 4703
rect 1974 4700 1975 4704
rect 1979 4700 1980 4704
rect 1994 4701 1995 4705
rect 1999 4701 2000 4705
rect 1994 4700 2000 4701
rect 1974 4699 1980 4700
rect 1934 4698 1940 4699
rect 111 4666 115 4667
rect 111 4661 115 4662
rect 159 4666 163 4667
rect 159 4661 163 4662
rect 295 4666 299 4667
rect 295 4661 299 4662
rect 431 4666 435 4667
rect 431 4661 435 4662
rect 567 4666 571 4667
rect 567 4661 571 4662
rect 703 4666 707 4667
rect 703 4661 707 4662
rect 112 4638 114 4661
rect 110 4637 116 4638
rect 160 4637 162 4661
rect 296 4637 298 4661
rect 432 4637 434 4661
rect 568 4637 570 4661
rect 704 4637 706 4661
rect 110 4633 111 4637
rect 115 4633 116 4637
rect 110 4632 116 4633
rect 158 4636 164 4637
rect 158 4632 159 4636
rect 163 4632 164 4636
rect 158 4631 164 4632
rect 294 4636 300 4637
rect 430 4636 436 4637
rect 566 4636 572 4637
rect 702 4636 708 4637
rect 294 4632 295 4636
rect 299 4632 300 4636
rect 294 4631 300 4632
rect 394 4635 400 4636
rect 394 4631 395 4635
rect 399 4631 400 4635
rect 430 4632 431 4636
rect 435 4632 436 4636
rect 430 4631 436 4632
rect 530 4635 536 4636
rect 530 4631 531 4635
rect 535 4631 536 4635
rect 566 4632 567 4636
rect 571 4632 572 4636
rect 566 4631 572 4632
rect 666 4635 672 4636
rect 666 4631 667 4635
rect 671 4631 672 4635
rect 702 4632 703 4636
rect 707 4632 708 4636
rect 702 4631 708 4632
rect 794 4635 800 4636
rect 794 4631 795 4635
rect 799 4631 800 4635
rect 394 4630 400 4631
rect 530 4630 536 4631
rect 666 4630 672 4631
rect 794 4630 800 4631
rect 130 4621 136 4622
rect 110 4620 116 4621
rect 110 4616 111 4620
rect 115 4616 116 4620
rect 130 4617 131 4621
rect 135 4617 136 4621
rect 130 4616 136 4617
rect 266 4621 272 4622
rect 266 4617 267 4621
rect 271 4617 272 4621
rect 266 4616 272 4617
rect 110 4615 116 4616
rect 112 4547 114 4615
rect 132 4547 134 4616
rect 268 4547 270 4616
rect 396 4572 398 4630
rect 402 4621 408 4622
rect 402 4617 403 4621
rect 407 4617 408 4621
rect 402 4616 408 4617
rect 394 4571 400 4572
rect 394 4567 395 4571
rect 399 4567 400 4571
rect 394 4566 400 4567
rect 404 4547 406 4616
rect 532 4572 534 4630
rect 538 4621 544 4622
rect 538 4617 539 4621
rect 543 4617 544 4621
rect 538 4616 544 4617
rect 530 4571 536 4572
rect 530 4567 531 4571
rect 535 4567 536 4571
rect 530 4566 536 4567
rect 540 4547 542 4616
rect 668 4572 670 4630
rect 674 4621 680 4622
rect 674 4617 675 4621
rect 679 4617 680 4621
rect 674 4616 680 4617
rect 666 4571 672 4572
rect 666 4567 667 4571
rect 671 4567 672 4571
rect 666 4566 672 4567
rect 676 4547 678 4616
rect 111 4546 115 4547
rect 111 4541 115 4542
rect 131 4546 135 4547
rect 131 4541 135 4542
rect 267 4546 271 4547
rect 267 4541 271 4542
rect 339 4546 343 4547
rect 339 4541 343 4542
rect 403 4546 407 4547
rect 403 4541 407 4542
rect 515 4546 519 4547
rect 515 4541 519 4542
rect 539 4546 543 4547
rect 539 4541 543 4542
rect 675 4546 679 4547
rect 675 4541 679 4542
rect 691 4546 695 4547
rect 691 4541 695 4542
rect 112 4481 114 4541
rect 110 4480 116 4481
rect 340 4480 342 4541
rect 516 4480 518 4541
rect 522 4527 528 4528
rect 522 4523 523 4527
rect 527 4523 528 4527
rect 522 4522 528 4523
rect 110 4476 111 4480
rect 115 4476 116 4480
rect 110 4475 116 4476
rect 338 4479 344 4480
rect 338 4475 339 4479
rect 343 4475 344 4479
rect 338 4474 344 4475
rect 514 4479 520 4480
rect 514 4475 515 4479
rect 519 4475 520 4479
rect 514 4474 520 4475
rect 366 4464 372 4465
rect 524 4464 526 4522
rect 692 4480 694 4541
rect 796 4536 798 4630
rect 804 4564 806 4698
rect 1936 4667 1938 4698
rect 1935 4666 1939 4667
rect 1935 4661 1939 4662
rect 1936 4638 1938 4661
rect 1934 4637 1940 4638
rect 1934 4633 1935 4637
rect 1939 4633 1940 4637
rect 1934 4632 1940 4633
rect 1934 4620 1940 4621
rect 1934 4616 1935 4620
rect 1939 4616 1940 4620
rect 1934 4615 1940 4616
rect 802 4563 808 4564
rect 802 4559 803 4563
rect 807 4559 808 4563
rect 802 4558 808 4559
rect 1936 4547 1938 4615
rect 1976 4607 1978 4699
rect 1996 4607 1998 4700
rect 2124 4656 2126 4714
rect 2130 4705 2136 4706
rect 2130 4701 2131 4705
rect 2135 4701 2136 4705
rect 2130 4700 2136 4701
rect 2122 4655 2128 4656
rect 2122 4651 2123 4655
rect 2127 4651 2128 4655
rect 2122 4650 2128 4651
rect 2132 4607 2134 4700
rect 2260 4656 2262 4714
rect 2266 4705 2272 4706
rect 2266 4701 2267 4705
rect 2271 4701 2272 4705
rect 2266 4700 2272 4701
rect 2258 4655 2264 4656
rect 2258 4651 2259 4655
rect 2263 4651 2264 4655
rect 2258 4650 2264 4651
rect 2268 4607 2270 4700
rect 2396 4656 2398 4714
rect 2402 4705 2408 4706
rect 2402 4701 2403 4705
rect 2407 4701 2408 4705
rect 2402 4700 2408 4701
rect 2394 4655 2400 4656
rect 2394 4651 2395 4655
rect 2399 4651 2400 4655
rect 2394 4650 2400 4651
rect 2404 4607 2406 4700
rect 2532 4656 2534 4714
rect 2538 4705 2544 4706
rect 2538 4701 2539 4705
rect 2543 4701 2544 4705
rect 2538 4700 2544 4701
rect 2530 4655 2536 4656
rect 2530 4651 2531 4655
rect 2535 4651 2536 4655
rect 2530 4650 2536 4651
rect 2442 4647 2448 4648
rect 2442 4643 2443 4647
rect 2447 4643 2448 4647
rect 2442 4642 2448 4643
rect 1975 4606 1979 4607
rect 1975 4601 1979 4602
rect 1995 4606 1999 4607
rect 1995 4601 1999 4602
rect 2131 4606 2135 4607
rect 2131 4601 2135 4602
rect 2267 4606 2271 4607
rect 2267 4601 2271 4602
rect 2323 4606 2327 4607
rect 2323 4601 2327 4602
rect 2403 4606 2407 4607
rect 2403 4601 2407 4602
rect 875 4546 879 4547
rect 875 4541 879 4542
rect 1059 4546 1063 4547
rect 1059 4541 1063 4542
rect 1243 4546 1247 4547
rect 1243 4541 1247 4542
rect 1427 4546 1431 4547
rect 1427 4541 1431 4542
rect 1619 4546 1623 4547
rect 1619 4541 1623 4542
rect 1787 4546 1791 4547
rect 1787 4541 1791 4542
rect 1935 4546 1939 4547
rect 1935 4541 1939 4542
rect 1976 4541 1978 4601
rect 794 4535 800 4536
rect 794 4531 795 4535
rect 799 4531 800 4535
rect 794 4530 800 4531
rect 698 4527 704 4528
rect 698 4523 699 4527
rect 703 4523 704 4527
rect 698 4522 704 4523
rect 690 4479 696 4480
rect 690 4475 691 4479
rect 695 4475 696 4479
rect 690 4474 696 4475
rect 542 4464 548 4465
rect 700 4464 702 4522
rect 876 4480 878 4541
rect 882 4527 888 4528
rect 882 4523 883 4527
rect 887 4523 888 4527
rect 882 4522 888 4523
rect 874 4479 880 4480
rect 874 4475 875 4479
rect 879 4475 880 4479
rect 874 4474 880 4475
rect 718 4464 724 4465
rect 884 4464 886 4522
rect 1060 4480 1062 4541
rect 1066 4527 1072 4528
rect 1066 4523 1067 4527
rect 1071 4523 1072 4527
rect 1066 4522 1072 4523
rect 1058 4479 1064 4480
rect 1058 4475 1059 4479
rect 1063 4475 1064 4479
rect 1058 4474 1064 4475
rect 902 4464 908 4465
rect 1068 4464 1070 4522
rect 1244 4480 1246 4541
rect 1418 4531 1424 4532
rect 1418 4527 1419 4531
rect 1423 4527 1424 4531
rect 1418 4526 1424 4527
rect 1242 4479 1248 4480
rect 1242 4475 1243 4479
rect 1247 4475 1248 4479
rect 1242 4474 1248 4475
rect 1086 4464 1092 4465
rect 1270 4464 1276 4465
rect 110 4463 116 4464
rect 110 4459 111 4463
rect 115 4459 116 4463
rect 366 4460 367 4464
rect 371 4460 372 4464
rect 366 4459 372 4460
rect 522 4463 528 4464
rect 522 4459 523 4463
rect 527 4459 528 4463
rect 542 4460 543 4464
rect 547 4460 548 4464
rect 542 4459 548 4460
rect 698 4463 704 4464
rect 698 4459 699 4463
rect 703 4459 704 4463
rect 718 4460 719 4464
rect 723 4460 724 4464
rect 718 4459 724 4460
rect 882 4463 888 4464
rect 882 4459 883 4463
rect 887 4459 888 4463
rect 902 4460 903 4464
rect 907 4460 908 4464
rect 902 4459 908 4460
rect 1066 4463 1072 4464
rect 1066 4459 1067 4463
rect 1071 4459 1072 4463
rect 1086 4460 1087 4464
rect 1091 4460 1092 4464
rect 1086 4459 1092 4460
rect 1178 4463 1184 4464
rect 1178 4459 1179 4463
rect 1183 4459 1184 4463
rect 1270 4460 1271 4464
rect 1275 4460 1276 4464
rect 1270 4459 1276 4460
rect 110 4458 116 4459
rect 112 4435 114 4458
rect 368 4435 370 4459
rect 522 4458 528 4459
rect 544 4435 546 4459
rect 698 4458 704 4459
rect 720 4435 722 4459
rect 882 4458 888 4459
rect 904 4435 906 4459
rect 1066 4458 1072 4459
rect 1088 4435 1090 4459
rect 1178 4458 1184 4459
rect 1180 4443 1182 4458
rect 1176 4441 1182 4443
rect 111 4434 115 4435
rect 111 4429 115 4430
rect 367 4434 371 4435
rect 367 4429 371 4430
rect 543 4434 547 4435
rect 543 4429 547 4430
rect 567 4434 571 4435
rect 567 4429 571 4430
rect 711 4434 715 4435
rect 711 4429 715 4430
rect 719 4434 723 4435
rect 719 4429 723 4430
rect 863 4434 867 4435
rect 863 4429 867 4430
rect 903 4434 907 4435
rect 903 4429 907 4430
rect 1023 4434 1027 4435
rect 1023 4429 1027 4430
rect 1087 4434 1091 4435
rect 1087 4429 1091 4430
rect 112 4406 114 4429
rect 110 4405 116 4406
rect 568 4405 570 4429
rect 712 4405 714 4429
rect 864 4405 866 4429
rect 1024 4405 1026 4429
rect 110 4401 111 4405
rect 115 4401 116 4405
rect 110 4400 116 4401
rect 566 4404 572 4405
rect 710 4404 716 4405
rect 566 4400 567 4404
rect 571 4400 572 4404
rect 566 4399 572 4400
rect 666 4403 672 4404
rect 666 4399 667 4403
rect 671 4399 672 4403
rect 710 4400 711 4404
rect 715 4400 716 4404
rect 710 4399 716 4400
rect 862 4404 868 4405
rect 1022 4404 1028 4405
rect 862 4400 863 4404
rect 867 4400 868 4404
rect 862 4399 868 4400
rect 962 4403 968 4404
rect 962 4399 963 4403
rect 967 4399 968 4403
rect 1022 4400 1023 4404
rect 1027 4400 1028 4404
rect 1022 4399 1028 4400
rect 1122 4403 1128 4404
rect 1122 4399 1123 4403
rect 1127 4399 1128 4403
rect 666 4398 672 4399
rect 962 4398 968 4399
rect 1122 4398 1128 4399
rect 538 4389 544 4390
rect 110 4388 116 4389
rect 110 4384 111 4388
rect 115 4384 116 4388
rect 538 4385 539 4389
rect 543 4385 544 4389
rect 538 4384 544 4385
rect 110 4383 116 4384
rect 112 4303 114 4383
rect 540 4303 542 4384
rect 668 4340 670 4398
rect 682 4389 688 4390
rect 682 4385 683 4389
rect 687 4385 688 4389
rect 682 4384 688 4385
rect 834 4389 840 4390
rect 834 4385 835 4389
rect 839 4385 840 4389
rect 834 4384 840 4385
rect 666 4339 672 4340
rect 666 4335 667 4339
rect 671 4335 672 4339
rect 666 4334 672 4335
rect 684 4303 686 4384
rect 836 4303 838 4384
rect 964 4340 966 4398
rect 994 4389 1000 4390
rect 994 4385 995 4389
rect 999 4385 1000 4389
rect 994 4384 1000 4385
rect 962 4339 968 4340
rect 962 4335 963 4339
rect 967 4335 968 4339
rect 962 4334 968 4335
rect 996 4303 998 4384
rect 1124 4340 1126 4398
rect 1154 4389 1160 4390
rect 1154 4385 1155 4389
rect 1159 4385 1160 4389
rect 1154 4384 1160 4385
rect 1122 4339 1128 4340
rect 1122 4335 1123 4339
rect 1127 4335 1128 4339
rect 1122 4334 1128 4335
rect 1156 4303 1158 4384
rect 1176 4332 1178 4441
rect 1272 4435 1274 4459
rect 1183 4434 1187 4435
rect 1183 4429 1187 4430
rect 1271 4434 1275 4435
rect 1271 4429 1275 4430
rect 1343 4434 1347 4435
rect 1343 4429 1347 4430
rect 1184 4405 1186 4429
rect 1344 4405 1346 4429
rect 1420 4411 1422 4526
rect 1428 4480 1430 4541
rect 1434 4527 1440 4528
rect 1434 4523 1435 4527
rect 1439 4523 1440 4527
rect 1434 4522 1440 4523
rect 1426 4479 1432 4480
rect 1426 4475 1427 4479
rect 1431 4475 1432 4479
rect 1426 4474 1432 4475
rect 1436 4464 1438 4522
rect 1620 4480 1622 4541
rect 1626 4527 1632 4528
rect 1626 4523 1627 4527
rect 1631 4523 1632 4527
rect 1626 4522 1632 4523
rect 1618 4479 1624 4480
rect 1618 4475 1619 4479
rect 1623 4475 1624 4479
rect 1618 4474 1624 4475
rect 1454 4464 1460 4465
rect 1628 4464 1630 4522
rect 1788 4480 1790 4541
rect 1794 4527 1800 4528
rect 1794 4523 1795 4527
rect 1799 4523 1800 4527
rect 1794 4522 1800 4523
rect 1786 4479 1792 4480
rect 1786 4475 1787 4479
rect 1791 4475 1792 4479
rect 1786 4474 1792 4475
rect 1646 4464 1652 4465
rect 1796 4464 1798 4522
rect 1936 4481 1938 4541
rect 1974 4540 1980 4541
rect 2324 4540 2326 4601
rect 1974 4536 1975 4540
rect 1979 4536 1980 4540
rect 1974 4535 1980 4536
rect 2322 4539 2328 4540
rect 2322 4535 2323 4539
rect 2327 4535 2328 4539
rect 2322 4534 2328 4535
rect 2350 4524 2356 4525
rect 2444 4524 2446 4642
rect 2540 4607 2542 4700
rect 2668 4656 2670 4714
rect 2674 4705 2680 4706
rect 2674 4701 2675 4705
rect 2679 4701 2680 4705
rect 2674 4700 2680 4701
rect 2666 4655 2672 4656
rect 2666 4651 2667 4655
rect 2671 4651 2672 4655
rect 2666 4650 2672 4651
rect 2676 4607 2678 4700
rect 2804 4656 2806 4714
rect 2810 4705 2816 4706
rect 2810 4701 2811 4705
rect 2815 4701 2816 4705
rect 2810 4700 2816 4701
rect 2802 4655 2808 4656
rect 2802 4651 2803 4655
rect 2807 4651 2808 4655
rect 2802 4650 2808 4651
rect 2812 4607 2814 4700
rect 2940 4656 2942 4714
rect 2946 4705 2952 4706
rect 2946 4701 2947 4705
rect 2951 4701 2952 4705
rect 2946 4700 2952 4701
rect 2938 4655 2944 4656
rect 2938 4651 2939 4655
rect 2943 4651 2944 4655
rect 2938 4650 2944 4651
rect 2948 4607 2950 4700
rect 3076 4656 3078 4714
rect 3082 4705 3088 4706
rect 3082 4701 3083 4705
rect 3087 4701 3088 4705
rect 3082 4700 3088 4701
rect 3074 4655 3080 4656
rect 3074 4651 3075 4655
rect 3079 4651 3080 4655
rect 3074 4650 3080 4651
rect 3084 4607 3086 4700
rect 3212 4656 3214 4714
rect 3218 4705 3224 4706
rect 3218 4701 3219 4705
rect 3223 4701 3224 4705
rect 3218 4700 3224 4701
rect 3370 4705 3376 4706
rect 3370 4701 3371 4705
rect 3375 4701 3376 4705
rect 3370 4700 3376 4701
rect 3514 4705 3520 4706
rect 3514 4701 3515 4705
rect 3519 4701 3520 4705
rect 3514 4700 3520 4701
rect 3210 4655 3216 4656
rect 3210 4651 3211 4655
rect 3215 4651 3216 4655
rect 3210 4650 3216 4651
rect 3220 4607 3222 4700
rect 3372 4607 3374 4700
rect 3516 4607 3518 4700
rect 2539 4606 2543 4607
rect 2539 4601 2543 4602
rect 2579 4606 2583 4607
rect 2579 4601 2583 4602
rect 2675 4606 2679 4607
rect 2675 4601 2679 4602
rect 2811 4606 2815 4607
rect 2811 4601 2815 4602
rect 2827 4606 2831 4607
rect 2827 4601 2831 4602
rect 2947 4606 2951 4607
rect 2947 4601 2951 4602
rect 3075 4606 3079 4607
rect 3075 4601 3079 4602
rect 3083 4606 3087 4607
rect 3083 4601 3087 4602
rect 3219 4606 3223 4607
rect 3219 4601 3223 4602
rect 3315 4606 3319 4607
rect 3315 4601 3319 4602
rect 3371 4606 3375 4607
rect 3371 4601 3375 4602
rect 3515 4606 3519 4607
rect 3515 4601 3519 4602
rect 3563 4606 3567 4607
rect 3563 4601 3567 4602
rect 2566 4591 2572 4592
rect 2566 4587 2567 4591
rect 2571 4587 2572 4591
rect 2566 4586 2572 4587
rect 2568 4532 2570 4586
rect 2580 4540 2582 4601
rect 2638 4591 2644 4592
rect 2638 4587 2639 4591
rect 2643 4587 2644 4591
rect 2638 4586 2644 4587
rect 2578 4539 2584 4540
rect 2578 4535 2579 4539
rect 2583 4535 2584 4539
rect 2578 4534 2584 4535
rect 2566 4531 2572 4532
rect 2566 4527 2567 4531
rect 2571 4527 2572 4531
rect 2566 4526 2572 4527
rect 2606 4524 2612 4525
rect 1974 4523 1980 4524
rect 1974 4519 1975 4523
rect 1979 4519 1980 4523
rect 2350 4520 2351 4524
rect 2355 4520 2356 4524
rect 2350 4519 2356 4520
rect 2442 4523 2448 4524
rect 2442 4519 2443 4523
rect 2447 4519 2448 4523
rect 2606 4520 2607 4524
rect 2611 4520 2612 4524
rect 2606 4519 2612 4520
rect 1974 4518 1980 4519
rect 1976 4487 1978 4518
rect 2352 4487 2354 4519
rect 2442 4518 2448 4519
rect 2608 4487 2610 4519
rect 1975 4486 1979 4487
rect 1975 4481 1979 4482
rect 2351 4486 2355 4487
rect 2351 4481 2355 4482
rect 2543 4486 2547 4487
rect 2543 4481 2547 4482
rect 2607 4486 2611 4487
rect 2607 4481 2611 4482
rect 1934 4480 1940 4481
rect 1934 4476 1935 4480
rect 1939 4476 1940 4480
rect 1934 4475 1940 4476
rect 1814 4464 1820 4465
rect 1434 4463 1440 4464
rect 1434 4459 1435 4463
rect 1439 4459 1440 4463
rect 1454 4460 1455 4464
rect 1459 4460 1460 4464
rect 1454 4459 1460 4460
rect 1626 4463 1632 4464
rect 1626 4459 1627 4463
rect 1631 4459 1632 4463
rect 1646 4460 1647 4464
rect 1651 4460 1652 4464
rect 1646 4459 1652 4460
rect 1794 4463 1800 4464
rect 1794 4459 1795 4463
rect 1799 4459 1800 4463
rect 1814 4460 1815 4464
rect 1819 4460 1820 4464
rect 1814 4459 1820 4460
rect 1910 4463 1916 4464
rect 1910 4459 1911 4463
rect 1915 4459 1916 4463
rect 1434 4458 1440 4459
rect 1456 4435 1458 4459
rect 1626 4458 1632 4459
rect 1648 4435 1650 4459
rect 1794 4458 1800 4459
rect 1816 4435 1818 4459
rect 1910 4458 1916 4459
rect 1934 4463 1940 4464
rect 1934 4459 1935 4463
rect 1939 4459 1940 4463
rect 1934 4458 1940 4459
rect 1976 4458 1978 4481
rect 1455 4434 1459 4435
rect 1455 4429 1459 4430
rect 1503 4434 1507 4435
rect 1503 4429 1507 4430
rect 1647 4434 1651 4435
rect 1647 4429 1651 4430
rect 1671 4434 1675 4435
rect 1671 4429 1675 4430
rect 1815 4434 1819 4435
rect 1815 4429 1819 4430
rect 1420 4409 1438 4411
rect 1182 4404 1188 4405
rect 1342 4404 1348 4405
rect 1436 4404 1438 4409
rect 1504 4405 1506 4429
rect 1672 4405 1674 4429
rect 1816 4405 1818 4429
rect 1502 4404 1508 4405
rect 1670 4404 1676 4405
rect 1814 4404 1820 4405
rect 1182 4400 1183 4404
rect 1187 4400 1188 4404
rect 1182 4399 1188 4400
rect 1278 4403 1284 4404
rect 1278 4399 1279 4403
rect 1283 4399 1284 4403
rect 1342 4400 1343 4404
rect 1347 4400 1348 4404
rect 1342 4399 1348 4400
rect 1434 4403 1440 4404
rect 1434 4399 1435 4403
rect 1439 4399 1440 4403
rect 1502 4400 1503 4404
rect 1507 4400 1508 4404
rect 1502 4399 1508 4400
rect 1594 4403 1600 4404
rect 1594 4399 1595 4403
rect 1599 4399 1600 4403
rect 1670 4400 1671 4404
rect 1675 4400 1676 4404
rect 1670 4399 1676 4400
rect 1770 4403 1776 4404
rect 1770 4399 1771 4403
rect 1775 4399 1776 4403
rect 1814 4400 1815 4404
rect 1819 4400 1820 4404
rect 1814 4399 1820 4400
rect 1278 4398 1284 4399
rect 1434 4398 1440 4399
rect 1594 4398 1600 4399
rect 1770 4398 1776 4399
rect 1174 4331 1180 4332
rect 1174 4327 1175 4331
rect 1179 4327 1180 4331
rect 1174 4326 1180 4327
rect 111 4302 115 4303
rect 111 4297 115 4298
rect 539 4302 543 4303
rect 539 4297 543 4298
rect 627 4302 631 4303
rect 627 4297 631 4298
rect 683 4302 687 4303
rect 683 4297 687 4298
rect 771 4302 775 4303
rect 771 4297 775 4298
rect 835 4302 839 4303
rect 835 4297 839 4298
rect 923 4302 927 4303
rect 923 4297 927 4298
rect 995 4302 999 4303
rect 1083 4302 1087 4303
rect 995 4297 999 4298
rect 1046 4299 1052 4300
rect 112 4237 114 4297
rect 110 4236 116 4237
rect 628 4236 630 4297
rect 772 4236 774 4297
rect 778 4283 784 4284
rect 778 4279 779 4283
rect 783 4279 784 4283
rect 778 4278 784 4279
rect 110 4232 111 4236
rect 115 4232 116 4236
rect 110 4231 116 4232
rect 626 4235 632 4236
rect 626 4231 627 4235
rect 631 4231 632 4235
rect 626 4230 632 4231
rect 770 4235 776 4236
rect 770 4231 771 4235
rect 775 4231 776 4235
rect 770 4230 776 4231
rect 654 4220 660 4221
rect 780 4220 782 4278
rect 924 4236 926 4297
rect 1046 4295 1047 4299
rect 1051 4295 1052 4299
rect 1083 4297 1087 4298
rect 1155 4302 1159 4303
rect 1155 4297 1159 4298
rect 1251 4302 1255 4303
rect 1251 4297 1255 4298
rect 1046 4294 1052 4295
rect 922 4235 928 4236
rect 922 4231 923 4235
rect 927 4231 928 4235
rect 922 4230 928 4231
rect 798 4220 804 4221
rect 950 4220 956 4221
rect 1048 4220 1050 4294
rect 1084 4236 1086 4297
rect 1206 4291 1212 4292
rect 1206 4287 1207 4291
rect 1211 4287 1212 4291
rect 1206 4286 1212 4287
rect 1082 4235 1088 4236
rect 1082 4231 1083 4235
rect 1087 4231 1088 4235
rect 1082 4230 1088 4231
rect 1110 4220 1116 4221
rect 1208 4220 1210 4286
rect 1252 4236 1254 4297
rect 1280 4288 1282 4398
rect 1314 4389 1320 4390
rect 1314 4385 1315 4389
rect 1319 4385 1320 4389
rect 1314 4384 1320 4385
rect 1474 4389 1480 4390
rect 1474 4385 1475 4389
rect 1479 4385 1480 4389
rect 1474 4384 1480 4385
rect 1316 4303 1318 4384
rect 1476 4303 1478 4384
rect 1542 4339 1548 4340
rect 1542 4335 1543 4339
rect 1547 4335 1548 4339
rect 1542 4334 1548 4335
rect 1315 4302 1319 4303
rect 1315 4297 1319 4298
rect 1419 4302 1423 4303
rect 1419 4297 1423 4298
rect 1475 4302 1479 4303
rect 1475 4297 1479 4298
rect 1278 4287 1284 4288
rect 1278 4283 1279 4287
rect 1283 4283 1284 4287
rect 1278 4282 1284 4283
rect 1420 4236 1422 4297
rect 1250 4235 1256 4236
rect 1250 4231 1251 4235
rect 1255 4231 1256 4235
rect 1250 4230 1256 4231
rect 1418 4235 1424 4236
rect 1418 4231 1419 4235
rect 1423 4231 1424 4235
rect 1418 4230 1424 4231
rect 1278 4220 1284 4221
rect 110 4219 116 4220
rect 110 4215 111 4219
rect 115 4215 116 4219
rect 654 4216 655 4220
rect 659 4216 660 4220
rect 654 4215 660 4216
rect 778 4219 784 4220
rect 778 4215 779 4219
rect 783 4215 784 4219
rect 798 4216 799 4220
rect 803 4216 804 4220
rect 798 4215 804 4216
rect 894 4219 900 4220
rect 894 4215 895 4219
rect 899 4215 900 4219
rect 950 4216 951 4220
rect 955 4216 956 4220
rect 950 4215 956 4216
rect 1046 4219 1052 4220
rect 1046 4215 1047 4219
rect 1051 4215 1052 4219
rect 1110 4216 1111 4220
rect 1115 4216 1116 4220
rect 1110 4215 1116 4216
rect 1206 4219 1212 4220
rect 1206 4215 1207 4219
rect 1211 4215 1212 4219
rect 1278 4216 1279 4220
rect 1283 4216 1284 4220
rect 1278 4215 1284 4216
rect 1446 4220 1452 4221
rect 1544 4220 1546 4334
rect 1596 4332 1598 4398
rect 1642 4389 1648 4390
rect 1642 4385 1643 4389
rect 1647 4385 1648 4389
rect 1642 4384 1648 4385
rect 1594 4331 1600 4332
rect 1594 4327 1595 4331
rect 1599 4327 1600 4331
rect 1594 4326 1600 4327
rect 1644 4303 1646 4384
rect 1772 4340 1774 4398
rect 1786 4389 1792 4390
rect 1786 4385 1787 4389
rect 1791 4385 1792 4389
rect 1786 4384 1792 4385
rect 1770 4339 1776 4340
rect 1770 4335 1771 4339
rect 1775 4335 1776 4339
rect 1770 4334 1776 4335
rect 1788 4303 1790 4384
rect 1912 4332 1914 4458
rect 1936 4435 1938 4458
rect 1974 4457 1980 4458
rect 2544 4457 2546 4481
rect 1974 4453 1975 4457
rect 1979 4453 1980 4457
rect 1974 4452 1980 4453
rect 2542 4456 2548 4457
rect 2640 4456 2642 4586
rect 2828 4540 2830 4601
rect 3066 4591 3072 4592
rect 3066 4587 3067 4591
rect 3071 4587 3072 4591
rect 3066 4586 3072 4587
rect 2826 4539 2832 4540
rect 2826 4535 2827 4539
rect 2831 4535 2832 4539
rect 2826 4534 2832 4535
rect 3068 4532 3070 4586
rect 3076 4540 3078 4601
rect 3316 4540 3318 4601
rect 3466 4591 3472 4592
rect 3466 4587 3467 4591
rect 3471 4587 3472 4591
rect 3466 4586 3472 4587
rect 3074 4539 3080 4540
rect 3074 4535 3075 4539
rect 3079 4535 3080 4539
rect 3074 4534 3080 4535
rect 3314 4539 3320 4540
rect 3314 4535 3315 4539
rect 3319 4535 3320 4539
rect 3314 4534 3320 4535
rect 3468 4532 3470 4586
rect 3564 4540 3566 4601
rect 3640 4592 3642 4714
rect 3650 4705 3656 4706
rect 3650 4701 3651 4705
rect 3655 4701 3656 4705
rect 3650 4700 3656 4701
rect 3652 4607 3654 4700
rect 3772 4648 3774 4714
rect 3798 4704 3804 4705
rect 3798 4700 3799 4704
rect 3803 4700 3804 4704
rect 3798 4699 3804 4700
rect 3770 4647 3776 4648
rect 3770 4643 3771 4647
rect 3775 4643 3776 4647
rect 3770 4642 3776 4643
rect 3800 4607 3802 4699
rect 3840 4635 3842 4719
rect 3984 4656 3986 4794
rect 4104 4771 4106 4795
rect 4328 4771 4330 4795
rect 4426 4794 4432 4795
rect 4536 4771 4538 4795
rect 4103 4770 4107 4771
rect 4103 4765 4107 4766
rect 4327 4770 4331 4771
rect 4327 4765 4331 4766
rect 4535 4770 4539 4771
rect 4535 4765 4539 4766
rect 4604 4756 4606 4858
rect 4632 4800 4634 4866
rect 4700 4816 4702 4877
rect 4752 4868 4754 4982
rect 4826 4973 4832 4974
rect 4826 4969 4827 4973
rect 4831 4969 4832 4973
rect 4826 4968 4832 4969
rect 4828 4883 4830 4968
rect 4952 4916 4954 4982
rect 4968 4924 4970 5058
rect 5128 5019 5130 5059
rect 5662 5058 5668 5059
rect 5664 5019 5666 5058
rect 5039 5018 5043 5019
rect 5039 5013 5043 5014
rect 5127 5018 5131 5019
rect 5127 5013 5131 5014
rect 5215 5018 5219 5019
rect 5215 5013 5219 5014
rect 5391 5018 5395 5019
rect 5391 5013 5395 5014
rect 5543 5018 5547 5019
rect 5543 5013 5547 5014
rect 5663 5018 5667 5019
rect 5663 5013 5667 5014
rect 5040 4989 5042 5013
rect 5216 4989 5218 5013
rect 5392 4989 5394 5013
rect 5544 4989 5546 5013
rect 5664 4990 5666 5013
rect 5662 4989 5668 4990
rect 5038 4988 5044 4989
rect 5214 4988 5220 4989
rect 5390 4988 5396 4989
rect 5038 4984 5039 4988
rect 5043 4984 5044 4988
rect 5038 4983 5044 4984
rect 5150 4987 5156 4988
rect 5150 4983 5151 4987
rect 5155 4983 5156 4987
rect 5214 4984 5215 4988
rect 5219 4984 5220 4988
rect 5214 4983 5220 4984
rect 5314 4987 5320 4988
rect 5314 4983 5315 4987
rect 5319 4983 5320 4987
rect 5390 4984 5391 4988
rect 5395 4984 5396 4988
rect 5390 4983 5396 4984
rect 5542 4988 5548 4989
rect 5542 4984 5543 4988
rect 5547 4984 5548 4988
rect 5542 4983 5548 4984
rect 5634 4987 5640 4988
rect 5634 4983 5635 4987
rect 5639 4983 5640 4987
rect 5662 4985 5663 4989
rect 5667 4985 5668 4989
rect 5662 4984 5668 4985
rect 5150 4982 5156 4983
rect 5314 4982 5320 4983
rect 5634 4982 5640 4983
rect 5010 4973 5016 4974
rect 5010 4969 5011 4973
rect 5015 4969 5016 4973
rect 5010 4968 5016 4969
rect 4966 4923 4972 4924
rect 4966 4919 4967 4923
rect 4971 4919 4972 4923
rect 4966 4918 4972 4919
rect 4950 4915 4956 4916
rect 4950 4911 4951 4915
rect 4955 4911 4956 4915
rect 4950 4910 4956 4911
rect 5012 4883 5014 4968
rect 5152 4924 5154 4982
rect 5186 4973 5192 4974
rect 5186 4969 5187 4973
rect 5191 4969 5192 4973
rect 5186 4968 5192 4969
rect 5150 4923 5156 4924
rect 5150 4919 5151 4923
rect 5155 4919 5156 4923
rect 5150 4918 5156 4919
rect 5188 4883 5190 4968
rect 5316 4924 5318 4982
rect 5362 4973 5368 4974
rect 5362 4969 5363 4973
rect 5367 4969 5368 4973
rect 5362 4968 5368 4969
rect 5514 4973 5520 4974
rect 5514 4969 5515 4973
rect 5519 4969 5520 4973
rect 5514 4968 5520 4969
rect 5314 4923 5320 4924
rect 5314 4919 5315 4923
rect 5319 4919 5320 4923
rect 5314 4918 5320 4919
rect 5364 4883 5366 4968
rect 5494 4915 5500 4916
rect 5494 4911 5495 4915
rect 5499 4911 5500 4915
rect 5494 4910 5500 4911
rect 4827 4882 4831 4883
rect 4827 4877 4831 4878
rect 4875 4882 4879 4883
rect 4875 4877 4879 4878
rect 5011 4882 5015 4883
rect 5011 4877 5015 4878
rect 5043 4882 5047 4883
rect 5043 4877 5047 4878
rect 5187 4882 5191 4883
rect 5187 4877 5191 4878
rect 5211 4882 5215 4883
rect 5211 4877 5215 4878
rect 5363 4882 5367 4883
rect 5363 4877 5367 4878
rect 5371 4882 5375 4883
rect 5371 4877 5375 4878
rect 4750 4867 4756 4868
rect 4750 4863 4751 4867
rect 4755 4863 4756 4867
rect 4750 4862 4756 4863
rect 4876 4816 4878 4877
rect 4882 4863 4888 4864
rect 4882 4859 4883 4863
rect 4887 4859 4888 4863
rect 4882 4858 4888 4859
rect 4698 4815 4704 4816
rect 4698 4811 4699 4815
rect 4703 4811 4704 4815
rect 4698 4810 4704 4811
rect 4874 4815 4880 4816
rect 4874 4811 4875 4815
rect 4879 4811 4880 4815
rect 4874 4810 4880 4811
rect 4726 4800 4732 4801
rect 4884 4800 4886 4858
rect 5044 4816 5046 4877
rect 5050 4863 5056 4864
rect 5050 4859 5051 4863
rect 5055 4859 5056 4863
rect 5050 4858 5056 4859
rect 5042 4815 5048 4816
rect 5042 4811 5043 4815
rect 5047 4811 5048 4815
rect 5042 4810 5048 4811
rect 4902 4800 4908 4801
rect 5052 4800 5054 4858
rect 5212 4816 5214 4877
rect 5330 4867 5336 4868
rect 5330 4863 5331 4867
rect 5335 4863 5336 4867
rect 5330 4862 5336 4863
rect 5210 4815 5216 4816
rect 5210 4811 5211 4815
rect 5215 4811 5216 4815
rect 5210 4810 5216 4811
rect 5070 4800 5076 4801
rect 5238 4800 5244 4801
rect 4630 4799 4636 4800
rect 4630 4795 4631 4799
rect 4635 4795 4636 4799
rect 4726 4796 4727 4800
rect 4731 4796 4732 4800
rect 4726 4795 4732 4796
rect 4882 4799 4888 4800
rect 4882 4795 4883 4799
rect 4887 4795 4888 4799
rect 4902 4796 4903 4800
rect 4907 4796 4908 4800
rect 4902 4795 4908 4796
rect 5050 4799 5056 4800
rect 5050 4795 5051 4799
rect 5055 4795 5056 4799
rect 5070 4796 5071 4800
rect 5075 4796 5076 4800
rect 5070 4795 5076 4796
rect 5166 4799 5172 4800
rect 5166 4795 5167 4799
rect 5171 4795 5172 4799
rect 5238 4796 5239 4800
rect 5243 4796 5244 4800
rect 5238 4795 5244 4796
rect 4630 4794 4636 4795
rect 4728 4771 4730 4795
rect 4882 4794 4888 4795
rect 4904 4771 4906 4795
rect 5050 4794 5056 4795
rect 5072 4771 5074 4795
rect 5166 4794 5172 4795
rect 4727 4770 4731 4771
rect 4727 4765 4731 4766
rect 4903 4770 4907 4771
rect 4903 4765 4907 4766
rect 4943 4770 4947 4771
rect 4943 4765 4947 4766
rect 5071 4770 5075 4771
rect 5071 4765 5075 4766
rect 5087 4770 5091 4771
rect 5087 4765 5091 4766
rect 4602 4755 4608 4756
rect 4602 4751 4603 4755
rect 4607 4751 4608 4755
rect 4602 4750 4608 4751
rect 4944 4741 4946 4765
rect 5088 4741 5090 4765
rect 4942 4740 4948 4741
rect 4942 4736 4943 4740
rect 4947 4736 4948 4740
rect 4942 4735 4948 4736
rect 5086 4740 5092 4741
rect 5086 4736 5087 4740
rect 5091 4736 5092 4740
rect 5086 4735 5092 4736
rect 4914 4725 4920 4726
rect 4914 4721 4915 4725
rect 4919 4721 4920 4725
rect 4914 4720 4920 4721
rect 5058 4725 5064 4726
rect 5058 4721 5059 4725
rect 5063 4721 5064 4725
rect 5058 4720 5064 4721
rect 3982 4655 3988 4656
rect 3982 4651 3983 4655
rect 3987 4651 3988 4655
rect 3982 4650 3988 4651
rect 4916 4635 4918 4720
rect 5060 4635 5062 4720
rect 5168 4676 5170 4794
rect 5240 4771 5242 4795
rect 5239 4770 5243 4771
rect 5239 4765 5243 4766
rect 5240 4741 5242 4765
rect 5238 4740 5244 4741
rect 5332 4740 5334 4862
rect 5372 4816 5374 4877
rect 5378 4863 5384 4864
rect 5378 4859 5379 4863
rect 5383 4859 5384 4863
rect 5378 4858 5384 4859
rect 5370 4815 5376 4816
rect 5370 4811 5371 4815
rect 5375 4811 5376 4815
rect 5370 4810 5376 4811
rect 5380 4800 5382 4858
rect 5398 4800 5404 4801
rect 5496 4800 5498 4910
rect 5516 4883 5518 4968
rect 5515 4882 5519 4883
rect 5515 4877 5519 4878
rect 5516 4816 5518 4877
rect 5636 4868 5638 4982
rect 5662 4972 5668 4973
rect 5662 4968 5663 4972
rect 5667 4968 5668 4972
rect 5662 4967 5668 4968
rect 5664 4883 5666 4967
rect 5663 4882 5667 4883
rect 5663 4877 5667 4878
rect 5634 4867 5640 4868
rect 5634 4863 5635 4867
rect 5639 4863 5640 4867
rect 5634 4862 5640 4863
rect 5664 4817 5666 4877
rect 5662 4816 5668 4817
rect 5514 4815 5520 4816
rect 5514 4811 5515 4815
rect 5519 4811 5520 4815
rect 5662 4812 5663 4816
rect 5667 4812 5668 4816
rect 5662 4811 5668 4812
rect 5514 4810 5520 4811
rect 5542 4800 5548 4801
rect 5378 4799 5384 4800
rect 5378 4795 5379 4799
rect 5383 4795 5384 4799
rect 5398 4796 5399 4800
rect 5403 4796 5404 4800
rect 5398 4795 5404 4796
rect 5494 4799 5500 4800
rect 5494 4795 5495 4799
rect 5499 4795 5500 4799
rect 5542 4796 5543 4800
rect 5547 4796 5548 4800
rect 5542 4795 5548 4796
rect 5638 4799 5644 4800
rect 5638 4795 5639 4799
rect 5643 4795 5644 4799
rect 5378 4794 5384 4795
rect 5400 4771 5402 4795
rect 5494 4794 5500 4795
rect 5544 4771 5546 4795
rect 5638 4794 5644 4795
rect 5662 4799 5668 4800
rect 5662 4795 5663 4799
rect 5667 4795 5668 4799
rect 5662 4794 5668 4795
rect 5399 4770 5403 4771
rect 5399 4765 5403 4766
rect 5543 4770 5547 4771
rect 5543 4765 5547 4766
rect 5400 4741 5402 4765
rect 5544 4741 5546 4765
rect 5398 4740 5404 4741
rect 5542 4740 5548 4741
rect 5238 4736 5239 4740
rect 5243 4736 5244 4740
rect 5238 4735 5244 4736
rect 5330 4739 5336 4740
rect 5330 4735 5331 4739
rect 5335 4735 5336 4739
rect 5398 4736 5399 4740
rect 5403 4736 5404 4740
rect 5398 4735 5404 4736
rect 5490 4739 5496 4740
rect 5490 4735 5491 4739
rect 5495 4735 5496 4739
rect 5542 4736 5543 4740
rect 5547 4736 5548 4740
rect 5542 4735 5548 4736
rect 5330 4734 5336 4735
rect 5490 4734 5496 4735
rect 5210 4725 5216 4726
rect 5210 4721 5211 4725
rect 5215 4721 5216 4725
rect 5210 4720 5216 4721
rect 5370 4725 5376 4726
rect 5370 4721 5371 4725
rect 5375 4721 5376 4725
rect 5370 4720 5376 4721
rect 5166 4675 5172 4676
rect 5166 4671 5167 4675
rect 5171 4671 5172 4675
rect 5166 4670 5172 4671
rect 5212 4635 5214 4720
rect 5372 4635 5374 4720
rect 5462 4675 5468 4676
rect 5462 4671 5463 4675
rect 5467 4671 5468 4675
rect 5462 4670 5468 4671
rect 3839 4634 3843 4635
rect 3839 4629 3843 4630
rect 4771 4634 4775 4635
rect 4771 4629 4775 4630
rect 4915 4634 4919 4635
rect 4915 4629 4919 4630
rect 4955 4634 4959 4635
rect 4955 4629 4959 4630
rect 5059 4634 5063 4635
rect 5059 4629 5063 4630
rect 5147 4634 5151 4635
rect 5147 4629 5151 4630
rect 5211 4634 5215 4635
rect 5211 4629 5215 4630
rect 5339 4634 5343 4635
rect 5339 4629 5343 4630
rect 5371 4634 5375 4635
rect 5371 4629 5375 4630
rect 3651 4606 3655 4607
rect 3651 4601 3655 4602
rect 3799 4606 3803 4607
rect 3799 4601 3803 4602
rect 3638 4591 3644 4592
rect 3638 4587 3639 4591
rect 3643 4587 3644 4591
rect 3638 4586 3644 4587
rect 3800 4541 3802 4601
rect 3840 4569 3842 4629
rect 3838 4568 3844 4569
rect 4772 4568 4774 4629
rect 4866 4615 4872 4616
rect 4866 4611 4867 4615
rect 4871 4611 4872 4615
rect 4866 4610 4872 4611
rect 4868 4573 4870 4610
rect 4867 4572 4871 4573
rect 4956 4568 4958 4629
rect 4962 4615 4968 4616
rect 4962 4611 4963 4615
rect 4967 4611 4968 4615
rect 4962 4610 4968 4611
rect 3838 4564 3839 4568
rect 3843 4564 3844 4568
rect 3838 4563 3844 4564
rect 4770 4567 4776 4568
rect 4867 4567 4871 4568
rect 4954 4567 4960 4568
rect 4770 4563 4771 4567
rect 4775 4563 4776 4567
rect 4770 4562 4776 4563
rect 4954 4563 4955 4567
rect 4959 4563 4960 4567
rect 4954 4562 4960 4563
rect 4798 4552 4804 4553
rect 4964 4552 4966 4610
rect 5148 4568 5150 4629
rect 5154 4615 5160 4616
rect 5154 4611 5155 4615
rect 5159 4611 5160 4615
rect 5154 4610 5160 4611
rect 5146 4567 5152 4568
rect 5146 4563 5147 4567
rect 5151 4563 5152 4567
rect 5146 4562 5152 4563
rect 4982 4552 4988 4553
rect 5156 4552 5158 4610
rect 5340 4568 5342 4629
rect 5346 4615 5352 4616
rect 5346 4611 5347 4615
rect 5351 4611 5352 4615
rect 5346 4610 5352 4611
rect 5338 4567 5344 4568
rect 5338 4563 5339 4567
rect 5343 4563 5344 4567
rect 5338 4562 5344 4563
rect 5174 4552 5180 4553
rect 5348 4552 5350 4610
rect 5423 4572 5427 4573
rect 5423 4567 5427 4568
rect 5366 4552 5372 4553
rect 3838 4551 3844 4552
rect 3838 4547 3839 4551
rect 3843 4547 3844 4551
rect 4798 4548 4799 4552
rect 4803 4548 4804 4552
rect 4798 4547 4804 4548
rect 4962 4551 4968 4552
rect 4962 4547 4963 4551
rect 4967 4547 4968 4551
rect 4982 4548 4983 4552
rect 4987 4548 4988 4552
rect 4982 4547 4988 4548
rect 5154 4551 5160 4552
rect 5154 4547 5155 4551
rect 5159 4547 5160 4551
rect 5174 4548 5175 4552
rect 5179 4548 5180 4552
rect 5174 4547 5180 4548
rect 5346 4551 5352 4552
rect 5346 4547 5347 4551
rect 5351 4547 5352 4551
rect 5366 4548 5367 4552
rect 5371 4548 5372 4552
rect 5366 4547 5372 4548
rect 3838 4546 3844 4547
rect 3798 4540 3804 4541
rect 3562 4539 3568 4540
rect 3562 4535 3563 4539
rect 3567 4535 3568 4539
rect 3798 4536 3799 4540
rect 3803 4536 3804 4540
rect 3798 4535 3804 4536
rect 3562 4534 3568 4535
rect 3066 4531 3072 4532
rect 3066 4527 3067 4531
rect 3071 4527 3072 4531
rect 3066 4526 3072 4527
rect 3466 4531 3472 4532
rect 3466 4527 3467 4531
rect 3471 4527 3472 4531
rect 3466 4526 3472 4527
rect 2854 4524 2860 4525
rect 3102 4524 3108 4525
rect 2854 4520 2855 4524
rect 2859 4520 2860 4524
rect 2854 4519 2860 4520
rect 2950 4523 2956 4524
rect 2950 4519 2951 4523
rect 2955 4519 2956 4523
rect 3102 4520 3103 4524
rect 3107 4520 3108 4524
rect 3102 4519 3108 4520
rect 3342 4524 3348 4525
rect 3342 4520 3343 4524
rect 3347 4520 3348 4524
rect 3342 4519 3348 4520
rect 3590 4524 3596 4525
rect 3590 4520 3591 4524
rect 3595 4520 3596 4524
rect 3590 4519 3596 4520
rect 3798 4523 3804 4524
rect 3798 4519 3799 4523
rect 3803 4519 3804 4523
rect 2856 4487 2858 4519
rect 2950 4518 2956 4519
rect 2783 4486 2787 4487
rect 2783 4481 2787 4482
rect 2855 4486 2859 4487
rect 2855 4481 2859 4482
rect 2784 4457 2786 4481
rect 2782 4456 2788 4457
rect 2542 4452 2543 4456
rect 2547 4452 2548 4456
rect 2542 4451 2548 4452
rect 2638 4455 2644 4456
rect 2638 4451 2639 4455
rect 2643 4451 2644 4455
rect 2782 4452 2783 4456
rect 2787 4452 2788 4456
rect 2782 4451 2788 4452
rect 2638 4450 2644 4451
rect 2514 4441 2520 4442
rect 1974 4440 1980 4441
rect 1974 4436 1975 4440
rect 1979 4436 1980 4440
rect 2514 4437 2515 4441
rect 2519 4437 2520 4441
rect 2514 4436 2520 4437
rect 2754 4441 2760 4442
rect 2754 4437 2755 4441
rect 2759 4437 2760 4441
rect 2754 4436 2760 4437
rect 1974 4435 1980 4436
rect 1935 4434 1939 4435
rect 1935 4429 1939 4430
rect 1936 4406 1938 4429
rect 1934 4405 1940 4406
rect 1926 4403 1932 4404
rect 1926 4399 1927 4403
rect 1931 4399 1932 4403
rect 1934 4401 1935 4405
rect 1939 4401 1940 4405
rect 1934 4400 1940 4401
rect 1926 4398 1932 4399
rect 1928 4348 1930 4398
rect 1934 4388 1940 4389
rect 1934 4384 1935 4388
rect 1939 4384 1940 4388
rect 1934 4383 1940 4384
rect 1926 4347 1932 4348
rect 1926 4343 1927 4347
rect 1931 4343 1932 4347
rect 1926 4342 1932 4343
rect 1910 4331 1916 4332
rect 1910 4327 1911 4331
rect 1915 4327 1916 4331
rect 1910 4326 1916 4327
rect 1936 4303 1938 4383
rect 1976 4363 1978 4435
rect 2516 4363 2518 4436
rect 2756 4363 2758 4436
rect 2952 4400 2954 4518
rect 3104 4487 3106 4519
rect 3344 4487 3346 4519
rect 3592 4487 3594 4519
rect 3798 4518 3804 4519
rect 3800 4487 3802 4518
rect 3840 4511 3842 4546
rect 4800 4511 4802 4547
rect 4962 4546 4968 4547
rect 4984 4511 4986 4547
rect 5154 4546 5160 4547
rect 5176 4511 5178 4547
rect 5346 4546 5352 4547
rect 5368 4511 5370 4547
rect 3839 4510 3843 4511
rect 3839 4505 3843 4506
rect 4487 4510 4491 4511
rect 4487 4505 4491 4506
rect 4671 4510 4675 4511
rect 4671 4505 4675 4506
rect 4799 4510 4803 4511
rect 4799 4505 4803 4506
rect 4879 4510 4883 4511
rect 4879 4505 4883 4506
rect 4983 4510 4987 4511
rect 4983 4505 4987 4506
rect 5095 4510 5099 4511
rect 5095 4505 5099 4506
rect 5175 4510 5179 4511
rect 5175 4505 5179 4506
rect 5327 4510 5331 4511
rect 5327 4505 5331 4506
rect 5367 4510 5371 4511
rect 5367 4505 5371 4506
rect 3015 4486 3019 4487
rect 3015 4481 3019 4482
rect 3103 4486 3107 4487
rect 3103 4481 3107 4482
rect 3247 4486 3251 4487
rect 3247 4481 3251 4482
rect 3343 4486 3347 4487
rect 3343 4481 3347 4482
rect 3471 4486 3475 4487
rect 3471 4481 3475 4482
rect 3591 4486 3595 4487
rect 3591 4481 3595 4482
rect 3679 4486 3683 4487
rect 3679 4481 3683 4482
rect 3799 4486 3803 4487
rect 3840 4482 3842 4505
rect 3799 4481 3803 4482
rect 3838 4481 3844 4482
rect 4488 4481 4490 4505
rect 4672 4481 4674 4505
rect 4880 4481 4882 4505
rect 5096 4481 5098 4505
rect 5328 4481 5330 4505
rect 3016 4457 3018 4481
rect 3248 4457 3250 4481
rect 3472 4457 3474 4481
rect 3680 4457 3682 4481
rect 3800 4458 3802 4481
rect 3838 4477 3839 4481
rect 3843 4477 3844 4481
rect 3838 4476 3844 4477
rect 4486 4480 4492 4481
rect 4486 4476 4487 4480
rect 4491 4476 4492 4480
rect 4486 4475 4492 4476
rect 4670 4480 4676 4481
rect 4670 4476 4671 4480
rect 4675 4476 4676 4480
rect 4670 4475 4676 4476
rect 4878 4480 4884 4481
rect 5094 4480 5100 4481
rect 4878 4476 4879 4480
rect 4883 4476 4884 4480
rect 4878 4475 4884 4476
rect 4978 4479 4984 4480
rect 4978 4475 4979 4479
rect 4983 4475 4984 4479
rect 5094 4476 5095 4480
rect 5099 4476 5100 4480
rect 5094 4475 5100 4476
rect 5326 4480 5332 4481
rect 5424 4480 5426 4567
rect 5464 4552 5466 4670
rect 5492 4668 5494 4734
rect 5514 4725 5520 4726
rect 5514 4721 5515 4725
rect 5519 4721 5520 4725
rect 5514 4720 5520 4721
rect 5490 4667 5496 4668
rect 5490 4663 5491 4667
rect 5495 4663 5496 4667
rect 5490 4662 5496 4663
rect 5516 4635 5518 4720
rect 5640 4676 5642 4794
rect 5664 4771 5666 4794
rect 5663 4770 5667 4771
rect 5663 4765 5667 4766
rect 5664 4742 5666 4765
rect 5662 4741 5668 4742
rect 5662 4737 5663 4741
rect 5667 4737 5668 4741
rect 5662 4736 5668 4737
rect 5662 4724 5668 4725
rect 5662 4720 5663 4724
rect 5667 4720 5668 4724
rect 5662 4719 5668 4720
rect 5638 4675 5644 4676
rect 5638 4671 5639 4675
rect 5643 4671 5644 4675
rect 5638 4670 5644 4671
rect 5664 4635 5666 4719
rect 5515 4634 5519 4635
rect 5515 4629 5519 4630
rect 5663 4634 5667 4635
rect 5663 4629 5667 4630
rect 5516 4568 5518 4629
rect 5664 4569 5666 4629
rect 5662 4568 5668 4569
rect 5514 4567 5520 4568
rect 5514 4563 5515 4567
rect 5519 4563 5520 4567
rect 5662 4564 5663 4568
rect 5667 4564 5668 4568
rect 5662 4563 5668 4564
rect 5514 4562 5520 4563
rect 5542 4552 5548 4553
rect 5462 4551 5468 4552
rect 5462 4547 5463 4551
rect 5467 4547 5468 4551
rect 5542 4548 5543 4552
rect 5547 4548 5548 4552
rect 5542 4547 5548 4548
rect 5642 4551 5648 4552
rect 5642 4547 5643 4551
rect 5647 4547 5648 4551
rect 5462 4546 5468 4547
rect 5544 4511 5546 4547
rect 5642 4546 5648 4547
rect 5662 4551 5668 4552
rect 5662 4547 5663 4551
rect 5667 4547 5668 4551
rect 5662 4546 5668 4547
rect 5543 4510 5547 4511
rect 5543 4505 5547 4506
rect 5544 4481 5546 4505
rect 5542 4480 5548 4481
rect 5326 4476 5327 4480
rect 5331 4476 5332 4480
rect 5326 4475 5332 4476
rect 5422 4479 5428 4480
rect 5422 4475 5423 4479
rect 5427 4475 5428 4479
rect 5542 4476 5543 4480
rect 5547 4476 5548 4480
rect 5542 4475 5548 4476
rect 5634 4479 5640 4480
rect 5634 4475 5635 4479
rect 5639 4475 5640 4479
rect 4978 4474 4984 4475
rect 5422 4474 5428 4475
rect 5634 4474 5640 4475
rect 4458 4465 4464 4466
rect 3838 4464 3844 4465
rect 3838 4460 3839 4464
rect 3843 4460 3844 4464
rect 4458 4461 4459 4465
rect 4463 4461 4464 4465
rect 4458 4460 4464 4461
rect 4642 4465 4648 4466
rect 4642 4461 4643 4465
rect 4647 4461 4648 4465
rect 4642 4460 4648 4461
rect 4850 4465 4856 4466
rect 4850 4461 4851 4465
rect 4855 4461 4856 4465
rect 4850 4460 4856 4461
rect 3838 4459 3844 4460
rect 3798 4457 3804 4458
rect 3014 4456 3020 4457
rect 3246 4456 3252 4457
rect 3470 4456 3476 4457
rect 3678 4456 3684 4457
rect 3014 4452 3015 4456
rect 3019 4452 3020 4456
rect 3014 4451 3020 4452
rect 3126 4455 3132 4456
rect 3126 4451 3127 4455
rect 3131 4451 3132 4455
rect 3246 4452 3247 4456
rect 3251 4452 3252 4456
rect 3246 4451 3252 4452
rect 3346 4455 3352 4456
rect 3346 4451 3347 4455
rect 3351 4451 3352 4455
rect 3470 4452 3471 4456
rect 3475 4452 3476 4456
rect 3470 4451 3476 4452
rect 3570 4455 3576 4456
rect 3570 4451 3571 4455
rect 3575 4451 3576 4455
rect 3678 4452 3679 4456
rect 3683 4452 3684 4456
rect 3678 4451 3684 4452
rect 3770 4455 3776 4456
rect 3770 4451 3771 4455
rect 3775 4451 3776 4455
rect 3798 4453 3799 4457
rect 3803 4453 3804 4457
rect 3798 4452 3804 4453
rect 3126 4450 3132 4451
rect 3346 4450 3352 4451
rect 3570 4450 3576 4451
rect 3770 4450 3776 4451
rect 2986 4441 2992 4442
rect 2986 4437 2987 4441
rect 2991 4437 2992 4441
rect 2986 4436 2992 4437
rect 2950 4399 2956 4400
rect 2950 4395 2951 4399
rect 2955 4395 2956 4399
rect 2950 4394 2956 4395
rect 2926 4383 2932 4384
rect 2926 4379 2927 4383
rect 2931 4379 2932 4383
rect 2926 4378 2932 4379
rect 1975 4362 1979 4363
rect 1975 4357 1979 4358
rect 1995 4362 1999 4363
rect 1995 4357 1999 4358
rect 2379 4362 2383 4363
rect 2379 4357 2383 4358
rect 2515 4362 2519 4363
rect 2515 4357 2519 4358
rect 2755 4362 2759 4363
rect 2755 4357 2759 4358
rect 2803 4362 2807 4363
rect 2803 4357 2807 4358
rect 1595 4302 1599 4303
rect 1595 4297 1599 4298
rect 1643 4302 1647 4303
rect 1643 4297 1647 4298
rect 1787 4302 1791 4303
rect 1787 4297 1791 4298
rect 1935 4302 1939 4303
rect 1935 4297 1939 4298
rect 1976 4297 1978 4357
rect 1596 4236 1598 4297
rect 1714 4291 1720 4292
rect 1714 4287 1715 4291
rect 1719 4287 1720 4291
rect 1714 4286 1720 4287
rect 1594 4235 1600 4236
rect 1594 4231 1595 4235
rect 1599 4231 1600 4235
rect 1594 4230 1600 4231
rect 1622 4220 1628 4221
rect 1716 4220 1718 4286
rect 1878 4279 1884 4280
rect 1878 4275 1879 4279
rect 1883 4275 1884 4279
rect 1878 4274 1884 4275
rect 1446 4216 1447 4220
rect 1451 4216 1452 4220
rect 1446 4215 1452 4216
rect 1542 4219 1548 4220
rect 1542 4215 1543 4219
rect 1547 4215 1548 4219
rect 1622 4216 1623 4220
rect 1627 4216 1628 4220
rect 1622 4215 1628 4216
rect 1714 4219 1720 4220
rect 1714 4215 1715 4219
rect 1719 4215 1720 4219
rect 110 4214 116 4215
rect 112 4187 114 4214
rect 656 4187 658 4215
rect 778 4214 784 4215
rect 800 4187 802 4215
rect 894 4214 900 4215
rect 896 4211 898 4214
rect 888 4209 898 4211
rect 111 4186 115 4187
rect 111 4181 115 4182
rect 519 4186 523 4187
rect 519 4181 523 4182
rect 655 4186 659 4187
rect 655 4181 659 4182
rect 703 4186 707 4187
rect 703 4181 707 4182
rect 799 4186 803 4187
rect 799 4181 803 4182
rect 112 4158 114 4181
rect 110 4157 116 4158
rect 520 4157 522 4181
rect 704 4157 706 4181
rect 110 4153 111 4157
rect 115 4153 116 4157
rect 110 4152 116 4153
rect 518 4156 524 4157
rect 518 4152 519 4156
rect 523 4152 524 4156
rect 518 4151 524 4152
rect 702 4156 708 4157
rect 702 4152 703 4156
rect 707 4152 708 4156
rect 702 4151 708 4152
rect 802 4155 808 4156
rect 802 4151 803 4155
rect 807 4151 808 4155
rect 802 4150 808 4151
rect 490 4141 496 4142
rect 110 4140 116 4141
rect 110 4136 111 4140
rect 115 4136 116 4140
rect 490 4137 491 4141
rect 495 4137 496 4141
rect 490 4136 496 4137
rect 674 4141 680 4142
rect 674 4137 675 4141
rect 679 4137 680 4141
rect 674 4136 680 4137
rect 110 4135 116 4136
rect 112 4075 114 4135
rect 492 4075 494 4136
rect 586 4127 592 4128
rect 586 4123 587 4127
rect 591 4123 592 4127
rect 586 4122 592 4123
rect 588 4092 590 4122
rect 586 4091 592 4092
rect 586 4087 587 4091
rect 591 4087 592 4091
rect 586 4086 592 4087
rect 676 4075 678 4136
rect 111 4074 115 4075
rect 111 4069 115 4070
rect 131 4074 135 4075
rect 131 4069 135 4070
rect 339 4074 343 4075
rect 339 4069 343 4070
rect 491 4074 495 4075
rect 491 4069 495 4070
rect 595 4074 599 4075
rect 595 4069 599 4070
rect 675 4074 679 4075
rect 675 4069 679 4070
rect 112 4009 114 4069
rect 110 4008 116 4009
rect 132 4008 134 4069
rect 340 4008 342 4069
rect 462 4063 468 4064
rect 462 4059 463 4063
rect 467 4059 468 4063
rect 462 4058 468 4059
rect 110 4004 111 4008
rect 115 4004 116 4008
rect 110 4003 116 4004
rect 130 4007 136 4008
rect 130 4003 131 4007
rect 135 4003 136 4007
rect 130 4002 136 4003
rect 338 4007 344 4008
rect 338 4003 339 4007
rect 343 4003 344 4007
rect 338 4002 344 4003
rect 158 3992 164 3993
rect 366 3992 372 3993
rect 464 3992 466 4058
rect 596 4008 598 4069
rect 804 4060 806 4150
rect 866 4141 872 4142
rect 866 4137 867 4141
rect 871 4137 872 4141
rect 866 4136 872 4137
rect 868 4075 870 4136
rect 888 4092 890 4209
rect 952 4187 954 4215
rect 1046 4214 1052 4215
rect 1112 4187 1114 4215
rect 1206 4214 1212 4215
rect 1280 4187 1282 4215
rect 1448 4187 1450 4215
rect 1542 4214 1548 4215
rect 1624 4187 1626 4215
rect 1714 4214 1720 4215
rect 895 4186 899 4187
rect 895 4181 899 4182
rect 951 4186 955 4187
rect 951 4181 955 4182
rect 1103 4186 1107 4187
rect 1103 4181 1107 4182
rect 1111 4186 1115 4187
rect 1111 4181 1115 4182
rect 1279 4186 1283 4187
rect 1279 4181 1283 4182
rect 1327 4186 1331 4187
rect 1327 4181 1331 4182
rect 1447 4186 1451 4187
rect 1447 4181 1451 4182
rect 1551 4186 1555 4187
rect 1551 4181 1555 4182
rect 1623 4186 1627 4187
rect 1623 4181 1627 4182
rect 1783 4186 1787 4187
rect 1783 4181 1787 4182
rect 896 4157 898 4181
rect 1104 4157 1106 4181
rect 1328 4157 1330 4181
rect 1552 4157 1554 4181
rect 1784 4157 1786 4181
rect 894 4156 900 4157
rect 1102 4156 1108 4157
rect 1326 4156 1332 4157
rect 1550 4156 1556 4157
rect 1782 4156 1788 4157
rect 1880 4156 1882 4274
rect 1936 4237 1938 4297
rect 1974 4296 1980 4297
rect 1996 4296 1998 4357
rect 2380 4296 2382 4357
rect 2386 4343 2392 4344
rect 2386 4339 2387 4343
rect 2391 4339 2392 4343
rect 2386 4338 2392 4339
rect 1974 4292 1975 4296
rect 1979 4292 1980 4296
rect 1974 4291 1980 4292
rect 1994 4295 2000 4296
rect 1994 4291 1995 4295
rect 1999 4291 2000 4295
rect 1994 4290 2000 4291
rect 2378 4295 2384 4296
rect 2378 4291 2379 4295
rect 2383 4291 2384 4295
rect 2378 4290 2384 4291
rect 2022 4280 2028 4281
rect 2388 4280 2390 4338
rect 2804 4296 2806 4357
rect 2802 4295 2808 4296
rect 2802 4291 2803 4295
rect 2807 4291 2808 4295
rect 2802 4290 2808 4291
rect 2406 4280 2412 4281
rect 2830 4280 2836 4281
rect 2928 4280 2930 4378
rect 2988 4363 2990 4436
rect 3128 4392 3130 4450
rect 3218 4441 3224 4442
rect 3218 4437 3219 4441
rect 3223 4437 3224 4441
rect 3218 4436 3224 4437
rect 3126 4391 3132 4392
rect 3126 4387 3127 4391
rect 3131 4387 3132 4391
rect 3126 4386 3132 4387
rect 3220 4363 3222 4436
rect 3348 4392 3350 4450
rect 3442 4441 3448 4442
rect 3442 4437 3443 4441
rect 3447 4437 3448 4441
rect 3442 4436 3448 4437
rect 3346 4391 3352 4392
rect 3346 4387 3347 4391
rect 3351 4387 3352 4391
rect 3346 4386 3352 4387
rect 3444 4363 3446 4436
rect 3572 4392 3574 4450
rect 3650 4441 3656 4442
rect 3650 4437 3651 4441
rect 3655 4437 3656 4441
rect 3650 4436 3656 4437
rect 3570 4391 3576 4392
rect 3570 4387 3571 4391
rect 3575 4387 3576 4391
rect 3570 4386 3576 4387
rect 3652 4363 3654 4436
rect 2987 4362 2991 4363
rect 2987 4357 2991 4358
rect 3219 4362 3223 4363
rect 3219 4357 3223 4358
rect 3235 4362 3239 4363
rect 3235 4357 3239 4358
rect 3443 4362 3447 4363
rect 3443 4357 3447 4358
rect 3651 4362 3655 4363
rect 3651 4357 3655 4358
rect 3236 4296 3238 4357
rect 3358 4351 3364 4352
rect 3358 4347 3359 4351
rect 3363 4347 3364 4351
rect 3358 4346 3364 4347
rect 3242 4343 3248 4344
rect 3242 4339 3243 4343
rect 3247 4339 3248 4343
rect 3242 4338 3248 4339
rect 3234 4295 3240 4296
rect 3234 4291 3235 4295
rect 3239 4291 3240 4295
rect 3234 4290 3240 4291
rect 1974 4279 1980 4280
rect 1974 4275 1975 4279
rect 1979 4275 1980 4279
rect 2022 4276 2023 4280
rect 2027 4276 2028 4280
rect 2022 4275 2028 4276
rect 2386 4279 2392 4280
rect 2386 4275 2387 4279
rect 2391 4275 2392 4279
rect 2406 4276 2407 4280
rect 2411 4276 2412 4280
rect 2406 4275 2412 4276
rect 2502 4279 2508 4280
rect 2502 4275 2503 4279
rect 2507 4275 2508 4279
rect 2830 4276 2831 4280
rect 2835 4276 2836 4280
rect 2830 4275 2836 4276
rect 2926 4279 2932 4280
rect 2926 4275 2927 4279
rect 2931 4275 2932 4279
rect 1974 4274 1980 4275
rect 1934 4236 1940 4237
rect 1934 4232 1935 4236
rect 1939 4232 1940 4236
rect 1934 4231 1940 4232
rect 1976 4223 1978 4274
rect 2024 4223 2026 4275
rect 2386 4274 2392 4275
rect 2408 4223 2410 4275
rect 2502 4274 2508 4275
rect 1975 4222 1979 4223
rect 1934 4219 1940 4220
rect 1934 4215 1935 4219
rect 1939 4215 1940 4219
rect 1975 4217 1979 4218
rect 2023 4222 2027 4223
rect 2023 4217 2027 4218
rect 2191 4222 2195 4223
rect 2191 4217 2195 4218
rect 2383 4222 2387 4223
rect 2383 4217 2387 4218
rect 2407 4222 2411 4223
rect 2407 4217 2411 4218
rect 1934 4214 1940 4215
rect 1936 4187 1938 4214
rect 1976 4194 1978 4217
rect 1974 4193 1980 4194
rect 2024 4193 2026 4217
rect 2192 4193 2194 4217
rect 2384 4193 2386 4217
rect 1974 4189 1975 4193
rect 1979 4189 1980 4193
rect 1974 4188 1980 4189
rect 2022 4192 2028 4193
rect 2190 4192 2196 4193
rect 2382 4192 2388 4193
rect 2022 4188 2023 4192
rect 2027 4188 2028 4192
rect 2022 4187 2028 4188
rect 2122 4191 2128 4192
rect 2122 4187 2123 4191
rect 2127 4187 2128 4191
rect 2190 4188 2191 4192
rect 2195 4188 2196 4192
rect 2190 4187 2196 4188
rect 2286 4191 2292 4192
rect 2286 4187 2287 4191
rect 2291 4187 2292 4191
rect 2382 4188 2383 4192
rect 2387 4188 2388 4192
rect 2382 4187 2388 4188
rect 2478 4191 2484 4192
rect 2478 4187 2479 4191
rect 2483 4187 2484 4191
rect 1935 4186 1939 4187
rect 2122 4186 2128 4187
rect 2286 4186 2292 4187
rect 2478 4186 2484 4187
rect 1935 4181 1939 4182
rect 1936 4158 1938 4181
rect 1994 4177 2000 4178
rect 1974 4176 1980 4177
rect 1974 4172 1975 4176
rect 1979 4172 1980 4176
rect 1994 4173 1995 4177
rect 1999 4173 2000 4177
rect 1994 4172 2000 4173
rect 1974 4171 1980 4172
rect 1934 4157 1940 4158
rect 894 4152 895 4156
rect 899 4152 900 4156
rect 894 4151 900 4152
rect 994 4155 1000 4156
rect 994 4151 995 4155
rect 999 4151 1000 4155
rect 1102 4152 1103 4156
rect 1107 4152 1108 4156
rect 1102 4151 1108 4152
rect 1202 4155 1208 4156
rect 1202 4151 1203 4155
rect 1207 4151 1208 4155
rect 1326 4152 1327 4156
rect 1331 4152 1332 4156
rect 1326 4151 1332 4152
rect 1418 4155 1424 4156
rect 1418 4151 1419 4155
rect 1423 4151 1424 4155
rect 1550 4152 1551 4156
rect 1555 4152 1556 4156
rect 1550 4151 1556 4152
rect 1650 4155 1656 4156
rect 1650 4151 1651 4155
rect 1655 4151 1656 4155
rect 1782 4152 1783 4156
rect 1787 4152 1788 4156
rect 1782 4151 1788 4152
rect 1878 4155 1884 4156
rect 1878 4151 1879 4155
rect 1883 4151 1884 4155
rect 1934 4153 1935 4157
rect 1939 4153 1940 4157
rect 1934 4152 1940 4153
rect 994 4150 1000 4151
rect 1202 4150 1208 4151
rect 1418 4150 1424 4151
rect 1650 4150 1656 4151
rect 1878 4150 1884 4151
rect 996 4092 998 4150
rect 1074 4141 1080 4142
rect 1074 4137 1075 4141
rect 1079 4137 1080 4141
rect 1074 4136 1080 4137
rect 886 4091 892 4092
rect 886 4087 887 4091
rect 891 4087 892 4091
rect 886 4086 892 4087
rect 994 4091 1000 4092
rect 994 4087 995 4091
rect 999 4087 1000 4091
rect 994 4086 1000 4087
rect 1076 4075 1078 4136
rect 1204 4092 1206 4150
rect 1298 4141 1304 4142
rect 1298 4137 1299 4141
rect 1303 4137 1304 4141
rect 1298 4136 1304 4137
rect 1202 4091 1208 4092
rect 1202 4087 1203 4091
rect 1207 4087 1208 4091
rect 1202 4086 1208 4087
rect 1300 4075 1302 4136
rect 1420 4128 1422 4150
rect 1522 4141 1528 4142
rect 1522 4137 1523 4141
rect 1527 4137 1528 4141
rect 1522 4136 1528 4137
rect 1418 4127 1424 4128
rect 1418 4123 1419 4127
rect 1423 4123 1424 4127
rect 1418 4122 1424 4123
rect 1524 4075 1526 4136
rect 1652 4092 1654 4150
rect 1754 4141 1760 4142
rect 1754 4137 1755 4141
rect 1759 4137 1760 4141
rect 1754 4136 1760 4137
rect 1934 4140 1940 4141
rect 1934 4136 1935 4140
rect 1939 4136 1940 4140
rect 1614 4091 1620 4092
rect 1614 4087 1615 4091
rect 1619 4087 1620 4091
rect 1614 4086 1620 4087
rect 1650 4091 1656 4092
rect 1650 4087 1651 4091
rect 1655 4087 1656 4091
rect 1650 4086 1656 4087
rect 867 4074 871 4075
rect 867 4069 871 4070
rect 875 4074 879 4075
rect 875 4069 879 4070
rect 1075 4074 1079 4075
rect 1075 4069 1079 4070
rect 1179 4074 1183 4075
rect 1179 4069 1183 4070
rect 1299 4074 1303 4075
rect 1299 4069 1303 4070
rect 1491 4074 1495 4075
rect 1491 4069 1495 4070
rect 1523 4074 1527 4075
rect 1523 4069 1527 4070
rect 794 4059 800 4060
rect 794 4055 795 4059
rect 799 4055 800 4059
rect 794 4054 800 4055
rect 802 4059 808 4060
rect 802 4055 803 4059
rect 807 4055 808 4059
rect 802 4054 808 4055
rect 594 4007 600 4008
rect 594 4003 595 4007
rect 599 4003 600 4007
rect 594 4002 600 4003
rect 796 4000 798 4054
rect 876 4008 878 4069
rect 1180 4008 1182 4069
rect 1186 4055 1192 4056
rect 1186 4051 1187 4055
rect 1191 4051 1192 4055
rect 1186 4050 1192 4051
rect 874 4007 880 4008
rect 874 4003 875 4007
rect 879 4003 880 4007
rect 874 4002 880 4003
rect 1178 4007 1184 4008
rect 1178 4003 1179 4007
rect 1183 4003 1184 4007
rect 1178 4002 1184 4003
rect 794 3999 800 4000
rect 794 3995 795 3999
rect 799 3995 800 3999
rect 794 3994 800 3995
rect 622 3992 628 3993
rect 110 3991 116 3992
rect 110 3987 111 3991
rect 115 3987 116 3991
rect 158 3988 159 3992
rect 163 3988 164 3992
rect 158 3987 164 3988
rect 254 3991 260 3992
rect 254 3987 255 3991
rect 259 3987 260 3991
rect 366 3988 367 3992
rect 371 3988 372 3992
rect 366 3987 372 3988
rect 462 3991 468 3992
rect 462 3987 463 3991
rect 467 3987 468 3991
rect 622 3988 623 3992
rect 627 3988 628 3992
rect 622 3987 628 3988
rect 902 3992 908 3993
rect 1188 3992 1190 4050
rect 1492 4008 1494 4069
rect 1586 4055 1592 4056
rect 1586 4051 1587 4055
rect 1591 4051 1592 4055
rect 1586 4050 1592 4051
rect 1588 4036 1590 4050
rect 1586 4035 1592 4036
rect 1586 4031 1587 4035
rect 1591 4031 1592 4035
rect 1586 4030 1592 4031
rect 1490 4007 1496 4008
rect 1490 4003 1491 4007
rect 1495 4003 1496 4007
rect 1490 4002 1496 4003
rect 1206 3992 1212 3993
rect 902 3988 903 3992
rect 907 3988 908 3992
rect 902 3987 908 3988
rect 1186 3991 1192 3992
rect 1186 3987 1187 3991
rect 1191 3987 1192 3991
rect 1206 3988 1207 3992
rect 1211 3988 1212 3992
rect 1206 3987 1212 3988
rect 1518 3992 1524 3993
rect 1616 3992 1618 4086
rect 1756 4075 1758 4136
rect 1934 4135 1940 4136
rect 1936 4075 1938 4135
rect 1976 4111 1978 4171
rect 1996 4111 1998 4172
rect 2124 4128 2126 4186
rect 2162 4177 2168 4178
rect 2162 4173 2163 4177
rect 2167 4173 2168 4177
rect 2162 4172 2168 4173
rect 2122 4127 2128 4128
rect 2122 4123 2123 4127
rect 2127 4123 2128 4127
rect 2122 4122 2128 4123
rect 2164 4111 2166 4172
rect 1975 4110 1979 4111
rect 1975 4105 1979 4106
rect 1995 4110 1999 4111
rect 1995 4105 1999 4106
rect 2075 4110 2079 4111
rect 2075 4105 2079 4106
rect 2163 4110 2167 4111
rect 2163 4105 2167 4106
rect 2259 4110 2263 4111
rect 2259 4105 2263 4106
rect 1755 4074 1759 4075
rect 1755 4069 1759 4070
rect 1787 4074 1791 4075
rect 1787 4069 1791 4070
rect 1935 4074 1939 4075
rect 1935 4069 1939 4070
rect 1788 4008 1790 4069
rect 1906 4059 1912 4060
rect 1906 4055 1907 4059
rect 1911 4055 1912 4059
rect 1906 4054 1912 4055
rect 1786 4007 1792 4008
rect 1786 4003 1787 4007
rect 1791 4003 1792 4007
rect 1786 4002 1792 4003
rect 1814 3992 1820 3993
rect 1518 3988 1519 3992
rect 1523 3988 1524 3992
rect 1518 3987 1524 3988
rect 1614 3991 1620 3992
rect 1614 3987 1615 3991
rect 1619 3987 1620 3991
rect 1814 3988 1815 3992
rect 1819 3988 1820 3992
rect 1814 3987 1820 3988
rect 110 3986 116 3987
rect 112 3959 114 3986
rect 160 3959 162 3987
rect 254 3986 260 3987
rect 111 3958 115 3959
rect 111 3953 115 3954
rect 159 3958 163 3959
rect 159 3953 163 3954
rect 112 3930 114 3953
rect 110 3929 116 3930
rect 160 3929 162 3953
rect 110 3925 111 3929
rect 115 3925 116 3929
rect 110 3924 116 3925
rect 158 3928 164 3929
rect 158 3924 159 3928
rect 163 3924 164 3928
rect 158 3923 164 3924
rect 130 3913 136 3914
rect 110 3912 116 3913
rect 110 3908 111 3912
rect 115 3908 116 3912
rect 130 3909 131 3913
rect 135 3909 136 3913
rect 130 3908 136 3909
rect 110 3907 116 3908
rect 112 3839 114 3907
rect 132 3839 134 3908
rect 256 3864 258 3986
rect 368 3959 370 3987
rect 462 3986 468 3987
rect 624 3959 626 3987
rect 904 3959 906 3987
rect 1186 3986 1192 3987
rect 1208 3959 1210 3987
rect 1520 3959 1522 3987
rect 1614 3986 1620 3987
rect 1816 3959 1818 3987
rect 343 3958 347 3959
rect 343 3953 347 3954
rect 367 3958 371 3959
rect 367 3953 371 3954
rect 567 3958 571 3959
rect 567 3953 571 3954
rect 623 3958 627 3959
rect 623 3953 627 3954
rect 807 3958 811 3959
rect 807 3953 811 3954
rect 903 3958 907 3959
rect 903 3953 907 3954
rect 1055 3958 1059 3959
rect 1055 3953 1059 3954
rect 1207 3958 1211 3959
rect 1207 3953 1211 3954
rect 1311 3958 1315 3959
rect 1311 3953 1315 3954
rect 1519 3958 1523 3959
rect 1519 3953 1523 3954
rect 1575 3958 1579 3959
rect 1575 3953 1579 3954
rect 1815 3958 1819 3959
rect 1815 3953 1819 3954
rect 344 3929 346 3953
rect 362 3943 368 3944
rect 362 3939 363 3943
rect 367 3939 368 3943
rect 362 3938 368 3939
rect 342 3928 348 3929
rect 274 3927 280 3928
rect 274 3923 275 3927
rect 279 3923 280 3927
rect 342 3924 343 3928
rect 347 3924 348 3928
rect 342 3923 348 3924
rect 274 3922 280 3923
rect 276 3864 278 3922
rect 314 3913 320 3914
rect 314 3909 315 3913
rect 319 3909 320 3913
rect 314 3908 320 3909
rect 254 3863 260 3864
rect 254 3859 255 3863
rect 259 3859 260 3863
rect 254 3858 260 3859
rect 274 3863 280 3864
rect 274 3859 275 3863
rect 279 3859 280 3863
rect 274 3858 280 3859
rect 316 3839 318 3908
rect 111 3838 115 3839
rect 111 3833 115 3834
rect 131 3838 135 3839
rect 131 3833 135 3834
rect 267 3838 271 3839
rect 267 3833 271 3834
rect 315 3838 319 3839
rect 315 3833 319 3834
rect 112 3773 114 3833
rect 110 3772 116 3773
rect 268 3772 270 3833
rect 364 3824 366 3938
rect 568 3929 570 3953
rect 808 3929 810 3953
rect 1056 3929 1058 3953
rect 1312 3929 1314 3953
rect 1576 3929 1578 3953
rect 1816 3929 1818 3953
rect 566 3928 572 3929
rect 806 3928 812 3929
rect 1054 3928 1060 3929
rect 438 3927 444 3928
rect 438 3923 439 3927
rect 443 3923 444 3927
rect 566 3924 567 3928
rect 571 3924 572 3928
rect 566 3923 572 3924
rect 694 3927 700 3928
rect 694 3923 695 3927
rect 699 3923 700 3927
rect 806 3924 807 3928
rect 811 3924 812 3928
rect 806 3923 812 3924
rect 942 3927 948 3928
rect 942 3923 943 3927
rect 947 3923 948 3927
rect 1054 3924 1055 3928
rect 1059 3924 1060 3928
rect 1054 3923 1060 3924
rect 1310 3928 1316 3929
rect 1310 3924 1311 3928
rect 1315 3924 1316 3928
rect 1310 3923 1316 3924
rect 1574 3928 1580 3929
rect 1574 3924 1575 3928
rect 1579 3924 1580 3928
rect 1574 3923 1580 3924
rect 1814 3928 1820 3929
rect 1908 3928 1910 4054
rect 1914 4035 1920 4036
rect 1914 4031 1915 4035
rect 1919 4031 1920 4035
rect 1914 4030 1920 4031
rect 1916 3992 1918 4030
rect 1936 4009 1938 4069
rect 1976 4045 1978 4105
rect 1974 4044 1980 4045
rect 2076 4044 2078 4105
rect 2260 4044 2262 4105
rect 2288 4096 2290 4186
rect 2354 4177 2360 4178
rect 2354 4173 2355 4177
rect 2359 4173 2360 4177
rect 2354 4172 2360 4173
rect 2356 4111 2358 4172
rect 2480 4120 2482 4186
rect 2504 4128 2506 4274
rect 2832 4223 2834 4275
rect 2926 4274 2932 4275
rect 2583 4222 2587 4223
rect 2583 4217 2587 4218
rect 2783 4222 2787 4223
rect 2783 4217 2787 4218
rect 2831 4222 2835 4223
rect 2831 4217 2835 4218
rect 2983 4222 2987 4223
rect 2983 4217 2987 4218
rect 2584 4193 2586 4217
rect 2784 4193 2786 4217
rect 2984 4193 2986 4217
rect 2582 4192 2588 4193
rect 2782 4192 2788 4193
rect 2982 4192 2988 4193
rect 3244 4192 3246 4338
rect 3262 4280 3268 4281
rect 3360 4280 3362 4346
rect 3652 4296 3654 4357
rect 3772 4348 3774 4450
rect 3798 4440 3804 4441
rect 3798 4436 3799 4440
rect 3803 4436 3804 4440
rect 3798 4435 3804 4436
rect 3800 4363 3802 4435
rect 3840 4375 3842 4459
rect 4460 4375 4462 4460
rect 4550 4415 4556 4416
rect 4550 4411 4551 4415
rect 4555 4411 4556 4415
rect 4550 4410 4556 4411
rect 3839 4374 3843 4375
rect 3839 4369 3843 4370
rect 3859 4374 3863 4375
rect 3859 4369 3863 4370
rect 3995 4374 3999 4375
rect 3995 4369 3999 4370
rect 4131 4374 4135 4375
rect 4131 4369 4135 4370
rect 4283 4374 4287 4375
rect 4283 4369 4287 4370
rect 4459 4374 4463 4375
rect 4459 4369 4463 4370
rect 4483 4374 4487 4375
rect 4483 4369 4487 4370
rect 3799 4362 3803 4363
rect 3778 4359 3784 4360
rect 3778 4355 3779 4359
rect 3783 4355 3784 4359
rect 3799 4357 3803 4358
rect 3778 4354 3784 4355
rect 3770 4347 3776 4348
rect 3770 4343 3771 4347
rect 3775 4343 3776 4347
rect 3770 4342 3776 4343
rect 3650 4295 3656 4296
rect 3650 4291 3651 4295
rect 3655 4291 3656 4295
rect 3650 4290 3656 4291
rect 3678 4280 3684 4281
rect 3780 4280 3782 4354
rect 3800 4297 3802 4357
rect 3840 4309 3842 4369
rect 3838 4308 3844 4309
rect 3860 4308 3862 4369
rect 3996 4308 3998 4369
rect 4002 4355 4008 4356
rect 4002 4351 4003 4355
rect 4007 4351 4008 4355
rect 4002 4350 4008 4351
rect 3838 4304 3839 4308
rect 3843 4304 3844 4308
rect 3838 4303 3844 4304
rect 3858 4307 3864 4308
rect 3858 4303 3859 4307
rect 3863 4303 3864 4307
rect 3858 4302 3864 4303
rect 3994 4307 4000 4308
rect 3994 4303 3995 4307
rect 3999 4303 4000 4307
rect 3994 4302 4000 4303
rect 3798 4296 3804 4297
rect 3798 4292 3799 4296
rect 3803 4292 3804 4296
rect 3886 4292 3892 4293
rect 4004 4292 4006 4350
rect 4132 4308 4134 4369
rect 4138 4355 4144 4356
rect 4138 4351 4139 4355
rect 4143 4351 4144 4355
rect 4138 4350 4144 4351
rect 4130 4307 4136 4308
rect 4130 4303 4131 4307
rect 4135 4303 4136 4307
rect 4130 4302 4136 4303
rect 4022 4292 4028 4293
rect 4140 4292 4142 4350
rect 4284 4308 4286 4369
rect 4378 4355 4384 4356
rect 4378 4351 4379 4355
rect 4383 4351 4384 4355
rect 4378 4350 4384 4351
rect 4282 4307 4288 4308
rect 4282 4303 4283 4307
rect 4287 4303 4288 4307
rect 4282 4302 4288 4303
rect 4158 4292 4164 4293
rect 4310 4292 4316 4293
rect 3798 4291 3804 4292
rect 3838 4291 3844 4292
rect 3838 4287 3839 4291
rect 3843 4287 3844 4291
rect 3886 4288 3887 4292
rect 3891 4288 3892 4292
rect 3886 4287 3892 4288
rect 4002 4291 4008 4292
rect 4002 4287 4003 4291
rect 4007 4287 4008 4291
rect 4022 4288 4023 4292
rect 4027 4288 4028 4292
rect 4022 4287 4028 4288
rect 4138 4291 4144 4292
rect 4138 4287 4139 4291
rect 4143 4287 4144 4291
rect 4158 4288 4159 4292
rect 4163 4288 4164 4292
rect 4158 4287 4164 4288
rect 4254 4291 4260 4292
rect 4254 4287 4255 4291
rect 4259 4287 4260 4291
rect 4310 4288 4311 4292
rect 4315 4288 4316 4292
rect 4310 4287 4316 4288
rect 3838 4286 3844 4287
rect 3262 4276 3263 4280
rect 3267 4276 3268 4280
rect 3262 4275 3268 4276
rect 3358 4279 3364 4280
rect 3358 4275 3359 4279
rect 3363 4275 3364 4279
rect 3678 4276 3679 4280
rect 3683 4276 3684 4280
rect 3678 4275 3684 4276
rect 3778 4279 3784 4280
rect 3778 4275 3779 4279
rect 3783 4275 3784 4279
rect 3264 4223 3266 4275
rect 3358 4274 3364 4275
rect 3680 4223 3682 4275
rect 3778 4274 3784 4275
rect 3798 4279 3804 4280
rect 3798 4275 3799 4279
rect 3803 4275 3804 4279
rect 3798 4274 3804 4275
rect 3800 4223 3802 4274
rect 3840 4263 3842 4286
rect 3888 4263 3890 4287
rect 4002 4286 4008 4287
rect 4024 4263 4026 4287
rect 4138 4286 4144 4287
rect 4160 4263 4162 4287
rect 4254 4286 4260 4287
rect 3839 4262 3843 4263
rect 3839 4257 3843 4258
rect 3887 4262 3891 4263
rect 3887 4257 3891 4258
rect 4023 4262 4027 4263
rect 4023 4257 4027 4258
rect 4159 4262 4163 4263
rect 4159 4257 4163 4258
rect 3840 4234 3842 4257
rect 3838 4233 3844 4234
rect 3888 4233 3890 4257
rect 4024 4233 4026 4257
rect 4160 4233 4162 4257
rect 3838 4229 3839 4233
rect 3843 4229 3844 4233
rect 3838 4228 3844 4229
rect 3886 4232 3892 4233
rect 4022 4232 4028 4233
rect 4158 4232 4164 4233
rect 3886 4228 3887 4232
rect 3891 4228 3892 4232
rect 3886 4227 3892 4228
rect 3986 4231 3992 4232
rect 3986 4227 3987 4231
rect 3991 4227 3992 4231
rect 4022 4228 4023 4232
rect 4027 4228 4028 4232
rect 4022 4227 4028 4228
rect 4122 4231 4128 4232
rect 4122 4227 4123 4231
rect 4127 4227 4128 4231
rect 4158 4228 4159 4232
rect 4163 4228 4164 4232
rect 4158 4227 4164 4228
rect 3986 4226 3992 4227
rect 4122 4226 4128 4227
rect 3263 4222 3267 4223
rect 3263 4217 3267 4218
rect 3679 4222 3683 4223
rect 3679 4217 3683 4218
rect 3799 4222 3803 4223
rect 3799 4217 3803 4218
rect 3858 4217 3864 4218
rect 3800 4194 3802 4217
rect 3838 4216 3844 4217
rect 3838 4212 3839 4216
rect 3843 4212 3844 4216
rect 3858 4213 3859 4217
rect 3863 4213 3864 4217
rect 3858 4212 3864 4213
rect 3838 4211 3844 4212
rect 3798 4193 3804 4194
rect 2582 4188 2583 4192
rect 2587 4188 2588 4192
rect 2582 4187 2588 4188
rect 2682 4191 2688 4192
rect 2682 4187 2683 4191
rect 2687 4187 2688 4191
rect 2782 4188 2783 4192
rect 2787 4188 2788 4192
rect 2782 4187 2788 4188
rect 2882 4191 2888 4192
rect 2882 4187 2883 4191
rect 2887 4187 2888 4191
rect 2982 4188 2983 4192
rect 2987 4188 2988 4192
rect 2982 4187 2988 4188
rect 3242 4191 3248 4192
rect 3242 4187 3243 4191
rect 3247 4187 3248 4191
rect 3798 4189 3799 4193
rect 3803 4189 3804 4193
rect 3798 4188 3804 4189
rect 2682 4186 2688 4187
rect 2882 4186 2888 4187
rect 3242 4186 3248 4187
rect 2554 4177 2560 4178
rect 2554 4173 2555 4177
rect 2559 4173 2560 4177
rect 2554 4172 2560 4173
rect 2502 4127 2508 4128
rect 2502 4123 2503 4127
rect 2507 4123 2508 4127
rect 2502 4122 2508 4123
rect 2478 4119 2484 4120
rect 2478 4115 2479 4119
rect 2483 4115 2484 4119
rect 2478 4114 2484 4115
rect 2556 4111 2558 4172
rect 2684 4128 2686 4186
rect 2754 4177 2760 4178
rect 2754 4173 2755 4177
rect 2759 4173 2760 4177
rect 2754 4172 2760 4173
rect 2566 4127 2572 4128
rect 2566 4123 2567 4127
rect 2571 4123 2572 4127
rect 2566 4122 2572 4123
rect 2682 4127 2688 4128
rect 2682 4123 2683 4127
rect 2687 4123 2688 4127
rect 2682 4122 2688 4123
rect 2355 4110 2359 4111
rect 2355 4105 2359 4106
rect 2443 4110 2447 4111
rect 2443 4105 2447 4106
rect 2555 4110 2559 4111
rect 2555 4105 2559 4106
rect 2286 4095 2292 4096
rect 2286 4091 2287 4095
rect 2291 4091 2292 4095
rect 2286 4090 2292 4091
rect 2444 4044 2446 4105
rect 2538 4091 2544 4092
rect 2538 4087 2539 4091
rect 2543 4087 2544 4091
rect 2538 4086 2544 4087
rect 2540 4064 2542 4086
rect 2538 4063 2544 4064
rect 2538 4059 2539 4063
rect 2543 4059 2544 4063
rect 2538 4058 2544 4059
rect 1974 4040 1975 4044
rect 1979 4040 1980 4044
rect 1974 4039 1980 4040
rect 2074 4043 2080 4044
rect 2074 4039 2075 4043
rect 2079 4039 2080 4043
rect 2074 4038 2080 4039
rect 2258 4043 2264 4044
rect 2258 4039 2259 4043
rect 2263 4039 2264 4043
rect 2258 4038 2264 4039
rect 2442 4043 2448 4044
rect 2442 4039 2443 4043
rect 2447 4039 2448 4043
rect 2442 4038 2448 4039
rect 2102 4028 2108 4029
rect 2286 4028 2292 4029
rect 1974 4027 1980 4028
rect 1974 4023 1975 4027
rect 1979 4023 1980 4027
rect 2102 4024 2103 4028
rect 2107 4024 2108 4028
rect 2102 4023 2108 4024
rect 2194 4027 2200 4028
rect 2194 4023 2195 4027
rect 2199 4023 2200 4027
rect 2286 4024 2287 4028
rect 2291 4024 2292 4028
rect 2286 4023 2292 4024
rect 2470 4028 2476 4029
rect 2568 4028 2570 4122
rect 2756 4111 2758 4172
rect 2884 4128 2886 4186
rect 2954 4177 2960 4178
rect 2954 4173 2955 4177
rect 2959 4173 2960 4177
rect 2954 4172 2960 4173
rect 3798 4176 3804 4177
rect 3798 4172 3799 4176
rect 3803 4172 3804 4176
rect 2882 4127 2888 4128
rect 2882 4123 2883 4127
rect 2887 4123 2888 4127
rect 2882 4122 2888 4123
rect 2956 4111 2958 4172
rect 3798 4171 3804 4172
rect 3800 4111 3802 4171
rect 3840 4111 3842 4211
rect 3860 4111 3862 4212
rect 3988 4168 3990 4226
rect 3994 4217 4000 4218
rect 3994 4213 3995 4217
rect 3999 4213 4000 4217
rect 3994 4212 4000 4213
rect 3986 4167 3992 4168
rect 3986 4163 3987 4167
rect 3991 4163 3992 4167
rect 3986 4162 3992 4163
rect 3996 4111 3998 4212
rect 4124 4168 4126 4226
rect 4130 4217 4136 4218
rect 4130 4213 4131 4217
rect 4135 4213 4136 4217
rect 4130 4212 4136 4213
rect 4122 4167 4128 4168
rect 4122 4163 4123 4167
rect 4127 4163 4128 4167
rect 4122 4162 4128 4163
rect 4132 4111 4134 4212
rect 4256 4160 4258 4286
rect 4312 4263 4314 4287
rect 4380 4277 4382 4350
rect 4484 4308 4486 4369
rect 4490 4355 4496 4356
rect 4490 4351 4491 4355
rect 4495 4351 4496 4355
rect 4490 4350 4496 4351
rect 4482 4307 4488 4308
rect 4482 4303 4483 4307
rect 4487 4303 4488 4307
rect 4482 4302 4488 4303
rect 4492 4292 4494 4350
rect 4510 4292 4516 4293
rect 4490 4291 4496 4292
rect 4490 4287 4491 4291
rect 4495 4287 4496 4291
rect 4510 4288 4511 4292
rect 4515 4288 4516 4292
rect 4510 4287 4516 4288
rect 4490 4286 4496 4287
rect 4379 4276 4383 4277
rect 4379 4271 4383 4272
rect 4512 4263 4514 4287
rect 4552 4280 4554 4410
rect 4644 4375 4646 4460
rect 4852 4375 4854 4460
rect 4980 4416 4982 4474
rect 5066 4465 5072 4466
rect 5066 4461 5067 4465
rect 5071 4461 5072 4465
rect 5066 4460 5072 4461
rect 5298 4465 5304 4466
rect 5298 4461 5299 4465
rect 5303 4461 5304 4465
rect 5298 4460 5304 4461
rect 5514 4465 5520 4466
rect 5514 4461 5515 4465
rect 5519 4461 5520 4465
rect 5514 4460 5520 4461
rect 4978 4415 4984 4416
rect 4978 4411 4979 4415
rect 4983 4411 4984 4415
rect 4978 4410 4984 4411
rect 5068 4375 5070 4460
rect 5300 4375 5302 4460
rect 5516 4375 5518 4460
rect 4643 4374 4647 4375
rect 4643 4369 4647 4370
rect 4715 4374 4719 4375
rect 4715 4369 4719 4370
rect 4851 4374 4855 4375
rect 4851 4369 4855 4370
rect 4979 4374 4983 4375
rect 4979 4369 4983 4370
rect 5067 4374 5071 4375
rect 5067 4369 5071 4370
rect 5251 4374 5255 4375
rect 5251 4369 5255 4370
rect 5299 4374 5303 4375
rect 5299 4369 5303 4370
rect 5515 4374 5519 4375
rect 5515 4369 5519 4370
rect 4716 4308 4718 4369
rect 4722 4355 4728 4356
rect 4722 4351 4723 4355
rect 4727 4351 4728 4355
rect 4722 4350 4728 4351
rect 4714 4307 4720 4308
rect 4714 4303 4715 4307
rect 4719 4303 4720 4307
rect 4714 4302 4720 4303
rect 4724 4292 4726 4350
rect 4980 4308 4982 4369
rect 4986 4355 4992 4356
rect 4986 4351 4987 4355
rect 4991 4351 4992 4355
rect 4986 4350 4992 4351
rect 4978 4307 4984 4308
rect 4978 4303 4979 4307
rect 4983 4303 4984 4307
rect 4978 4302 4984 4303
rect 4742 4292 4748 4293
rect 4988 4292 4990 4350
rect 5252 4308 5254 4369
rect 5258 4355 5264 4356
rect 5258 4351 5259 4355
rect 5263 4351 5264 4355
rect 5258 4350 5264 4351
rect 5250 4307 5256 4308
rect 5250 4303 5251 4307
rect 5255 4303 5256 4307
rect 5250 4302 5256 4303
rect 5006 4292 5012 4293
rect 5260 4292 5262 4350
rect 5516 4308 5518 4369
rect 5636 4360 5638 4474
rect 5644 4416 5646 4546
rect 5664 4511 5666 4546
rect 5663 4510 5667 4511
rect 5663 4505 5667 4506
rect 5664 4482 5666 4505
rect 5662 4481 5668 4482
rect 5662 4477 5663 4481
rect 5667 4477 5668 4481
rect 5662 4476 5668 4477
rect 5662 4464 5668 4465
rect 5662 4460 5663 4464
rect 5667 4460 5668 4464
rect 5662 4459 5668 4460
rect 5642 4415 5648 4416
rect 5642 4411 5643 4415
rect 5647 4411 5648 4415
rect 5642 4410 5648 4411
rect 5664 4375 5666 4459
rect 5663 4374 5667 4375
rect 5663 4369 5667 4370
rect 5634 4359 5640 4360
rect 5634 4355 5635 4359
rect 5639 4355 5640 4359
rect 5634 4354 5640 4355
rect 5664 4309 5666 4369
rect 5662 4308 5668 4309
rect 5514 4307 5520 4308
rect 5514 4303 5515 4307
rect 5519 4303 5520 4307
rect 5662 4304 5663 4308
rect 5667 4304 5668 4308
rect 5662 4303 5668 4304
rect 5514 4302 5520 4303
rect 5278 4292 5284 4293
rect 4722 4291 4728 4292
rect 4722 4287 4723 4291
rect 4727 4287 4728 4291
rect 4742 4288 4743 4292
rect 4747 4288 4748 4292
rect 4742 4287 4748 4288
rect 4986 4291 4992 4292
rect 4986 4287 4987 4291
rect 4991 4287 4992 4291
rect 5006 4288 5007 4292
rect 5011 4288 5012 4292
rect 5006 4287 5012 4288
rect 5258 4291 5264 4292
rect 5258 4287 5259 4291
rect 5263 4287 5264 4291
rect 5278 4288 5279 4292
rect 5283 4288 5284 4292
rect 5278 4287 5284 4288
rect 5542 4292 5548 4293
rect 5542 4288 5543 4292
rect 5547 4288 5548 4292
rect 5542 4287 5548 4288
rect 5638 4291 5644 4292
rect 5638 4287 5639 4291
rect 5643 4287 5644 4291
rect 4722 4286 4728 4287
rect 4550 4279 4556 4280
rect 4550 4275 4551 4279
rect 4555 4275 4556 4279
rect 4550 4274 4556 4275
rect 4744 4263 4746 4287
rect 4986 4286 4992 4287
rect 5008 4263 5010 4287
rect 5258 4286 5264 4287
rect 5280 4263 5282 4287
rect 5367 4276 5371 4277
rect 5367 4271 5371 4272
rect 4303 4262 4307 4263
rect 4303 4257 4307 4258
rect 4311 4262 4315 4263
rect 4311 4257 4315 4258
rect 4503 4262 4507 4263
rect 4503 4257 4507 4258
rect 4511 4262 4515 4263
rect 4511 4257 4515 4258
rect 4735 4262 4739 4263
rect 4735 4257 4739 4258
rect 4743 4262 4747 4263
rect 4743 4257 4747 4258
rect 4999 4262 5003 4263
rect 4999 4257 5003 4258
rect 5007 4262 5011 4263
rect 5007 4257 5011 4258
rect 5271 4262 5275 4263
rect 5271 4257 5275 4258
rect 5279 4262 5283 4263
rect 5279 4257 5283 4258
rect 4304 4233 4306 4257
rect 4504 4233 4506 4257
rect 4736 4233 4738 4257
rect 5000 4233 5002 4257
rect 5272 4233 5274 4257
rect 4302 4232 4308 4233
rect 4502 4232 4508 4233
rect 4302 4228 4303 4232
rect 4307 4228 4308 4232
rect 4302 4227 4308 4228
rect 4446 4231 4452 4232
rect 4446 4227 4447 4231
rect 4451 4227 4452 4231
rect 4502 4228 4503 4232
rect 4507 4228 4508 4232
rect 4502 4227 4508 4228
rect 4734 4232 4740 4233
rect 4734 4228 4735 4232
rect 4739 4228 4740 4232
rect 4734 4227 4740 4228
rect 4998 4232 5004 4233
rect 5270 4232 5276 4233
rect 5368 4232 5370 4271
rect 5544 4263 5546 4287
rect 5638 4286 5644 4287
rect 5662 4291 5668 4292
rect 5662 4287 5663 4291
rect 5667 4287 5668 4291
rect 5662 4286 5668 4287
rect 5543 4262 5547 4263
rect 5543 4257 5547 4258
rect 5544 4233 5546 4257
rect 5542 4232 5548 4233
rect 4998 4228 4999 4232
rect 5003 4228 5004 4232
rect 4998 4227 5004 4228
rect 5098 4231 5104 4232
rect 5098 4227 5099 4231
rect 5103 4227 5104 4231
rect 5270 4228 5271 4232
rect 5275 4228 5276 4232
rect 5270 4227 5276 4228
rect 5366 4231 5372 4232
rect 5366 4227 5367 4231
rect 5371 4227 5372 4231
rect 5542 4228 5543 4232
rect 5547 4228 5548 4232
rect 5542 4227 5548 4228
rect 4446 4226 4452 4227
rect 5098 4226 5104 4227
rect 5366 4226 5372 4227
rect 4274 4217 4280 4218
rect 4274 4213 4275 4217
rect 4279 4213 4280 4217
rect 4274 4212 4280 4213
rect 4254 4159 4260 4160
rect 4254 4155 4255 4159
rect 4259 4155 4260 4159
rect 4254 4154 4260 4155
rect 4276 4111 4278 4212
rect 4448 4168 4450 4226
rect 4474 4217 4480 4218
rect 4474 4213 4475 4217
rect 4479 4213 4480 4217
rect 4474 4212 4480 4213
rect 4706 4217 4712 4218
rect 4706 4213 4707 4217
rect 4711 4213 4712 4217
rect 4706 4212 4712 4213
rect 4970 4217 4976 4218
rect 4970 4213 4971 4217
rect 4975 4213 4976 4217
rect 4970 4212 4976 4213
rect 4446 4167 4452 4168
rect 4446 4163 4447 4167
rect 4451 4163 4452 4167
rect 4446 4162 4452 4163
rect 4476 4111 4478 4212
rect 4708 4111 4710 4212
rect 4972 4111 4974 4212
rect 5100 4168 5102 4226
rect 5242 4217 5248 4218
rect 5242 4213 5243 4217
rect 5247 4213 5248 4217
rect 5242 4212 5248 4213
rect 5514 4217 5520 4218
rect 5514 4213 5515 4217
rect 5519 4213 5520 4217
rect 5514 4212 5520 4213
rect 5098 4167 5104 4168
rect 5098 4163 5099 4167
rect 5103 4163 5104 4167
rect 5098 4162 5104 4163
rect 5244 4111 5246 4212
rect 5516 4111 5518 4212
rect 5640 4168 5642 4286
rect 5664 4263 5666 4286
rect 5663 4262 5667 4263
rect 5663 4257 5667 4258
rect 5664 4234 5666 4257
rect 5662 4233 5668 4234
rect 5662 4229 5663 4233
rect 5667 4229 5668 4233
rect 5662 4228 5668 4229
rect 5662 4216 5668 4217
rect 5662 4212 5663 4216
rect 5667 4212 5668 4216
rect 5662 4211 5668 4212
rect 5638 4167 5644 4168
rect 5638 4163 5639 4167
rect 5643 4163 5644 4167
rect 5638 4162 5644 4163
rect 5664 4111 5666 4211
rect 2619 4110 2623 4111
rect 2619 4105 2623 4106
rect 2755 4110 2759 4111
rect 2755 4105 2759 4106
rect 2787 4110 2791 4111
rect 2787 4105 2791 4106
rect 2955 4110 2959 4111
rect 2955 4105 2959 4106
rect 3131 4110 3135 4111
rect 3131 4105 3135 4106
rect 3799 4110 3803 4111
rect 3799 4105 3803 4106
rect 3839 4110 3843 4111
rect 3839 4105 3843 4106
rect 3859 4110 3863 4111
rect 3859 4105 3863 4106
rect 3995 4110 3999 4111
rect 3995 4105 3999 4106
rect 4131 4110 4135 4111
rect 4131 4105 4135 4106
rect 4275 4110 4279 4111
rect 4275 4105 4279 4106
rect 4475 4110 4479 4111
rect 4475 4105 4479 4106
rect 4563 4110 4567 4111
rect 4563 4105 4567 4106
rect 4699 4110 4703 4111
rect 4699 4105 4703 4106
rect 4707 4110 4711 4111
rect 4707 4105 4711 4106
rect 4835 4110 4839 4111
rect 4835 4105 4839 4106
rect 4971 4110 4975 4111
rect 4971 4105 4975 4106
rect 5107 4110 5111 4111
rect 5107 4105 5111 4106
rect 5243 4110 5247 4111
rect 5243 4105 5247 4106
rect 5379 4110 5383 4111
rect 5379 4105 5383 4106
rect 5515 4110 5519 4111
rect 5515 4105 5519 4106
rect 5663 4110 5667 4111
rect 5663 4105 5667 4106
rect 2620 4044 2622 4105
rect 2746 4095 2752 4096
rect 2746 4091 2747 4095
rect 2751 4091 2752 4095
rect 2746 4090 2752 4091
rect 2738 4063 2744 4064
rect 2738 4059 2739 4063
rect 2743 4059 2744 4063
rect 2738 4058 2744 4059
rect 2618 4043 2624 4044
rect 2618 4039 2619 4043
rect 2623 4039 2624 4043
rect 2618 4038 2624 4039
rect 2646 4028 2652 4029
rect 2470 4024 2471 4028
rect 2475 4024 2476 4028
rect 2470 4023 2476 4024
rect 2566 4027 2572 4028
rect 2566 4023 2567 4027
rect 2571 4023 2572 4027
rect 2646 4024 2647 4028
rect 2651 4024 2652 4028
rect 2740 4028 2742 4058
rect 2748 4036 2750 4090
rect 2788 4044 2790 4105
rect 2956 4044 2958 4105
rect 3078 4099 3084 4100
rect 3078 4095 3079 4099
rect 3083 4095 3084 4099
rect 3078 4094 3084 4095
rect 2786 4043 2792 4044
rect 2786 4039 2787 4043
rect 2791 4039 2792 4043
rect 2786 4038 2792 4039
rect 2954 4043 2960 4044
rect 2954 4039 2955 4043
rect 2959 4039 2960 4043
rect 2954 4038 2960 4039
rect 2746 4035 2752 4036
rect 2746 4031 2747 4035
rect 2751 4031 2752 4035
rect 2746 4030 2752 4031
rect 2814 4028 2820 4029
rect 2740 4027 2748 4028
rect 2740 4025 2743 4027
rect 2646 4023 2652 4024
rect 2742 4023 2743 4025
rect 2747 4023 2748 4027
rect 2814 4024 2815 4028
rect 2819 4024 2820 4028
rect 2814 4023 2820 4024
rect 2982 4028 2988 4029
rect 3080 4028 3082 4094
rect 3132 4044 3134 4105
rect 3138 4091 3144 4092
rect 3138 4087 3139 4091
rect 3143 4087 3144 4091
rect 3138 4086 3144 4087
rect 3130 4043 3136 4044
rect 3130 4039 3131 4043
rect 3135 4039 3136 4043
rect 3130 4038 3136 4039
rect 2982 4024 2983 4028
rect 2987 4024 2988 4028
rect 2982 4023 2988 4024
rect 3078 4027 3084 4028
rect 3078 4023 3079 4027
rect 3083 4023 3084 4027
rect 1974 4022 1980 4023
rect 1934 4008 1940 4009
rect 1934 4004 1935 4008
rect 1939 4004 1940 4008
rect 1934 4003 1940 4004
rect 1914 3991 1920 3992
rect 1914 3987 1915 3991
rect 1919 3987 1920 3991
rect 1914 3986 1920 3987
rect 1934 3991 1940 3992
rect 1976 3991 1978 4022
rect 2104 3991 2106 4023
rect 2194 4022 2200 4023
rect 1934 3987 1935 3991
rect 1939 3987 1940 3991
rect 1934 3986 1940 3987
rect 1975 3990 1979 3991
rect 1936 3959 1938 3986
rect 1975 3985 1979 3986
rect 2103 3990 2107 3991
rect 2103 3985 2107 3986
rect 2127 3990 2131 3991
rect 2127 3985 2131 3986
rect 1976 3962 1978 3985
rect 1974 3961 1980 3962
rect 2128 3961 2130 3985
rect 1935 3958 1939 3959
rect 1974 3957 1975 3961
rect 1979 3957 1980 3961
rect 1974 3956 1980 3957
rect 2126 3960 2132 3961
rect 2126 3956 2127 3960
rect 2131 3956 2132 3960
rect 2126 3955 2132 3956
rect 1935 3953 1939 3954
rect 1936 3930 1938 3953
rect 2098 3945 2104 3946
rect 1974 3944 1980 3945
rect 1974 3940 1975 3944
rect 1979 3940 1980 3944
rect 2098 3941 2099 3945
rect 2103 3941 2104 3945
rect 2098 3940 2104 3941
rect 1974 3939 1980 3940
rect 1934 3929 1940 3930
rect 1814 3924 1815 3928
rect 1819 3924 1820 3928
rect 1814 3923 1820 3924
rect 1906 3927 1912 3928
rect 1906 3923 1907 3927
rect 1911 3923 1912 3927
rect 1934 3925 1935 3929
rect 1939 3925 1940 3929
rect 1934 3924 1940 3925
rect 438 3922 444 3923
rect 694 3922 700 3923
rect 942 3922 948 3923
rect 1906 3922 1912 3923
rect 440 3864 442 3922
rect 538 3913 544 3914
rect 538 3909 539 3913
rect 543 3909 544 3913
rect 538 3908 544 3909
rect 438 3863 444 3864
rect 438 3859 439 3863
rect 443 3859 444 3863
rect 438 3858 444 3859
rect 540 3839 542 3908
rect 696 3864 698 3922
rect 778 3913 784 3914
rect 778 3909 779 3913
rect 783 3909 784 3913
rect 778 3908 784 3909
rect 694 3863 700 3864
rect 694 3859 695 3863
rect 699 3859 700 3863
rect 694 3858 700 3859
rect 780 3839 782 3908
rect 944 3864 946 3922
rect 1026 3913 1032 3914
rect 1026 3909 1027 3913
rect 1031 3909 1032 3913
rect 1026 3908 1032 3909
rect 1282 3913 1288 3914
rect 1282 3909 1283 3913
rect 1287 3909 1288 3913
rect 1282 3908 1288 3909
rect 1546 3913 1552 3914
rect 1546 3909 1547 3913
rect 1551 3909 1552 3913
rect 1546 3908 1552 3909
rect 1786 3913 1792 3914
rect 1786 3909 1787 3913
rect 1791 3909 1792 3913
rect 1786 3908 1792 3909
rect 1934 3912 1940 3913
rect 1934 3908 1935 3912
rect 1939 3908 1940 3912
rect 942 3863 948 3864
rect 942 3859 943 3863
rect 947 3859 948 3863
rect 942 3858 948 3859
rect 1028 3839 1030 3908
rect 1284 3839 1286 3908
rect 1378 3863 1384 3864
rect 1378 3859 1379 3863
rect 1383 3859 1384 3863
rect 1378 3858 1384 3859
rect 475 3838 479 3839
rect 475 3833 479 3834
rect 539 3838 543 3839
rect 539 3833 543 3834
rect 707 3838 711 3839
rect 707 3833 711 3834
rect 779 3838 783 3839
rect 779 3833 783 3834
rect 963 3838 967 3839
rect 963 3833 967 3834
rect 1027 3838 1031 3839
rect 1027 3833 1031 3834
rect 1235 3838 1239 3839
rect 1235 3833 1239 3834
rect 1283 3838 1287 3839
rect 1283 3833 1287 3834
rect 362 3823 368 3824
rect 362 3819 363 3823
rect 367 3819 368 3823
rect 362 3818 368 3819
rect 476 3772 478 3833
rect 482 3819 488 3820
rect 482 3815 483 3819
rect 487 3815 488 3819
rect 482 3814 488 3815
rect 110 3768 111 3772
rect 115 3768 116 3772
rect 110 3767 116 3768
rect 266 3771 272 3772
rect 266 3767 267 3771
rect 271 3767 272 3771
rect 266 3766 272 3767
rect 474 3771 480 3772
rect 474 3767 475 3771
rect 479 3767 480 3771
rect 474 3766 480 3767
rect 294 3756 300 3757
rect 484 3756 486 3814
rect 708 3772 710 3833
rect 714 3819 720 3820
rect 714 3815 715 3819
rect 719 3815 720 3819
rect 714 3814 720 3815
rect 706 3771 712 3772
rect 706 3767 707 3771
rect 711 3767 712 3771
rect 706 3766 712 3767
rect 502 3756 508 3757
rect 716 3756 718 3814
rect 964 3772 966 3833
rect 970 3819 976 3820
rect 970 3815 971 3819
rect 975 3815 976 3819
rect 970 3814 976 3815
rect 962 3771 968 3772
rect 962 3767 963 3771
rect 967 3767 968 3771
rect 962 3766 968 3767
rect 734 3756 740 3757
rect 972 3756 974 3814
rect 1236 3772 1238 3833
rect 1242 3819 1248 3820
rect 1242 3815 1243 3819
rect 1247 3815 1248 3819
rect 1242 3814 1248 3815
rect 1234 3771 1240 3772
rect 1234 3767 1235 3771
rect 1239 3767 1240 3771
rect 1234 3766 1240 3767
rect 990 3756 996 3757
rect 1244 3756 1246 3814
rect 1380 3764 1382 3858
rect 1548 3839 1550 3908
rect 1788 3839 1790 3908
rect 1934 3907 1940 3908
rect 1936 3839 1938 3907
rect 1976 3871 1978 3939
rect 2100 3871 2102 3940
rect 2196 3896 2198 4022
rect 2288 3991 2290 4023
rect 2472 3991 2474 4023
rect 2566 4022 2572 4023
rect 2648 3991 2650 4023
rect 2742 4022 2748 4023
rect 2816 3991 2818 4023
rect 2984 3991 2986 4023
rect 3078 4022 3084 4023
rect 2287 3990 2291 3991
rect 2287 3985 2291 3986
rect 2311 3990 2315 3991
rect 2311 3985 2315 3986
rect 2471 3990 2475 3991
rect 2471 3985 2475 3986
rect 2487 3990 2491 3991
rect 2487 3985 2491 3986
rect 2647 3990 2651 3991
rect 2647 3985 2651 3986
rect 2663 3990 2667 3991
rect 2663 3985 2667 3986
rect 2815 3990 2819 3991
rect 2815 3985 2819 3986
rect 2831 3990 2835 3991
rect 2831 3985 2835 3986
rect 2983 3990 2987 3991
rect 2983 3985 2987 3986
rect 2999 3990 3003 3991
rect 2999 3985 3003 3986
rect 2312 3961 2314 3985
rect 2488 3961 2490 3985
rect 2664 3961 2666 3985
rect 2832 3961 2834 3985
rect 3000 3961 3002 3985
rect 2310 3960 2316 3961
rect 2310 3956 2311 3960
rect 2315 3956 2316 3960
rect 2310 3955 2316 3956
rect 2486 3960 2492 3961
rect 2662 3960 2668 3961
rect 2486 3956 2487 3960
rect 2491 3956 2492 3960
rect 2486 3955 2492 3956
rect 2578 3959 2584 3960
rect 2578 3955 2579 3959
rect 2583 3955 2584 3959
rect 2662 3956 2663 3960
rect 2667 3956 2668 3960
rect 2662 3955 2668 3956
rect 2830 3960 2836 3961
rect 2998 3960 3004 3961
rect 3140 3960 3142 4086
rect 3800 4045 3802 4105
rect 3840 4045 3842 4105
rect 3798 4044 3804 4045
rect 3798 4040 3799 4044
rect 3803 4040 3804 4044
rect 3798 4039 3804 4040
rect 3838 4044 3844 4045
rect 4564 4044 4566 4105
rect 4700 4044 4702 4105
rect 4706 4091 4712 4092
rect 4706 4087 4707 4091
rect 4711 4087 4712 4091
rect 4706 4086 4712 4087
rect 3838 4040 3839 4044
rect 3843 4040 3844 4044
rect 3838 4039 3844 4040
rect 4562 4043 4568 4044
rect 4562 4039 4563 4043
rect 4567 4039 4568 4043
rect 4562 4038 4568 4039
rect 4698 4043 4704 4044
rect 4698 4039 4699 4043
rect 4703 4039 4704 4043
rect 4698 4038 4704 4039
rect 3158 4028 3164 4029
rect 4590 4028 4596 4029
rect 4708 4028 4710 4086
rect 4836 4044 4838 4105
rect 4842 4091 4848 4092
rect 4842 4087 4843 4091
rect 4847 4087 4848 4091
rect 4842 4086 4848 4087
rect 4834 4043 4840 4044
rect 4834 4039 4835 4043
rect 4839 4039 4840 4043
rect 4834 4038 4840 4039
rect 4726 4028 4732 4029
rect 4844 4028 4846 4086
rect 4972 4044 4974 4105
rect 5090 4103 5096 4104
rect 5090 4099 5091 4103
rect 5095 4099 5096 4103
rect 5090 4098 5096 4099
rect 4970 4043 4976 4044
rect 4970 4039 4971 4043
rect 4975 4039 4976 4043
rect 4970 4038 4976 4039
rect 4862 4028 4868 4029
rect 4998 4028 5004 4029
rect 5092 4028 5094 4098
rect 5108 4044 5110 4105
rect 5230 4099 5236 4100
rect 5230 4095 5231 4099
rect 5235 4095 5236 4099
rect 5230 4094 5236 4095
rect 5202 4091 5208 4092
rect 5202 4087 5203 4091
rect 5207 4087 5208 4091
rect 5202 4086 5208 4087
rect 5204 4064 5206 4086
rect 5202 4063 5208 4064
rect 5202 4059 5203 4063
rect 5207 4059 5208 4063
rect 5202 4058 5208 4059
rect 5106 4043 5112 4044
rect 5106 4039 5107 4043
rect 5111 4039 5112 4043
rect 5106 4038 5112 4039
rect 5134 4028 5140 4029
rect 5232 4028 5234 4094
rect 5244 4044 5246 4105
rect 5338 4091 5344 4092
rect 5338 4087 5339 4091
rect 5343 4087 5344 4091
rect 5338 4086 5344 4087
rect 5340 4056 5342 4086
rect 5366 4063 5372 4064
rect 5366 4059 5367 4063
rect 5371 4059 5372 4063
rect 5366 4058 5372 4059
rect 5338 4055 5344 4056
rect 5338 4051 5339 4055
rect 5343 4051 5344 4055
rect 5338 4050 5344 4051
rect 5242 4043 5248 4044
rect 5242 4039 5243 4043
rect 5247 4039 5248 4043
rect 5242 4038 5248 4039
rect 5270 4028 5276 4029
rect 5368 4028 5370 4058
rect 5380 4044 5382 4105
rect 5422 4095 5428 4096
rect 5422 4091 5423 4095
rect 5427 4091 5428 4095
rect 5422 4090 5428 4091
rect 5378 4043 5384 4044
rect 5378 4039 5379 4043
rect 5383 4039 5384 4043
rect 5378 4038 5384 4039
rect 5406 4028 5412 4029
rect 3158 4024 3159 4028
rect 3163 4024 3164 4028
rect 3158 4023 3164 4024
rect 3798 4027 3804 4028
rect 3798 4023 3799 4027
rect 3803 4023 3804 4027
rect 3160 3991 3162 4023
rect 3798 4022 3804 4023
rect 3838 4027 3844 4028
rect 3838 4023 3839 4027
rect 3843 4023 3844 4027
rect 4590 4024 4591 4028
rect 4595 4024 4596 4028
rect 4590 4023 4596 4024
rect 4706 4027 4712 4028
rect 4706 4023 4707 4027
rect 4711 4023 4712 4027
rect 4726 4024 4727 4028
rect 4731 4024 4732 4028
rect 4726 4023 4732 4024
rect 4842 4027 4848 4028
rect 4842 4023 4843 4027
rect 4847 4023 4848 4027
rect 4862 4024 4863 4028
rect 4867 4024 4868 4028
rect 4862 4023 4868 4024
rect 4958 4027 4964 4028
rect 4958 4023 4959 4027
rect 4963 4023 4964 4027
rect 4998 4024 4999 4028
rect 5003 4024 5004 4028
rect 4998 4023 5004 4024
rect 5090 4027 5096 4028
rect 5090 4023 5091 4027
rect 5095 4023 5096 4027
rect 5134 4024 5135 4028
rect 5139 4024 5140 4028
rect 5134 4023 5140 4024
rect 5230 4027 5236 4028
rect 5230 4023 5231 4027
rect 5235 4023 5236 4027
rect 5270 4024 5271 4028
rect 5275 4024 5276 4028
rect 5270 4023 5276 4024
rect 5366 4027 5372 4028
rect 5366 4023 5367 4027
rect 5371 4023 5372 4027
rect 5406 4024 5407 4028
rect 5411 4024 5412 4028
rect 5406 4023 5412 4024
rect 3838 4022 3844 4023
rect 3800 3991 3802 4022
rect 3159 3990 3163 3991
rect 3159 3985 3163 3986
rect 3175 3990 3179 3991
rect 3175 3985 3179 3986
rect 3351 3990 3355 3991
rect 3351 3985 3355 3986
rect 3799 3990 3803 3991
rect 3799 3985 3803 3986
rect 3176 3961 3178 3985
rect 3352 3961 3354 3985
rect 3800 3962 3802 3985
rect 3840 3979 3842 4022
rect 4592 3979 4594 4023
rect 4706 4022 4712 4023
rect 4728 3979 4730 4023
rect 4842 4022 4848 4023
rect 4864 3979 4866 4023
rect 4958 4022 4964 4023
rect 3839 3978 3843 3979
rect 3839 3973 3843 3974
rect 4359 3978 4363 3979
rect 4359 3973 4363 3974
rect 4543 3978 4547 3979
rect 4543 3973 4547 3974
rect 4591 3978 4595 3979
rect 4591 3973 4595 3974
rect 4727 3978 4731 3979
rect 4727 3973 4731 3974
rect 4735 3978 4739 3979
rect 4735 3973 4739 3974
rect 4863 3978 4867 3979
rect 4863 3973 4867 3974
rect 4927 3978 4931 3979
rect 4927 3973 4931 3974
rect 3798 3961 3804 3962
rect 3174 3960 3180 3961
rect 3350 3960 3356 3961
rect 2830 3956 2831 3960
rect 2835 3956 2836 3960
rect 2830 3955 2836 3956
rect 2926 3959 2932 3960
rect 2926 3955 2927 3959
rect 2931 3955 2932 3959
rect 2998 3956 2999 3960
rect 3003 3956 3004 3960
rect 2998 3955 3004 3956
rect 3138 3959 3144 3960
rect 3138 3955 3139 3959
rect 3143 3955 3144 3959
rect 3174 3956 3175 3960
rect 3179 3956 3180 3960
rect 3174 3955 3180 3956
rect 3266 3959 3272 3960
rect 3266 3955 3267 3959
rect 3271 3955 3272 3959
rect 3350 3956 3351 3960
rect 3355 3956 3356 3960
rect 3350 3955 3356 3956
rect 3446 3959 3452 3960
rect 3446 3955 3447 3959
rect 3451 3955 3452 3959
rect 3798 3957 3799 3961
rect 3803 3957 3804 3961
rect 3798 3956 3804 3957
rect 2578 3954 2584 3955
rect 2926 3954 2932 3955
rect 3138 3954 3144 3955
rect 3266 3954 3272 3955
rect 3446 3954 3452 3955
rect 2282 3945 2288 3946
rect 2282 3941 2283 3945
rect 2287 3941 2288 3945
rect 2282 3940 2288 3941
rect 2458 3945 2464 3946
rect 2458 3941 2459 3945
rect 2463 3941 2464 3945
rect 2458 3940 2464 3941
rect 2194 3895 2200 3896
rect 2194 3891 2195 3895
rect 2199 3891 2200 3895
rect 2194 3890 2200 3891
rect 2284 3871 2286 3940
rect 2460 3871 2462 3940
rect 1975 3870 1979 3871
rect 1975 3865 1979 3866
rect 2099 3870 2103 3871
rect 2099 3865 2103 3866
rect 2283 3870 2287 3871
rect 2283 3865 2287 3866
rect 2291 3870 2295 3871
rect 2291 3865 2295 3866
rect 2459 3870 2463 3871
rect 2459 3865 2463 3866
rect 2523 3870 2527 3871
rect 2523 3865 2527 3866
rect 1515 3838 1519 3839
rect 1515 3833 1519 3834
rect 1547 3838 1551 3839
rect 1547 3833 1551 3834
rect 1787 3838 1791 3839
rect 1787 3833 1791 3834
rect 1935 3838 1939 3839
rect 1935 3833 1939 3834
rect 1516 3772 1518 3833
rect 1610 3819 1616 3820
rect 1610 3815 1611 3819
rect 1615 3815 1616 3819
rect 1610 3814 1616 3815
rect 1612 3796 1614 3814
rect 1610 3795 1616 3796
rect 1610 3791 1611 3795
rect 1615 3791 1616 3795
rect 1610 3790 1616 3791
rect 1788 3772 1790 3833
rect 1854 3823 1860 3824
rect 1854 3819 1855 3823
rect 1859 3819 1860 3823
rect 1854 3818 1860 3819
rect 1514 3771 1520 3772
rect 1514 3767 1515 3771
rect 1519 3767 1520 3771
rect 1514 3766 1520 3767
rect 1786 3771 1792 3772
rect 1786 3767 1787 3771
rect 1791 3767 1792 3771
rect 1786 3766 1792 3767
rect 1378 3763 1384 3764
rect 1378 3759 1379 3763
rect 1383 3759 1384 3763
rect 1378 3758 1384 3759
rect 1262 3756 1268 3757
rect 110 3755 116 3756
rect 110 3751 111 3755
rect 115 3751 116 3755
rect 294 3752 295 3756
rect 299 3752 300 3756
rect 294 3751 300 3752
rect 482 3755 488 3756
rect 482 3751 483 3755
rect 487 3751 488 3755
rect 502 3752 503 3756
rect 507 3752 508 3756
rect 502 3751 508 3752
rect 714 3755 720 3756
rect 714 3751 715 3755
rect 719 3751 720 3755
rect 734 3752 735 3756
rect 739 3752 740 3756
rect 734 3751 740 3752
rect 970 3755 976 3756
rect 970 3751 971 3755
rect 975 3751 976 3755
rect 990 3752 991 3756
rect 995 3752 996 3756
rect 990 3751 996 3752
rect 1242 3755 1248 3756
rect 1242 3751 1243 3755
rect 1247 3751 1248 3755
rect 1262 3752 1263 3756
rect 1267 3752 1268 3756
rect 1262 3751 1268 3752
rect 1542 3756 1548 3757
rect 1542 3752 1543 3756
rect 1547 3752 1548 3756
rect 1542 3751 1548 3752
rect 1814 3756 1820 3757
rect 1814 3752 1815 3756
rect 1819 3752 1820 3756
rect 1814 3751 1820 3752
rect 110 3750 116 3751
rect 112 3723 114 3750
rect 296 3723 298 3751
rect 482 3750 488 3751
rect 504 3723 506 3751
rect 714 3750 720 3751
rect 698 3739 704 3740
rect 698 3735 699 3739
rect 703 3735 704 3739
rect 698 3734 704 3735
rect 111 3722 115 3723
rect 111 3717 115 3718
rect 295 3722 299 3723
rect 295 3717 299 3718
rect 503 3722 507 3723
rect 503 3717 507 3718
rect 631 3722 635 3723
rect 631 3717 635 3718
rect 112 3694 114 3717
rect 110 3693 116 3694
rect 632 3693 634 3717
rect 110 3689 111 3693
rect 115 3689 116 3693
rect 110 3688 116 3689
rect 630 3692 636 3693
rect 630 3688 631 3692
rect 635 3688 636 3692
rect 630 3687 636 3688
rect 602 3677 608 3678
rect 110 3676 116 3677
rect 110 3672 111 3676
rect 115 3672 116 3676
rect 602 3673 603 3677
rect 607 3673 608 3677
rect 602 3672 608 3673
rect 110 3671 116 3672
rect 112 3599 114 3671
rect 604 3599 606 3672
rect 700 3628 702 3734
rect 736 3723 738 3751
rect 970 3750 976 3751
rect 992 3723 994 3751
rect 1242 3750 1248 3751
rect 1264 3723 1266 3751
rect 1544 3723 1546 3751
rect 1816 3723 1818 3751
rect 735 3722 739 3723
rect 735 3717 739 3718
rect 775 3722 779 3723
rect 775 3717 779 3718
rect 927 3722 931 3723
rect 927 3717 931 3718
rect 991 3722 995 3723
rect 991 3717 995 3718
rect 1087 3722 1091 3723
rect 1087 3717 1091 3718
rect 1255 3722 1259 3723
rect 1255 3717 1259 3718
rect 1263 3722 1267 3723
rect 1263 3717 1267 3718
rect 1423 3722 1427 3723
rect 1423 3717 1427 3718
rect 1543 3722 1547 3723
rect 1543 3717 1547 3718
rect 1591 3722 1595 3723
rect 1591 3717 1595 3718
rect 1759 3722 1763 3723
rect 1759 3717 1763 3718
rect 1815 3722 1819 3723
rect 1815 3717 1819 3718
rect 776 3693 778 3717
rect 928 3693 930 3717
rect 1088 3693 1090 3717
rect 1256 3693 1258 3717
rect 1424 3693 1426 3717
rect 1592 3693 1594 3717
rect 1760 3693 1762 3717
rect 774 3692 780 3693
rect 730 3691 736 3692
rect 730 3687 731 3691
rect 735 3687 736 3691
rect 774 3688 775 3692
rect 779 3688 780 3692
rect 774 3687 780 3688
rect 926 3692 932 3693
rect 1086 3692 1092 3693
rect 1254 3692 1260 3693
rect 1422 3692 1428 3693
rect 1590 3692 1596 3693
rect 1758 3692 1764 3693
rect 1856 3692 1858 3818
rect 1910 3795 1916 3796
rect 1910 3791 1911 3795
rect 1915 3791 1916 3795
rect 1910 3790 1916 3791
rect 1912 3756 1914 3790
rect 1936 3773 1938 3833
rect 1976 3805 1978 3865
rect 1974 3804 1980 3805
rect 2292 3804 2294 3865
rect 2524 3804 2526 3865
rect 2580 3864 2582 3954
rect 2634 3945 2640 3946
rect 2634 3941 2635 3945
rect 2639 3941 2640 3945
rect 2634 3940 2640 3941
rect 2802 3945 2808 3946
rect 2802 3941 2803 3945
rect 2807 3941 2808 3945
rect 2802 3940 2808 3941
rect 2636 3871 2638 3940
rect 2730 3923 2736 3924
rect 2730 3919 2731 3923
rect 2735 3919 2736 3923
rect 2730 3918 2736 3919
rect 2732 3896 2734 3918
rect 2730 3895 2736 3896
rect 2730 3891 2731 3895
rect 2735 3891 2736 3895
rect 2730 3890 2736 3891
rect 2804 3871 2806 3940
rect 2928 3896 2930 3954
rect 2970 3945 2976 3946
rect 2970 3941 2971 3945
rect 2975 3941 2976 3945
rect 2970 3940 2976 3941
rect 3146 3945 3152 3946
rect 3146 3941 3147 3945
rect 3151 3941 3152 3945
rect 3146 3940 3152 3941
rect 2926 3895 2932 3896
rect 2926 3891 2927 3895
rect 2931 3891 2932 3895
rect 2926 3890 2932 3891
rect 2972 3871 2974 3940
rect 3148 3871 3150 3940
rect 3268 3924 3270 3954
rect 3322 3945 3328 3946
rect 3322 3941 3323 3945
rect 3327 3941 3328 3945
rect 3322 3940 3328 3941
rect 3266 3923 3272 3924
rect 3266 3919 3267 3923
rect 3271 3919 3272 3923
rect 3266 3918 3272 3919
rect 3282 3895 3288 3896
rect 3282 3891 3283 3895
rect 3287 3891 3288 3895
rect 3282 3890 3288 3891
rect 2635 3870 2639 3871
rect 2635 3865 2639 3866
rect 2739 3870 2743 3871
rect 2739 3865 2743 3866
rect 2803 3870 2807 3871
rect 2803 3865 2807 3866
rect 2947 3870 2951 3871
rect 2947 3865 2951 3866
rect 2971 3870 2975 3871
rect 2971 3865 2975 3866
rect 3147 3870 3151 3871
rect 3147 3865 3151 3866
rect 3155 3870 3159 3871
rect 3155 3865 3159 3866
rect 2578 3863 2584 3864
rect 2578 3859 2579 3863
rect 2583 3859 2584 3863
rect 2578 3858 2584 3859
rect 2530 3851 2536 3852
rect 2530 3847 2531 3851
rect 2535 3847 2536 3851
rect 2530 3846 2536 3847
rect 1974 3800 1975 3804
rect 1979 3800 1980 3804
rect 1974 3799 1980 3800
rect 2290 3803 2296 3804
rect 2290 3799 2291 3803
rect 2295 3799 2296 3803
rect 2290 3798 2296 3799
rect 2522 3803 2528 3804
rect 2522 3799 2523 3803
rect 2527 3799 2528 3803
rect 2522 3798 2528 3799
rect 2318 3788 2324 3789
rect 2532 3788 2534 3846
rect 2740 3804 2742 3865
rect 2938 3855 2944 3856
rect 2938 3851 2939 3855
rect 2943 3851 2944 3855
rect 2938 3850 2944 3851
rect 2738 3803 2744 3804
rect 2738 3799 2739 3803
rect 2743 3799 2744 3803
rect 2738 3798 2744 3799
rect 2940 3796 2942 3850
rect 2948 3804 2950 3865
rect 2954 3851 2960 3852
rect 2954 3847 2955 3851
rect 2959 3847 2960 3851
rect 2954 3846 2960 3847
rect 2946 3803 2952 3804
rect 2946 3799 2947 3803
rect 2951 3799 2952 3803
rect 2946 3798 2952 3799
rect 2938 3795 2944 3796
rect 2938 3791 2939 3795
rect 2943 3791 2944 3795
rect 2938 3790 2944 3791
rect 2550 3788 2556 3789
rect 2766 3788 2772 3789
rect 2956 3788 2958 3846
rect 3156 3804 3158 3865
rect 3162 3851 3168 3852
rect 3162 3847 3163 3851
rect 3167 3847 3168 3851
rect 3162 3846 3168 3847
rect 3154 3803 3160 3804
rect 3154 3799 3155 3803
rect 3159 3799 3160 3803
rect 3154 3798 3160 3799
rect 2974 3788 2980 3789
rect 3164 3788 3166 3846
rect 3182 3788 3188 3789
rect 3284 3788 3286 3890
rect 3324 3871 3326 3940
rect 3448 3888 3450 3954
rect 3840 3950 3842 3973
rect 3838 3949 3844 3950
rect 4360 3949 4362 3973
rect 4544 3949 4546 3973
rect 4736 3949 4738 3973
rect 4928 3949 4930 3973
rect 3838 3945 3839 3949
rect 3843 3945 3844 3949
rect 3798 3944 3804 3945
rect 3838 3944 3844 3945
rect 4358 3948 4364 3949
rect 4542 3948 4548 3949
rect 4734 3948 4740 3949
rect 4926 3948 4932 3949
rect 4358 3944 4359 3948
rect 4363 3944 4364 3948
rect 3798 3940 3799 3944
rect 3803 3940 3804 3944
rect 4358 3943 4364 3944
rect 4470 3947 4476 3948
rect 4470 3943 4471 3947
rect 4475 3943 4476 3947
rect 4542 3944 4543 3948
rect 4547 3944 4548 3948
rect 4542 3943 4548 3944
rect 4642 3947 4648 3948
rect 4642 3943 4643 3947
rect 4647 3943 4648 3947
rect 4734 3944 4735 3948
rect 4739 3944 4740 3948
rect 4734 3943 4740 3944
rect 4826 3947 4832 3948
rect 4826 3943 4827 3947
rect 4831 3943 4832 3947
rect 4926 3944 4927 3948
rect 4931 3944 4932 3948
rect 4926 3943 4932 3944
rect 4470 3942 4476 3943
rect 4642 3942 4648 3943
rect 4826 3942 4832 3943
rect 3798 3939 3804 3940
rect 3446 3887 3452 3888
rect 3446 3883 3447 3887
rect 3451 3883 3452 3887
rect 3446 3882 3452 3883
rect 3800 3871 3802 3939
rect 4330 3933 4336 3934
rect 3838 3932 3844 3933
rect 3838 3928 3839 3932
rect 3843 3928 3844 3932
rect 4330 3929 4331 3933
rect 4335 3929 4336 3933
rect 4330 3928 4336 3929
rect 3838 3927 3844 3928
rect 3323 3870 3327 3871
rect 3323 3865 3327 3866
rect 3355 3870 3359 3871
rect 3355 3865 3359 3866
rect 3563 3870 3567 3871
rect 3563 3865 3567 3866
rect 3799 3870 3803 3871
rect 3799 3865 3803 3866
rect 3356 3804 3358 3865
rect 3390 3855 3396 3856
rect 3390 3851 3391 3855
rect 3395 3851 3396 3855
rect 3390 3850 3396 3851
rect 3354 3803 3360 3804
rect 3354 3799 3355 3803
rect 3359 3799 3360 3803
rect 3354 3798 3360 3799
rect 3382 3788 3388 3789
rect 1974 3787 1980 3788
rect 1974 3783 1975 3787
rect 1979 3783 1980 3787
rect 2318 3784 2319 3788
rect 2323 3784 2324 3788
rect 2318 3783 2324 3784
rect 2530 3787 2536 3788
rect 2530 3783 2531 3787
rect 2535 3783 2536 3787
rect 2550 3784 2551 3788
rect 2555 3784 2556 3788
rect 2550 3783 2556 3784
rect 2646 3787 2652 3788
rect 2646 3783 2647 3787
rect 2651 3783 2652 3787
rect 2766 3784 2767 3788
rect 2771 3784 2772 3788
rect 2766 3783 2772 3784
rect 2954 3787 2960 3788
rect 2954 3783 2955 3787
rect 2959 3783 2960 3787
rect 2974 3784 2975 3788
rect 2979 3784 2980 3788
rect 2974 3783 2980 3784
rect 3162 3787 3168 3788
rect 3162 3783 3163 3787
rect 3167 3783 3168 3787
rect 3182 3784 3183 3788
rect 3187 3784 3188 3788
rect 3182 3783 3188 3784
rect 3282 3787 3288 3788
rect 3282 3783 3283 3787
rect 3287 3783 3288 3787
rect 3382 3784 3383 3788
rect 3387 3784 3388 3788
rect 3382 3783 3388 3784
rect 1974 3782 1980 3783
rect 1934 3772 1940 3773
rect 1934 3768 1935 3772
rect 1939 3768 1940 3772
rect 1934 3767 1940 3768
rect 1910 3755 1916 3756
rect 1910 3751 1911 3755
rect 1915 3751 1916 3755
rect 1910 3750 1916 3751
rect 1934 3755 1940 3756
rect 1976 3755 1978 3782
rect 2320 3755 2322 3783
rect 2530 3782 2536 3783
rect 2552 3755 2554 3783
rect 2646 3782 2652 3783
rect 2648 3779 2650 3782
rect 2640 3777 2650 3779
rect 1934 3751 1935 3755
rect 1939 3751 1940 3755
rect 1934 3750 1940 3751
rect 1975 3754 1979 3755
rect 1936 3723 1938 3750
rect 1975 3749 1979 3750
rect 2319 3754 2323 3755
rect 2319 3749 2323 3750
rect 2407 3754 2411 3755
rect 2407 3749 2411 3750
rect 2551 3754 2555 3755
rect 2551 3749 2555 3750
rect 1976 3726 1978 3749
rect 1974 3725 1980 3726
rect 2408 3725 2410 3749
rect 1935 3722 1939 3723
rect 1974 3721 1975 3725
rect 1979 3721 1980 3725
rect 1974 3720 1980 3721
rect 2406 3724 2412 3725
rect 2406 3720 2407 3724
rect 2411 3720 2412 3724
rect 2406 3719 2412 3720
rect 2502 3723 2508 3724
rect 2502 3719 2503 3723
rect 2507 3719 2508 3723
rect 2502 3718 2508 3719
rect 1935 3717 1939 3718
rect 1936 3694 1938 3717
rect 2378 3709 2384 3710
rect 1974 3708 1980 3709
rect 1974 3704 1975 3708
rect 1979 3704 1980 3708
rect 2378 3705 2379 3709
rect 2383 3705 2384 3709
rect 2378 3704 2384 3705
rect 1974 3703 1980 3704
rect 1934 3693 1940 3694
rect 926 3688 927 3692
rect 931 3688 932 3692
rect 926 3687 932 3688
rect 1026 3691 1032 3692
rect 1026 3687 1027 3691
rect 1031 3687 1032 3691
rect 1086 3688 1087 3692
rect 1091 3688 1092 3692
rect 1086 3687 1092 3688
rect 1186 3691 1192 3692
rect 1186 3687 1187 3691
rect 1191 3687 1192 3691
rect 1254 3688 1255 3692
rect 1259 3688 1260 3692
rect 1254 3687 1260 3688
rect 1346 3691 1352 3692
rect 1346 3687 1347 3691
rect 1351 3687 1352 3691
rect 1422 3688 1423 3692
rect 1427 3688 1428 3692
rect 1422 3687 1428 3688
rect 1522 3691 1528 3692
rect 1522 3687 1523 3691
rect 1527 3687 1528 3691
rect 1590 3688 1591 3692
rect 1595 3688 1596 3692
rect 1590 3687 1596 3688
rect 1690 3691 1696 3692
rect 1690 3687 1691 3691
rect 1695 3687 1696 3691
rect 1758 3688 1759 3692
rect 1763 3688 1764 3692
rect 1758 3687 1764 3688
rect 1854 3691 1860 3692
rect 1854 3687 1855 3691
rect 1859 3687 1860 3691
rect 1934 3689 1935 3693
rect 1939 3689 1940 3693
rect 1934 3688 1940 3689
rect 730 3686 736 3687
rect 1026 3686 1032 3687
rect 1186 3686 1192 3687
rect 1346 3686 1352 3687
rect 1522 3686 1528 3687
rect 1690 3686 1696 3687
rect 1854 3686 1860 3687
rect 732 3628 734 3686
rect 746 3677 752 3678
rect 746 3673 747 3677
rect 751 3673 752 3677
rect 746 3672 752 3673
rect 898 3677 904 3678
rect 898 3673 899 3677
rect 903 3673 904 3677
rect 898 3672 904 3673
rect 698 3627 704 3628
rect 698 3623 699 3627
rect 703 3623 704 3627
rect 698 3622 704 3623
rect 730 3627 736 3628
rect 730 3623 731 3627
rect 735 3623 736 3627
rect 730 3622 736 3623
rect 748 3599 750 3672
rect 900 3599 902 3672
rect 1028 3628 1030 3686
rect 1058 3677 1064 3678
rect 1058 3673 1059 3677
rect 1063 3673 1064 3677
rect 1058 3672 1064 3673
rect 1026 3627 1032 3628
rect 1026 3623 1027 3627
rect 1031 3623 1032 3627
rect 1026 3622 1032 3623
rect 1060 3599 1062 3672
rect 1188 3628 1190 3686
rect 1226 3677 1232 3678
rect 1226 3673 1227 3677
rect 1231 3673 1232 3677
rect 1226 3672 1232 3673
rect 1186 3627 1192 3628
rect 1186 3623 1187 3627
rect 1191 3623 1192 3627
rect 1186 3622 1192 3623
rect 1228 3599 1230 3672
rect 111 3598 115 3599
rect 111 3593 115 3594
rect 603 3598 607 3599
rect 603 3593 607 3594
rect 747 3598 751 3599
rect 747 3593 751 3594
rect 779 3598 783 3599
rect 779 3593 783 3594
rect 899 3598 903 3599
rect 899 3593 903 3594
rect 915 3598 919 3599
rect 915 3593 919 3594
rect 1051 3598 1055 3599
rect 1051 3593 1055 3594
rect 1059 3598 1063 3599
rect 1059 3593 1063 3594
rect 1187 3598 1191 3599
rect 1187 3593 1191 3594
rect 1227 3598 1231 3599
rect 1227 3593 1231 3594
rect 1323 3598 1327 3599
rect 1323 3593 1327 3594
rect 112 3533 114 3593
rect 110 3532 116 3533
rect 780 3532 782 3593
rect 916 3532 918 3593
rect 922 3579 928 3580
rect 922 3575 923 3579
rect 927 3575 928 3579
rect 922 3574 928 3575
rect 110 3528 111 3532
rect 115 3528 116 3532
rect 110 3527 116 3528
rect 778 3531 784 3532
rect 778 3527 779 3531
rect 783 3527 784 3531
rect 778 3526 784 3527
rect 914 3531 920 3532
rect 914 3527 915 3531
rect 919 3527 920 3531
rect 914 3526 920 3527
rect 806 3516 812 3517
rect 924 3516 926 3574
rect 1052 3532 1054 3593
rect 1058 3579 1064 3580
rect 1058 3575 1059 3579
rect 1063 3575 1064 3579
rect 1058 3574 1064 3575
rect 1050 3531 1056 3532
rect 1050 3527 1051 3531
rect 1055 3527 1056 3531
rect 1050 3526 1056 3527
rect 942 3516 948 3517
rect 1060 3516 1062 3574
rect 1188 3532 1190 3593
rect 1194 3579 1200 3580
rect 1194 3575 1195 3579
rect 1199 3575 1200 3579
rect 1194 3574 1200 3575
rect 1186 3531 1192 3532
rect 1186 3527 1187 3531
rect 1191 3527 1192 3531
rect 1186 3526 1192 3527
rect 1078 3516 1084 3517
rect 1196 3516 1198 3574
rect 1324 3532 1326 3593
rect 1348 3592 1350 3686
rect 1394 3677 1400 3678
rect 1394 3673 1395 3677
rect 1399 3673 1400 3677
rect 1394 3672 1400 3673
rect 1396 3599 1398 3672
rect 1524 3628 1526 3686
rect 1562 3677 1568 3678
rect 1562 3673 1563 3677
rect 1567 3673 1568 3677
rect 1562 3672 1568 3673
rect 1522 3627 1528 3628
rect 1522 3623 1523 3627
rect 1527 3623 1528 3627
rect 1522 3622 1528 3623
rect 1564 3599 1566 3672
rect 1692 3628 1694 3686
rect 1730 3677 1736 3678
rect 1730 3673 1731 3677
rect 1735 3673 1736 3677
rect 1730 3672 1736 3673
rect 1934 3676 1940 3677
rect 1934 3672 1935 3676
rect 1939 3672 1940 3676
rect 1690 3627 1696 3628
rect 1690 3623 1691 3627
rect 1695 3623 1696 3627
rect 1690 3622 1696 3623
rect 1732 3599 1734 3672
rect 1934 3671 1940 3672
rect 1850 3619 1856 3620
rect 1850 3615 1851 3619
rect 1855 3615 1856 3619
rect 1850 3614 1856 3615
rect 1395 3598 1399 3599
rect 1395 3593 1399 3594
rect 1459 3598 1463 3599
rect 1459 3593 1463 3594
rect 1563 3598 1567 3599
rect 1563 3593 1567 3594
rect 1595 3598 1599 3599
rect 1595 3593 1599 3594
rect 1731 3598 1735 3599
rect 1731 3593 1735 3594
rect 1346 3591 1352 3592
rect 1346 3587 1347 3591
rect 1351 3587 1352 3591
rect 1346 3586 1352 3587
rect 1370 3591 1376 3592
rect 1370 3587 1371 3591
rect 1375 3587 1376 3591
rect 1370 3586 1376 3587
rect 1330 3579 1336 3580
rect 1330 3575 1331 3579
rect 1335 3575 1336 3579
rect 1330 3574 1336 3575
rect 1322 3531 1328 3532
rect 1322 3527 1323 3531
rect 1327 3527 1328 3531
rect 1322 3526 1328 3527
rect 1214 3516 1220 3517
rect 1332 3516 1334 3574
rect 1350 3516 1356 3517
rect 110 3515 116 3516
rect 110 3511 111 3515
rect 115 3511 116 3515
rect 806 3512 807 3516
rect 811 3512 812 3516
rect 806 3511 812 3512
rect 922 3515 928 3516
rect 922 3511 923 3515
rect 927 3511 928 3515
rect 942 3512 943 3516
rect 947 3512 948 3516
rect 942 3511 948 3512
rect 1058 3515 1064 3516
rect 1058 3511 1059 3515
rect 1063 3511 1064 3515
rect 1078 3512 1079 3516
rect 1083 3512 1084 3516
rect 1078 3511 1084 3512
rect 1194 3515 1200 3516
rect 1194 3511 1195 3515
rect 1199 3511 1200 3515
rect 1214 3512 1215 3516
rect 1219 3512 1220 3516
rect 1214 3511 1220 3512
rect 1330 3515 1336 3516
rect 1330 3511 1331 3515
rect 1335 3511 1336 3515
rect 1350 3512 1351 3516
rect 1355 3512 1356 3516
rect 1350 3511 1356 3512
rect 110 3510 116 3511
rect 112 3463 114 3510
rect 808 3463 810 3511
rect 922 3510 928 3511
rect 944 3463 946 3511
rect 1058 3510 1064 3511
rect 1080 3463 1082 3511
rect 1194 3510 1200 3511
rect 1216 3463 1218 3511
rect 1330 3510 1336 3511
rect 1352 3463 1354 3511
rect 111 3462 115 3463
rect 111 3457 115 3458
rect 727 3462 731 3463
rect 727 3457 731 3458
rect 807 3462 811 3463
rect 807 3457 811 3458
rect 863 3462 867 3463
rect 863 3457 867 3458
rect 943 3462 947 3463
rect 943 3457 947 3458
rect 999 3462 1003 3463
rect 999 3457 1003 3458
rect 1079 3462 1083 3463
rect 1079 3457 1083 3458
rect 1135 3462 1139 3463
rect 1135 3457 1139 3458
rect 1215 3462 1219 3463
rect 1215 3457 1219 3458
rect 1271 3462 1275 3463
rect 1271 3457 1275 3458
rect 1351 3462 1355 3463
rect 1351 3457 1355 3458
rect 112 3434 114 3457
rect 110 3433 116 3434
rect 728 3433 730 3457
rect 864 3433 866 3457
rect 1000 3433 1002 3457
rect 1136 3433 1138 3457
rect 1272 3433 1274 3457
rect 110 3429 111 3433
rect 115 3429 116 3433
rect 110 3428 116 3429
rect 726 3432 732 3433
rect 862 3432 868 3433
rect 998 3432 1004 3433
rect 726 3428 727 3432
rect 731 3428 732 3432
rect 726 3427 732 3428
rect 826 3431 832 3432
rect 826 3427 827 3431
rect 831 3427 832 3431
rect 862 3428 863 3432
rect 867 3428 868 3432
rect 862 3427 868 3428
rect 962 3431 968 3432
rect 962 3427 963 3431
rect 967 3427 968 3431
rect 998 3428 999 3432
rect 1003 3428 1004 3432
rect 998 3427 1004 3428
rect 1134 3432 1140 3433
rect 1270 3432 1276 3433
rect 1372 3432 1374 3586
rect 1460 3532 1462 3593
rect 1596 3532 1598 3593
rect 1602 3579 1608 3580
rect 1602 3575 1603 3579
rect 1607 3575 1608 3579
rect 1602 3574 1608 3575
rect 1458 3531 1464 3532
rect 1458 3527 1459 3531
rect 1463 3527 1464 3531
rect 1458 3526 1464 3527
rect 1594 3531 1600 3532
rect 1594 3527 1595 3531
rect 1599 3527 1600 3531
rect 1594 3526 1600 3527
rect 1486 3516 1492 3517
rect 1604 3516 1606 3574
rect 1732 3532 1734 3593
rect 1738 3579 1744 3580
rect 1738 3575 1739 3579
rect 1743 3575 1744 3579
rect 1738 3574 1744 3575
rect 1730 3531 1736 3532
rect 1730 3527 1731 3531
rect 1735 3527 1736 3531
rect 1730 3526 1736 3527
rect 1622 3516 1628 3517
rect 1740 3516 1742 3574
rect 1758 3516 1764 3517
rect 1852 3516 1854 3614
rect 1936 3599 1938 3671
rect 1976 3635 1978 3703
rect 2380 3635 2382 3704
rect 1975 3634 1979 3635
rect 1975 3629 1979 3630
rect 2379 3634 2383 3635
rect 2379 3629 2383 3630
rect 2411 3634 2415 3635
rect 2411 3629 2415 3630
rect 1935 3598 1939 3599
rect 1935 3593 1939 3594
rect 1936 3533 1938 3593
rect 1976 3569 1978 3629
rect 1974 3568 1980 3569
rect 2412 3568 2414 3629
rect 2504 3620 2506 3718
rect 2618 3709 2624 3710
rect 2618 3705 2619 3709
rect 2623 3705 2624 3709
rect 2618 3704 2624 3705
rect 2620 3635 2622 3704
rect 2640 3660 2642 3777
rect 2768 3755 2770 3783
rect 2954 3782 2960 3783
rect 2976 3755 2978 3783
rect 3162 3782 3168 3783
rect 3184 3755 3186 3783
rect 3282 3782 3288 3783
rect 3384 3755 3386 3783
rect 2647 3754 2651 3755
rect 2647 3749 2651 3750
rect 2767 3754 2771 3755
rect 2767 3749 2771 3750
rect 2871 3754 2875 3755
rect 2871 3749 2875 3750
rect 2975 3754 2979 3755
rect 2975 3749 2979 3750
rect 3087 3754 3091 3755
rect 3087 3749 3091 3750
rect 3183 3754 3187 3755
rect 3183 3749 3187 3750
rect 3295 3754 3299 3755
rect 3295 3749 3299 3750
rect 3383 3754 3387 3755
rect 3383 3749 3387 3750
rect 2648 3725 2650 3749
rect 2872 3725 2874 3749
rect 3088 3725 3090 3749
rect 3296 3725 3298 3749
rect 2646 3724 2652 3725
rect 2870 3724 2876 3725
rect 3086 3724 3092 3725
rect 3294 3724 3300 3725
rect 3392 3724 3394 3850
rect 3564 3804 3566 3865
rect 3570 3851 3576 3852
rect 3570 3847 3571 3851
rect 3575 3847 3576 3851
rect 3570 3846 3576 3847
rect 3562 3803 3568 3804
rect 3562 3799 3563 3803
rect 3567 3799 3568 3803
rect 3562 3798 3568 3799
rect 3572 3788 3574 3846
rect 3800 3805 3802 3865
rect 3840 3859 3842 3927
rect 4332 3859 4334 3928
rect 4426 3915 4432 3916
rect 4426 3911 4427 3915
rect 4431 3911 4432 3915
rect 4426 3910 4432 3911
rect 4428 3884 4430 3910
rect 4472 3884 4474 3942
rect 4514 3933 4520 3934
rect 4514 3929 4515 3933
rect 4519 3929 4520 3933
rect 4514 3928 4520 3929
rect 4426 3883 4432 3884
rect 4426 3879 4427 3883
rect 4431 3879 4432 3883
rect 4426 3878 4432 3879
rect 4470 3883 4476 3884
rect 4470 3879 4471 3883
rect 4475 3879 4476 3883
rect 4470 3878 4476 3879
rect 4516 3859 4518 3928
rect 3839 3858 3843 3859
rect 3839 3853 3843 3854
rect 4051 3858 4055 3859
rect 4051 3853 4055 3854
rect 4267 3858 4271 3859
rect 4267 3853 4271 3854
rect 4331 3858 4335 3859
rect 4331 3853 4335 3854
rect 4483 3858 4487 3859
rect 4483 3853 4487 3854
rect 4515 3858 4519 3859
rect 4515 3853 4519 3854
rect 3798 3804 3804 3805
rect 3798 3800 3799 3804
rect 3803 3800 3804 3804
rect 3798 3799 3804 3800
rect 3840 3793 3842 3853
rect 3838 3792 3844 3793
rect 4052 3792 4054 3853
rect 4268 3792 4270 3853
rect 4474 3843 4480 3844
rect 4474 3839 4475 3843
rect 4479 3839 4480 3843
rect 4474 3838 4480 3839
rect 3590 3788 3596 3789
rect 3838 3788 3839 3792
rect 3843 3788 3844 3792
rect 3570 3787 3576 3788
rect 3570 3783 3571 3787
rect 3575 3783 3576 3787
rect 3590 3784 3591 3788
rect 3595 3784 3596 3788
rect 3590 3783 3596 3784
rect 3798 3787 3804 3788
rect 3838 3787 3844 3788
rect 4050 3791 4056 3792
rect 4050 3787 4051 3791
rect 4055 3787 4056 3791
rect 3798 3783 3799 3787
rect 3803 3783 3804 3787
rect 4050 3786 4056 3787
rect 4266 3791 4272 3792
rect 4266 3787 4267 3791
rect 4271 3787 4272 3791
rect 4266 3786 4272 3787
rect 4476 3784 4478 3838
rect 4484 3792 4486 3853
rect 4644 3844 4646 3942
rect 4706 3933 4712 3934
rect 4706 3929 4707 3933
rect 4711 3929 4712 3933
rect 4706 3928 4712 3929
rect 4708 3859 4710 3928
rect 4828 3916 4830 3942
rect 4898 3933 4904 3934
rect 4898 3929 4899 3933
rect 4903 3929 4904 3933
rect 4898 3928 4904 3929
rect 4826 3915 4832 3916
rect 4826 3911 4827 3915
rect 4831 3911 4832 3915
rect 4826 3910 4832 3911
rect 4900 3859 4902 3928
rect 4960 3884 4962 4022
rect 5000 3979 5002 4023
rect 5090 4022 5096 4023
rect 5136 3979 5138 4023
rect 5230 4022 5236 4023
rect 5272 3979 5274 4023
rect 5366 4022 5372 4023
rect 5408 3979 5410 4023
rect 4999 3978 5003 3979
rect 4999 3973 5003 3974
rect 5127 3978 5131 3979
rect 5127 3973 5131 3974
rect 5135 3978 5139 3979
rect 5135 3973 5139 3974
rect 5271 3978 5275 3979
rect 5271 3973 5275 3974
rect 5327 3978 5331 3979
rect 5327 3973 5331 3974
rect 5407 3978 5411 3979
rect 5407 3973 5411 3974
rect 5128 3949 5130 3973
rect 5328 3949 5330 3973
rect 5126 3948 5132 3949
rect 5022 3947 5028 3948
rect 5022 3943 5023 3947
rect 5027 3943 5028 3947
rect 5126 3944 5127 3948
rect 5131 3944 5132 3948
rect 5126 3943 5132 3944
rect 5326 3948 5332 3949
rect 5424 3948 5426 4090
rect 5498 4055 5504 4056
rect 5498 4051 5499 4055
rect 5503 4051 5504 4055
rect 5498 4050 5504 4051
rect 5500 4028 5502 4050
rect 5516 4044 5518 4105
rect 5664 4045 5666 4105
rect 5662 4044 5668 4045
rect 5514 4043 5520 4044
rect 5514 4039 5515 4043
rect 5519 4039 5520 4043
rect 5662 4040 5663 4044
rect 5667 4040 5668 4044
rect 5662 4039 5668 4040
rect 5514 4038 5520 4039
rect 5542 4028 5548 4029
rect 5498 4027 5504 4028
rect 5498 4023 5499 4027
rect 5503 4023 5504 4027
rect 5542 4024 5543 4028
rect 5547 4024 5548 4028
rect 5542 4023 5548 4024
rect 5638 4027 5644 4028
rect 5638 4023 5639 4027
rect 5643 4023 5644 4027
rect 5498 4022 5504 4023
rect 5544 3979 5546 4023
rect 5638 4022 5644 4023
rect 5662 4027 5668 4028
rect 5662 4023 5663 4027
rect 5667 4023 5668 4027
rect 5662 4022 5668 4023
rect 5527 3978 5531 3979
rect 5527 3973 5531 3974
rect 5543 3978 5547 3979
rect 5543 3973 5547 3974
rect 5528 3949 5530 3973
rect 5526 3948 5532 3949
rect 5326 3944 5327 3948
rect 5331 3944 5332 3948
rect 5326 3943 5332 3944
rect 5422 3947 5428 3948
rect 5422 3943 5423 3947
rect 5427 3943 5428 3947
rect 5526 3944 5527 3948
rect 5531 3944 5532 3948
rect 5526 3943 5532 3944
rect 5618 3947 5624 3948
rect 5618 3943 5619 3947
rect 5623 3943 5624 3947
rect 5022 3942 5028 3943
rect 5422 3942 5428 3943
rect 5618 3942 5624 3943
rect 4958 3883 4964 3884
rect 4958 3879 4959 3883
rect 4963 3879 4964 3883
rect 4958 3878 4964 3879
rect 5024 3876 5026 3942
rect 5098 3933 5104 3934
rect 5098 3929 5099 3933
rect 5103 3929 5104 3933
rect 5098 3928 5104 3929
rect 5298 3933 5304 3934
rect 5298 3929 5299 3933
rect 5303 3929 5304 3933
rect 5298 3928 5304 3929
rect 5498 3933 5504 3934
rect 5498 3929 5499 3933
rect 5503 3929 5504 3933
rect 5498 3928 5504 3929
rect 5034 3883 5040 3884
rect 5034 3879 5035 3883
rect 5039 3879 5040 3883
rect 5034 3878 5040 3879
rect 5022 3875 5028 3876
rect 5022 3871 5023 3875
rect 5027 3871 5028 3875
rect 5022 3870 5028 3871
rect 4699 3858 4703 3859
rect 4699 3853 4703 3854
rect 4707 3858 4711 3859
rect 4707 3853 4711 3854
rect 4899 3858 4903 3859
rect 4899 3853 4903 3854
rect 4907 3858 4911 3859
rect 4907 3853 4911 3854
rect 4634 3843 4640 3844
rect 4634 3839 4635 3843
rect 4639 3839 4640 3843
rect 4634 3838 4640 3839
rect 4642 3843 4648 3844
rect 4642 3839 4643 3843
rect 4647 3839 4648 3843
rect 4642 3838 4648 3839
rect 4482 3791 4488 3792
rect 4482 3787 4483 3791
rect 4487 3787 4488 3791
rect 4482 3786 4488 3787
rect 4636 3784 4638 3838
rect 4700 3792 4702 3853
rect 4908 3792 4910 3853
rect 4698 3791 4704 3792
rect 4698 3787 4699 3791
rect 4703 3787 4704 3791
rect 4698 3786 4704 3787
rect 4906 3791 4912 3792
rect 4906 3787 4907 3791
rect 4911 3787 4912 3791
rect 4906 3786 4912 3787
rect 3570 3782 3576 3783
rect 3592 3755 3594 3783
rect 3798 3782 3804 3783
rect 4474 3783 4480 3784
rect 3800 3755 3802 3782
rect 4474 3779 4475 3783
rect 4479 3779 4480 3783
rect 4474 3778 4480 3779
rect 4634 3783 4640 3784
rect 4634 3779 4635 3783
rect 4639 3779 4640 3783
rect 4634 3778 4640 3779
rect 4078 3776 4084 3777
rect 4294 3776 4300 3777
rect 3838 3775 3844 3776
rect 3838 3771 3839 3775
rect 3843 3771 3844 3775
rect 4078 3772 4079 3776
rect 4083 3772 4084 3776
rect 4078 3771 4084 3772
rect 4170 3775 4176 3776
rect 4170 3771 4171 3775
rect 4175 3771 4176 3775
rect 4294 3772 4295 3776
rect 4299 3772 4300 3776
rect 4294 3771 4300 3772
rect 4510 3776 4516 3777
rect 4510 3772 4511 3776
rect 4515 3772 4516 3776
rect 4510 3771 4516 3772
rect 4726 3776 4732 3777
rect 4726 3772 4727 3776
rect 4731 3772 4732 3776
rect 4726 3771 4732 3772
rect 4934 3776 4940 3777
rect 5036 3776 5038 3878
rect 5100 3859 5102 3928
rect 5300 3859 5302 3928
rect 5500 3859 5502 3928
rect 5099 3858 5103 3859
rect 5099 3853 5103 3854
rect 5115 3858 5119 3859
rect 5115 3853 5119 3854
rect 5299 3858 5303 3859
rect 5299 3853 5303 3854
rect 5323 3858 5327 3859
rect 5323 3853 5327 3854
rect 5499 3858 5503 3859
rect 5499 3853 5503 3854
rect 5515 3858 5519 3859
rect 5515 3853 5519 3854
rect 5098 3843 5104 3844
rect 5098 3839 5099 3843
rect 5103 3839 5104 3843
rect 5098 3838 5104 3839
rect 5100 3784 5102 3838
rect 5116 3792 5118 3853
rect 5324 3792 5326 3853
rect 5446 3847 5452 3848
rect 5446 3843 5447 3847
rect 5451 3843 5452 3847
rect 5446 3842 5452 3843
rect 5114 3791 5120 3792
rect 5114 3787 5115 3791
rect 5119 3787 5120 3791
rect 5114 3786 5120 3787
rect 5322 3791 5328 3792
rect 5322 3787 5323 3791
rect 5327 3787 5328 3791
rect 5322 3786 5328 3787
rect 5098 3783 5104 3784
rect 5098 3779 5099 3783
rect 5103 3779 5104 3783
rect 5098 3778 5104 3779
rect 5142 3776 5148 3777
rect 4934 3772 4935 3776
rect 4939 3772 4940 3776
rect 4934 3771 4940 3772
rect 5034 3775 5040 3776
rect 5034 3771 5035 3775
rect 5039 3771 5040 3775
rect 5142 3772 5143 3776
rect 5147 3772 5148 3776
rect 5142 3771 5148 3772
rect 5350 3776 5356 3777
rect 5448 3776 5450 3842
rect 5516 3792 5518 3853
rect 5620 3844 5622 3942
rect 5640 3884 5642 4022
rect 5664 3979 5666 4022
rect 5663 3978 5667 3979
rect 5663 3973 5667 3974
rect 5664 3950 5666 3973
rect 5662 3949 5668 3950
rect 5662 3945 5663 3949
rect 5667 3945 5668 3949
rect 5662 3944 5668 3945
rect 5662 3932 5668 3933
rect 5662 3928 5663 3932
rect 5667 3928 5668 3932
rect 5662 3927 5668 3928
rect 5638 3883 5644 3884
rect 5638 3879 5639 3883
rect 5643 3879 5644 3883
rect 5638 3878 5644 3879
rect 5664 3859 5666 3927
rect 5663 3858 5667 3859
rect 5663 3853 5667 3854
rect 5618 3843 5624 3844
rect 5618 3839 5619 3843
rect 5623 3839 5624 3843
rect 5618 3838 5624 3839
rect 5664 3793 5666 3853
rect 5662 3792 5668 3793
rect 5514 3791 5520 3792
rect 5514 3787 5515 3791
rect 5519 3787 5520 3791
rect 5662 3788 5663 3792
rect 5667 3788 5668 3792
rect 5662 3787 5668 3788
rect 5514 3786 5520 3787
rect 5542 3776 5548 3777
rect 5350 3772 5351 3776
rect 5355 3772 5356 3776
rect 5350 3771 5356 3772
rect 5446 3775 5452 3776
rect 5446 3771 5447 3775
rect 5451 3771 5452 3775
rect 5542 3772 5543 3776
rect 5547 3772 5548 3776
rect 5542 3771 5548 3772
rect 5662 3775 5668 3776
rect 5662 3771 5663 3775
rect 5667 3771 5668 3775
rect 3838 3770 3844 3771
rect 3495 3754 3499 3755
rect 3495 3749 3499 3750
rect 3591 3754 3595 3755
rect 3591 3749 3595 3750
rect 3679 3754 3683 3755
rect 3679 3749 3683 3750
rect 3799 3754 3803 3755
rect 3799 3749 3803 3750
rect 3496 3725 3498 3749
rect 3680 3725 3682 3749
rect 3800 3726 3802 3749
rect 3798 3725 3804 3726
rect 3494 3724 3500 3725
rect 3678 3724 3684 3725
rect 2646 3720 2647 3724
rect 2651 3720 2652 3724
rect 2646 3719 2652 3720
rect 2742 3723 2748 3724
rect 2742 3719 2743 3723
rect 2747 3719 2748 3723
rect 2870 3720 2871 3724
rect 2875 3720 2876 3724
rect 2870 3719 2876 3720
rect 2970 3723 2976 3724
rect 2970 3719 2971 3723
rect 2975 3719 2976 3723
rect 3086 3720 3087 3724
rect 3091 3720 3092 3724
rect 3086 3719 3092 3720
rect 3186 3723 3192 3724
rect 3186 3719 3187 3723
rect 3191 3719 3192 3723
rect 3294 3720 3295 3724
rect 3299 3720 3300 3724
rect 3294 3719 3300 3720
rect 3390 3723 3396 3724
rect 3390 3719 3391 3723
rect 3395 3719 3396 3723
rect 3494 3720 3495 3724
rect 3499 3720 3500 3724
rect 3494 3719 3500 3720
rect 3590 3723 3596 3724
rect 3590 3719 3591 3723
rect 3595 3719 3596 3723
rect 3678 3720 3679 3724
rect 3683 3720 3684 3724
rect 3678 3719 3684 3720
rect 3770 3723 3776 3724
rect 3770 3719 3771 3723
rect 3775 3719 3776 3723
rect 3798 3721 3799 3725
rect 3803 3721 3804 3725
rect 3798 3720 3804 3721
rect 3840 3719 3842 3770
rect 4080 3719 4082 3771
rect 4170 3770 4176 3771
rect 2742 3718 2748 3719
rect 2970 3718 2976 3719
rect 3186 3718 3192 3719
rect 3390 3718 3396 3719
rect 3590 3718 3596 3719
rect 3770 3718 3776 3719
rect 3839 3718 3843 3719
rect 2638 3659 2644 3660
rect 2638 3655 2639 3659
rect 2643 3655 2644 3659
rect 2638 3654 2644 3655
rect 2744 3652 2746 3718
rect 2842 3709 2848 3710
rect 2842 3705 2843 3709
rect 2847 3705 2848 3709
rect 2842 3704 2848 3705
rect 2742 3651 2748 3652
rect 2742 3647 2743 3651
rect 2747 3647 2748 3651
rect 2742 3646 2748 3647
rect 2844 3635 2846 3704
rect 2938 3687 2944 3688
rect 2938 3683 2939 3687
rect 2943 3683 2944 3687
rect 2938 3682 2944 3683
rect 2940 3660 2942 3682
rect 2972 3660 2974 3718
rect 3058 3709 3064 3710
rect 3058 3705 3059 3709
rect 3063 3705 3064 3709
rect 3058 3704 3064 3705
rect 2938 3659 2944 3660
rect 2938 3655 2939 3659
rect 2943 3655 2944 3659
rect 2938 3654 2944 3655
rect 2970 3659 2976 3660
rect 2970 3655 2971 3659
rect 2975 3655 2976 3659
rect 2970 3654 2976 3655
rect 3060 3635 3062 3704
rect 3188 3660 3190 3718
rect 3266 3709 3272 3710
rect 3266 3705 3267 3709
rect 3271 3705 3272 3709
rect 3266 3704 3272 3705
rect 3466 3709 3472 3710
rect 3466 3705 3467 3709
rect 3471 3705 3472 3709
rect 3466 3704 3472 3705
rect 3186 3659 3192 3660
rect 3186 3655 3187 3659
rect 3191 3655 3192 3659
rect 3186 3654 3192 3655
rect 3268 3635 3270 3704
rect 3468 3635 3470 3704
rect 3592 3688 3594 3718
rect 3650 3709 3656 3710
rect 3650 3705 3651 3709
rect 3655 3705 3656 3709
rect 3650 3704 3656 3705
rect 3590 3687 3596 3688
rect 3590 3683 3591 3687
rect 3595 3683 3596 3687
rect 3590 3682 3596 3683
rect 3652 3635 3654 3704
rect 3772 3652 3774 3718
rect 3839 3713 3843 3714
rect 3887 3718 3891 3719
rect 3887 3713 3891 3714
rect 4055 3718 4059 3719
rect 4055 3713 4059 3714
rect 4079 3718 4083 3719
rect 4079 3713 4083 3714
rect 3798 3708 3804 3709
rect 3798 3704 3799 3708
rect 3803 3704 3804 3708
rect 3798 3703 3804 3704
rect 3770 3651 3776 3652
rect 3770 3647 3771 3651
rect 3775 3647 3776 3651
rect 3770 3646 3776 3647
rect 3800 3635 3802 3703
rect 3840 3690 3842 3713
rect 3838 3689 3844 3690
rect 3888 3689 3890 3713
rect 4056 3689 4058 3713
rect 3838 3685 3839 3689
rect 3843 3685 3844 3689
rect 3838 3684 3844 3685
rect 3886 3688 3892 3689
rect 4054 3688 4060 3689
rect 3886 3684 3887 3688
rect 3891 3684 3892 3688
rect 3886 3683 3892 3684
rect 3982 3687 3988 3688
rect 3982 3683 3983 3687
rect 3987 3683 3988 3687
rect 4054 3684 4055 3688
rect 4059 3684 4060 3688
rect 4054 3683 4060 3684
rect 3982 3682 3988 3683
rect 3858 3673 3864 3674
rect 3838 3672 3844 3673
rect 3838 3668 3839 3672
rect 3843 3668 3844 3672
rect 3858 3669 3859 3673
rect 3863 3669 3864 3673
rect 3858 3668 3864 3669
rect 3838 3667 3844 3668
rect 2547 3634 2551 3635
rect 2547 3629 2551 3630
rect 2619 3634 2623 3635
rect 2619 3629 2623 3630
rect 2683 3634 2687 3635
rect 2683 3629 2687 3630
rect 2843 3634 2847 3635
rect 2843 3629 2847 3630
rect 3059 3634 3063 3635
rect 3059 3629 3063 3630
rect 3267 3634 3271 3635
rect 3267 3629 3271 3630
rect 3467 3634 3471 3635
rect 3467 3629 3471 3630
rect 3651 3634 3655 3635
rect 3651 3629 3655 3630
rect 3799 3634 3803 3635
rect 3799 3629 3803 3630
rect 2502 3619 2508 3620
rect 2502 3615 2503 3619
rect 2507 3615 2508 3619
rect 2502 3614 2508 3615
rect 2548 3568 2550 3629
rect 2554 3615 2560 3616
rect 2554 3611 2555 3615
rect 2559 3611 2560 3615
rect 2554 3610 2560 3611
rect 1974 3564 1975 3568
rect 1979 3564 1980 3568
rect 1974 3563 1980 3564
rect 2410 3567 2416 3568
rect 2410 3563 2411 3567
rect 2415 3563 2416 3567
rect 2410 3562 2416 3563
rect 2546 3567 2552 3568
rect 2546 3563 2547 3567
rect 2551 3563 2552 3567
rect 2546 3562 2552 3563
rect 2438 3552 2444 3553
rect 2556 3552 2558 3610
rect 2684 3568 2686 3629
rect 2690 3615 2696 3616
rect 2690 3611 2691 3615
rect 2695 3611 2696 3615
rect 2690 3610 2696 3611
rect 2682 3567 2688 3568
rect 2682 3563 2683 3567
rect 2687 3563 2688 3567
rect 2682 3562 2688 3563
rect 2574 3552 2580 3553
rect 2692 3552 2694 3610
rect 3778 3591 3784 3592
rect 3778 3587 3779 3591
rect 3783 3587 3784 3591
rect 3778 3586 3784 3587
rect 2710 3552 2716 3553
rect 1974 3551 1980 3552
rect 1974 3547 1975 3551
rect 1979 3547 1980 3551
rect 2438 3548 2439 3552
rect 2443 3548 2444 3552
rect 2438 3547 2444 3548
rect 2554 3551 2560 3552
rect 2554 3547 2555 3551
rect 2559 3547 2560 3551
rect 2574 3548 2575 3552
rect 2579 3548 2580 3552
rect 2574 3547 2580 3548
rect 2690 3551 2696 3552
rect 2690 3547 2691 3551
rect 2695 3547 2696 3551
rect 2710 3548 2711 3552
rect 2715 3548 2716 3552
rect 2710 3547 2716 3548
rect 2806 3551 2812 3552
rect 2806 3547 2807 3551
rect 2811 3547 2812 3551
rect 1974 3546 1980 3547
rect 1934 3532 1940 3533
rect 1934 3528 1935 3532
rect 1939 3528 1940 3532
rect 1934 3527 1940 3528
rect 1446 3515 1452 3516
rect 1446 3511 1447 3515
rect 1451 3511 1452 3515
rect 1486 3512 1487 3516
rect 1491 3512 1492 3516
rect 1486 3511 1492 3512
rect 1602 3515 1608 3516
rect 1602 3511 1603 3515
rect 1607 3511 1608 3515
rect 1622 3512 1623 3516
rect 1627 3512 1628 3516
rect 1622 3511 1628 3512
rect 1738 3515 1744 3516
rect 1738 3511 1739 3515
rect 1743 3511 1744 3515
rect 1758 3512 1759 3516
rect 1763 3512 1764 3516
rect 1758 3511 1764 3512
rect 1850 3515 1856 3516
rect 1850 3511 1851 3515
rect 1855 3511 1856 3515
rect 1446 3510 1452 3511
rect 1407 3462 1411 3463
rect 1407 3457 1411 3458
rect 1408 3433 1410 3457
rect 1406 3432 1412 3433
rect 1134 3428 1135 3432
rect 1139 3428 1140 3432
rect 1134 3427 1140 3428
rect 1234 3431 1240 3432
rect 1234 3427 1235 3431
rect 1239 3427 1240 3431
rect 1270 3428 1271 3432
rect 1275 3428 1276 3432
rect 1270 3427 1276 3428
rect 1370 3431 1376 3432
rect 1370 3427 1371 3431
rect 1375 3427 1376 3431
rect 1406 3428 1407 3432
rect 1411 3428 1412 3432
rect 1406 3427 1412 3428
rect 826 3426 832 3427
rect 962 3426 968 3427
rect 1234 3426 1240 3427
rect 1370 3426 1376 3427
rect 698 3417 704 3418
rect 110 3416 116 3417
rect 110 3412 111 3416
rect 115 3412 116 3416
rect 698 3413 699 3417
rect 703 3413 704 3417
rect 698 3412 704 3413
rect 110 3411 116 3412
rect 112 3347 114 3411
rect 700 3347 702 3412
rect 828 3368 830 3426
rect 834 3417 840 3418
rect 834 3413 835 3417
rect 839 3413 840 3417
rect 834 3412 840 3413
rect 826 3367 832 3368
rect 826 3363 827 3367
rect 831 3363 832 3367
rect 826 3362 832 3363
rect 836 3347 838 3412
rect 964 3368 966 3426
rect 970 3417 976 3418
rect 970 3413 971 3417
rect 975 3413 976 3417
rect 970 3412 976 3413
rect 1106 3417 1112 3418
rect 1106 3413 1107 3417
rect 1111 3413 1112 3417
rect 1106 3412 1112 3413
rect 962 3367 968 3368
rect 962 3363 963 3367
rect 967 3363 968 3367
rect 962 3362 968 3363
rect 874 3359 880 3360
rect 874 3355 875 3359
rect 879 3355 880 3359
rect 874 3354 880 3355
rect 111 3346 115 3347
rect 111 3341 115 3342
rect 699 3346 703 3347
rect 699 3341 703 3342
rect 755 3346 759 3347
rect 755 3341 759 3342
rect 835 3346 839 3347
rect 835 3341 839 3342
rect 112 3281 114 3341
rect 110 3280 116 3281
rect 756 3280 758 3341
rect 110 3276 111 3280
rect 115 3276 116 3280
rect 110 3275 116 3276
rect 754 3279 760 3280
rect 754 3275 755 3279
rect 759 3275 760 3279
rect 754 3274 760 3275
rect 782 3264 788 3265
rect 876 3264 878 3354
rect 972 3347 974 3412
rect 1108 3347 1110 3412
rect 1236 3368 1238 3426
rect 1242 3417 1248 3418
rect 1242 3413 1243 3417
rect 1247 3413 1248 3417
rect 1242 3412 1248 3413
rect 1378 3417 1384 3418
rect 1378 3413 1379 3417
rect 1383 3413 1384 3417
rect 1378 3412 1384 3413
rect 1234 3367 1240 3368
rect 1234 3363 1235 3367
rect 1239 3363 1240 3367
rect 1234 3362 1240 3363
rect 1244 3347 1246 3412
rect 1380 3347 1382 3412
rect 1448 3368 1450 3510
rect 1488 3463 1490 3511
rect 1602 3510 1608 3511
rect 1624 3463 1626 3511
rect 1738 3510 1744 3511
rect 1760 3463 1762 3511
rect 1850 3510 1856 3511
rect 1934 3515 1940 3516
rect 1934 3511 1935 3515
rect 1939 3511 1940 3515
rect 1934 3510 1940 3511
rect 1936 3463 1938 3510
rect 1976 3483 1978 3546
rect 2440 3483 2442 3547
rect 2554 3546 2560 3547
rect 2576 3483 2578 3547
rect 2690 3546 2696 3547
rect 2712 3483 2714 3547
rect 2806 3546 2812 3547
rect 1975 3482 1979 3483
rect 1975 3477 1979 3478
rect 2439 3482 2443 3483
rect 2439 3477 2443 3478
rect 2575 3482 2579 3483
rect 2575 3477 2579 3478
rect 2599 3482 2603 3483
rect 2599 3477 2603 3478
rect 2711 3482 2715 3483
rect 2711 3477 2715 3478
rect 1487 3462 1491 3463
rect 1487 3457 1491 3458
rect 1543 3462 1547 3463
rect 1543 3457 1547 3458
rect 1623 3462 1627 3463
rect 1623 3457 1627 3458
rect 1679 3462 1683 3463
rect 1679 3457 1683 3458
rect 1759 3462 1763 3463
rect 1759 3457 1763 3458
rect 1815 3462 1819 3463
rect 1815 3457 1819 3458
rect 1935 3462 1939 3463
rect 1935 3457 1939 3458
rect 1544 3433 1546 3457
rect 1680 3433 1682 3457
rect 1816 3433 1818 3457
rect 1936 3434 1938 3457
rect 1976 3454 1978 3477
rect 1974 3453 1980 3454
rect 2600 3453 2602 3477
rect 1974 3449 1975 3453
rect 1979 3449 1980 3453
rect 1974 3448 1980 3449
rect 2598 3452 2604 3453
rect 2598 3448 2599 3452
rect 2603 3448 2604 3452
rect 2598 3447 2604 3448
rect 2698 3451 2704 3452
rect 2698 3447 2699 3451
rect 2703 3447 2704 3451
rect 2698 3446 2704 3447
rect 2570 3437 2576 3438
rect 1974 3436 1980 3437
rect 1934 3433 1940 3434
rect 1542 3432 1548 3433
rect 1678 3432 1684 3433
rect 1814 3432 1820 3433
rect 1506 3431 1512 3432
rect 1506 3427 1507 3431
rect 1511 3427 1512 3431
rect 1542 3428 1543 3432
rect 1547 3428 1548 3432
rect 1542 3427 1548 3428
rect 1642 3431 1648 3432
rect 1642 3427 1643 3431
rect 1647 3427 1648 3431
rect 1678 3428 1679 3432
rect 1683 3428 1684 3432
rect 1678 3427 1684 3428
rect 1778 3431 1784 3432
rect 1778 3427 1779 3431
rect 1783 3427 1784 3431
rect 1814 3428 1815 3432
rect 1819 3428 1820 3432
rect 1814 3427 1820 3428
rect 1906 3431 1912 3432
rect 1906 3427 1907 3431
rect 1911 3427 1912 3431
rect 1934 3429 1935 3433
rect 1939 3429 1940 3433
rect 1974 3432 1975 3436
rect 1979 3432 1980 3436
rect 2570 3433 2571 3437
rect 2575 3433 2576 3437
rect 2570 3432 2576 3433
rect 1974 3431 1980 3432
rect 1934 3428 1940 3429
rect 1506 3426 1512 3427
rect 1642 3426 1648 3427
rect 1778 3426 1784 3427
rect 1906 3426 1912 3427
rect 1508 3368 1510 3426
rect 1514 3417 1520 3418
rect 1514 3413 1515 3417
rect 1519 3413 1520 3417
rect 1514 3412 1520 3413
rect 1446 3367 1452 3368
rect 1446 3363 1447 3367
rect 1451 3363 1452 3367
rect 1446 3362 1452 3363
rect 1506 3367 1512 3368
rect 1506 3363 1507 3367
rect 1511 3363 1512 3367
rect 1506 3362 1512 3363
rect 1516 3347 1518 3412
rect 1644 3368 1646 3426
rect 1650 3417 1656 3418
rect 1650 3413 1651 3417
rect 1655 3413 1656 3417
rect 1650 3412 1656 3413
rect 1642 3367 1648 3368
rect 1642 3363 1643 3367
rect 1647 3363 1648 3367
rect 1642 3362 1648 3363
rect 1652 3347 1654 3412
rect 1780 3368 1782 3426
rect 1786 3417 1792 3418
rect 1786 3413 1787 3417
rect 1791 3413 1792 3417
rect 1786 3412 1792 3413
rect 1778 3367 1784 3368
rect 1778 3363 1779 3367
rect 1783 3363 1784 3367
rect 1778 3362 1784 3363
rect 1788 3347 1790 3412
rect 891 3346 895 3347
rect 891 3341 895 3342
rect 971 3346 975 3347
rect 971 3341 975 3342
rect 1035 3346 1039 3347
rect 1035 3341 1039 3342
rect 1107 3346 1111 3347
rect 1107 3341 1111 3342
rect 1187 3346 1191 3347
rect 1187 3341 1191 3342
rect 1243 3346 1247 3347
rect 1243 3341 1247 3342
rect 1339 3346 1343 3347
rect 1339 3341 1343 3342
rect 1379 3346 1383 3347
rect 1379 3341 1383 3342
rect 1491 3346 1495 3347
rect 1491 3341 1495 3342
rect 1515 3346 1519 3347
rect 1515 3341 1519 3342
rect 1651 3346 1655 3347
rect 1651 3341 1655 3342
rect 1787 3346 1791 3347
rect 1787 3341 1791 3342
rect 892 3280 894 3341
rect 1018 3331 1024 3332
rect 1018 3327 1019 3331
rect 1023 3327 1024 3331
rect 1018 3326 1024 3327
rect 890 3279 896 3280
rect 890 3275 891 3279
rect 895 3275 896 3279
rect 890 3274 896 3275
rect 1020 3272 1022 3326
rect 1036 3280 1038 3341
rect 1158 3339 1164 3340
rect 1158 3335 1159 3339
rect 1163 3335 1164 3339
rect 1158 3334 1164 3335
rect 1130 3327 1136 3328
rect 1130 3323 1131 3327
rect 1135 3323 1136 3327
rect 1130 3322 1136 3323
rect 1034 3279 1040 3280
rect 1034 3275 1035 3279
rect 1039 3275 1040 3279
rect 1034 3274 1040 3275
rect 1018 3271 1024 3272
rect 1018 3267 1019 3271
rect 1023 3267 1024 3271
rect 1018 3266 1024 3267
rect 918 3264 924 3265
rect 1062 3264 1068 3265
rect 110 3263 116 3264
rect 110 3259 111 3263
rect 115 3259 116 3263
rect 782 3260 783 3264
rect 787 3260 788 3264
rect 782 3259 788 3260
rect 874 3263 880 3264
rect 874 3259 875 3263
rect 879 3259 880 3263
rect 918 3260 919 3264
rect 923 3260 924 3264
rect 918 3259 924 3260
rect 1010 3263 1016 3264
rect 1010 3259 1011 3263
rect 1015 3259 1016 3263
rect 1062 3260 1063 3264
rect 1067 3260 1068 3264
rect 1062 3259 1068 3260
rect 110 3258 116 3259
rect 112 3235 114 3258
rect 784 3235 786 3259
rect 874 3258 880 3259
rect 920 3235 922 3259
rect 1010 3258 1016 3259
rect 111 3234 115 3235
rect 111 3229 115 3230
rect 391 3234 395 3235
rect 391 3229 395 3230
rect 647 3234 651 3235
rect 647 3229 651 3230
rect 783 3234 787 3235
rect 783 3229 787 3230
rect 919 3234 923 3235
rect 919 3229 923 3230
rect 927 3234 931 3235
rect 927 3229 931 3230
rect 112 3206 114 3229
rect 110 3205 116 3206
rect 392 3205 394 3229
rect 648 3205 650 3229
rect 928 3205 930 3229
rect 110 3201 111 3205
rect 115 3201 116 3205
rect 110 3200 116 3201
rect 390 3204 396 3205
rect 646 3204 652 3205
rect 926 3204 932 3205
rect 390 3200 391 3204
rect 395 3200 396 3204
rect 390 3199 396 3200
rect 490 3203 496 3204
rect 490 3199 491 3203
rect 495 3199 496 3203
rect 646 3200 647 3204
rect 651 3200 652 3204
rect 646 3199 652 3200
rect 742 3203 748 3204
rect 742 3199 743 3203
rect 747 3199 748 3203
rect 926 3200 927 3204
rect 931 3200 932 3204
rect 926 3199 932 3200
rect 490 3198 496 3199
rect 742 3198 748 3199
rect 362 3189 368 3190
rect 110 3188 116 3189
rect 110 3184 111 3188
rect 115 3184 116 3188
rect 362 3185 363 3189
rect 367 3185 368 3189
rect 362 3184 368 3185
rect 110 3183 116 3184
rect 112 3111 114 3183
rect 364 3111 366 3184
rect 111 3110 115 3111
rect 111 3105 115 3106
rect 131 3110 135 3111
rect 131 3105 135 3106
rect 307 3110 311 3111
rect 307 3105 311 3106
rect 363 3110 367 3111
rect 363 3105 367 3106
rect 112 3045 114 3105
rect 110 3044 116 3045
rect 132 3044 134 3105
rect 308 3044 310 3105
rect 430 3099 436 3100
rect 430 3095 431 3099
rect 435 3095 436 3099
rect 492 3096 494 3198
rect 618 3189 624 3190
rect 618 3185 619 3189
rect 623 3185 624 3189
rect 618 3184 624 3185
rect 620 3111 622 3184
rect 744 3132 746 3198
rect 898 3189 904 3190
rect 898 3185 899 3189
rect 903 3185 904 3189
rect 898 3184 904 3185
rect 742 3131 748 3132
rect 742 3127 743 3131
rect 747 3127 748 3131
rect 742 3126 748 3127
rect 900 3111 902 3184
rect 1012 3140 1014 3258
rect 1064 3235 1066 3259
rect 1063 3234 1067 3235
rect 1063 3229 1067 3230
rect 1132 3220 1134 3322
rect 1160 3264 1162 3334
rect 1188 3280 1190 3341
rect 1340 3280 1342 3341
rect 1462 3335 1468 3336
rect 1462 3331 1463 3335
rect 1467 3331 1468 3335
rect 1462 3330 1468 3331
rect 1434 3327 1440 3328
rect 1434 3323 1435 3327
rect 1439 3323 1440 3327
rect 1434 3322 1440 3323
rect 1186 3279 1192 3280
rect 1186 3275 1187 3279
rect 1191 3275 1192 3279
rect 1186 3274 1192 3275
rect 1338 3279 1344 3280
rect 1338 3275 1339 3279
rect 1343 3275 1344 3279
rect 1338 3274 1344 3275
rect 1214 3264 1220 3265
rect 1158 3263 1164 3264
rect 1158 3259 1159 3263
rect 1163 3259 1164 3263
rect 1214 3260 1215 3264
rect 1219 3260 1220 3264
rect 1214 3259 1220 3260
rect 1366 3264 1372 3265
rect 1366 3260 1367 3264
rect 1371 3260 1372 3264
rect 1366 3259 1372 3260
rect 1158 3258 1164 3259
rect 1216 3235 1218 3259
rect 1368 3235 1370 3259
rect 1215 3234 1219 3235
rect 1215 3229 1219 3230
rect 1223 3234 1227 3235
rect 1223 3229 1227 3230
rect 1367 3234 1371 3235
rect 1367 3229 1371 3230
rect 1130 3219 1136 3220
rect 1130 3215 1131 3219
rect 1135 3215 1136 3219
rect 1130 3214 1136 3215
rect 1224 3205 1226 3229
rect 1436 3220 1438 3322
rect 1464 3264 1466 3330
rect 1492 3280 1494 3341
rect 1652 3280 1654 3341
rect 1658 3327 1664 3328
rect 1658 3323 1659 3327
rect 1663 3323 1664 3327
rect 1658 3322 1664 3323
rect 1490 3279 1496 3280
rect 1490 3275 1491 3279
rect 1495 3275 1496 3279
rect 1490 3274 1496 3275
rect 1650 3279 1656 3280
rect 1650 3275 1651 3279
rect 1655 3275 1656 3279
rect 1650 3274 1656 3275
rect 1518 3264 1524 3265
rect 1660 3264 1662 3322
rect 1788 3280 1790 3341
rect 1908 3336 1910 3426
rect 1934 3416 1940 3417
rect 1934 3412 1935 3416
rect 1939 3412 1940 3416
rect 1934 3411 1940 3412
rect 1936 3347 1938 3411
rect 1976 3363 1978 3431
rect 2572 3363 2574 3432
rect 1975 3362 1979 3363
rect 1975 3357 1979 3358
rect 2531 3362 2535 3363
rect 2531 3357 2535 3358
rect 2571 3362 2575 3363
rect 2571 3357 2575 3358
rect 1935 3346 1939 3347
rect 1935 3341 1939 3342
rect 1906 3335 1912 3336
rect 1906 3331 1907 3335
rect 1911 3331 1912 3335
rect 1906 3330 1912 3331
rect 1794 3327 1800 3328
rect 1794 3323 1795 3327
rect 1799 3323 1800 3327
rect 1794 3322 1800 3323
rect 1786 3279 1792 3280
rect 1786 3275 1787 3279
rect 1791 3275 1792 3279
rect 1786 3274 1792 3275
rect 1678 3264 1684 3265
rect 1796 3264 1798 3322
rect 1936 3281 1938 3341
rect 1976 3297 1978 3357
rect 1974 3296 1980 3297
rect 2532 3296 2534 3357
rect 2700 3348 2702 3446
rect 2794 3437 2800 3438
rect 2794 3433 2795 3437
rect 2799 3433 2800 3437
rect 2794 3432 2800 3433
rect 2796 3363 2798 3432
rect 2808 3388 2810 3546
rect 2823 3482 2827 3483
rect 2823 3477 2827 3478
rect 3047 3482 3051 3483
rect 3047 3477 3051 3478
rect 3263 3482 3267 3483
rect 3263 3477 3267 3478
rect 3479 3482 3483 3483
rect 3479 3477 3483 3478
rect 3679 3482 3683 3483
rect 3679 3477 3683 3478
rect 2824 3453 2826 3477
rect 3048 3453 3050 3477
rect 3264 3453 3266 3477
rect 3480 3453 3482 3477
rect 3680 3453 3682 3477
rect 2822 3452 2828 3453
rect 3046 3452 3052 3453
rect 3262 3452 3268 3453
rect 3478 3452 3484 3453
rect 3678 3452 3684 3453
rect 3780 3452 3782 3586
rect 3800 3569 3802 3629
rect 3840 3607 3842 3667
rect 3860 3607 3862 3668
rect 3984 3660 3986 3682
rect 4026 3673 4032 3674
rect 4026 3669 4027 3673
rect 4031 3669 4032 3673
rect 4026 3668 4032 3669
rect 3982 3659 3988 3660
rect 3982 3655 3983 3659
rect 3987 3655 3988 3659
rect 3982 3654 3988 3655
rect 3954 3623 3960 3624
rect 3954 3619 3955 3623
rect 3959 3619 3960 3623
rect 3954 3618 3960 3619
rect 3839 3606 3843 3607
rect 3839 3601 3843 3602
rect 3859 3606 3863 3607
rect 3859 3601 3863 3602
rect 3798 3568 3804 3569
rect 3798 3564 3799 3568
rect 3803 3564 3804 3568
rect 3798 3563 3804 3564
rect 3798 3551 3804 3552
rect 3798 3547 3799 3551
rect 3803 3547 3804 3551
rect 3798 3546 3804 3547
rect 3800 3483 3802 3546
rect 3840 3541 3842 3601
rect 3838 3540 3844 3541
rect 3860 3540 3862 3601
rect 3956 3597 3958 3618
rect 4028 3607 4030 3668
rect 4172 3624 4174 3770
rect 4296 3719 4298 3771
rect 4512 3719 4514 3771
rect 4728 3719 4730 3771
rect 4936 3719 4938 3771
rect 5034 3770 5040 3771
rect 5144 3719 5146 3771
rect 5352 3719 5354 3771
rect 5446 3770 5452 3771
rect 5544 3719 5546 3771
rect 5662 3770 5668 3771
rect 5664 3719 5666 3770
rect 4247 3718 4251 3719
rect 4247 3713 4251 3714
rect 4295 3718 4299 3719
rect 4295 3713 4299 3714
rect 4439 3718 4443 3719
rect 4439 3713 4443 3714
rect 4511 3718 4515 3719
rect 4511 3713 4515 3714
rect 4631 3718 4635 3719
rect 4631 3713 4635 3714
rect 4727 3718 4731 3719
rect 4727 3713 4731 3714
rect 4935 3718 4939 3719
rect 4935 3713 4939 3714
rect 5143 3718 5147 3719
rect 5143 3713 5147 3714
rect 5351 3718 5355 3719
rect 5351 3713 5355 3714
rect 5543 3718 5547 3719
rect 5543 3713 5547 3714
rect 5663 3718 5667 3719
rect 5663 3713 5667 3714
rect 4248 3689 4250 3713
rect 4440 3689 4442 3713
rect 4632 3689 4634 3713
rect 5664 3690 5666 3713
rect 5662 3689 5668 3690
rect 4246 3688 4252 3689
rect 4182 3687 4188 3688
rect 4182 3683 4183 3687
rect 4187 3683 4188 3687
rect 4246 3684 4247 3688
rect 4251 3684 4252 3688
rect 4246 3683 4252 3684
rect 4438 3688 4444 3689
rect 4630 3688 4636 3689
rect 4438 3684 4439 3688
rect 4443 3684 4444 3688
rect 4438 3683 4444 3684
rect 4566 3687 4572 3688
rect 4566 3683 4567 3687
rect 4571 3683 4572 3687
rect 4630 3684 4631 3688
rect 4635 3684 4636 3688
rect 4630 3683 4636 3684
rect 4722 3687 4728 3688
rect 4722 3683 4723 3687
rect 4727 3683 4728 3687
rect 5662 3685 5663 3689
rect 5667 3685 5668 3689
rect 5662 3684 5668 3685
rect 4182 3682 4188 3683
rect 4566 3682 4572 3683
rect 4722 3682 4728 3683
rect 4184 3624 4186 3682
rect 4218 3673 4224 3674
rect 4218 3669 4219 3673
rect 4223 3669 4224 3673
rect 4218 3668 4224 3669
rect 4410 3673 4416 3674
rect 4410 3669 4411 3673
rect 4415 3669 4416 3673
rect 4410 3668 4416 3669
rect 4170 3623 4176 3624
rect 4170 3619 4171 3623
rect 4175 3619 4176 3623
rect 4170 3618 4176 3619
rect 4182 3623 4188 3624
rect 4182 3619 4183 3623
rect 4187 3619 4188 3623
rect 4182 3618 4188 3619
rect 4220 3607 4222 3668
rect 4412 3607 4414 3668
rect 4568 3624 4570 3682
rect 4602 3673 4608 3674
rect 4602 3669 4603 3673
rect 4607 3669 4608 3673
rect 4602 3668 4608 3669
rect 4566 3623 4572 3624
rect 4566 3619 4567 3623
rect 4571 3619 4572 3623
rect 4566 3618 4572 3619
rect 4604 3607 4606 3668
rect 3995 3606 3999 3607
rect 3995 3601 3999 3602
rect 4027 3606 4031 3607
rect 4027 3601 4031 3602
rect 4131 3606 4135 3607
rect 4131 3601 4135 3602
rect 4219 3606 4223 3607
rect 4219 3601 4223 3602
rect 4267 3606 4271 3607
rect 4267 3601 4271 3602
rect 4403 3606 4407 3607
rect 4403 3601 4407 3602
rect 4411 3606 4415 3607
rect 4411 3601 4415 3602
rect 4539 3606 4543 3607
rect 4539 3601 4543 3602
rect 4603 3606 4607 3607
rect 4603 3601 4607 3602
rect 4675 3606 4679 3607
rect 4675 3601 4679 3602
rect 3955 3596 3959 3597
rect 3955 3591 3959 3592
rect 3996 3540 3998 3601
rect 4002 3587 4008 3588
rect 4002 3583 4003 3587
rect 4007 3583 4008 3587
rect 4002 3582 4008 3583
rect 3838 3536 3839 3540
rect 3843 3536 3844 3540
rect 3838 3535 3844 3536
rect 3858 3539 3864 3540
rect 3858 3535 3859 3539
rect 3863 3535 3864 3539
rect 3858 3534 3864 3535
rect 3994 3539 4000 3540
rect 3994 3535 3995 3539
rect 3999 3535 4000 3539
rect 3994 3534 4000 3535
rect 3886 3524 3892 3525
rect 4004 3524 4006 3582
rect 4132 3540 4134 3601
rect 4138 3587 4144 3588
rect 4138 3583 4139 3587
rect 4143 3583 4144 3587
rect 4138 3582 4144 3583
rect 4130 3539 4136 3540
rect 4130 3535 4131 3539
rect 4135 3535 4136 3539
rect 4130 3534 4136 3535
rect 4022 3524 4028 3525
rect 4140 3524 4142 3582
rect 4268 3540 4270 3601
rect 4274 3587 4280 3588
rect 4274 3583 4275 3587
rect 4279 3583 4280 3587
rect 4274 3582 4280 3583
rect 4266 3539 4272 3540
rect 4266 3535 4267 3539
rect 4271 3535 4272 3539
rect 4266 3534 4272 3535
rect 4158 3524 4164 3525
rect 4276 3524 4278 3582
rect 4404 3540 4406 3601
rect 4527 3596 4531 3597
rect 4527 3591 4531 3592
rect 4410 3587 4416 3588
rect 4410 3583 4411 3587
rect 4415 3583 4416 3587
rect 4410 3582 4416 3583
rect 4402 3539 4408 3540
rect 4402 3535 4403 3539
rect 4407 3535 4408 3539
rect 4402 3534 4408 3535
rect 4294 3524 4300 3525
rect 4412 3524 4414 3582
rect 4430 3524 4436 3525
rect 4528 3524 4530 3591
rect 4540 3540 4542 3601
rect 4676 3540 4678 3601
rect 4724 3600 4726 3682
rect 5662 3672 5668 3673
rect 5662 3668 5663 3672
rect 5667 3668 5668 3672
rect 5662 3667 5668 3668
rect 5664 3607 5666 3667
rect 4811 3606 4815 3607
rect 4811 3601 4815 3602
rect 4947 3606 4951 3607
rect 4947 3601 4951 3602
rect 5083 3606 5087 3607
rect 5083 3601 5087 3602
rect 5663 3606 5667 3607
rect 5663 3601 5667 3602
rect 4722 3599 4728 3600
rect 4722 3595 4723 3599
rect 4727 3595 4728 3599
rect 4722 3594 4728 3595
rect 4682 3587 4688 3588
rect 4682 3583 4683 3587
rect 4687 3583 4688 3587
rect 4682 3582 4688 3583
rect 4538 3539 4544 3540
rect 4538 3535 4539 3539
rect 4543 3535 4544 3539
rect 4538 3534 4544 3535
rect 4674 3539 4680 3540
rect 4674 3535 4675 3539
rect 4679 3535 4680 3539
rect 4674 3534 4680 3535
rect 4566 3524 4572 3525
rect 4684 3524 4686 3582
rect 4812 3540 4814 3601
rect 4818 3587 4824 3588
rect 4818 3583 4819 3587
rect 4823 3583 4824 3587
rect 4818 3582 4824 3583
rect 4810 3539 4816 3540
rect 4810 3535 4811 3539
rect 4815 3535 4816 3539
rect 4810 3534 4816 3535
rect 4702 3524 4708 3525
rect 4820 3524 4822 3582
rect 4948 3540 4950 3601
rect 4954 3587 4960 3588
rect 4954 3583 4955 3587
rect 4959 3583 4960 3587
rect 4954 3582 4960 3583
rect 4946 3539 4952 3540
rect 4946 3535 4947 3539
rect 4951 3535 4952 3539
rect 4946 3534 4952 3535
rect 4838 3524 4844 3525
rect 4956 3524 4958 3582
rect 5084 3540 5086 3601
rect 5090 3587 5096 3588
rect 5090 3583 5091 3587
rect 5095 3583 5096 3587
rect 5090 3582 5096 3583
rect 5082 3539 5088 3540
rect 5082 3535 5083 3539
rect 5087 3535 5088 3539
rect 5082 3534 5088 3535
rect 4974 3524 4980 3525
rect 5092 3524 5094 3582
rect 5664 3541 5666 3601
rect 5662 3540 5668 3541
rect 5662 3536 5663 3540
rect 5667 3536 5668 3540
rect 5662 3535 5668 3536
rect 5110 3524 5116 3525
rect 3838 3523 3844 3524
rect 3838 3519 3839 3523
rect 3843 3519 3844 3523
rect 3886 3520 3887 3524
rect 3891 3520 3892 3524
rect 3886 3519 3892 3520
rect 4002 3523 4008 3524
rect 4002 3519 4003 3523
rect 4007 3519 4008 3523
rect 4022 3520 4023 3524
rect 4027 3520 4028 3524
rect 4022 3519 4028 3520
rect 4138 3523 4144 3524
rect 4138 3519 4139 3523
rect 4143 3519 4144 3523
rect 4158 3520 4159 3524
rect 4163 3520 4164 3524
rect 4158 3519 4164 3520
rect 4274 3523 4280 3524
rect 4274 3519 4275 3523
rect 4279 3519 4280 3523
rect 4294 3520 4295 3524
rect 4299 3520 4300 3524
rect 4294 3519 4300 3520
rect 4410 3523 4416 3524
rect 4410 3519 4411 3523
rect 4415 3519 4416 3523
rect 4430 3520 4431 3524
rect 4435 3520 4436 3524
rect 4430 3519 4436 3520
rect 4526 3523 4532 3524
rect 4526 3519 4527 3523
rect 4531 3519 4532 3523
rect 4566 3520 4567 3524
rect 4571 3520 4572 3524
rect 4566 3519 4572 3520
rect 4682 3523 4688 3524
rect 4682 3519 4683 3523
rect 4687 3519 4688 3523
rect 4702 3520 4703 3524
rect 4707 3520 4708 3524
rect 4702 3519 4708 3520
rect 4818 3523 4824 3524
rect 4818 3519 4819 3523
rect 4823 3519 4824 3523
rect 4838 3520 4839 3524
rect 4843 3520 4844 3524
rect 4838 3519 4844 3520
rect 4954 3523 4960 3524
rect 4954 3519 4955 3523
rect 4959 3519 4960 3523
rect 4974 3520 4975 3524
rect 4979 3520 4980 3524
rect 4974 3519 4980 3520
rect 5090 3523 5096 3524
rect 5090 3519 5091 3523
rect 5095 3519 5096 3523
rect 5110 3520 5111 3524
rect 5115 3520 5116 3524
rect 5110 3519 5116 3520
rect 5206 3523 5212 3524
rect 5206 3519 5207 3523
rect 5211 3519 5212 3523
rect 3838 3518 3844 3519
rect 3840 3487 3842 3518
rect 3888 3487 3890 3519
rect 4002 3518 4008 3519
rect 4024 3487 4026 3519
rect 4138 3518 4144 3519
rect 4160 3487 4162 3519
rect 4274 3518 4280 3519
rect 4296 3487 4298 3519
rect 4410 3518 4416 3519
rect 4432 3487 4434 3519
rect 4526 3518 4532 3519
rect 4568 3487 4570 3519
rect 4682 3518 4688 3519
rect 4704 3487 4706 3519
rect 4818 3518 4824 3519
rect 4840 3487 4842 3519
rect 4954 3518 4960 3519
rect 4898 3487 4904 3488
rect 4976 3487 4978 3519
rect 5090 3518 5096 3519
rect 5112 3487 5114 3519
rect 5206 3518 5212 3519
rect 5662 3523 5668 3524
rect 5662 3519 5663 3523
rect 5667 3519 5668 3523
rect 5662 3518 5668 3519
rect 5208 3488 5210 3518
rect 5206 3487 5212 3488
rect 5664 3487 5666 3518
rect 3839 3486 3843 3487
rect 3799 3482 3803 3483
rect 3839 3481 3843 3482
rect 3887 3486 3891 3487
rect 3887 3481 3891 3482
rect 4023 3486 4027 3487
rect 4023 3481 4027 3482
rect 4159 3486 4163 3487
rect 4159 3481 4163 3482
rect 4295 3486 4299 3487
rect 4295 3481 4299 3482
rect 4431 3486 4435 3487
rect 4431 3481 4435 3482
rect 4567 3486 4571 3487
rect 4567 3481 4571 3482
rect 4703 3486 4707 3487
rect 4703 3481 4707 3482
rect 4831 3486 4835 3487
rect 4831 3481 4835 3482
rect 4839 3486 4843 3487
rect 4898 3483 4899 3487
rect 4903 3483 4904 3487
rect 4898 3482 4904 3483
rect 4967 3486 4971 3487
rect 4839 3481 4843 3482
rect 3799 3477 3803 3478
rect 3800 3454 3802 3477
rect 3840 3458 3842 3481
rect 3838 3457 3844 3458
rect 4832 3457 4834 3481
rect 3798 3453 3804 3454
rect 2822 3448 2823 3452
rect 2827 3448 2828 3452
rect 2822 3447 2828 3448
rect 2914 3451 2920 3452
rect 2914 3447 2915 3451
rect 2919 3447 2920 3451
rect 3046 3448 3047 3452
rect 3051 3448 3052 3452
rect 3046 3447 3052 3448
rect 3146 3451 3152 3452
rect 3146 3447 3147 3451
rect 3151 3447 3152 3451
rect 3262 3448 3263 3452
rect 3267 3448 3268 3452
rect 3262 3447 3268 3448
rect 3362 3451 3368 3452
rect 3362 3447 3363 3451
rect 3367 3447 3368 3451
rect 3478 3448 3479 3452
rect 3483 3448 3484 3452
rect 3478 3447 3484 3448
rect 3598 3451 3604 3452
rect 3598 3447 3599 3451
rect 3603 3447 3604 3451
rect 3678 3448 3679 3452
rect 3683 3448 3684 3452
rect 3678 3447 3684 3448
rect 3778 3451 3784 3452
rect 3778 3447 3779 3451
rect 3783 3447 3784 3451
rect 3798 3449 3799 3453
rect 3803 3449 3804 3453
rect 3838 3453 3839 3457
rect 3843 3453 3844 3457
rect 3838 3452 3844 3453
rect 4830 3456 4836 3457
rect 4830 3452 4831 3456
rect 4835 3452 4836 3456
rect 4830 3451 4836 3452
rect 3798 3448 3804 3449
rect 2914 3446 2920 3447
rect 3146 3446 3152 3447
rect 3362 3446 3368 3447
rect 3598 3446 3604 3447
rect 3778 3446 3784 3447
rect 2806 3387 2812 3388
rect 2806 3383 2807 3387
rect 2811 3383 2812 3387
rect 2806 3382 2812 3383
rect 2916 3380 2918 3446
rect 3018 3437 3024 3438
rect 3018 3433 3019 3437
rect 3023 3433 3024 3437
rect 3018 3432 3024 3433
rect 2914 3379 2920 3380
rect 2914 3375 2915 3379
rect 2919 3375 2920 3379
rect 2914 3374 2920 3375
rect 3020 3363 3022 3432
rect 3148 3388 3150 3446
rect 3234 3437 3240 3438
rect 3234 3433 3235 3437
rect 3239 3433 3240 3437
rect 3234 3432 3240 3433
rect 3114 3387 3120 3388
rect 3114 3383 3115 3387
rect 3119 3383 3120 3387
rect 3114 3382 3120 3383
rect 3146 3387 3152 3388
rect 3146 3383 3147 3387
rect 3151 3383 3152 3387
rect 3146 3382 3152 3383
rect 2715 3362 2719 3363
rect 2715 3357 2719 3358
rect 2795 3362 2799 3363
rect 2795 3357 2799 3358
rect 2899 3362 2903 3363
rect 2899 3357 2903 3358
rect 3019 3362 3023 3363
rect 3019 3357 3023 3358
rect 3083 3362 3087 3363
rect 3083 3357 3087 3358
rect 2698 3347 2704 3348
rect 2698 3343 2699 3347
rect 2703 3343 2704 3347
rect 2698 3342 2704 3343
rect 2716 3296 2718 3357
rect 2900 3296 2902 3357
rect 3070 3347 3076 3348
rect 3070 3343 3071 3347
rect 3075 3343 3076 3347
rect 3070 3342 3076 3343
rect 1974 3292 1975 3296
rect 1979 3292 1980 3296
rect 1974 3291 1980 3292
rect 2530 3295 2536 3296
rect 2530 3291 2531 3295
rect 2535 3291 2536 3295
rect 2530 3290 2536 3291
rect 2714 3295 2720 3296
rect 2714 3291 2715 3295
rect 2719 3291 2720 3295
rect 2714 3290 2720 3291
rect 2898 3295 2904 3296
rect 2898 3291 2899 3295
rect 2903 3291 2904 3295
rect 2898 3290 2904 3291
rect 1934 3280 1940 3281
rect 2558 3280 2564 3281
rect 2742 3280 2748 3281
rect 1934 3276 1935 3280
rect 1939 3276 1940 3280
rect 1934 3275 1940 3276
rect 1974 3279 1980 3280
rect 1974 3275 1975 3279
rect 1979 3275 1980 3279
rect 2558 3276 2559 3280
rect 2563 3276 2564 3280
rect 2558 3275 2564 3276
rect 2654 3279 2660 3280
rect 2654 3275 2655 3279
rect 2659 3275 2660 3279
rect 2742 3276 2743 3280
rect 2747 3276 2748 3280
rect 2742 3275 2748 3276
rect 2926 3280 2932 3281
rect 2926 3276 2927 3280
rect 2931 3276 2932 3280
rect 2926 3275 2932 3276
rect 1974 3274 1980 3275
rect 1814 3264 1820 3265
rect 1462 3263 1468 3264
rect 1462 3259 1463 3263
rect 1467 3259 1468 3263
rect 1518 3260 1519 3264
rect 1523 3260 1524 3264
rect 1518 3259 1524 3260
rect 1658 3263 1664 3264
rect 1658 3259 1659 3263
rect 1663 3259 1664 3263
rect 1678 3260 1679 3264
rect 1683 3260 1684 3264
rect 1678 3259 1684 3260
rect 1794 3263 1800 3264
rect 1794 3259 1795 3263
rect 1799 3259 1800 3263
rect 1814 3260 1815 3264
rect 1819 3260 1820 3264
rect 1814 3259 1820 3260
rect 1910 3263 1916 3264
rect 1910 3259 1911 3263
rect 1915 3259 1916 3263
rect 1462 3258 1468 3259
rect 1520 3235 1522 3259
rect 1658 3258 1664 3259
rect 1680 3235 1682 3259
rect 1794 3258 1800 3259
rect 1816 3235 1818 3259
rect 1910 3258 1916 3259
rect 1934 3263 1940 3264
rect 1934 3259 1935 3263
rect 1939 3259 1940 3263
rect 1934 3258 1940 3259
rect 1519 3234 1523 3235
rect 1519 3229 1523 3230
rect 1527 3234 1531 3235
rect 1527 3229 1531 3230
rect 1679 3234 1683 3235
rect 1679 3229 1683 3230
rect 1815 3234 1819 3235
rect 1815 3229 1819 3230
rect 1434 3219 1440 3220
rect 1434 3215 1435 3219
rect 1439 3215 1440 3219
rect 1434 3214 1440 3215
rect 1528 3205 1530 3229
rect 1816 3205 1818 3229
rect 1222 3204 1228 3205
rect 1018 3203 1024 3204
rect 1018 3199 1019 3203
rect 1023 3199 1024 3203
rect 1222 3200 1223 3204
rect 1227 3200 1228 3204
rect 1222 3199 1228 3200
rect 1526 3204 1532 3205
rect 1526 3200 1527 3204
rect 1531 3200 1532 3204
rect 1526 3199 1532 3200
rect 1814 3204 1820 3205
rect 1814 3200 1815 3204
rect 1819 3200 1820 3204
rect 1814 3199 1820 3200
rect 1018 3198 1024 3199
rect 1010 3139 1016 3140
rect 1010 3135 1011 3139
rect 1015 3135 1016 3139
rect 1010 3134 1016 3135
rect 1020 3132 1022 3198
rect 1194 3189 1200 3190
rect 1194 3185 1195 3189
rect 1199 3185 1200 3189
rect 1194 3184 1200 3185
rect 1498 3189 1504 3190
rect 1498 3185 1499 3189
rect 1503 3185 1504 3189
rect 1498 3184 1504 3185
rect 1786 3189 1792 3190
rect 1786 3185 1787 3189
rect 1791 3185 1792 3189
rect 1786 3184 1792 3185
rect 1026 3139 1032 3140
rect 1026 3135 1027 3139
rect 1031 3135 1032 3139
rect 1026 3134 1032 3135
rect 1018 3131 1024 3132
rect 1018 3127 1019 3131
rect 1023 3127 1024 3131
rect 1018 3126 1024 3127
rect 507 3110 511 3111
rect 507 3105 511 3106
rect 619 3110 623 3111
rect 619 3105 623 3106
rect 707 3110 711 3111
rect 707 3105 711 3106
rect 899 3110 903 3111
rect 899 3105 903 3106
rect 430 3094 436 3095
rect 490 3095 496 3096
rect 110 3040 111 3044
rect 115 3040 116 3044
rect 110 3039 116 3040
rect 130 3043 136 3044
rect 130 3039 131 3043
rect 135 3039 136 3043
rect 130 3038 136 3039
rect 306 3043 312 3044
rect 306 3039 307 3043
rect 311 3039 312 3043
rect 306 3038 312 3039
rect 158 3028 164 3029
rect 334 3028 340 3029
rect 432 3028 434 3094
rect 490 3091 491 3095
rect 495 3091 496 3095
rect 490 3090 496 3091
rect 498 3087 504 3088
rect 498 3083 499 3087
rect 503 3083 504 3087
rect 498 3082 504 3083
rect 500 3036 502 3082
rect 508 3044 510 3105
rect 708 3044 710 3105
rect 802 3091 808 3092
rect 802 3087 803 3091
rect 807 3087 808 3091
rect 802 3086 808 3087
rect 506 3043 512 3044
rect 506 3039 507 3043
rect 511 3039 512 3043
rect 506 3038 512 3039
rect 706 3043 712 3044
rect 706 3039 707 3043
rect 711 3039 712 3043
rect 706 3038 712 3039
rect 498 3035 504 3036
rect 498 3031 499 3035
rect 503 3031 504 3035
rect 498 3030 504 3031
rect 534 3028 540 3029
rect 110 3027 116 3028
rect 110 3023 111 3027
rect 115 3023 116 3027
rect 158 3024 159 3028
rect 163 3024 164 3028
rect 158 3023 164 3024
rect 250 3027 256 3028
rect 250 3023 251 3027
rect 255 3023 256 3027
rect 334 3024 335 3028
rect 339 3024 340 3028
rect 334 3023 340 3024
rect 430 3027 436 3028
rect 430 3023 431 3027
rect 435 3023 436 3027
rect 534 3024 535 3028
rect 539 3024 540 3028
rect 534 3023 540 3024
rect 734 3028 740 3029
rect 734 3024 735 3028
rect 739 3024 740 3028
rect 734 3023 740 3024
rect 110 3022 116 3023
rect 112 2995 114 3022
rect 160 2995 162 3023
rect 250 3022 256 3023
rect 111 2994 115 2995
rect 111 2989 115 2990
rect 159 2994 163 2995
rect 159 2989 163 2990
rect 112 2966 114 2989
rect 110 2965 116 2966
rect 160 2965 162 2989
rect 110 2961 111 2965
rect 115 2961 116 2965
rect 110 2960 116 2961
rect 158 2964 164 2965
rect 158 2960 159 2964
rect 163 2960 164 2964
rect 158 2959 164 2960
rect 130 2949 136 2950
rect 110 2948 116 2949
rect 110 2944 111 2948
rect 115 2944 116 2948
rect 130 2945 131 2949
rect 135 2945 136 2949
rect 130 2944 136 2945
rect 110 2943 116 2944
rect 112 2879 114 2943
rect 132 2879 134 2944
rect 252 2900 254 3022
rect 336 2995 338 3023
rect 430 3022 436 3023
rect 536 2995 538 3023
rect 736 2995 738 3023
rect 295 2994 299 2995
rect 295 2989 299 2990
rect 335 2994 339 2995
rect 335 2989 339 2990
rect 431 2994 435 2995
rect 431 2989 435 2990
rect 535 2994 539 2995
rect 535 2989 539 2990
rect 567 2994 571 2995
rect 567 2989 571 2990
rect 703 2994 707 2995
rect 703 2989 707 2990
rect 735 2994 739 2995
rect 735 2989 739 2990
rect 296 2965 298 2989
rect 432 2965 434 2989
rect 568 2965 570 2989
rect 704 2965 706 2989
rect 294 2964 300 2965
rect 430 2964 436 2965
rect 566 2964 572 2965
rect 702 2964 708 2965
rect 804 2964 806 3086
rect 900 3044 902 3105
rect 906 3091 912 3092
rect 906 3087 907 3091
rect 911 3087 912 3091
rect 906 3086 912 3087
rect 898 3043 904 3044
rect 898 3039 899 3043
rect 903 3039 904 3043
rect 898 3038 904 3039
rect 908 3028 910 3086
rect 926 3028 932 3029
rect 1028 3028 1030 3134
rect 1196 3111 1198 3184
rect 1500 3111 1502 3184
rect 1574 3139 1580 3140
rect 1574 3135 1575 3139
rect 1579 3135 1580 3139
rect 1574 3134 1580 3135
rect 1091 3110 1095 3111
rect 1091 3105 1095 3106
rect 1195 3110 1199 3111
rect 1195 3105 1199 3106
rect 1275 3110 1279 3111
rect 1275 3105 1279 3106
rect 1451 3110 1455 3111
rect 1451 3105 1455 3106
rect 1499 3110 1503 3111
rect 1499 3105 1503 3106
rect 1092 3044 1094 3105
rect 1266 3095 1272 3096
rect 1266 3091 1267 3095
rect 1271 3091 1272 3095
rect 1266 3090 1272 3091
rect 1090 3043 1096 3044
rect 1090 3039 1091 3043
rect 1095 3039 1096 3043
rect 1090 3038 1096 3039
rect 1268 3036 1270 3090
rect 1276 3044 1278 3105
rect 1282 3091 1288 3092
rect 1282 3087 1283 3091
rect 1287 3087 1288 3091
rect 1282 3086 1288 3087
rect 1274 3043 1280 3044
rect 1274 3039 1275 3043
rect 1279 3039 1280 3043
rect 1274 3038 1280 3039
rect 1266 3035 1272 3036
rect 1266 3031 1267 3035
rect 1271 3031 1272 3035
rect 1266 3030 1272 3031
rect 1118 3028 1124 3029
rect 1284 3028 1286 3086
rect 1452 3044 1454 3105
rect 1458 3091 1464 3092
rect 1458 3087 1459 3091
rect 1463 3087 1464 3091
rect 1458 3086 1464 3087
rect 1450 3043 1456 3044
rect 1450 3039 1451 3043
rect 1455 3039 1456 3043
rect 1450 3038 1456 3039
rect 1302 3028 1308 3029
rect 1460 3028 1462 3086
rect 1478 3028 1484 3029
rect 1576 3028 1578 3134
rect 1788 3111 1790 3184
rect 1912 3140 1914 3258
rect 1936 3235 1938 3258
rect 1976 3251 1978 3274
rect 2560 3251 2562 3275
rect 2654 3274 2660 3275
rect 1975 3250 1979 3251
rect 1975 3245 1979 3246
rect 2023 3250 2027 3251
rect 2023 3245 2027 3246
rect 2255 3250 2259 3251
rect 2255 3245 2259 3246
rect 2503 3250 2507 3251
rect 2503 3245 2507 3246
rect 2559 3250 2563 3251
rect 2559 3245 2563 3246
rect 1935 3234 1939 3235
rect 1935 3229 1939 3230
rect 1936 3206 1938 3229
rect 1976 3222 1978 3245
rect 1974 3221 1980 3222
rect 2024 3221 2026 3245
rect 2256 3221 2258 3245
rect 2504 3221 2506 3245
rect 1974 3217 1975 3221
rect 1979 3217 1980 3221
rect 1974 3216 1980 3217
rect 2022 3220 2028 3221
rect 2254 3220 2260 3221
rect 2502 3220 2508 3221
rect 2022 3216 2023 3220
rect 2027 3216 2028 3220
rect 2022 3215 2028 3216
rect 2142 3219 2148 3220
rect 2142 3215 2143 3219
rect 2147 3215 2148 3219
rect 2254 3216 2255 3220
rect 2259 3216 2260 3220
rect 2254 3215 2260 3216
rect 2346 3219 2352 3220
rect 2346 3215 2347 3219
rect 2351 3215 2352 3219
rect 2502 3216 2503 3220
rect 2507 3216 2508 3220
rect 2502 3215 2508 3216
rect 2594 3219 2600 3220
rect 2594 3215 2595 3219
rect 2599 3215 2600 3219
rect 2142 3214 2148 3215
rect 2346 3214 2352 3215
rect 2594 3214 2600 3215
rect 1934 3205 1940 3206
rect 1994 3205 2000 3206
rect 1926 3203 1932 3204
rect 1926 3199 1927 3203
rect 1931 3199 1932 3203
rect 1934 3201 1935 3205
rect 1939 3201 1940 3205
rect 1934 3200 1940 3201
rect 1974 3204 1980 3205
rect 1974 3200 1975 3204
rect 1979 3200 1980 3204
rect 1994 3201 1995 3205
rect 1999 3201 2000 3205
rect 1994 3200 2000 3201
rect 1974 3199 1980 3200
rect 1926 3198 1932 3199
rect 1928 3156 1930 3198
rect 1934 3188 1940 3189
rect 1934 3184 1935 3188
rect 1939 3184 1940 3188
rect 1934 3183 1940 3184
rect 1926 3155 1932 3156
rect 1926 3151 1927 3155
rect 1931 3151 1932 3155
rect 1926 3150 1932 3151
rect 1910 3139 1916 3140
rect 1910 3135 1911 3139
rect 1915 3135 1916 3139
rect 1910 3134 1916 3135
rect 1936 3111 1938 3183
rect 1976 3139 1978 3199
rect 1996 3139 1998 3200
rect 2144 3156 2146 3214
rect 2226 3205 2232 3206
rect 2226 3201 2227 3205
rect 2231 3201 2232 3205
rect 2226 3200 2232 3201
rect 2142 3155 2148 3156
rect 2142 3151 2143 3155
rect 2147 3151 2148 3155
rect 2142 3150 2148 3151
rect 2228 3139 2230 3200
rect 1975 3138 1979 3139
rect 1975 3133 1979 3134
rect 1995 3138 1999 3139
rect 1995 3133 1999 3134
rect 2227 3138 2231 3139
rect 2227 3133 2231 3134
rect 1627 3110 1631 3111
rect 1627 3105 1631 3106
rect 1787 3110 1791 3111
rect 1787 3105 1791 3106
rect 1935 3110 1939 3111
rect 1935 3105 1939 3106
rect 1628 3044 1630 3105
rect 1788 3044 1790 3105
rect 1936 3045 1938 3105
rect 1976 3073 1978 3133
rect 2348 3096 2350 3214
rect 2474 3205 2480 3206
rect 2474 3201 2475 3205
rect 2479 3201 2480 3205
rect 2474 3200 2480 3201
rect 2476 3139 2478 3200
rect 2475 3138 2479 3139
rect 2475 3133 2479 3134
rect 2483 3138 2487 3139
rect 2483 3133 2487 3134
rect 2346 3095 2352 3096
rect 2346 3091 2347 3095
rect 2351 3091 2352 3095
rect 2346 3090 2352 3091
rect 1974 3072 1980 3073
rect 2484 3072 2486 3133
rect 2596 3124 2598 3214
rect 2656 3156 2658 3274
rect 2744 3251 2746 3275
rect 2928 3251 2930 3275
rect 2743 3250 2747 3251
rect 2743 3245 2747 3246
rect 2927 3250 2931 3251
rect 2927 3245 2931 3246
rect 2975 3250 2979 3251
rect 2975 3245 2979 3246
rect 2744 3221 2746 3245
rect 2976 3221 2978 3245
rect 2742 3220 2748 3221
rect 2974 3220 2980 3221
rect 3072 3220 3074 3342
rect 3084 3296 3086 3357
rect 3090 3343 3096 3344
rect 3090 3339 3091 3343
rect 3095 3339 3096 3343
rect 3090 3338 3096 3339
rect 3082 3295 3088 3296
rect 3082 3291 3083 3295
rect 3087 3291 3088 3295
rect 3082 3290 3088 3291
rect 3092 3280 3094 3338
rect 3116 3304 3118 3382
rect 3236 3363 3238 3432
rect 3364 3388 3366 3446
rect 3450 3437 3456 3438
rect 3450 3433 3451 3437
rect 3455 3433 3456 3437
rect 3450 3432 3456 3433
rect 3362 3387 3368 3388
rect 3362 3383 3363 3387
rect 3367 3383 3368 3387
rect 3362 3382 3368 3383
rect 3452 3363 3454 3432
rect 3600 3388 3602 3446
rect 4802 3441 4808 3442
rect 3838 3440 3844 3441
rect 3650 3437 3656 3438
rect 3650 3433 3651 3437
rect 3655 3433 3656 3437
rect 3650 3432 3656 3433
rect 3798 3436 3804 3437
rect 3798 3432 3799 3436
rect 3803 3432 3804 3436
rect 3838 3436 3839 3440
rect 3843 3436 3844 3440
rect 4802 3437 4803 3441
rect 4807 3437 4808 3441
rect 4802 3436 4808 3437
rect 3838 3435 3844 3436
rect 3598 3387 3604 3388
rect 3598 3383 3599 3387
rect 3603 3383 3604 3387
rect 3598 3382 3604 3383
rect 3652 3363 3654 3432
rect 3798 3431 3804 3432
rect 3800 3363 3802 3431
rect 3840 3375 3842 3435
rect 4804 3375 4806 3436
rect 4900 3392 4902 3482
rect 4967 3481 4971 3482
rect 4975 3486 4979 3487
rect 4975 3481 4979 3482
rect 5103 3486 5107 3487
rect 5103 3481 5107 3482
rect 5111 3486 5115 3487
rect 5206 3483 5207 3487
rect 5211 3483 5212 3487
rect 5206 3482 5212 3483
rect 5239 3486 5243 3487
rect 5111 3481 5115 3482
rect 5239 3481 5243 3482
rect 5375 3486 5379 3487
rect 5375 3481 5379 3482
rect 5663 3486 5667 3487
rect 5663 3481 5667 3482
rect 4968 3457 4970 3481
rect 5104 3457 5106 3481
rect 5240 3457 5242 3481
rect 5376 3457 5378 3481
rect 5664 3458 5666 3481
rect 5662 3457 5668 3458
rect 4966 3456 4972 3457
rect 5102 3456 5108 3457
rect 5238 3456 5244 3457
rect 5374 3456 5380 3457
rect 4930 3455 4936 3456
rect 4930 3451 4931 3455
rect 4935 3451 4936 3455
rect 4966 3452 4967 3456
rect 4971 3452 4972 3456
rect 4966 3451 4972 3452
rect 5066 3455 5072 3456
rect 5066 3451 5067 3455
rect 5071 3451 5072 3455
rect 5102 3452 5103 3456
rect 5107 3452 5108 3456
rect 5102 3451 5108 3452
rect 5202 3455 5208 3456
rect 5202 3451 5203 3455
rect 5207 3451 5208 3455
rect 5238 3452 5239 3456
rect 5243 3452 5244 3456
rect 5238 3451 5244 3452
rect 5338 3455 5344 3456
rect 5338 3451 5339 3455
rect 5343 3451 5344 3455
rect 5374 3452 5375 3456
rect 5379 3452 5380 3456
rect 5374 3451 5380 3452
rect 5470 3455 5476 3456
rect 5470 3451 5471 3455
rect 5475 3451 5476 3455
rect 5662 3453 5663 3457
rect 5667 3453 5668 3457
rect 5662 3452 5668 3453
rect 4930 3450 4936 3451
rect 5066 3450 5072 3451
rect 5202 3450 5208 3451
rect 5338 3450 5344 3451
rect 5470 3450 5476 3451
rect 4932 3392 4934 3450
rect 4938 3441 4944 3442
rect 4938 3437 4939 3441
rect 4943 3437 4944 3441
rect 4938 3436 4944 3437
rect 4898 3391 4904 3392
rect 4898 3387 4899 3391
rect 4903 3387 4904 3391
rect 4898 3386 4904 3387
rect 4930 3391 4936 3392
rect 4930 3387 4931 3391
rect 4935 3387 4936 3391
rect 4930 3386 4936 3387
rect 4940 3375 4942 3436
rect 5068 3392 5070 3450
rect 5074 3441 5080 3442
rect 5074 3437 5075 3441
rect 5079 3437 5080 3441
rect 5074 3436 5080 3437
rect 5066 3391 5072 3392
rect 5066 3387 5067 3391
rect 5071 3387 5072 3391
rect 5066 3386 5072 3387
rect 5076 3375 5078 3436
rect 5204 3392 5206 3450
rect 5210 3441 5216 3442
rect 5210 3437 5211 3441
rect 5215 3437 5216 3441
rect 5210 3436 5216 3437
rect 5202 3391 5208 3392
rect 5202 3387 5203 3391
rect 5207 3387 5208 3391
rect 5202 3386 5208 3387
rect 5212 3375 5214 3436
rect 5340 3392 5342 3450
rect 5346 3441 5352 3442
rect 5346 3437 5347 3441
rect 5351 3437 5352 3441
rect 5346 3436 5352 3437
rect 5338 3391 5344 3392
rect 5338 3387 5339 3391
rect 5343 3387 5344 3391
rect 5338 3386 5344 3387
rect 5348 3375 5350 3436
rect 3839 3374 3843 3375
rect 3839 3369 3843 3370
rect 3859 3374 3863 3375
rect 3859 3369 3863 3370
rect 4139 3374 4143 3375
rect 4139 3369 4143 3370
rect 4427 3374 4431 3375
rect 4427 3369 4431 3370
rect 4691 3374 4695 3375
rect 4691 3369 4695 3370
rect 4803 3374 4807 3375
rect 4803 3369 4807 3370
rect 4939 3374 4943 3375
rect 4939 3369 4943 3370
rect 5075 3374 5079 3375
rect 5075 3369 5079 3370
rect 5179 3374 5183 3375
rect 5179 3369 5183 3370
rect 5211 3374 5215 3375
rect 5211 3369 5215 3370
rect 5347 3374 5351 3375
rect 5347 3369 5351 3370
rect 5427 3374 5431 3375
rect 5427 3369 5431 3370
rect 3235 3362 3239 3363
rect 3235 3357 3239 3358
rect 3267 3362 3271 3363
rect 3267 3357 3271 3358
rect 3451 3362 3455 3363
rect 3451 3357 3455 3358
rect 3651 3362 3655 3363
rect 3651 3357 3655 3358
rect 3799 3362 3803 3363
rect 3799 3357 3803 3358
rect 3114 3303 3120 3304
rect 3114 3299 3115 3303
rect 3119 3299 3120 3303
rect 3114 3298 3120 3299
rect 3268 3296 3270 3357
rect 3274 3343 3280 3344
rect 3274 3339 3275 3343
rect 3279 3339 3280 3343
rect 3274 3338 3280 3339
rect 3266 3295 3272 3296
rect 3266 3291 3267 3295
rect 3271 3291 3272 3295
rect 3266 3290 3272 3291
rect 3110 3280 3116 3281
rect 3276 3280 3278 3338
rect 3800 3297 3802 3357
rect 3840 3309 3842 3369
rect 3838 3308 3844 3309
rect 3860 3308 3862 3369
rect 4140 3308 4142 3369
rect 4262 3363 4268 3364
rect 4262 3359 4263 3363
rect 4267 3359 4268 3363
rect 4262 3358 4268 3359
rect 4146 3355 4152 3356
rect 4146 3351 4147 3355
rect 4151 3351 4152 3355
rect 4146 3350 4152 3351
rect 3838 3304 3839 3308
rect 3843 3304 3844 3308
rect 3838 3303 3844 3304
rect 3858 3307 3864 3308
rect 3858 3303 3859 3307
rect 3863 3303 3864 3307
rect 3858 3302 3864 3303
rect 4138 3307 4144 3308
rect 4138 3303 4139 3307
rect 4143 3303 4144 3307
rect 4138 3302 4144 3303
rect 3798 3296 3804 3297
rect 3798 3292 3799 3296
rect 3803 3292 3804 3296
rect 3886 3292 3892 3293
rect 3798 3291 3804 3292
rect 3838 3291 3844 3292
rect 3838 3287 3839 3291
rect 3843 3287 3844 3291
rect 3886 3288 3887 3292
rect 3891 3288 3892 3292
rect 3886 3287 3892 3288
rect 3838 3286 3844 3287
rect 3294 3280 3300 3281
rect 3090 3279 3096 3280
rect 3090 3275 3091 3279
rect 3095 3275 3096 3279
rect 3110 3276 3111 3280
rect 3115 3276 3116 3280
rect 3110 3275 3116 3276
rect 3274 3279 3280 3280
rect 3274 3275 3275 3279
rect 3279 3275 3280 3279
rect 3294 3276 3295 3280
rect 3299 3276 3300 3280
rect 3294 3275 3300 3276
rect 3402 3279 3408 3280
rect 3402 3275 3403 3279
rect 3407 3275 3408 3279
rect 3090 3274 3096 3275
rect 3112 3251 3114 3275
rect 3274 3274 3280 3275
rect 3296 3251 3298 3275
rect 3402 3274 3408 3275
rect 3798 3279 3804 3280
rect 3798 3275 3799 3279
rect 3803 3275 3804 3279
rect 3798 3274 3804 3275
rect 3111 3250 3115 3251
rect 3111 3245 3115 3246
rect 3207 3250 3211 3251
rect 3207 3245 3211 3246
rect 3295 3250 3299 3251
rect 3295 3245 3299 3246
rect 3208 3221 3210 3245
rect 3206 3220 3212 3221
rect 2742 3216 2743 3220
rect 2747 3216 2748 3220
rect 2742 3215 2748 3216
rect 2854 3219 2860 3220
rect 2854 3215 2855 3219
rect 2859 3215 2860 3219
rect 2974 3216 2975 3220
rect 2979 3216 2980 3220
rect 2974 3215 2980 3216
rect 3070 3219 3076 3220
rect 3070 3215 3071 3219
rect 3075 3215 3076 3219
rect 3206 3216 3207 3220
rect 3211 3216 3212 3220
rect 3206 3215 3212 3216
rect 3298 3219 3304 3220
rect 3298 3215 3299 3219
rect 3303 3215 3304 3219
rect 2854 3214 2860 3215
rect 3070 3214 3076 3215
rect 3298 3214 3304 3215
rect 2714 3205 2720 3206
rect 2714 3201 2715 3205
rect 2719 3201 2720 3205
rect 2714 3200 2720 3201
rect 2654 3155 2660 3156
rect 2654 3151 2655 3155
rect 2659 3151 2660 3155
rect 2654 3150 2660 3151
rect 2716 3139 2718 3200
rect 2856 3156 2858 3214
rect 2946 3205 2952 3206
rect 2946 3201 2947 3205
rect 2951 3201 2952 3205
rect 2946 3200 2952 3201
rect 3178 3205 3184 3206
rect 3178 3201 3179 3205
rect 3183 3201 3184 3205
rect 3178 3200 3184 3201
rect 2854 3155 2860 3156
rect 2854 3151 2855 3155
rect 2859 3151 2860 3155
rect 2854 3150 2860 3151
rect 2898 3147 2904 3148
rect 2898 3143 2899 3147
rect 2903 3143 2904 3147
rect 2898 3142 2904 3143
rect 2715 3138 2719 3139
rect 2715 3133 2719 3134
rect 2779 3138 2783 3139
rect 2779 3133 2783 3134
rect 2594 3123 2600 3124
rect 2594 3119 2595 3123
rect 2599 3119 2600 3123
rect 2594 3118 2600 3119
rect 2780 3072 2782 3133
rect 2874 3119 2880 3120
rect 2874 3115 2875 3119
rect 2879 3115 2880 3119
rect 2874 3114 2880 3115
rect 2876 3080 2878 3114
rect 2874 3079 2880 3080
rect 2874 3075 2875 3079
rect 2879 3075 2880 3079
rect 2874 3074 2880 3075
rect 1974 3068 1975 3072
rect 1979 3068 1980 3072
rect 1974 3067 1980 3068
rect 2482 3071 2488 3072
rect 2482 3067 2483 3071
rect 2487 3067 2488 3071
rect 2482 3066 2488 3067
rect 2778 3071 2784 3072
rect 2778 3067 2779 3071
rect 2783 3067 2784 3071
rect 2778 3066 2784 3067
rect 2510 3056 2516 3057
rect 2806 3056 2812 3057
rect 2900 3056 2902 3142
rect 2948 3139 2950 3200
rect 3180 3139 3182 3200
rect 2947 3138 2951 3139
rect 2947 3133 2951 3134
rect 3075 3138 3079 3139
rect 3075 3133 3079 3134
rect 3179 3138 3183 3139
rect 3179 3133 3183 3134
rect 3076 3072 3078 3133
rect 3300 3124 3302 3214
rect 3404 3156 3406 3274
rect 3800 3251 3802 3274
rect 3447 3250 3451 3251
rect 3447 3245 3451 3246
rect 3799 3250 3803 3251
rect 3799 3245 3803 3246
rect 3448 3221 3450 3245
rect 3800 3222 3802 3245
rect 3840 3239 3842 3286
rect 3888 3239 3890 3287
rect 3839 3238 3843 3239
rect 3839 3233 3843 3234
rect 3887 3238 3891 3239
rect 3887 3233 3891 3234
rect 3911 3238 3915 3239
rect 3911 3233 3915 3234
rect 3798 3221 3804 3222
rect 3446 3220 3452 3221
rect 3446 3216 3447 3220
rect 3451 3216 3452 3220
rect 3446 3215 3452 3216
rect 3542 3219 3548 3220
rect 3542 3215 3543 3219
rect 3547 3215 3548 3219
rect 3798 3217 3799 3221
rect 3803 3217 3804 3221
rect 3798 3216 3804 3217
rect 3542 3214 3548 3215
rect 3418 3205 3424 3206
rect 3418 3201 3419 3205
rect 3423 3201 3424 3205
rect 3418 3200 3424 3201
rect 3402 3155 3408 3156
rect 3402 3151 3403 3155
rect 3407 3151 3408 3155
rect 3402 3150 3408 3151
rect 3420 3139 3422 3200
rect 3544 3148 3546 3214
rect 3840 3210 3842 3233
rect 3838 3209 3844 3210
rect 3912 3209 3914 3233
rect 3838 3205 3839 3209
rect 3843 3205 3844 3209
rect 3798 3204 3804 3205
rect 3838 3204 3844 3205
rect 3910 3208 3916 3209
rect 4148 3208 4150 3350
rect 4166 3292 4172 3293
rect 4264 3292 4266 3358
rect 4428 3308 4430 3369
rect 4522 3355 4528 3356
rect 4522 3351 4523 3355
rect 4527 3351 4528 3355
rect 4522 3350 4528 3351
rect 4524 3325 4526 3350
rect 4523 3324 4527 3325
rect 4523 3319 4527 3320
rect 4692 3308 4694 3369
rect 4698 3355 4704 3356
rect 4698 3351 4699 3355
rect 4703 3351 4704 3355
rect 4698 3350 4704 3351
rect 4426 3307 4432 3308
rect 4426 3303 4427 3307
rect 4431 3303 4432 3307
rect 4426 3302 4432 3303
rect 4690 3307 4696 3308
rect 4690 3303 4691 3307
rect 4695 3303 4696 3307
rect 4690 3302 4696 3303
rect 4454 3292 4460 3293
rect 4700 3292 4702 3350
rect 4940 3308 4942 3369
rect 5059 3324 5063 3325
rect 5059 3319 5063 3320
rect 4938 3307 4944 3308
rect 4938 3303 4939 3307
rect 4943 3303 4944 3307
rect 4938 3302 4944 3303
rect 4718 3292 4724 3293
rect 4966 3292 4972 3293
rect 5060 3292 5062 3319
rect 5180 3308 5182 3369
rect 5302 3363 5308 3364
rect 5302 3359 5303 3363
rect 5307 3359 5308 3363
rect 5302 3358 5308 3359
rect 5178 3307 5184 3308
rect 5178 3303 5179 3307
rect 5183 3303 5184 3307
rect 5178 3302 5184 3303
rect 5206 3292 5212 3293
rect 5304 3292 5306 3358
rect 5418 3351 5424 3352
rect 5418 3347 5419 3351
rect 5423 3347 5424 3351
rect 5418 3346 5424 3347
rect 5420 3300 5422 3346
rect 5428 3308 5430 3369
rect 5472 3360 5474 3450
rect 5662 3440 5668 3441
rect 5662 3436 5663 3440
rect 5667 3436 5668 3440
rect 5662 3435 5668 3436
rect 5664 3375 5666 3435
rect 5663 3374 5667 3375
rect 5663 3369 5667 3370
rect 5470 3359 5476 3360
rect 5470 3355 5471 3359
rect 5475 3355 5476 3359
rect 5470 3354 5476 3355
rect 5664 3309 5666 3369
rect 5662 3308 5668 3309
rect 5426 3307 5432 3308
rect 5426 3303 5427 3307
rect 5431 3303 5432 3307
rect 5662 3304 5663 3308
rect 5667 3304 5668 3308
rect 5662 3303 5668 3304
rect 5426 3302 5432 3303
rect 5418 3299 5424 3300
rect 5418 3295 5419 3299
rect 5423 3295 5424 3299
rect 5418 3294 5424 3295
rect 5454 3292 5460 3293
rect 4166 3288 4167 3292
rect 4171 3288 4172 3292
rect 4166 3287 4172 3288
rect 4262 3291 4268 3292
rect 4262 3287 4263 3291
rect 4267 3287 4268 3291
rect 4454 3288 4455 3292
rect 4459 3288 4460 3292
rect 4454 3287 4460 3288
rect 4698 3291 4704 3292
rect 4698 3287 4699 3291
rect 4703 3287 4704 3291
rect 4718 3288 4719 3292
rect 4723 3288 4724 3292
rect 4718 3287 4724 3288
rect 4818 3291 4824 3292
rect 4818 3287 4819 3291
rect 4823 3287 4824 3291
rect 4966 3288 4967 3292
rect 4971 3288 4972 3292
rect 4966 3287 4972 3288
rect 5058 3291 5064 3292
rect 5058 3287 5059 3291
rect 5063 3287 5064 3291
rect 5206 3288 5207 3292
rect 5211 3288 5212 3292
rect 5206 3287 5212 3288
rect 5302 3291 5308 3292
rect 5302 3287 5303 3291
rect 5307 3287 5308 3291
rect 5454 3288 5455 3292
rect 5459 3288 5460 3292
rect 5454 3287 5460 3288
rect 5662 3291 5668 3292
rect 5662 3287 5663 3291
rect 5667 3287 5668 3291
rect 4168 3239 4170 3287
rect 4262 3286 4268 3287
rect 4456 3239 4458 3287
rect 4698 3286 4704 3287
rect 4720 3239 4722 3287
rect 4818 3286 4824 3287
rect 4167 3238 4171 3239
rect 4167 3233 4171 3234
rect 4183 3238 4187 3239
rect 4183 3233 4187 3234
rect 4439 3238 4443 3239
rect 4439 3233 4443 3234
rect 4455 3238 4459 3239
rect 4455 3233 4459 3234
rect 4687 3238 4691 3239
rect 4687 3233 4691 3234
rect 4719 3238 4723 3239
rect 4719 3233 4723 3234
rect 4184 3209 4186 3233
rect 4440 3209 4442 3233
rect 4688 3209 4690 3233
rect 4182 3208 4188 3209
rect 3910 3204 3911 3208
rect 3915 3204 3916 3208
rect 3798 3200 3799 3204
rect 3803 3200 3804 3204
rect 3910 3203 3916 3204
rect 4146 3207 4152 3208
rect 4146 3203 4147 3207
rect 4151 3203 4152 3207
rect 4182 3204 4183 3208
rect 4187 3204 4188 3208
rect 4182 3203 4188 3204
rect 4438 3208 4444 3209
rect 4686 3208 4692 3209
rect 4438 3204 4439 3208
rect 4443 3204 4444 3208
rect 4438 3203 4444 3204
rect 4534 3207 4540 3208
rect 4534 3203 4535 3207
rect 4539 3203 4540 3207
rect 4686 3204 4687 3208
rect 4691 3204 4692 3208
rect 4686 3203 4692 3204
rect 4778 3207 4784 3208
rect 4778 3203 4779 3207
rect 4783 3203 4784 3207
rect 4146 3202 4152 3203
rect 4534 3202 4540 3203
rect 4778 3202 4784 3203
rect 3798 3199 3804 3200
rect 3542 3147 3548 3148
rect 3542 3143 3543 3147
rect 3547 3143 3548 3147
rect 3542 3142 3548 3143
rect 3800 3139 3802 3199
rect 3882 3193 3888 3194
rect 3838 3192 3844 3193
rect 3838 3188 3839 3192
rect 3843 3188 3844 3192
rect 3882 3189 3883 3193
rect 3887 3189 3888 3193
rect 3882 3188 3888 3189
rect 4154 3193 4160 3194
rect 4154 3189 4155 3193
rect 4159 3189 4160 3193
rect 4154 3188 4160 3189
rect 4410 3193 4416 3194
rect 4410 3189 4411 3193
rect 4415 3189 4416 3193
rect 4410 3188 4416 3189
rect 3838 3187 3844 3188
rect 3371 3138 3375 3139
rect 3371 3133 3375 3134
rect 3419 3138 3423 3139
rect 3419 3133 3423 3134
rect 3651 3138 3655 3139
rect 3651 3133 3655 3134
rect 3799 3138 3803 3139
rect 3799 3133 3803 3134
rect 3298 3123 3304 3124
rect 3298 3119 3299 3123
rect 3303 3119 3304 3123
rect 3298 3118 3304 3119
rect 3214 3079 3220 3080
rect 3214 3075 3215 3079
rect 3219 3075 3220 3079
rect 3214 3074 3220 3075
rect 3074 3071 3080 3072
rect 3074 3067 3075 3071
rect 3079 3067 3080 3071
rect 3074 3066 3080 3067
rect 3102 3056 3108 3057
rect 1974 3055 1980 3056
rect 1974 3051 1975 3055
rect 1979 3051 1980 3055
rect 2510 3052 2511 3056
rect 2515 3052 2516 3056
rect 2510 3051 2516 3052
rect 2606 3055 2612 3056
rect 2606 3051 2607 3055
rect 2611 3051 2612 3055
rect 2806 3052 2807 3056
rect 2811 3052 2812 3056
rect 2806 3051 2812 3052
rect 2898 3055 2904 3056
rect 2898 3051 2899 3055
rect 2903 3051 2904 3055
rect 3102 3052 3103 3056
rect 3107 3052 3108 3056
rect 3102 3051 3108 3052
rect 1974 3050 1980 3051
rect 1934 3044 1940 3045
rect 1626 3043 1632 3044
rect 1626 3039 1627 3043
rect 1631 3039 1632 3043
rect 1626 3038 1632 3039
rect 1786 3043 1792 3044
rect 1786 3039 1787 3043
rect 1791 3039 1792 3043
rect 1934 3040 1935 3044
rect 1939 3040 1940 3044
rect 1934 3039 1940 3040
rect 1786 3038 1792 3039
rect 1654 3028 1660 3029
rect 906 3027 912 3028
rect 906 3023 907 3027
rect 911 3023 912 3027
rect 926 3024 927 3028
rect 931 3024 932 3028
rect 926 3023 932 3024
rect 1026 3027 1032 3028
rect 1026 3023 1027 3027
rect 1031 3023 1032 3027
rect 1118 3024 1119 3028
rect 1123 3024 1124 3028
rect 1118 3023 1124 3024
rect 1282 3027 1288 3028
rect 1282 3023 1283 3027
rect 1287 3023 1288 3027
rect 1302 3024 1303 3028
rect 1307 3024 1308 3028
rect 1302 3023 1308 3024
rect 1458 3027 1464 3028
rect 1458 3023 1459 3027
rect 1463 3023 1464 3027
rect 1478 3024 1479 3028
rect 1483 3024 1484 3028
rect 1478 3023 1484 3024
rect 1574 3027 1580 3028
rect 1574 3023 1575 3027
rect 1579 3023 1580 3027
rect 1654 3024 1655 3028
rect 1659 3024 1660 3028
rect 1654 3023 1660 3024
rect 1814 3028 1820 3029
rect 1814 3024 1815 3028
rect 1819 3024 1820 3028
rect 1814 3023 1820 3024
rect 1934 3027 1940 3028
rect 1934 3023 1935 3027
rect 1939 3023 1940 3027
rect 906 3022 912 3023
rect 928 2995 930 3023
rect 1026 3022 1032 3023
rect 1120 2995 1122 3023
rect 1282 3022 1288 3023
rect 1304 2995 1306 3023
rect 1458 3022 1464 3023
rect 1480 2995 1482 3023
rect 1574 3022 1580 3023
rect 1656 2995 1658 3023
rect 1816 2995 1818 3023
rect 1934 3022 1940 3023
rect 1936 2995 1938 3022
rect 1976 3019 1978 3050
rect 2512 3019 2514 3051
rect 2606 3050 2612 3051
rect 1975 3018 1979 3019
rect 1975 3013 1979 3014
rect 2191 3018 2195 3019
rect 2191 3013 2195 3014
rect 2351 3018 2355 3019
rect 2351 3013 2355 3014
rect 2511 3018 2515 3019
rect 2511 3013 2515 3014
rect 2519 3018 2523 3019
rect 2519 3013 2523 3014
rect 927 2994 931 2995
rect 927 2989 931 2990
rect 1119 2994 1123 2995
rect 1119 2989 1123 2990
rect 1303 2994 1307 2995
rect 1303 2989 1307 2990
rect 1479 2994 1483 2995
rect 1479 2989 1483 2990
rect 1655 2994 1659 2995
rect 1655 2989 1659 2990
rect 1815 2994 1819 2995
rect 1815 2989 1819 2990
rect 1935 2994 1939 2995
rect 1976 2990 1978 3013
rect 1935 2989 1939 2990
rect 1974 2989 1980 2990
rect 2192 2989 2194 3013
rect 2352 2989 2354 3013
rect 2520 2989 2522 3013
rect 1936 2966 1938 2989
rect 1974 2985 1975 2989
rect 1979 2985 1980 2989
rect 1974 2984 1980 2985
rect 2190 2988 2196 2989
rect 2350 2988 2356 2989
rect 2518 2988 2524 2989
rect 2190 2984 2191 2988
rect 2195 2984 2196 2988
rect 2190 2983 2196 2984
rect 2286 2987 2292 2988
rect 2286 2983 2287 2987
rect 2291 2983 2292 2987
rect 2350 2984 2351 2988
rect 2355 2984 2356 2988
rect 2350 2983 2356 2984
rect 2446 2987 2452 2988
rect 2446 2983 2447 2987
rect 2451 2983 2452 2987
rect 2518 2984 2519 2988
rect 2523 2984 2524 2988
rect 2518 2983 2524 2984
rect 2286 2982 2292 2983
rect 2446 2982 2452 2983
rect 2162 2973 2168 2974
rect 1974 2972 1980 2973
rect 1974 2968 1975 2972
rect 1979 2968 1980 2972
rect 2162 2969 2163 2973
rect 2167 2969 2168 2973
rect 2162 2968 2168 2969
rect 1974 2967 1980 2968
rect 1934 2965 1940 2966
rect 294 2960 295 2964
rect 299 2960 300 2964
rect 294 2959 300 2960
rect 394 2963 400 2964
rect 394 2959 395 2963
rect 399 2959 400 2963
rect 430 2960 431 2964
rect 435 2960 436 2964
rect 430 2959 436 2960
rect 530 2963 536 2964
rect 530 2959 531 2963
rect 535 2959 536 2963
rect 566 2960 567 2964
rect 571 2960 572 2964
rect 566 2959 572 2960
rect 658 2963 664 2964
rect 658 2959 659 2963
rect 663 2959 664 2963
rect 702 2960 703 2964
rect 707 2960 708 2964
rect 702 2959 708 2960
rect 802 2963 808 2964
rect 802 2959 803 2963
rect 807 2959 808 2963
rect 1934 2961 1935 2965
rect 1939 2961 1940 2965
rect 1934 2960 1940 2961
rect 394 2958 400 2959
rect 530 2958 536 2959
rect 658 2958 664 2959
rect 802 2958 808 2959
rect 266 2949 272 2950
rect 266 2945 267 2949
rect 271 2945 272 2949
rect 266 2944 272 2945
rect 250 2899 256 2900
rect 250 2895 251 2899
rect 255 2895 256 2899
rect 250 2894 256 2895
rect 268 2879 270 2944
rect 396 2900 398 2958
rect 402 2949 408 2950
rect 402 2945 403 2949
rect 407 2945 408 2949
rect 402 2944 408 2945
rect 394 2899 400 2900
rect 394 2895 395 2899
rect 399 2895 400 2899
rect 394 2894 400 2895
rect 404 2879 406 2944
rect 532 2900 534 2958
rect 538 2949 544 2950
rect 538 2945 539 2949
rect 543 2945 544 2949
rect 538 2944 544 2945
rect 530 2899 536 2900
rect 530 2895 531 2899
rect 535 2895 536 2899
rect 530 2894 536 2895
rect 540 2879 542 2944
rect 111 2878 115 2879
rect 111 2873 115 2874
rect 131 2878 135 2879
rect 131 2873 135 2874
rect 227 2878 231 2879
rect 227 2873 231 2874
rect 267 2878 271 2879
rect 267 2873 271 2874
rect 363 2878 367 2879
rect 363 2873 367 2874
rect 403 2878 407 2879
rect 403 2873 407 2874
rect 499 2878 503 2879
rect 499 2873 503 2874
rect 539 2878 543 2879
rect 539 2873 543 2874
rect 635 2878 639 2879
rect 635 2873 639 2874
rect 112 2813 114 2873
rect 110 2812 116 2813
rect 228 2812 230 2873
rect 364 2812 366 2873
rect 370 2859 376 2860
rect 370 2855 371 2859
rect 375 2855 376 2859
rect 370 2854 376 2855
rect 110 2808 111 2812
rect 115 2808 116 2812
rect 110 2807 116 2808
rect 226 2811 232 2812
rect 226 2807 227 2811
rect 231 2807 232 2811
rect 226 2806 232 2807
rect 362 2811 368 2812
rect 362 2807 363 2811
rect 367 2807 368 2811
rect 362 2806 368 2807
rect 254 2796 260 2797
rect 372 2796 374 2854
rect 500 2812 502 2873
rect 506 2859 512 2860
rect 506 2855 507 2859
rect 511 2855 512 2859
rect 506 2854 512 2855
rect 498 2811 504 2812
rect 498 2807 499 2811
rect 503 2807 504 2811
rect 498 2806 504 2807
rect 390 2796 396 2797
rect 508 2796 510 2854
rect 636 2812 638 2873
rect 660 2872 662 2958
rect 674 2949 680 2950
rect 674 2945 675 2949
rect 679 2945 680 2949
rect 674 2944 680 2945
rect 1934 2948 1940 2949
rect 1934 2944 1935 2948
rect 1939 2944 1940 2948
rect 676 2879 678 2944
rect 1934 2943 1940 2944
rect 758 2899 764 2900
rect 758 2895 759 2899
rect 763 2895 764 2899
rect 758 2894 764 2895
rect 675 2878 679 2879
rect 675 2873 679 2874
rect 658 2871 664 2872
rect 658 2867 659 2871
rect 663 2867 664 2871
rect 658 2866 664 2867
rect 634 2811 640 2812
rect 634 2807 635 2811
rect 639 2807 640 2811
rect 634 2806 640 2807
rect 526 2796 532 2797
rect 110 2795 116 2796
rect 110 2791 111 2795
rect 115 2791 116 2795
rect 254 2792 255 2796
rect 259 2792 260 2796
rect 254 2791 260 2792
rect 370 2795 376 2796
rect 370 2791 371 2795
rect 375 2791 376 2795
rect 390 2792 391 2796
rect 395 2792 396 2796
rect 390 2791 396 2792
rect 506 2795 512 2796
rect 506 2791 507 2795
rect 511 2791 512 2795
rect 526 2792 527 2796
rect 531 2792 532 2796
rect 526 2791 532 2792
rect 662 2796 668 2797
rect 760 2796 762 2894
rect 1936 2879 1938 2943
rect 1976 2903 1978 2967
rect 2164 2903 2166 2968
rect 2258 2951 2264 2952
rect 2258 2947 2259 2951
rect 2263 2947 2264 2951
rect 2258 2946 2264 2947
rect 2260 2924 2262 2946
rect 2258 2923 2264 2924
rect 2258 2919 2259 2923
rect 2263 2919 2264 2923
rect 2258 2918 2264 2919
rect 1975 2902 1979 2903
rect 1975 2897 1979 2898
rect 1995 2902 1999 2903
rect 1995 2897 1999 2898
rect 2131 2902 2135 2903
rect 2131 2897 2135 2898
rect 2163 2902 2167 2903
rect 2163 2897 2167 2898
rect 2267 2902 2271 2903
rect 2267 2897 2271 2898
rect 771 2878 775 2879
rect 771 2873 775 2874
rect 1935 2878 1939 2879
rect 1935 2873 1939 2874
rect 772 2812 774 2873
rect 894 2863 900 2864
rect 894 2859 895 2863
rect 899 2859 900 2863
rect 894 2858 900 2859
rect 770 2811 776 2812
rect 770 2807 771 2811
rect 775 2807 776 2811
rect 770 2806 776 2807
rect 798 2796 804 2797
rect 662 2792 663 2796
rect 667 2792 668 2796
rect 662 2791 668 2792
rect 758 2795 764 2796
rect 758 2791 759 2795
rect 763 2791 764 2795
rect 798 2792 799 2796
rect 803 2792 804 2796
rect 798 2791 804 2792
rect 110 2790 116 2791
rect 112 2763 114 2790
rect 256 2763 258 2791
rect 370 2790 376 2791
rect 392 2763 394 2791
rect 506 2790 512 2791
rect 528 2763 530 2791
rect 664 2763 666 2791
rect 758 2790 764 2791
rect 800 2763 802 2791
rect 111 2762 115 2763
rect 111 2757 115 2758
rect 255 2762 259 2763
rect 255 2757 259 2758
rect 375 2762 379 2763
rect 375 2757 379 2758
rect 391 2762 395 2763
rect 391 2757 395 2758
rect 527 2762 531 2763
rect 527 2757 531 2758
rect 575 2762 579 2763
rect 575 2757 579 2758
rect 663 2762 667 2763
rect 663 2757 667 2758
rect 799 2762 803 2763
rect 799 2757 803 2758
rect 112 2734 114 2757
rect 110 2733 116 2734
rect 376 2733 378 2757
rect 576 2733 578 2757
rect 800 2733 802 2757
rect 110 2729 111 2733
rect 115 2729 116 2733
rect 110 2728 116 2729
rect 374 2732 380 2733
rect 574 2732 580 2733
rect 798 2732 804 2733
rect 896 2732 898 2858
rect 1936 2813 1938 2873
rect 1976 2837 1978 2897
rect 1974 2836 1980 2837
rect 1996 2836 1998 2897
rect 2090 2883 2096 2884
rect 2090 2879 2091 2883
rect 2095 2879 2096 2883
rect 2090 2878 2096 2879
rect 2092 2856 2094 2878
rect 2090 2855 2096 2856
rect 2090 2851 2091 2855
rect 2095 2851 2096 2855
rect 2090 2850 2096 2851
rect 2132 2836 2134 2897
rect 2138 2883 2144 2884
rect 2138 2879 2139 2883
rect 2143 2879 2144 2883
rect 2138 2878 2144 2879
rect 1974 2832 1975 2836
rect 1979 2832 1980 2836
rect 1974 2831 1980 2832
rect 1994 2835 2000 2836
rect 1994 2831 1995 2835
rect 1999 2831 2000 2835
rect 1994 2830 2000 2831
rect 2130 2835 2136 2836
rect 2130 2831 2131 2835
rect 2135 2831 2136 2835
rect 2130 2830 2136 2831
rect 2022 2820 2028 2821
rect 2140 2820 2142 2878
rect 2268 2836 2270 2897
rect 2288 2888 2290 2982
rect 2322 2973 2328 2974
rect 2322 2969 2323 2973
rect 2327 2969 2328 2973
rect 2322 2968 2328 2969
rect 2324 2903 2326 2968
rect 2448 2952 2450 2982
rect 2490 2973 2496 2974
rect 2490 2969 2491 2973
rect 2495 2969 2496 2973
rect 2490 2968 2496 2969
rect 2446 2951 2452 2952
rect 2446 2947 2447 2951
rect 2451 2947 2452 2951
rect 2446 2946 2452 2947
rect 2492 2903 2494 2968
rect 2608 2924 2610 3050
rect 2808 3019 2810 3051
rect 2898 3050 2904 3051
rect 3104 3019 3106 3051
rect 2703 3018 2707 3019
rect 2703 3013 2707 3014
rect 2807 3018 2811 3019
rect 2807 3013 2811 3014
rect 2903 3018 2907 3019
rect 2903 3013 2907 3014
rect 3103 3018 3107 3019
rect 3103 3013 3107 3014
rect 3119 3018 3123 3019
rect 3119 3013 3123 3014
rect 2704 2989 2706 3013
rect 2904 2989 2906 3013
rect 3120 2989 3122 3013
rect 2702 2988 2708 2989
rect 2902 2988 2908 2989
rect 3118 2988 3124 2989
rect 3216 2988 3218 3074
rect 3372 3072 3374 3133
rect 3378 3119 3384 3120
rect 3378 3115 3379 3119
rect 3383 3115 3384 3119
rect 3378 3114 3384 3115
rect 3370 3071 3376 3072
rect 3370 3067 3371 3071
rect 3375 3067 3376 3071
rect 3370 3066 3376 3067
rect 3380 3056 3382 3114
rect 3652 3072 3654 3133
rect 3658 3119 3664 3120
rect 3658 3115 3659 3119
rect 3663 3115 3664 3119
rect 3658 3114 3664 3115
rect 3650 3071 3656 3072
rect 3650 3067 3651 3071
rect 3655 3067 3656 3071
rect 3650 3066 3656 3067
rect 3398 3056 3404 3057
rect 3660 3056 3662 3114
rect 3800 3073 3802 3133
rect 3840 3123 3842 3187
rect 3884 3123 3886 3188
rect 4050 3143 4056 3144
rect 4050 3139 4051 3143
rect 4055 3139 4056 3143
rect 4050 3138 4056 3139
rect 3839 3122 3843 3123
rect 3839 3117 3843 3118
rect 3883 3122 3887 3123
rect 3883 3117 3887 3118
rect 3931 3122 3935 3123
rect 3931 3117 3935 3118
rect 3798 3072 3804 3073
rect 3798 3068 3799 3072
rect 3803 3068 3804 3072
rect 3798 3067 3804 3068
rect 3840 3057 3842 3117
rect 3678 3056 3684 3057
rect 3838 3056 3844 3057
rect 3932 3056 3934 3117
rect 3378 3055 3384 3056
rect 3378 3051 3379 3055
rect 3383 3051 3384 3055
rect 3398 3052 3399 3056
rect 3403 3052 3404 3056
rect 3398 3051 3404 3052
rect 3658 3055 3664 3056
rect 3658 3051 3659 3055
rect 3663 3051 3664 3055
rect 3678 3052 3679 3056
rect 3683 3052 3684 3056
rect 3678 3051 3684 3052
rect 3770 3055 3776 3056
rect 3770 3051 3771 3055
rect 3775 3051 3776 3055
rect 3378 3050 3384 3051
rect 3400 3019 3402 3051
rect 3658 3050 3664 3051
rect 3680 3019 3682 3051
rect 3770 3050 3776 3051
rect 3798 3055 3804 3056
rect 3798 3051 3799 3055
rect 3803 3051 3804 3055
rect 3838 3052 3839 3056
rect 3843 3052 3844 3056
rect 3838 3051 3844 3052
rect 3930 3055 3936 3056
rect 3930 3051 3931 3055
rect 3935 3051 3936 3055
rect 3798 3050 3804 3051
rect 3930 3050 3936 3051
rect 3335 3018 3339 3019
rect 3335 3013 3339 3014
rect 3399 3018 3403 3019
rect 3399 3013 3403 3014
rect 3559 3018 3563 3019
rect 3559 3013 3563 3014
rect 3679 3018 3683 3019
rect 3679 3013 3683 3014
rect 3336 2989 3338 3013
rect 3560 2989 3562 3013
rect 3334 2988 3340 2989
rect 3558 2988 3564 2989
rect 2638 2987 2644 2988
rect 2638 2983 2639 2987
rect 2643 2983 2644 2987
rect 2702 2984 2703 2988
rect 2707 2984 2708 2988
rect 2702 2983 2708 2984
rect 2794 2987 2800 2988
rect 2794 2983 2795 2987
rect 2799 2983 2800 2987
rect 2902 2984 2903 2988
rect 2907 2984 2908 2988
rect 2902 2983 2908 2984
rect 3002 2987 3008 2988
rect 3002 2983 3003 2987
rect 3007 2983 3008 2987
rect 3118 2984 3119 2988
rect 3123 2984 3124 2988
rect 3118 2983 3124 2984
rect 3214 2987 3220 2988
rect 3214 2983 3215 2987
rect 3219 2983 3220 2987
rect 3334 2984 3335 2988
rect 3339 2984 3340 2988
rect 3334 2983 3340 2984
rect 3426 2987 3432 2988
rect 3426 2983 3427 2987
rect 3431 2983 3432 2987
rect 3558 2984 3559 2988
rect 3563 2984 3564 2988
rect 3558 2983 3564 2984
rect 3650 2987 3656 2988
rect 3650 2983 3651 2987
rect 3655 2983 3656 2987
rect 2638 2982 2644 2983
rect 2794 2982 2800 2983
rect 3002 2982 3008 2983
rect 3214 2982 3220 2983
rect 3426 2982 3432 2983
rect 3650 2982 3656 2983
rect 2640 2924 2642 2982
rect 2674 2973 2680 2974
rect 2674 2969 2675 2973
rect 2679 2969 2680 2973
rect 2674 2968 2680 2969
rect 2606 2923 2612 2924
rect 2606 2919 2607 2923
rect 2611 2919 2612 2923
rect 2606 2918 2612 2919
rect 2638 2923 2644 2924
rect 2638 2919 2639 2923
rect 2643 2919 2644 2923
rect 2638 2918 2644 2919
rect 2676 2903 2678 2968
rect 2796 2916 2798 2982
rect 2874 2973 2880 2974
rect 2874 2969 2875 2973
rect 2879 2969 2880 2973
rect 2874 2968 2880 2969
rect 2794 2915 2800 2916
rect 2794 2911 2795 2915
rect 2799 2911 2800 2915
rect 2794 2910 2800 2911
rect 2876 2903 2878 2968
rect 3004 2924 3006 2982
rect 3090 2973 3096 2974
rect 3090 2969 3091 2973
rect 3095 2969 3096 2973
rect 3090 2968 3096 2969
rect 3306 2973 3312 2974
rect 3306 2969 3307 2973
rect 3311 2969 3312 2973
rect 3306 2968 3312 2969
rect 2958 2923 2964 2924
rect 2958 2919 2959 2923
rect 2963 2919 2964 2923
rect 2958 2918 2964 2919
rect 3002 2923 3008 2924
rect 3002 2919 3003 2923
rect 3007 2919 3008 2923
rect 3002 2918 3008 2919
rect 2323 2902 2327 2903
rect 2323 2897 2327 2898
rect 2403 2902 2407 2903
rect 2403 2897 2407 2898
rect 2491 2902 2495 2903
rect 2491 2897 2495 2898
rect 2539 2902 2543 2903
rect 2539 2897 2543 2898
rect 2675 2902 2679 2903
rect 2675 2897 2679 2898
rect 2683 2902 2687 2903
rect 2683 2897 2687 2898
rect 2835 2902 2839 2903
rect 2835 2897 2839 2898
rect 2875 2902 2879 2903
rect 2875 2897 2879 2898
rect 2286 2887 2292 2888
rect 2286 2883 2287 2887
rect 2291 2883 2292 2887
rect 2286 2882 2292 2883
rect 2404 2836 2406 2897
rect 2410 2883 2416 2884
rect 2410 2879 2411 2883
rect 2415 2879 2416 2883
rect 2410 2878 2416 2879
rect 2266 2835 2272 2836
rect 2266 2831 2267 2835
rect 2271 2831 2272 2835
rect 2266 2830 2272 2831
rect 2402 2835 2408 2836
rect 2402 2831 2403 2835
rect 2407 2831 2408 2835
rect 2402 2830 2408 2831
rect 2158 2820 2164 2821
rect 2294 2820 2300 2821
rect 2412 2820 2414 2878
rect 2540 2836 2542 2897
rect 2546 2883 2552 2884
rect 2546 2879 2547 2883
rect 2551 2879 2552 2883
rect 2546 2878 2552 2879
rect 2538 2835 2544 2836
rect 2538 2831 2539 2835
rect 2543 2831 2544 2835
rect 2538 2830 2544 2831
rect 2430 2820 2436 2821
rect 2548 2820 2550 2878
rect 2662 2855 2668 2856
rect 2662 2851 2663 2855
rect 2667 2851 2668 2855
rect 2662 2850 2668 2851
rect 2566 2820 2572 2821
rect 2664 2820 2666 2850
rect 2684 2836 2686 2897
rect 2718 2887 2724 2888
rect 2718 2883 2719 2887
rect 2723 2883 2724 2887
rect 2718 2882 2724 2883
rect 2682 2835 2688 2836
rect 2682 2831 2683 2835
rect 2687 2831 2688 2835
rect 2682 2830 2688 2831
rect 2710 2820 2716 2821
rect 1974 2819 1980 2820
rect 1974 2815 1975 2819
rect 1979 2815 1980 2819
rect 2022 2816 2023 2820
rect 2027 2816 2028 2820
rect 2022 2815 2028 2816
rect 2138 2819 2144 2820
rect 2138 2815 2139 2819
rect 2143 2815 2144 2819
rect 2158 2816 2159 2820
rect 2163 2816 2164 2820
rect 2158 2815 2164 2816
rect 2250 2819 2256 2820
rect 2250 2815 2251 2819
rect 2255 2815 2256 2819
rect 2294 2816 2295 2820
rect 2299 2816 2300 2820
rect 2294 2815 2300 2816
rect 2410 2819 2416 2820
rect 2410 2815 2411 2819
rect 2415 2815 2416 2819
rect 2430 2816 2431 2820
rect 2435 2816 2436 2820
rect 2430 2815 2436 2816
rect 2546 2819 2552 2820
rect 2546 2815 2547 2819
rect 2551 2815 2552 2819
rect 2566 2816 2567 2820
rect 2571 2816 2572 2820
rect 2566 2815 2572 2816
rect 2662 2819 2668 2820
rect 2662 2815 2663 2819
rect 2667 2815 2668 2819
rect 2710 2816 2711 2820
rect 2715 2816 2716 2820
rect 2710 2815 2716 2816
rect 1974 2814 1980 2815
rect 1934 2812 1940 2813
rect 1934 2808 1935 2812
rect 1939 2808 1940 2812
rect 1934 2807 1940 2808
rect 1934 2795 1940 2796
rect 1934 2791 1935 2795
rect 1939 2791 1940 2795
rect 1934 2790 1940 2791
rect 918 2779 924 2780
rect 918 2775 919 2779
rect 923 2775 924 2779
rect 918 2774 924 2775
rect 374 2728 375 2732
rect 379 2728 380 2732
rect 374 2727 380 2728
rect 474 2731 480 2732
rect 474 2727 475 2731
rect 479 2727 480 2731
rect 574 2728 575 2732
rect 579 2728 580 2732
rect 574 2727 580 2728
rect 674 2731 680 2732
rect 674 2727 675 2731
rect 679 2727 680 2731
rect 798 2728 799 2732
rect 803 2728 804 2732
rect 798 2727 804 2728
rect 894 2731 900 2732
rect 894 2727 895 2731
rect 899 2727 900 2731
rect 474 2726 480 2727
rect 674 2726 680 2727
rect 894 2726 900 2727
rect 346 2717 352 2718
rect 110 2716 116 2717
rect 110 2712 111 2716
rect 115 2712 116 2716
rect 346 2713 347 2717
rect 351 2713 352 2717
rect 346 2712 352 2713
rect 110 2711 116 2712
rect 112 2651 114 2711
rect 348 2651 350 2712
rect 476 2668 478 2726
rect 546 2717 552 2718
rect 546 2713 547 2717
rect 551 2713 552 2717
rect 546 2712 552 2713
rect 474 2667 480 2668
rect 474 2663 475 2667
rect 479 2663 480 2667
rect 474 2662 480 2663
rect 506 2659 512 2660
rect 506 2655 507 2659
rect 511 2655 512 2659
rect 506 2654 512 2655
rect 111 2650 115 2651
rect 111 2645 115 2646
rect 347 2650 351 2651
rect 347 2645 351 2646
rect 387 2650 391 2651
rect 387 2645 391 2646
rect 112 2585 114 2645
rect 110 2584 116 2585
rect 388 2584 390 2645
rect 110 2580 111 2584
rect 115 2580 116 2584
rect 110 2579 116 2580
rect 386 2583 392 2584
rect 386 2579 387 2583
rect 391 2579 392 2583
rect 386 2578 392 2579
rect 414 2568 420 2569
rect 508 2568 510 2654
rect 548 2651 550 2712
rect 676 2668 678 2726
rect 770 2717 776 2718
rect 770 2713 771 2717
rect 775 2713 776 2717
rect 770 2712 776 2713
rect 674 2667 680 2668
rect 674 2663 675 2667
rect 679 2663 680 2667
rect 674 2662 680 2663
rect 772 2651 774 2712
rect 920 2668 922 2774
rect 1936 2763 1938 2790
rect 1976 2787 1978 2814
rect 2024 2787 2026 2815
rect 2138 2814 2144 2815
rect 2160 2787 2162 2815
rect 2250 2814 2256 2815
rect 1975 2786 1979 2787
rect 1975 2781 1979 2782
rect 2023 2786 2027 2787
rect 2023 2781 2027 2782
rect 2159 2786 2163 2787
rect 2159 2781 2163 2782
rect 1039 2762 1043 2763
rect 1039 2757 1043 2758
rect 1295 2762 1299 2763
rect 1295 2757 1299 2758
rect 1567 2762 1571 2763
rect 1567 2757 1571 2758
rect 1815 2762 1819 2763
rect 1815 2757 1819 2758
rect 1935 2762 1939 2763
rect 1976 2758 1978 2781
rect 1935 2757 1939 2758
rect 1974 2757 1980 2758
rect 2024 2757 2026 2781
rect 2160 2757 2162 2781
rect 1040 2733 1042 2757
rect 1296 2733 1298 2757
rect 1568 2733 1570 2757
rect 1816 2733 1818 2757
rect 1936 2734 1938 2757
rect 1974 2753 1975 2757
rect 1979 2753 1980 2757
rect 1974 2752 1980 2753
rect 2022 2756 2028 2757
rect 2158 2756 2164 2757
rect 2022 2752 2023 2756
rect 2027 2752 2028 2756
rect 2022 2751 2028 2752
rect 2114 2755 2120 2756
rect 2114 2751 2115 2755
rect 2119 2751 2120 2755
rect 2158 2752 2159 2756
rect 2163 2752 2164 2756
rect 2158 2751 2164 2752
rect 2114 2750 2120 2751
rect 1994 2741 2000 2742
rect 1974 2740 1980 2741
rect 1974 2736 1975 2740
rect 1979 2736 1980 2740
rect 1994 2737 1995 2741
rect 1999 2737 2000 2741
rect 1994 2736 2000 2737
rect 1974 2735 1980 2736
rect 1934 2733 1940 2734
rect 1038 2732 1044 2733
rect 1038 2728 1039 2732
rect 1043 2728 1044 2732
rect 1038 2727 1044 2728
rect 1294 2732 1300 2733
rect 1566 2732 1572 2733
rect 1814 2732 1820 2733
rect 1294 2728 1295 2732
rect 1299 2728 1300 2732
rect 1294 2727 1300 2728
rect 1386 2731 1392 2732
rect 1386 2727 1387 2731
rect 1391 2727 1392 2731
rect 1566 2728 1567 2732
rect 1571 2728 1572 2732
rect 1566 2727 1572 2728
rect 1658 2731 1664 2732
rect 1658 2727 1659 2731
rect 1663 2727 1664 2731
rect 1814 2728 1815 2732
rect 1819 2728 1820 2732
rect 1814 2727 1820 2728
rect 1910 2731 1916 2732
rect 1910 2727 1911 2731
rect 1915 2727 1916 2731
rect 1934 2729 1935 2733
rect 1939 2729 1940 2733
rect 1934 2728 1940 2729
rect 1386 2726 1392 2727
rect 1658 2726 1664 2727
rect 1910 2726 1916 2727
rect 1010 2717 1016 2718
rect 1010 2713 1011 2717
rect 1015 2713 1016 2717
rect 1010 2712 1016 2713
rect 1266 2717 1272 2718
rect 1266 2713 1267 2717
rect 1271 2713 1272 2717
rect 1266 2712 1272 2713
rect 918 2667 924 2668
rect 918 2663 919 2667
rect 923 2663 924 2667
rect 918 2662 924 2663
rect 1012 2651 1014 2712
rect 1268 2651 1270 2712
rect 539 2650 543 2651
rect 539 2645 543 2646
rect 547 2650 551 2651
rect 547 2645 551 2646
rect 699 2650 703 2651
rect 699 2645 703 2646
rect 771 2650 775 2651
rect 771 2645 775 2646
rect 867 2650 871 2651
rect 867 2645 871 2646
rect 1011 2650 1015 2651
rect 1011 2645 1015 2646
rect 1035 2650 1039 2651
rect 1035 2645 1039 2646
rect 1203 2650 1207 2651
rect 1203 2645 1207 2646
rect 1267 2650 1271 2651
rect 1267 2645 1271 2646
rect 1371 2650 1375 2651
rect 1388 2648 1390 2726
rect 1538 2717 1544 2718
rect 1538 2713 1539 2717
rect 1543 2713 1544 2717
rect 1538 2712 1544 2713
rect 1540 2651 1542 2712
rect 1539 2650 1543 2651
rect 1371 2645 1375 2646
rect 1386 2647 1392 2648
rect 540 2584 542 2645
rect 662 2639 668 2640
rect 662 2635 663 2639
rect 667 2635 668 2639
rect 662 2634 668 2635
rect 634 2631 640 2632
rect 634 2627 635 2631
rect 639 2627 640 2631
rect 634 2626 640 2627
rect 538 2583 544 2584
rect 538 2579 539 2583
rect 543 2579 544 2583
rect 538 2578 544 2579
rect 566 2568 572 2569
rect 110 2567 116 2568
rect 110 2563 111 2567
rect 115 2563 116 2567
rect 414 2564 415 2568
rect 419 2564 420 2568
rect 414 2563 420 2564
rect 506 2567 512 2568
rect 506 2563 507 2567
rect 511 2563 512 2567
rect 566 2564 567 2568
rect 571 2564 572 2568
rect 566 2563 572 2564
rect 110 2562 116 2563
rect 112 2539 114 2562
rect 416 2539 418 2563
rect 506 2562 512 2563
rect 568 2539 570 2563
rect 111 2538 115 2539
rect 111 2533 115 2534
rect 327 2538 331 2539
rect 327 2533 331 2534
rect 415 2538 419 2539
rect 415 2533 419 2534
rect 535 2538 539 2539
rect 535 2533 539 2534
rect 567 2538 571 2539
rect 567 2533 571 2534
rect 112 2510 114 2533
rect 110 2509 116 2510
rect 328 2509 330 2533
rect 536 2509 538 2533
rect 110 2505 111 2509
rect 115 2505 116 2509
rect 110 2504 116 2505
rect 326 2508 332 2509
rect 534 2508 540 2509
rect 636 2508 638 2626
rect 664 2568 666 2634
rect 700 2584 702 2645
rect 854 2635 860 2636
rect 854 2631 855 2635
rect 859 2631 860 2635
rect 854 2630 860 2631
rect 698 2583 704 2584
rect 698 2579 699 2583
rect 703 2579 704 2583
rect 698 2578 704 2579
rect 856 2576 858 2630
rect 868 2584 870 2645
rect 1036 2584 1038 2645
rect 1158 2643 1164 2644
rect 1158 2639 1159 2643
rect 1163 2639 1164 2643
rect 1158 2638 1164 2639
rect 866 2583 872 2584
rect 866 2579 867 2583
rect 871 2579 872 2583
rect 866 2578 872 2579
rect 1034 2583 1040 2584
rect 1034 2579 1035 2583
rect 1039 2579 1040 2583
rect 1034 2578 1040 2579
rect 854 2575 860 2576
rect 854 2571 855 2575
rect 859 2571 860 2575
rect 854 2570 860 2571
rect 726 2568 732 2569
rect 894 2568 900 2569
rect 662 2567 668 2568
rect 662 2563 663 2567
rect 667 2563 668 2567
rect 726 2564 727 2568
rect 731 2564 732 2568
rect 726 2563 732 2564
rect 822 2567 828 2568
rect 822 2563 823 2567
rect 827 2563 828 2567
rect 894 2564 895 2568
rect 899 2564 900 2568
rect 894 2563 900 2564
rect 1062 2568 1068 2569
rect 1160 2568 1162 2638
rect 1204 2584 1206 2645
rect 1372 2584 1374 2645
rect 1386 2643 1387 2647
rect 1391 2643 1392 2647
rect 1539 2645 1543 2646
rect 1386 2642 1392 2643
rect 1494 2639 1500 2640
rect 1494 2635 1495 2639
rect 1499 2635 1500 2639
rect 1494 2634 1500 2635
rect 1466 2631 1472 2632
rect 1466 2627 1467 2631
rect 1471 2627 1472 2631
rect 1466 2626 1472 2627
rect 1468 2604 1470 2626
rect 1466 2603 1472 2604
rect 1466 2599 1467 2603
rect 1471 2599 1472 2603
rect 1466 2598 1472 2599
rect 1202 2583 1208 2584
rect 1202 2579 1203 2583
rect 1207 2579 1208 2583
rect 1202 2578 1208 2579
rect 1370 2583 1376 2584
rect 1370 2579 1371 2583
rect 1375 2579 1376 2583
rect 1370 2578 1376 2579
rect 1230 2568 1236 2569
rect 1398 2568 1404 2569
rect 1496 2568 1498 2634
rect 1540 2584 1542 2645
rect 1660 2636 1662 2726
rect 1786 2717 1792 2718
rect 1786 2713 1787 2717
rect 1791 2713 1792 2717
rect 1786 2712 1792 2713
rect 1788 2651 1790 2712
rect 1912 2660 1914 2726
rect 1934 2716 1940 2717
rect 1934 2712 1935 2716
rect 1939 2712 1940 2716
rect 1934 2711 1940 2712
rect 1910 2659 1916 2660
rect 1910 2655 1911 2659
rect 1915 2655 1916 2659
rect 1910 2654 1916 2655
rect 1936 2651 1938 2711
rect 1976 2667 1978 2735
rect 1996 2667 1998 2736
rect 2116 2668 2118 2750
rect 2130 2741 2136 2742
rect 2130 2737 2131 2741
rect 2135 2737 2136 2741
rect 2130 2736 2136 2737
rect 2114 2667 2120 2668
rect 2132 2667 2134 2736
rect 2252 2692 2254 2814
rect 2296 2787 2298 2815
rect 2410 2814 2416 2815
rect 2432 2787 2434 2815
rect 2546 2814 2552 2815
rect 2568 2787 2570 2815
rect 2662 2814 2668 2815
rect 2712 2787 2714 2815
rect 2295 2786 2299 2787
rect 2295 2781 2299 2782
rect 2303 2786 2307 2787
rect 2303 2781 2307 2782
rect 2431 2786 2435 2787
rect 2431 2781 2435 2782
rect 2463 2786 2467 2787
rect 2463 2781 2467 2782
rect 2567 2786 2571 2787
rect 2567 2781 2571 2782
rect 2623 2786 2627 2787
rect 2623 2781 2627 2782
rect 2711 2786 2715 2787
rect 2711 2781 2715 2782
rect 2304 2757 2306 2781
rect 2464 2757 2466 2781
rect 2624 2757 2626 2781
rect 2302 2756 2308 2757
rect 2462 2756 2468 2757
rect 2622 2756 2628 2757
rect 2720 2756 2722 2882
rect 2836 2836 2838 2897
rect 2842 2883 2848 2884
rect 2842 2879 2843 2883
rect 2847 2879 2848 2883
rect 2842 2878 2848 2879
rect 2834 2835 2840 2836
rect 2834 2831 2835 2835
rect 2839 2831 2840 2835
rect 2834 2830 2840 2831
rect 2844 2820 2846 2878
rect 2862 2820 2868 2821
rect 2960 2820 2962 2918
rect 3092 2903 3094 2968
rect 3308 2903 3310 2968
rect 2995 2902 2999 2903
rect 2995 2897 2999 2898
rect 3091 2902 3095 2903
rect 3091 2897 3095 2898
rect 3155 2902 3159 2903
rect 3155 2897 3159 2898
rect 3307 2902 3311 2903
rect 3307 2897 3311 2898
rect 3315 2902 3319 2903
rect 3315 2897 3319 2898
rect 2996 2836 2998 2897
rect 3146 2887 3152 2888
rect 3146 2883 3147 2887
rect 3151 2883 3152 2887
rect 3146 2882 3152 2883
rect 2994 2835 3000 2836
rect 2994 2831 2995 2835
rect 2999 2831 3000 2835
rect 2994 2830 3000 2831
rect 3148 2828 3150 2882
rect 3156 2836 3158 2897
rect 3306 2887 3312 2888
rect 3306 2883 3307 2887
rect 3311 2883 3312 2887
rect 3306 2882 3312 2883
rect 3154 2835 3160 2836
rect 3154 2831 3155 2835
rect 3159 2831 3160 2835
rect 3154 2830 3160 2831
rect 3308 2828 3310 2882
rect 3316 2836 3318 2897
rect 3428 2888 3430 2982
rect 3530 2973 3536 2974
rect 3530 2969 3531 2973
rect 3535 2969 3536 2973
rect 3530 2968 3536 2969
rect 3532 2903 3534 2968
rect 3652 2916 3654 2982
rect 3772 2924 3774 3050
rect 3800 3019 3802 3050
rect 3958 3040 3964 3041
rect 4052 3040 4054 3138
rect 4156 3123 4158 3188
rect 4412 3123 4414 3188
rect 4131 3122 4135 3123
rect 4131 3117 4135 3118
rect 4155 3122 4159 3123
rect 4155 3117 4159 3118
rect 4331 3122 4335 3123
rect 4331 3117 4335 3118
rect 4411 3122 4415 3123
rect 4411 3117 4415 3118
rect 4523 3122 4527 3123
rect 4523 3117 4527 3118
rect 4094 3107 4100 3108
rect 4094 3103 4095 3107
rect 4099 3103 4100 3107
rect 4094 3102 4100 3103
rect 3838 3039 3844 3040
rect 3838 3035 3839 3039
rect 3843 3035 3844 3039
rect 3958 3036 3959 3040
rect 3963 3036 3964 3040
rect 3958 3035 3964 3036
rect 4050 3039 4056 3040
rect 4050 3035 4051 3039
rect 4055 3035 4056 3039
rect 3838 3034 3844 3035
rect 3799 3018 3803 3019
rect 3799 3013 3803 3014
rect 3800 2990 3802 3013
rect 3798 2989 3804 2990
rect 3798 2985 3799 2989
rect 3803 2985 3804 2989
rect 3840 2987 3842 3034
rect 3960 2987 3962 3035
rect 4050 3034 4056 3035
rect 3798 2984 3804 2985
rect 3839 2986 3843 2987
rect 3839 2981 3843 2982
rect 3959 2986 3963 2987
rect 3959 2981 3963 2982
rect 3999 2986 4003 2987
rect 3999 2981 4003 2982
rect 3798 2972 3804 2973
rect 3798 2968 3799 2972
rect 3803 2968 3804 2972
rect 3798 2967 3804 2968
rect 3770 2923 3776 2924
rect 3770 2919 3771 2923
rect 3775 2919 3776 2923
rect 3770 2918 3776 2919
rect 3650 2915 3656 2916
rect 3650 2911 3651 2915
rect 3655 2911 3656 2915
rect 3650 2910 3656 2911
rect 3800 2903 3802 2967
rect 3840 2958 3842 2981
rect 3838 2957 3844 2958
rect 4000 2957 4002 2981
rect 3838 2953 3839 2957
rect 3843 2953 3844 2957
rect 3838 2952 3844 2953
rect 3998 2956 4004 2957
rect 4096 2956 4098 3102
rect 4132 3056 4134 3117
rect 4226 3103 4232 3104
rect 4226 3098 4227 3103
rect 4231 3098 4232 3103
rect 4227 3095 4231 3096
rect 4332 3056 4334 3117
rect 4338 3103 4344 3104
rect 4338 3099 4339 3103
rect 4343 3099 4344 3103
rect 4338 3098 4344 3099
rect 4130 3055 4136 3056
rect 4130 3051 4131 3055
rect 4135 3051 4136 3055
rect 4130 3050 4136 3051
rect 4330 3055 4336 3056
rect 4330 3051 4331 3055
rect 4335 3051 4336 3055
rect 4330 3050 4336 3051
rect 4158 3040 4164 3041
rect 4340 3040 4342 3098
rect 4524 3056 4526 3117
rect 4536 3108 4538 3202
rect 4658 3193 4664 3194
rect 4658 3189 4659 3193
rect 4663 3189 4664 3193
rect 4658 3188 4664 3189
rect 4660 3123 4662 3188
rect 4780 3136 4782 3202
rect 4820 3144 4822 3286
rect 4968 3239 4970 3287
rect 5058 3286 5064 3287
rect 5208 3239 5210 3287
rect 5302 3286 5308 3287
rect 5456 3239 5458 3287
rect 5662 3286 5668 3287
rect 5664 3239 5666 3286
rect 4935 3238 4939 3239
rect 4935 3233 4939 3234
rect 4967 3238 4971 3239
rect 4967 3233 4971 3234
rect 5191 3238 5195 3239
rect 5191 3233 5195 3234
rect 5207 3238 5211 3239
rect 5207 3233 5211 3234
rect 5455 3238 5459 3239
rect 5455 3233 5459 3234
rect 5663 3238 5667 3239
rect 5663 3233 5667 3234
rect 4936 3209 4938 3233
rect 5192 3209 5194 3233
rect 5664 3210 5666 3233
rect 5662 3209 5668 3210
rect 4934 3208 4940 3209
rect 5190 3208 5196 3209
rect 4934 3204 4935 3208
rect 4939 3204 4940 3208
rect 4934 3203 4940 3204
rect 5030 3207 5036 3208
rect 5030 3203 5031 3207
rect 5035 3203 5036 3207
rect 5190 3204 5191 3208
rect 5195 3204 5196 3208
rect 5190 3203 5196 3204
rect 5286 3207 5292 3208
rect 5286 3203 5287 3207
rect 5291 3203 5292 3207
rect 5662 3205 5663 3209
rect 5667 3205 5668 3209
rect 5662 3204 5668 3205
rect 5030 3202 5036 3203
rect 5286 3202 5292 3203
rect 4906 3193 4912 3194
rect 4906 3189 4907 3193
rect 4911 3189 4912 3193
rect 4906 3188 4912 3189
rect 4818 3143 4824 3144
rect 4818 3139 4819 3143
rect 4823 3139 4824 3143
rect 4818 3138 4824 3139
rect 4778 3135 4784 3136
rect 4778 3131 4779 3135
rect 4783 3131 4784 3135
rect 4778 3130 4784 3131
rect 4908 3123 4910 3188
rect 5032 3144 5034 3202
rect 5162 3193 5168 3194
rect 5162 3189 5163 3193
rect 5167 3189 5168 3193
rect 5162 3188 5168 3189
rect 5030 3143 5036 3144
rect 5030 3139 5031 3143
rect 5035 3139 5036 3143
rect 5030 3138 5036 3139
rect 5164 3123 5166 3188
rect 5288 3136 5290 3202
rect 5662 3192 5668 3193
rect 5662 3188 5663 3192
rect 5667 3188 5668 3192
rect 5662 3187 5668 3188
rect 5286 3135 5292 3136
rect 5286 3131 5287 3135
rect 5291 3131 5292 3135
rect 5286 3130 5292 3131
rect 5664 3123 5666 3187
rect 4659 3122 4663 3123
rect 4659 3117 4663 3118
rect 4715 3122 4719 3123
rect 4715 3117 4719 3118
rect 4907 3122 4911 3123
rect 4907 3117 4911 3118
rect 4915 3122 4919 3123
rect 4915 3117 4919 3118
rect 5163 3122 5167 3123
rect 5163 3117 5167 3118
rect 5663 3122 5667 3123
rect 5663 3117 5667 3118
rect 4534 3107 4540 3108
rect 4534 3103 4535 3107
rect 4539 3103 4540 3107
rect 4534 3102 4540 3103
rect 4716 3056 4718 3117
rect 4722 3103 4728 3104
rect 4722 3099 4723 3103
rect 4727 3099 4728 3103
rect 4722 3098 4728 3099
rect 4522 3055 4528 3056
rect 4522 3051 4523 3055
rect 4527 3051 4528 3055
rect 4522 3050 4528 3051
rect 4714 3055 4720 3056
rect 4714 3051 4715 3055
rect 4719 3051 4720 3055
rect 4714 3050 4720 3051
rect 4358 3040 4364 3041
rect 4550 3040 4556 3041
rect 4724 3040 4726 3098
rect 4916 3056 4918 3117
rect 4922 3103 4928 3104
rect 4922 3099 4923 3103
rect 4927 3099 4928 3103
rect 4922 3098 4928 3099
rect 5039 3100 5043 3101
rect 4914 3055 4920 3056
rect 4914 3051 4915 3055
rect 4919 3051 4920 3055
rect 4914 3050 4920 3051
rect 4742 3040 4748 3041
rect 4924 3040 4926 3098
rect 5039 3095 5043 3096
rect 4942 3040 4948 3041
rect 5040 3040 5042 3095
rect 5664 3057 5666 3117
rect 5662 3056 5668 3057
rect 5662 3052 5663 3056
rect 5667 3052 5668 3056
rect 5662 3051 5668 3052
rect 4158 3036 4159 3040
rect 4163 3036 4164 3040
rect 4158 3035 4164 3036
rect 4338 3039 4344 3040
rect 4338 3035 4339 3039
rect 4343 3035 4344 3039
rect 4358 3036 4359 3040
rect 4363 3036 4364 3040
rect 4358 3035 4364 3036
rect 4466 3039 4472 3040
rect 4466 3035 4467 3039
rect 4471 3035 4472 3039
rect 4550 3036 4551 3040
rect 4555 3036 4556 3040
rect 4550 3035 4556 3036
rect 4722 3039 4728 3040
rect 4722 3035 4723 3039
rect 4727 3035 4728 3039
rect 4742 3036 4743 3040
rect 4747 3036 4748 3040
rect 4742 3035 4748 3036
rect 4922 3039 4928 3040
rect 4922 3035 4923 3039
rect 4927 3035 4928 3039
rect 4942 3036 4943 3040
rect 4947 3036 4948 3040
rect 4942 3035 4948 3036
rect 5038 3039 5044 3040
rect 5038 3035 5039 3039
rect 5043 3035 5044 3039
rect 4160 2987 4162 3035
rect 4338 3034 4344 3035
rect 4360 2987 4362 3035
rect 4466 3034 4472 3035
rect 4159 2986 4163 2987
rect 4159 2981 4163 2982
rect 4335 2986 4339 2987
rect 4335 2981 4339 2982
rect 4359 2986 4363 2987
rect 4359 2981 4363 2982
rect 4160 2957 4162 2981
rect 4336 2957 4338 2981
rect 4158 2956 4164 2957
rect 3998 2952 3999 2956
rect 4003 2952 4004 2956
rect 3998 2951 4004 2952
rect 4094 2955 4100 2956
rect 4094 2951 4095 2955
rect 4099 2951 4100 2955
rect 4158 2952 4159 2956
rect 4163 2952 4164 2956
rect 4158 2951 4164 2952
rect 4334 2956 4340 2957
rect 4334 2952 4335 2956
rect 4339 2952 4340 2956
rect 4334 2951 4340 2952
rect 4442 2955 4448 2956
rect 4442 2951 4443 2955
rect 4447 2951 4448 2955
rect 4094 2950 4100 2951
rect 4442 2950 4448 2951
rect 3970 2941 3976 2942
rect 3838 2940 3844 2941
rect 3838 2936 3839 2940
rect 3843 2936 3844 2940
rect 3970 2937 3971 2941
rect 3975 2937 3976 2941
rect 3970 2936 3976 2937
rect 4130 2941 4136 2942
rect 4130 2937 4131 2941
rect 4135 2937 4136 2941
rect 4130 2936 4136 2937
rect 4306 2941 4312 2942
rect 4306 2937 4307 2941
rect 4311 2937 4312 2941
rect 4306 2936 4312 2937
rect 3838 2935 3844 2936
rect 3531 2902 3535 2903
rect 3531 2897 3535 2898
rect 3799 2902 3803 2903
rect 3799 2897 3803 2898
rect 3426 2887 3432 2888
rect 3426 2883 3427 2887
rect 3431 2883 3432 2887
rect 3426 2882 3432 2883
rect 3800 2837 3802 2897
rect 3840 2859 3842 2935
rect 3972 2859 3974 2936
rect 3982 2891 3988 2892
rect 3982 2887 3983 2891
rect 3987 2887 3988 2891
rect 3982 2886 3988 2887
rect 3839 2858 3843 2859
rect 3839 2853 3843 2854
rect 3859 2858 3863 2859
rect 3859 2853 3863 2854
rect 3971 2858 3975 2859
rect 3971 2853 3975 2854
rect 3798 2836 3804 2837
rect 3314 2835 3320 2836
rect 3314 2831 3315 2835
rect 3319 2831 3320 2835
rect 3798 2832 3799 2836
rect 3803 2832 3804 2836
rect 3798 2831 3804 2832
rect 3314 2830 3320 2831
rect 3146 2827 3152 2828
rect 3146 2823 3147 2827
rect 3151 2823 3152 2827
rect 3146 2822 3152 2823
rect 3306 2827 3312 2828
rect 3306 2823 3307 2827
rect 3311 2823 3312 2827
rect 3306 2822 3312 2823
rect 3022 2820 3028 2821
rect 3182 2820 3188 2821
rect 2842 2819 2848 2820
rect 2842 2815 2843 2819
rect 2847 2815 2848 2819
rect 2862 2816 2863 2820
rect 2867 2816 2868 2820
rect 2862 2815 2868 2816
rect 2958 2819 2964 2820
rect 2958 2815 2959 2819
rect 2963 2815 2964 2819
rect 3022 2816 3023 2820
rect 3027 2816 3028 2820
rect 3022 2815 3028 2816
rect 3118 2819 3124 2820
rect 3118 2815 3119 2819
rect 3123 2815 3124 2819
rect 3182 2816 3183 2820
rect 3187 2816 3188 2820
rect 3182 2815 3188 2816
rect 3342 2820 3348 2821
rect 3342 2816 3343 2820
rect 3347 2816 3348 2820
rect 3342 2815 3348 2816
rect 3798 2819 3804 2820
rect 3798 2815 3799 2819
rect 3803 2815 3804 2819
rect 2842 2814 2848 2815
rect 2864 2787 2866 2815
rect 2958 2814 2964 2815
rect 3024 2787 3026 2815
rect 3118 2814 3124 2815
rect 2783 2786 2787 2787
rect 2783 2781 2787 2782
rect 2863 2786 2867 2787
rect 2863 2781 2867 2782
rect 2943 2786 2947 2787
rect 2943 2781 2947 2782
rect 3023 2786 3027 2787
rect 3023 2781 3027 2782
rect 3103 2786 3107 2787
rect 3103 2781 3107 2782
rect 2784 2757 2786 2781
rect 2944 2757 2946 2781
rect 3104 2757 3106 2781
rect 2782 2756 2788 2757
rect 2942 2756 2948 2757
rect 3102 2756 3108 2757
rect 2258 2755 2264 2756
rect 2258 2751 2259 2755
rect 2263 2751 2264 2755
rect 2302 2752 2303 2756
rect 2307 2752 2308 2756
rect 2302 2751 2308 2752
rect 2402 2755 2408 2756
rect 2402 2751 2403 2755
rect 2407 2751 2408 2755
rect 2462 2752 2463 2756
rect 2467 2752 2468 2756
rect 2462 2751 2468 2752
rect 2558 2755 2564 2756
rect 2558 2751 2559 2755
rect 2563 2751 2564 2755
rect 2622 2752 2623 2756
rect 2627 2752 2628 2756
rect 2622 2751 2628 2752
rect 2718 2755 2724 2756
rect 2718 2751 2719 2755
rect 2723 2751 2724 2755
rect 2782 2752 2783 2756
rect 2787 2752 2788 2756
rect 2782 2751 2788 2752
rect 2874 2755 2880 2756
rect 2874 2751 2875 2755
rect 2879 2751 2880 2755
rect 2942 2752 2943 2756
rect 2947 2752 2948 2756
rect 2942 2751 2948 2752
rect 3034 2755 3040 2756
rect 3034 2751 3035 2755
rect 3039 2751 3040 2755
rect 3102 2752 3103 2756
rect 3107 2752 3108 2756
rect 3102 2751 3108 2752
rect 2258 2750 2264 2751
rect 2402 2750 2408 2751
rect 2558 2750 2564 2751
rect 2718 2750 2724 2751
rect 2874 2750 2880 2751
rect 3034 2750 3040 2751
rect 2260 2692 2262 2750
rect 2274 2741 2280 2742
rect 2274 2737 2275 2741
rect 2279 2737 2280 2741
rect 2274 2736 2280 2737
rect 2250 2691 2256 2692
rect 2250 2687 2251 2691
rect 2255 2687 2256 2691
rect 2250 2686 2256 2687
rect 2258 2691 2264 2692
rect 2258 2687 2259 2691
rect 2263 2687 2264 2691
rect 2258 2686 2264 2687
rect 2276 2667 2278 2736
rect 2404 2692 2406 2750
rect 2434 2741 2440 2742
rect 2434 2737 2435 2741
rect 2439 2737 2440 2741
rect 2434 2736 2440 2737
rect 2402 2691 2408 2692
rect 2402 2687 2403 2691
rect 2407 2687 2408 2691
rect 2402 2686 2408 2687
rect 2436 2667 2438 2736
rect 2560 2684 2562 2750
rect 2594 2741 2600 2742
rect 2594 2737 2595 2741
rect 2599 2737 2600 2741
rect 2594 2736 2600 2737
rect 2754 2741 2760 2742
rect 2754 2737 2755 2741
rect 2759 2737 2760 2741
rect 2754 2736 2760 2737
rect 2558 2683 2564 2684
rect 2558 2679 2559 2683
rect 2563 2679 2564 2683
rect 2558 2678 2564 2679
rect 2596 2667 2598 2736
rect 2756 2667 2758 2736
rect 2822 2691 2828 2692
rect 2822 2687 2823 2691
rect 2827 2687 2828 2691
rect 2822 2686 2828 2687
rect 1975 2666 1979 2667
rect 1975 2661 1979 2662
rect 1995 2666 1999 2667
rect 2114 2663 2115 2667
rect 2119 2663 2120 2667
rect 2114 2662 2120 2663
rect 2131 2666 2135 2667
rect 1995 2661 1999 2662
rect 2131 2661 2135 2662
rect 2275 2666 2279 2667
rect 2275 2661 2279 2662
rect 2435 2666 2439 2667
rect 2435 2661 2439 2662
rect 2595 2666 2599 2667
rect 2595 2661 2599 2662
rect 2699 2666 2703 2667
rect 2699 2661 2703 2662
rect 2755 2666 2759 2667
rect 2755 2661 2759 2662
rect 1715 2650 1719 2651
rect 1715 2645 1719 2646
rect 1787 2650 1791 2651
rect 1787 2645 1791 2646
rect 1935 2650 1939 2651
rect 1935 2645 1939 2646
rect 1658 2635 1664 2636
rect 1658 2631 1659 2635
rect 1663 2631 1664 2635
rect 1658 2630 1664 2631
rect 1716 2584 1718 2645
rect 1722 2631 1728 2632
rect 1722 2627 1723 2631
rect 1727 2627 1728 2631
rect 1722 2626 1728 2627
rect 1538 2583 1544 2584
rect 1538 2579 1539 2583
rect 1543 2579 1544 2583
rect 1538 2578 1544 2579
rect 1714 2583 1720 2584
rect 1714 2579 1715 2583
rect 1719 2579 1720 2583
rect 1714 2578 1720 2579
rect 1566 2568 1572 2569
rect 1724 2568 1726 2626
rect 1838 2603 1844 2604
rect 1838 2599 1839 2603
rect 1843 2599 1844 2603
rect 1838 2598 1844 2599
rect 1742 2568 1748 2569
rect 1840 2568 1842 2598
rect 1936 2585 1938 2645
rect 1976 2601 1978 2661
rect 1974 2600 1980 2601
rect 2700 2600 2702 2661
rect 2794 2647 2800 2648
rect 2794 2643 2795 2647
rect 2799 2643 2800 2647
rect 2794 2642 2800 2643
rect 1974 2596 1975 2600
rect 1979 2596 1980 2600
rect 1974 2595 1980 2596
rect 2698 2599 2704 2600
rect 2698 2595 2699 2599
rect 2703 2595 2704 2599
rect 2698 2594 2704 2595
rect 1934 2584 1940 2585
rect 2726 2584 2732 2585
rect 1934 2580 1935 2584
rect 1939 2580 1940 2584
rect 1934 2579 1940 2580
rect 1974 2583 1980 2584
rect 1974 2579 1975 2583
rect 1979 2579 1980 2583
rect 2726 2580 2727 2584
rect 2731 2580 2732 2584
rect 2726 2579 2732 2580
rect 1974 2578 1980 2579
rect 1062 2564 1063 2568
rect 1067 2564 1068 2568
rect 1062 2563 1068 2564
rect 1158 2567 1164 2568
rect 1158 2563 1159 2567
rect 1163 2563 1164 2567
rect 1230 2564 1231 2568
rect 1235 2564 1236 2568
rect 1230 2563 1236 2564
rect 1326 2567 1332 2568
rect 1326 2563 1327 2567
rect 1331 2563 1332 2567
rect 1398 2564 1399 2568
rect 1403 2564 1404 2568
rect 1398 2563 1404 2564
rect 1494 2567 1500 2568
rect 1494 2563 1495 2567
rect 1499 2563 1500 2567
rect 1566 2564 1567 2568
rect 1571 2564 1572 2568
rect 1566 2563 1572 2564
rect 1722 2567 1728 2568
rect 1722 2563 1723 2567
rect 1727 2563 1728 2567
rect 1742 2564 1743 2568
rect 1747 2564 1748 2568
rect 1742 2563 1748 2564
rect 1838 2567 1844 2568
rect 1838 2563 1839 2567
rect 1843 2563 1844 2567
rect 662 2562 668 2563
rect 728 2539 730 2563
rect 822 2562 828 2563
rect 727 2538 731 2539
rect 727 2533 731 2534
rect 735 2538 739 2539
rect 735 2533 739 2534
rect 736 2509 738 2533
rect 734 2508 740 2509
rect 326 2504 327 2508
rect 331 2504 332 2508
rect 326 2503 332 2504
rect 426 2507 432 2508
rect 426 2503 427 2507
rect 431 2503 432 2507
rect 534 2504 535 2508
rect 539 2504 540 2508
rect 534 2503 540 2504
rect 634 2507 640 2508
rect 634 2503 635 2507
rect 639 2503 640 2507
rect 734 2504 735 2508
rect 739 2504 740 2508
rect 734 2503 740 2504
rect 426 2502 432 2503
rect 634 2502 640 2503
rect 298 2493 304 2494
rect 110 2492 116 2493
rect 110 2488 111 2492
rect 115 2488 116 2492
rect 298 2489 299 2493
rect 303 2489 304 2493
rect 298 2488 304 2489
rect 110 2487 116 2488
rect 112 2423 114 2487
rect 300 2423 302 2488
rect 428 2444 430 2502
rect 506 2493 512 2494
rect 506 2489 507 2493
rect 511 2489 512 2493
rect 506 2488 512 2489
rect 706 2493 712 2494
rect 706 2489 707 2493
rect 711 2489 712 2493
rect 706 2488 712 2489
rect 426 2443 432 2444
rect 426 2439 427 2443
rect 431 2439 432 2443
rect 426 2438 432 2439
rect 508 2423 510 2488
rect 708 2423 710 2488
rect 824 2444 826 2562
rect 896 2539 898 2563
rect 1064 2539 1066 2563
rect 1158 2562 1164 2563
rect 1232 2539 1234 2563
rect 1326 2562 1332 2563
rect 895 2538 899 2539
rect 895 2533 899 2534
rect 919 2538 923 2539
rect 919 2533 923 2534
rect 1063 2538 1067 2539
rect 1063 2533 1067 2534
rect 1095 2538 1099 2539
rect 1095 2533 1099 2534
rect 1231 2538 1235 2539
rect 1231 2533 1235 2534
rect 1271 2538 1275 2539
rect 1271 2533 1275 2534
rect 920 2509 922 2533
rect 1096 2509 1098 2533
rect 1272 2509 1274 2533
rect 918 2508 924 2509
rect 1094 2508 1100 2509
rect 1270 2508 1276 2509
rect 918 2504 919 2508
rect 923 2504 924 2508
rect 918 2503 924 2504
rect 1030 2507 1036 2508
rect 1030 2503 1031 2507
rect 1035 2503 1036 2507
rect 1094 2504 1095 2508
rect 1099 2504 1100 2508
rect 1094 2503 1100 2504
rect 1186 2507 1192 2508
rect 1186 2503 1187 2507
rect 1191 2503 1192 2507
rect 1270 2504 1271 2508
rect 1275 2504 1276 2508
rect 1270 2503 1276 2504
rect 1030 2502 1036 2503
rect 1186 2502 1192 2503
rect 890 2493 896 2494
rect 890 2489 891 2493
rect 895 2489 896 2493
rect 890 2488 896 2489
rect 822 2443 828 2444
rect 822 2439 823 2443
rect 827 2439 828 2443
rect 822 2438 828 2439
rect 892 2423 894 2488
rect 1032 2444 1034 2502
rect 1066 2493 1072 2494
rect 1066 2489 1067 2493
rect 1071 2489 1072 2493
rect 1066 2488 1072 2489
rect 1030 2443 1036 2444
rect 1030 2439 1031 2443
rect 1035 2439 1036 2443
rect 1030 2438 1036 2439
rect 1068 2423 1070 2488
rect 111 2422 115 2423
rect 111 2417 115 2418
rect 131 2422 135 2423
rect 131 2417 135 2418
rect 299 2422 303 2423
rect 299 2417 303 2418
rect 403 2422 407 2423
rect 403 2417 407 2418
rect 507 2422 511 2423
rect 507 2417 511 2418
rect 691 2422 695 2423
rect 691 2417 695 2418
rect 707 2422 711 2423
rect 707 2417 711 2418
rect 891 2422 895 2423
rect 891 2417 895 2418
rect 971 2422 975 2423
rect 971 2417 975 2418
rect 1067 2422 1071 2423
rect 1067 2417 1071 2418
rect 112 2357 114 2417
rect 110 2356 116 2357
rect 132 2356 134 2417
rect 226 2403 232 2404
rect 226 2399 227 2403
rect 231 2399 232 2403
rect 226 2398 232 2399
rect 228 2376 230 2398
rect 226 2375 232 2376
rect 226 2371 227 2375
rect 231 2371 232 2375
rect 226 2370 232 2371
rect 404 2356 406 2417
rect 518 2407 524 2408
rect 518 2403 519 2407
rect 523 2403 524 2407
rect 518 2402 524 2403
rect 110 2352 111 2356
rect 115 2352 116 2356
rect 110 2351 116 2352
rect 130 2355 136 2356
rect 130 2351 131 2355
rect 135 2351 136 2355
rect 130 2350 136 2351
rect 402 2355 408 2356
rect 402 2351 403 2355
rect 407 2351 408 2355
rect 402 2350 408 2351
rect 158 2340 164 2341
rect 110 2339 116 2340
rect 110 2335 111 2339
rect 115 2335 116 2339
rect 158 2336 159 2340
rect 163 2336 164 2340
rect 158 2335 164 2336
rect 430 2340 436 2341
rect 430 2336 431 2340
rect 435 2336 436 2340
rect 430 2335 436 2336
rect 110 2334 116 2335
rect 112 2295 114 2334
rect 160 2295 162 2335
rect 432 2295 434 2335
rect 111 2294 115 2295
rect 111 2289 115 2290
rect 159 2294 163 2295
rect 159 2289 163 2290
rect 423 2294 427 2295
rect 423 2289 427 2290
rect 431 2294 435 2295
rect 431 2289 435 2290
rect 112 2266 114 2289
rect 110 2265 116 2266
rect 160 2265 162 2289
rect 424 2265 426 2289
rect 110 2261 111 2265
rect 115 2261 116 2265
rect 110 2260 116 2261
rect 158 2264 164 2265
rect 158 2260 159 2264
rect 163 2260 164 2264
rect 158 2259 164 2260
rect 422 2264 428 2265
rect 520 2264 522 2402
rect 692 2356 694 2417
rect 698 2403 704 2404
rect 698 2399 699 2403
rect 703 2399 704 2403
rect 698 2398 704 2399
rect 690 2355 696 2356
rect 690 2351 691 2355
rect 695 2351 696 2355
rect 690 2350 696 2351
rect 700 2340 702 2398
rect 814 2375 820 2376
rect 814 2371 815 2375
rect 819 2371 820 2375
rect 814 2370 820 2371
rect 718 2340 724 2341
rect 816 2340 818 2370
rect 972 2356 974 2417
rect 1188 2408 1190 2502
rect 1242 2493 1248 2494
rect 1242 2489 1243 2493
rect 1247 2489 1248 2493
rect 1242 2488 1248 2489
rect 1244 2423 1246 2488
rect 1328 2444 1330 2562
rect 1400 2539 1402 2563
rect 1494 2562 1500 2563
rect 1568 2539 1570 2563
rect 1722 2562 1728 2563
rect 1744 2539 1746 2563
rect 1838 2562 1844 2563
rect 1934 2567 1940 2568
rect 1934 2563 1935 2567
rect 1939 2563 1940 2567
rect 1934 2562 1940 2563
rect 1936 2539 1938 2562
rect 1976 2555 1978 2578
rect 2728 2555 2730 2579
rect 1975 2554 1979 2555
rect 1975 2549 1979 2550
rect 2607 2554 2611 2555
rect 2607 2549 2611 2550
rect 2727 2554 2731 2555
rect 2727 2549 2731 2550
rect 2759 2554 2763 2555
rect 2759 2549 2763 2550
rect 1399 2538 1403 2539
rect 1399 2533 1403 2534
rect 1439 2538 1443 2539
rect 1439 2533 1443 2534
rect 1567 2538 1571 2539
rect 1567 2533 1571 2534
rect 1607 2538 1611 2539
rect 1607 2533 1611 2534
rect 1743 2538 1747 2539
rect 1743 2533 1747 2534
rect 1775 2538 1779 2539
rect 1775 2533 1779 2534
rect 1935 2538 1939 2539
rect 1935 2533 1939 2534
rect 1440 2509 1442 2533
rect 1608 2509 1610 2533
rect 1776 2509 1778 2533
rect 1936 2510 1938 2533
rect 1976 2526 1978 2549
rect 1974 2525 1980 2526
rect 2608 2525 2610 2549
rect 2760 2525 2762 2549
rect 2796 2540 2798 2642
rect 2824 2584 2826 2686
rect 2876 2684 2878 2750
rect 2914 2741 2920 2742
rect 2914 2737 2915 2741
rect 2919 2737 2920 2741
rect 2914 2736 2920 2737
rect 2874 2683 2880 2684
rect 2874 2679 2875 2683
rect 2879 2679 2880 2683
rect 2874 2678 2880 2679
rect 2916 2667 2918 2736
rect 2835 2666 2839 2667
rect 2835 2661 2839 2662
rect 2915 2666 2919 2667
rect 2915 2661 2919 2662
rect 2971 2666 2975 2667
rect 2971 2661 2975 2662
rect 2836 2600 2838 2661
rect 2972 2600 2974 2661
rect 3036 2660 3038 2750
rect 3074 2741 3080 2742
rect 3074 2737 3075 2741
rect 3079 2737 3080 2741
rect 3074 2736 3080 2737
rect 3076 2667 3078 2736
rect 3120 2692 3122 2814
rect 3184 2787 3186 2815
rect 3344 2787 3346 2815
rect 3798 2814 3804 2815
rect 3800 2787 3802 2814
rect 3840 2793 3842 2853
rect 3838 2792 3844 2793
rect 3860 2792 3862 2853
rect 3954 2839 3960 2840
rect 3954 2835 3955 2839
rect 3959 2835 3960 2839
rect 3954 2834 3960 2835
rect 3838 2788 3839 2792
rect 3843 2788 3844 2792
rect 3838 2787 3844 2788
rect 3858 2791 3864 2792
rect 3858 2787 3859 2791
rect 3863 2787 3864 2791
rect 3183 2786 3187 2787
rect 3183 2781 3187 2782
rect 3343 2786 3347 2787
rect 3343 2781 3347 2782
rect 3799 2786 3803 2787
rect 3858 2786 3864 2787
rect 3799 2781 3803 2782
rect 3800 2758 3802 2781
rect 3886 2776 3892 2777
rect 3838 2775 3844 2776
rect 3838 2771 3839 2775
rect 3843 2771 3844 2775
rect 3886 2772 3887 2776
rect 3891 2772 3892 2776
rect 3886 2771 3892 2772
rect 3838 2770 3844 2771
rect 3798 2757 3804 2758
rect 3198 2755 3204 2756
rect 3198 2751 3199 2755
rect 3203 2751 3204 2755
rect 3798 2753 3799 2757
rect 3803 2753 3804 2757
rect 3798 2752 3804 2753
rect 3198 2750 3204 2751
rect 3118 2691 3124 2692
rect 3118 2687 3119 2691
rect 3123 2687 3124 2691
rect 3118 2686 3124 2687
rect 3200 2684 3202 2750
rect 3798 2740 3804 2741
rect 3798 2736 3799 2740
rect 3803 2736 3804 2740
rect 3798 2735 3804 2736
rect 3840 2735 3842 2770
rect 3888 2735 3890 2771
rect 3956 2744 3958 2834
rect 3984 2776 3986 2886
rect 4132 2859 4134 2936
rect 4308 2859 4310 2936
rect 4011 2858 4015 2859
rect 4011 2853 4015 2854
rect 4131 2858 4135 2859
rect 4131 2853 4135 2854
rect 4211 2858 4215 2859
rect 4211 2853 4215 2854
rect 4307 2858 4311 2859
rect 4307 2853 4311 2854
rect 4435 2858 4439 2859
rect 4435 2853 4439 2854
rect 4012 2792 4014 2853
rect 4202 2843 4208 2844
rect 4202 2839 4203 2843
rect 4207 2839 4208 2843
rect 4202 2838 4208 2839
rect 4010 2791 4016 2792
rect 4010 2787 4011 2791
rect 4015 2787 4016 2791
rect 4010 2786 4016 2787
rect 4204 2784 4206 2838
rect 4212 2792 4214 2853
rect 4436 2792 4438 2853
rect 4444 2844 4446 2950
rect 4468 2892 4470 3034
rect 4552 2987 4554 3035
rect 4722 3034 4728 3035
rect 4744 2987 4746 3035
rect 4922 3034 4928 3035
rect 4944 2987 4946 3035
rect 5038 3034 5044 3035
rect 5662 3039 5668 3040
rect 5662 3035 5663 3039
rect 5667 3035 5668 3039
rect 5662 3034 5668 3035
rect 5664 2987 5666 3034
rect 4519 2986 4523 2987
rect 4519 2981 4523 2982
rect 4551 2986 4555 2987
rect 4551 2981 4555 2982
rect 4719 2986 4723 2987
rect 4719 2981 4723 2982
rect 4743 2986 4747 2987
rect 4743 2981 4747 2982
rect 4927 2986 4931 2987
rect 4927 2981 4931 2982
rect 4943 2986 4947 2987
rect 4943 2981 4947 2982
rect 5135 2986 5139 2987
rect 5135 2981 5139 2982
rect 5351 2986 5355 2987
rect 5351 2981 5355 2982
rect 5543 2986 5547 2987
rect 5543 2981 5547 2982
rect 5663 2986 5667 2987
rect 5663 2981 5667 2982
rect 4520 2957 4522 2981
rect 4720 2957 4722 2981
rect 4928 2957 4930 2981
rect 5136 2957 5138 2981
rect 5352 2957 5354 2981
rect 5544 2957 5546 2981
rect 5664 2958 5666 2981
rect 5662 2957 5668 2958
rect 4518 2956 4524 2957
rect 4718 2956 4724 2957
rect 4926 2956 4932 2957
rect 5134 2956 5140 2957
rect 5350 2956 5356 2957
rect 5542 2956 5548 2957
rect 4518 2952 4519 2956
rect 4523 2952 4524 2956
rect 4518 2951 4524 2952
rect 4618 2955 4624 2956
rect 4618 2951 4619 2955
rect 4623 2951 4624 2955
rect 4718 2952 4719 2956
rect 4723 2952 4724 2956
rect 4718 2951 4724 2952
rect 4818 2955 4824 2956
rect 4818 2951 4819 2955
rect 4823 2951 4824 2955
rect 4926 2952 4927 2956
rect 4931 2952 4932 2956
rect 4926 2951 4932 2952
rect 5018 2955 5024 2956
rect 5018 2951 5019 2955
rect 5023 2951 5024 2955
rect 5134 2952 5135 2956
rect 5139 2952 5140 2956
rect 5134 2951 5140 2952
rect 5286 2955 5292 2956
rect 5286 2951 5287 2955
rect 5291 2951 5292 2955
rect 5350 2952 5351 2956
rect 5355 2952 5356 2956
rect 5350 2951 5356 2952
rect 5482 2955 5488 2956
rect 5482 2951 5483 2955
rect 5487 2951 5488 2955
rect 5542 2952 5543 2956
rect 5547 2952 5548 2956
rect 5542 2951 5548 2952
rect 5634 2955 5640 2956
rect 5634 2951 5635 2955
rect 5639 2951 5640 2955
rect 5662 2953 5663 2957
rect 5667 2953 5668 2957
rect 5662 2952 5668 2953
rect 4618 2950 4624 2951
rect 4818 2950 4824 2951
rect 5018 2950 5024 2951
rect 5286 2950 5292 2951
rect 5482 2950 5488 2951
rect 5634 2950 5640 2951
rect 4490 2941 4496 2942
rect 4490 2937 4491 2941
rect 4495 2937 4496 2941
rect 4490 2936 4496 2937
rect 4466 2891 4472 2892
rect 4466 2887 4467 2891
rect 4471 2887 4472 2891
rect 4466 2886 4472 2887
rect 4492 2859 4494 2936
rect 4620 2892 4622 2950
rect 4690 2941 4696 2942
rect 4690 2937 4691 2941
rect 4695 2937 4696 2941
rect 4690 2936 4696 2937
rect 4618 2891 4624 2892
rect 4618 2887 4619 2891
rect 4623 2887 4624 2891
rect 4618 2886 4624 2887
rect 4692 2859 4694 2936
rect 4820 2892 4822 2950
rect 4898 2941 4904 2942
rect 4898 2937 4899 2941
rect 4903 2937 4904 2941
rect 4898 2936 4904 2937
rect 4818 2891 4824 2892
rect 4818 2887 4819 2891
rect 4823 2887 4824 2891
rect 4818 2886 4824 2887
rect 4900 2859 4902 2936
rect 5020 2884 5022 2950
rect 5106 2941 5112 2942
rect 5106 2937 5107 2941
rect 5111 2937 5112 2941
rect 5106 2936 5112 2937
rect 5018 2883 5024 2884
rect 5018 2879 5019 2883
rect 5023 2879 5024 2883
rect 5018 2878 5024 2879
rect 5108 2859 5110 2936
rect 5288 2892 5290 2950
rect 5322 2941 5328 2942
rect 5322 2937 5323 2941
rect 5327 2937 5328 2941
rect 5322 2936 5328 2937
rect 5286 2891 5292 2892
rect 5286 2887 5287 2891
rect 5291 2887 5292 2891
rect 5286 2886 5292 2887
rect 5324 2859 5326 2936
rect 5484 2892 5486 2950
rect 5514 2941 5520 2942
rect 5514 2937 5515 2941
rect 5519 2937 5520 2941
rect 5514 2936 5520 2937
rect 5482 2891 5488 2892
rect 5482 2887 5483 2891
rect 5487 2887 5488 2891
rect 5482 2886 5488 2887
rect 5374 2883 5380 2884
rect 5374 2879 5375 2883
rect 5379 2879 5380 2883
rect 5374 2878 5380 2879
rect 4491 2858 4495 2859
rect 4491 2853 4495 2854
rect 4691 2858 4695 2859
rect 4691 2853 4695 2854
rect 4899 2858 4903 2859
rect 4899 2853 4903 2854
rect 4963 2858 4967 2859
rect 4963 2853 4967 2854
rect 5107 2858 5111 2859
rect 5107 2853 5111 2854
rect 5251 2858 5255 2859
rect 5251 2853 5255 2854
rect 5323 2858 5327 2859
rect 5323 2853 5327 2854
rect 4442 2843 4448 2844
rect 4442 2839 4443 2843
rect 4447 2839 4448 2843
rect 4442 2838 4448 2839
rect 4692 2792 4694 2853
rect 4698 2839 4704 2840
rect 4698 2835 4699 2839
rect 4703 2835 4704 2839
rect 4698 2834 4704 2835
rect 4210 2791 4216 2792
rect 4210 2787 4211 2791
rect 4215 2787 4216 2791
rect 4210 2786 4216 2787
rect 4434 2791 4440 2792
rect 4434 2787 4435 2791
rect 4439 2787 4440 2791
rect 4434 2786 4440 2787
rect 4690 2791 4696 2792
rect 4690 2787 4691 2791
rect 4695 2787 4696 2791
rect 4690 2786 4696 2787
rect 4202 2783 4208 2784
rect 4202 2779 4203 2783
rect 4207 2779 4208 2783
rect 4202 2778 4208 2779
rect 4038 2776 4044 2777
rect 3982 2775 3988 2776
rect 3982 2771 3983 2775
rect 3987 2771 3988 2775
rect 4038 2772 4039 2776
rect 4043 2772 4044 2776
rect 4038 2771 4044 2772
rect 4238 2776 4244 2777
rect 4238 2772 4239 2776
rect 4243 2772 4244 2776
rect 4238 2771 4244 2772
rect 4462 2776 4468 2777
rect 4700 2776 4702 2834
rect 4964 2792 4966 2853
rect 4970 2839 4976 2840
rect 4970 2835 4971 2839
rect 4975 2835 4976 2839
rect 4970 2834 4976 2835
rect 4962 2791 4968 2792
rect 4962 2787 4963 2791
rect 4967 2787 4968 2791
rect 4962 2786 4968 2787
rect 4718 2776 4724 2777
rect 4972 2776 4974 2834
rect 5252 2792 5254 2853
rect 5250 2791 5256 2792
rect 5250 2787 5251 2791
rect 5255 2787 5256 2791
rect 5250 2786 5256 2787
rect 4990 2776 4996 2777
rect 4462 2772 4463 2776
rect 4467 2772 4468 2776
rect 4462 2771 4468 2772
rect 4698 2775 4704 2776
rect 4698 2771 4699 2775
rect 4703 2771 4704 2775
rect 4718 2772 4719 2776
rect 4723 2772 4724 2776
rect 4718 2771 4724 2772
rect 4970 2775 4976 2776
rect 4970 2771 4971 2775
rect 4975 2771 4976 2775
rect 4990 2772 4991 2776
rect 4995 2772 4996 2776
rect 4990 2771 4996 2772
rect 5278 2776 5284 2777
rect 5376 2776 5378 2878
rect 5516 2859 5518 2936
rect 5515 2858 5519 2859
rect 5515 2853 5519 2854
rect 5390 2843 5396 2844
rect 5390 2839 5391 2843
rect 5395 2839 5396 2843
rect 5390 2838 5396 2839
rect 5278 2772 5279 2776
rect 5283 2772 5284 2776
rect 5278 2771 5284 2772
rect 5374 2775 5380 2776
rect 5374 2771 5375 2775
rect 5379 2771 5380 2775
rect 3982 2770 3988 2771
rect 3954 2743 3960 2744
rect 3954 2739 3955 2743
rect 3959 2739 3960 2743
rect 3954 2738 3960 2739
rect 4040 2735 4042 2771
rect 4062 2743 4068 2744
rect 4062 2739 4063 2743
rect 4067 2739 4068 2743
rect 4062 2738 4068 2739
rect 3198 2683 3204 2684
rect 3198 2679 3199 2683
rect 3203 2679 3204 2683
rect 3198 2678 3204 2679
rect 3800 2667 3802 2735
rect 3839 2734 3843 2735
rect 3839 2729 3843 2730
rect 3887 2734 3891 2735
rect 3887 2729 3891 2730
rect 3967 2734 3971 2735
rect 3967 2729 3971 2730
rect 4039 2734 4043 2735
rect 4039 2729 4043 2730
rect 3840 2706 3842 2729
rect 3838 2705 3844 2706
rect 3968 2705 3970 2729
rect 3838 2701 3839 2705
rect 3843 2701 3844 2705
rect 3838 2700 3844 2701
rect 3966 2704 3972 2705
rect 4064 2704 4066 2738
rect 4240 2735 4242 2771
rect 4464 2735 4466 2771
rect 4698 2770 4704 2771
rect 4720 2735 4722 2771
rect 4970 2770 4976 2771
rect 4992 2735 4994 2771
rect 5280 2735 5282 2771
rect 5374 2770 5380 2771
rect 4223 2734 4227 2735
rect 4223 2729 4227 2730
rect 4239 2734 4243 2735
rect 4239 2729 4243 2730
rect 4463 2734 4467 2735
rect 4463 2729 4467 2730
rect 4527 2734 4531 2735
rect 4527 2729 4531 2730
rect 4719 2734 4723 2735
rect 4719 2729 4723 2730
rect 4863 2734 4867 2735
rect 4863 2729 4867 2730
rect 4991 2734 4995 2735
rect 4991 2729 4995 2730
rect 5215 2734 5219 2735
rect 5215 2729 5219 2730
rect 5279 2734 5283 2735
rect 5279 2729 5283 2730
rect 4224 2705 4226 2729
rect 4362 2719 4368 2720
rect 4362 2715 4363 2719
rect 4367 2715 4368 2719
rect 4362 2714 4368 2715
rect 4222 2704 4228 2705
rect 3966 2700 3967 2704
rect 3971 2700 3972 2704
rect 3966 2699 3972 2700
rect 4062 2703 4068 2704
rect 4062 2699 4063 2703
rect 4067 2699 4068 2703
rect 4222 2700 4223 2704
rect 4227 2700 4228 2704
rect 4222 2699 4228 2700
rect 4062 2698 4068 2699
rect 3938 2689 3944 2690
rect 3838 2688 3844 2689
rect 3838 2684 3839 2688
rect 3843 2684 3844 2688
rect 3938 2685 3939 2689
rect 3943 2685 3944 2689
rect 3938 2684 3944 2685
rect 4194 2689 4200 2690
rect 4194 2685 4195 2689
rect 4199 2685 4200 2689
rect 4194 2684 4200 2685
rect 3838 2683 3844 2684
rect 3075 2666 3079 2667
rect 3075 2661 3079 2662
rect 3799 2666 3803 2667
rect 3799 2661 3803 2662
rect 3034 2659 3040 2660
rect 3034 2655 3035 2659
rect 3039 2655 3040 2659
rect 3034 2654 3040 2655
rect 2978 2647 2984 2648
rect 2978 2643 2979 2647
rect 2983 2643 2984 2647
rect 2978 2642 2984 2643
rect 2834 2599 2840 2600
rect 2834 2595 2835 2599
rect 2839 2595 2840 2599
rect 2834 2594 2840 2595
rect 2970 2599 2976 2600
rect 2970 2595 2971 2599
rect 2975 2595 2976 2599
rect 2970 2594 2976 2595
rect 2862 2584 2868 2585
rect 2980 2584 2982 2642
rect 3800 2601 3802 2661
rect 3840 2623 3842 2683
rect 3940 2623 3942 2684
rect 4186 2631 4192 2632
rect 4186 2627 4187 2631
rect 4191 2627 4192 2631
rect 4186 2626 4192 2627
rect 3839 2622 3843 2623
rect 3839 2617 3843 2618
rect 3891 2622 3895 2623
rect 3891 2617 3895 2618
rect 3939 2622 3943 2623
rect 3939 2617 3943 2618
rect 4067 2622 4071 2623
rect 4067 2617 4071 2618
rect 3798 2600 3804 2601
rect 3798 2596 3799 2600
rect 3803 2596 3804 2600
rect 3798 2595 3804 2596
rect 2998 2584 3004 2585
rect 2822 2583 2828 2584
rect 2822 2579 2823 2583
rect 2827 2579 2828 2583
rect 2862 2580 2863 2584
rect 2867 2580 2868 2584
rect 2862 2579 2868 2580
rect 2978 2583 2984 2584
rect 2978 2579 2979 2583
rect 2983 2579 2984 2583
rect 2998 2580 2999 2584
rect 3003 2580 3004 2584
rect 2998 2579 3004 2580
rect 3094 2583 3100 2584
rect 3094 2579 3095 2583
rect 3099 2579 3100 2583
rect 2822 2578 2828 2579
rect 2864 2555 2866 2579
rect 2978 2578 2984 2579
rect 3000 2555 3002 2579
rect 3094 2578 3100 2579
rect 3798 2583 3804 2584
rect 3798 2579 3799 2583
rect 3803 2579 3804 2583
rect 3798 2578 3804 2579
rect 2863 2554 2867 2555
rect 2863 2549 2867 2550
rect 2911 2554 2915 2555
rect 2911 2549 2915 2550
rect 2999 2554 3003 2555
rect 2999 2549 3003 2550
rect 3063 2554 3067 2555
rect 3063 2549 3067 2550
rect 2794 2539 2800 2540
rect 2794 2535 2795 2539
rect 2799 2535 2800 2539
rect 2794 2534 2800 2535
rect 2912 2525 2914 2549
rect 3064 2525 3066 2549
rect 1974 2521 1975 2525
rect 1979 2521 1980 2525
rect 1974 2520 1980 2521
rect 2606 2524 2612 2525
rect 2758 2524 2764 2525
rect 2606 2520 2607 2524
rect 2611 2520 2612 2524
rect 2606 2519 2612 2520
rect 2702 2523 2708 2524
rect 2702 2519 2703 2523
rect 2707 2519 2708 2523
rect 2758 2520 2759 2524
rect 2763 2520 2764 2524
rect 2758 2519 2764 2520
rect 2910 2524 2916 2525
rect 3062 2524 3068 2525
rect 2910 2520 2911 2524
rect 2915 2520 2916 2524
rect 2910 2519 2916 2520
rect 3002 2523 3008 2524
rect 3002 2519 3003 2523
rect 3007 2519 3008 2523
rect 3062 2520 3063 2524
rect 3067 2520 3068 2524
rect 3062 2519 3068 2520
rect 2702 2518 2708 2519
rect 3002 2518 3008 2519
rect 1934 2509 1940 2510
rect 2578 2509 2584 2510
rect 1438 2508 1444 2509
rect 1606 2508 1612 2509
rect 1774 2508 1780 2509
rect 1370 2507 1376 2508
rect 1370 2503 1371 2507
rect 1375 2503 1376 2507
rect 1438 2504 1439 2508
rect 1443 2504 1444 2508
rect 1438 2503 1444 2504
rect 1538 2507 1544 2508
rect 1538 2503 1539 2507
rect 1543 2503 1544 2507
rect 1606 2504 1607 2508
rect 1611 2504 1612 2508
rect 1606 2503 1612 2504
rect 1706 2507 1712 2508
rect 1706 2503 1707 2507
rect 1711 2503 1712 2507
rect 1774 2504 1775 2508
rect 1779 2504 1780 2508
rect 1774 2503 1780 2504
rect 1866 2507 1872 2508
rect 1866 2503 1867 2507
rect 1871 2503 1872 2507
rect 1934 2505 1935 2509
rect 1939 2505 1940 2509
rect 1934 2504 1940 2505
rect 1974 2508 1980 2509
rect 1974 2504 1975 2508
rect 1979 2504 1980 2508
rect 2578 2505 2579 2509
rect 2583 2505 2584 2509
rect 2578 2504 2584 2505
rect 1974 2503 1980 2504
rect 1370 2502 1376 2503
rect 1538 2502 1544 2503
rect 1706 2502 1712 2503
rect 1866 2502 1872 2503
rect 1372 2444 1374 2502
rect 1410 2493 1416 2494
rect 1410 2489 1411 2493
rect 1415 2489 1416 2493
rect 1410 2488 1416 2489
rect 1326 2443 1332 2444
rect 1326 2439 1327 2443
rect 1331 2439 1332 2443
rect 1326 2438 1332 2439
rect 1370 2443 1376 2444
rect 1370 2439 1371 2443
rect 1375 2439 1376 2443
rect 1370 2438 1376 2439
rect 1412 2423 1414 2488
rect 1540 2444 1542 2502
rect 1578 2493 1584 2494
rect 1578 2489 1579 2493
rect 1583 2489 1584 2493
rect 1578 2488 1584 2489
rect 1538 2443 1544 2444
rect 1538 2439 1539 2443
rect 1543 2439 1544 2443
rect 1538 2438 1544 2439
rect 1580 2423 1582 2488
rect 1708 2444 1710 2502
rect 1746 2493 1752 2494
rect 1746 2489 1747 2493
rect 1751 2489 1752 2493
rect 1746 2488 1752 2489
rect 1706 2443 1712 2444
rect 1706 2439 1707 2443
rect 1711 2439 1712 2443
rect 1706 2438 1712 2439
rect 1748 2423 1750 2488
rect 1243 2422 1247 2423
rect 1243 2417 1247 2418
rect 1251 2422 1255 2423
rect 1251 2417 1255 2418
rect 1411 2422 1415 2423
rect 1411 2417 1415 2418
rect 1531 2422 1535 2423
rect 1531 2417 1535 2418
rect 1579 2422 1583 2423
rect 1579 2417 1583 2418
rect 1747 2422 1751 2423
rect 1747 2417 1751 2418
rect 1787 2422 1791 2423
rect 1787 2417 1791 2418
rect 1186 2407 1192 2408
rect 1186 2403 1187 2407
rect 1191 2403 1192 2407
rect 1186 2402 1192 2403
rect 1252 2356 1254 2417
rect 1258 2403 1264 2404
rect 1258 2399 1259 2403
rect 1263 2399 1264 2403
rect 1258 2398 1264 2399
rect 970 2355 976 2356
rect 970 2351 971 2355
rect 975 2351 976 2355
rect 970 2350 976 2351
rect 1250 2355 1256 2356
rect 1250 2351 1251 2355
rect 1255 2351 1256 2355
rect 1250 2350 1256 2351
rect 998 2340 1004 2341
rect 1260 2340 1262 2398
rect 1532 2356 1534 2417
rect 1788 2356 1790 2417
rect 1868 2416 1870 2502
rect 1934 2492 1940 2493
rect 1934 2488 1935 2492
rect 1939 2488 1940 2492
rect 1934 2487 1940 2488
rect 1936 2423 1938 2487
rect 1976 2427 1978 2503
rect 2580 2427 2582 2504
rect 2704 2460 2706 2518
rect 2730 2509 2736 2510
rect 2730 2505 2731 2509
rect 2735 2505 2736 2509
rect 2730 2504 2736 2505
rect 2882 2509 2888 2510
rect 2882 2505 2883 2509
rect 2887 2505 2888 2509
rect 2882 2504 2888 2505
rect 2690 2459 2696 2460
rect 2690 2455 2691 2459
rect 2695 2455 2696 2459
rect 2690 2454 2696 2455
rect 2702 2459 2708 2460
rect 2702 2455 2703 2459
rect 2707 2455 2708 2459
rect 2702 2454 2708 2455
rect 1975 2426 1979 2427
rect 1935 2422 1939 2423
rect 1975 2421 1979 2422
rect 1995 2426 1999 2427
rect 1995 2421 1999 2422
rect 2275 2426 2279 2427
rect 2275 2421 2279 2422
rect 2571 2426 2575 2427
rect 2571 2421 2575 2422
rect 2579 2426 2583 2427
rect 2579 2421 2583 2422
rect 1935 2417 1939 2418
rect 1866 2415 1872 2416
rect 1866 2411 1867 2415
rect 1871 2411 1872 2415
rect 1866 2410 1872 2411
rect 1914 2411 1920 2412
rect 1914 2407 1915 2411
rect 1919 2407 1920 2411
rect 1914 2406 1920 2407
rect 1794 2403 1800 2404
rect 1794 2399 1795 2403
rect 1799 2399 1800 2403
rect 1794 2398 1800 2399
rect 1530 2355 1536 2356
rect 1530 2351 1531 2355
rect 1535 2351 1536 2355
rect 1530 2350 1536 2351
rect 1786 2355 1792 2356
rect 1786 2351 1787 2355
rect 1791 2351 1792 2355
rect 1786 2350 1792 2351
rect 1278 2340 1284 2341
rect 1558 2340 1564 2341
rect 1796 2340 1798 2398
rect 1814 2340 1820 2341
rect 1916 2340 1918 2406
rect 1936 2357 1938 2417
rect 1976 2361 1978 2421
rect 1974 2360 1980 2361
rect 1996 2360 1998 2421
rect 2276 2360 2278 2421
rect 2572 2360 2574 2421
rect 2578 2407 2584 2408
rect 2578 2403 2579 2407
rect 2583 2403 2584 2407
rect 2578 2402 2584 2403
rect 1934 2356 1940 2357
rect 1934 2352 1935 2356
rect 1939 2352 1940 2356
rect 1974 2356 1975 2360
rect 1979 2356 1980 2360
rect 1974 2355 1980 2356
rect 1994 2359 2000 2360
rect 1994 2355 1995 2359
rect 1999 2355 2000 2359
rect 1994 2354 2000 2355
rect 2274 2359 2280 2360
rect 2274 2355 2275 2359
rect 2279 2355 2280 2359
rect 2274 2354 2280 2355
rect 2570 2359 2576 2360
rect 2570 2355 2571 2359
rect 2575 2355 2576 2359
rect 2570 2354 2576 2355
rect 1934 2351 1940 2352
rect 2022 2344 2028 2345
rect 2302 2344 2308 2345
rect 2580 2344 2582 2402
rect 2598 2344 2604 2345
rect 2692 2344 2694 2454
rect 2732 2427 2734 2504
rect 2884 2427 2886 2504
rect 2731 2426 2735 2427
rect 2731 2421 2735 2422
rect 2859 2426 2863 2427
rect 2859 2421 2863 2422
rect 2883 2426 2887 2427
rect 2883 2421 2887 2422
rect 2702 2415 2708 2416
rect 2702 2411 2703 2415
rect 2707 2411 2708 2415
rect 2702 2410 2708 2411
rect 1974 2343 1980 2344
rect 698 2339 704 2340
rect 698 2335 699 2339
rect 703 2335 704 2339
rect 718 2336 719 2340
rect 723 2336 724 2340
rect 718 2335 724 2336
rect 814 2339 820 2340
rect 814 2335 815 2339
rect 819 2335 820 2339
rect 998 2336 999 2340
rect 1003 2336 1004 2340
rect 998 2335 1004 2336
rect 1258 2339 1264 2340
rect 1258 2335 1259 2339
rect 1263 2335 1264 2339
rect 1278 2336 1279 2340
rect 1283 2336 1284 2340
rect 1278 2335 1284 2336
rect 1374 2339 1380 2340
rect 1374 2335 1375 2339
rect 1379 2335 1380 2339
rect 1558 2336 1559 2340
rect 1563 2336 1564 2340
rect 1558 2335 1564 2336
rect 1794 2339 1800 2340
rect 1794 2335 1795 2339
rect 1799 2335 1800 2339
rect 1814 2336 1815 2340
rect 1819 2336 1820 2340
rect 1814 2335 1820 2336
rect 1914 2339 1920 2340
rect 1914 2335 1915 2339
rect 1919 2335 1920 2339
rect 698 2334 704 2335
rect 720 2295 722 2335
rect 814 2334 820 2335
rect 1000 2295 1002 2335
rect 1258 2334 1264 2335
rect 1280 2295 1282 2335
rect 1374 2334 1380 2335
rect 711 2294 715 2295
rect 711 2289 715 2290
rect 719 2294 723 2295
rect 719 2289 723 2290
rect 999 2294 1003 2295
rect 999 2289 1003 2290
rect 1279 2294 1283 2295
rect 1279 2289 1283 2290
rect 1295 2294 1299 2295
rect 1295 2289 1299 2290
rect 712 2265 714 2289
rect 1000 2265 1002 2289
rect 1296 2265 1298 2289
rect 710 2264 716 2265
rect 998 2264 1004 2265
rect 1294 2264 1300 2265
rect 422 2260 423 2264
rect 427 2260 428 2264
rect 422 2259 428 2260
rect 518 2263 524 2264
rect 518 2259 519 2263
rect 523 2259 524 2263
rect 710 2260 711 2264
rect 715 2260 716 2264
rect 710 2259 716 2260
rect 810 2263 816 2264
rect 810 2259 811 2263
rect 815 2259 816 2263
rect 998 2260 999 2264
rect 1003 2260 1004 2264
rect 998 2259 1004 2260
rect 1094 2263 1100 2264
rect 1094 2259 1095 2263
rect 1099 2259 1100 2263
rect 1294 2260 1295 2264
rect 1299 2260 1300 2264
rect 1294 2259 1300 2260
rect 518 2258 524 2259
rect 810 2258 816 2259
rect 1094 2258 1100 2259
rect 130 2249 136 2250
rect 110 2248 116 2249
rect 110 2244 111 2248
rect 115 2244 116 2248
rect 130 2245 131 2249
rect 135 2245 136 2249
rect 130 2244 136 2245
rect 394 2249 400 2250
rect 394 2245 395 2249
rect 399 2245 400 2249
rect 394 2244 400 2245
rect 682 2249 688 2250
rect 682 2245 683 2249
rect 687 2245 688 2249
rect 682 2244 688 2245
rect 110 2243 116 2244
rect 112 2171 114 2243
rect 132 2171 134 2244
rect 250 2199 256 2200
rect 250 2195 251 2199
rect 255 2195 256 2199
rect 250 2194 256 2195
rect 111 2170 115 2171
rect 111 2165 115 2166
rect 131 2170 135 2171
rect 131 2165 135 2166
rect 112 2105 114 2165
rect 110 2104 116 2105
rect 132 2104 134 2165
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 130 2103 136 2104
rect 130 2099 131 2103
rect 135 2099 136 2103
rect 130 2098 136 2099
rect 158 2088 164 2089
rect 252 2088 254 2194
rect 396 2171 398 2244
rect 684 2171 686 2244
rect 812 2200 814 2258
rect 970 2249 976 2250
rect 970 2245 971 2249
rect 975 2245 976 2249
rect 970 2244 976 2245
rect 810 2199 816 2200
rect 810 2195 811 2199
rect 815 2195 816 2199
rect 810 2194 816 2195
rect 972 2171 974 2244
rect 395 2170 399 2171
rect 395 2165 399 2166
rect 403 2170 407 2171
rect 403 2165 407 2166
rect 683 2170 687 2171
rect 683 2165 687 2166
rect 731 2170 735 2171
rect 731 2165 735 2166
rect 971 2170 975 2171
rect 971 2165 975 2166
rect 1083 2170 1087 2171
rect 1083 2165 1087 2166
rect 404 2104 406 2165
rect 526 2159 532 2160
rect 526 2155 527 2159
rect 531 2155 532 2159
rect 526 2154 532 2155
rect 498 2151 504 2152
rect 498 2147 499 2151
rect 503 2147 504 2151
rect 498 2146 504 2147
rect 500 2116 502 2146
rect 498 2115 504 2116
rect 498 2111 499 2115
rect 503 2111 504 2115
rect 498 2110 504 2111
rect 402 2103 408 2104
rect 402 2099 403 2103
rect 407 2099 408 2103
rect 402 2098 408 2099
rect 430 2088 436 2089
rect 528 2088 530 2154
rect 732 2104 734 2165
rect 738 2151 744 2152
rect 738 2147 739 2151
rect 743 2147 744 2151
rect 738 2146 744 2147
rect 730 2103 736 2104
rect 730 2099 731 2103
rect 735 2099 736 2103
rect 730 2098 736 2099
rect 110 2087 116 2088
rect 110 2083 111 2087
rect 115 2083 116 2087
rect 158 2084 159 2088
rect 163 2084 164 2088
rect 158 2083 164 2084
rect 250 2087 256 2088
rect 250 2083 251 2087
rect 255 2083 256 2087
rect 430 2084 431 2088
rect 435 2084 436 2088
rect 430 2083 436 2084
rect 526 2087 532 2088
rect 526 2083 527 2087
rect 531 2083 532 2087
rect 110 2082 116 2083
rect 112 2055 114 2082
rect 160 2055 162 2083
rect 250 2082 256 2083
rect 432 2055 434 2083
rect 526 2082 532 2083
rect 111 2054 115 2055
rect 111 2049 115 2050
rect 159 2054 163 2055
rect 159 2049 163 2050
rect 223 2054 227 2055
rect 223 2049 227 2050
rect 383 2054 387 2055
rect 383 2049 387 2050
rect 431 2054 435 2055
rect 431 2049 435 2050
rect 559 2054 563 2055
rect 559 2049 563 2050
rect 112 2026 114 2049
rect 110 2025 116 2026
rect 224 2025 226 2049
rect 384 2025 386 2049
rect 560 2025 562 2049
rect 110 2021 111 2025
rect 115 2021 116 2025
rect 110 2020 116 2021
rect 222 2024 228 2025
rect 382 2024 388 2025
rect 222 2020 223 2024
rect 227 2020 228 2024
rect 222 2019 228 2020
rect 322 2023 328 2024
rect 322 2019 323 2023
rect 327 2019 328 2023
rect 382 2020 383 2024
rect 387 2020 388 2024
rect 382 2019 388 2020
rect 558 2024 564 2025
rect 740 2024 742 2146
rect 854 2115 860 2116
rect 854 2111 855 2115
rect 859 2111 860 2115
rect 854 2110 860 2111
rect 758 2088 764 2089
rect 856 2088 858 2110
rect 1084 2104 1086 2165
rect 1096 2156 1098 2258
rect 1266 2249 1272 2250
rect 1266 2245 1267 2249
rect 1271 2245 1272 2249
rect 1266 2244 1272 2245
rect 1268 2171 1270 2244
rect 1376 2200 1378 2334
rect 1560 2295 1562 2335
rect 1794 2334 1800 2335
rect 1816 2295 1818 2335
rect 1914 2334 1920 2335
rect 1934 2339 1940 2340
rect 1934 2335 1935 2339
rect 1939 2335 1940 2339
rect 1974 2339 1975 2343
rect 1979 2339 1980 2343
rect 2022 2340 2023 2344
rect 2027 2340 2028 2344
rect 2022 2339 2028 2340
rect 2114 2343 2120 2344
rect 2114 2339 2115 2343
rect 2119 2339 2120 2343
rect 2302 2340 2303 2344
rect 2307 2340 2308 2344
rect 2302 2339 2308 2340
rect 2578 2343 2584 2344
rect 2578 2339 2579 2343
rect 2583 2339 2584 2343
rect 2598 2340 2599 2344
rect 2603 2340 2604 2344
rect 2598 2339 2604 2340
rect 2690 2343 2696 2344
rect 2690 2339 2691 2343
rect 2695 2339 2696 2343
rect 1974 2338 1980 2339
rect 1934 2334 1940 2335
rect 1936 2295 1938 2334
rect 1976 2303 1978 2338
rect 2024 2303 2026 2339
rect 2114 2338 2120 2339
rect 1975 2302 1979 2303
rect 1975 2297 1979 2298
rect 2023 2302 2027 2303
rect 2023 2297 2027 2298
rect 1559 2294 1563 2295
rect 1559 2289 1563 2290
rect 1815 2294 1819 2295
rect 1815 2289 1819 2290
rect 1935 2294 1939 2295
rect 1935 2289 1939 2290
rect 1936 2266 1938 2289
rect 1976 2274 1978 2297
rect 1974 2273 1980 2274
rect 2024 2273 2026 2297
rect 1974 2269 1975 2273
rect 1979 2269 1980 2273
rect 1974 2268 1980 2269
rect 2022 2272 2028 2273
rect 2022 2268 2023 2272
rect 2027 2268 2028 2272
rect 2022 2267 2028 2268
rect 1934 2265 1940 2266
rect 1386 2263 1392 2264
rect 1386 2259 1387 2263
rect 1391 2259 1392 2263
rect 1934 2261 1935 2265
rect 1939 2261 1940 2265
rect 1934 2260 1940 2261
rect 1386 2258 1392 2259
rect 1374 2199 1380 2200
rect 1374 2195 1375 2199
rect 1379 2195 1380 2199
rect 1374 2194 1380 2195
rect 1388 2192 1390 2258
rect 1994 2257 2000 2258
rect 1974 2256 1980 2257
rect 1974 2252 1975 2256
rect 1979 2252 1980 2256
rect 1994 2253 1995 2257
rect 1999 2253 2000 2257
rect 1994 2252 2000 2253
rect 1974 2251 1980 2252
rect 1934 2248 1940 2249
rect 1934 2244 1935 2248
rect 1939 2244 1940 2248
rect 1934 2243 1940 2244
rect 1386 2191 1392 2192
rect 1386 2187 1387 2191
rect 1391 2187 1392 2191
rect 1386 2186 1392 2187
rect 1936 2171 1938 2243
rect 1976 2183 1978 2251
rect 1996 2183 1998 2252
rect 2116 2208 2118 2338
rect 2304 2303 2306 2339
rect 2578 2338 2584 2339
rect 2600 2303 2602 2339
rect 2690 2338 2696 2339
rect 2159 2302 2163 2303
rect 2159 2297 2163 2298
rect 2295 2302 2299 2303
rect 2295 2297 2299 2298
rect 2303 2302 2307 2303
rect 2303 2297 2307 2298
rect 2447 2302 2451 2303
rect 2447 2297 2451 2298
rect 2599 2302 2603 2303
rect 2599 2297 2603 2298
rect 2607 2302 2611 2303
rect 2607 2297 2611 2298
rect 2160 2273 2162 2297
rect 2296 2273 2298 2297
rect 2448 2273 2450 2297
rect 2608 2273 2610 2297
rect 2158 2272 2164 2273
rect 2294 2272 2300 2273
rect 2122 2271 2128 2272
rect 2122 2267 2123 2271
rect 2127 2267 2128 2271
rect 2158 2268 2159 2272
rect 2163 2268 2164 2272
rect 2158 2267 2164 2268
rect 2258 2271 2264 2272
rect 2258 2267 2259 2271
rect 2263 2267 2264 2271
rect 2294 2268 2295 2272
rect 2299 2268 2300 2272
rect 2294 2267 2300 2268
rect 2446 2272 2452 2273
rect 2606 2272 2612 2273
rect 2704 2272 2706 2410
rect 2860 2360 2862 2421
rect 3004 2412 3006 2518
rect 3034 2509 3040 2510
rect 3034 2505 3035 2509
rect 3039 2505 3040 2509
rect 3034 2504 3040 2505
rect 3036 2427 3038 2504
rect 3096 2460 3098 2578
rect 3800 2555 3802 2578
rect 3840 2557 3842 2617
rect 3838 2556 3844 2557
rect 3892 2556 3894 2617
rect 3986 2603 3992 2604
rect 3986 2599 3987 2603
rect 3991 2599 3992 2603
rect 3986 2598 3992 2599
rect 3223 2554 3227 2555
rect 3223 2549 3227 2550
rect 3799 2554 3803 2555
rect 3838 2552 3839 2556
rect 3843 2552 3844 2556
rect 3838 2551 3844 2552
rect 3890 2555 3896 2556
rect 3890 2551 3891 2555
rect 3895 2551 3896 2555
rect 3890 2550 3896 2551
rect 3799 2549 3803 2550
rect 3224 2525 3226 2549
rect 3800 2526 3802 2549
rect 3918 2540 3924 2541
rect 3838 2539 3844 2540
rect 3838 2535 3839 2539
rect 3843 2535 3844 2539
rect 3918 2536 3919 2540
rect 3923 2536 3924 2540
rect 3918 2535 3924 2536
rect 3838 2534 3844 2535
rect 3798 2525 3804 2526
rect 3222 2524 3228 2525
rect 3162 2523 3168 2524
rect 3162 2519 3163 2523
rect 3167 2519 3168 2523
rect 3222 2520 3223 2524
rect 3227 2520 3228 2524
rect 3222 2519 3228 2520
rect 3318 2523 3324 2524
rect 3318 2519 3319 2523
rect 3323 2519 3324 2523
rect 3798 2521 3799 2525
rect 3803 2521 3804 2525
rect 3798 2520 3804 2521
rect 3162 2518 3168 2519
rect 3318 2518 3324 2519
rect 3164 2460 3166 2518
rect 3194 2509 3200 2510
rect 3194 2505 3195 2509
rect 3199 2505 3200 2509
rect 3194 2504 3200 2505
rect 3094 2459 3100 2460
rect 3094 2455 3095 2459
rect 3099 2455 3100 2459
rect 3094 2454 3100 2455
rect 3162 2459 3168 2460
rect 3162 2455 3163 2459
rect 3167 2455 3168 2459
rect 3162 2454 3168 2455
rect 3196 2427 3198 2504
rect 3320 2452 3322 2518
rect 3798 2508 3804 2509
rect 3798 2504 3799 2508
rect 3803 2504 3804 2508
rect 3840 2507 3842 2534
rect 3920 2507 3922 2535
rect 3798 2503 3804 2504
rect 3839 2506 3843 2507
rect 3318 2451 3324 2452
rect 3318 2447 3319 2451
rect 3323 2447 3324 2451
rect 3318 2446 3324 2447
rect 3800 2427 3802 2503
rect 3839 2501 3843 2502
rect 3887 2506 3891 2507
rect 3887 2501 3891 2502
rect 3919 2506 3923 2507
rect 3919 2501 3923 2502
rect 3840 2478 3842 2501
rect 3838 2477 3844 2478
rect 3888 2477 3890 2501
rect 3838 2473 3839 2477
rect 3843 2473 3844 2477
rect 3838 2472 3844 2473
rect 3886 2476 3892 2477
rect 3988 2476 3990 2598
rect 4068 2556 4070 2617
rect 4074 2603 4080 2604
rect 4074 2599 4075 2603
rect 4079 2599 4080 2603
rect 4074 2598 4080 2599
rect 4066 2555 4072 2556
rect 4066 2551 4067 2555
rect 4071 2551 4072 2555
rect 4066 2550 4072 2551
rect 4076 2540 4078 2598
rect 4094 2540 4100 2541
rect 4188 2540 4190 2626
rect 4196 2623 4198 2684
rect 4195 2622 4199 2623
rect 4195 2617 4199 2618
rect 4267 2622 4271 2623
rect 4267 2617 4271 2618
rect 4268 2556 4270 2617
rect 4364 2608 4366 2714
rect 4528 2705 4530 2729
rect 4864 2705 4866 2729
rect 5216 2705 5218 2729
rect 4526 2704 4532 2705
rect 4862 2704 4868 2705
rect 5214 2704 5220 2705
rect 4422 2703 4428 2704
rect 4422 2699 4423 2703
rect 4427 2699 4428 2703
rect 4526 2700 4527 2704
rect 4531 2700 4532 2704
rect 4526 2699 4532 2700
rect 4626 2703 4632 2704
rect 4626 2699 4627 2703
rect 4631 2699 4632 2703
rect 4862 2700 4863 2704
rect 4867 2700 4868 2704
rect 4862 2699 4868 2700
rect 4982 2703 4988 2704
rect 4982 2699 4983 2703
rect 4987 2699 4988 2703
rect 5214 2700 5215 2704
rect 5219 2700 5220 2704
rect 5214 2699 5220 2700
rect 4422 2698 4428 2699
rect 4626 2698 4632 2699
rect 4982 2698 4988 2699
rect 4424 2640 4426 2698
rect 4498 2689 4504 2690
rect 4498 2685 4499 2689
rect 4503 2685 4504 2689
rect 4498 2684 4504 2685
rect 4422 2639 4428 2640
rect 4422 2635 4423 2639
rect 4427 2635 4428 2639
rect 4422 2634 4428 2635
rect 4500 2623 4502 2684
rect 4628 2640 4630 2698
rect 4834 2689 4840 2690
rect 4834 2685 4835 2689
rect 4839 2685 4840 2689
rect 4834 2684 4840 2685
rect 4626 2639 4632 2640
rect 4626 2635 4627 2639
rect 4631 2635 4632 2639
rect 4626 2634 4632 2635
rect 4836 2623 4838 2684
rect 4984 2640 4986 2698
rect 5186 2689 5192 2690
rect 5186 2685 5187 2689
rect 5191 2685 5192 2689
rect 5186 2684 5192 2685
rect 4982 2639 4988 2640
rect 4982 2635 4983 2639
rect 4987 2635 4988 2639
rect 4982 2634 4988 2635
rect 5188 2623 5190 2684
rect 4491 2622 4495 2623
rect 4491 2617 4495 2618
rect 4499 2622 4503 2623
rect 4499 2617 4503 2618
rect 4731 2622 4735 2623
rect 4731 2617 4735 2618
rect 4835 2622 4839 2623
rect 4835 2617 4839 2618
rect 4995 2622 4999 2623
rect 4995 2617 4999 2618
rect 5187 2622 5191 2623
rect 5187 2617 5191 2618
rect 5267 2622 5271 2623
rect 5267 2617 5271 2618
rect 4362 2607 4368 2608
rect 4362 2603 4363 2607
rect 4367 2603 4368 2607
rect 4362 2602 4368 2603
rect 4492 2556 4494 2617
rect 4498 2603 4504 2604
rect 4498 2599 4499 2603
rect 4503 2599 4504 2603
rect 4498 2598 4504 2599
rect 4266 2555 4272 2556
rect 4266 2551 4267 2555
rect 4271 2551 4272 2555
rect 4266 2550 4272 2551
rect 4490 2555 4496 2556
rect 4490 2551 4491 2555
rect 4495 2551 4496 2555
rect 4490 2550 4496 2551
rect 4294 2540 4300 2541
rect 4500 2540 4502 2598
rect 4732 2556 4734 2617
rect 4738 2603 4744 2604
rect 4738 2599 4739 2603
rect 4743 2599 4744 2603
rect 4738 2598 4744 2599
rect 4730 2555 4736 2556
rect 4730 2551 4731 2555
rect 4735 2551 4736 2555
rect 4730 2550 4736 2551
rect 4518 2540 4524 2541
rect 4740 2540 4742 2598
rect 4996 2556 4998 2617
rect 5002 2603 5008 2604
rect 5002 2599 5003 2603
rect 5007 2599 5008 2603
rect 5002 2598 5008 2599
rect 4994 2555 5000 2556
rect 4994 2551 4995 2555
rect 4999 2551 5000 2555
rect 4994 2550 5000 2551
rect 4758 2540 4764 2541
rect 5004 2540 5006 2598
rect 5268 2556 5270 2617
rect 5266 2555 5272 2556
rect 5266 2551 5267 2555
rect 5271 2551 5272 2555
rect 5266 2550 5272 2551
rect 5022 2540 5028 2541
rect 5294 2540 5300 2541
rect 5392 2540 5394 2838
rect 5516 2792 5518 2853
rect 5636 2844 5638 2950
rect 5662 2940 5668 2941
rect 5662 2936 5663 2940
rect 5667 2936 5668 2940
rect 5662 2935 5668 2936
rect 5664 2859 5666 2935
rect 5663 2858 5667 2859
rect 5663 2853 5667 2854
rect 5634 2843 5640 2844
rect 5634 2839 5635 2843
rect 5639 2839 5640 2843
rect 5634 2838 5640 2839
rect 5664 2793 5666 2853
rect 5662 2792 5668 2793
rect 5514 2791 5520 2792
rect 5514 2787 5515 2791
rect 5519 2787 5520 2791
rect 5662 2788 5663 2792
rect 5667 2788 5668 2792
rect 5662 2787 5668 2788
rect 5514 2786 5520 2787
rect 5542 2776 5548 2777
rect 5542 2772 5543 2776
rect 5547 2772 5548 2776
rect 5542 2771 5548 2772
rect 5642 2775 5648 2776
rect 5642 2771 5643 2775
rect 5647 2771 5648 2775
rect 5544 2735 5546 2771
rect 5642 2770 5648 2771
rect 5662 2775 5668 2776
rect 5662 2771 5663 2775
rect 5667 2771 5668 2775
rect 5662 2770 5668 2771
rect 5543 2734 5547 2735
rect 5543 2729 5547 2730
rect 5544 2705 5546 2729
rect 5542 2704 5548 2705
rect 5542 2700 5543 2704
rect 5547 2700 5548 2704
rect 5542 2699 5548 2700
rect 5634 2703 5640 2704
rect 5634 2699 5635 2703
rect 5639 2699 5640 2703
rect 5634 2698 5640 2699
rect 5514 2689 5520 2690
rect 5514 2685 5515 2689
rect 5519 2685 5520 2689
rect 5514 2684 5520 2685
rect 5516 2623 5518 2684
rect 5515 2622 5519 2623
rect 5515 2617 5519 2618
rect 5442 2607 5448 2608
rect 5442 2603 5443 2607
rect 5447 2603 5448 2607
rect 5442 2602 5448 2603
rect 4074 2539 4080 2540
rect 4074 2535 4075 2539
rect 4079 2535 4080 2539
rect 4094 2536 4095 2540
rect 4099 2536 4100 2540
rect 4094 2535 4100 2536
rect 4186 2539 4192 2540
rect 4186 2535 4187 2539
rect 4191 2535 4192 2539
rect 4294 2536 4295 2540
rect 4299 2536 4300 2540
rect 4294 2535 4300 2536
rect 4498 2539 4504 2540
rect 4498 2535 4499 2539
rect 4503 2535 4504 2539
rect 4518 2536 4519 2540
rect 4523 2536 4524 2540
rect 4518 2535 4524 2536
rect 4738 2539 4744 2540
rect 4738 2535 4739 2539
rect 4743 2535 4744 2539
rect 4758 2536 4759 2540
rect 4763 2536 4764 2540
rect 4758 2535 4764 2536
rect 5002 2539 5008 2540
rect 5002 2535 5003 2539
rect 5007 2535 5008 2539
rect 5022 2536 5023 2540
rect 5027 2536 5028 2540
rect 5022 2535 5028 2536
rect 5114 2539 5120 2540
rect 5114 2535 5115 2539
rect 5119 2535 5120 2539
rect 5294 2536 5295 2540
rect 5299 2536 5300 2540
rect 5294 2535 5300 2536
rect 5390 2539 5396 2540
rect 5390 2535 5391 2539
rect 5395 2535 5396 2539
rect 4074 2534 4080 2535
rect 4096 2507 4098 2535
rect 4186 2534 4192 2535
rect 4296 2507 4298 2535
rect 4498 2534 4504 2535
rect 4520 2507 4522 2535
rect 4738 2534 4744 2535
rect 4760 2507 4762 2535
rect 5002 2534 5008 2535
rect 5024 2507 5026 2535
rect 5114 2534 5120 2535
rect 4087 2506 4091 2507
rect 4087 2501 4091 2502
rect 4095 2506 4099 2507
rect 4095 2501 4099 2502
rect 4295 2506 4299 2507
rect 4295 2501 4299 2502
rect 4319 2506 4323 2507
rect 4319 2501 4323 2502
rect 4519 2506 4523 2507
rect 4519 2501 4523 2502
rect 4567 2506 4571 2507
rect 4567 2501 4571 2502
rect 4759 2506 4763 2507
rect 4759 2501 4763 2502
rect 4823 2506 4827 2507
rect 4823 2501 4827 2502
rect 5023 2506 5027 2507
rect 5023 2501 5027 2502
rect 5087 2506 5091 2507
rect 5087 2501 5091 2502
rect 4088 2477 4090 2501
rect 4320 2477 4322 2501
rect 4568 2477 4570 2501
rect 4824 2477 4826 2501
rect 5088 2477 5090 2501
rect 4086 2476 4092 2477
rect 4318 2476 4324 2477
rect 4566 2476 4572 2477
rect 4822 2476 4828 2477
rect 5086 2476 5092 2477
rect 3886 2472 3887 2476
rect 3891 2472 3892 2476
rect 3886 2471 3892 2472
rect 3986 2475 3992 2476
rect 3986 2471 3987 2475
rect 3991 2471 3992 2475
rect 4086 2472 4087 2476
rect 4091 2472 4092 2476
rect 4086 2471 4092 2472
rect 4182 2475 4188 2476
rect 4182 2471 4183 2475
rect 4187 2471 4188 2475
rect 4318 2472 4319 2476
rect 4323 2472 4324 2476
rect 4318 2471 4324 2472
rect 4438 2475 4444 2476
rect 4438 2471 4439 2475
rect 4443 2471 4444 2475
rect 4566 2472 4567 2476
rect 4571 2472 4572 2476
rect 4566 2471 4572 2472
rect 4710 2475 4716 2476
rect 4710 2471 4711 2475
rect 4715 2471 4716 2475
rect 4822 2472 4823 2476
rect 4827 2472 4828 2476
rect 4822 2471 4828 2472
rect 4974 2475 4980 2476
rect 4974 2471 4975 2475
rect 4979 2471 4980 2475
rect 5086 2472 5087 2476
rect 5091 2472 5092 2476
rect 5086 2471 5092 2472
rect 3986 2470 3992 2471
rect 4182 2470 4188 2471
rect 4438 2470 4444 2471
rect 4710 2470 4716 2471
rect 4974 2470 4980 2471
rect 3858 2461 3864 2462
rect 3838 2460 3844 2461
rect 3838 2456 3839 2460
rect 3843 2456 3844 2460
rect 3858 2457 3859 2461
rect 3863 2457 3864 2461
rect 3858 2456 3864 2457
rect 4058 2461 4064 2462
rect 4058 2457 4059 2461
rect 4063 2457 4064 2461
rect 4058 2456 4064 2457
rect 3838 2455 3844 2456
rect 3035 2426 3039 2427
rect 3035 2421 3039 2422
rect 3147 2426 3151 2427
rect 3147 2421 3151 2422
rect 3195 2426 3199 2427
rect 3195 2421 3199 2422
rect 3435 2426 3439 2427
rect 3435 2421 3439 2422
rect 3799 2426 3803 2427
rect 3799 2421 3803 2422
rect 3002 2411 3008 2412
rect 3002 2407 3003 2411
rect 3007 2407 3008 2411
rect 3002 2406 3008 2407
rect 3148 2360 3150 2421
rect 3154 2407 3160 2408
rect 3154 2403 3155 2407
rect 3159 2403 3160 2407
rect 3154 2402 3160 2403
rect 2858 2359 2864 2360
rect 2858 2355 2859 2359
rect 2863 2355 2864 2359
rect 2858 2354 2864 2355
rect 3146 2359 3152 2360
rect 3146 2355 3147 2359
rect 3151 2355 3152 2359
rect 3146 2354 3152 2355
rect 2886 2344 2892 2345
rect 3156 2344 3158 2402
rect 3436 2360 3438 2421
rect 3442 2407 3448 2408
rect 3442 2403 3443 2407
rect 3447 2403 3448 2407
rect 3442 2402 3448 2403
rect 3434 2359 3440 2360
rect 3434 2355 3435 2359
rect 3439 2355 3440 2359
rect 3434 2354 3440 2355
rect 3174 2344 3180 2345
rect 3444 2344 3446 2402
rect 3790 2379 3796 2380
rect 3790 2375 3791 2379
rect 3795 2375 3796 2379
rect 3790 2374 3796 2375
rect 3462 2344 3468 2345
rect 2886 2340 2887 2344
rect 2891 2340 2892 2344
rect 2886 2339 2892 2340
rect 3154 2343 3160 2344
rect 3154 2339 3155 2343
rect 3159 2339 3160 2343
rect 3174 2340 3175 2344
rect 3179 2340 3180 2344
rect 3174 2339 3180 2340
rect 3442 2343 3448 2344
rect 3442 2339 3443 2343
rect 3447 2339 3448 2343
rect 3462 2340 3463 2344
rect 3467 2340 3468 2344
rect 3462 2339 3468 2340
rect 3558 2343 3564 2344
rect 3558 2339 3559 2343
rect 3563 2339 3564 2343
rect 2888 2303 2890 2339
rect 3154 2338 3160 2339
rect 3176 2303 3178 2339
rect 3442 2338 3448 2339
rect 3464 2303 3466 2339
rect 3558 2338 3564 2339
rect 2767 2302 2771 2303
rect 2767 2297 2771 2298
rect 2887 2302 2891 2303
rect 2887 2297 2891 2298
rect 2927 2302 2931 2303
rect 2927 2297 2931 2298
rect 3079 2302 3083 2303
rect 3079 2297 3083 2298
rect 3175 2302 3179 2303
rect 3175 2297 3179 2298
rect 3231 2302 3235 2303
rect 3231 2297 3235 2298
rect 3383 2302 3387 2303
rect 3383 2297 3387 2298
rect 3463 2302 3467 2303
rect 3463 2297 3467 2298
rect 3543 2302 3547 2303
rect 3543 2297 3547 2298
rect 2768 2273 2770 2297
rect 2928 2273 2930 2297
rect 3080 2273 3082 2297
rect 3232 2273 3234 2297
rect 3384 2273 3386 2297
rect 3544 2273 3546 2297
rect 2766 2272 2772 2273
rect 2926 2272 2932 2273
rect 3078 2272 3084 2273
rect 3230 2272 3236 2273
rect 3382 2272 3388 2273
rect 3542 2272 3548 2273
rect 2446 2268 2447 2272
rect 2451 2268 2452 2272
rect 2446 2267 2452 2268
rect 2538 2271 2544 2272
rect 2538 2267 2539 2271
rect 2543 2267 2544 2271
rect 2606 2268 2607 2272
rect 2611 2268 2612 2272
rect 2606 2267 2612 2268
rect 2702 2271 2708 2272
rect 2702 2267 2703 2271
rect 2707 2267 2708 2271
rect 2766 2268 2767 2272
rect 2771 2268 2772 2272
rect 2766 2267 2772 2268
rect 2858 2271 2864 2272
rect 2858 2267 2859 2271
rect 2863 2267 2864 2271
rect 2926 2268 2927 2272
rect 2931 2268 2932 2272
rect 2926 2267 2932 2268
rect 3018 2271 3024 2272
rect 3018 2267 3019 2271
rect 3023 2267 3024 2271
rect 3078 2268 3079 2272
rect 3083 2268 3084 2272
rect 3078 2267 3084 2268
rect 3174 2271 3180 2272
rect 3174 2267 3175 2271
rect 3179 2267 3180 2271
rect 3230 2268 3231 2272
rect 3235 2268 3236 2272
rect 3230 2267 3236 2268
rect 3326 2271 3332 2272
rect 3326 2267 3327 2271
rect 3331 2267 3332 2271
rect 3382 2268 3383 2272
rect 3387 2268 3388 2272
rect 3382 2267 3388 2268
rect 3478 2271 3484 2272
rect 3478 2267 3479 2271
rect 3483 2267 3484 2271
rect 3542 2268 3543 2272
rect 3547 2268 3548 2272
rect 3542 2267 3548 2268
rect 2122 2266 2128 2267
rect 2258 2266 2264 2267
rect 2538 2266 2544 2267
rect 2702 2266 2708 2267
rect 2858 2266 2864 2267
rect 3018 2266 3024 2267
rect 3174 2266 3180 2267
rect 3326 2266 3332 2267
rect 3478 2266 3484 2267
rect 2124 2208 2126 2266
rect 2130 2257 2136 2258
rect 2130 2253 2131 2257
rect 2135 2253 2136 2257
rect 2130 2252 2136 2253
rect 2114 2207 2120 2208
rect 2114 2203 2115 2207
rect 2119 2203 2120 2207
rect 2114 2202 2120 2203
rect 2122 2207 2128 2208
rect 2122 2203 2123 2207
rect 2127 2203 2128 2207
rect 2122 2202 2128 2203
rect 2132 2183 2134 2252
rect 2260 2208 2262 2266
rect 2266 2257 2272 2258
rect 2266 2253 2267 2257
rect 2271 2253 2272 2257
rect 2266 2252 2272 2253
rect 2418 2257 2424 2258
rect 2418 2253 2419 2257
rect 2423 2253 2424 2257
rect 2418 2252 2424 2253
rect 2258 2207 2264 2208
rect 2258 2203 2259 2207
rect 2263 2203 2264 2207
rect 2258 2202 2264 2203
rect 2268 2183 2270 2252
rect 2420 2183 2422 2252
rect 1975 2182 1979 2183
rect 1975 2177 1979 2178
rect 1995 2182 1999 2183
rect 1995 2177 1999 2178
rect 2131 2182 2135 2183
rect 2131 2177 2135 2178
rect 2267 2182 2271 2183
rect 2267 2177 2271 2178
rect 2331 2182 2335 2183
rect 2331 2177 2335 2178
rect 2419 2182 2423 2183
rect 2419 2177 2423 2178
rect 2531 2182 2535 2183
rect 2531 2177 2535 2178
rect 1267 2170 1271 2171
rect 1267 2165 1271 2166
rect 1443 2170 1447 2171
rect 1443 2165 1447 2166
rect 1787 2170 1791 2171
rect 1787 2165 1791 2166
rect 1935 2170 1939 2171
rect 1935 2165 1939 2166
rect 1094 2155 1100 2156
rect 1094 2151 1095 2155
rect 1099 2151 1100 2155
rect 1094 2150 1100 2151
rect 1444 2104 1446 2165
rect 1450 2151 1456 2152
rect 1450 2147 1451 2151
rect 1455 2147 1456 2151
rect 1450 2146 1456 2147
rect 1082 2103 1088 2104
rect 1082 2099 1083 2103
rect 1087 2099 1088 2103
rect 1082 2098 1088 2099
rect 1442 2103 1448 2104
rect 1442 2099 1443 2103
rect 1447 2099 1448 2103
rect 1442 2098 1448 2099
rect 1110 2088 1116 2089
rect 1452 2088 1454 2146
rect 1788 2104 1790 2165
rect 1936 2105 1938 2165
rect 1976 2117 1978 2177
rect 2118 2155 2124 2156
rect 2118 2151 2119 2155
rect 2123 2151 2124 2155
rect 2118 2150 2124 2151
rect 1974 2116 1980 2117
rect 1974 2112 1975 2116
rect 1979 2112 1980 2116
rect 1974 2111 1980 2112
rect 1934 2104 1940 2105
rect 1786 2103 1792 2104
rect 1786 2099 1787 2103
rect 1791 2099 1792 2103
rect 1934 2100 1935 2104
rect 1939 2100 1940 2104
rect 1934 2099 1940 2100
rect 1974 2099 1980 2100
rect 1786 2098 1792 2099
rect 1974 2095 1975 2099
rect 1979 2095 1980 2099
rect 1974 2094 1980 2095
rect 1470 2088 1476 2089
rect 1814 2088 1820 2089
rect 758 2084 759 2088
rect 763 2084 764 2088
rect 758 2083 764 2084
rect 854 2087 860 2088
rect 854 2083 855 2087
rect 859 2083 860 2087
rect 1110 2084 1111 2088
rect 1115 2084 1116 2088
rect 1110 2083 1116 2084
rect 1450 2087 1456 2088
rect 1450 2083 1451 2087
rect 1455 2083 1456 2087
rect 1470 2084 1471 2088
rect 1475 2084 1476 2088
rect 1470 2083 1476 2084
rect 1566 2087 1572 2088
rect 1566 2083 1567 2087
rect 1571 2083 1572 2087
rect 1814 2084 1815 2088
rect 1819 2084 1820 2088
rect 1814 2083 1820 2084
rect 1910 2087 1916 2088
rect 1910 2083 1911 2087
rect 1915 2083 1916 2087
rect 760 2055 762 2083
rect 854 2082 860 2083
rect 1112 2055 1114 2083
rect 1450 2082 1456 2083
rect 1472 2055 1474 2083
rect 1566 2082 1572 2083
rect 751 2054 755 2055
rect 751 2049 755 2050
rect 759 2054 763 2055
rect 759 2049 763 2050
rect 959 2054 963 2055
rect 959 2049 963 2050
rect 1111 2054 1115 2055
rect 1111 2049 1115 2050
rect 1167 2054 1171 2055
rect 1167 2049 1171 2050
rect 1383 2054 1387 2055
rect 1383 2049 1387 2050
rect 1471 2054 1475 2055
rect 1471 2049 1475 2050
rect 752 2025 754 2049
rect 960 2025 962 2049
rect 1168 2025 1170 2049
rect 1384 2025 1386 2049
rect 750 2024 756 2025
rect 958 2024 964 2025
rect 1166 2024 1172 2025
rect 1382 2024 1388 2025
rect 558 2020 559 2024
rect 563 2020 564 2024
rect 558 2019 564 2020
rect 738 2023 744 2024
rect 738 2019 739 2023
rect 743 2019 744 2023
rect 750 2020 751 2024
rect 755 2020 756 2024
rect 750 2019 756 2020
rect 842 2023 848 2024
rect 842 2019 843 2023
rect 847 2019 848 2023
rect 958 2020 959 2024
rect 963 2020 964 2024
rect 958 2019 964 2020
rect 1054 2023 1060 2024
rect 1054 2019 1055 2023
rect 1059 2019 1060 2023
rect 1166 2020 1167 2024
rect 1171 2020 1172 2024
rect 1166 2019 1172 2020
rect 1258 2023 1264 2024
rect 1258 2019 1259 2023
rect 1263 2019 1264 2023
rect 1382 2020 1383 2024
rect 1387 2020 1388 2024
rect 1382 2019 1388 2020
rect 1482 2023 1488 2024
rect 1482 2019 1483 2023
rect 1487 2019 1488 2023
rect 322 2018 328 2019
rect 738 2018 744 2019
rect 842 2018 848 2019
rect 1054 2018 1060 2019
rect 1258 2018 1264 2019
rect 1482 2018 1488 2019
rect 194 2009 200 2010
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 194 2005 195 2009
rect 199 2005 200 2009
rect 194 2004 200 2005
rect 110 2003 116 2004
rect 112 1935 114 2003
rect 196 1935 198 2004
rect 324 1960 326 2018
rect 354 2009 360 2010
rect 354 2005 355 2009
rect 359 2005 360 2009
rect 354 2004 360 2005
rect 530 2009 536 2010
rect 530 2005 531 2009
rect 535 2005 536 2009
rect 530 2004 536 2005
rect 722 2009 728 2010
rect 722 2005 723 2009
rect 727 2005 728 2009
rect 722 2004 728 2005
rect 314 1959 320 1960
rect 314 1955 315 1959
rect 319 1955 320 1959
rect 314 1954 320 1955
rect 322 1959 328 1960
rect 322 1955 323 1959
rect 327 1955 328 1959
rect 322 1954 328 1955
rect 111 1934 115 1935
rect 111 1929 115 1930
rect 195 1934 199 1935
rect 195 1929 199 1930
rect 112 1869 114 1929
rect 110 1868 116 1869
rect 196 1868 198 1929
rect 110 1864 111 1868
rect 115 1864 116 1868
rect 110 1863 116 1864
rect 194 1867 200 1868
rect 194 1863 195 1867
rect 199 1863 200 1867
rect 194 1862 200 1863
rect 222 1852 228 1853
rect 316 1852 318 1954
rect 356 1935 358 2004
rect 532 1935 534 2004
rect 724 1935 726 2004
rect 355 1934 359 1935
rect 355 1929 359 1930
rect 387 1934 391 1935
rect 387 1929 391 1930
rect 531 1934 535 1935
rect 531 1929 535 1930
rect 595 1934 599 1935
rect 595 1929 599 1930
rect 723 1934 727 1935
rect 723 1929 727 1930
rect 819 1934 823 1935
rect 819 1929 823 1930
rect 388 1868 390 1929
rect 506 1923 512 1924
rect 506 1919 507 1923
rect 511 1919 512 1923
rect 506 1918 512 1919
rect 386 1867 392 1868
rect 386 1863 387 1867
rect 391 1863 392 1867
rect 386 1862 392 1863
rect 414 1852 420 1853
rect 508 1852 510 1918
rect 574 1911 580 1912
rect 574 1907 575 1911
rect 579 1907 580 1911
rect 574 1906 580 1907
rect 110 1851 116 1852
rect 110 1847 111 1851
rect 115 1847 116 1851
rect 222 1848 223 1852
rect 227 1848 228 1852
rect 222 1847 228 1848
rect 314 1851 320 1852
rect 314 1847 315 1851
rect 319 1847 320 1851
rect 414 1848 415 1852
rect 419 1848 420 1852
rect 414 1847 420 1848
rect 506 1851 512 1852
rect 506 1847 507 1851
rect 511 1847 512 1851
rect 110 1846 116 1847
rect 112 1807 114 1846
rect 224 1807 226 1847
rect 314 1846 320 1847
rect 416 1807 418 1847
rect 506 1846 512 1847
rect 111 1806 115 1807
rect 111 1801 115 1802
rect 159 1806 163 1807
rect 159 1801 163 1802
rect 223 1806 227 1807
rect 223 1801 227 1802
rect 303 1806 307 1807
rect 303 1801 307 1802
rect 415 1806 419 1807
rect 415 1801 419 1802
rect 479 1806 483 1807
rect 479 1801 483 1802
rect 112 1778 114 1801
rect 110 1777 116 1778
rect 160 1777 162 1801
rect 304 1777 306 1801
rect 480 1777 482 1801
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 110 1772 116 1773
rect 158 1776 164 1777
rect 302 1776 308 1777
rect 478 1776 484 1777
rect 576 1776 578 1906
rect 596 1868 598 1929
rect 820 1868 822 1929
rect 844 1928 846 2018
rect 930 2009 936 2010
rect 930 2005 931 2009
rect 935 2005 936 2009
rect 930 2004 936 2005
rect 932 1935 934 2004
rect 1026 1987 1032 1988
rect 1026 1983 1027 1987
rect 1031 1983 1032 1987
rect 1026 1982 1032 1983
rect 1028 1960 1030 1982
rect 1026 1959 1032 1960
rect 1026 1955 1027 1959
rect 1031 1955 1032 1959
rect 1026 1954 1032 1955
rect 1056 1952 1058 2018
rect 1138 2009 1144 2010
rect 1138 2005 1139 2009
rect 1143 2005 1144 2009
rect 1138 2004 1144 2005
rect 1054 1951 1060 1952
rect 1054 1947 1055 1951
rect 1059 1947 1060 1951
rect 1054 1946 1060 1947
rect 1140 1935 1142 2004
rect 1234 2003 1240 2004
rect 1234 1999 1235 2003
rect 1239 1999 1240 2003
rect 1234 1998 1240 1999
rect 1236 1960 1238 1998
rect 1260 1988 1262 2018
rect 1354 2009 1360 2010
rect 1354 2005 1355 2009
rect 1359 2005 1360 2009
rect 1354 2004 1360 2005
rect 1258 1987 1264 1988
rect 1258 1983 1259 1987
rect 1263 1983 1264 1987
rect 1258 1982 1264 1983
rect 1234 1959 1240 1960
rect 1234 1955 1235 1959
rect 1239 1955 1240 1959
rect 1234 1954 1240 1955
rect 1356 1935 1358 2004
rect 931 1934 935 1935
rect 931 1929 935 1930
rect 1051 1934 1055 1935
rect 1051 1929 1055 1930
rect 1139 1934 1143 1935
rect 1139 1929 1143 1930
rect 1283 1934 1287 1935
rect 1283 1929 1287 1930
rect 1355 1934 1359 1935
rect 1355 1929 1359 1930
rect 842 1927 848 1928
rect 842 1923 843 1927
rect 847 1923 848 1927
rect 842 1922 848 1923
rect 826 1915 832 1916
rect 826 1911 827 1915
rect 831 1911 832 1915
rect 826 1910 832 1911
rect 594 1867 600 1868
rect 594 1863 595 1867
rect 599 1863 600 1867
rect 594 1862 600 1863
rect 818 1867 824 1868
rect 818 1863 819 1867
rect 823 1863 824 1867
rect 818 1862 824 1863
rect 622 1852 628 1853
rect 828 1852 830 1910
rect 1052 1868 1054 1929
rect 1058 1915 1064 1916
rect 1058 1911 1059 1915
rect 1063 1911 1064 1915
rect 1058 1910 1064 1911
rect 1050 1867 1056 1868
rect 1050 1863 1051 1867
rect 1055 1863 1056 1867
rect 1050 1862 1056 1863
rect 846 1852 852 1853
rect 1060 1852 1062 1910
rect 1284 1868 1286 1929
rect 1484 1920 1486 2018
rect 1568 2004 1570 2082
rect 1816 2055 1818 2083
rect 1910 2082 1916 2083
rect 1934 2087 1940 2088
rect 1934 2083 1935 2087
rect 1939 2083 1940 2087
rect 1934 2082 1940 2083
rect 1607 2054 1611 2055
rect 1607 2049 1611 2050
rect 1815 2054 1819 2055
rect 1815 2049 1819 2050
rect 1608 2025 1610 2049
rect 1816 2025 1818 2049
rect 1606 2024 1612 2025
rect 1814 2024 1820 2025
rect 1606 2020 1607 2024
rect 1611 2020 1612 2024
rect 1606 2019 1612 2020
rect 1702 2023 1708 2024
rect 1702 2019 1703 2023
rect 1707 2019 1708 2023
rect 1814 2020 1815 2024
rect 1819 2020 1820 2024
rect 1814 2019 1820 2020
rect 1702 2018 1708 2019
rect 1578 2009 1584 2010
rect 1578 2005 1579 2009
rect 1583 2005 1584 2009
rect 1578 2004 1584 2005
rect 1566 2003 1572 2004
rect 1566 1999 1567 2003
rect 1571 1999 1572 2003
rect 1566 1998 1572 1999
rect 1580 1935 1582 2004
rect 1674 2003 1680 2004
rect 1674 1999 1675 2003
rect 1679 1999 1680 2003
rect 1674 1998 1680 1999
rect 1676 1960 1678 1998
rect 1674 1959 1680 1960
rect 1674 1955 1675 1959
rect 1679 1955 1680 1959
rect 1674 1954 1680 1955
rect 1704 1952 1706 2018
rect 1786 2009 1792 2010
rect 1786 2005 1787 2009
rect 1791 2005 1792 2009
rect 1786 2004 1792 2005
rect 1702 1951 1708 1952
rect 1702 1947 1703 1951
rect 1707 1947 1708 1951
rect 1702 1946 1708 1947
rect 1788 1935 1790 2004
rect 1912 1960 1914 2082
rect 1936 2055 1938 2082
rect 1976 2063 1978 2094
rect 1975 2062 1979 2063
rect 1975 2057 1979 2058
rect 2023 2062 2027 2063
rect 2023 2057 2027 2058
rect 1935 2054 1939 2055
rect 1935 2049 1939 2050
rect 1936 2026 1938 2049
rect 1976 2034 1978 2057
rect 1974 2033 1980 2034
rect 2024 2033 2026 2057
rect 1974 2029 1975 2033
rect 1979 2029 1980 2033
rect 1974 2028 1980 2029
rect 2022 2032 2028 2033
rect 2120 2032 2122 2150
rect 2132 2116 2134 2177
rect 2332 2116 2334 2177
rect 2338 2163 2344 2164
rect 2338 2159 2339 2163
rect 2343 2159 2344 2163
rect 2338 2158 2344 2159
rect 2130 2115 2136 2116
rect 2130 2111 2131 2115
rect 2135 2111 2136 2115
rect 2130 2110 2136 2111
rect 2330 2115 2336 2116
rect 2330 2111 2331 2115
rect 2335 2111 2336 2115
rect 2330 2110 2336 2111
rect 2158 2100 2164 2101
rect 2340 2100 2342 2158
rect 2532 2116 2534 2177
rect 2540 2176 2542 2266
rect 2578 2257 2584 2258
rect 2578 2253 2579 2257
rect 2583 2253 2584 2257
rect 2578 2252 2584 2253
rect 2738 2257 2744 2258
rect 2738 2253 2739 2257
rect 2743 2253 2744 2257
rect 2738 2252 2744 2253
rect 2580 2183 2582 2252
rect 2740 2183 2742 2252
rect 2850 2207 2856 2208
rect 2850 2203 2851 2207
rect 2855 2203 2856 2207
rect 2850 2202 2856 2203
rect 2579 2182 2583 2183
rect 2579 2177 2583 2178
rect 2731 2182 2735 2183
rect 2731 2177 2735 2178
rect 2739 2182 2743 2183
rect 2739 2177 2743 2178
rect 2538 2175 2544 2176
rect 2538 2171 2539 2175
rect 2543 2171 2544 2175
rect 2538 2170 2544 2171
rect 2538 2163 2544 2164
rect 2538 2159 2539 2163
rect 2543 2159 2544 2163
rect 2538 2158 2544 2159
rect 2530 2115 2536 2116
rect 2530 2111 2531 2115
rect 2535 2111 2536 2115
rect 2530 2110 2536 2111
rect 2358 2100 2364 2101
rect 2540 2100 2542 2158
rect 2732 2116 2734 2177
rect 2738 2163 2744 2164
rect 2738 2159 2739 2163
rect 2743 2159 2744 2163
rect 2738 2158 2744 2159
rect 2730 2115 2736 2116
rect 2730 2111 2731 2115
rect 2735 2111 2736 2115
rect 2730 2110 2736 2111
rect 2558 2100 2564 2101
rect 2740 2100 2742 2158
rect 2758 2100 2764 2101
rect 2852 2100 2854 2202
rect 2860 2200 2862 2266
rect 2898 2257 2904 2258
rect 2898 2253 2899 2257
rect 2903 2253 2904 2257
rect 2898 2252 2904 2253
rect 2858 2199 2864 2200
rect 2858 2195 2859 2199
rect 2863 2195 2864 2199
rect 2858 2194 2864 2195
rect 2900 2183 2902 2252
rect 2899 2182 2903 2183
rect 2899 2177 2903 2178
rect 2923 2182 2927 2183
rect 2923 2177 2927 2178
rect 2924 2116 2926 2177
rect 3020 2168 3022 2266
rect 3050 2257 3056 2258
rect 3050 2253 3051 2257
rect 3055 2253 3056 2257
rect 3050 2252 3056 2253
rect 3052 2183 3054 2252
rect 3146 2239 3152 2240
rect 3146 2235 3147 2239
rect 3151 2235 3152 2239
rect 3146 2234 3152 2235
rect 3148 2208 3150 2234
rect 3146 2207 3152 2208
rect 3146 2203 3147 2207
rect 3151 2203 3152 2207
rect 3146 2202 3152 2203
rect 3176 2200 3178 2266
rect 3202 2257 3208 2258
rect 3202 2253 3203 2257
rect 3207 2253 3208 2257
rect 3202 2252 3208 2253
rect 3174 2199 3180 2200
rect 3174 2195 3175 2199
rect 3179 2195 3180 2199
rect 3174 2194 3180 2195
rect 3204 2183 3206 2252
rect 3328 2240 3330 2266
rect 3354 2257 3360 2258
rect 3354 2253 3355 2257
rect 3359 2253 3360 2257
rect 3354 2252 3360 2253
rect 3326 2239 3332 2240
rect 3326 2235 3327 2239
rect 3331 2235 3332 2239
rect 3326 2234 3332 2235
rect 3356 2183 3358 2252
rect 3422 2207 3428 2208
rect 3422 2203 3423 2207
rect 3427 2203 3428 2207
rect 3422 2202 3428 2203
rect 3051 2182 3055 2183
rect 3051 2177 3055 2178
rect 3115 2182 3119 2183
rect 3115 2177 3119 2178
rect 3203 2182 3207 2183
rect 3203 2177 3207 2178
rect 3299 2182 3303 2183
rect 3299 2177 3303 2178
rect 3355 2182 3359 2183
rect 3355 2177 3359 2178
rect 3018 2167 3024 2168
rect 3018 2163 3019 2167
rect 3023 2163 3024 2167
rect 3018 2162 3024 2163
rect 3116 2116 3118 2177
rect 3122 2163 3128 2164
rect 3122 2159 3123 2163
rect 3127 2159 3128 2163
rect 3122 2158 3128 2159
rect 2922 2115 2928 2116
rect 2922 2111 2923 2115
rect 2927 2111 2928 2115
rect 2922 2110 2928 2111
rect 3114 2115 3120 2116
rect 3114 2111 3115 2115
rect 3119 2111 3120 2115
rect 3114 2110 3120 2111
rect 2950 2100 2956 2101
rect 3124 2100 3126 2158
rect 3300 2116 3302 2177
rect 3298 2115 3304 2116
rect 3298 2111 3299 2115
rect 3303 2111 3304 2115
rect 3298 2110 3304 2111
rect 3142 2100 3148 2101
rect 3326 2100 3332 2101
rect 3424 2100 3426 2202
rect 3480 2200 3482 2266
rect 3514 2257 3520 2258
rect 3514 2253 3515 2257
rect 3519 2253 3520 2257
rect 3514 2252 3520 2253
rect 3478 2199 3484 2200
rect 3478 2195 3479 2199
rect 3483 2195 3484 2199
rect 3478 2194 3484 2195
rect 3516 2183 3518 2252
rect 3560 2208 3562 2338
rect 3679 2302 3683 2303
rect 3679 2297 3683 2298
rect 3680 2273 3682 2297
rect 3678 2272 3684 2273
rect 3792 2272 3794 2374
rect 3800 2361 3802 2421
rect 3840 2395 3842 2455
rect 3860 2395 3862 2456
rect 4060 2395 4062 2456
rect 4184 2404 4186 2470
rect 4387 2468 4391 2469
rect 4387 2463 4391 2464
rect 4290 2461 4296 2462
rect 4290 2457 4291 2461
rect 4295 2457 4296 2461
rect 4290 2456 4296 2457
rect 4210 2411 4216 2412
rect 4210 2407 4211 2411
rect 4215 2407 4216 2411
rect 4210 2406 4216 2407
rect 4182 2403 4188 2404
rect 4182 2399 4183 2403
rect 4187 2399 4188 2403
rect 4182 2398 4188 2399
rect 3839 2394 3843 2395
rect 3839 2389 3843 2390
rect 3859 2394 3863 2395
rect 3859 2389 3863 2390
rect 4059 2394 4063 2395
rect 4059 2389 4063 2390
rect 4091 2394 4095 2395
rect 4091 2389 4095 2390
rect 3798 2360 3804 2361
rect 3798 2356 3799 2360
rect 3803 2356 3804 2360
rect 3798 2355 3804 2356
rect 3798 2343 3804 2344
rect 3798 2339 3799 2343
rect 3803 2339 3804 2343
rect 3798 2338 3804 2339
rect 3800 2303 3802 2338
rect 3840 2329 3842 2389
rect 3838 2328 3844 2329
rect 3860 2328 3862 2389
rect 4092 2328 4094 2389
rect 4098 2375 4104 2376
rect 4098 2371 4099 2375
rect 4103 2371 4104 2375
rect 4098 2370 4104 2371
rect 3838 2324 3839 2328
rect 3843 2324 3844 2328
rect 3838 2323 3844 2324
rect 3858 2327 3864 2328
rect 3858 2323 3859 2327
rect 3863 2323 3864 2327
rect 3858 2322 3864 2323
rect 4090 2327 4096 2328
rect 4090 2323 4091 2327
rect 4095 2323 4096 2327
rect 4090 2322 4096 2323
rect 3886 2312 3892 2313
rect 4100 2312 4102 2370
rect 4118 2312 4124 2313
rect 4212 2312 4214 2406
rect 4292 2395 4294 2456
rect 4388 2412 4390 2463
rect 4440 2412 4442 2470
rect 4538 2461 4544 2462
rect 4538 2457 4539 2461
rect 4543 2457 4544 2461
rect 4538 2456 4544 2457
rect 4386 2411 4392 2412
rect 4386 2407 4387 2411
rect 4391 2407 4392 2411
rect 4386 2406 4392 2407
rect 4438 2411 4444 2412
rect 4438 2407 4439 2411
rect 4443 2407 4444 2411
rect 4438 2406 4444 2407
rect 4540 2395 4542 2456
rect 4712 2412 4714 2470
rect 4794 2461 4800 2462
rect 4794 2457 4795 2461
rect 4799 2457 4800 2461
rect 4794 2456 4800 2457
rect 4710 2411 4716 2412
rect 4710 2407 4711 2411
rect 4715 2407 4716 2411
rect 4710 2406 4716 2407
rect 4796 2395 4798 2456
rect 4976 2412 4978 2470
rect 5116 2469 5118 2534
rect 5296 2507 5298 2535
rect 5390 2534 5396 2535
rect 5295 2506 5299 2507
rect 5295 2501 5299 2502
rect 5351 2506 5355 2507
rect 5351 2501 5355 2502
rect 5352 2477 5354 2501
rect 5350 2476 5356 2477
rect 5444 2476 5446 2602
rect 5516 2556 5518 2617
rect 5636 2608 5638 2698
rect 5644 2640 5646 2770
rect 5664 2735 5666 2770
rect 5663 2734 5667 2735
rect 5663 2729 5667 2730
rect 5664 2706 5666 2729
rect 5662 2705 5668 2706
rect 5662 2701 5663 2705
rect 5667 2701 5668 2705
rect 5662 2700 5668 2701
rect 5662 2688 5668 2689
rect 5662 2684 5663 2688
rect 5667 2684 5668 2688
rect 5662 2683 5668 2684
rect 5642 2639 5648 2640
rect 5642 2635 5643 2639
rect 5647 2635 5648 2639
rect 5642 2634 5648 2635
rect 5664 2623 5666 2683
rect 5663 2622 5667 2623
rect 5663 2617 5667 2618
rect 5634 2607 5640 2608
rect 5634 2603 5635 2607
rect 5639 2603 5640 2607
rect 5634 2602 5640 2603
rect 5664 2557 5666 2617
rect 5662 2556 5668 2557
rect 5514 2555 5520 2556
rect 5514 2551 5515 2555
rect 5519 2551 5520 2555
rect 5662 2552 5663 2556
rect 5667 2552 5668 2556
rect 5662 2551 5668 2552
rect 5514 2550 5520 2551
rect 5542 2540 5548 2541
rect 5542 2536 5543 2540
rect 5547 2536 5548 2540
rect 5542 2535 5548 2536
rect 5634 2539 5640 2540
rect 5634 2535 5635 2539
rect 5639 2535 5640 2539
rect 5544 2507 5546 2535
rect 5634 2534 5640 2535
rect 5662 2539 5668 2540
rect 5662 2535 5663 2539
rect 5667 2535 5668 2539
rect 5662 2534 5668 2535
rect 5543 2506 5547 2507
rect 5543 2501 5547 2502
rect 5350 2472 5351 2476
rect 5355 2472 5356 2476
rect 5350 2471 5356 2472
rect 5442 2475 5448 2476
rect 5442 2471 5443 2475
rect 5447 2471 5448 2475
rect 5442 2470 5448 2471
rect 5115 2468 5119 2469
rect 5115 2463 5119 2464
rect 5058 2461 5064 2462
rect 5058 2457 5059 2461
rect 5063 2457 5064 2461
rect 5058 2456 5064 2457
rect 5322 2461 5328 2462
rect 5322 2457 5323 2461
rect 5327 2457 5328 2461
rect 5322 2456 5328 2457
rect 4974 2411 4980 2412
rect 4974 2407 4975 2411
rect 4979 2407 4980 2411
rect 4974 2406 4980 2407
rect 5060 2395 5062 2456
rect 5324 2395 5326 2456
rect 5406 2411 5412 2412
rect 5406 2407 5407 2411
rect 5411 2407 5412 2411
rect 5406 2406 5412 2407
rect 4291 2394 4295 2395
rect 4291 2389 4295 2390
rect 4339 2394 4343 2395
rect 4339 2389 4343 2390
rect 4539 2394 4543 2395
rect 4539 2389 4543 2390
rect 4579 2394 4583 2395
rect 4579 2389 4583 2390
rect 4795 2394 4799 2395
rect 4795 2389 4799 2390
rect 4811 2394 4815 2395
rect 4811 2389 4815 2390
rect 5043 2394 5047 2395
rect 5043 2389 5047 2390
rect 5059 2394 5063 2395
rect 5059 2389 5063 2390
rect 5283 2394 5287 2395
rect 5283 2389 5287 2390
rect 5323 2394 5327 2395
rect 5323 2389 5327 2390
rect 4340 2328 4342 2389
rect 4580 2328 4582 2389
rect 4586 2375 4592 2376
rect 4586 2371 4587 2375
rect 4591 2371 4592 2375
rect 4586 2370 4592 2371
rect 4338 2327 4344 2328
rect 4338 2323 4339 2327
rect 4343 2323 4344 2327
rect 4338 2322 4344 2323
rect 4578 2327 4584 2328
rect 4578 2323 4579 2327
rect 4583 2323 4584 2327
rect 4578 2322 4584 2323
rect 4366 2312 4372 2313
rect 4588 2312 4590 2370
rect 4812 2328 4814 2389
rect 4818 2375 4824 2376
rect 4818 2371 4819 2375
rect 4823 2371 4824 2375
rect 4818 2370 4824 2371
rect 4810 2327 4816 2328
rect 4810 2323 4811 2327
rect 4815 2323 4816 2327
rect 4810 2322 4816 2323
rect 4606 2312 4612 2313
rect 4820 2312 4822 2370
rect 5044 2328 5046 2389
rect 5050 2375 5056 2376
rect 5050 2371 5051 2375
rect 5055 2371 5056 2375
rect 5050 2370 5056 2371
rect 5042 2327 5048 2328
rect 5042 2323 5043 2327
rect 5047 2323 5048 2327
rect 5042 2322 5048 2323
rect 4838 2312 4844 2313
rect 5052 2312 5054 2370
rect 5284 2328 5286 2389
rect 5282 2327 5288 2328
rect 5282 2323 5283 2327
rect 5287 2323 5288 2327
rect 5282 2322 5288 2323
rect 5070 2312 5076 2313
rect 5310 2312 5316 2313
rect 5408 2312 5410 2406
rect 5515 2394 5519 2395
rect 5515 2389 5519 2390
rect 5498 2379 5504 2380
rect 5498 2375 5499 2379
rect 5503 2375 5504 2379
rect 5498 2374 5504 2375
rect 3838 2311 3844 2312
rect 3838 2307 3839 2311
rect 3843 2307 3844 2311
rect 3886 2308 3887 2312
rect 3891 2308 3892 2312
rect 3886 2307 3892 2308
rect 4098 2311 4104 2312
rect 4098 2307 4099 2311
rect 4103 2307 4104 2311
rect 4118 2308 4119 2312
rect 4123 2308 4124 2312
rect 4118 2307 4124 2308
rect 4210 2311 4216 2312
rect 4210 2307 4211 2311
rect 4215 2307 4216 2311
rect 4366 2308 4367 2312
rect 4371 2308 4372 2312
rect 4366 2307 4372 2308
rect 4586 2311 4592 2312
rect 4586 2307 4587 2311
rect 4591 2307 4592 2311
rect 4606 2308 4607 2312
rect 4611 2308 4612 2312
rect 4606 2307 4612 2308
rect 4818 2311 4824 2312
rect 4818 2307 4819 2311
rect 4823 2307 4824 2311
rect 4838 2308 4839 2312
rect 4843 2308 4844 2312
rect 4838 2307 4844 2308
rect 5050 2311 5056 2312
rect 5050 2307 5051 2311
rect 5055 2307 5056 2311
rect 5070 2308 5071 2312
rect 5075 2308 5076 2312
rect 5070 2307 5076 2308
rect 5166 2311 5172 2312
rect 5166 2307 5167 2311
rect 5171 2307 5172 2311
rect 5310 2308 5311 2312
rect 5315 2308 5316 2312
rect 5310 2307 5316 2308
rect 5406 2311 5412 2312
rect 5406 2307 5407 2311
rect 5411 2307 5412 2311
rect 3838 2306 3844 2307
rect 3799 2302 3803 2303
rect 3799 2297 3803 2298
rect 3800 2274 3802 2297
rect 3798 2273 3804 2274
rect 3642 2271 3648 2272
rect 3642 2267 3643 2271
rect 3647 2267 3648 2271
rect 3678 2268 3679 2272
rect 3683 2268 3684 2272
rect 3678 2267 3684 2268
rect 3790 2271 3796 2272
rect 3790 2267 3791 2271
rect 3795 2267 3796 2271
rect 3798 2269 3799 2273
rect 3803 2269 3804 2273
rect 3798 2268 3804 2269
rect 3642 2266 3648 2267
rect 3790 2266 3796 2267
rect 3644 2208 3646 2266
rect 3840 2259 3842 2306
rect 3888 2259 3890 2307
rect 4098 2306 4104 2307
rect 4120 2259 4122 2307
rect 4210 2306 4216 2307
rect 4368 2259 4370 2307
rect 4586 2306 4592 2307
rect 4608 2259 4610 2307
rect 4818 2306 4824 2307
rect 4840 2259 4842 2307
rect 5050 2306 5056 2307
rect 5072 2259 5074 2307
rect 5166 2306 5172 2307
rect 3839 2258 3843 2259
rect 3650 2257 3656 2258
rect 3650 2253 3651 2257
rect 3655 2253 3656 2257
rect 3650 2252 3656 2253
rect 3798 2256 3804 2257
rect 3798 2252 3799 2256
rect 3803 2252 3804 2256
rect 3839 2253 3843 2254
rect 3887 2258 3891 2259
rect 3887 2253 3891 2254
rect 4119 2258 4123 2259
rect 4119 2253 4123 2254
rect 4367 2258 4371 2259
rect 4367 2253 4371 2254
rect 4591 2258 4595 2259
rect 4591 2253 4595 2254
rect 4607 2258 4611 2259
rect 4607 2253 4611 2254
rect 4727 2258 4731 2259
rect 4727 2253 4731 2254
rect 4839 2258 4843 2259
rect 4839 2253 4843 2254
rect 4863 2258 4867 2259
rect 4863 2253 4867 2254
rect 4999 2258 5003 2259
rect 4999 2253 5003 2254
rect 5071 2258 5075 2259
rect 5071 2253 5075 2254
rect 5135 2258 5139 2259
rect 5135 2253 5139 2254
rect 3558 2207 3564 2208
rect 3558 2203 3559 2207
rect 3563 2203 3564 2207
rect 3558 2202 3564 2203
rect 3642 2207 3648 2208
rect 3642 2203 3643 2207
rect 3647 2203 3648 2207
rect 3642 2202 3648 2203
rect 3652 2183 3654 2252
rect 3798 2251 3804 2252
rect 3800 2183 3802 2251
rect 3840 2230 3842 2253
rect 3838 2229 3844 2230
rect 4592 2229 4594 2253
rect 4728 2229 4730 2253
rect 4864 2229 4866 2253
rect 5000 2229 5002 2253
rect 5136 2229 5138 2253
rect 3838 2225 3839 2229
rect 3843 2225 3844 2229
rect 3838 2224 3844 2225
rect 4590 2228 4596 2229
rect 4726 2228 4732 2229
rect 4862 2228 4868 2229
rect 4998 2228 5004 2229
rect 5134 2228 5140 2229
rect 4590 2224 4591 2228
rect 4595 2224 4596 2228
rect 4590 2223 4596 2224
rect 4690 2227 4696 2228
rect 4690 2223 4691 2227
rect 4695 2223 4696 2227
rect 4726 2224 4727 2228
rect 4731 2224 4732 2228
rect 4726 2223 4732 2224
rect 4826 2227 4832 2228
rect 4826 2223 4827 2227
rect 4831 2223 4832 2227
rect 4862 2224 4863 2228
rect 4867 2224 4868 2228
rect 4862 2223 4868 2224
rect 4962 2227 4968 2228
rect 4962 2223 4963 2227
rect 4967 2223 4968 2227
rect 4998 2224 4999 2228
rect 5003 2224 5004 2228
rect 4998 2223 5004 2224
rect 5098 2227 5104 2228
rect 5098 2223 5099 2227
rect 5103 2223 5104 2227
rect 5134 2224 5135 2228
rect 5139 2224 5140 2228
rect 5134 2223 5140 2224
rect 4690 2222 4696 2223
rect 4826 2222 4832 2223
rect 4962 2222 4968 2223
rect 5098 2222 5104 2223
rect 4562 2213 4568 2214
rect 3838 2212 3844 2213
rect 3838 2208 3839 2212
rect 3843 2208 3844 2212
rect 4562 2209 4563 2213
rect 4567 2209 4568 2213
rect 4562 2208 4568 2209
rect 3838 2207 3844 2208
rect 3483 2182 3487 2183
rect 3483 2177 3487 2178
rect 3515 2182 3519 2183
rect 3515 2177 3519 2178
rect 3651 2182 3655 2183
rect 3651 2177 3655 2178
rect 3799 2182 3803 2183
rect 3799 2177 3803 2178
rect 3484 2116 3486 2177
rect 3578 2163 3584 2164
rect 3578 2159 3579 2163
rect 3583 2159 3584 2163
rect 3578 2158 3584 2159
rect 3482 2115 3488 2116
rect 3482 2111 3483 2115
rect 3487 2111 3488 2115
rect 3482 2110 3488 2111
rect 3510 2100 3516 2101
rect 2158 2096 2159 2100
rect 2163 2096 2164 2100
rect 2158 2095 2164 2096
rect 2338 2099 2344 2100
rect 2338 2095 2339 2099
rect 2343 2095 2344 2099
rect 2358 2096 2359 2100
rect 2363 2096 2364 2100
rect 2358 2095 2364 2096
rect 2538 2099 2544 2100
rect 2538 2095 2539 2099
rect 2543 2095 2544 2099
rect 2558 2096 2559 2100
rect 2563 2096 2564 2100
rect 2558 2095 2564 2096
rect 2738 2099 2744 2100
rect 2738 2095 2739 2099
rect 2743 2095 2744 2099
rect 2758 2096 2759 2100
rect 2763 2096 2764 2100
rect 2758 2095 2764 2096
rect 2850 2099 2856 2100
rect 2850 2095 2851 2099
rect 2855 2095 2856 2099
rect 2950 2096 2951 2100
rect 2955 2096 2956 2100
rect 2950 2095 2956 2096
rect 3122 2099 3128 2100
rect 3122 2095 3123 2099
rect 3127 2095 3128 2099
rect 3142 2096 3143 2100
rect 3147 2096 3148 2100
rect 3142 2095 3148 2096
rect 3238 2099 3244 2100
rect 3238 2095 3239 2099
rect 3243 2095 3244 2099
rect 3326 2096 3327 2100
rect 3331 2096 3332 2100
rect 3326 2095 3332 2096
rect 3422 2099 3428 2100
rect 3422 2095 3423 2099
rect 3427 2095 3428 2099
rect 3510 2096 3511 2100
rect 3515 2096 3516 2100
rect 3510 2095 3516 2096
rect 2160 2063 2162 2095
rect 2338 2094 2344 2095
rect 2360 2063 2362 2095
rect 2538 2094 2544 2095
rect 2560 2063 2562 2095
rect 2738 2094 2744 2095
rect 2760 2063 2762 2095
rect 2850 2094 2856 2095
rect 2952 2063 2954 2095
rect 3122 2094 3128 2095
rect 3144 2063 3146 2095
rect 3238 2094 3244 2095
rect 2159 2062 2163 2063
rect 2159 2057 2163 2058
rect 2279 2062 2283 2063
rect 2279 2057 2283 2058
rect 2359 2062 2363 2063
rect 2359 2057 2363 2058
rect 2551 2062 2555 2063
rect 2551 2057 2555 2058
rect 2559 2062 2563 2063
rect 2559 2057 2563 2058
rect 2759 2062 2763 2063
rect 2759 2057 2763 2058
rect 2799 2062 2803 2063
rect 2799 2057 2803 2058
rect 2951 2062 2955 2063
rect 2951 2057 2955 2058
rect 3031 2062 3035 2063
rect 3031 2057 3035 2058
rect 3143 2062 3147 2063
rect 3143 2057 3147 2058
rect 2280 2033 2282 2057
rect 2552 2033 2554 2057
rect 2800 2033 2802 2057
rect 3032 2033 3034 2057
rect 2278 2032 2284 2033
rect 2550 2032 2556 2033
rect 2798 2032 2804 2033
rect 3030 2032 3036 2033
rect 2022 2028 2023 2032
rect 2027 2028 2028 2032
rect 2022 2027 2028 2028
rect 2118 2031 2124 2032
rect 2118 2027 2119 2031
rect 2123 2027 2124 2031
rect 2278 2028 2279 2032
rect 2283 2028 2284 2032
rect 2278 2027 2284 2028
rect 2374 2031 2380 2032
rect 2374 2027 2375 2031
rect 2379 2027 2380 2031
rect 2550 2028 2551 2032
rect 2555 2028 2556 2032
rect 2550 2027 2556 2028
rect 2646 2031 2652 2032
rect 2646 2027 2647 2031
rect 2651 2027 2652 2031
rect 2798 2028 2799 2032
rect 2803 2028 2804 2032
rect 2798 2027 2804 2028
rect 2890 2031 2896 2032
rect 2890 2027 2891 2031
rect 2895 2027 2896 2031
rect 3030 2028 3031 2032
rect 3035 2028 3036 2032
rect 3030 2027 3036 2028
rect 3122 2031 3128 2032
rect 3122 2027 3123 2031
rect 3127 2027 3128 2031
rect 2118 2026 2124 2027
rect 2374 2026 2380 2027
rect 2646 2026 2652 2027
rect 2890 2026 2896 2027
rect 3122 2026 3128 2027
rect 1934 2025 1940 2026
rect 1934 2021 1935 2025
rect 1939 2021 1940 2025
rect 1934 2020 1940 2021
rect 1994 2017 2000 2018
rect 1974 2016 1980 2017
rect 1974 2012 1975 2016
rect 1979 2012 1980 2016
rect 1994 2013 1995 2017
rect 1999 2013 2000 2017
rect 1994 2012 2000 2013
rect 2250 2017 2256 2018
rect 2250 2013 2251 2017
rect 2255 2013 2256 2017
rect 2250 2012 2256 2013
rect 1974 2011 1980 2012
rect 1934 2008 1940 2009
rect 1934 2004 1935 2008
rect 1939 2004 1940 2008
rect 1934 2003 1940 2004
rect 1910 1959 1916 1960
rect 1910 1955 1911 1959
rect 1915 1955 1916 1959
rect 1910 1954 1916 1955
rect 1936 1935 1938 2003
rect 1976 1939 1978 2011
rect 1996 1939 1998 2012
rect 2252 1939 2254 2012
rect 2376 1960 2378 2026
rect 2522 2017 2528 2018
rect 2522 2013 2523 2017
rect 2527 2013 2528 2017
rect 2522 2012 2528 2013
rect 2442 1967 2448 1968
rect 2442 1963 2443 1967
rect 2447 1963 2448 1967
rect 2442 1962 2448 1963
rect 2374 1959 2380 1960
rect 2374 1955 2375 1959
rect 2379 1955 2380 1959
rect 2374 1954 2380 1955
rect 1975 1938 1979 1939
rect 1523 1934 1527 1935
rect 1523 1929 1527 1930
rect 1579 1934 1583 1935
rect 1579 1929 1583 1930
rect 1771 1934 1775 1935
rect 1771 1929 1775 1930
rect 1787 1934 1791 1935
rect 1787 1929 1791 1930
rect 1935 1934 1939 1935
rect 1975 1933 1979 1934
rect 1995 1938 1999 1939
rect 1995 1933 1999 1934
rect 2251 1938 2255 1939
rect 2251 1933 2255 1934
rect 2315 1938 2319 1939
rect 2315 1933 2319 1934
rect 1935 1929 1939 1930
rect 1474 1919 1480 1920
rect 1474 1915 1475 1919
rect 1479 1915 1480 1919
rect 1474 1914 1480 1915
rect 1482 1919 1488 1920
rect 1482 1915 1483 1919
rect 1487 1915 1488 1919
rect 1482 1914 1488 1915
rect 1282 1867 1288 1868
rect 1282 1863 1283 1867
rect 1287 1863 1288 1867
rect 1282 1862 1288 1863
rect 1476 1860 1478 1914
rect 1524 1868 1526 1929
rect 1772 1868 1774 1929
rect 1778 1915 1784 1916
rect 1778 1911 1779 1915
rect 1783 1911 1784 1915
rect 1778 1910 1784 1911
rect 1522 1867 1528 1868
rect 1522 1863 1523 1867
rect 1527 1863 1528 1867
rect 1522 1862 1528 1863
rect 1770 1867 1776 1868
rect 1770 1863 1771 1867
rect 1775 1863 1776 1867
rect 1770 1862 1776 1863
rect 1474 1859 1480 1860
rect 1474 1855 1475 1859
rect 1479 1855 1480 1859
rect 1474 1854 1480 1855
rect 1078 1852 1084 1853
rect 1310 1852 1316 1853
rect 1550 1852 1556 1853
rect 1780 1852 1782 1910
rect 1936 1869 1938 1929
rect 1976 1873 1978 1933
rect 1974 1872 1980 1873
rect 1996 1872 1998 1933
rect 2206 1923 2212 1924
rect 2206 1919 2207 1923
rect 2211 1919 2212 1923
rect 2206 1918 2212 1919
rect 1934 1868 1940 1869
rect 1934 1864 1935 1868
rect 1939 1864 1940 1868
rect 1974 1868 1975 1872
rect 1979 1868 1980 1872
rect 1974 1867 1980 1868
rect 1994 1871 2000 1872
rect 1994 1867 1995 1871
rect 1999 1867 2000 1871
rect 1994 1866 2000 1867
rect 1934 1863 1940 1864
rect 2022 1856 2028 1857
rect 1974 1855 1980 1856
rect 1798 1852 1804 1853
rect 622 1848 623 1852
rect 627 1848 628 1852
rect 622 1847 628 1848
rect 826 1851 832 1852
rect 826 1847 827 1851
rect 831 1847 832 1851
rect 846 1848 847 1852
rect 851 1848 852 1852
rect 846 1847 852 1848
rect 1058 1851 1064 1852
rect 1058 1847 1059 1851
rect 1063 1847 1064 1851
rect 1078 1848 1079 1852
rect 1083 1848 1084 1852
rect 1078 1847 1084 1848
rect 1170 1851 1176 1852
rect 1170 1847 1171 1851
rect 1175 1847 1176 1851
rect 1310 1848 1311 1852
rect 1315 1848 1316 1852
rect 1310 1847 1316 1848
rect 1406 1851 1412 1852
rect 1406 1847 1407 1851
rect 1411 1847 1412 1851
rect 1550 1848 1551 1852
rect 1555 1848 1556 1852
rect 1550 1847 1556 1848
rect 1778 1851 1784 1852
rect 1778 1847 1779 1851
rect 1783 1847 1784 1851
rect 1798 1848 1799 1852
rect 1803 1848 1804 1852
rect 1798 1847 1804 1848
rect 1934 1851 1940 1852
rect 1934 1847 1935 1851
rect 1939 1847 1940 1851
rect 1974 1851 1975 1855
rect 1979 1851 1980 1855
rect 2022 1852 2023 1856
rect 2027 1852 2028 1856
rect 2022 1851 2028 1852
rect 1974 1850 1980 1851
rect 624 1807 626 1847
rect 826 1846 832 1847
rect 848 1807 850 1847
rect 1058 1846 1064 1847
rect 1080 1807 1082 1847
rect 1170 1846 1176 1847
rect 623 1806 627 1807
rect 623 1801 627 1802
rect 655 1806 659 1807
rect 655 1801 659 1802
rect 831 1806 835 1807
rect 831 1801 835 1802
rect 847 1806 851 1807
rect 847 1801 851 1802
rect 1007 1806 1011 1807
rect 1007 1801 1011 1802
rect 1079 1806 1083 1807
rect 1079 1801 1083 1802
rect 656 1777 658 1801
rect 832 1777 834 1801
rect 1008 1777 1010 1801
rect 654 1776 660 1777
rect 830 1776 836 1777
rect 1006 1776 1012 1777
rect 158 1772 159 1776
rect 163 1772 164 1776
rect 158 1771 164 1772
rect 266 1775 272 1776
rect 266 1771 267 1775
rect 271 1771 272 1775
rect 302 1772 303 1776
rect 307 1772 308 1776
rect 302 1771 308 1772
rect 418 1775 424 1776
rect 418 1771 419 1775
rect 423 1771 424 1775
rect 478 1772 479 1776
rect 483 1772 484 1776
rect 478 1771 484 1772
rect 574 1775 580 1776
rect 574 1771 575 1775
rect 579 1771 580 1775
rect 654 1772 655 1776
rect 659 1772 660 1776
rect 654 1771 660 1772
rect 770 1775 776 1776
rect 770 1771 771 1775
rect 775 1771 776 1775
rect 830 1772 831 1776
rect 835 1772 836 1776
rect 830 1771 836 1772
rect 926 1775 932 1776
rect 926 1771 927 1775
rect 931 1771 932 1775
rect 1006 1772 1007 1776
rect 1011 1772 1012 1776
rect 1006 1771 1012 1772
rect 1098 1775 1104 1776
rect 1098 1771 1099 1775
rect 1103 1771 1104 1775
rect 266 1770 272 1771
rect 418 1770 424 1771
rect 574 1770 580 1771
rect 770 1770 776 1771
rect 926 1770 932 1771
rect 1098 1770 1104 1771
rect 130 1761 136 1762
rect 110 1760 116 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 130 1757 131 1761
rect 135 1757 136 1761
rect 130 1756 136 1757
rect 110 1755 116 1756
rect 112 1691 114 1755
rect 132 1691 134 1756
rect 268 1712 270 1770
rect 274 1761 280 1762
rect 274 1757 275 1761
rect 279 1757 280 1761
rect 274 1756 280 1757
rect 250 1711 256 1712
rect 250 1707 251 1711
rect 255 1707 256 1711
rect 250 1706 256 1707
rect 266 1711 272 1712
rect 266 1707 267 1711
rect 271 1707 272 1711
rect 266 1706 272 1707
rect 111 1690 115 1691
rect 111 1685 115 1686
rect 131 1690 135 1691
rect 131 1685 135 1686
rect 112 1625 114 1685
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 110 1619 116 1620
rect 110 1607 116 1608
rect 110 1603 111 1607
rect 115 1603 116 1607
rect 110 1602 116 1603
rect 112 1559 114 1602
rect 111 1558 115 1559
rect 111 1553 115 1554
rect 159 1558 163 1559
rect 159 1553 163 1554
rect 112 1530 114 1553
rect 110 1529 116 1530
rect 160 1529 162 1553
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 158 1528 164 1529
rect 252 1528 254 1706
rect 276 1691 278 1756
rect 420 1712 422 1770
rect 450 1761 456 1762
rect 450 1757 451 1761
rect 455 1757 456 1761
rect 450 1756 456 1757
rect 626 1761 632 1762
rect 626 1757 627 1761
rect 631 1757 632 1761
rect 626 1756 632 1757
rect 418 1711 424 1712
rect 418 1707 419 1711
rect 423 1707 424 1711
rect 418 1706 424 1707
rect 452 1691 454 1756
rect 628 1691 630 1756
rect 722 1739 728 1740
rect 722 1735 723 1739
rect 727 1735 728 1739
rect 722 1734 728 1735
rect 724 1712 726 1734
rect 772 1712 774 1770
rect 802 1761 808 1762
rect 802 1757 803 1761
rect 807 1757 808 1761
rect 802 1756 808 1757
rect 722 1711 728 1712
rect 722 1707 723 1711
rect 727 1707 728 1711
rect 722 1706 728 1707
rect 770 1711 776 1712
rect 770 1707 771 1711
rect 775 1707 776 1711
rect 770 1706 776 1707
rect 804 1691 806 1756
rect 275 1690 279 1691
rect 275 1685 279 1686
rect 451 1690 455 1691
rect 451 1685 455 1686
rect 627 1690 631 1691
rect 627 1685 631 1686
rect 803 1690 807 1691
rect 803 1685 807 1686
rect 875 1690 879 1691
rect 875 1685 879 1686
rect 876 1624 878 1685
rect 928 1676 930 1770
rect 978 1761 984 1762
rect 978 1757 979 1761
rect 983 1757 984 1761
rect 978 1756 984 1757
rect 980 1691 982 1756
rect 1100 1740 1102 1770
rect 1154 1761 1160 1762
rect 1154 1757 1155 1761
rect 1159 1757 1160 1761
rect 1154 1756 1160 1757
rect 1098 1739 1104 1740
rect 1098 1735 1099 1739
rect 1103 1735 1104 1739
rect 1098 1734 1104 1735
rect 1156 1691 1158 1756
rect 1172 1704 1174 1846
rect 1312 1807 1314 1847
rect 1406 1846 1412 1847
rect 1183 1806 1187 1807
rect 1183 1801 1187 1802
rect 1311 1806 1315 1807
rect 1311 1801 1315 1802
rect 1359 1806 1363 1807
rect 1359 1801 1363 1802
rect 1184 1777 1186 1801
rect 1360 1777 1362 1801
rect 1182 1776 1188 1777
rect 1358 1776 1364 1777
rect 1182 1772 1183 1776
rect 1187 1772 1188 1776
rect 1182 1771 1188 1772
rect 1290 1775 1296 1776
rect 1290 1771 1291 1775
rect 1295 1771 1296 1775
rect 1358 1772 1359 1776
rect 1363 1772 1364 1776
rect 1358 1771 1364 1772
rect 1290 1770 1296 1771
rect 1170 1703 1176 1704
rect 1170 1699 1171 1703
rect 1175 1699 1176 1703
rect 1170 1698 1176 1699
rect 979 1690 983 1691
rect 979 1685 983 1686
rect 1011 1690 1015 1691
rect 1011 1685 1015 1686
rect 1147 1690 1151 1691
rect 1147 1685 1151 1686
rect 1155 1690 1159 1691
rect 1155 1685 1159 1686
rect 1283 1690 1287 1691
rect 1283 1685 1287 1686
rect 926 1675 932 1676
rect 926 1671 927 1675
rect 931 1671 932 1675
rect 926 1670 932 1671
rect 1012 1624 1014 1685
rect 1148 1624 1150 1685
rect 1266 1679 1272 1680
rect 1266 1675 1267 1679
rect 1271 1675 1272 1679
rect 1266 1674 1272 1675
rect 1242 1671 1248 1672
rect 1242 1667 1243 1671
rect 1247 1667 1248 1671
rect 1242 1666 1248 1667
rect 1244 1644 1246 1666
rect 1242 1643 1248 1644
rect 1242 1639 1243 1643
rect 1247 1639 1248 1643
rect 1242 1638 1248 1639
rect 874 1623 880 1624
rect 874 1619 875 1623
rect 879 1619 880 1623
rect 874 1618 880 1619
rect 1010 1623 1016 1624
rect 1010 1619 1011 1623
rect 1015 1619 1016 1623
rect 1010 1618 1016 1619
rect 1146 1623 1152 1624
rect 1146 1619 1147 1623
rect 1151 1619 1152 1623
rect 1146 1618 1152 1619
rect 902 1608 908 1609
rect 1038 1608 1044 1609
rect 1174 1608 1180 1609
rect 1268 1608 1270 1674
rect 1284 1624 1286 1685
rect 1292 1676 1294 1770
rect 1330 1761 1336 1762
rect 1330 1757 1331 1761
rect 1335 1757 1336 1761
rect 1330 1756 1336 1757
rect 1332 1691 1334 1756
rect 1408 1712 1410 1846
rect 1552 1807 1554 1847
rect 1778 1846 1784 1847
rect 1800 1807 1802 1847
rect 1934 1846 1940 1847
rect 1936 1807 1938 1846
rect 1976 1823 1978 1850
rect 2024 1823 2026 1851
rect 1975 1822 1979 1823
rect 1975 1817 1979 1818
rect 2023 1822 2027 1823
rect 2023 1817 2027 1818
rect 2111 1822 2115 1823
rect 2111 1817 2115 1818
rect 1535 1806 1539 1807
rect 1535 1801 1539 1802
rect 1551 1806 1555 1807
rect 1551 1801 1555 1802
rect 1711 1806 1715 1807
rect 1711 1801 1715 1802
rect 1799 1806 1803 1807
rect 1799 1801 1803 1802
rect 1935 1806 1939 1807
rect 1935 1801 1939 1802
rect 1536 1777 1538 1801
rect 1712 1777 1714 1801
rect 1936 1778 1938 1801
rect 1976 1794 1978 1817
rect 1974 1793 1980 1794
rect 2112 1793 2114 1817
rect 1974 1789 1975 1793
rect 1979 1789 1980 1793
rect 1974 1788 1980 1789
rect 2110 1792 2116 1793
rect 2208 1792 2210 1918
rect 2316 1872 2318 1933
rect 2322 1919 2328 1920
rect 2322 1915 2323 1919
rect 2327 1915 2328 1919
rect 2322 1914 2328 1915
rect 2314 1871 2320 1872
rect 2314 1867 2315 1871
rect 2319 1867 2320 1871
rect 2314 1866 2320 1867
rect 2324 1856 2326 1914
rect 2342 1856 2348 1857
rect 2444 1856 2446 1962
rect 2524 1939 2526 2012
rect 2648 1960 2650 2026
rect 2770 2017 2776 2018
rect 2770 2013 2771 2017
rect 2775 2013 2776 2017
rect 2770 2012 2776 2013
rect 2646 1959 2652 1960
rect 2646 1955 2647 1959
rect 2651 1955 2652 1959
rect 2646 1954 2652 1955
rect 2772 1939 2774 2012
rect 2866 2003 2872 2004
rect 2866 1999 2867 2003
rect 2871 1999 2872 2003
rect 2866 1998 2872 1999
rect 2868 1968 2870 1998
rect 2866 1967 2872 1968
rect 2866 1963 2867 1967
rect 2871 1963 2872 1967
rect 2866 1962 2872 1963
rect 2523 1938 2527 1939
rect 2523 1933 2527 1934
rect 2619 1938 2623 1939
rect 2619 1933 2623 1934
rect 2771 1938 2775 1939
rect 2771 1933 2775 1934
rect 2620 1872 2622 1933
rect 2892 1924 2894 2026
rect 3002 2017 3008 2018
rect 3002 2013 3003 2017
rect 3007 2013 3008 2017
rect 3002 2012 3008 2013
rect 3004 1939 3006 2012
rect 3124 2004 3126 2026
rect 3226 2017 3232 2018
rect 3226 2013 3227 2017
rect 3231 2013 3232 2017
rect 3226 2012 3232 2013
rect 3122 2003 3128 2004
rect 3122 1999 3123 2003
rect 3127 1999 3128 2003
rect 3122 1998 3128 1999
rect 3228 1939 3230 2012
rect 3240 1968 3242 2094
rect 3328 2063 3330 2095
rect 3422 2094 3428 2095
rect 3512 2063 3514 2095
rect 3255 2062 3259 2063
rect 3255 2057 3259 2058
rect 3327 2062 3331 2063
rect 3327 2057 3331 2058
rect 3479 2062 3483 2063
rect 3479 2057 3483 2058
rect 3511 2062 3515 2063
rect 3511 2057 3515 2058
rect 3256 2033 3258 2057
rect 3480 2033 3482 2057
rect 3254 2032 3260 2033
rect 3478 2032 3484 2033
rect 3580 2032 3582 2158
rect 3652 2116 3654 2177
rect 3774 2175 3780 2176
rect 3774 2171 3775 2175
rect 3779 2171 3780 2175
rect 3774 2170 3780 2171
rect 3658 2163 3664 2164
rect 3658 2159 3659 2163
rect 3663 2159 3664 2163
rect 3658 2158 3664 2159
rect 3650 2115 3656 2116
rect 3650 2111 3651 2115
rect 3655 2111 3656 2115
rect 3650 2110 3656 2111
rect 3660 2100 3662 2158
rect 3678 2100 3684 2101
rect 3776 2100 3778 2170
rect 3800 2117 3802 2177
rect 3840 2131 3842 2207
rect 4564 2131 4566 2208
rect 4692 2164 4694 2222
rect 4698 2213 4704 2214
rect 4698 2209 4699 2213
rect 4703 2209 4704 2213
rect 4698 2208 4704 2209
rect 4690 2163 4696 2164
rect 4690 2159 4691 2163
rect 4695 2159 4696 2163
rect 4690 2158 4696 2159
rect 4700 2131 4702 2208
rect 4828 2164 4830 2222
rect 4834 2213 4840 2214
rect 4834 2209 4835 2213
rect 4839 2209 4840 2213
rect 4834 2208 4840 2209
rect 4826 2163 4832 2164
rect 4826 2159 4827 2163
rect 4831 2159 4832 2163
rect 4826 2158 4832 2159
rect 4836 2131 4838 2208
rect 4964 2164 4966 2222
rect 4970 2213 4976 2214
rect 4970 2209 4971 2213
rect 4975 2209 4976 2213
rect 4970 2208 4976 2209
rect 4962 2163 4968 2164
rect 4962 2159 4963 2163
rect 4967 2159 4968 2163
rect 4962 2158 4968 2159
rect 4972 2131 4974 2208
rect 5100 2164 5102 2222
rect 5106 2213 5112 2214
rect 5106 2209 5107 2213
rect 5111 2209 5112 2213
rect 5106 2208 5112 2209
rect 5098 2163 5104 2164
rect 5098 2159 5099 2163
rect 5103 2159 5104 2163
rect 5098 2158 5104 2159
rect 5108 2131 5110 2208
rect 5168 2156 5170 2306
rect 5312 2259 5314 2307
rect 5406 2306 5412 2307
rect 5271 2258 5275 2259
rect 5271 2253 5275 2254
rect 5311 2258 5315 2259
rect 5311 2253 5315 2254
rect 5407 2258 5411 2259
rect 5407 2253 5411 2254
rect 5272 2229 5274 2253
rect 5408 2229 5410 2253
rect 5270 2228 5276 2229
rect 5406 2228 5412 2229
rect 5500 2228 5502 2374
rect 5516 2328 5518 2389
rect 5636 2380 5638 2534
rect 5664 2507 5666 2534
rect 5663 2506 5667 2507
rect 5663 2501 5667 2502
rect 5664 2478 5666 2501
rect 5662 2477 5668 2478
rect 5662 2473 5663 2477
rect 5667 2473 5668 2477
rect 5662 2472 5668 2473
rect 5662 2460 5668 2461
rect 5662 2456 5663 2460
rect 5667 2456 5668 2460
rect 5662 2455 5668 2456
rect 5664 2395 5666 2455
rect 5663 2394 5667 2395
rect 5663 2389 5667 2390
rect 5634 2379 5640 2380
rect 5634 2375 5635 2379
rect 5639 2375 5640 2379
rect 5634 2374 5640 2375
rect 5664 2329 5666 2389
rect 5662 2328 5668 2329
rect 5514 2327 5520 2328
rect 5514 2323 5515 2327
rect 5519 2323 5520 2327
rect 5662 2324 5663 2328
rect 5667 2324 5668 2328
rect 5662 2323 5668 2324
rect 5514 2322 5520 2323
rect 5542 2312 5548 2313
rect 5542 2308 5543 2312
rect 5547 2308 5548 2312
rect 5542 2307 5548 2308
rect 5634 2311 5640 2312
rect 5634 2307 5635 2311
rect 5639 2307 5640 2311
rect 5544 2259 5546 2307
rect 5634 2306 5640 2307
rect 5662 2311 5668 2312
rect 5662 2307 5663 2311
rect 5667 2307 5668 2311
rect 5662 2306 5668 2307
rect 5543 2258 5547 2259
rect 5543 2253 5547 2254
rect 5544 2229 5546 2253
rect 5542 2228 5548 2229
rect 5234 2227 5240 2228
rect 5234 2223 5235 2227
rect 5239 2223 5240 2227
rect 5270 2224 5271 2228
rect 5275 2224 5276 2228
rect 5270 2223 5276 2224
rect 5370 2227 5376 2228
rect 5370 2223 5371 2227
rect 5375 2223 5376 2227
rect 5406 2224 5407 2228
rect 5411 2224 5412 2228
rect 5406 2223 5412 2224
rect 5498 2227 5504 2228
rect 5498 2223 5499 2227
rect 5503 2223 5504 2227
rect 5542 2224 5543 2228
rect 5547 2224 5548 2228
rect 5542 2223 5548 2224
rect 5234 2222 5240 2223
rect 5370 2222 5376 2223
rect 5498 2222 5504 2223
rect 5236 2164 5238 2222
rect 5242 2213 5248 2214
rect 5242 2209 5243 2213
rect 5247 2209 5248 2213
rect 5242 2208 5248 2209
rect 5234 2163 5240 2164
rect 5234 2159 5235 2163
rect 5239 2159 5240 2163
rect 5234 2158 5240 2159
rect 5166 2155 5172 2156
rect 5166 2151 5167 2155
rect 5171 2151 5172 2155
rect 5166 2150 5172 2151
rect 5244 2131 5246 2208
rect 5372 2164 5374 2222
rect 5378 2213 5384 2214
rect 5378 2209 5379 2213
rect 5383 2209 5384 2213
rect 5378 2208 5384 2209
rect 5514 2213 5520 2214
rect 5514 2209 5515 2213
rect 5519 2209 5520 2213
rect 5514 2208 5520 2209
rect 5370 2163 5376 2164
rect 5370 2159 5371 2163
rect 5375 2159 5376 2163
rect 5370 2158 5376 2159
rect 5380 2131 5382 2208
rect 5516 2131 5518 2208
rect 5636 2164 5638 2306
rect 5664 2259 5666 2306
rect 5663 2258 5667 2259
rect 5663 2253 5667 2254
rect 5664 2230 5666 2253
rect 5662 2229 5668 2230
rect 5642 2227 5648 2228
rect 5642 2223 5643 2227
rect 5647 2223 5648 2227
rect 5662 2225 5663 2229
rect 5667 2225 5668 2229
rect 5662 2224 5668 2225
rect 5642 2222 5648 2223
rect 5634 2163 5640 2164
rect 5634 2159 5635 2163
rect 5639 2159 5640 2163
rect 5634 2158 5640 2159
rect 3839 2130 3843 2131
rect 3839 2125 3843 2126
rect 4563 2130 4567 2131
rect 4563 2125 4567 2126
rect 4699 2130 4703 2131
rect 4699 2125 4703 2126
rect 4835 2130 4839 2131
rect 4835 2125 4839 2126
rect 4955 2130 4959 2131
rect 4955 2125 4959 2126
rect 4971 2130 4975 2131
rect 4971 2125 4975 2126
rect 5091 2130 5095 2131
rect 5091 2125 5095 2126
rect 5107 2130 5111 2131
rect 5107 2125 5111 2126
rect 5227 2130 5231 2131
rect 5227 2125 5231 2126
rect 5243 2130 5247 2131
rect 5243 2125 5247 2126
rect 5379 2130 5383 2131
rect 5379 2125 5383 2126
rect 5515 2130 5519 2131
rect 5515 2125 5519 2126
rect 3798 2116 3804 2117
rect 3798 2112 3799 2116
rect 3803 2112 3804 2116
rect 3798 2111 3804 2112
rect 3658 2099 3664 2100
rect 3658 2095 3659 2099
rect 3663 2095 3664 2099
rect 3678 2096 3679 2100
rect 3683 2096 3684 2100
rect 3678 2095 3684 2096
rect 3774 2099 3780 2100
rect 3774 2095 3775 2099
rect 3779 2095 3780 2099
rect 3658 2094 3664 2095
rect 3680 2063 3682 2095
rect 3774 2094 3780 2095
rect 3798 2099 3804 2100
rect 3798 2095 3799 2099
rect 3803 2095 3804 2099
rect 3798 2094 3804 2095
rect 3800 2063 3802 2094
rect 3840 2065 3842 2125
rect 3838 2064 3844 2065
rect 4956 2064 4958 2125
rect 5082 2115 5088 2116
rect 5082 2111 5083 2115
rect 5087 2111 5088 2115
rect 5082 2110 5088 2111
rect 3679 2062 3683 2063
rect 3679 2057 3683 2058
rect 3799 2062 3803 2063
rect 3838 2060 3839 2064
rect 3843 2060 3844 2064
rect 3838 2059 3844 2060
rect 4954 2063 4960 2064
rect 4954 2059 4955 2063
rect 4959 2059 4960 2063
rect 4954 2058 4960 2059
rect 3799 2057 3803 2058
rect 3680 2033 3682 2057
rect 3800 2034 3802 2057
rect 5084 2056 5086 2110
rect 5092 2064 5094 2125
rect 5228 2064 5230 2125
rect 5350 2123 5356 2124
rect 5350 2119 5351 2123
rect 5355 2119 5356 2123
rect 5350 2118 5356 2119
rect 5090 2063 5096 2064
rect 5090 2059 5091 2063
rect 5095 2059 5096 2063
rect 5090 2058 5096 2059
rect 5226 2063 5232 2064
rect 5226 2059 5227 2063
rect 5231 2059 5232 2063
rect 5226 2058 5232 2059
rect 5082 2055 5088 2056
rect 5082 2051 5083 2055
rect 5087 2051 5088 2055
rect 5082 2050 5088 2051
rect 4982 2048 4988 2049
rect 5118 2048 5124 2049
rect 3838 2047 3844 2048
rect 3838 2043 3839 2047
rect 3843 2043 3844 2047
rect 4982 2044 4983 2048
rect 4987 2044 4988 2048
rect 4982 2043 4988 2044
rect 5074 2047 5080 2048
rect 5074 2043 5075 2047
rect 5079 2043 5080 2047
rect 5118 2044 5119 2048
rect 5123 2044 5124 2048
rect 5118 2043 5124 2044
rect 5254 2048 5260 2049
rect 5352 2048 5354 2118
rect 5410 2115 5416 2116
rect 5410 2111 5411 2115
rect 5415 2111 5416 2115
rect 5410 2110 5416 2111
rect 5254 2044 5255 2048
rect 5259 2044 5260 2048
rect 5254 2043 5260 2044
rect 5350 2047 5356 2048
rect 5350 2043 5351 2047
rect 5355 2043 5356 2047
rect 3838 2042 3844 2043
rect 3798 2033 3804 2034
rect 3678 2032 3684 2033
rect 3254 2028 3255 2032
rect 3259 2028 3260 2032
rect 3254 2027 3260 2028
rect 3350 2031 3356 2032
rect 3350 2027 3351 2031
rect 3355 2027 3356 2031
rect 3478 2028 3479 2032
rect 3483 2028 3484 2032
rect 3478 2027 3484 2028
rect 3578 2031 3584 2032
rect 3578 2027 3579 2031
rect 3583 2027 3584 2031
rect 3678 2028 3679 2032
rect 3683 2028 3684 2032
rect 3678 2027 3684 2028
rect 3770 2031 3776 2032
rect 3770 2027 3771 2031
rect 3775 2027 3776 2031
rect 3798 2029 3799 2033
rect 3803 2029 3804 2033
rect 3798 2028 3804 2029
rect 3350 2026 3356 2027
rect 3578 2026 3584 2027
rect 3770 2026 3776 2027
rect 3238 1967 3244 1968
rect 3238 1963 3239 1967
rect 3243 1963 3244 1967
rect 3238 1962 3244 1963
rect 3352 1960 3354 2026
rect 3450 2017 3456 2018
rect 3450 2013 3451 2017
rect 3455 2013 3456 2017
rect 3450 2012 3456 2013
rect 3650 2017 3656 2018
rect 3650 2013 3651 2017
rect 3655 2013 3656 2017
rect 3650 2012 3656 2013
rect 3350 1959 3356 1960
rect 3350 1955 3351 1959
rect 3355 1955 3356 1959
rect 3350 1954 3356 1955
rect 3452 1939 3454 2012
rect 3546 1999 3552 2000
rect 3546 1995 3547 1999
rect 3551 1995 3552 1999
rect 3546 1994 3552 1995
rect 3548 1968 3550 1994
rect 3546 1967 3552 1968
rect 3546 1963 3547 1967
rect 3551 1963 3552 1967
rect 3546 1962 3552 1963
rect 3652 1939 3654 2012
rect 3772 2000 3774 2026
rect 3840 2019 3842 2042
rect 4984 2019 4986 2043
rect 5074 2042 5080 2043
rect 3839 2018 3843 2019
rect 3798 2016 3804 2017
rect 3798 2012 3799 2016
rect 3803 2012 3804 2016
rect 3839 2013 3843 2014
rect 4727 2018 4731 2019
rect 4727 2013 4731 2014
rect 4863 2018 4867 2019
rect 4863 2013 4867 2014
rect 4983 2018 4987 2019
rect 4983 2013 4987 2014
rect 5007 2018 5011 2019
rect 5007 2013 5011 2014
rect 3798 2011 3804 2012
rect 3770 1999 3776 2000
rect 3770 1995 3771 1999
rect 3775 1995 3776 1999
rect 3770 1994 3776 1995
rect 3770 1967 3776 1968
rect 3770 1963 3771 1967
rect 3775 1963 3776 1967
rect 3770 1962 3776 1963
rect 2899 1938 2903 1939
rect 2899 1933 2903 1934
rect 3003 1938 3007 1939
rect 3003 1933 3007 1934
rect 3163 1938 3167 1939
rect 3163 1933 3167 1934
rect 3227 1938 3231 1939
rect 3227 1933 3231 1934
rect 3419 1938 3423 1939
rect 3419 1933 3423 1934
rect 3451 1938 3455 1939
rect 3451 1933 3455 1934
rect 3651 1938 3655 1939
rect 3651 1933 3655 1934
rect 2890 1923 2896 1924
rect 2890 1919 2891 1923
rect 2895 1919 2896 1923
rect 2890 1918 2896 1919
rect 2900 1872 2902 1933
rect 2906 1919 2912 1920
rect 2906 1915 2907 1919
rect 2911 1915 2912 1919
rect 2906 1914 2912 1915
rect 2618 1871 2624 1872
rect 2618 1867 2619 1871
rect 2623 1867 2624 1871
rect 2618 1866 2624 1867
rect 2898 1871 2904 1872
rect 2898 1867 2899 1871
rect 2903 1867 2904 1871
rect 2898 1866 2904 1867
rect 2646 1856 2652 1857
rect 2908 1856 2910 1914
rect 3164 1872 3166 1933
rect 3170 1919 3176 1920
rect 3170 1915 3171 1919
rect 3175 1915 3176 1919
rect 3170 1914 3176 1915
rect 3162 1871 3168 1872
rect 3162 1867 3163 1871
rect 3167 1867 3168 1871
rect 3162 1866 3168 1867
rect 2926 1856 2932 1857
rect 3172 1856 3174 1914
rect 3420 1872 3422 1933
rect 3534 1923 3540 1924
rect 3534 1919 3535 1923
rect 3539 1919 3540 1923
rect 3534 1918 3540 1919
rect 3418 1871 3424 1872
rect 3418 1867 3419 1871
rect 3423 1867 3424 1871
rect 3418 1866 3424 1867
rect 3190 1856 3196 1857
rect 3446 1856 3452 1857
rect 2322 1855 2328 1856
rect 2322 1851 2323 1855
rect 2327 1851 2328 1855
rect 2342 1852 2343 1856
rect 2347 1852 2348 1856
rect 2342 1851 2348 1852
rect 2442 1855 2448 1856
rect 2442 1851 2443 1855
rect 2447 1851 2448 1855
rect 2646 1852 2647 1856
rect 2651 1852 2652 1856
rect 2646 1851 2652 1852
rect 2906 1855 2912 1856
rect 2906 1851 2907 1855
rect 2911 1851 2912 1855
rect 2926 1852 2927 1856
rect 2931 1852 2932 1856
rect 2926 1851 2932 1852
rect 3170 1855 3176 1856
rect 3170 1851 3171 1855
rect 3175 1851 3176 1855
rect 3190 1852 3191 1856
rect 3195 1852 3196 1856
rect 3190 1851 3196 1852
rect 3286 1855 3292 1856
rect 3286 1851 3287 1855
rect 3291 1851 3292 1855
rect 3446 1852 3447 1856
rect 3451 1852 3452 1856
rect 3446 1851 3452 1852
rect 2322 1850 2328 1851
rect 2344 1823 2346 1851
rect 2442 1850 2448 1851
rect 2648 1823 2650 1851
rect 2906 1850 2912 1851
rect 2928 1823 2930 1851
rect 3170 1850 3176 1851
rect 3192 1823 3194 1851
rect 3286 1850 3292 1851
rect 2343 1822 2347 1823
rect 2343 1817 2347 1818
rect 2391 1822 2395 1823
rect 2391 1817 2395 1818
rect 2647 1822 2651 1823
rect 2647 1817 2651 1818
rect 2663 1822 2667 1823
rect 2663 1817 2667 1818
rect 2927 1822 2931 1823
rect 2927 1817 2931 1818
rect 3183 1822 3187 1823
rect 3183 1817 3187 1818
rect 3191 1822 3195 1823
rect 3191 1817 3195 1818
rect 2392 1793 2394 1817
rect 2664 1793 2666 1817
rect 2928 1793 2930 1817
rect 3184 1793 3186 1817
rect 2390 1792 2396 1793
rect 2662 1792 2668 1793
rect 2926 1792 2932 1793
rect 3182 1792 3188 1793
rect 2110 1788 2111 1792
rect 2115 1788 2116 1792
rect 2110 1787 2116 1788
rect 2206 1791 2212 1792
rect 2206 1787 2207 1791
rect 2211 1787 2212 1791
rect 2390 1788 2391 1792
rect 2395 1788 2396 1792
rect 2390 1787 2396 1788
rect 2486 1791 2492 1792
rect 2486 1787 2487 1791
rect 2491 1787 2492 1791
rect 2662 1788 2663 1792
rect 2667 1788 2668 1792
rect 2662 1787 2668 1788
rect 2754 1791 2760 1792
rect 2754 1787 2755 1791
rect 2759 1787 2760 1791
rect 2926 1788 2927 1792
rect 2931 1788 2932 1792
rect 2926 1787 2932 1788
rect 3018 1791 3024 1792
rect 3018 1787 3019 1791
rect 3023 1787 3024 1791
rect 3182 1788 3183 1792
rect 3187 1788 3188 1792
rect 3182 1787 3188 1788
rect 3278 1791 3284 1792
rect 3278 1787 3279 1791
rect 3283 1787 3284 1791
rect 2206 1786 2212 1787
rect 2486 1786 2492 1787
rect 2754 1786 2760 1787
rect 3018 1786 3024 1787
rect 3278 1786 3284 1787
rect 1934 1777 1940 1778
rect 2082 1777 2088 1778
rect 1534 1776 1540 1777
rect 1710 1776 1716 1777
rect 1470 1775 1476 1776
rect 1470 1771 1471 1775
rect 1475 1771 1476 1775
rect 1534 1772 1535 1776
rect 1539 1772 1540 1776
rect 1534 1771 1540 1772
rect 1646 1775 1652 1776
rect 1646 1771 1647 1775
rect 1651 1771 1652 1775
rect 1710 1772 1711 1776
rect 1715 1772 1716 1776
rect 1710 1771 1716 1772
rect 1806 1775 1812 1776
rect 1806 1771 1807 1775
rect 1811 1771 1812 1775
rect 1934 1773 1935 1777
rect 1939 1773 1940 1777
rect 1934 1772 1940 1773
rect 1974 1776 1980 1777
rect 1974 1772 1975 1776
rect 1979 1772 1980 1776
rect 2082 1773 2083 1777
rect 2087 1773 2088 1777
rect 2082 1772 2088 1773
rect 2362 1777 2368 1778
rect 2362 1773 2363 1777
rect 2367 1773 2368 1777
rect 2362 1772 2368 1773
rect 1974 1771 1980 1772
rect 1470 1770 1476 1771
rect 1646 1770 1652 1771
rect 1806 1770 1812 1771
rect 1472 1712 1474 1770
rect 1506 1761 1512 1762
rect 1506 1757 1507 1761
rect 1511 1757 1512 1761
rect 1506 1756 1512 1757
rect 1406 1711 1412 1712
rect 1406 1707 1407 1711
rect 1411 1707 1412 1711
rect 1406 1706 1412 1707
rect 1470 1711 1476 1712
rect 1470 1707 1471 1711
rect 1475 1707 1476 1711
rect 1470 1706 1476 1707
rect 1508 1691 1510 1756
rect 1648 1712 1650 1770
rect 1682 1761 1688 1762
rect 1682 1757 1683 1761
rect 1687 1757 1688 1761
rect 1682 1756 1688 1757
rect 1646 1711 1652 1712
rect 1646 1707 1647 1711
rect 1651 1707 1652 1711
rect 1646 1706 1652 1707
rect 1684 1691 1686 1756
rect 1808 1704 1810 1770
rect 1934 1760 1940 1761
rect 1934 1756 1935 1760
rect 1939 1756 1940 1760
rect 1934 1755 1940 1756
rect 1806 1703 1812 1704
rect 1806 1699 1807 1703
rect 1811 1699 1812 1703
rect 1806 1698 1812 1699
rect 1936 1691 1938 1755
rect 1331 1690 1335 1691
rect 1331 1685 1335 1686
rect 1419 1690 1423 1691
rect 1419 1685 1423 1686
rect 1507 1690 1511 1691
rect 1507 1685 1511 1686
rect 1555 1690 1559 1691
rect 1555 1685 1559 1686
rect 1683 1690 1687 1691
rect 1683 1685 1687 1686
rect 1935 1690 1939 1691
rect 1935 1685 1939 1686
rect 1290 1675 1296 1676
rect 1290 1671 1291 1675
rect 1295 1671 1296 1675
rect 1290 1670 1296 1671
rect 1420 1624 1422 1685
rect 1426 1671 1432 1672
rect 1426 1667 1427 1671
rect 1431 1667 1432 1671
rect 1426 1666 1432 1667
rect 1282 1623 1288 1624
rect 1282 1619 1283 1623
rect 1287 1619 1288 1623
rect 1282 1618 1288 1619
rect 1418 1623 1424 1624
rect 1418 1619 1419 1623
rect 1423 1619 1424 1623
rect 1418 1618 1424 1619
rect 1310 1608 1316 1609
rect 1428 1608 1430 1666
rect 1556 1624 1558 1685
rect 1562 1671 1568 1672
rect 1562 1667 1563 1671
rect 1567 1667 1568 1671
rect 1562 1666 1568 1667
rect 1554 1623 1560 1624
rect 1554 1619 1555 1623
rect 1559 1619 1560 1623
rect 1554 1618 1560 1619
rect 1446 1608 1452 1609
rect 1564 1608 1566 1666
rect 1678 1643 1684 1644
rect 1678 1639 1679 1643
rect 1683 1639 1684 1643
rect 1678 1638 1684 1639
rect 1582 1608 1588 1609
rect 1680 1608 1682 1638
rect 1936 1625 1938 1685
rect 1976 1679 1978 1771
rect 2084 1679 2086 1772
rect 2364 1679 2366 1772
rect 2488 1720 2490 1786
rect 2634 1777 2640 1778
rect 2634 1773 2635 1777
rect 2639 1773 2640 1777
rect 2634 1772 2640 1773
rect 2610 1727 2616 1728
rect 2610 1723 2611 1727
rect 2615 1723 2616 1727
rect 2610 1722 2616 1723
rect 2486 1719 2492 1720
rect 2486 1715 2487 1719
rect 2491 1715 2492 1719
rect 2486 1714 2492 1715
rect 1975 1678 1979 1679
rect 1975 1673 1979 1674
rect 2083 1678 2087 1679
rect 2083 1673 2087 1674
rect 2219 1678 2223 1679
rect 2219 1673 2223 1674
rect 2355 1678 2359 1679
rect 2355 1673 2359 1674
rect 2363 1678 2367 1679
rect 2363 1673 2367 1674
rect 2491 1678 2495 1679
rect 2491 1673 2495 1674
rect 1934 1624 1940 1625
rect 1934 1620 1935 1624
rect 1939 1620 1940 1624
rect 1934 1619 1940 1620
rect 1976 1613 1978 1673
rect 1974 1612 1980 1613
rect 2084 1612 2086 1673
rect 2178 1659 2184 1660
rect 2178 1655 2179 1659
rect 2183 1655 2184 1659
rect 2178 1654 2184 1655
rect 1974 1608 1975 1612
rect 1979 1608 1980 1612
rect 902 1604 903 1608
rect 907 1604 908 1608
rect 902 1603 908 1604
rect 998 1607 1004 1608
rect 998 1603 999 1607
rect 1003 1603 1004 1607
rect 1038 1604 1039 1608
rect 1043 1604 1044 1608
rect 1038 1603 1044 1604
rect 1134 1607 1140 1608
rect 1134 1603 1135 1607
rect 1139 1603 1140 1607
rect 1174 1604 1175 1608
rect 1179 1604 1180 1608
rect 1174 1603 1180 1604
rect 1266 1607 1272 1608
rect 1266 1603 1267 1607
rect 1271 1603 1272 1607
rect 1310 1604 1311 1608
rect 1315 1604 1316 1608
rect 1310 1603 1316 1604
rect 1426 1607 1432 1608
rect 1426 1603 1427 1607
rect 1431 1603 1432 1607
rect 1446 1604 1447 1608
rect 1451 1604 1452 1608
rect 1446 1603 1452 1604
rect 1562 1607 1568 1608
rect 1562 1603 1563 1607
rect 1567 1603 1568 1607
rect 1582 1604 1583 1608
rect 1587 1604 1588 1608
rect 1582 1603 1588 1604
rect 1678 1607 1684 1608
rect 1678 1603 1679 1607
rect 1683 1603 1684 1607
rect 904 1559 906 1603
rect 998 1602 1004 1603
rect 391 1558 395 1559
rect 391 1553 395 1554
rect 631 1558 635 1559
rect 631 1553 635 1554
rect 871 1558 875 1559
rect 871 1553 875 1554
rect 903 1558 907 1559
rect 903 1553 907 1554
rect 392 1529 394 1553
rect 632 1529 634 1553
rect 872 1529 874 1553
rect 390 1528 396 1529
rect 630 1528 636 1529
rect 870 1528 876 1529
rect 158 1524 159 1528
rect 163 1524 164 1528
rect 158 1523 164 1524
rect 250 1527 256 1528
rect 250 1523 251 1527
rect 255 1523 256 1527
rect 390 1524 391 1528
rect 395 1524 396 1528
rect 390 1523 396 1524
rect 518 1527 524 1528
rect 518 1523 519 1527
rect 523 1523 524 1527
rect 630 1524 631 1528
rect 635 1524 636 1528
rect 630 1523 636 1524
rect 730 1527 736 1528
rect 730 1523 731 1527
rect 735 1523 736 1527
rect 870 1524 871 1528
rect 875 1524 876 1528
rect 870 1523 876 1524
rect 990 1527 996 1528
rect 990 1523 991 1527
rect 995 1523 996 1527
rect 250 1522 256 1523
rect 518 1522 524 1523
rect 730 1522 736 1523
rect 990 1522 996 1523
rect 130 1513 136 1514
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 130 1509 131 1513
rect 135 1509 136 1513
rect 130 1508 136 1509
rect 362 1513 368 1514
rect 362 1509 363 1513
rect 367 1509 368 1513
rect 362 1508 368 1509
rect 110 1507 116 1508
rect 112 1435 114 1507
rect 132 1435 134 1508
rect 364 1435 366 1508
rect 458 1507 464 1508
rect 458 1503 459 1507
rect 463 1503 464 1507
rect 458 1502 464 1503
rect 460 1464 462 1502
rect 520 1464 522 1522
rect 602 1513 608 1514
rect 602 1509 603 1513
rect 607 1509 608 1513
rect 602 1508 608 1509
rect 458 1463 464 1464
rect 458 1459 459 1463
rect 463 1459 464 1463
rect 458 1458 464 1459
rect 518 1463 524 1464
rect 518 1459 519 1463
rect 523 1459 524 1463
rect 518 1458 524 1459
rect 454 1455 460 1456
rect 454 1451 455 1455
rect 459 1451 460 1455
rect 454 1450 460 1451
rect 111 1434 115 1435
rect 111 1429 115 1430
rect 131 1434 135 1435
rect 131 1429 135 1430
rect 331 1434 335 1435
rect 331 1429 335 1430
rect 363 1434 367 1435
rect 363 1429 367 1430
rect 112 1369 114 1429
rect 110 1368 116 1369
rect 132 1368 134 1429
rect 254 1419 260 1420
rect 254 1415 255 1419
rect 259 1415 260 1419
rect 254 1414 260 1415
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 130 1367 136 1368
rect 130 1363 131 1367
rect 135 1363 136 1367
rect 130 1362 136 1363
rect 158 1352 164 1353
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 158 1348 159 1352
rect 163 1348 164 1352
rect 158 1347 164 1348
rect 110 1346 116 1347
rect 112 1323 114 1346
rect 160 1323 162 1347
rect 111 1322 115 1323
rect 111 1317 115 1318
rect 159 1322 163 1323
rect 159 1317 163 1318
rect 112 1294 114 1317
rect 110 1293 116 1294
rect 160 1293 162 1317
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 158 1292 164 1293
rect 256 1292 258 1414
rect 332 1368 334 1429
rect 338 1415 344 1416
rect 338 1411 339 1415
rect 343 1411 344 1415
rect 338 1410 344 1411
rect 330 1367 336 1368
rect 330 1363 331 1367
rect 335 1363 336 1367
rect 330 1362 336 1363
rect 340 1352 342 1410
rect 358 1352 364 1353
rect 456 1352 458 1450
rect 604 1435 606 1508
rect 555 1434 559 1435
rect 555 1429 559 1430
rect 603 1434 607 1435
rect 603 1429 607 1430
rect 556 1368 558 1429
rect 732 1420 734 1522
rect 842 1513 848 1514
rect 842 1509 843 1513
rect 847 1509 848 1513
rect 842 1508 848 1509
rect 844 1435 846 1508
rect 779 1434 783 1435
rect 779 1429 783 1430
rect 843 1434 847 1435
rect 843 1429 847 1430
rect 730 1419 736 1420
rect 650 1415 656 1416
rect 650 1411 651 1415
rect 655 1411 656 1415
rect 730 1415 731 1419
rect 735 1415 736 1419
rect 730 1414 736 1415
rect 650 1410 656 1411
rect 652 1396 654 1410
rect 650 1395 656 1396
rect 650 1391 651 1395
rect 655 1391 656 1395
rect 650 1390 656 1391
rect 780 1368 782 1429
rect 992 1420 994 1522
rect 1000 1508 1002 1602
rect 1040 1559 1042 1603
rect 1134 1602 1140 1603
rect 1039 1558 1043 1559
rect 1039 1553 1043 1554
rect 1111 1558 1115 1559
rect 1111 1553 1115 1554
rect 1112 1529 1114 1553
rect 1110 1528 1116 1529
rect 1110 1524 1111 1528
rect 1115 1524 1116 1528
rect 1110 1523 1116 1524
rect 1082 1513 1088 1514
rect 1082 1509 1083 1513
rect 1087 1509 1088 1513
rect 1082 1508 1088 1509
rect 998 1507 1004 1508
rect 998 1503 999 1507
rect 1003 1503 1004 1507
rect 998 1502 1004 1503
rect 1084 1435 1086 1508
rect 1136 1464 1138 1602
rect 1176 1559 1178 1603
rect 1266 1602 1272 1603
rect 1312 1559 1314 1603
rect 1426 1602 1432 1603
rect 1448 1559 1450 1603
rect 1562 1602 1568 1603
rect 1584 1559 1586 1603
rect 1678 1602 1684 1603
rect 1934 1607 1940 1608
rect 1974 1607 1980 1608
rect 2082 1611 2088 1612
rect 2082 1607 2083 1611
rect 2087 1607 2088 1611
rect 1934 1603 1935 1607
rect 1939 1603 1940 1607
rect 2082 1606 2088 1607
rect 1934 1602 1940 1603
rect 1936 1559 1938 1602
rect 2110 1596 2116 1597
rect 1974 1595 1980 1596
rect 1974 1591 1975 1595
rect 1979 1591 1980 1595
rect 2110 1592 2111 1596
rect 2115 1592 2116 1596
rect 2110 1591 2116 1592
rect 1974 1590 1980 1591
rect 1976 1563 1978 1590
rect 2112 1563 2114 1591
rect 1975 1562 1979 1563
rect 1175 1558 1179 1559
rect 1175 1553 1179 1554
rect 1311 1558 1315 1559
rect 1311 1553 1315 1554
rect 1351 1558 1355 1559
rect 1351 1553 1355 1554
rect 1447 1558 1451 1559
rect 1447 1553 1451 1554
rect 1583 1558 1587 1559
rect 1583 1553 1587 1554
rect 1935 1558 1939 1559
rect 1975 1557 1979 1558
rect 2111 1562 2115 1563
rect 2111 1557 2115 1558
rect 2143 1562 2147 1563
rect 2143 1557 2147 1558
rect 1935 1553 1939 1554
rect 1352 1529 1354 1553
rect 1936 1530 1938 1553
rect 1976 1534 1978 1557
rect 1974 1533 1980 1534
rect 2144 1533 2146 1557
rect 2180 1548 2182 1654
rect 2220 1612 2222 1673
rect 2226 1659 2232 1660
rect 2226 1655 2227 1659
rect 2231 1655 2232 1659
rect 2226 1654 2232 1655
rect 2218 1611 2224 1612
rect 2218 1607 2219 1611
rect 2223 1607 2224 1611
rect 2218 1606 2224 1607
rect 2228 1596 2230 1654
rect 2356 1612 2358 1673
rect 2362 1659 2368 1660
rect 2362 1655 2363 1659
rect 2367 1655 2368 1659
rect 2362 1654 2368 1655
rect 2354 1611 2360 1612
rect 2354 1607 2355 1611
rect 2359 1607 2360 1611
rect 2354 1606 2360 1607
rect 2246 1596 2252 1597
rect 2364 1596 2366 1654
rect 2492 1612 2494 1673
rect 2498 1659 2504 1660
rect 2498 1655 2499 1659
rect 2503 1655 2504 1659
rect 2498 1654 2504 1655
rect 2490 1611 2496 1612
rect 2490 1607 2491 1611
rect 2495 1607 2496 1611
rect 2490 1606 2496 1607
rect 2382 1596 2388 1597
rect 2500 1596 2502 1654
rect 2518 1596 2524 1597
rect 2612 1596 2614 1722
rect 2636 1679 2638 1772
rect 2627 1678 2631 1679
rect 2627 1673 2631 1674
rect 2635 1678 2639 1679
rect 2635 1673 2639 1674
rect 2628 1612 2630 1673
rect 2756 1664 2758 1786
rect 2898 1777 2904 1778
rect 2898 1773 2899 1777
rect 2903 1773 2904 1777
rect 2898 1772 2904 1773
rect 2900 1679 2902 1772
rect 3020 1720 3022 1786
rect 3154 1777 3160 1778
rect 3154 1773 3155 1777
rect 3159 1773 3160 1777
rect 3154 1772 3160 1773
rect 3018 1719 3024 1720
rect 3018 1715 3019 1719
rect 3023 1715 3024 1719
rect 3018 1714 3024 1715
rect 3156 1679 3158 1772
rect 3280 1720 3282 1786
rect 3288 1728 3290 1850
rect 3448 1823 3450 1851
rect 3439 1822 3443 1823
rect 3439 1817 3443 1818
rect 3447 1822 3451 1823
rect 3447 1817 3451 1818
rect 3440 1793 3442 1817
rect 3438 1792 3444 1793
rect 3536 1792 3538 1918
rect 3652 1872 3654 1933
rect 3658 1919 3664 1920
rect 3658 1915 3659 1919
rect 3663 1915 3664 1919
rect 3658 1914 3664 1915
rect 3650 1871 3656 1872
rect 3650 1867 3651 1871
rect 3655 1867 3656 1871
rect 3650 1866 3656 1867
rect 3660 1856 3662 1914
rect 3678 1856 3684 1857
rect 3772 1856 3774 1962
rect 3800 1939 3802 2011
rect 3840 1990 3842 2013
rect 3838 1989 3844 1990
rect 4728 1989 4730 2013
rect 4864 1989 4866 2013
rect 5008 1989 5010 2013
rect 3838 1985 3839 1989
rect 3843 1985 3844 1989
rect 3838 1984 3844 1985
rect 4726 1988 4732 1989
rect 4862 1988 4868 1989
rect 5006 1988 5012 1989
rect 4726 1984 4727 1988
rect 4731 1984 4732 1988
rect 4726 1983 4732 1984
rect 4826 1987 4832 1988
rect 4826 1983 4827 1987
rect 4831 1983 4832 1987
rect 4862 1984 4863 1988
rect 4867 1984 4868 1988
rect 4862 1983 4868 1984
rect 4970 1987 4976 1988
rect 4970 1983 4971 1987
rect 4975 1983 4976 1987
rect 5006 1984 5007 1988
rect 5011 1984 5012 1988
rect 5006 1983 5012 1984
rect 4826 1982 4832 1983
rect 4970 1982 4976 1983
rect 4698 1973 4704 1974
rect 3838 1972 3844 1973
rect 3838 1968 3839 1972
rect 3843 1968 3844 1972
rect 4698 1969 4699 1973
rect 4703 1969 4704 1973
rect 4698 1968 4704 1969
rect 3838 1967 3844 1968
rect 3799 1938 3803 1939
rect 3799 1933 3803 1934
rect 3800 1873 3802 1933
rect 3840 1907 3842 1967
rect 4700 1907 4702 1968
rect 4828 1924 4830 1982
rect 4834 1973 4840 1974
rect 4834 1969 4835 1973
rect 4839 1969 4840 1973
rect 4834 1968 4840 1969
rect 4826 1923 4832 1924
rect 4826 1919 4827 1923
rect 4831 1919 4832 1923
rect 4826 1918 4832 1919
rect 4836 1907 4838 1968
rect 3839 1906 3843 1907
rect 3839 1901 3843 1902
rect 4275 1906 4279 1907
rect 4275 1901 4279 1902
rect 4499 1906 4503 1907
rect 4499 1901 4503 1902
rect 4699 1906 4703 1907
rect 4699 1901 4703 1902
rect 4731 1906 4735 1907
rect 4731 1901 4735 1902
rect 4835 1906 4839 1907
rect 4835 1901 4839 1902
rect 3798 1872 3804 1873
rect 3798 1868 3799 1872
rect 3803 1868 3804 1872
rect 3798 1867 3804 1868
rect 3658 1855 3664 1856
rect 3658 1851 3659 1855
rect 3663 1851 3664 1855
rect 3678 1852 3679 1856
rect 3683 1852 3684 1856
rect 3678 1851 3684 1852
rect 3770 1855 3776 1856
rect 3770 1851 3771 1855
rect 3775 1851 3776 1855
rect 3658 1850 3664 1851
rect 3680 1823 3682 1851
rect 3770 1850 3776 1851
rect 3798 1855 3804 1856
rect 3798 1851 3799 1855
rect 3803 1851 3804 1855
rect 3798 1850 3804 1851
rect 3800 1823 3802 1850
rect 3840 1841 3842 1901
rect 3838 1840 3844 1841
rect 4276 1840 4278 1901
rect 4490 1891 4496 1892
rect 4490 1887 4491 1891
rect 4495 1887 4496 1891
rect 4490 1886 4496 1887
rect 3838 1836 3839 1840
rect 3843 1836 3844 1840
rect 3838 1835 3844 1836
rect 4274 1839 4280 1840
rect 4274 1835 4275 1839
rect 4279 1835 4280 1839
rect 4274 1834 4280 1835
rect 4492 1832 4494 1886
rect 4500 1840 4502 1901
rect 4506 1887 4512 1888
rect 4506 1883 4507 1887
rect 4511 1883 4512 1887
rect 4506 1882 4512 1883
rect 4498 1839 4504 1840
rect 4498 1835 4499 1839
rect 4503 1835 4504 1839
rect 4498 1834 4504 1835
rect 4490 1831 4496 1832
rect 4490 1827 4491 1831
rect 4495 1827 4496 1831
rect 4490 1826 4496 1827
rect 4302 1824 4308 1825
rect 4508 1824 4510 1882
rect 4732 1840 4734 1901
rect 4972 1892 4974 1982
rect 4978 1973 4984 1974
rect 4978 1969 4979 1973
rect 4983 1969 4984 1973
rect 4978 1968 4984 1969
rect 4980 1907 4982 1968
rect 5076 1924 5078 2042
rect 5120 2019 5122 2043
rect 5256 2019 5258 2043
rect 5350 2042 5356 2043
rect 5119 2018 5123 2019
rect 5119 2013 5123 2014
rect 5159 2018 5163 2019
rect 5159 2013 5163 2014
rect 5255 2018 5259 2019
rect 5255 2013 5259 2014
rect 5319 2018 5323 2019
rect 5319 2013 5323 2014
rect 5160 1989 5162 2013
rect 5320 1989 5322 2013
rect 5158 1988 5164 1989
rect 5318 1988 5324 1989
rect 5412 1988 5414 2110
rect 5487 2018 5491 2019
rect 5487 2013 5491 2014
rect 5488 1989 5490 2013
rect 5486 1988 5492 1989
rect 5158 1984 5159 1988
rect 5163 1984 5164 1988
rect 5158 1983 5164 1984
rect 5250 1987 5256 1988
rect 5250 1983 5251 1987
rect 5255 1983 5256 1987
rect 5318 1984 5319 1988
rect 5323 1984 5324 1988
rect 5318 1983 5324 1984
rect 5410 1987 5416 1988
rect 5410 1983 5411 1987
rect 5415 1983 5416 1987
rect 5486 1984 5487 1988
rect 5491 1984 5492 1988
rect 5486 1983 5492 1984
rect 5582 1987 5588 1988
rect 5582 1983 5583 1987
rect 5587 1983 5588 1987
rect 5250 1982 5256 1983
rect 5410 1982 5416 1983
rect 5582 1982 5588 1983
rect 5130 1973 5136 1974
rect 5130 1969 5131 1973
rect 5135 1969 5136 1973
rect 5130 1968 5136 1969
rect 5074 1923 5080 1924
rect 5074 1919 5075 1923
rect 5079 1919 5080 1923
rect 5074 1918 5080 1919
rect 5132 1907 5134 1968
rect 5252 1916 5254 1982
rect 5290 1973 5296 1974
rect 5290 1969 5291 1973
rect 5295 1969 5296 1973
rect 5290 1968 5296 1969
rect 5458 1973 5464 1974
rect 5458 1969 5459 1973
rect 5463 1969 5464 1973
rect 5458 1968 5464 1969
rect 5250 1915 5256 1916
rect 5250 1911 5251 1915
rect 5255 1911 5256 1915
rect 5250 1910 5256 1911
rect 5292 1907 5294 1968
rect 5358 1923 5364 1924
rect 5358 1919 5359 1923
rect 5363 1919 5364 1923
rect 5358 1918 5364 1919
rect 4979 1906 4983 1907
rect 4979 1901 4983 1902
rect 5131 1906 5135 1907
rect 5131 1901 5135 1902
rect 5235 1906 5239 1907
rect 5235 1901 5239 1902
rect 5291 1906 5295 1907
rect 5291 1901 5295 1902
rect 4970 1891 4976 1892
rect 4738 1887 4744 1888
rect 4738 1883 4739 1887
rect 4743 1883 4744 1887
rect 4970 1887 4971 1891
rect 4975 1887 4976 1891
rect 4970 1886 4976 1887
rect 4738 1882 4744 1883
rect 4730 1839 4736 1840
rect 4730 1835 4731 1839
rect 4735 1835 4736 1839
rect 4730 1834 4736 1835
rect 4526 1824 4532 1825
rect 4740 1824 4742 1882
rect 4980 1840 4982 1901
rect 5236 1840 5238 1901
rect 5338 1891 5344 1892
rect 5338 1887 5339 1891
rect 5343 1887 5344 1891
rect 5338 1886 5344 1887
rect 4978 1839 4984 1840
rect 4978 1835 4979 1839
rect 4983 1835 4984 1839
rect 4978 1834 4984 1835
rect 5234 1839 5240 1840
rect 5234 1835 5235 1839
rect 5239 1835 5240 1839
rect 5234 1834 5240 1835
rect 4758 1824 4764 1825
rect 5006 1824 5012 1825
rect 3838 1823 3844 1824
rect 3679 1822 3683 1823
rect 3679 1817 3683 1818
rect 3799 1822 3803 1823
rect 3838 1819 3839 1823
rect 3843 1819 3844 1823
rect 4302 1820 4303 1824
rect 4307 1820 4308 1824
rect 4302 1819 4308 1820
rect 4506 1823 4512 1824
rect 4506 1819 4507 1823
rect 4511 1819 4512 1823
rect 4526 1820 4527 1824
rect 4531 1820 4532 1824
rect 4526 1819 4532 1820
rect 4738 1823 4744 1824
rect 4738 1819 4739 1823
rect 4743 1819 4744 1823
rect 4758 1820 4759 1824
rect 4763 1820 4764 1824
rect 4758 1819 4764 1820
rect 4858 1823 4864 1824
rect 4858 1819 4859 1823
rect 4863 1819 4864 1823
rect 5006 1820 5007 1824
rect 5011 1820 5012 1824
rect 5006 1819 5012 1820
rect 5262 1824 5268 1825
rect 5262 1820 5263 1824
rect 5267 1820 5268 1824
rect 5262 1819 5268 1820
rect 3838 1818 3844 1819
rect 3799 1817 3803 1818
rect 3680 1793 3682 1817
rect 3800 1794 3802 1817
rect 3798 1793 3804 1794
rect 3678 1792 3684 1793
rect 3438 1788 3439 1792
rect 3443 1788 3444 1792
rect 3438 1787 3444 1788
rect 3534 1791 3540 1792
rect 3534 1787 3535 1791
rect 3539 1787 3540 1791
rect 3678 1788 3679 1792
rect 3683 1788 3684 1792
rect 3678 1787 3684 1788
rect 3770 1791 3776 1792
rect 3770 1787 3771 1791
rect 3775 1787 3776 1791
rect 3798 1789 3799 1793
rect 3803 1789 3804 1793
rect 3798 1788 3804 1789
rect 3840 1787 3842 1818
rect 4304 1787 4306 1819
rect 4506 1818 4512 1819
rect 4528 1787 4530 1819
rect 4738 1818 4744 1819
rect 4760 1787 4762 1819
rect 4858 1818 4864 1819
rect 3534 1786 3540 1787
rect 3770 1786 3776 1787
rect 3839 1786 3843 1787
rect 3410 1777 3416 1778
rect 3410 1773 3411 1777
rect 3415 1773 3416 1777
rect 3410 1772 3416 1773
rect 3650 1777 3656 1778
rect 3650 1773 3651 1777
rect 3655 1773 3656 1777
rect 3650 1772 3656 1773
rect 3286 1727 3292 1728
rect 3286 1723 3287 1727
rect 3291 1723 3292 1727
rect 3286 1722 3292 1723
rect 3278 1719 3284 1720
rect 3278 1715 3279 1719
rect 3283 1715 3284 1719
rect 3278 1714 3284 1715
rect 3412 1679 3414 1772
rect 3652 1679 3654 1772
rect 3772 1720 3774 1786
rect 3839 1781 3843 1782
rect 3887 1786 3891 1787
rect 3887 1781 3891 1782
rect 4087 1786 4091 1787
rect 4087 1781 4091 1782
rect 4303 1786 4307 1787
rect 4303 1781 4307 1782
rect 4343 1786 4347 1787
rect 4343 1781 4347 1782
rect 4527 1786 4531 1787
rect 4527 1781 4531 1782
rect 4623 1786 4627 1787
rect 4623 1781 4627 1782
rect 4759 1786 4763 1787
rect 4759 1781 4763 1782
rect 3798 1776 3804 1777
rect 3798 1772 3799 1776
rect 3803 1772 3804 1776
rect 3798 1771 3804 1772
rect 3770 1719 3776 1720
rect 3770 1715 3771 1719
rect 3775 1715 3776 1719
rect 3770 1714 3776 1715
rect 3800 1679 3802 1771
rect 3840 1758 3842 1781
rect 3838 1757 3844 1758
rect 3888 1757 3890 1781
rect 4088 1757 4090 1781
rect 4344 1757 4346 1781
rect 4624 1757 4626 1781
rect 3838 1753 3839 1757
rect 3843 1753 3844 1757
rect 3838 1752 3844 1753
rect 3886 1756 3892 1757
rect 4086 1756 4092 1757
rect 4342 1756 4348 1757
rect 4622 1756 4628 1757
rect 3886 1752 3887 1756
rect 3891 1752 3892 1756
rect 3886 1751 3892 1752
rect 3982 1755 3988 1756
rect 3982 1751 3983 1755
rect 3987 1751 3988 1755
rect 4086 1752 4087 1756
rect 4091 1752 4092 1756
rect 4086 1751 4092 1752
rect 4222 1755 4228 1756
rect 4222 1751 4223 1755
rect 4227 1751 4228 1755
rect 4342 1752 4343 1756
rect 4347 1752 4348 1756
rect 4342 1751 4348 1752
rect 4434 1755 4440 1756
rect 4434 1751 4435 1755
rect 4439 1751 4440 1755
rect 4622 1752 4623 1756
rect 4627 1752 4628 1756
rect 4622 1751 4628 1752
rect 4714 1755 4720 1756
rect 4714 1751 4715 1755
rect 4719 1751 4720 1755
rect 3982 1750 3988 1751
rect 4222 1750 4228 1751
rect 4434 1750 4440 1751
rect 4714 1750 4720 1751
rect 3858 1741 3864 1742
rect 3838 1740 3844 1741
rect 3838 1736 3839 1740
rect 3843 1736 3844 1740
rect 3858 1737 3859 1741
rect 3863 1737 3864 1741
rect 3858 1736 3864 1737
rect 3838 1735 3844 1736
rect 2771 1678 2775 1679
rect 2771 1673 2775 1674
rect 2899 1678 2903 1679
rect 2899 1673 2903 1674
rect 2915 1678 2919 1679
rect 2915 1673 2919 1674
rect 3155 1678 3159 1679
rect 3155 1673 3159 1674
rect 3411 1678 3415 1679
rect 3411 1673 3415 1674
rect 3651 1678 3655 1679
rect 3651 1673 3655 1674
rect 3799 1678 3803 1679
rect 3799 1673 3803 1674
rect 2754 1663 2760 1664
rect 2754 1659 2755 1663
rect 2759 1659 2760 1663
rect 2754 1658 2760 1659
rect 2772 1612 2774 1673
rect 2778 1659 2784 1660
rect 2778 1655 2779 1659
rect 2783 1655 2784 1659
rect 2778 1654 2784 1655
rect 2626 1611 2632 1612
rect 2626 1607 2627 1611
rect 2631 1607 2632 1611
rect 2626 1606 2632 1607
rect 2770 1611 2776 1612
rect 2770 1607 2771 1611
rect 2775 1607 2776 1611
rect 2770 1606 2776 1607
rect 2654 1596 2660 1597
rect 2780 1596 2782 1654
rect 2916 1612 2918 1673
rect 2922 1659 2928 1660
rect 2922 1655 2923 1659
rect 2927 1655 2928 1659
rect 2922 1654 2928 1655
rect 2914 1611 2920 1612
rect 2914 1607 2915 1611
rect 2919 1607 2920 1611
rect 2914 1606 2920 1607
rect 2798 1596 2804 1597
rect 2924 1596 2926 1654
rect 3800 1613 3802 1673
rect 3840 1671 3842 1735
rect 3860 1671 3862 1736
rect 3984 1728 3986 1750
rect 4058 1741 4064 1742
rect 4058 1737 4059 1741
rect 4063 1737 4064 1741
rect 4058 1736 4064 1737
rect 3982 1727 3988 1728
rect 3982 1723 3983 1727
rect 3987 1723 3988 1727
rect 3982 1722 3988 1723
rect 3978 1691 3984 1692
rect 3978 1687 3979 1691
rect 3983 1687 3984 1691
rect 3978 1686 3984 1687
rect 3839 1670 3843 1671
rect 3839 1665 3843 1666
rect 3859 1670 3863 1671
rect 3859 1665 3863 1666
rect 3798 1612 3804 1613
rect 3798 1608 3799 1612
rect 3803 1608 3804 1612
rect 3798 1607 3804 1608
rect 3840 1605 3842 1665
rect 3838 1604 3844 1605
rect 3860 1604 3862 1665
rect 3838 1600 3839 1604
rect 3843 1600 3844 1604
rect 3838 1599 3844 1600
rect 3858 1603 3864 1604
rect 3858 1599 3859 1603
rect 3863 1599 3864 1603
rect 3858 1598 3864 1599
rect 2942 1596 2948 1597
rect 2226 1595 2232 1596
rect 2226 1591 2227 1595
rect 2231 1591 2232 1595
rect 2246 1592 2247 1596
rect 2251 1592 2252 1596
rect 2246 1591 2252 1592
rect 2362 1595 2368 1596
rect 2362 1591 2363 1595
rect 2367 1591 2368 1595
rect 2382 1592 2383 1596
rect 2387 1592 2388 1596
rect 2382 1591 2388 1592
rect 2498 1595 2504 1596
rect 2498 1591 2499 1595
rect 2503 1591 2504 1595
rect 2518 1592 2519 1596
rect 2523 1592 2524 1596
rect 2518 1591 2524 1592
rect 2610 1595 2616 1596
rect 2610 1591 2611 1595
rect 2615 1591 2616 1595
rect 2654 1592 2655 1596
rect 2659 1592 2660 1596
rect 2654 1591 2660 1592
rect 2778 1595 2784 1596
rect 2778 1591 2779 1595
rect 2783 1591 2784 1595
rect 2798 1592 2799 1596
rect 2803 1592 2804 1596
rect 2798 1591 2804 1592
rect 2922 1595 2928 1596
rect 2922 1591 2923 1595
rect 2927 1591 2928 1595
rect 2942 1592 2943 1596
rect 2947 1592 2948 1596
rect 2942 1591 2948 1592
rect 3038 1595 3044 1596
rect 3038 1591 3039 1595
rect 3043 1591 3044 1595
rect 2226 1590 2232 1591
rect 2248 1563 2250 1591
rect 2362 1590 2368 1591
rect 2384 1563 2386 1591
rect 2498 1590 2504 1591
rect 2520 1563 2522 1591
rect 2610 1590 2616 1591
rect 2656 1563 2658 1591
rect 2778 1590 2784 1591
rect 2800 1563 2802 1591
rect 2922 1590 2928 1591
rect 2944 1563 2946 1591
rect 3038 1590 3044 1591
rect 3798 1595 3804 1596
rect 3798 1591 3799 1595
rect 3803 1591 3804 1595
rect 3798 1590 3804 1591
rect 2247 1562 2251 1563
rect 2247 1557 2251 1558
rect 2279 1562 2283 1563
rect 2279 1557 2283 1558
rect 2383 1562 2387 1563
rect 2383 1557 2387 1558
rect 2415 1562 2419 1563
rect 2415 1557 2419 1558
rect 2519 1562 2523 1563
rect 2519 1557 2523 1558
rect 2551 1562 2555 1563
rect 2551 1557 2555 1558
rect 2655 1562 2659 1563
rect 2655 1557 2659 1558
rect 2687 1562 2691 1563
rect 2687 1557 2691 1558
rect 2799 1562 2803 1563
rect 2799 1557 2803 1558
rect 2823 1562 2827 1563
rect 2823 1557 2827 1558
rect 2943 1562 2947 1563
rect 2943 1557 2947 1558
rect 2959 1562 2963 1563
rect 2959 1557 2963 1558
rect 2178 1547 2184 1548
rect 2178 1543 2179 1547
rect 2183 1543 2184 1547
rect 2178 1542 2184 1543
rect 2280 1533 2282 1557
rect 2416 1533 2418 1557
rect 2552 1533 2554 1557
rect 2688 1533 2690 1557
rect 2824 1533 2826 1557
rect 2960 1533 2962 1557
rect 1934 1529 1940 1530
rect 1350 1528 1356 1529
rect 1350 1524 1351 1528
rect 1355 1524 1356 1528
rect 1350 1523 1356 1524
rect 1442 1527 1448 1528
rect 1442 1523 1443 1527
rect 1447 1523 1448 1527
rect 1934 1525 1935 1529
rect 1939 1525 1940 1529
rect 1974 1529 1975 1533
rect 1979 1529 1980 1533
rect 1974 1528 1980 1529
rect 2142 1532 2148 1533
rect 2142 1528 2143 1532
rect 2147 1528 2148 1532
rect 2142 1527 2148 1528
rect 2278 1532 2284 1533
rect 2414 1532 2420 1533
rect 2550 1532 2556 1533
rect 2686 1532 2692 1533
rect 2822 1532 2828 1533
rect 2958 1532 2964 1533
rect 2278 1528 2279 1532
rect 2283 1528 2284 1532
rect 2278 1527 2284 1528
rect 2374 1531 2380 1532
rect 2374 1527 2375 1531
rect 2379 1527 2380 1531
rect 2414 1528 2415 1532
rect 2419 1528 2420 1532
rect 2414 1527 2420 1528
rect 2514 1531 2520 1532
rect 2514 1527 2515 1531
rect 2519 1527 2520 1531
rect 2550 1528 2551 1532
rect 2555 1528 2556 1532
rect 2550 1527 2556 1528
rect 2650 1531 2656 1532
rect 2650 1527 2651 1531
rect 2655 1527 2656 1531
rect 2686 1528 2687 1532
rect 2691 1528 2692 1532
rect 2686 1527 2692 1528
rect 2786 1531 2792 1532
rect 2786 1527 2787 1531
rect 2791 1527 2792 1531
rect 2822 1528 2823 1532
rect 2827 1528 2828 1532
rect 2822 1527 2828 1528
rect 2914 1531 2920 1532
rect 2914 1527 2915 1531
rect 2919 1527 2920 1531
rect 2958 1528 2959 1532
rect 2963 1528 2964 1532
rect 2958 1527 2964 1528
rect 2374 1526 2380 1527
rect 2514 1526 2520 1527
rect 2650 1526 2656 1527
rect 2786 1526 2792 1527
rect 2914 1526 2920 1527
rect 1934 1524 1940 1525
rect 1442 1522 1448 1523
rect 1322 1513 1328 1514
rect 1322 1509 1323 1513
rect 1327 1509 1328 1513
rect 1322 1508 1328 1509
rect 1134 1463 1140 1464
rect 1134 1459 1135 1463
rect 1139 1459 1140 1463
rect 1134 1458 1140 1459
rect 1324 1435 1326 1508
rect 1444 1456 1446 1522
rect 2114 1517 2120 1518
rect 1974 1516 1980 1517
rect 1934 1512 1940 1513
rect 1934 1508 1935 1512
rect 1939 1508 1940 1512
rect 1974 1512 1975 1516
rect 1979 1512 1980 1516
rect 2114 1513 2115 1517
rect 2119 1513 2120 1517
rect 2114 1512 2120 1513
rect 2250 1517 2256 1518
rect 2250 1513 2251 1517
rect 2255 1513 2256 1517
rect 2250 1512 2256 1513
rect 1974 1511 1980 1512
rect 1934 1507 1940 1508
rect 1442 1455 1448 1456
rect 1442 1451 1443 1455
rect 1447 1451 1448 1455
rect 1442 1450 1448 1451
rect 1936 1435 1938 1507
rect 1976 1435 1978 1511
rect 2116 1435 2118 1512
rect 2252 1435 2254 1512
rect 2346 1491 2352 1492
rect 2346 1487 2347 1491
rect 2351 1487 2352 1491
rect 2346 1486 2352 1487
rect 2348 1468 2350 1486
rect 2346 1467 2352 1468
rect 2346 1463 2347 1467
rect 2351 1463 2352 1467
rect 2346 1462 2352 1463
rect 2376 1460 2378 1526
rect 2386 1517 2392 1518
rect 2386 1513 2387 1517
rect 2391 1513 2392 1517
rect 2386 1512 2392 1513
rect 2374 1459 2380 1460
rect 2374 1455 2375 1459
rect 2379 1455 2380 1459
rect 2374 1454 2380 1455
rect 2388 1435 2390 1512
rect 2516 1468 2518 1526
rect 2522 1517 2528 1518
rect 2522 1513 2523 1517
rect 2527 1513 2528 1517
rect 2522 1512 2528 1513
rect 2514 1467 2520 1468
rect 2514 1463 2515 1467
rect 2519 1463 2520 1467
rect 2514 1462 2520 1463
rect 2524 1435 2526 1512
rect 2652 1468 2654 1526
rect 2658 1517 2664 1518
rect 2658 1513 2659 1517
rect 2663 1513 2664 1517
rect 2658 1512 2664 1513
rect 2650 1467 2656 1468
rect 2650 1463 2651 1467
rect 2655 1463 2656 1467
rect 2650 1462 2656 1463
rect 2660 1435 2662 1512
rect 2788 1468 2790 1526
rect 2794 1517 2800 1518
rect 2794 1513 2795 1517
rect 2799 1513 2800 1517
rect 2794 1512 2800 1513
rect 2786 1467 2792 1468
rect 2786 1463 2787 1467
rect 2791 1463 2792 1467
rect 2786 1462 2792 1463
rect 2796 1435 2798 1512
rect 2916 1492 2918 1526
rect 2930 1517 2936 1518
rect 2930 1513 2931 1517
rect 2935 1513 2936 1517
rect 2930 1512 2936 1513
rect 2914 1491 2920 1492
rect 2914 1487 2915 1491
rect 2919 1487 2920 1491
rect 2914 1486 2920 1487
rect 2814 1459 2820 1460
rect 2814 1455 2815 1459
rect 2819 1455 2820 1459
rect 2814 1454 2820 1455
rect 1003 1434 1007 1435
rect 1003 1429 1007 1430
rect 1083 1434 1087 1435
rect 1083 1429 1087 1430
rect 1323 1434 1327 1435
rect 1323 1429 1327 1430
rect 1935 1434 1939 1435
rect 1935 1429 1939 1430
rect 1975 1434 1979 1435
rect 1975 1429 1979 1430
rect 2099 1434 2103 1435
rect 2099 1429 2103 1430
rect 2115 1434 2119 1435
rect 2115 1429 2119 1430
rect 2243 1434 2247 1435
rect 2243 1429 2247 1430
rect 2251 1434 2255 1435
rect 2251 1429 2255 1430
rect 2387 1434 2391 1435
rect 2387 1429 2391 1430
rect 2523 1434 2527 1435
rect 2523 1429 2527 1430
rect 2539 1434 2543 1435
rect 2539 1429 2543 1430
rect 2659 1434 2663 1435
rect 2659 1429 2663 1430
rect 2691 1434 2695 1435
rect 2691 1429 2695 1430
rect 2795 1434 2799 1435
rect 2795 1429 2799 1430
rect 990 1419 996 1420
rect 990 1415 991 1419
rect 995 1415 996 1419
rect 990 1414 996 1415
rect 1004 1368 1006 1429
rect 1126 1395 1132 1396
rect 1126 1391 1127 1395
rect 1131 1391 1132 1395
rect 1126 1390 1132 1391
rect 554 1367 560 1368
rect 554 1363 555 1367
rect 559 1363 560 1367
rect 554 1362 560 1363
rect 778 1367 784 1368
rect 778 1363 779 1367
rect 783 1363 784 1367
rect 778 1362 784 1363
rect 1002 1367 1008 1368
rect 1002 1363 1003 1367
rect 1007 1363 1008 1367
rect 1002 1362 1008 1363
rect 582 1352 588 1353
rect 806 1352 812 1353
rect 1030 1352 1036 1353
rect 1128 1352 1130 1390
rect 1936 1369 1938 1429
rect 1976 1369 1978 1429
rect 1934 1368 1940 1369
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 1934 1363 1940 1364
rect 1974 1368 1980 1369
rect 2100 1368 2102 1429
rect 2194 1415 2200 1416
rect 2194 1411 2195 1415
rect 2199 1411 2200 1415
rect 2194 1410 2200 1411
rect 1974 1364 1975 1368
rect 1979 1364 1980 1368
rect 1974 1363 1980 1364
rect 2098 1367 2104 1368
rect 2098 1363 2099 1367
rect 2103 1363 2104 1367
rect 2098 1362 2104 1363
rect 2126 1352 2132 1353
rect 338 1351 344 1352
rect 338 1347 339 1351
rect 343 1347 344 1351
rect 358 1348 359 1352
rect 363 1348 364 1352
rect 358 1347 364 1348
rect 454 1351 460 1352
rect 454 1347 455 1351
rect 459 1347 460 1351
rect 582 1348 583 1352
rect 587 1348 588 1352
rect 582 1347 588 1348
rect 674 1351 680 1352
rect 674 1347 675 1351
rect 679 1347 680 1351
rect 806 1348 807 1352
rect 811 1348 812 1352
rect 806 1347 812 1348
rect 902 1351 908 1352
rect 902 1347 903 1351
rect 907 1347 908 1351
rect 1030 1348 1031 1352
rect 1035 1348 1036 1352
rect 1030 1347 1036 1348
rect 1126 1351 1132 1352
rect 1126 1347 1127 1351
rect 1131 1347 1132 1351
rect 338 1346 344 1347
rect 360 1323 362 1347
rect 454 1346 460 1347
rect 584 1323 586 1347
rect 674 1346 680 1347
rect 359 1322 363 1323
rect 359 1317 363 1318
rect 367 1322 371 1323
rect 367 1317 371 1318
rect 583 1322 587 1323
rect 583 1317 587 1318
rect 607 1322 611 1323
rect 607 1317 611 1318
rect 368 1293 370 1317
rect 608 1293 610 1317
rect 366 1292 372 1293
rect 606 1292 612 1293
rect 158 1288 159 1292
rect 163 1288 164 1292
rect 158 1287 164 1288
rect 254 1291 260 1292
rect 254 1287 255 1291
rect 259 1287 260 1291
rect 366 1288 367 1292
rect 371 1288 372 1292
rect 366 1287 372 1288
rect 462 1291 468 1292
rect 462 1287 463 1291
rect 467 1287 468 1291
rect 606 1288 607 1292
rect 611 1288 612 1292
rect 606 1287 612 1288
rect 254 1286 260 1287
rect 462 1286 468 1287
rect 130 1277 136 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 130 1273 131 1277
rect 135 1273 136 1277
rect 130 1272 136 1273
rect 338 1277 344 1278
rect 338 1273 339 1277
rect 343 1273 344 1277
rect 338 1272 344 1273
rect 110 1271 116 1272
rect 112 1199 114 1271
rect 132 1199 134 1272
rect 250 1227 256 1228
rect 250 1223 251 1227
rect 255 1223 256 1227
rect 250 1222 256 1223
rect 111 1198 115 1199
rect 111 1193 115 1194
rect 131 1198 135 1199
rect 131 1193 135 1194
rect 112 1133 114 1193
rect 110 1132 116 1133
rect 132 1132 134 1193
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 130 1131 136 1132
rect 130 1127 131 1131
rect 135 1127 136 1131
rect 130 1126 136 1127
rect 158 1116 164 1117
rect 252 1116 254 1222
rect 340 1199 342 1272
rect 275 1198 279 1199
rect 275 1193 279 1194
rect 339 1198 343 1199
rect 339 1193 343 1194
rect 443 1198 447 1199
rect 443 1193 447 1194
rect 266 1183 272 1184
rect 266 1179 267 1183
rect 271 1179 272 1183
rect 266 1178 272 1179
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 158 1112 159 1116
rect 163 1112 164 1116
rect 158 1111 164 1112
rect 250 1115 256 1116
rect 250 1111 251 1115
rect 255 1111 256 1115
rect 110 1110 116 1111
rect 112 1079 114 1110
rect 160 1079 162 1111
rect 250 1110 256 1111
rect 111 1078 115 1079
rect 111 1073 115 1074
rect 159 1078 163 1079
rect 159 1073 163 1074
rect 175 1078 179 1079
rect 175 1073 179 1074
rect 112 1050 114 1073
rect 110 1049 116 1050
rect 176 1049 178 1073
rect 110 1045 111 1049
rect 115 1045 116 1049
rect 110 1044 116 1045
rect 174 1048 180 1049
rect 268 1048 270 1178
rect 276 1132 278 1193
rect 370 1179 376 1180
rect 370 1175 371 1179
rect 375 1175 376 1179
rect 370 1174 376 1175
rect 372 1156 374 1174
rect 370 1155 376 1156
rect 370 1151 371 1155
rect 375 1151 376 1155
rect 370 1150 376 1151
rect 444 1132 446 1193
rect 464 1184 466 1286
rect 578 1277 584 1278
rect 578 1273 579 1277
rect 583 1273 584 1277
rect 578 1272 584 1273
rect 580 1199 582 1272
rect 676 1228 678 1346
rect 808 1323 810 1347
rect 902 1346 908 1347
rect 807 1322 811 1323
rect 807 1317 811 1318
rect 847 1322 851 1323
rect 847 1317 851 1318
rect 848 1293 850 1317
rect 846 1292 852 1293
rect 702 1291 708 1292
rect 702 1287 703 1291
rect 707 1287 708 1291
rect 846 1288 847 1292
rect 851 1288 852 1292
rect 846 1287 852 1288
rect 702 1286 708 1287
rect 674 1227 680 1228
rect 674 1223 675 1227
rect 679 1223 680 1227
rect 674 1222 680 1223
rect 704 1220 706 1286
rect 818 1277 824 1278
rect 818 1273 819 1277
rect 823 1273 824 1277
rect 818 1272 824 1273
rect 702 1219 708 1220
rect 702 1215 703 1219
rect 707 1215 708 1219
rect 702 1214 708 1215
rect 820 1199 822 1272
rect 904 1228 906 1346
rect 1032 1323 1034 1347
rect 1126 1346 1132 1347
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 1934 1346 1940 1347
rect 1974 1351 1980 1352
rect 1974 1347 1975 1351
rect 1979 1347 1980 1351
rect 2126 1348 2127 1352
rect 2131 1348 2132 1352
rect 2126 1347 2132 1348
rect 1974 1346 1980 1347
rect 1936 1323 1938 1346
rect 1031 1322 1035 1323
rect 1031 1317 1035 1318
rect 1087 1322 1091 1323
rect 1087 1317 1091 1318
rect 1935 1322 1939 1323
rect 1976 1319 1978 1346
rect 2128 1319 2130 1347
rect 2196 1320 2198 1410
rect 2244 1368 2246 1429
rect 2250 1415 2256 1416
rect 2250 1411 2251 1415
rect 2255 1411 2256 1415
rect 2250 1410 2256 1411
rect 2242 1367 2248 1368
rect 2242 1363 2243 1367
rect 2247 1363 2248 1367
rect 2242 1362 2248 1363
rect 2252 1352 2254 1410
rect 2388 1368 2390 1429
rect 2394 1415 2400 1416
rect 2394 1411 2395 1415
rect 2399 1411 2400 1415
rect 2394 1410 2400 1411
rect 2386 1367 2392 1368
rect 2386 1363 2387 1367
rect 2391 1363 2392 1367
rect 2386 1362 2392 1363
rect 2270 1352 2276 1353
rect 2396 1352 2398 1410
rect 2540 1368 2542 1429
rect 2546 1415 2552 1416
rect 2546 1411 2547 1415
rect 2551 1411 2552 1415
rect 2546 1410 2552 1411
rect 2538 1367 2544 1368
rect 2538 1363 2539 1367
rect 2543 1363 2544 1367
rect 2538 1362 2544 1363
rect 2414 1352 2420 1353
rect 2548 1352 2550 1410
rect 2692 1368 2694 1429
rect 2698 1415 2704 1416
rect 2698 1411 2699 1415
rect 2703 1411 2704 1415
rect 2698 1410 2704 1411
rect 2690 1367 2696 1368
rect 2690 1363 2691 1367
rect 2695 1363 2696 1367
rect 2690 1362 2696 1363
rect 2566 1352 2572 1353
rect 2700 1352 2702 1410
rect 2718 1352 2724 1353
rect 2816 1352 2818 1454
rect 2932 1435 2934 1512
rect 3040 1468 3042 1590
rect 3800 1563 3802 1590
rect 3886 1588 3892 1589
rect 3980 1588 3982 1686
rect 4060 1671 4062 1736
rect 4224 1692 4226 1750
rect 4314 1741 4320 1742
rect 4314 1737 4315 1741
rect 4319 1737 4320 1741
rect 4314 1736 4320 1737
rect 4222 1691 4228 1692
rect 4222 1687 4223 1691
rect 4227 1687 4228 1691
rect 4222 1686 4228 1687
rect 4316 1671 4318 1736
rect 3995 1670 3999 1671
rect 3995 1665 3999 1666
rect 4059 1670 4063 1671
rect 4059 1665 4063 1666
rect 4139 1670 4143 1671
rect 4139 1665 4143 1666
rect 4315 1670 4319 1671
rect 4315 1665 4319 1666
rect 4323 1670 4327 1671
rect 4323 1665 4327 1666
rect 3996 1604 3998 1665
rect 4002 1651 4008 1652
rect 4002 1647 4003 1651
rect 4007 1647 4008 1651
rect 4002 1646 4008 1647
rect 3994 1603 4000 1604
rect 3994 1599 3995 1603
rect 3999 1599 4000 1603
rect 3994 1598 4000 1599
rect 3838 1587 3844 1588
rect 3838 1583 3839 1587
rect 3843 1583 3844 1587
rect 3886 1584 3887 1588
rect 3891 1584 3892 1588
rect 3886 1583 3892 1584
rect 3978 1587 3984 1588
rect 3978 1583 3979 1587
rect 3983 1583 3984 1587
rect 3838 1582 3844 1583
rect 3095 1562 3099 1563
rect 3095 1557 3099 1558
rect 3231 1562 3235 1563
rect 3231 1557 3235 1558
rect 3799 1562 3803 1563
rect 3799 1557 3803 1558
rect 3096 1533 3098 1557
rect 3232 1533 3234 1557
rect 3800 1534 3802 1557
rect 3840 1555 3842 1582
rect 3888 1555 3890 1583
rect 3978 1582 3984 1583
rect 3839 1554 3843 1555
rect 3839 1549 3843 1550
rect 3887 1554 3891 1555
rect 3887 1549 3891 1550
rect 3798 1533 3804 1534
rect 3094 1532 3100 1533
rect 3230 1532 3236 1533
rect 3058 1531 3064 1532
rect 3058 1527 3059 1531
rect 3063 1527 3064 1531
rect 3094 1528 3095 1532
rect 3099 1528 3100 1532
rect 3094 1527 3100 1528
rect 3194 1531 3200 1532
rect 3194 1527 3195 1531
rect 3199 1527 3200 1531
rect 3230 1528 3231 1532
rect 3235 1528 3236 1532
rect 3230 1527 3236 1528
rect 3322 1531 3328 1532
rect 3322 1527 3323 1531
rect 3327 1527 3328 1531
rect 3798 1529 3799 1533
rect 3803 1529 3804 1533
rect 3798 1528 3804 1529
rect 3058 1526 3064 1527
rect 3194 1526 3200 1527
rect 3322 1526 3328 1527
rect 3840 1526 3842 1549
rect 3060 1468 3062 1526
rect 3066 1517 3072 1518
rect 3066 1513 3067 1517
rect 3071 1513 3072 1517
rect 3066 1512 3072 1513
rect 3038 1467 3044 1468
rect 3038 1463 3039 1467
rect 3043 1463 3044 1467
rect 3038 1462 3044 1463
rect 3058 1467 3064 1468
rect 3058 1463 3059 1467
rect 3063 1463 3064 1467
rect 3058 1462 3064 1463
rect 3068 1435 3070 1512
rect 3196 1468 3198 1526
rect 3202 1517 3208 1518
rect 3202 1513 3203 1517
rect 3207 1513 3208 1517
rect 3202 1512 3208 1513
rect 3194 1467 3200 1468
rect 3194 1463 3195 1467
rect 3199 1463 3200 1467
rect 3194 1462 3200 1463
rect 3204 1435 3206 1512
rect 2851 1434 2855 1435
rect 2851 1429 2855 1430
rect 2931 1434 2935 1435
rect 2931 1429 2935 1430
rect 3011 1434 3015 1435
rect 3011 1429 3015 1430
rect 3067 1434 3071 1435
rect 3067 1429 3071 1430
rect 3171 1434 3175 1435
rect 3171 1429 3175 1430
rect 3203 1434 3207 1435
rect 3203 1429 3207 1430
rect 2852 1368 2854 1429
rect 3012 1368 3014 1429
rect 3172 1368 3174 1429
rect 3324 1420 3326 1526
rect 3838 1525 3844 1526
rect 3888 1525 3890 1549
rect 3838 1521 3839 1525
rect 3843 1521 3844 1525
rect 3838 1520 3844 1521
rect 3886 1524 3892 1525
rect 4004 1524 4006 1646
rect 4140 1604 4142 1665
rect 4262 1659 4268 1660
rect 4262 1655 4263 1659
rect 4267 1655 4268 1659
rect 4262 1654 4268 1655
rect 4146 1651 4152 1652
rect 4146 1647 4147 1651
rect 4151 1647 4152 1651
rect 4146 1646 4152 1647
rect 4138 1603 4144 1604
rect 4138 1599 4139 1603
rect 4143 1599 4144 1603
rect 4138 1598 4144 1599
rect 4022 1588 4028 1589
rect 4148 1588 4150 1646
rect 4166 1588 4172 1589
rect 4264 1588 4266 1654
rect 4324 1604 4326 1665
rect 4436 1656 4438 1750
rect 4594 1741 4600 1742
rect 4594 1737 4595 1741
rect 4599 1737 4600 1741
rect 4594 1736 4600 1737
rect 4596 1671 4598 1736
rect 4716 1684 4718 1750
rect 4860 1692 4862 1818
rect 5008 1787 5010 1819
rect 5264 1787 5266 1819
rect 4927 1786 4931 1787
rect 4927 1781 4931 1782
rect 5007 1786 5011 1787
rect 5007 1781 5011 1782
rect 5247 1786 5251 1787
rect 5247 1781 5251 1782
rect 5263 1786 5267 1787
rect 5263 1781 5267 1782
rect 4928 1757 4930 1781
rect 5248 1757 5250 1781
rect 4926 1756 4932 1757
rect 5246 1756 5252 1757
rect 5340 1756 5342 1886
rect 5360 1824 5362 1918
rect 5460 1907 5462 1968
rect 5459 1906 5463 1907
rect 5459 1901 5463 1902
rect 5499 1906 5503 1907
rect 5499 1901 5503 1902
rect 5500 1840 5502 1901
rect 5584 1892 5586 1982
rect 5644 1933 5646 2222
rect 5662 2212 5668 2213
rect 5662 2208 5663 2212
rect 5667 2208 5668 2212
rect 5662 2207 5668 2208
rect 5664 2131 5666 2207
rect 5663 2130 5667 2131
rect 5663 2125 5667 2126
rect 5664 2065 5666 2125
rect 5662 2064 5668 2065
rect 5662 2060 5663 2064
rect 5667 2060 5668 2064
rect 5662 2059 5668 2060
rect 5662 2047 5668 2048
rect 5662 2043 5663 2047
rect 5667 2043 5668 2047
rect 5662 2042 5668 2043
rect 5664 2019 5666 2042
rect 5663 2018 5667 2019
rect 5663 2013 5667 2014
rect 5664 1990 5666 2013
rect 5662 1989 5668 1990
rect 5662 1985 5663 1989
rect 5667 1985 5668 1989
rect 5662 1984 5668 1985
rect 5662 1972 5668 1973
rect 5662 1968 5663 1972
rect 5667 1968 5668 1972
rect 5662 1967 5668 1968
rect 5644 1931 5650 1933
rect 5648 1924 5650 1931
rect 5646 1923 5652 1924
rect 5646 1919 5647 1923
rect 5651 1919 5652 1923
rect 5646 1918 5652 1919
rect 5664 1907 5666 1967
rect 5663 1906 5667 1907
rect 5663 1901 5667 1902
rect 5582 1891 5588 1892
rect 5582 1887 5583 1891
rect 5587 1887 5588 1891
rect 5582 1886 5588 1887
rect 5664 1841 5666 1901
rect 5662 1840 5668 1841
rect 5498 1839 5504 1840
rect 5498 1835 5499 1839
rect 5503 1835 5504 1839
rect 5662 1836 5663 1840
rect 5667 1836 5668 1840
rect 5662 1835 5668 1836
rect 5498 1834 5504 1835
rect 5526 1824 5532 1825
rect 5358 1823 5364 1824
rect 5358 1819 5359 1823
rect 5363 1819 5364 1823
rect 5526 1820 5527 1824
rect 5531 1820 5532 1824
rect 5526 1819 5532 1820
rect 5622 1823 5628 1824
rect 5622 1819 5623 1823
rect 5627 1819 5628 1823
rect 5358 1818 5364 1819
rect 5528 1787 5530 1819
rect 5622 1818 5628 1819
rect 5662 1823 5668 1824
rect 5662 1819 5663 1823
rect 5667 1819 5668 1823
rect 5662 1818 5668 1819
rect 5527 1786 5531 1787
rect 5527 1781 5531 1782
rect 5543 1786 5547 1787
rect 5543 1781 5547 1782
rect 5544 1757 5546 1781
rect 5542 1756 5548 1757
rect 4926 1752 4927 1756
rect 4931 1752 4932 1756
rect 4926 1751 4932 1752
rect 5022 1755 5028 1756
rect 5022 1751 5023 1755
rect 5027 1751 5028 1755
rect 5246 1752 5247 1756
rect 5251 1752 5252 1756
rect 5246 1751 5252 1752
rect 5338 1755 5344 1756
rect 5338 1751 5339 1755
rect 5343 1751 5344 1755
rect 5542 1752 5543 1756
rect 5547 1752 5548 1756
rect 5542 1751 5548 1752
rect 5022 1750 5028 1751
rect 5338 1750 5344 1751
rect 4898 1741 4904 1742
rect 4898 1737 4899 1741
rect 4903 1737 4904 1741
rect 4898 1736 4904 1737
rect 4858 1691 4864 1692
rect 4858 1687 4859 1691
rect 4863 1687 4864 1691
rect 4858 1686 4864 1687
rect 4714 1683 4720 1684
rect 4714 1679 4715 1683
rect 4719 1679 4720 1683
rect 4714 1678 4720 1679
rect 4900 1671 4902 1736
rect 5024 1684 5026 1750
rect 5218 1741 5224 1742
rect 5218 1737 5219 1741
rect 5223 1737 5224 1741
rect 5218 1736 5224 1737
rect 5514 1741 5520 1742
rect 5514 1737 5515 1741
rect 5519 1737 5520 1741
rect 5514 1736 5520 1737
rect 5022 1683 5028 1684
rect 5022 1679 5023 1683
rect 5027 1679 5028 1683
rect 5022 1678 5028 1679
rect 5220 1671 5222 1736
rect 5394 1691 5400 1692
rect 5394 1687 5395 1691
rect 5399 1687 5400 1691
rect 5394 1686 5400 1687
rect 4531 1670 4535 1671
rect 4531 1665 4535 1666
rect 4595 1670 4599 1671
rect 4595 1665 4599 1666
rect 4763 1670 4767 1671
rect 4763 1665 4767 1666
rect 4899 1670 4903 1671
rect 4899 1665 4903 1666
rect 5011 1670 5015 1671
rect 5011 1665 5015 1666
rect 5219 1670 5223 1671
rect 5219 1665 5223 1666
rect 5275 1670 5279 1671
rect 5275 1665 5279 1666
rect 4434 1655 4440 1656
rect 4434 1651 4435 1655
rect 4439 1651 4440 1655
rect 4434 1650 4440 1651
rect 4532 1604 4534 1665
rect 4538 1651 4544 1652
rect 4538 1647 4539 1651
rect 4543 1647 4544 1651
rect 4538 1646 4544 1647
rect 4322 1603 4328 1604
rect 4322 1599 4323 1603
rect 4327 1599 4328 1603
rect 4322 1598 4328 1599
rect 4530 1603 4536 1604
rect 4530 1599 4531 1603
rect 4535 1599 4536 1603
rect 4530 1598 4536 1599
rect 4350 1588 4356 1589
rect 4540 1588 4542 1646
rect 4764 1604 4766 1665
rect 4770 1651 4776 1652
rect 4770 1647 4771 1651
rect 4775 1647 4776 1651
rect 4770 1646 4776 1647
rect 4762 1603 4768 1604
rect 4762 1599 4763 1603
rect 4767 1599 4768 1603
rect 4762 1598 4768 1599
rect 4558 1588 4564 1589
rect 4772 1588 4774 1646
rect 5012 1604 5014 1665
rect 5018 1651 5024 1652
rect 5018 1647 5019 1651
rect 5023 1647 5024 1651
rect 5018 1646 5024 1647
rect 5010 1603 5016 1604
rect 5010 1599 5011 1603
rect 5015 1599 5016 1603
rect 5010 1598 5016 1599
rect 4790 1588 4796 1589
rect 5020 1588 5022 1646
rect 5276 1604 5278 1665
rect 5274 1603 5280 1604
rect 5274 1599 5275 1603
rect 5279 1599 5280 1603
rect 5274 1598 5280 1599
rect 5038 1588 5044 1589
rect 5302 1588 5308 1589
rect 5396 1588 5398 1686
rect 5516 1671 5518 1736
rect 5624 1692 5626 1818
rect 5664 1787 5666 1818
rect 5663 1786 5667 1787
rect 5663 1781 5667 1782
rect 5664 1758 5666 1781
rect 5662 1757 5668 1758
rect 5634 1755 5640 1756
rect 5634 1751 5635 1755
rect 5639 1751 5640 1755
rect 5662 1753 5663 1757
rect 5667 1753 5668 1757
rect 5662 1752 5668 1753
rect 5634 1750 5640 1751
rect 5622 1691 5628 1692
rect 5622 1687 5623 1691
rect 5627 1687 5628 1691
rect 5622 1686 5628 1687
rect 5515 1670 5519 1671
rect 5515 1665 5519 1666
rect 5402 1655 5408 1656
rect 5402 1651 5403 1655
rect 5407 1651 5408 1655
rect 5402 1650 5408 1651
rect 4022 1584 4023 1588
rect 4027 1584 4028 1588
rect 4022 1583 4028 1584
rect 4146 1587 4152 1588
rect 4146 1583 4147 1587
rect 4151 1583 4152 1587
rect 4166 1584 4167 1588
rect 4171 1584 4172 1588
rect 4166 1583 4172 1584
rect 4262 1587 4268 1588
rect 4262 1583 4263 1587
rect 4267 1583 4268 1587
rect 4350 1584 4351 1588
rect 4355 1584 4356 1588
rect 4350 1583 4356 1584
rect 4538 1587 4544 1588
rect 4538 1583 4539 1587
rect 4543 1583 4544 1587
rect 4558 1584 4559 1588
rect 4563 1584 4564 1588
rect 4558 1583 4564 1584
rect 4770 1587 4776 1588
rect 4770 1583 4771 1587
rect 4775 1583 4776 1587
rect 4790 1584 4791 1588
rect 4795 1584 4796 1588
rect 4790 1583 4796 1584
rect 5018 1587 5024 1588
rect 5018 1583 5019 1587
rect 5023 1583 5024 1587
rect 5038 1584 5039 1588
rect 5043 1584 5044 1588
rect 5038 1583 5044 1584
rect 5130 1587 5136 1588
rect 5130 1583 5131 1587
rect 5135 1583 5136 1587
rect 5302 1584 5303 1588
rect 5307 1584 5308 1588
rect 5302 1583 5308 1584
rect 5394 1587 5400 1588
rect 5394 1583 5395 1587
rect 5399 1583 5400 1587
rect 4024 1555 4026 1583
rect 4146 1582 4152 1583
rect 4168 1555 4170 1583
rect 4262 1582 4268 1583
rect 4352 1555 4354 1583
rect 4538 1582 4544 1583
rect 4560 1555 4562 1583
rect 4770 1582 4776 1583
rect 4792 1555 4794 1583
rect 5018 1582 5024 1583
rect 5040 1555 5042 1583
rect 5130 1582 5136 1583
rect 4023 1554 4027 1555
rect 4023 1549 4027 1550
rect 4111 1554 4115 1555
rect 4111 1549 4115 1550
rect 4167 1554 4171 1555
rect 4167 1549 4171 1550
rect 4343 1554 4347 1555
rect 4343 1549 4347 1550
rect 4351 1554 4355 1555
rect 4351 1549 4355 1550
rect 4559 1554 4563 1555
rect 4559 1549 4563 1550
rect 4575 1554 4579 1555
rect 4575 1549 4579 1550
rect 4791 1554 4795 1555
rect 4791 1549 4795 1550
rect 4815 1554 4819 1555
rect 4815 1549 4819 1550
rect 5039 1554 5043 1555
rect 5039 1549 5043 1550
rect 5063 1554 5067 1555
rect 5063 1549 5067 1550
rect 4112 1525 4114 1549
rect 4344 1525 4346 1549
rect 4576 1525 4578 1549
rect 4816 1525 4818 1549
rect 5064 1525 5066 1549
rect 4110 1524 4116 1525
rect 4342 1524 4348 1525
rect 3886 1520 3887 1524
rect 3891 1520 3892 1524
rect 3886 1519 3892 1520
rect 4002 1523 4008 1524
rect 4002 1519 4003 1523
rect 4007 1519 4008 1523
rect 4110 1520 4111 1524
rect 4115 1520 4116 1524
rect 4110 1519 4116 1520
rect 4206 1523 4212 1524
rect 4206 1519 4207 1523
rect 4211 1519 4212 1523
rect 4342 1520 4343 1524
rect 4347 1520 4348 1524
rect 4342 1519 4348 1520
rect 4574 1524 4580 1525
rect 4814 1524 4820 1525
rect 5062 1524 5068 1525
rect 4574 1520 4575 1524
rect 4579 1520 4580 1524
rect 4574 1519 4580 1520
rect 4702 1523 4708 1524
rect 4702 1519 4703 1523
rect 4707 1519 4708 1523
rect 4814 1520 4815 1524
rect 4819 1520 4820 1524
rect 4814 1519 4820 1520
rect 4950 1523 4956 1524
rect 4950 1519 4951 1523
rect 4955 1519 4956 1523
rect 5062 1520 5063 1524
rect 5067 1520 5068 1524
rect 5062 1519 5068 1520
rect 4002 1518 4008 1519
rect 4206 1518 4212 1519
rect 4702 1518 4708 1519
rect 4950 1518 4956 1519
rect 3798 1516 3804 1517
rect 3798 1512 3799 1516
rect 3803 1512 3804 1516
rect 3798 1511 3804 1512
rect 3800 1435 3802 1511
rect 3858 1509 3864 1510
rect 3838 1508 3844 1509
rect 3838 1504 3839 1508
rect 3843 1504 3844 1508
rect 3858 1505 3859 1509
rect 3863 1505 3864 1509
rect 3858 1504 3864 1505
rect 4082 1509 4088 1510
rect 4082 1505 4083 1509
rect 4087 1505 4088 1509
rect 4082 1504 4088 1505
rect 4208 1504 4210 1518
rect 4314 1509 4320 1510
rect 4314 1505 4315 1509
rect 4319 1505 4320 1509
rect 4314 1504 4320 1505
rect 4546 1509 4552 1510
rect 4546 1505 4547 1509
rect 4551 1505 4552 1509
rect 4546 1504 4552 1505
rect 3838 1503 3844 1504
rect 3840 1443 3842 1503
rect 3860 1443 3862 1504
rect 3954 1503 3960 1504
rect 3954 1499 3955 1503
rect 3959 1499 3960 1503
rect 3954 1498 3960 1499
rect 3956 1460 3958 1498
rect 3954 1459 3960 1460
rect 3954 1455 3955 1459
rect 3959 1455 3960 1459
rect 3954 1454 3960 1455
rect 4084 1443 4086 1504
rect 4206 1503 4212 1504
rect 4206 1499 4207 1503
rect 4211 1499 4212 1503
rect 4206 1498 4212 1499
rect 4202 1459 4208 1460
rect 4202 1455 4203 1459
rect 4207 1455 4208 1459
rect 4202 1454 4208 1455
rect 3839 1442 3843 1443
rect 3839 1437 3843 1438
rect 3859 1442 3863 1443
rect 3859 1437 3863 1438
rect 4083 1442 4087 1443
rect 4083 1437 4087 1438
rect 3799 1434 3803 1435
rect 3799 1429 3803 1430
rect 3322 1419 3328 1420
rect 3322 1415 3323 1419
rect 3327 1415 3328 1419
rect 3322 1414 3328 1415
rect 3800 1369 3802 1429
rect 3840 1377 3842 1437
rect 3838 1376 3844 1377
rect 3860 1376 3862 1437
rect 3982 1427 3988 1428
rect 3982 1423 3983 1427
rect 3987 1423 3988 1427
rect 3982 1422 3988 1423
rect 3838 1372 3839 1376
rect 3843 1372 3844 1376
rect 3838 1371 3844 1372
rect 3858 1375 3864 1376
rect 3858 1371 3859 1375
rect 3863 1371 3864 1375
rect 3858 1370 3864 1371
rect 3798 1368 3804 1369
rect 2850 1367 2856 1368
rect 2850 1363 2851 1367
rect 2855 1363 2856 1367
rect 2850 1362 2856 1363
rect 3010 1367 3016 1368
rect 3010 1363 3011 1367
rect 3015 1363 3016 1367
rect 3010 1362 3016 1363
rect 3170 1367 3176 1368
rect 3170 1363 3171 1367
rect 3175 1363 3176 1367
rect 3798 1364 3799 1368
rect 3803 1364 3804 1368
rect 3798 1363 3804 1364
rect 3170 1362 3176 1363
rect 3886 1360 3892 1361
rect 3838 1359 3844 1360
rect 3838 1355 3839 1359
rect 3843 1355 3844 1359
rect 3886 1356 3887 1360
rect 3891 1356 3892 1360
rect 3886 1355 3892 1356
rect 3838 1354 3844 1355
rect 2878 1352 2884 1353
rect 2250 1351 2256 1352
rect 2250 1347 2251 1351
rect 2255 1347 2256 1351
rect 2270 1348 2271 1352
rect 2275 1348 2276 1352
rect 2270 1347 2276 1348
rect 2394 1351 2400 1352
rect 2394 1347 2395 1351
rect 2399 1347 2400 1351
rect 2414 1348 2415 1352
rect 2419 1348 2420 1352
rect 2414 1347 2420 1348
rect 2546 1351 2552 1352
rect 2546 1347 2547 1351
rect 2551 1347 2552 1351
rect 2566 1348 2567 1352
rect 2571 1348 2572 1352
rect 2566 1347 2572 1348
rect 2698 1351 2704 1352
rect 2698 1347 2699 1351
rect 2703 1347 2704 1351
rect 2718 1348 2719 1352
rect 2723 1348 2724 1352
rect 2718 1347 2724 1348
rect 2814 1351 2820 1352
rect 2814 1347 2815 1351
rect 2819 1347 2820 1351
rect 2878 1348 2879 1352
rect 2883 1348 2884 1352
rect 2878 1347 2884 1348
rect 3038 1352 3044 1353
rect 3038 1348 3039 1352
rect 3043 1348 3044 1352
rect 3038 1347 3044 1348
rect 3198 1352 3204 1353
rect 3198 1348 3199 1352
rect 3203 1348 3204 1352
rect 3198 1347 3204 1348
rect 3798 1351 3804 1352
rect 3798 1347 3799 1351
rect 3803 1347 3804 1351
rect 2250 1346 2256 1347
rect 2194 1319 2200 1320
rect 2272 1319 2274 1347
rect 2394 1346 2400 1347
rect 2416 1319 2418 1347
rect 2546 1346 2552 1347
rect 2568 1319 2570 1347
rect 2698 1346 2704 1347
rect 2720 1319 2722 1347
rect 2814 1346 2820 1347
rect 2880 1319 2882 1347
rect 2886 1319 2892 1320
rect 3040 1319 3042 1347
rect 3200 1319 3202 1347
rect 3798 1346 3804 1347
rect 3800 1319 3802 1346
rect 3840 1331 3842 1354
rect 3888 1331 3890 1355
rect 3839 1330 3843 1331
rect 3839 1325 3843 1326
rect 3887 1330 3891 1331
rect 3887 1325 3891 1326
rect 1935 1317 1939 1318
rect 1975 1318 1979 1319
rect 1088 1293 1090 1317
rect 1936 1294 1938 1317
rect 1975 1313 1979 1314
rect 2023 1318 2027 1319
rect 2023 1313 2027 1314
rect 2127 1318 2131 1319
rect 2127 1313 2131 1314
rect 2175 1318 2179 1319
rect 2194 1315 2195 1319
rect 2199 1315 2200 1319
rect 2194 1314 2200 1315
rect 2271 1318 2275 1319
rect 2175 1313 2179 1314
rect 2271 1313 2275 1314
rect 2367 1318 2371 1319
rect 2367 1313 2371 1314
rect 2415 1318 2419 1319
rect 2415 1313 2419 1314
rect 2567 1318 2571 1319
rect 2567 1313 2571 1314
rect 2575 1318 2579 1319
rect 2575 1313 2579 1314
rect 2719 1318 2723 1319
rect 2719 1313 2723 1314
rect 2791 1318 2795 1319
rect 2791 1313 2795 1314
rect 2879 1318 2883 1319
rect 2886 1315 2887 1319
rect 2891 1315 2892 1319
rect 2886 1314 2892 1315
rect 3015 1318 3019 1319
rect 2879 1313 2883 1314
rect 1934 1293 1940 1294
rect 1086 1292 1092 1293
rect 970 1291 976 1292
rect 970 1287 971 1291
rect 975 1287 976 1291
rect 1086 1288 1087 1292
rect 1091 1288 1092 1292
rect 1086 1287 1092 1288
rect 1178 1291 1184 1292
rect 1178 1287 1179 1291
rect 1183 1287 1184 1291
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 1976 1290 1978 1313
rect 1934 1288 1940 1289
rect 1974 1289 1980 1290
rect 2024 1289 2026 1313
rect 2176 1289 2178 1313
rect 2368 1289 2370 1313
rect 2576 1289 2578 1313
rect 2792 1289 2794 1313
rect 970 1286 976 1287
rect 1178 1286 1184 1287
rect 972 1228 974 1286
rect 1058 1277 1064 1278
rect 1058 1273 1059 1277
rect 1063 1273 1064 1277
rect 1058 1272 1064 1273
rect 902 1227 908 1228
rect 902 1223 903 1227
rect 907 1223 908 1227
rect 902 1222 908 1223
rect 970 1227 976 1228
rect 970 1223 971 1227
rect 975 1223 976 1227
rect 970 1222 976 1223
rect 1060 1199 1062 1272
rect 579 1198 583 1199
rect 579 1193 583 1194
rect 603 1198 607 1199
rect 603 1193 607 1194
rect 763 1198 767 1199
rect 763 1193 767 1194
rect 819 1198 823 1199
rect 819 1193 823 1194
rect 923 1198 927 1199
rect 923 1193 927 1194
rect 1059 1198 1063 1199
rect 1059 1193 1063 1194
rect 1075 1198 1079 1199
rect 1075 1193 1079 1194
rect 462 1183 468 1184
rect 462 1179 463 1183
rect 467 1179 468 1183
rect 462 1178 468 1179
rect 604 1132 606 1193
rect 610 1179 616 1180
rect 610 1175 611 1179
rect 615 1175 616 1179
rect 610 1174 616 1175
rect 274 1131 280 1132
rect 274 1127 275 1131
rect 279 1127 280 1131
rect 274 1126 280 1127
rect 442 1131 448 1132
rect 442 1127 443 1131
rect 447 1127 448 1131
rect 442 1126 448 1127
rect 602 1131 608 1132
rect 602 1127 603 1131
rect 607 1127 608 1131
rect 602 1126 608 1127
rect 302 1116 308 1117
rect 470 1116 476 1117
rect 612 1116 614 1174
rect 726 1155 732 1156
rect 726 1151 727 1155
rect 731 1151 732 1155
rect 726 1150 732 1151
rect 630 1116 636 1117
rect 728 1116 730 1150
rect 764 1132 766 1193
rect 914 1183 920 1184
rect 914 1179 915 1183
rect 919 1179 920 1183
rect 914 1178 920 1179
rect 762 1131 768 1132
rect 762 1127 763 1131
rect 767 1127 768 1131
rect 762 1126 768 1127
rect 916 1124 918 1178
rect 924 1132 926 1193
rect 1076 1132 1078 1193
rect 1180 1192 1182 1286
rect 1974 1285 1975 1289
rect 1979 1285 1980 1289
rect 1974 1284 1980 1285
rect 2022 1288 2028 1289
rect 2022 1284 2023 1288
rect 2027 1284 2028 1288
rect 2022 1283 2028 1284
rect 2174 1288 2180 1289
rect 2366 1288 2372 1289
rect 2574 1288 2580 1289
rect 2790 1288 2796 1289
rect 2888 1288 2890 1314
rect 3015 1313 3019 1314
rect 3039 1318 3043 1319
rect 3039 1313 3043 1314
rect 3199 1318 3203 1319
rect 3199 1313 3203 1314
rect 3239 1318 3243 1319
rect 3239 1313 3243 1314
rect 3471 1318 3475 1319
rect 3471 1313 3475 1314
rect 3679 1318 3683 1319
rect 3679 1313 3683 1314
rect 3799 1318 3803 1319
rect 3799 1313 3803 1314
rect 3016 1289 3018 1313
rect 3240 1289 3242 1313
rect 3472 1289 3474 1313
rect 3680 1289 3682 1313
rect 3800 1290 3802 1313
rect 3840 1302 3842 1325
rect 3838 1301 3844 1302
rect 3888 1301 3890 1325
rect 3838 1297 3839 1301
rect 3843 1297 3844 1301
rect 3838 1296 3844 1297
rect 3886 1300 3892 1301
rect 3984 1300 3986 1422
rect 4084 1376 4086 1437
rect 4090 1423 4096 1424
rect 4090 1419 4091 1423
rect 4095 1419 4096 1423
rect 4090 1418 4096 1419
rect 4082 1375 4088 1376
rect 4082 1371 4083 1375
rect 4087 1371 4088 1375
rect 4082 1370 4088 1371
rect 4092 1360 4094 1418
rect 4110 1360 4116 1361
rect 4204 1360 4206 1454
rect 4316 1443 4318 1504
rect 4418 1503 4424 1504
rect 4418 1499 4419 1503
rect 4423 1499 4424 1503
rect 4418 1498 4424 1499
rect 4410 1495 4416 1496
rect 4410 1491 4411 1495
rect 4415 1491 4416 1495
rect 4410 1490 4416 1491
rect 4412 1460 4414 1490
rect 4410 1459 4416 1460
rect 4410 1455 4411 1459
rect 4415 1455 4416 1459
rect 4410 1454 4416 1455
rect 4315 1442 4319 1443
rect 4315 1437 4319 1438
rect 4323 1442 4327 1443
rect 4323 1437 4327 1438
rect 4324 1376 4326 1437
rect 4420 1428 4422 1498
rect 4548 1443 4550 1504
rect 4704 1460 4706 1518
rect 4786 1509 4792 1510
rect 4786 1505 4787 1509
rect 4791 1505 4792 1509
rect 4786 1504 4792 1505
rect 4702 1459 4708 1460
rect 4702 1455 4703 1459
rect 4707 1455 4708 1459
rect 4702 1454 4708 1455
rect 4788 1443 4790 1504
rect 4952 1460 4954 1518
rect 5034 1509 5040 1510
rect 5034 1505 5035 1509
rect 5039 1505 5040 1509
rect 5034 1504 5040 1505
rect 4950 1459 4956 1460
rect 4950 1455 4951 1459
rect 4955 1455 4956 1459
rect 4950 1454 4956 1455
rect 5036 1443 5038 1504
rect 5132 1496 5134 1582
rect 5304 1555 5306 1583
rect 5394 1582 5400 1583
rect 5303 1554 5307 1555
rect 5303 1549 5307 1550
rect 5311 1554 5315 1555
rect 5311 1549 5315 1550
rect 5312 1525 5314 1549
rect 5310 1524 5316 1525
rect 5404 1524 5406 1650
rect 5516 1604 5518 1665
rect 5636 1656 5638 1750
rect 5662 1740 5668 1741
rect 5662 1736 5663 1740
rect 5667 1736 5668 1740
rect 5662 1735 5668 1736
rect 5664 1671 5666 1735
rect 5663 1670 5667 1671
rect 5663 1665 5667 1666
rect 5634 1655 5640 1656
rect 5634 1651 5635 1655
rect 5639 1651 5640 1655
rect 5634 1650 5640 1651
rect 5664 1605 5666 1665
rect 5662 1604 5668 1605
rect 5514 1603 5520 1604
rect 5514 1599 5515 1603
rect 5519 1599 5520 1603
rect 5662 1600 5663 1604
rect 5667 1600 5668 1604
rect 5662 1599 5668 1600
rect 5514 1598 5520 1599
rect 5542 1588 5548 1589
rect 5542 1584 5543 1588
rect 5547 1584 5548 1588
rect 5542 1583 5548 1584
rect 5638 1587 5644 1588
rect 5638 1583 5639 1587
rect 5643 1583 5644 1587
rect 5544 1555 5546 1583
rect 5638 1582 5644 1583
rect 5662 1587 5668 1588
rect 5662 1583 5663 1587
rect 5667 1583 5668 1587
rect 5662 1582 5668 1583
rect 5543 1554 5547 1555
rect 5543 1549 5547 1550
rect 5544 1525 5546 1549
rect 5542 1524 5548 1525
rect 5154 1523 5160 1524
rect 5154 1519 5155 1523
rect 5159 1519 5160 1523
rect 5310 1520 5311 1524
rect 5315 1520 5316 1524
rect 5310 1519 5316 1520
rect 5402 1523 5408 1524
rect 5402 1519 5403 1523
rect 5407 1519 5408 1523
rect 5542 1520 5543 1524
rect 5547 1520 5548 1524
rect 5542 1519 5548 1520
rect 5154 1518 5160 1519
rect 5402 1518 5408 1519
rect 5156 1504 5158 1518
rect 5282 1509 5288 1510
rect 5282 1505 5283 1509
rect 5287 1505 5288 1509
rect 5282 1504 5288 1505
rect 5514 1509 5520 1510
rect 5514 1505 5515 1509
rect 5519 1505 5520 1509
rect 5514 1504 5520 1505
rect 5154 1503 5160 1504
rect 5154 1499 5155 1503
rect 5159 1499 5160 1503
rect 5154 1498 5160 1499
rect 5130 1495 5136 1496
rect 5130 1491 5131 1495
rect 5135 1491 5136 1495
rect 5130 1490 5136 1491
rect 5284 1443 5286 1504
rect 5516 1443 5518 1504
rect 5640 1460 5642 1582
rect 5664 1555 5666 1582
rect 5663 1554 5667 1555
rect 5663 1549 5667 1550
rect 5664 1526 5666 1549
rect 5662 1525 5668 1526
rect 5662 1521 5663 1525
rect 5667 1521 5668 1525
rect 5662 1520 5668 1521
rect 5662 1508 5668 1509
rect 5662 1504 5663 1508
rect 5667 1504 5668 1508
rect 5662 1503 5668 1504
rect 5638 1459 5644 1460
rect 5638 1455 5639 1459
rect 5643 1455 5644 1459
rect 5638 1454 5644 1455
rect 5542 1451 5548 1452
rect 5542 1447 5543 1451
rect 5547 1447 5548 1451
rect 5542 1446 5548 1447
rect 4547 1442 4551 1443
rect 4547 1437 4551 1438
rect 4771 1442 4775 1443
rect 4771 1437 4775 1438
rect 4787 1442 4791 1443
rect 4787 1437 4791 1438
rect 4987 1442 4991 1443
rect 4987 1437 4991 1438
rect 5035 1442 5039 1443
rect 5035 1437 5039 1438
rect 5203 1442 5207 1443
rect 5203 1437 5207 1438
rect 5283 1442 5287 1443
rect 5283 1437 5287 1438
rect 5419 1442 5423 1443
rect 5419 1437 5423 1438
rect 5515 1442 5519 1443
rect 5515 1437 5519 1438
rect 4418 1427 4424 1428
rect 4418 1423 4419 1427
rect 4423 1423 4424 1427
rect 4418 1422 4424 1423
rect 4548 1376 4550 1437
rect 4554 1423 4560 1424
rect 4554 1419 4555 1423
rect 4559 1419 4560 1423
rect 4554 1418 4560 1419
rect 4322 1375 4328 1376
rect 4322 1371 4323 1375
rect 4327 1371 4328 1375
rect 4322 1370 4328 1371
rect 4546 1375 4552 1376
rect 4546 1371 4547 1375
rect 4551 1371 4552 1375
rect 4546 1370 4552 1371
rect 4350 1360 4356 1361
rect 4556 1360 4558 1418
rect 4772 1376 4774 1437
rect 4778 1423 4784 1424
rect 4778 1419 4779 1423
rect 4783 1419 4784 1423
rect 4778 1418 4784 1419
rect 4770 1375 4776 1376
rect 4770 1371 4771 1375
rect 4775 1371 4776 1375
rect 4770 1370 4776 1371
rect 4574 1360 4580 1361
rect 4780 1360 4782 1418
rect 4988 1376 4990 1437
rect 4994 1423 5000 1424
rect 4994 1419 4995 1423
rect 4999 1419 5000 1423
rect 4994 1418 5000 1419
rect 4986 1375 4992 1376
rect 4986 1371 4987 1375
rect 4991 1371 4992 1375
rect 4986 1370 4992 1371
rect 4798 1360 4804 1361
rect 4996 1360 4998 1418
rect 5204 1376 5206 1437
rect 5210 1423 5216 1424
rect 5210 1419 5211 1423
rect 5215 1419 5216 1423
rect 5210 1418 5216 1419
rect 5202 1375 5208 1376
rect 5202 1371 5203 1375
rect 5207 1371 5208 1375
rect 5202 1370 5208 1371
rect 5014 1360 5020 1361
rect 5212 1360 5214 1418
rect 5420 1376 5422 1437
rect 5534 1427 5540 1428
rect 5534 1423 5535 1427
rect 5539 1423 5540 1427
rect 5534 1422 5540 1423
rect 5418 1375 5424 1376
rect 5418 1371 5419 1375
rect 5423 1371 5424 1375
rect 5418 1370 5424 1371
rect 5230 1360 5236 1361
rect 5446 1360 5452 1361
rect 4090 1359 4096 1360
rect 4090 1355 4091 1359
rect 4095 1355 4096 1359
rect 4110 1356 4111 1360
rect 4115 1356 4116 1360
rect 4110 1355 4116 1356
rect 4202 1359 4208 1360
rect 4202 1355 4203 1359
rect 4207 1355 4208 1359
rect 4350 1356 4351 1360
rect 4355 1356 4356 1360
rect 4350 1355 4356 1356
rect 4554 1359 4560 1360
rect 4554 1355 4555 1359
rect 4559 1355 4560 1359
rect 4574 1356 4575 1360
rect 4579 1356 4580 1360
rect 4574 1355 4580 1356
rect 4778 1359 4784 1360
rect 4778 1355 4779 1359
rect 4783 1355 4784 1359
rect 4798 1356 4799 1360
rect 4803 1356 4804 1360
rect 4798 1355 4804 1356
rect 4994 1359 5000 1360
rect 4994 1355 4995 1359
rect 4999 1355 5000 1359
rect 5014 1356 5015 1360
rect 5019 1356 5020 1360
rect 5014 1355 5020 1356
rect 5210 1359 5216 1360
rect 5210 1355 5211 1359
rect 5215 1355 5216 1359
rect 5230 1356 5231 1360
rect 5235 1356 5236 1360
rect 5230 1355 5236 1356
rect 5322 1359 5328 1360
rect 5322 1355 5323 1359
rect 5327 1355 5328 1359
rect 5446 1356 5447 1360
rect 5451 1356 5452 1360
rect 5446 1355 5452 1356
rect 4090 1354 4096 1355
rect 4112 1331 4114 1355
rect 4202 1354 4208 1355
rect 4352 1331 4354 1355
rect 4554 1354 4560 1355
rect 4576 1331 4578 1355
rect 4778 1354 4784 1355
rect 4800 1331 4802 1355
rect 4994 1354 5000 1355
rect 5016 1331 5018 1355
rect 5210 1354 5216 1355
rect 5232 1331 5234 1355
rect 5322 1354 5328 1355
rect 4111 1330 4115 1331
rect 4111 1325 4115 1326
rect 4119 1330 4123 1331
rect 4119 1325 4123 1326
rect 4351 1330 4355 1331
rect 4351 1325 4355 1326
rect 4391 1330 4395 1331
rect 4391 1325 4395 1326
rect 4575 1330 4579 1331
rect 4575 1325 4579 1326
rect 4671 1330 4675 1331
rect 4671 1325 4675 1326
rect 4799 1330 4803 1331
rect 4799 1325 4803 1326
rect 4967 1330 4971 1331
rect 4967 1325 4971 1326
rect 5015 1330 5019 1331
rect 5015 1325 5019 1326
rect 5231 1330 5235 1331
rect 5231 1325 5235 1326
rect 5263 1330 5267 1331
rect 5263 1325 5267 1326
rect 4120 1301 4122 1325
rect 4392 1301 4394 1325
rect 4672 1301 4674 1325
rect 4968 1301 4970 1325
rect 5264 1301 5266 1325
rect 4118 1300 4124 1301
rect 4390 1300 4396 1301
rect 4670 1300 4676 1301
rect 4966 1300 4972 1301
rect 5262 1300 5268 1301
rect 3886 1296 3887 1300
rect 3891 1296 3892 1300
rect 3886 1295 3892 1296
rect 3982 1299 3988 1300
rect 3982 1295 3983 1299
rect 3987 1295 3988 1299
rect 4118 1296 4119 1300
rect 4123 1296 4124 1300
rect 4118 1295 4124 1296
rect 4218 1299 4224 1300
rect 4218 1295 4219 1299
rect 4223 1295 4224 1299
rect 4390 1296 4391 1300
rect 4395 1296 4396 1300
rect 4390 1295 4396 1296
rect 4490 1299 4496 1300
rect 4490 1295 4491 1299
rect 4495 1295 4496 1299
rect 4670 1296 4671 1300
rect 4675 1296 4676 1300
rect 4670 1295 4676 1296
rect 4766 1299 4772 1300
rect 4766 1295 4767 1299
rect 4771 1295 4772 1299
rect 4966 1296 4967 1300
rect 4971 1296 4972 1300
rect 4966 1295 4972 1296
rect 5066 1299 5072 1300
rect 5066 1295 5067 1299
rect 5071 1295 5072 1299
rect 5262 1296 5263 1300
rect 5267 1296 5268 1300
rect 5262 1295 5268 1296
rect 3982 1294 3988 1295
rect 4218 1294 4224 1295
rect 4490 1294 4496 1295
rect 4766 1294 4772 1295
rect 5066 1294 5072 1295
rect 3798 1289 3804 1290
rect 3014 1288 3020 1289
rect 3238 1288 3244 1289
rect 3470 1288 3476 1289
rect 2174 1284 2175 1288
rect 2179 1284 2180 1288
rect 2174 1283 2180 1284
rect 2310 1287 2316 1288
rect 2310 1283 2311 1287
rect 2315 1283 2316 1287
rect 2366 1284 2367 1288
rect 2371 1284 2372 1288
rect 2366 1283 2372 1284
rect 2466 1287 2472 1288
rect 2466 1283 2467 1287
rect 2471 1283 2472 1287
rect 2574 1284 2575 1288
rect 2579 1284 2580 1288
rect 2574 1283 2580 1284
rect 2674 1287 2680 1288
rect 2674 1283 2675 1287
rect 2679 1283 2680 1287
rect 2790 1284 2791 1288
rect 2795 1284 2796 1288
rect 2790 1283 2796 1284
rect 2886 1287 2892 1288
rect 2886 1283 2887 1287
rect 2891 1283 2892 1287
rect 3014 1284 3015 1288
rect 3019 1284 3020 1288
rect 3014 1283 3020 1284
rect 3114 1287 3120 1288
rect 3114 1283 3115 1287
rect 3119 1283 3120 1287
rect 3238 1284 3239 1288
rect 3243 1284 3244 1288
rect 3238 1283 3244 1284
rect 3334 1287 3340 1288
rect 3334 1283 3335 1287
rect 3339 1283 3340 1287
rect 3470 1284 3471 1288
rect 3475 1284 3476 1288
rect 3470 1283 3476 1284
rect 3678 1288 3684 1289
rect 3678 1284 3679 1288
rect 3683 1284 3684 1288
rect 3678 1283 3684 1284
rect 3790 1287 3796 1288
rect 3790 1283 3791 1287
rect 3795 1283 3796 1287
rect 3798 1285 3799 1289
rect 3803 1285 3804 1289
rect 3858 1285 3864 1286
rect 3798 1284 3804 1285
rect 3838 1284 3844 1285
rect 2310 1282 2316 1283
rect 2466 1282 2472 1283
rect 2674 1282 2680 1283
rect 2886 1282 2892 1283
rect 3114 1282 3120 1283
rect 3334 1282 3340 1283
rect 3790 1282 3796 1283
rect 1934 1276 1940 1277
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 1994 1273 2000 1274
rect 1934 1271 1940 1272
rect 1974 1272 1980 1273
rect 1914 1223 1920 1224
rect 1914 1219 1915 1223
rect 1919 1219 1920 1223
rect 1914 1218 1920 1219
rect 1219 1198 1223 1199
rect 1219 1193 1223 1194
rect 1363 1198 1367 1199
rect 1363 1193 1367 1194
rect 1507 1198 1511 1199
rect 1507 1193 1511 1194
rect 1651 1198 1655 1199
rect 1651 1193 1655 1194
rect 1787 1198 1791 1199
rect 1787 1193 1791 1194
rect 1178 1191 1184 1192
rect 1178 1187 1179 1191
rect 1183 1187 1184 1191
rect 1178 1186 1184 1187
rect 1220 1132 1222 1193
rect 1334 1187 1340 1188
rect 1334 1183 1335 1187
rect 1339 1183 1340 1187
rect 1334 1182 1340 1183
rect 1226 1179 1232 1180
rect 1226 1175 1227 1179
rect 1231 1175 1232 1179
rect 1226 1174 1232 1175
rect 922 1131 928 1132
rect 922 1127 923 1131
rect 927 1127 928 1131
rect 922 1126 928 1127
rect 1074 1131 1080 1132
rect 1074 1127 1075 1131
rect 1079 1127 1080 1131
rect 1074 1126 1080 1127
rect 1218 1131 1224 1132
rect 1218 1127 1219 1131
rect 1223 1127 1224 1131
rect 1218 1126 1224 1127
rect 914 1123 920 1124
rect 914 1119 915 1123
rect 919 1119 920 1123
rect 914 1118 920 1119
rect 790 1116 796 1117
rect 950 1116 956 1117
rect 302 1112 303 1116
rect 307 1112 308 1116
rect 302 1111 308 1112
rect 398 1115 404 1116
rect 398 1111 399 1115
rect 403 1111 404 1115
rect 470 1112 471 1116
rect 475 1112 476 1116
rect 470 1111 476 1112
rect 610 1115 616 1116
rect 610 1111 611 1115
rect 615 1111 616 1115
rect 630 1112 631 1116
rect 635 1112 636 1116
rect 630 1111 636 1112
rect 726 1115 732 1116
rect 726 1111 727 1115
rect 731 1111 732 1115
rect 790 1112 791 1116
rect 795 1112 796 1116
rect 790 1111 796 1112
rect 886 1115 892 1116
rect 886 1111 887 1115
rect 891 1111 892 1115
rect 950 1112 951 1116
rect 955 1112 956 1116
rect 950 1111 956 1112
rect 1102 1116 1108 1117
rect 1228 1116 1230 1174
rect 1246 1116 1252 1117
rect 1102 1112 1103 1116
rect 1107 1112 1108 1116
rect 1102 1111 1108 1112
rect 1226 1115 1232 1116
rect 1226 1111 1227 1115
rect 1231 1111 1232 1115
rect 1246 1112 1247 1116
rect 1251 1112 1252 1116
rect 1246 1111 1252 1112
rect 304 1079 306 1111
rect 398 1110 404 1111
rect 303 1078 307 1079
rect 303 1073 307 1074
rect 174 1044 175 1048
rect 179 1044 180 1048
rect 174 1043 180 1044
rect 266 1047 272 1048
rect 266 1043 267 1047
rect 271 1043 272 1047
rect 266 1042 272 1043
rect 146 1033 152 1034
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 146 1029 147 1033
rect 151 1029 152 1033
rect 146 1028 152 1029
rect 386 1033 392 1034
rect 386 1029 387 1033
rect 391 1029 392 1033
rect 386 1028 392 1029
rect 110 1027 116 1028
rect 112 959 114 1027
rect 148 959 150 1028
rect 318 983 324 984
rect 318 979 319 983
rect 323 979 324 983
rect 318 978 324 979
rect 111 958 115 959
rect 111 953 115 954
rect 147 958 151 959
rect 147 953 151 954
rect 195 958 199 959
rect 195 953 199 954
rect 112 893 114 953
rect 110 892 116 893
rect 196 892 198 953
rect 110 888 111 892
rect 115 888 116 892
rect 110 887 116 888
rect 194 891 200 892
rect 194 887 195 891
rect 199 887 200 891
rect 194 886 200 887
rect 222 876 228 877
rect 320 876 322 978
rect 388 959 390 1028
rect 400 984 402 1110
rect 472 1079 474 1111
rect 610 1110 616 1111
rect 632 1079 634 1111
rect 726 1110 732 1111
rect 792 1079 794 1111
rect 886 1110 892 1111
rect 415 1078 419 1079
rect 415 1073 419 1074
rect 471 1078 475 1079
rect 471 1073 475 1074
rect 631 1078 635 1079
rect 631 1073 635 1074
rect 639 1078 643 1079
rect 639 1073 643 1074
rect 791 1078 795 1079
rect 791 1073 795 1074
rect 855 1078 859 1079
rect 855 1073 859 1074
rect 416 1049 418 1073
rect 640 1049 642 1073
rect 856 1049 858 1073
rect 414 1048 420 1049
rect 638 1048 644 1049
rect 854 1048 860 1049
rect 414 1044 415 1048
rect 419 1044 420 1048
rect 414 1043 420 1044
rect 514 1047 520 1048
rect 514 1043 515 1047
rect 519 1043 520 1047
rect 638 1044 639 1048
rect 643 1044 644 1048
rect 638 1043 644 1044
rect 734 1047 740 1048
rect 734 1043 735 1047
rect 739 1043 740 1047
rect 854 1044 855 1048
rect 859 1044 860 1048
rect 854 1043 860 1044
rect 514 1042 520 1043
rect 734 1042 740 1043
rect 516 984 518 1042
rect 610 1033 616 1034
rect 610 1029 611 1033
rect 615 1029 616 1033
rect 610 1028 616 1029
rect 398 983 404 984
rect 398 979 399 983
rect 403 979 404 983
rect 398 978 404 979
rect 514 983 520 984
rect 514 979 515 983
rect 519 979 520 983
rect 514 978 520 979
rect 612 959 614 1028
rect 387 958 391 959
rect 387 953 391 954
rect 419 958 423 959
rect 419 953 423 954
rect 611 958 615 959
rect 611 953 615 954
rect 667 958 671 959
rect 667 953 671 954
rect 420 892 422 953
rect 538 947 544 948
rect 538 943 539 947
rect 543 943 544 947
rect 538 942 544 943
rect 426 939 432 940
rect 426 935 427 939
rect 431 935 432 939
rect 426 934 432 935
rect 418 891 424 892
rect 418 887 419 891
rect 423 887 424 891
rect 418 886 424 887
rect 110 875 116 876
rect 110 871 111 875
rect 115 871 116 875
rect 222 872 223 876
rect 227 872 228 876
rect 222 871 228 872
rect 318 875 324 876
rect 318 871 319 875
rect 323 871 324 875
rect 110 870 116 871
rect 112 823 114 870
rect 224 823 226 871
rect 318 870 324 871
rect 111 822 115 823
rect 111 817 115 818
rect 223 822 227 823
rect 223 817 227 818
rect 112 794 114 817
rect 110 793 116 794
rect 224 793 226 817
rect 110 789 111 793
rect 115 789 116 793
rect 110 788 116 789
rect 222 792 228 793
rect 428 792 430 934
rect 446 876 452 877
rect 540 876 542 942
rect 668 892 670 953
rect 736 944 738 1042
rect 826 1033 832 1034
rect 826 1029 827 1033
rect 831 1029 832 1033
rect 826 1028 832 1029
rect 828 959 830 1028
rect 888 984 890 1110
rect 952 1079 954 1111
rect 1104 1079 1106 1111
rect 1226 1110 1232 1111
rect 1248 1079 1250 1111
rect 951 1078 955 1079
rect 951 1073 955 1074
rect 1055 1078 1059 1079
rect 1055 1073 1059 1074
rect 1103 1078 1107 1079
rect 1103 1073 1107 1074
rect 1239 1078 1243 1079
rect 1239 1073 1243 1074
rect 1247 1078 1251 1079
rect 1247 1073 1251 1074
rect 1056 1049 1058 1073
rect 1240 1049 1242 1073
rect 1054 1048 1060 1049
rect 1238 1048 1244 1049
rect 1336 1048 1338 1182
rect 1364 1132 1366 1193
rect 1370 1179 1376 1180
rect 1370 1175 1371 1179
rect 1375 1175 1376 1179
rect 1370 1174 1376 1175
rect 1362 1131 1368 1132
rect 1362 1127 1363 1131
rect 1367 1127 1368 1131
rect 1362 1126 1368 1127
rect 1372 1116 1374 1174
rect 1508 1132 1510 1193
rect 1514 1179 1520 1180
rect 1514 1175 1515 1179
rect 1519 1175 1520 1179
rect 1514 1174 1520 1175
rect 1506 1131 1512 1132
rect 1506 1127 1507 1131
rect 1511 1127 1512 1131
rect 1506 1126 1512 1127
rect 1390 1116 1396 1117
rect 1516 1116 1518 1174
rect 1652 1132 1654 1193
rect 1658 1179 1664 1180
rect 1658 1175 1659 1179
rect 1663 1175 1664 1179
rect 1658 1174 1664 1175
rect 1650 1131 1656 1132
rect 1650 1127 1651 1131
rect 1655 1127 1656 1131
rect 1650 1126 1656 1127
rect 1534 1116 1540 1117
rect 1660 1116 1662 1174
rect 1788 1132 1790 1193
rect 1794 1179 1800 1180
rect 1794 1175 1795 1179
rect 1799 1175 1800 1179
rect 1794 1174 1800 1175
rect 1786 1131 1792 1132
rect 1786 1127 1787 1131
rect 1791 1127 1792 1131
rect 1786 1126 1792 1127
rect 1678 1116 1684 1117
rect 1796 1116 1798 1174
rect 1814 1116 1820 1117
rect 1916 1116 1918 1218
rect 1936 1199 1938 1271
rect 1974 1268 1975 1272
rect 1979 1268 1980 1272
rect 1994 1269 1995 1273
rect 1999 1269 2000 1273
rect 1994 1268 2000 1269
rect 2146 1273 2152 1274
rect 2146 1269 2147 1273
rect 2151 1269 2152 1273
rect 2146 1268 2152 1269
rect 1974 1267 1980 1268
rect 1976 1199 1978 1267
rect 1996 1199 1998 1268
rect 2148 1199 2150 1268
rect 2312 1224 2314 1282
rect 2338 1273 2344 1274
rect 2338 1269 2339 1273
rect 2343 1269 2344 1273
rect 2338 1268 2344 1269
rect 2310 1223 2316 1224
rect 2310 1219 2311 1223
rect 2315 1219 2316 1223
rect 2310 1218 2316 1219
rect 2340 1199 2342 1268
rect 2468 1224 2470 1282
rect 2546 1273 2552 1274
rect 2546 1269 2547 1273
rect 2551 1269 2552 1273
rect 2546 1268 2552 1269
rect 2466 1223 2472 1224
rect 2466 1219 2467 1223
rect 2471 1219 2472 1223
rect 2466 1218 2472 1219
rect 2548 1199 2550 1268
rect 2676 1224 2678 1282
rect 2762 1273 2768 1274
rect 2762 1269 2763 1273
rect 2767 1269 2768 1273
rect 2762 1268 2768 1269
rect 2986 1273 2992 1274
rect 2986 1269 2987 1273
rect 2991 1269 2992 1273
rect 2986 1268 2992 1269
rect 2674 1223 2680 1224
rect 2674 1219 2675 1223
rect 2679 1219 2680 1223
rect 2674 1218 2680 1219
rect 2764 1199 2766 1268
rect 2988 1199 2990 1268
rect 3116 1224 3118 1282
rect 3210 1273 3216 1274
rect 3210 1269 3211 1273
rect 3215 1269 3216 1273
rect 3210 1268 3216 1269
rect 3114 1223 3120 1224
rect 3114 1219 3115 1223
rect 3119 1219 3120 1223
rect 3114 1218 3120 1219
rect 3212 1199 3214 1268
rect 1935 1198 1939 1199
rect 1935 1193 1939 1194
rect 1975 1198 1979 1199
rect 1975 1193 1979 1194
rect 1995 1198 1999 1199
rect 1995 1193 1999 1194
rect 2147 1198 2151 1199
rect 2147 1193 2151 1194
rect 2339 1198 2343 1199
rect 2339 1193 2343 1194
rect 2547 1198 2551 1199
rect 2547 1193 2551 1194
rect 2723 1198 2727 1199
rect 2723 1193 2727 1194
rect 2763 1198 2767 1199
rect 2763 1193 2767 1194
rect 2899 1198 2903 1199
rect 2899 1193 2903 1194
rect 2987 1198 2991 1199
rect 2987 1193 2991 1194
rect 3083 1198 3087 1199
rect 3083 1193 3087 1194
rect 3211 1198 3215 1199
rect 3211 1193 3215 1194
rect 3275 1198 3279 1199
rect 3275 1193 3279 1194
rect 1936 1133 1938 1193
rect 1976 1133 1978 1193
rect 1934 1132 1940 1133
rect 1934 1128 1935 1132
rect 1939 1128 1940 1132
rect 1934 1127 1940 1128
rect 1974 1132 1980 1133
rect 2724 1132 2726 1193
rect 2818 1179 2824 1180
rect 2818 1175 2819 1179
rect 2823 1175 2824 1179
rect 2818 1174 2824 1175
rect 2820 1160 2822 1174
rect 2818 1159 2824 1160
rect 2818 1155 2819 1159
rect 2823 1155 2824 1159
rect 2818 1154 2824 1155
rect 2900 1132 2902 1193
rect 2906 1179 2912 1180
rect 2906 1175 2907 1179
rect 2911 1175 2912 1179
rect 2906 1174 2912 1175
rect 1974 1128 1975 1132
rect 1979 1128 1980 1132
rect 1974 1127 1980 1128
rect 2722 1131 2728 1132
rect 2722 1127 2723 1131
rect 2727 1127 2728 1131
rect 2722 1126 2728 1127
rect 2898 1131 2904 1132
rect 2898 1127 2899 1131
rect 2903 1127 2904 1131
rect 2898 1126 2904 1127
rect 2750 1116 2756 1117
rect 2908 1116 2910 1174
rect 3084 1132 3086 1193
rect 3202 1159 3208 1160
rect 3202 1155 3203 1159
rect 3207 1155 3208 1159
rect 3202 1154 3208 1155
rect 3082 1131 3088 1132
rect 3082 1127 3083 1131
rect 3087 1127 3088 1131
rect 3082 1126 3088 1127
rect 2926 1116 2932 1117
rect 3110 1116 3116 1117
rect 3204 1116 3206 1154
rect 3276 1132 3278 1193
rect 3336 1184 3338 1282
rect 3442 1273 3448 1274
rect 3442 1269 3443 1273
rect 3447 1269 3448 1273
rect 3442 1268 3448 1269
rect 3650 1273 3656 1274
rect 3650 1269 3651 1273
rect 3655 1269 3656 1273
rect 3650 1268 3656 1269
rect 3444 1199 3446 1268
rect 3582 1223 3588 1224
rect 3582 1219 3583 1223
rect 3587 1219 3588 1223
rect 3582 1218 3588 1219
rect 3584 1203 3586 1218
rect 3584 1201 3590 1203
rect 3443 1198 3447 1199
rect 3443 1193 3447 1194
rect 3467 1198 3471 1199
rect 3467 1193 3471 1194
rect 3334 1183 3340 1184
rect 3334 1179 3335 1183
rect 3339 1179 3340 1183
rect 3334 1178 3340 1179
rect 3468 1132 3470 1193
rect 3274 1131 3280 1132
rect 3274 1127 3275 1131
rect 3279 1127 3280 1131
rect 3274 1126 3280 1127
rect 3466 1131 3472 1132
rect 3466 1127 3467 1131
rect 3471 1127 3472 1131
rect 3466 1126 3472 1127
rect 3302 1116 3308 1117
rect 1370 1115 1376 1116
rect 1370 1111 1371 1115
rect 1375 1111 1376 1115
rect 1390 1112 1391 1116
rect 1395 1112 1396 1116
rect 1390 1111 1396 1112
rect 1514 1115 1520 1116
rect 1514 1111 1515 1115
rect 1519 1111 1520 1115
rect 1534 1112 1535 1116
rect 1539 1112 1540 1116
rect 1534 1111 1540 1112
rect 1658 1115 1664 1116
rect 1658 1111 1659 1115
rect 1663 1111 1664 1115
rect 1678 1112 1679 1116
rect 1683 1112 1684 1116
rect 1678 1111 1684 1112
rect 1794 1115 1800 1116
rect 1794 1111 1795 1115
rect 1799 1111 1800 1115
rect 1814 1112 1815 1116
rect 1819 1112 1820 1116
rect 1814 1111 1820 1112
rect 1914 1115 1920 1116
rect 1914 1111 1915 1115
rect 1919 1111 1920 1115
rect 1370 1110 1376 1111
rect 1392 1079 1394 1111
rect 1514 1110 1520 1111
rect 1536 1079 1538 1111
rect 1658 1110 1664 1111
rect 1680 1079 1682 1111
rect 1794 1110 1800 1111
rect 1816 1079 1818 1111
rect 1914 1110 1920 1111
rect 1934 1115 1940 1116
rect 1934 1111 1935 1115
rect 1939 1111 1940 1115
rect 1934 1110 1940 1111
rect 1974 1115 1980 1116
rect 1974 1111 1975 1115
rect 1979 1111 1980 1115
rect 2750 1112 2751 1116
rect 2755 1112 2756 1116
rect 2750 1111 2756 1112
rect 2906 1115 2912 1116
rect 2906 1111 2907 1115
rect 2911 1111 2912 1115
rect 2926 1112 2927 1116
rect 2931 1112 2932 1116
rect 2926 1111 2932 1112
rect 3018 1115 3024 1116
rect 3018 1111 3019 1115
rect 3023 1111 3024 1115
rect 3110 1112 3111 1116
rect 3115 1112 3116 1116
rect 3110 1111 3116 1112
rect 3202 1115 3208 1116
rect 3202 1111 3203 1115
rect 3207 1111 3208 1115
rect 3302 1112 3303 1116
rect 3307 1112 3308 1116
rect 3302 1111 3308 1112
rect 3494 1116 3500 1117
rect 3588 1116 3590 1201
rect 3652 1199 3654 1268
rect 3792 1236 3794 1282
rect 3838 1280 3839 1284
rect 3843 1280 3844 1284
rect 3858 1281 3859 1285
rect 3863 1281 3864 1285
rect 3858 1280 3864 1281
rect 4090 1285 4096 1286
rect 4090 1281 4091 1285
rect 4095 1281 4096 1285
rect 4090 1280 4096 1281
rect 3838 1279 3844 1280
rect 3798 1272 3804 1273
rect 3798 1268 3799 1272
rect 3803 1268 3804 1272
rect 3798 1267 3804 1268
rect 3790 1235 3796 1236
rect 3790 1231 3791 1235
rect 3795 1231 3796 1235
rect 3790 1230 3796 1231
rect 3800 1199 3802 1267
rect 3840 1199 3842 1279
rect 3860 1199 3862 1280
rect 4092 1199 4094 1280
rect 4220 1236 4222 1294
rect 4362 1285 4368 1286
rect 4362 1281 4363 1285
rect 4367 1281 4368 1285
rect 4362 1280 4368 1281
rect 4134 1235 4140 1236
rect 4134 1231 4135 1235
rect 4139 1231 4140 1235
rect 4134 1230 4140 1231
rect 4218 1235 4224 1236
rect 4218 1231 4219 1235
rect 4223 1231 4224 1235
rect 4218 1230 4224 1231
rect 3651 1198 3655 1199
rect 3651 1193 3655 1194
rect 3799 1198 3803 1199
rect 3799 1193 3803 1194
rect 3839 1198 3843 1199
rect 3839 1193 3843 1194
rect 3859 1198 3863 1199
rect 3859 1193 3863 1194
rect 4011 1198 4015 1199
rect 4011 1193 4015 1194
rect 4091 1198 4095 1199
rect 4091 1193 4095 1194
rect 3642 1183 3648 1184
rect 3642 1179 3643 1183
rect 3647 1179 3648 1183
rect 3642 1178 3648 1179
rect 3644 1124 3646 1178
rect 3652 1132 3654 1193
rect 3670 1183 3676 1184
rect 3670 1179 3671 1183
rect 3675 1179 3676 1183
rect 3670 1178 3676 1179
rect 3650 1131 3656 1132
rect 3650 1127 3651 1131
rect 3655 1127 3656 1131
rect 3650 1126 3656 1127
rect 3642 1123 3648 1124
rect 3642 1119 3643 1123
rect 3647 1119 3648 1123
rect 3642 1118 3648 1119
rect 3494 1112 3495 1116
rect 3499 1112 3500 1116
rect 3494 1111 3500 1112
rect 3586 1115 3592 1116
rect 3586 1111 3587 1115
rect 3591 1111 3592 1115
rect 1974 1110 1980 1111
rect 1936 1079 1938 1110
rect 1391 1078 1395 1079
rect 1391 1073 1395 1074
rect 1423 1078 1427 1079
rect 1423 1073 1427 1074
rect 1535 1078 1539 1079
rect 1535 1073 1539 1074
rect 1607 1078 1611 1079
rect 1607 1073 1611 1074
rect 1679 1078 1683 1079
rect 1679 1073 1683 1074
rect 1791 1078 1795 1079
rect 1791 1073 1795 1074
rect 1815 1078 1819 1079
rect 1815 1073 1819 1074
rect 1935 1078 1939 1079
rect 1976 1075 1978 1110
rect 2752 1075 2754 1111
rect 2906 1110 2912 1111
rect 2928 1075 2930 1111
rect 3018 1110 3024 1111
rect 1935 1073 1939 1074
rect 1975 1074 1979 1075
rect 1424 1049 1426 1073
rect 1608 1049 1610 1073
rect 1792 1049 1794 1073
rect 1936 1050 1938 1073
rect 1975 1069 1979 1070
rect 2559 1074 2563 1075
rect 2559 1069 2563 1070
rect 2751 1074 2755 1075
rect 2751 1069 2755 1070
rect 2927 1074 2931 1075
rect 2927 1069 2931 1070
rect 2951 1074 2955 1075
rect 2951 1069 2955 1070
rect 1934 1049 1940 1050
rect 1422 1048 1428 1049
rect 1606 1048 1612 1049
rect 1790 1048 1796 1049
rect 954 1047 960 1048
rect 954 1043 955 1047
rect 959 1043 960 1047
rect 1054 1044 1055 1048
rect 1059 1044 1060 1048
rect 1054 1043 1060 1044
rect 1154 1047 1160 1048
rect 1154 1043 1155 1047
rect 1159 1043 1160 1047
rect 1238 1044 1239 1048
rect 1243 1044 1244 1048
rect 1238 1043 1244 1044
rect 1334 1047 1340 1048
rect 1334 1043 1335 1047
rect 1339 1043 1340 1047
rect 1422 1044 1423 1048
rect 1427 1044 1428 1048
rect 1422 1043 1428 1044
rect 1518 1047 1524 1048
rect 1518 1043 1519 1047
rect 1523 1043 1524 1047
rect 1606 1044 1607 1048
rect 1611 1044 1612 1048
rect 1606 1043 1612 1044
rect 1702 1047 1708 1048
rect 1702 1043 1703 1047
rect 1707 1043 1708 1047
rect 1790 1044 1791 1048
rect 1795 1044 1796 1048
rect 1790 1043 1796 1044
rect 1886 1047 1892 1048
rect 1886 1043 1887 1047
rect 1891 1043 1892 1047
rect 1934 1045 1935 1049
rect 1939 1045 1940 1049
rect 1976 1046 1978 1069
rect 1934 1044 1940 1045
rect 1974 1045 1980 1046
rect 2560 1045 2562 1069
rect 2752 1045 2754 1069
rect 2952 1045 2954 1069
rect 954 1042 960 1043
rect 1154 1042 1160 1043
rect 1334 1042 1340 1043
rect 1518 1042 1524 1043
rect 1702 1042 1708 1043
rect 1886 1042 1892 1043
rect 956 984 958 1042
rect 1026 1033 1032 1034
rect 1026 1029 1027 1033
rect 1031 1029 1032 1033
rect 1026 1028 1032 1029
rect 886 983 892 984
rect 886 979 887 983
rect 891 979 892 983
rect 886 978 892 979
rect 954 983 960 984
rect 954 979 955 983
rect 959 979 960 983
rect 954 978 960 979
rect 1028 959 1030 1028
rect 827 958 831 959
rect 827 953 831 954
rect 931 958 935 959
rect 931 953 935 954
rect 1027 958 1031 959
rect 1027 953 1031 954
rect 734 943 740 944
rect 734 939 735 943
rect 739 939 740 943
rect 734 938 740 939
rect 932 892 934 953
rect 1156 944 1158 1042
rect 1210 1033 1216 1034
rect 1210 1029 1211 1033
rect 1215 1029 1216 1033
rect 1210 1028 1216 1029
rect 1394 1033 1400 1034
rect 1394 1029 1395 1033
rect 1399 1029 1400 1033
rect 1394 1028 1400 1029
rect 1212 959 1214 1028
rect 1396 959 1398 1028
rect 1490 1011 1496 1012
rect 1490 1007 1491 1011
rect 1495 1007 1496 1011
rect 1490 1006 1496 1007
rect 1492 984 1494 1006
rect 1490 983 1496 984
rect 1490 979 1491 983
rect 1495 979 1496 983
rect 1490 978 1496 979
rect 1520 976 1522 1042
rect 1578 1033 1584 1034
rect 1578 1029 1579 1033
rect 1583 1029 1584 1033
rect 1578 1028 1584 1029
rect 1518 975 1524 976
rect 1518 971 1519 975
rect 1523 971 1524 975
rect 1518 970 1524 971
rect 1580 959 1582 1028
rect 1704 1012 1706 1042
rect 1762 1033 1768 1034
rect 1762 1029 1763 1033
rect 1767 1029 1768 1033
rect 1762 1028 1768 1029
rect 1702 1011 1708 1012
rect 1702 1007 1703 1011
rect 1707 1007 1708 1011
rect 1702 1006 1708 1007
rect 1764 959 1766 1028
rect 1888 976 1890 1042
rect 1974 1041 1975 1045
rect 1979 1041 1980 1045
rect 1974 1040 1980 1041
rect 2558 1044 2564 1045
rect 2750 1044 2756 1045
rect 2950 1044 2956 1045
rect 2558 1040 2559 1044
rect 2563 1040 2564 1044
rect 2558 1039 2564 1040
rect 2650 1043 2656 1044
rect 2650 1039 2651 1043
rect 2655 1039 2656 1043
rect 2750 1040 2751 1044
rect 2755 1040 2756 1044
rect 2750 1039 2756 1040
rect 2842 1043 2848 1044
rect 2842 1039 2843 1043
rect 2847 1039 2848 1043
rect 2950 1040 2951 1044
rect 2955 1040 2956 1044
rect 2950 1039 2956 1040
rect 2650 1038 2656 1039
rect 2842 1038 2848 1039
rect 1934 1032 1940 1033
rect 1934 1028 1935 1032
rect 1939 1028 1940 1032
rect 2530 1029 2536 1030
rect 1934 1027 1940 1028
rect 1974 1028 1980 1029
rect 1906 983 1912 984
rect 1906 979 1907 983
rect 1911 979 1912 983
rect 1906 978 1912 979
rect 1886 975 1892 976
rect 1886 971 1887 975
rect 1891 971 1892 975
rect 1886 970 1892 971
rect 1211 958 1215 959
rect 1211 953 1215 954
rect 1219 958 1223 959
rect 1219 953 1223 954
rect 1395 958 1399 959
rect 1395 953 1399 954
rect 1515 958 1519 959
rect 1515 953 1519 954
rect 1579 958 1583 959
rect 1579 953 1583 954
rect 1763 958 1767 959
rect 1763 953 1767 954
rect 1787 958 1791 959
rect 1787 953 1791 954
rect 1154 943 1160 944
rect 938 939 944 940
rect 938 935 939 939
rect 943 935 944 939
rect 1154 939 1155 943
rect 1159 939 1160 943
rect 1154 938 1160 939
rect 938 934 944 935
rect 666 891 672 892
rect 666 887 667 891
rect 671 887 672 891
rect 666 886 672 887
rect 930 891 936 892
rect 930 887 931 891
rect 935 887 936 891
rect 930 886 936 887
rect 694 876 700 877
rect 940 876 942 934
rect 1220 892 1222 953
rect 1516 892 1518 953
rect 1522 939 1528 940
rect 1522 935 1523 939
rect 1527 935 1528 939
rect 1522 934 1528 935
rect 1218 891 1224 892
rect 1218 887 1219 891
rect 1223 887 1224 891
rect 1218 886 1224 887
rect 1514 891 1520 892
rect 1514 887 1515 891
rect 1519 887 1520 891
rect 1514 886 1520 887
rect 958 876 964 877
rect 1246 876 1252 877
rect 1524 876 1526 934
rect 1788 892 1790 953
rect 1786 891 1792 892
rect 1786 887 1787 891
rect 1791 887 1792 891
rect 1786 886 1792 887
rect 1542 876 1548 877
rect 1814 876 1820 877
rect 1908 876 1910 978
rect 1936 959 1938 1027
rect 1974 1024 1975 1028
rect 1979 1024 1980 1028
rect 2530 1025 2531 1029
rect 2535 1025 2536 1029
rect 2530 1024 2536 1025
rect 1974 1023 1980 1024
rect 1976 963 1978 1023
rect 2532 963 2534 1024
rect 2626 1011 2632 1012
rect 2626 1007 2627 1011
rect 2631 1007 2632 1011
rect 2626 1006 2632 1007
rect 2628 980 2630 1006
rect 2626 979 2632 980
rect 2626 975 2627 979
rect 2631 975 2632 979
rect 2626 974 2632 975
rect 1975 962 1979 963
rect 1935 958 1939 959
rect 1975 957 1979 958
rect 1995 962 1999 963
rect 1995 957 1999 958
rect 2219 962 2223 963
rect 2219 957 2223 958
rect 2467 962 2471 963
rect 2467 957 2471 958
rect 2531 962 2535 963
rect 2531 957 2535 958
rect 1935 953 1939 954
rect 1936 893 1938 953
rect 1976 897 1978 957
rect 1986 943 1992 944
rect 1986 939 1987 943
rect 1991 939 1992 943
rect 1986 938 1992 939
rect 1974 896 1980 897
rect 1934 892 1940 893
rect 1934 888 1935 892
rect 1939 888 1940 892
rect 1974 892 1975 896
rect 1979 892 1980 896
rect 1974 891 1980 892
rect 1988 888 1990 938
rect 1996 896 1998 957
rect 2220 896 2222 957
rect 2342 951 2348 952
rect 2342 947 2343 951
rect 2347 947 2348 951
rect 2342 946 2348 947
rect 2314 943 2320 944
rect 2314 939 2315 943
rect 2319 939 2320 943
rect 2314 938 2320 939
rect 1994 895 2000 896
rect 1994 891 1995 895
rect 1999 891 2000 895
rect 1994 890 2000 891
rect 2218 895 2224 896
rect 2218 891 2219 895
rect 2223 891 2224 895
rect 2218 890 2224 891
rect 1934 887 1940 888
rect 1986 887 1992 888
rect 1986 883 1987 887
rect 1991 883 1992 887
rect 1986 882 1992 883
rect 2022 880 2028 881
rect 1974 879 1980 880
rect 446 872 447 876
rect 451 872 452 876
rect 446 871 452 872
rect 538 875 544 876
rect 538 871 539 875
rect 543 871 544 875
rect 694 872 695 876
rect 699 872 700 876
rect 694 871 700 872
rect 938 875 944 876
rect 938 871 939 875
rect 943 871 944 875
rect 958 872 959 876
rect 963 872 964 876
rect 958 871 964 872
rect 1054 875 1060 876
rect 1054 871 1055 875
rect 1059 871 1060 875
rect 1246 872 1247 876
rect 1251 872 1252 876
rect 1246 871 1252 872
rect 1522 875 1528 876
rect 1522 871 1523 875
rect 1527 871 1528 875
rect 1542 872 1543 876
rect 1547 872 1548 876
rect 1542 871 1548 872
rect 1638 875 1644 876
rect 1638 871 1639 875
rect 1643 871 1644 875
rect 1814 872 1815 876
rect 1819 872 1820 876
rect 1814 871 1820 872
rect 1906 875 1912 876
rect 1906 871 1907 875
rect 1911 871 1912 875
rect 448 823 450 871
rect 538 870 544 871
rect 538 859 544 860
rect 538 855 539 859
rect 543 855 544 859
rect 538 854 544 855
rect 447 822 451 823
rect 447 817 451 818
rect 448 793 450 817
rect 446 792 452 793
rect 222 788 223 792
rect 227 788 228 792
rect 222 787 228 788
rect 426 791 432 792
rect 426 787 427 791
rect 431 787 432 791
rect 446 788 447 792
rect 451 788 452 792
rect 446 787 452 788
rect 426 786 432 787
rect 194 777 200 778
rect 110 776 116 777
rect 110 772 111 776
rect 115 772 116 776
rect 194 773 195 777
rect 199 773 200 777
rect 194 772 200 773
rect 418 777 424 778
rect 418 773 419 777
rect 423 773 424 777
rect 418 772 424 773
rect 110 771 116 772
rect 112 703 114 771
rect 196 703 198 772
rect 420 703 422 772
rect 540 728 542 854
rect 696 823 698 871
rect 938 870 944 871
rect 960 823 962 871
rect 1054 870 1060 871
rect 1056 860 1058 870
rect 1054 859 1060 860
rect 1054 855 1055 859
rect 1059 855 1060 859
rect 1054 854 1060 855
rect 1248 823 1250 871
rect 1522 870 1528 871
rect 1544 823 1546 871
rect 1638 870 1644 871
rect 663 822 667 823
rect 663 817 667 818
rect 695 822 699 823
rect 695 817 699 818
rect 879 822 883 823
rect 879 817 883 818
rect 959 822 963 823
rect 959 817 963 818
rect 1087 822 1091 823
rect 1087 817 1091 818
rect 1247 822 1251 823
rect 1247 817 1251 818
rect 1295 822 1299 823
rect 1295 817 1299 818
rect 1511 822 1515 823
rect 1511 817 1515 818
rect 1543 822 1547 823
rect 1543 817 1547 818
rect 664 793 666 817
rect 880 793 882 817
rect 1088 793 1090 817
rect 1296 793 1298 817
rect 1512 793 1514 817
rect 662 792 668 793
rect 878 792 884 793
rect 1086 792 1092 793
rect 1294 792 1300 793
rect 1510 792 1516 793
rect 546 791 552 792
rect 546 787 547 791
rect 551 787 552 791
rect 662 788 663 792
rect 667 788 668 792
rect 662 787 668 788
rect 762 791 768 792
rect 762 787 763 791
rect 767 787 768 791
rect 878 788 879 792
rect 883 788 884 792
rect 878 787 884 788
rect 974 791 980 792
rect 974 787 975 791
rect 979 787 980 791
rect 1086 788 1087 792
rect 1091 788 1092 792
rect 1086 787 1092 788
rect 1178 791 1184 792
rect 1178 787 1179 791
rect 1183 787 1184 791
rect 1294 788 1295 792
rect 1299 788 1300 792
rect 1294 787 1300 788
rect 1386 791 1392 792
rect 1386 787 1387 791
rect 1391 787 1392 791
rect 1510 788 1511 792
rect 1515 788 1516 792
rect 1510 787 1516 788
rect 1606 791 1612 792
rect 1606 787 1607 791
rect 1611 787 1612 791
rect 546 786 552 787
rect 762 786 768 787
rect 974 786 980 787
rect 1178 786 1184 787
rect 1386 786 1392 787
rect 1606 786 1612 787
rect 548 728 550 786
rect 634 777 640 778
rect 634 773 635 777
rect 639 773 640 777
rect 634 772 640 773
rect 538 727 544 728
rect 538 723 539 727
rect 543 723 544 727
rect 538 722 544 723
rect 546 727 552 728
rect 546 723 547 727
rect 551 723 552 727
rect 546 722 552 723
rect 562 719 568 720
rect 562 715 563 719
rect 567 715 568 719
rect 562 714 568 715
rect 111 702 115 703
rect 111 697 115 698
rect 131 702 135 703
rect 131 697 135 698
rect 195 702 199 703
rect 195 697 199 698
rect 275 702 279 703
rect 275 697 279 698
rect 419 702 423 703
rect 419 697 423 698
rect 443 702 447 703
rect 443 697 447 698
rect 112 637 114 697
rect 110 636 116 637
rect 132 636 134 697
rect 254 687 260 688
rect 254 683 255 687
rect 259 683 260 687
rect 254 682 260 683
rect 110 632 111 636
rect 115 632 116 636
rect 110 631 116 632
rect 130 635 136 636
rect 130 631 131 635
rect 135 631 136 635
rect 130 630 136 631
rect 158 620 164 621
rect 110 619 116 620
rect 110 615 111 619
rect 115 615 116 619
rect 158 616 159 620
rect 163 616 164 620
rect 158 615 164 616
rect 110 614 116 615
rect 112 579 114 614
rect 160 579 162 615
rect 111 578 115 579
rect 111 573 115 574
rect 159 578 163 579
rect 159 573 163 574
rect 112 550 114 573
rect 110 549 116 550
rect 160 549 162 573
rect 110 545 111 549
rect 115 545 116 549
rect 110 544 116 545
rect 158 548 164 549
rect 256 548 258 682
rect 276 636 278 697
rect 282 683 288 684
rect 282 679 283 683
rect 287 679 288 683
rect 282 678 288 679
rect 274 635 280 636
rect 274 631 275 635
rect 279 631 280 635
rect 274 630 280 631
rect 284 620 286 678
rect 444 636 446 697
rect 450 683 456 684
rect 450 679 451 683
rect 455 679 456 683
rect 450 678 456 679
rect 442 635 448 636
rect 442 631 443 635
rect 447 631 448 635
rect 442 630 448 631
rect 302 620 308 621
rect 452 620 454 678
rect 470 620 476 621
rect 564 620 566 714
rect 636 703 638 772
rect 764 728 766 786
rect 850 777 856 778
rect 850 773 851 777
rect 855 773 856 777
rect 850 772 856 773
rect 762 727 768 728
rect 762 723 763 727
rect 767 723 768 727
rect 762 722 768 723
rect 852 703 854 772
rect 611 702 615 703
rect 611 697 615 698
rect 635 702 639 703
rect 635 697 639 698
rect 771 702 775 703
rect 771 697 775 698
rect 851 702 855 703
rect 851 697 855 698
rect 923 702 927 703
rect 923 697 927 698
rect 612 636 614 697
rect 762 687 768 688
rect 762 683 763 687
rect 767 683 768 687
rect 762 682 768 683
rect 610 635 616 636
rect 610 631 611 635
rect 615 631 616 635
rect 610 630 616 631
rect 764 628 766 682
rect 772 636 774 697
rect 910 687 916 688
rect 910 683 911 687
rect 915 683 916 687
rect 910 682 916 683
rect 770 635 776 636
rect 770 631 771 635
rect 775 631 776 635
rect 770 630 776 631
rect 912 628 914 682
rect 924 636 926 697
rect 976 688 978 786
rect 1058 777 1064 778
rect 1058 773 1059 777
rect 1063 773 1064 777
rect 1058 772 1064 773
rect 1060 703 1062 772
rect 1059 702 1063 703
rect 1059 697 1063 698
rect 1075 702 1079 703
rect 1075 697 1079 698
rect 974 687 980 688
rect 974 683 975 687
rect 979 683 980 687
rect 974 682 980 683
rect 1076 636 1078 697
rect 1180 688 1182 786
rect 1266 777 1272 778
rect 1266 773 1267 777
rect 1271 773 1272 777
rect 1266 772 1272 773
rect 1268 703 1270 772
rect 1388 720 1390 786
rect 1482 777 1488 778
rect 1482 773 1483 777
rect 1487 773 1488 777
rect 1482 772 1488 773
rect 1386 719 1392 720
rect 1386 715 1387 719
rect 1391 715 1392 719
rect 1386 714 1392 715
rect 1484 703 1486 772
rect 1608 720 1610 786
rect 1640 728 1642 870
rect 1816 823 1818 871
rect 1906 870 1912 871
rect 1934 875 1940 876
rect 1934 871 1935 875
rect 1939 871 1940 875
rect 1974 875 1975 879
rect 1979 875 1980 879
rect 2022 876 2023 880
rect 2027 876 2028 880
rect 2022 875 2028 876
rect 2246 880 2252 881
rect 2246 876 2247 880
rect 2251 876 2252 880
rect 2246 875 2252 876
rect 1974 874 1980 875
rect 1934 870 1940 871
rect 1936 823 1938 870
rect 1976 851 1978 874
rect 2024 851 2026 875
rect 2248 851 2250 875
rect 1975 850 1979 851
rect 1975 845 1979 846
rect 2023 850 2027 851
rect 2023 845 2027 846
rect 2223 850 2227 851
rect 2223 845 2227 846
rect 2247 850 2251 851
rect 2247 845 2251 846
rect 1815 822 1819 823
rect 1815 817 1819 818
rect 1935 822 1939 823
rect 1976 822 1978 845
rect 1935 817 1939 818
rect 1974 821 1980 822
rect 2224 821 2226 845
rect 1974 817 1975 821
rect 1979 817 1980 821
rect 1936 794 1938 817
rect 1974 816 1980 817
rect 2222 820 2228 821
rect 2316 820 2318 938
rect 2344 880 2346 946
rect 2468 896 2470 957
rect 2652 948 2654 1038
rect 2722 1029 2728 1030
rect 2722 1025 2723 1029
rect 2727 1025 2728 1029
rect 2722 1024 2728 1025
rect 2724 963 2726 1024
rect 2844 1012 2846 1038
rect 2922 1029 2928 1030
rect 2922 1025 2923 1029
rect 2927 1025 2928 1029
rect 2922 1024 2928 1025
rect 2842 1011 2848 1012
rect 2842 1007 2843 1011
rect 2847 1007 2848 1011
rect 2842 1006 2848 1007
rect 2924 963 2926 1024
rect 3020 980 3022 1110
rect 3112 1075 3114 1111
rect 3202 1110 3208 1111
rect 3304 1075 3306 1111
rect 3496 1075 3498 1111
rect 3586 1110 3592 1111
rect 3111 1074 3115 1075
rect 3111 1069 3115 1070
rect 3151 1074 3155 1075
rect 3151 1069 3155 1070
rect 3303 1074 3307 1075
rect 3303 1069 3307 1070
rect 3359 1074 3363 1075
rect 3359 1069 3363 1070
rect 3495 1074 3499 1075
rect 3495 1069 3499 1070
rect 3575 1074 3579 1075
rect 3575 1069 3579 1070
rect 3152 1045 3154 1069
rect 3360 1045 3362 1069
rect 3576 1045 3578 1069
rect 3150 1044 3156 1045
rect 3358 1044 3364 1045
rect 3574 1044 3580 1045
rect 3672 1044 3674 1178
rect 3800 1133 3802 1193
rect 3840 1133 3842 1193
rect 3798 1132 3804 1133
rect 3798 1128 3799 1132
rect 3803 1128 3804 1132
rect 3798 1127 3804 1128
rect 3838 1132 3844 1133
rect 4012 1132 4014 1193
rect 3838 1128 3839 1132
rect 3843 1128 3844 1132
rect 3838 1127 3844 1128
rect 4010 1131 4016 1132
rect 4010 1127 4011 1131
rect 4015 1127 4016 1131
rect 4010 1126 4016 1127
rect 3678 1116 3684 1117
rect 4038 1116 4044 1117
rect 4136 1116 4138 1230
rect 4364 1199 4366 1280
rect 4492 1236 4494 1294
rect 4642 1285 4648 1286
rect 4642 1281 4643 1285
rect 4647 1281 4648 1285
rect 4642 1280 4648 1281
rect 4490 1235 4496 1236
rect 4490 1231 4491 1235
rect 4495 1231 4496 1235
rect 4490 1230 4496 1231
rect 4644 1199 4646 1280
rect 4211 1198 4215 1199
rect 4211 1193 4215 1194
rect 4363 1198 4367 1199
rect 4363 1193 4367 1194
rect 4435 1198 4439 1199
rect 4435 1193 4439 1194
rect 4643 1198 4647 1199
rect 4643 1193 4647 1194
rect 4691 1198 4695 1199
rect 4691 1193 4695 1194
rect 4212 1132 4214 1193
rect 4334 1187 4340 1188
rect 4334 1183 4335 1187
rect 4339 1183 4340 1187
rect 4334 1182 4340 1183
rect 4218 1179 4224 1180
rect 4218 1175 4219 1179
rect 4223 1175 4224 1179
rect 4218 1174 4224 1175
rect 4210 1131 4216 1132
rect 4210 1127 4211 1131
rect 4215 1127 4216 1131
rect 4210 1126 4216 1127
rect 3678 1112 3679 1116
rect 3683 1112 3684 1116
rect 3678 1111 3684 1112
rect 3798 1115 3804 1116
rect 3798 1111 3799 1115
rect 3803 1111 3804 1115
rect 3680 1075 3682 1111
rect 3798 1110 3804 1111
rect 3838 1115 3844 1116
rect 3838 1111 3839 1115
rect 3843 1111 3844 1115
rect 4038 1112 4039 1116
rect 4043 1112 4044 1116
rect 4038 1111 4044 1112
rect 4134 1115 4140 1116
rect 4134 1111 4135 1115
rect 4139 1111 4140 1115
rect 3838 1110 3844 1111
rect 3800 1075 3802 1110
rect 3840 1075 3842 1110
rect 4040 1075 4042 1111
rect 4134 1110 4140 1111
rect 3679 1074 3683 1075
rect 3679 1069 3683 1070
rect 3799 1074 3803 1075
rect 3799 1069 3803 1070
rect 3839 1074 3843 1075
rect 3839 1069 3843 1070
rect 4039 1074 4043 1075
rect 4039 1069 4043 1070
rect 4095 1074 4099 1075
rect 4095 1069 4099 1070
rect 3800 1046 3802 1069
rect 3840 1046 3842 1069
rect 3798 1045 3804 1046
rect 3050 1043 3056 1044
rect 3050 1039 3051 1043
rect 3055 1039 3056 1043
rect 3150 1040 3151 1044
rect 3155 1040 3156 1044
rect 3150 1039 3156 1040
rect 3242 1043 3248 1044
rect 3242 1039 3243 1043
rect 3247 1039 3248 1043
rect 3358 1040 3359 1044
rect 3363 1040 3364 1044
rect 3358 1039 3364 1040
rect 3458 1043 3464 1044
rect 3458 1039 3459 1043
rect 3463 1039 3464 1043
rect 3574 1040 3575 1044
rect 3579 1040 3580 1044
rect 3574 1039 3580 1040
rect 3670 1043 3676 1044
rect 3670 1039 3671 1043
rect 3675 1039 3676 1043
rect 3798 1041 3799 1045
rect 3803 1041 3804 1045
rect 3798 1040 3804 1041
rect 3838 1045 3844 1046
rect 4096 1045 4098 1069
rect 3838 1041 3839 1045
rect 3843 1041 3844 1045
rect 3838 1040 3844 1041
rect 4094 1044 4100 1045
rect 4220 1044 4222 1174
rect 4238 1116 4244 1117
rect 4336 1116 4338 1182
rect 4436 1132 4438 1193
rect 4682 1183 4688 1184
rect 4682 1179 4683 1183
rect 4687 1179 4688 1183
rect 4682 1178 4688 1179
rect 4434 1131 4440 1132
rect 4434 1127 4435 1131
rect 4439 1127 4440 1131
rect 4434 1126 4440 1127
rect 4684 1124 4686 1178
rect 4692 1132 4694 1193
rect 4768 1184 4770 1294
rect 4938 1285 4944 1286
rect 4938 1281 4939 1285
rect 4943 1281 4944 1285
rect 4938 1280 4944 1281
rect 4940 1199 4942 1280
rect 5068 1236 5070 1294
rect 5234 1285 5240 1286
rect 5234 1281 5235 1285
rect 5239 1281 5240 1285
rect 5234 1280 5240 1281
rect 5066 1235 5072 1236
rect 5066 1231 5067 1235
rect 5071 1231 5072 1235
rect 5066 1230 5072 1231
rect 5236 1199 5238 1280
rect 5324 1228 5326 1354
rect 5448 1331 5450 1355
rect 5447 1330 5451 1331
rect 5447 1325 5451 1326
rect 5354 1299 5360 1300
rect 5354 1295 5355 1299
rect 5359 1295 5360 1299
rect 5354 1294 5360 1295
rect 5322 1227 5328 1228
rect 5322 1223 5323 1227
rect 5327 1223 5328 1227
rect 5322 1222 5328 1223
rect 4939 1198 4943 1199
rect 4939 1193 4943 1194
rect 4963 1198 4967 1199
rect 4963 1193 4967 1194
rect 5235 1198 5239 1199
rect 5235 1193 5239 1194
rect 5251 1198 5255 1199
rect 5251 1193 5255 1194
rect 4766 1183 4772 1184
rect 4766 1179 4767 1183
rect 4771 1179 4772 1183
rect 4766 1178 4772 1179
rect 4964 1132 4966 1193
rect 4970 1179 4976 1180
rect 4970 1175 4971 1179
rect 4975 1175 4976 1179
rect 4970 1174 4976 1175
rect 4690 1131 4696 1132
rect 4690 1127 4691 1131
rect 4695 1127 4696 1131
rect 4690 1126 4696 1127
rect 4962 1131 4968 1132
rect 4962 1127 4963 1131
rect 4967 1127 4968 1131
rect 4962 1126 4968 1127
rect 4682 1123 4688 1124
rect 4682 1119 4683 1123
rect 4687 1119 4688 1123
rect 4682 1118 4688 1119
rect 4462 1116 4468 1117
rect 4718 1116 4724 1117
rect 4972 1116 4974 1174
rect 5252 1132 5254 1193
rect 5356 1184 5358 1294
rect 5514 1285 5520 1286
rect 5514 1281 5515 1285
rect 5519 1281 5520 1285
rect 5514 1280 5520 1281
rect 5516 1199 5518 1280
rect 5515 1198 5519 1199
rect 5515 1193 5519 1194
rect 5354 1183 5360 1184
rect 5354 1179 5355 1183
rect 5359 1179 5360 1183
rect 5354 1178 5360 1179
rect 5516 1132 5518 1193
rect 5250 1131 5256 1132
rect 5250 1127 5251 1131
rect 5255 1127 5256 1131
rect 5250 1126 5256 1127
rect 5514 1131 5520 1132
rect 5514 1127 5515 1131
rect 5519 1127 5520 1131
rect 5514 1126 5520 1127
rect 4990 1116 4996 1117
rect 4238 1112 4239 1116
rect 4243 1112 4244 1116
rect 4238 1111 4244 1112
rect 4334 1115 4340 1116
rect 4334 1111 4335 1115
rect 4339 1111 4340 1115
rect 4462 1112 4463 1116
rect 4467 1112 4468 1116
rect 4462 1111 4468 1112
rect 4578 1115 4584 1116
rect 4578 1111 4579 1115
rect 4583 1111 4584 1115
rect 4718 1112 4719 1116
rect 4723 1112 4724 1116
rect 4718 1111 4724 1112
rect 4970 1115 4976 1116
rect 4970 1111 4971 1115
rect 4975 1111 4976 1115
rect 4990 1112 4991 1116
rect 4995 1112 4996 1116
rect 4990 1111 4996 1112
rect 5278 1116 5284 1117
rect 5278 1112 5279 1116
rect 5283 1112 5284 1116
rect 5278 1111 5284 1112
rect 5374 1115 5380 1116
rect 5374 1111 5375 1115
rect 5379 1111 5380 1115
rect 4240 1075 4242 1111
rect 4334 1110 4340 1111
rect 4464 1075 4466 1111
rect 4578 1110 4584 1111
rect 4239 1074 4243 1075
rect 4239 1069 4243 1070
rect 4391 1074 4395 1075
rect 4391 1069 4395 1070
rect 4463 1074 4467 1075
rect 4463 1069 4467 1070
rect 4392 1045 4394 1069
rect 4390 1044 4396 1045
rect 4094 1040 4095 1044
rect 4099 1040 4100 1044
rect 4094 1039 4100 1040
rect 4218 1043 4224 1044
rect 4218 1039 4219 1043
rect 4223 1039 4224 1043
rect 4390 1040 4391 1044
rect 4395 1040 4396 1044
rect 4390 1039 4396 1040
rect 4482 1043 4488 1044
rect 4482 1039 4483 1043
rect 4487 1039 4488 1043
rect 3050 1038 3056 1039
rect 3242 1038 3248 1039
rect 3458 1038 3464 1039
rect 3670 1038 3676 1039
rect 4218 1038 4224 1039
rect 4482 1038 4488 1039
rect 3052 980 3054 1038
rect 3122 1029 3128 1030
rect 3122 1025 3123 1029
rect 3127 1025 3128 1029
rect 3122 1024 3128 1025
rect 3018 979 3024 980
rect 3018 975 3019 979
rect 3023 975 3024 979
rect 3018 974 3024 975
rect 3050 979 3056 980
rect 3050 975 3051 979
rect 3055 975 3056 979
rect 3050 974 3056 975
rect 3124 963 3126 1024
rect 3244 972 3246 1038
rect 3330 1029 3336 1030
rect 3330 1025 3331 1029
rect 3335 1025 3336 1029
rect 3330 1024 3336 1025
rect 3242 971 3248 972
rect 3242 967 3243 971
rect 3247 967 3248 971
rect 3242 966 3248 967
rect 3332 963 3334 1024
rect 3460 980 3462 1038
rect 3546 1029 3552 1030
rect 4066 1029 4072 1030
rect 3546 1025 3547 1029
rect 3551 1025 3552 1029
rect 3546 1024 3552 1025
rect 3798 1028 3804 1029
rect 3798 1024 3799 1028
rect 3803 1024 3804 1028
rect 3458 979 3464 980
rect 3458 975 3459 979
rect 3463 975 3464 979
rect 3458 974 3464 975
rect 3530 971 3536 972
rect 3530 967 3531 971
rect 3535 967 3536 971
rect 3530 966 3536 967
rect 2707 962 2711 963
rect 2707 957 2711 958
rect 2723 962 2727 963
rect 2723 957 2727 958
rect 2923 962 2927 963
rect 2923 957 2927 958
rect 2939 962 2943 963
rect 2939 957 2943 958
rect 3123 962 3127 963
rect 3123 957 3127 958
rect 3171 962 3175 963
rect 3171 957 3175 958
rect 3331 962 3335 963
rect 3331 957 3335 958
rect 3411 962 3415 963
rect 3411 957 3415 958
rect 2650 947 2656 948
rect 2650 943 2651 947
rect 2655 943 2656 947
rect 2650 942 2656 943
rect 2708 896 2710 957
rect 2714 943 2720 944
rect 2714 939 2715 943
rect 2719 939 2720 943
rect 2714 938 2720 939
rect 2466 895 2472 896
rect 2466 891 2467 895
rect 2471 891 2472 895
rect 2466 890 2472 891
rect 2706 895 2712 896
rect 2706 891 2707 895
rect 2711 891 2712 895
rect 2706 890 2712 891
rect 2494 880 2500 881
rect 2716 880 2718 938
rect 2940 896 2942 957
rect 3034 943 3040 944
rect 3034 939 3035 943
rect 3039 939 3040 943
rect 3034 938 3040 939
rect 3036 904 3038 938
rect 3034 903 3040 904
rect 3034 899 3035 903
rect 3039 899 3040 903
rect 3034 898 3040 899
rect 3172 896 3174 957
rect 3178 943 3184 944
rect 3178 939 3179 943
rect 3183 939 3184 943
rect 3178 938 3184 939
rect 2938 895 2944 896
rect 2938 891 2939 895
rect 2943 891 2944 895
rect 2938 890 2944 891
rect 3170 895 3176 896
rect 3170 891 3171 895
rect 3175 891 3176 895
rect 3170 890 3176 891
rect 2734 880 2740 881
rect 2966 880 2972 881
rect 3180 880 3182 938
rect 3206 903 3212 904
rect 3206 899 3207 903
rect 3211 899 3212 903
rect 3206 898 3212 899
rect 3198 880 3204 881
rect 2342 879 2348 880
rect 2342 875 2343 879
rect 2347 875 2348 879
rect 2494 876 2495 880
rect 2499 876 2500 880
rect 2494 875 2500 876
rect 2714 879 2720 880
rect 2714 875 2715 879
rect 2719 875 2720 879
rect 2734 876 2735 880
rect 2739 876 2740 880
rect 2734 875 2740 876
rect 2830 879 2836 880
rect 2830 875 2831 879
rect 2835 875 2836 879
rect 2966 876 2967 880
rect 2971 876 2972 880
rect 2966 875 2972 876
rect 3178 879 3184 880
rect 3178 875 3179 879
rect 3183 875 3184 879
rect 3198 876 3199 880
rect 3203 876 3204 880
rect 3198 875 3204 876
rect 2342 874 2348 875
rect 2496 851 2498 875
rect 2714 874 2720 875
rect 2736 851 2738 875
rect 2830 874 2836 875
rect 2439 850 2443 851
rect 2439 845 2443 846
rect 2495 850 2499 851
rect 2495 845 2499 846
rect 2663 850 2667 851
rect 2663 845 2667 846
rect 2735 850 2739 851
rect 2735 845 2739 846
rect 2440 821 2442 845
rect 2664 821 2666 845
rect 2438 820 2444 821
rect 2662 820 2668 821
rect 2222 816 2223 820
rect 2227 816 2228 820
rect 2222 815 2228 816
rect 2314 819 2320 820
rect 2314 815 2315 819
rect 2319 815 2320 819
rect 2438 816 2439 820
rect 2443 816 2444 820
rect 2438 815 2444 816
rect 2534 819 2540 820
rect 2534 815 2535 819
rect 2539 815 2540 819
rect 2662 816 2663 820
rect 2667 816 2668 820
rect 2662 815 2668 816
rect 2758 819 2764 820
rect 2758 815 2759 819
rect 2763 815 2764 819
rect 2314 814 2320 815
rect 2534 814 2540 815
rect 2758 814 2764 815
rect 2194 805 2200 806
rect 1974 804 1980 805
rect 1974 800 1975 804
rect 1979 800 1980 804
rect 2194 801 2195 805
rect 2199 801 2200 805
rect 2194 800 2200 801
rect 2410 805 2416 806
rect 2410 801 2411 805
rect 2415 801 2416 805
rect 2410 800 2416 801
rect 1974 799 1980 800
rect 1934 793 1940 794
rect 1934 789 1935 793
rect 1939 789 1940 793
rect 1934 788 1940 789
rect 1934 776 1940 777
rect 1934 772 1935 776
rect 1939 772 1940 776
rect 1934 771 1940 772
rect 1638 727 1644 728
rect 1638 723 1639 727
rect 1643 723 1644 727
rect 1638 722 1644 723
rect 1606 719 1612 720
rect 1606 715 1607 719
rect 1611 715 1612 719
rect 1606 714 1612 715
rect 1936 703 1938 771
rect 1976 723 1978 799
rect 2196 723 2198 800
rect 2412 723 2414 800
rect 2536 748 2538 814
rect 2634 805 2640 806
rect 2634 801 2635 805
rect 2639 801 2640 805
rect 2634 800 2640 801
rect 2534 747 2540 748
rect 2534 743 2535 747
rect 2539 743 2540 747
rect 2534 742 2540 743
rect 2636 723 2638 800
rect 2760 748 2762 814
rect 2832 756 2834 874
rect 2968 851 2970 875
rect 3178 874 3184 875
rect 3200 851 3202 875
rect 2887 850 2891 851
rect 2887 845 2891 846
rect 2967 850 2971 851
rect 2967 845 2971 846
rect 3111 850 3115 851
rect 3111 845 3115 846
rect 3199 850 3203 851
rect 3199 845 3203 846
rect 2888 821 2890 845
rect 3112 821 3114 845
rect 2886 820 2892 821
rect 3110 820 3116 821
rect 3208 820 3210 898
rect 3412 896 3414 957
rect 3418 943 3424 944
rect 3418 939 3419 943
rect 3423 939 3424 943
rect 3418 938 3424 939
rect 3410 895 3416 896
rect 3410 891 3411 895
rect 3415 891 3416 895
rect 3410 890 3416 891
rect 3420 880 3422 938
rect 3438 880 3444 881
rect 3532 880 3534 966
rect 3548 963 3550 1024
rect 3798 1023 3804 1024
rect 3838 1028 3844 1029
rect 3838 1024 3839 1028
rect 3843 1024 3844 1028
rect 4066 1025 4067 1029
rect 4071 1025 4072 1029
rect 4066 1024 4072 1025
rect 4362 1029 4368 1030
rect 4362 1025 4363 1029
rect 4367 1025 4368 1029
rect 4362 1024 4368 1025
rect 3838 1023 3844 1024
rect 3800 963 3802 1023
rect 3547 962 3551 963
rect 3547 957 3551 958
rect 3799 962 3803 963
rect 3840 959 3842 1023
rect 4068 959 4070 1024
rect 4274 979 4280 980
rect 4274 975 4275 979
rect 4279 975 4280 979
rect 4274 974 4280 975
rect 3799 957 3803 958
rect 3839 958 3843 959
rect 3800 897 3802 957
rect 3839 953 3843 954
rect 3931 958 3935 959
rect 3931 953 3935 954
rect 4067 958 4071 959
rect 4067 953 4071 954
rect 4155 958 4159 959
rect 4155 953 4159 954
rect 3798 896 3804 897
rect 3798 892 3799 896
rect 3803 892 3804 896
rect 3840 893 3842 953
rect 3798 891 3804 892
rect 3838 892 3844 893
rect 3932 892 3934 953
rect 3982 943 3988 944
rect 3982 939 3983 943
rect 3987 939 3988 943
rect 3982 938 3988 939
rect 3838 888 3839 892
rect 3843 888 3844 892
rect 3838 887 3844 888
rect 3930 891 3936 892
rect 3930 887 3931 891
rect 3935 887 3936 891
rect 3930 886 3936 887
rect 3418 879 3424 880
rect 3418 875 3419 879
rect 3423 875 3424 879
rect 3438 876 3439 880
rect 3443 876 3444 880
rect 3438 875 3444 876
rect 3530 879 3536 880
rect 3530 875 3531 879
rect 3535 875 3536 879
rect 3418 874 3424 875
rect 3440 851 3442 875
rect 3530 874 3536 875
rect 3798 879 3804 880
rect 3798 875 3799 879
rect 3803 875 3804 879
rect 3958 876 3964 877
rect 3798 874 3804 875
rect 3838 875 3844 876
rect 3800 851 3802 874
rect 3838 871 3839 875
rect 3843 871 3844 875
rect 3958 872 3959 876
rect 3963 872 3964 876
rect 3958 871 3964 872
rect 3838 870 3844 871
rect 3335 850 3339 851
rect 3335 845 3339 846
rect 3439 850 3443 851
rect 3439 845 3443 846
rect 3559 850 3563 851
rect 3559 845 3563 846
rect 3799 850 3803 851
rect 3840 847 3842 870
rect 3960 847 3962 871
rect 3799 845 3803 846
rect 3839 846 3843 847
rect 3336 821 3338 845
rect 3560 821 3562 845
rect 3800 822 3802 845
rect 3839 841 3843 842
rect 3887 846 3891 847
rect 3887 841 3891 842
rect 3959 846 3963 847
rect 3959 841 3963 842
rect 3798 821 3804 822
rect 3334 820 3340 821
rect 3558 820 3564 821
rect 2886 816 2887 820
rect 2891 816 2892 820
rect 2886 815 2892 816
rect 2978 819 2984 820
rect 2978 815 2979 819
rect 2983 815 2984 819
rect 3110 816 3111 820
rect 3115 816 3116 820
rect 3110 815 3116 816
rect 3206 819 3212 820
rect 3206 815 3207 819
rect 3211 815 3212 819
rect 3334 816 3335 820
rect 3339 816 3340 820
rect 3334 815 3340 816
rect 3430 819 3436 820
rect 3430 815 3431 819
rect 3435 815 3436 819
rect 3558 816 3559 820
rect 3563 816 3564 820
rect 3558 815 3564 816
rect 3650 819 3656 820
rect 3650 815 3651 819
rect 3655 815 3656 819
rect 3798 817 3799 821
rect 3803 817 3804 821
rect 3840 818 3842 841
rect 3798 816 3804 817
rect 3838 817 3844 818
rect 3888 817 3890 841
rect 2978 814 2984 815
rect 3206 814 3212 815
rect 3430 814 3436 815
rect 3650 814 3656 815
rect 2858 805 2864 806
rect 2858 801 2859 805
rect 2863 801 2864 805
rect 2858 800 2864 801
rect 2830 755 2836 756
rect 2830 751 2831 755
rect 2835 751 2836 755
rect 2830 750 2836 751
rect 2758 747 2764 748
rect 2758 743 2759 747
rect 2763 743 2764 747
rect 2758 742 2764 743
rect 2860 723 2862 800
rect 2980 748 2982 814
rect 3082 805 3088 806
rect 3082 801 3083 805
rect 3087 801 3088 805
rect 3082 800 3088 801
rect 3306 805 3312 806
rect 3306 801 3307 805
rect 3311 801 3312 805
rect 3306 800 3312 801
rect 2978 747 2984 748
rect 2978 743 2979 747
rect 2983 743 2984 747
rect 2978 742 2984 743
rect 3084 723 3086 800
rect 3178 783 3184 784
rect 3178 779 3179 783
rect 3183 779 3184 783
rect 3178 778 3184 779
rect 3180 756 3182 778
rect 3178 755 3184 756
rect 3178 751 3179 755
rect 3183 751 3184 755
rect 3178 750 3184 751
rect 3308 723 3310 800
rect 3432 784 3434 814
rect 3530 805 3536 806
rect 3530 801 3531 805
rect 3535 801 3536 805
rect 3530 800 3536 801
rect 3430 783 3436 784
rect 3430 779 3431 783
rect 3435 779 3436 783
rect 3430 778 3436 779
rect 3506 755 3512 756
rect 3506 751 3507 755
rect 3511 751 3512 755
rect 3506 750 3512 751
rect 1975 722 1979 723
rect 1975 717 1979 718
rect 2195 722 2199 723
rect 2195 717 2199 718
rect 2411 722 2415 723
rect 2411 717 2415 718
rect 2635 722 2639 723
rect 2635 717 2639 718
rect 2859 722 2863 723
rect 2859 717 2863 718
rect 3083 722 3087 723
rect 3083 717 3087 718
rect 3307 722 3311 723
rect 3307 717 3311 718
rect 3379 722 3383 723
rect 3379 717 3383 718
rect 1219 702 1223 703
rect 1219 697 1223 698
rect 1267 702 1271 703
rect 1267 697 1271 698
rect 1363 702 1367 703
rect 1363 697 1367 698
rect 1483 702 1487 703
rect 1483 697 1487 698
rect 1507 702 1511 703
rect 1507 697 1511 698
rect 1651 702 1655 703
rect 1651 697 1655 698
rect 1787 702 1791 703
rect 1787 697 1791 698
rect 1935 702 1939 703
rect 1935 697 1939 698
rect 1178 687 1184 688
rect 1178 683 1179 687
rect 1183 683 1184 687
rect 1178 682 1184 683
rect 1220 636 1222 697
rect 1226 683 1232 684
rect 1226 679 1227 683
rect 1231 679 1232 683
rect 1226 678 1232 679
rect 922 635 928 636
rect 922 631 923 635
rect 927 631 928 635
rect 922 630 928 631
rect 1074 635 1080 636
rect 1074 631 1075 635
rect 1079 631 1080 635
rect 1074 630 1080 631
rect 1218 635 1224 636
rect 1218 631 1219 635
rect 1223 631 1224 635
rect 1218 630 1224 631
rect 762 627 768 628
rect 762 623 763 627
rect 767 623 768 627
rect 762 622 768 623
rect 910 627 916 628
rect 910 623 911 627
rect 915 623 916 627
rect 910 622 916 623
rect 638 620 644 621
rect 798 620 804 621
rect 282 619 288 620
rect 282 615 283 619
rect 287 615 288 619
rect 302 616 303 620
rect 307 616 308 620
rect 302 615 308 616
rect 450 619 456 620
rect 450 615 451 619
rect 455 615 456 619
rect 470 616 471 620
rect 475 616 476 620
rect 470 615 476 616
rect 562 619 568 620
rect 562 615 563 619
rect 567 615 568 619
rect 638 616 639 620
rect 643 616 644 620
rect 638 615 644 616
rect 734 619 740 620
rect 734 615 735 619
rect 739 615 740 619
rect 798 616 799 620
rect 803 616 804 620
rect 798 615 804 616
rect 950 620 956 621
rect 950 616 951 620
rect 955 616 956 620
rect 950 615 956 616
rect 1102 620 1108 621
rect 1228 620 1230 678
rect 1364 636 1366 697
rect 1370 683 1376 684
rect 1370 679 1371 683
rect 1375 679 1376 683
rect 1370 678 1376 679
rect 1362 635 1368 636
rect 1362 631 1363 635
rect 1367 631 1368 635
rect 1362 630 1368 631
rect 1246 620 1252 621
rect 1372 620 1374 678
rect 1508 636 1510 697
rect 1514 683 1520 684
rect 1514 679 1515 683
rect 1519 679 1520 683
rect 1514 678 1520 679
rect 1506 635 1512 636
rect 1506 631 1507 635
rect 1511 631 1512 635
rect 1506 630 1512 631
rect 1390 620 1396 621
rect 1516 620 1518 678
rect 1652 636 1654 697
rect 1658 683 1664 684
rect 1658 679 1659 683
rect 1663 679 1664 683
rect 1658 678 1664 679
rect 1650 635 1656 636
rect 1650 631 1651 635
rect 1655 631 1656 635
rect 1650 630 1656 631
rect 1534 620 1540 621
rect 1660 620 1662 678
rect 1788 636 1790 697
rect 1794 683 1800 684
rect 1794 679 1795 683
rect 1799 679 1800 683
rect 1794 678 1800 679
rect 1786 635 1792 636
rect 1786 631 1787 635
rect 1791 631 1792 635
rect 1786 630 1792 631
rect 1678 620 1684 621
rect 1796 620 1798 678
rect 1936 637 1938 697
rect 1976 657 1978 717
rect 1974 656 1980 657
rect 3380 656 3382 717
rect 3474 703 3480 704
rect 3474 699 3475 703
rect 3479 699 3480 703
rect 3474 698 3480 699
rect 3476 664 3478 698
rect 3474 663 3480 664
rect 3474 659 3475 663
rect 3479 659 3480 663
rect 3474 658 3480 659
rect 1974 652 1975 656
rect 1979 652 1980 656
rect 1974 651 1980 652
rect 3378 655 3384 656
rect 3378 651 3379 655
rect 3383 651 3384 655
rect 3378 650 3384 651
rect 3406 640 3412 641
rect 3508 640 3510 750
rect 3532 723 3534 800
rect 3652 748 3654 814
rect 3838 813 3839 817
rect 3843 813 3844 817
rect 3838 812 3844 813
rect 3886 816 3892 817
rect 3984 816 3986 938
rect 4156 892 4158 953
rect 4162 939 4168 940
rect 4162 935 4163 939
rect 4167 935 4168 939
rect 4162 934 4168 935
rect 4154 891 4160 892
rect 4154 887 4155 891
rect 4159 887 4160 891
rect 4154 886 4160 887
rect 4164 876 4166 934
rect 4182 876 4188 877
rect 4276 876 4278 974
rect 4364 959 4366 1024
rect 4363 958 4367 959
rect 4363 953 4367 954
rect 4379 958 4383 959
rect 4379 953 4383 954
rect 4380 892 4382 953
rect 4484 944 4486 1038
rect 4580 980 4582 1110
rect 4720 1075 4722 1111
rect 4970 1110 4976 1111
rect 4992 1075 4994 1111
rect 5280 1075 5282 1111
rect 5374 1110 5380 1111
rect 4687 1074 4691 1075
rect 4687 1069 4691 1070
rect 4719 1074 4723 1075
rect 4719 1069 4723 1070
rect 4975 1074 4979 1075
rect 4975 1069 4979 1070
rect 4991 1074 4995 1075
rect 4991 1069 4995 1070
rect 5263 1074 5267 1075
rect 5263 1069 5267 1070
rect 5279 1074 5283 1075
rect 5279 1069 5283 1070
rect 4688 1045 4690 1069
rect 4976 1045 4978 1069
rect 5264 1045 5266 1069
rect 4686 1044 4692 1045
rect 4974 1044 4980 1045
rect 5262 1044 5268 1045
rect 4686 1040 4687 1044
rect 4691 1040 4692 1044
rect 4686 1039 4692 1040
rect 4778 1043 4784 1044
rect 4778 1039 4779 1043
rect 4783 1039 4784 1043
rect 4974 1040 4975 1044
rect 4979 1040 4980 1044
rect 4974 1039 4980 1040
rect 5074 1043 5080 1044
rect 5074 1039 5075 1043
rect 5079 1039 5080 1043
rect 5262 1040 5263 1044
rect 5267 1040 5268 1044
rect 5262 1039 5268 1040
rect 5354 1043 5360 1044
rect 5354 1039 5355 1043
rect 5359 1039 5360 1043
rect 4778 1038 4784 1039
rect 5074 1038 5080 1039
rect 5354 1038 5360 1039
rect 4658 1029 4664 1030
rect 4658 1025 4659 1029
rect 4663 1025 4664 1029
rect 4658 1024 4664 1025
rect 4578 979 4584 980
rect 4578 975 4579 979
rect 4583 975 4584 979
rect 4578 974 4584 975
rect 4660 959 4662 1024
rect 4780 972 4782 1038
rect 4946 1029 4952 1030
rect 4946 1025 4947 1029
rect 4951 1025 4952 1029
rect 4946 1024 4952 1025
rect 4778 971 4784 972
rect 4778 967 4779 971
rect 4783 967 4784 971
rect 4778 966 4784 967
rect 4948 959 4950 1024
rect 5076 980 5078 1038
rect 5234 1029 5240 1030
rect 5234 1025 5235 1029
rect 5239 1025 5240 1029
rect 5234 1024 5240 1025
rect 5074 979 5080 980
rect 5074 975 5075 979
rect 5079 975 5080 979
rect 5074 974 5080 975
rect 5236 959 5238 1024
rect 4595 958 4599 959
rect 4595 953 4599 954
rect 4659 958 4663 959
rect 4659 953 4663 954
rect 4811 958 4815 959
rect 4811 953 4815 954
rect 4947 958 4951 959
rect 4947 953 4951 954
rect 5027 958 5031 959
rect 5027 953 5031 954
rect 5235 958 5239 959
rect 5235 953 5239 954
rect 5243 958 5247 959
rect 5243 953 5247 954
rect 4482 943 4488 944
rect 4482 939 4483 943
rect 4487 939 4488 943
rect 4482 938 4488 939
rect 4596 892 4598 953
rect 4602 939 4608 940
rect 4602 935 4603 939
rect 4607 935 4608 939
rect 4602 934 4608 935
rect 4378 891 4384 892
rect 4378 887 4379 891
rect 4383 887 4384 891
rect 4378 886 4384 887
rect 4594 891 4600 892
rect 4594 887 4595 891
rect 4599 887 4600 891
rect 4594 886 4600 887
rect 4406 876 4412 877
rect 4604 876 4606 934
rect 4812 892 4814 953
rect 4818 939 4824 940
rect 4818 935 4819 939
rect 4823 935 4824 939
rect 4818 934 4824 935
rect 4810 891 4816 892
rect 4810 887 4811 891
rect 4815 887 4816 891
rect 4810 886 4816 887
rect 4622 876 4628 877
rect 4820 876 4822 934
rect 5028 892 5030 953
rect 5244 892 5246 953
rect 5356 944 5358 1038
rect 5376 972 5378 1110
rect 5514 1029 5520 1030
rect 5514 1025 5515 1029
rect 5519 1025 5520 1029
rect 5514 1024 5520 1025
rect 5374 971 5380 972
rect 5374 967 5375 971
rect 5379 967 5380 971
rect 5374 966 5380 967
rect 5516 959 5518 1024
rect 5467 958 5471 959
rect 5467 953 5471 954
rect 5515 958 5519 959
rect 5515 953 5519 954
rect 5354 943 5360 944
rect 5354 939 5355 943
rect 5359 939 5360 943
rect 5354 938 5360 939
rect 5468 892 5470 953
rect 5536 916 5538 1422
rect 5544 1360 5546 1446
rect 5664 1443 5666 1503
rect 5663 1442 5667 1443
rect 5663 1437 5667 1438
rect 5664 1377 5666 1437
rect 5662 1376 5668 1377
rect 5662 1372 5663 1376
rect 5667 1372 5668 1376
rect 5662 1371 5668 1372
rect 5542 1359 5548 1360
rect 5542 1355 5543 1359
rect 5547 1355 5548 1359
rect 5542 1354 5548 1355
rect 5662 1359 5668 1360
rect 5662 1355 5663 1359
rect 5667 1355 5668 1359
rect 5662 1354 5668 1355
rect 5664 1331 5666 1354
rect 5543 1330 5547 1331
rect 5543 1325 5547 1326
rect 5663 1330 5667 1331
rect 5663 1325 5667 1326
rect 5544 1301 5546 1325
rect 5664 1302 5666 1325
rect 5662 1301 5668 1302
rect 5542 1300 5548 1301
rect 5542 1296 5543 1300
rect 5547 1296 5548 1300
rect 5542 1295 5548 1296
rect 5634 1299 5640 1300
rect 5634 1295 5635 1299
rect 5639 1295 5640 1299
rect 5662 1297 5663 1301
rect 5667 1297 5668 1301
rect 5662 1296 5668 1297
rect 5634 1294 5640 1295
rect 5636 1184 5638 1294
rect 5662 1284 5668 1285
rect 5662 1280 5663 1284
rect 5667 1280 5668 1284
rect 5662 1279 5668 1280
rect 5664 1199 5666 1279
rect 5663 1198 5667 1199
rect 5663 1193 5667 1194
rect 5634 1183 5640 1184
rect 5634 1179 5635 1183
rect 5639 1179 5640 1183
rect 5634 1178 5640 1179
rect 5664 1133 5666 1193
rect 5662 1132 5668 1133
rect 5662 1128 5663 1132
rect 5667 1128 5668 1132
rect 5662 1127 5668 1128
rect 5542 1116 5548 1117
rect 5542 1112 5543 1116
rect 5547 1112 5548 1116
rect 5542 1111 5548 1112
rect 5638 1115 5644 1116
rect 5638 1111 5639 1115
rect 5643 1111 5644 1115
rect 5544 1075 5546 1111
rect 5638 1110 5644 1111
rect 5662 1115 5668 1116
rect 5662 1111 5663 1115
rect 5667 1111 5668 1115
rect 5662 1110 5668 1111
rect 5543 1074 5547 1075
rect 5543 1069 5547 1070
rect 5544 1045 5546 1069
rect 5542 1044 5548 1045
rect 5542 1040 5543 1044
rect 5547 1040 5548 1044
rect 5542 1039 5548 1040
rect 5640 980 5642 1110
rect 5664 1075 5666 1110
rect 5663 1074 5667 1075
rect 5663 1069 5667 1070
rect 5664 1046 5666 1069
rect 5662 1045 5668 1046
rect 5662 1041 5663 1045
rect 5667 1041 5668 1045
rect 5662 1040 5668 1041
rect 5646 1035 5652 1036
rect 5646 1031 5647 1035
rect 5651 1031 5652 1035
rect 5646 1030 5652 1031
rect 5638 979 5644 980
rect 5638 975 5639 979
rect 5643 975 5644 979
rect 5638 974 5644 975
rect 5598 943 5604 944
rect 5598 939 5599 943
rect 5603 939 5604 943
rect 5598 938 5604 939
rect 5534 915 5540 916
rect 5534 911 5535 915
rect 5539 911 5540 915
rect 5534 910 5540 911
rect 5590 915 5596 916
rect 5590 911 5591 915
rect 5595 911 5596 915
rect 5590 910 5596 911
rect 5026 891 5032 892
rect 5026 887 5027 891
rect 5031 887 5032 891
rect 5026 886 5032 887
rect 5242 891 5248 892
rect 5242 887 5243 891
rect 5247 887 5248 891
rect 5242 886 5248 887
rect 5466 891 5472 892
rect 5466 887 5467 891
rect 5471 887 5472 891
rect 5466 886 5472 887
rect 4838 876 4844 877
rect 5054 876 5060 877
rect 5270 876 5276 877
rect 4162 875 4168 876
rect 4162 871 4163 875
rect 4167 871 4168 875
rect 4182 872 4183 876
rect 4187 872 4188 876
rect 4182 871 4188 872
rect 4274 875 4280 876
rect 4274 871 4275 875
rect 4279 871 4280 875
rect 4406 872 4407 876
rect 4411 872 4412 876
rect 4406 871 4412 872
rect 4602 875 4608 876
rect 4602 871 4603 875
rect 4607 871 4608 875
rect 4622 872 4623 876
rect 4627 872 4628 876
rect 4622 871 4628 872
rect 4818 875 4824 876
rect 4818 871 4819 875
rect 4823 871 4824 875
rect 4838 872 4839 876
rect 4843 872 4844 876
rect 4838 871 4844 872
rect 4930 875 4936 876
rect 4930 871 4931 875
rect 4935 871 4936 875
rect 5054 872 5055 876
rect 5059 872 5060 876
rect 5054 871 5060 872
rect 5154 875 5160 876
rect 5154 871 5155 875
rect 5159 871 5160 875
rect 5270 872 5271 876
rect 5275 872 5276 876
rect 5270 871 5276 872
rect 5494 876 5500 877
rect 5592 876 5594 910
rect 5494 872 5495 876
rect 5499 872 5500 876
rect 5494 871 5500 872
rect 5590 875 5596 876
rect 5590 871 5591 875
rect 5595 871 5596 875
rect 4162 870 4168 871
rect 4184 847 4186 871
rect 4274 870 4280 871
rect 4408 847 4410 871
rect 4602 870 4608 871
rect 4624 847 4626 871
rect 4818 870 4824 871
rect 4840 847 4842 871
rect 4930 870 4936 871
rect 4111 846 4115 847
rect 4111 841 4115 842
rect 4183 846 4187 847
rect 4183 841 4187 842
rect 4343 846 4347 847
rect 4343 841 4347 842
rect 4407 846 4411 847
rect 4407 841 4411 842
rect 4575 846 4579 847
rect 4575 841 4579 842
rect 4623 846 4627 847
rect 4623 841 4627 842
rect 4799 846 4803 847
rect 4799 841 4803 842
rect 4839 846 4843 847
rect 4839 841 4843 842
rect 4112 817 4114 841
rect 4344 817 4346 841
rect 4576 817 4578 841
rect 4800 817 4802 841
rect 4110 816 4116 817
rect 4342 816 4348 817
rect 3886 812 3887 816
rect 3891 812 3892 816
rect 3886 811 3892 812
rect 3982 815 3988 816
rect 3982 811 3983 815
rect 3987 811 3988 815
rect 4110 812 4111 816
rect 4115 812 4116 816
rect 4110 811 4116 812
rect 4206 815 4212 816
rect 4206 811 4207 815
rect 4211 811 4212 815
rect 4342 812 4343 816
rect 4347 812 4348 816
rect 4342 811 4348 812
rect 4574 816 4580 817
rect 4798 816 4804 817
rect 4574 812 4575 816
rect 4579 812 4580 816
rect 4574 811 4580 812
rect 4674 815 4680 816
rect 4674 811 4675 815
rect 4679 811 4680 815
rect 4798 812 4799 816
rect 4803 812 4804 816
rect 4798 811 4804 812
rect 4890 815 4896 816
rect 4890 811 4891 815
rect 4895 811 4896 815
rect 3982 810 3988 811
rect 4206 810 4212 811
rect 4674 810 4680 811
rect 4890 810 4896 811
rect 3798 804 3804 805
rect 3798 800 3799 804
rect 3803 800 3804 804
rect 3858 801 3864 802
rect 3798 799 3804 800
rect 3838 800 3844 801
rect 3650 747 3656 748
rect 3650 743 3651 747
rect 3655 743 3656 747
rect 3650 742 3656 743
rect 3800 723 3802 799
rect 3838 796 3839 800
rect 3843 796 3844 800
rect 3858 797 3859 801
rect 3863 797 3864 801
rect 3858 796 3864 797
rect 4082 801 4088 802
rect 4082 797 4083 801
rect 4087 797 4088 801
rect 4082 796 4088 797
rect 3838 795 3844 796
rect 3840 735 3842 795
rect 3860 735 3862 796
rect 3954 783 3960 784
rect 3954 779 3955 783
rect 3959 779 3960 783
rect 3954 778 3960 779
rect 3956 752 3958 778
rect 3954 751 3960 752
rect 3954 747 3955 751
rect 3959 747 3960 751
rect 3954 746 3960 747
rect 4084 735 4086 796
rect 4208 784 4210 810
rect 4314 801 4320 802
rect 4314 797 4315 801
rect 4319 797 4320 801
rect 4314 796 4320 797
rect 4546 801 4552 802
rect 4546 797 4547 801
rect 4551 797 4552 801
rect 4546 796 4552 797
rect 4206 783 4212 784
rect 4206 779 4207 783
rect 4211 779 4212 783
rect 4206 778 4212 779
rect 4202 751 4208 752
rect 4202 747 4203 751
rect 4207 747 4208 751
rect 4202 746 4208 747
rect 3839 734 3843 735
rect 3839 729 3843 730
rect 3859 734 3863 735
rect 3859 729 3863 730
rect 4083 734 4087 735
rect 4083 729 4087 730
rect 3515 722 3519 723
rect 3515 717 3519 718
rect 3531 722 3535 723
rect 3531 717 3535 718
rect 3651 722 3655 723
rect 3651 717 3655 718
rect 3799 722 3803 723
rect 3799 717 3803 718
rect 3516 656 3518 717
rect 3638 663 3644 664
rect 3638 659 3639 663
rect 3643 659 3644 663
rect 3638 658 3644 659
rect 3514 655 3520 656
rect 3514 651 3515 655
rect 3519 651 3520 655
rect 3514 650 3520 651
rect 3542 640 3548 641
rect 3640 640 3642 658
rect 3652 656 3654 717
rect 3774 707 3780 708
rect 3774 703 3775 707
rect 3779 703 3780 707
rect 3774 702 3780 703
rect 3650 655 3656 656
rect 3650 651 3651 655
rect 3655 651 3656 655
rect 3650 650 3656 651
rect 3678 640 3684 641
rect 1974 639 1980 640
rect 1934 636 1940 637
rect 1934 632 1935 636
rect 1939 632 1940 636
rect 1974 635 1975 639
rect 1979 635 1980 639
rect 3406 636 3407 640
rect 3411 636 3412 640
rect 3406 635 3412 636
rect 3506 639 3512 640
rect 3506 635 3507 639
rect 3511 635 3512 639
rect 3542 636 3543 640
rect 3547 636 3548 640
rect 3542 635 3548 636
rect 3638 639 3644 640
rect 3638 635 3639 639
rect 3643 635 3644 639
rect 3678 636 3679 640
rect 3683 636 3684 640
rect 3678 635 3684 636
rect 1974 634 1980 635
rect 1934 631 1940 632
rect 1814 620 1820 621
rect 1102 616 1103 620
rect 1107 616 1108 620
rect 1102 615 1108 616
rect 1226 619 1232 620
rect 1226 615 1227 619
rect 1231 615 1232 619
rect 1246 616 1247 620
rect 1251 616 1252 620
rect 1246 615 1252 616
rect 1370 619 1376 620
rect 1370 615 1371 619
rect 1375 615 1376 619
rect 1390 616 1391 620
rect 1395 616 1396 620
rect 1390 615 1396 616
rect 1514 619 1520 620
rect 1514 615 1515 619
rect 1519 615 1520 619
rect 1534 616 1535 620
rect 1539 616 1540 620
rect 1534 615 1540 616
rect 1658 619 1664 620
rect 1658 615 1659 619
rect 1663 615 1664 619
rect 1678 616 1679 620
rect 1683 616 1684 620
rect 1678 615 1684 616
rect 1794 619 1800 620
rect 1794 615 1795 619
rect 1799 615 1800 619
rect 1814 616 1815 620
rect 1819 616 1820 620
rect 1814 615 1820 616
rect 1910 619 1916 620
rect 1910 615 1911 619
rect 1915 615 1916 619
rect 282 614 288 615
rect 304 579 306 615
rect 450 614 456 615
rect 472 579 474 615
rect 562 614 568 615
rect 640 579 642 615
rect 734 614 740 615
rect 303 578 307 579
rect 303 573 307 574
rect 375 578 379 579
rect 375 573 379 574
rect 471 578 475 579
rect 471 573 475 574
rect 599 578 603 579
rect 599 573 603 574
rect 639 578 643 579
rect 639 573 643 574
rect 376 549 378 573
rect 600 549 602 573
rect 374 548 380 549
rect 598 548 604 549
rect 158 544 159 548
rect 163 544 164 548
rect 158 543 164 544
rect 254 547 260 548
rect 254 543 255 547
rect 259 543 260 547
rect 374 544 375 548
rect 379 544 380 548
rect 374 543 380 544
rect 466 547 472 548
rect 466 543 467 547
rect 471 543 472 547
rect 598 544 599 548
rect 603 544 604 548
rect 598 543 604 544
rect 698 547 704 548
rect 698 543 699 547
rect 703 543 704 547
rect 254 542 260 543
rect 466 542 472 543
rect 698 542 704 543
rect 130 533 136 534
rect 110 532 116 533
rect 110 528 111 532
rect 115 528 116 532
rect 130 529 131 533
rect 135 529 136 533
rect 130 528 136 529
rect 346 533 352 534
rect 346 529 347 533
rect 351 529 352 533
rect 346 528 352 529
rect 110 527 116 528
rect 112 467 114 527
rect 132 467 134 528
rect 348 467 350 528
rect 468 476 470 542
rect 570 533 576 534
rect 570 529 571 533
rect 575 529 576 533
rect 570 528 576 529
rect 466 475 472 476
rect 466 471 467 475
rect 471 471 472 475
rect 466 470 472 471
rect 572 467 574 528
rect 700 484 702 542
rect 736 492 738 614
rect 800 579 802 615
rect 952 579 954 615
rect 1104 579 1106 615
rect 1226 614 1232 615
rect 1248 579 1250 615
rect 1370 614 1376 615
rect 1392 579 1394 615
rect 1514 614 1520 615
rect 1536 579 1538 615
rect 1658 614 1664 615
rect 1680 579 1682 615
rect 1794 614 1800 615
rect 1816 579 1818 615
rect 1910 614 1916 615
rect 1934 619 1940 620
rect 1934 615 1935 619
rect 1939 615 1940 619
rect 1934 614 1940 615
rect 799 578 803 579
rect 799 573 803 574
rect 807 578 811 579
rect 807 573 811 574
rect 951 578 955 579
rect 951 573 955 574
rect 999 578 1003 579
rect 999 573 1003 574
rect 1103 578 1107 579
rect 1103 573 1107 574
rect 1175 578 1179 579
rect 1175 573 1179 574
rect 1247 578 1251 579
rect 1247 573 1251 574
rect 1343 578 1347 579
rect 1343 573 1347 574
rect 1391 578 1395 579
rect 1391 573 1395 574
rect 1511 578 1515 579
rect 1511 573 1515 574
rect 1535 578 1539 579
rect 1535 573 1539 574
rect 1671 578 1675 579
rect 1671 573 1675 574
rect 1679 578 1683 579
rect 1679 573 1683 574
rect 1815 578 1819 579
rect 1815 573 1819 574
rect 808 549 810 573
rect 1000 549 1002 573
rect 1176 549 1178 573
rect 1344 549 1346 573
rect 1512 549 1514 573
rect 1672 549 1674 573
rect 1816 549 1818 573
rect 806 548 812 549
rect 998 548 1004 549
rect 1174 548 1180 549
rect 1342 548 1348 549
rect 1510 548 1516 549
rect 1670 548 1676 549
rect 1814 548 1820 549
rect 806 544 807 548
rect 811 544 812 548
rect 806 543 812 544
rect 934 547 940 548
rect 934 543 935 547
rect 939 543 940 547
rect 998 544 999 548
rect 1003 544 1004 548
rect 998 543 1004 544
rect 1094 547 1100 548
rect 1094 543 1095 547
rect 1099 543 1100 547
rect 1174 544 1175 548
rect 1179 544 1180 548
rect 1174 543 1180 544
rect 1274 547 1280 548
rect 1274 543 1275 547
rect 1279 543 1280 547
rect 1342 544 1343 548
rect 1347 544 1348 548
rect 1342 543 1348 544
rect 1442 547 1448 548
rect 1442 543 1443 547
rect 1447 543 1448 547
rect 1510 544 1511 548
rect 1515 544 1516 548
rect 1510 543 1516 544
rect 1610 547 1616 548
rect 1610 543 1611 547
rect 1615 543 1616 547
rect 1670 544 1671 548
rect 1675 544 1676 548
rect 1670 543 1676 544
rect 1770 547 1776 548
rect 1770 543 1771 547
rect 1775 543 1776 547
rect 1814 544 1815 548
rect 1819 544 1820 548
rect 1814 543 1820 544
rect 934 542 940 543
rect 1094 542 1100 543
rect 1274 542 1280 543
rect 1442 542 1448 543
rect 1610 542 1616 543
rect 1770 542 1776 543
rect 778 533 784 534
rect 778 529 779 533
rect 783 529 784 533
rect 778 528 784 529
rect 734 491 740 492
rect 734 487 735 491
rect 739 487 740 491
rect 734 486 740 487
rect 698 483 704 484
rect 698 479 699 483
rect 703 479 704 483
rect 698 478 704 479
rect 780 467 782 528
rect 936 484 938 542
rect 970 533 976 534
rect 970 529 971 533
rect 975 529 976 533
rect 970 528 976 529
rect 934 483 940 484
rect 934 479 935 483
rect 939 479 940 483
rect 934 478 940 479
rect 972 467 974 528
rect 111 466 115 467
rect 111 461 115 462
rect 131 466 135 467
rect 131 461 135 462
rect 195 466 199 467
rect 195 461 199 462
rect 347 466 351 467
rect 347 461 351 462
rect 475 466 479 467
rect 475 461 479 462
rect 571 466 575 467
rect 571 461 575 462
rect 755 466 759 467
rect 755 461 759 462
rect 779 466 783 467
rect 779 461 783 462
rect 971 466 975 467
rect 971 461 975 462
rect 1043 466 1047 467
rect 1043 461 1047 462
rect 112 401 114 461
rect 110 400 116 401
rect 196 400 198 461
rect 476 400 478 461
rect 598 451 604 452
rect 598 447 599 451
rect 603 447 604 451
rect 598 446 604 447
rect 110 396 111 400
rect 115 396 116 400
rect 110 395 116 396
rect 194 399 200 400
rect 194 395 195 399
rect 199 395 200 399
rect 194 394 200 395
rect 474 399 480 400
rect 474 395 475 399
rect 479 395 480 399
rect 474 394 480 395
rect 222 384 228 385
rect 110 383 116 384
rect 110 379 111 383
rect 115 379 116 383
rect 222 380 223 384
rect 227 380 228 384
rect 222 379 228 380
rect 502 384 508 385
rect 502 380 503 384
rect 507 380 508 384
rect 502 379 508 380
rect 110 378 116 379
rect 112 355 114 378
rect 224 355 226 379
rect 504 355 506 379
rect 111 354 115 355
rect 111 349 115 350
rect 223 354 227 355
rect 223 349 227 350
rect 311 354 315 355
rect 311 349 315 350
rect 503 354 507 355
rect 503 349 507 350
rect 112 326 114 349
rect 110 325 116 326
rect 312 325 314 349
rect 504 325 506 349
rect 110 321 111 325
rect 115 321 116 325
rect 110 320 116 321
rect 310 324 316 325
rect 502 324 508 325
rect 600 324 602 446
rect 756 400 758 461
rect 1044 400 1046 461
rect 1096 452 1098 542
rect 1146 533 1152 534
rect 1146 529 1147 533
rect 1151 529 1152 533
rect 1146 528 1152 529
rect 1148 467 1150 528
rect 1276 484 1278 542
rect 1314 533 1320 534
rect 1314 529 1315 533
rect 1319 529 1320 533
rect 1314 528 1320 529
rect 1274 483 1280 484
rect 1274 479 1275 483
rect 1279 479 1280 483
rect 1274 478 1280 479
rect 1316 467 1318 528
rect 1444 484 1446 542
rect 1482 533 1488 534
rect 1482 529 1483 533
rect 1487 529 1488 533
rect 1482 528 1488 529
rect 1442 483 1448 484
rect 1442 479 1443 483
rect 1447 479 1448 483
rect 1442 478 1448 479
rect 1484 467 1486 528
rect 1612 484 1614 542
rect 1642 533 1648 534
rect 1642 529 1643 533
rect 1647 529 1648 533
rect 1642 528 1648 529
rect 1610 483 1616 484
rect 1610 479 1611 483
rect 1615 479 1616 483
rect 1610 478 1616 479
rect 1644 467 1646 528
rect 1772 484 1774 542
rect 1786 533 1792 534
rect 1786 529 1787 533
rect 1791 529 1792 533
rect 1786 528 1792 529
rect 1770 483 1776 484
rect 1770 479 1771 483
rect 1775 479 1776 483
rect 1770 478 1776 479
rect 1788 467 1790 528
rect 1912 476 1914 614
rect 1936 579 1938 614
rect 1976 603 1978 634
rect 3408 603 3410 635
rect 3506 634 3512 635
rect 3544 603 3546 635
rect 3638 634 3644 635
rect 3680 603 3682 635
rect 1975 602 1979 603
rect 1975 597 1979 598
rect 3271 602 3275 603
rect 3271 597 3275 598
rect 3407 602 3411 603
rect 3407 597 3411 598
rect 3543 602 3547 603
rect 3543 597 3547 598
rect 3679 602 3683 603
rect 3679 597 3683 598
rect 1935 578 1939 579
rect 1976 574 1978 597
rect 1935 573 1939 574
rect 1974 573 1980 574
rect 3272 573 3274 597
rect 3408 573 3410 597
rect 3544 573 3546 597
rect 3680 573 3682 597
rect 1936 550 1938 573
rect 1974 569 1975 573
rect 1979 569 1980 573
rect 1974 568 1980 569
rect 3270 572 3276 573
rect 3406 572 3412 573
rect 3542 572 3548 573
rect 3678 572 3684 573
rect 3776 572 3778 702
rect 3800 657 3802 717
rect 3840 669 3842 729
rect 3838 668 3844 669
rect 3860 668 3862 729
rect 3982 719 3988 720
rect 3982 715 3983 719
rect 3987 715 3988 719
rect 3982 714 3988 715
rect 3838 664 3839 668
rect 3843 664 3844 668
rect 3838 663 3844 664
rect 3858 667 3864 668
rect 3858 663 3859 667
rect 3863 663 3864 667
rect 3858 662 3864 663
rect 3798 656 3804 657
rect 3798 652 3799 656
rect 3803 652 3804 656
rect 3886 652 3892 653
rect 3798 651 3804 652
rect 3838 651 3844 652
rect 3838 647 3839 651
rect 3843 647 3844 651
rect 3886 648 3887 652
rect 3891 648 3892 652
rect 3886 647 3892 648
rect 3838 646 3844 647
rect 3798 639 3804 640
rect 3798 635 3799 639
rect 3803 635 3804 639
rect 3798 634 3804 635
rect 3800 603 3802 634
rect 3840 615 3842 646
rect 3888 615 3890 647
rect 3839 614 3843 615
rect 3839 609 3843 610
rect 3887 614 3891 615
rect 3887 609 3891 610
rect 3799 602 3803 603
rect 3799 597 3803 598
rect 3800 574 3802 597
rect 3840 586 3842 609
rect 3838 585 3844 586
rect 3888 585 3890 609
rect 3838 581 3839 585
rect 3843 581 3844 585
rect 3838 580 3844 581
rect 3886 584 3892 585
rect 3984 584 3986 714
rect 4084 668 4086 729
rect 4090 715 4096 716
rect 4090 711 4091 715
rect 4095 711 4096 715
rect 4090 710 4096 711
rect 4082 667 4088 668
rect 4082 663 4083 667
rect 4087 663 4088 667
rect 4082 662 4088 663
rect 4092 652 4094 710
rect 4110 652 4116 653
rect 4204 652 4206 746
rect 4316 735 4318 796
rect 4548 735 4550 796
rect 4676 752 4678 810
rect 4770 801 4776 802
rect 4770 797 4771 801
rect 4775 797 4776 801
rect 4770 796 4776 797
rect 4674 751 4680 752
rect 4674 747 4675 751
rect 4679 747 4680 751
rect 4674 746 4680 747
rect 4650 735 4656 736
rect 4772 735 4774 796
rect 4315 734 4319 735
rect 4315 729 4319 730
rect 4323 734 4327 735
rect 4323 729 4327 730
rect 4547 734 4551 735
rect 4547 729 4551 730
rect 4555 734 4559 735
rect 4650 731 4651 735
rect 4655 731 4656 735
rect 4650 730 4656 731
rect 4771 734 4775 735
rect 4555 729 4559 730
rect 4324 668 4326 729
rect 4556 668 4558 729
rect 4652 716 4654 730
rect 4771 729 4775 730
rect 4779 734 4783 735
rect 4779 729 4783 730
rect 4678 723 4684 724
rect 4678 719 4679 723
rect 4683 719 4684 723
rect 4678 718 4684 719
rect 4650 715 4656 716
rect 4650 711 4651 715
rect 4655 711 4656 715
rect 4650 710 4656 711
rect 4322 667 4328 668
rect 4322 663 4323 667
rect 4327 663 4328 667
rect 4322 662 4328 663
rect 4554 667 4560 668
rect 4554 663 4555 667
rect 4559 663 4560 667
rect 4554 662 4560 663
rect 4350 652 4356 653
rect 4582 652 4588 653
rect 4680 652 4682 718
rect 4780 668 4782 729
rect 4892 720 4894 810
rect 4932 744 4934 870
rect 5056 847 5058 871
rect 5154 870 5160 871
rect 5031 846 5035 847
rect 5031 841 5035 842
rect 5055 846 5059 847
rect 5055 841 5059 842
rect 5032 817 5034 841
rect 5030 816 5036 817
rect 5030 812 5031 816
rect 5035 812 5036 816
rect 5030 811 5036 812
rect 5122 815 5128 816
rect 5122 811 5123 815
rect 5127 811 5128 815
rect 5122 810 5128 811
rect 5002 801 5008 802
rect 5002 797 5003 801
rect 5007 797 5008 801
rect 5002 796 5008 797
rect 4930 743 4936 744
rect 4930 739 4931 743
rect 4935 739 4936 743
rect 4930 738 4936 739
rect 5004 735 5006 796
rect 5124 736 5126 810
rect 5156 752 5158 870
rect 5272 847 5274 871
rect 5496 847 5498 871
rect 5590 870 5596 871
rect 5263 846 5267 847
rect 5263 841 5267 842
rect 5271 846 5275 847
rect 5271 841 5275 842
rect 5495 846 5499 847
rect 5495 841 5499 842
rect 5264 817 5266 841
rect 5496 817 5498 841
rect 5262 816 5268 817
rect 5494 816 5500 817
rect 5262 812 5263 816
rect 5267 812 5268 816
rect 5262 811 5268 812
rect 5354 815 5360 816
rect 5354 811 5355 815
rect 5359 811 5360 815
rect 5494 812 5495 816
rect 5499 812 5500 816
rect 5494 811 5500 812
rect 5591 815 5597 816
rect 5591 811 5592 815
rect 5596 814 5597 815
rect 5600 814 5602 938
rect 5596 812 5602 814
rect 5596 811 5597 812
rect 5354 810 5360 811
rect 5591 810 5597 811
rect 5234 801 5240 802
rect 5234 797 5235 801
rect 5239 797 5240 801
rect 5234 796 5240 797
rect 5154 751 5160 752
rect 5154 747 5155 751
rect 5159 747 5160 751
rect 5154 746 5160 747
rect 5122 735 5128 736
rect 5236 735 5238 796
rect 5356 744 5358 810
rect 5466 801 5472 802
rect 5466 797 5467 801
rect 5471 797 5472 801
rect 5466 796 5472 797
rect 5354 743 5360 744
rect 5354 739 5355 743
rect 5359 739 5360 743
rect 5354 738 5360 739
rect 5468 735 5470 796
rect 5648 752 5650 1030
rect 5662 1028 5668 1029
rect 5662 1024 5663 1028
rect 5667 1024 5668 1028
rect 5662 1023 5668 1024
rect 5664 959 5666 1023
rect 5663 958 5667 959
rect 5663 953 5667 954
rect 5664 893 5666 953
rect 5662 892 5668 893
rect 5662 888 5663 892
rect 5667 888 5668 892
rect 5662 887 5668 888
rect 5662 875 5668 876
rect 5662 871 5663 875
rect 5667 871 5668 875
rect 5662 870 5668 871
rect 5664 847 5666 870
rect 5663 846 5667 847
rect 5663 841 5667 842
rect 5664 818 5666 841
rect 5662 817 5668 818
rect 5662 813 5663 817
rect 5667 813 5668 817
rect 5662 812 5668 813
rect 5662 800 5668 801
rect 5662 796 5663 800
rect 5667 796 5668 800
rect 5662 795 5668 796
rect 5646 751 5652 752
rect 5646 747 5647 751
rect 5651 747 5652 751
rect 5646 746 5652 747
rect 5664 735 5666 795
rect 5003 734 5007 735
rect 5122 731 5123 735
rect 5127 731 5128 735
rect 5122 730 5128 731
rect 5227 734 5231 735
rect 5003 729 5007 730
rect 5227 729 5231 730
rect 5235 734 5239 735
rect 5235 729 5239 730
rect 5459 734 5463 735
rect 5459 729 5463 730
rect 5467 734 5471 735
rect 5467 729 5471 730
rect 5663 734 5667 735
rect 5663 729 5667 730
rect 4890 719 4896 720
rect 4890 715 4891 719
rect 4895 715 4896 719
rect 4890 714 4896 715
rect 5004 668 5006 729
rect 5010 715 5016 716
rect 5010 711 5011 715
rect 5015 711 5016 715
rect 5010 710 5016 711
rect 4778 667 4784 668
rect 4778 663 4779 667
rect 4783 663 4784 667
rect 4778 662 4784 663
rect 5002 667 5008 668
rect 5002 663 5003 667
rect 5007 663 5008 667
rect 5002 662 5008 663
rect 4806 652 4812 653
rect 5012 652 5014 710
rect 5228 668 5230 729
rect 5234 715 5240 716
rect 5234 711 5235 715
rect 5239 711 5240 715
rect 5234 710 5240 711
rect 5226 667 5232 668
rect 5226 663 5227 667
rect 5231 663 5232 667
rect 5226 662 5232 663
rect 5030 652 5036 653
rect 5236 652 5238 710
rect 5460 668 5462 729
rect 5638 719 5644 720
rect 5638 715 5639 719
rect 5643 715 5644 719
rect 5638 714 5644 715
rect 5458 667 5464 668
rect 5458 663 5459 667
rect 5463 663 5464 667
rect 5458 662 5464 663
rect 5254 652 5260 653
rect 5486 652 5492 653
rect 4090 651 4096 652
rect 4090 647 4091 651
rect 4095 647 4096 651
rect 4110 648 4111 652
rect 4115 648 4116 652
rect 4110 647 4116 648
rect 4202 651 4208 652
rect 4202 647 4203 651
rect 4207 647 4208 651
rect 4350 648 4351 652
rect 4355 648 4356 652
rect 4350 647 4356 648
rect 4446 651 4452 652
rect 4446 647 4447 651
rect 4451 647 4452 651
rect 4582 648 4583 652
rect 4587 648 4588 652
rect 4582 647 4588 648
rect 4678 651 4684 652
rect 4678 647 4679 651
rect 4683 647 4684 651
rect 4806 648 4807 652
rect 4811 648 4812 652
rect 4806 647 4812 648
rect 5010 651 5016 652
rect 5010 647 5011 651
rect 5015 647 5016 651
rect 5030 648 5031 652
rect 5035 648 5036 652
rect 5030 647 5036 648
rect 5234 651 5240 652
rect 5234 647 5235 651
rect 5239 647 5240 651
rect 5254 648 5255 652
rect 5259 648 5260 652
rect 5254 647 5260 648
rect 5346 651 5352 652
rect 5346 647 5347 651
rect 5351 647 5352 651
rect 5486 648 5487 652
rect 5491 648 5492 652
rect 5486 647 5492 648
rect 5582 651 5588 652
rect 5582 647 5583 651
rect 5587 647 5588 651
rect 4090 646 4096 647
rect 4112 615 4114 647
rect 4202 646 4208 647
rect 4352 615 4354 647
rect 4446 646 4452 647
rect 4111 614 4115 615
rect 4111 609 4115 610
rect 4143 614 4147 615
rect 4143 609 4147 610
rect 4351 614 4355 615
rect 4351 609 4355 610
rect 4407 614 4411 615
rect 4407 609 4411 610
rect 4144 585 4146 609
rect 4408 585 4410 609
rect 4142 584 4148 585
rect 4406 584 4412 585
rect 3886 580 3887 584
rect 3891 580 3892 584
rect 3886 579 3892 580
rect 3982 583 3988 584
rect 3982 579 3983 583
rect 3987 579 3988 583
rect 4142 580 4143 584
rect 4147 580 4148 584
rect 4142 579 4148 580
rect 4238 583 4244 584
rect 4238 579 4239 583
rect 4243 579 4244 583
rect 4406 580 4407 584
rect 4411 580 4412 584
rect 4406 579 4412 580
rect 3982 578 3988 579
rect 4238 578 4244 579
rect 3798 573 3804 574
rect 3270 568 3271 572
rect 3275 568 3276 572
rect 3270 567 3276 568
rect 3370 571 3376 572
rect 3370 567 3371 571
rect 3375 567 3376 571
rect 3406 568 3407 572
rect 3411 568 3412 572
rect 3406 567 3412 568
rect 3506 571 3512 572
rect 3506 567 3507 571
rect 3511 567 3512 571
rect 3542 568 3543 572
rect 3547 568 3548 572
rect 3542 567 3548 568
rect 3642 571 3648 572
rect 3642 567 3643 571
rect 3647 567 3648 571
rect 3678 568 3679 572
rect 3683 568 3684 572
rect 3678 567 3684 568
rect 3774 571 3780 572
rect 3774 567 3775 571
rect 3779 567 3780 571
rect 3798 569 3799 573
rect 3803 569 3804 573
rect 3858 569 3864 570
rect 3798 568 3804 569
rect 3838 568 3844 569
rect 3370 566 3376 567
rect 3506 566 3512 567
rect 3642 566 3648 567
rect 3774 566 3780 567
rect 3242 557 3248 558
rect 1974 556 1980 557
rect 1974 552 1975 556
rect 1979 552 1980 556
rect 3242 553 3243 557
rect 3247 553 3248 557
rect 3242 552 3248 553
rect 1974 551 1980 552
rect 1934 549 1940 550
rect 1926 547 1932 548
rect 1926 543 1927 547
rect 1931 543 1932 547
rect 1934 545 1935 549
rect 1939 545 1940 549
rect 1934 544 1940 545
rect 1926 542 1932 543
rect 1910 475 1916 476
rect 1910 471 1911 475
rect 1915 471 1916 475
rect 1910 470 1916 471
rect 1147 466 1151 467
rect 1147 461 1151 462
rect 1315 466 1319 467
rect 1315 461 1319 462
rect 1331 466 1335 467
rect 1331 461 1335 462
rect 1483 466 1487 467
rect 1483 461 1487 462
rect 1643 466 1647 467
rect 1643 461 1647 462
rect 1787 466 1791 467
rect 1787 461 1791 462
rect 1094 451 1100 452
rect 1094 447 1095 451
rect 1099 447 1100 451
rect 1094 446 1100 447
rect 1332 400 1334 461
rect 1928 456 1930 542
rect 1934 532 1940 533
rect 1934 528 1935 532
rect 1939 528 1940 532
rect 1934 527 1940 528
rect 1936 467 1938 527
rect 1976 471 1978 551
rect 3244 471 3246 552
rect 3372 508 3374 566
rect 3378 557 3384 558
rect 3378 553 3379 557
rect 3383 553 3384 557
rect 3378 552 3384 553
rect 3370 507 3376 508
rect 3370 503 3371 507
rect 3375 503 3376 507
rect 3370 502 3376 503
rect 3380 471 3382 552
rect 3508 508 3510 566
rect 3514 557 3520 558
rect 3514 553 3515 557
rect 3519 553 3520 557
rect 3514 552 3520 553
rect 3506 507 3512 508
rect 3506 503 3507 507
rect 3511 503 3512 507
rect 3506 502 3512 503
rect 3516 471 3518 552
rect 3644 508 3646 566
rect 3838 564 3839 568
rect 3843 564 3844 568
rect 3858 565 3859 569
rect 3863 565 3864 569
rect 3858 564 3864 565
rect 4114 569 4120 570
rect 4114 565 4115 569
rect 4119 565 4120 569
rect 4114 564 4120 565
rect 3838 563 3844 564
rect 3650 557 3656 558
rect 3650 553 3651 557
rect 3655 553 3656 557
rect 3650 552 3656 553
rect 3798 556 3804 557
rect 3798 552 3799 556
rect 3803 552 3804 556
rect 3642 507 3648 508
rect 3642 503 3643 507
rect 3647 503 3648 507
rect 3642 502 3648 503
rect 3652 471 3654 552
rect 3798 551 3804 552
rect 3658 499 3664 500
rect 3658 495 3659 499
rect 3663 495 3664 499
rect 3658 494 3664 495
rect 1975 470 1979 471
rect 1935 466 1939 467
rect 1975 465 1979 466
rect 1995 470 1999 471
rect 1995 465 1999 466
rect 2155 470 2159 471
rect 2155 465 2159 466
rect 2347 470 2351 471
rect 2347 465 2351 466
rect 2539 470 2543 471
rect 2539 465 2543 466
rect 2739 470 2743 471
rect 2739 465 2743 466
rect 2931 470 2935 471
rect 2931 465 2935 466
rect 3131 470 3135 471
rect 3131 465 3135 466
rect 3243 470 3247 471
rect 3243 465 3247 466
rect 3331 470 3335 471
rect 3331 465 3335 466
rect 3379 470 3383 471
rect 3379 465 3383 466
rect 3515 470 3519 471
rect 3515 465 3519 466
rect 3531 470 3535 471
rect 3531 465 3535 466
rect 3651 470 3655 471
rect 3651 465 3655 466
rect 1935 461 1939 462
rect 1926 455 1932 456
rect 1926 451 1927 455
rect 1931 451 1932 455
rect 1926 450 1932 451
rect 1338 447 1344 448
rect 1338 443 1339 447
rect 1343 443 1344 447
rect 1338 442 1344 443
rect 754 399 760 400
rect 754 395 755 399
rect 759 395 760 399
rect 754 394 760 395
rect 1042 399 1048 400
rect 1042 395 1043 399
rect 1047 395 1048 399
rect 1042 394 1048 395
rect 1330 399 1336 400
rect 1330 395 1331 399
rect 1335 395 1336 399
rect 1330 394 1336 395
rect 782 384 788 385
rect 1070 384 1076 385
rect 1340 384 1342 442
rect 1936 401 1938 461
rect 1976 405 1978 465
rect 1974 404 1980 405
rect 1996 404 1998 465
rect 2156 404 2158 465
rect 2162 451 2168 452
rect 2162 447 2163 451
rect 2167 447 2168 451
rect 2162 446 2168 447
rect 1934 400 1940 401
rect 1934 396 1935 400
rect 1939 396 1940 400
rect 1974 400 1975 404
rect 1979 400 1980 404
rect 1974 399 1980 400
rect 1994 403 2000 404
rect 1994 399 1995 403
rect 1999 399 2000 403
rect 1994 398 2000 399
rect 2154 403 2160 404
rect 2154 399 2155 403
rect 2159 399 2160 403
rect 2154 398 2160 399
rect 1934 395 1940 396
rect 2022 388 2028 389
rect 2164 388 2166 446
rect 2348 404 2350 465
rect 2354 451 2360 452
rect 2354 447 2355 451
rect 2359 447 2360 451
rect 2354 446 2360 447
rect 2346 403 2352 404
rect 2346 399 2347 403
rect 2351 399 2352 403
rect 2346 398 2352 399
rect 2182 388 2188 389
rect 2356 388 2358 446
rect 2540 404 2542 465
rect 2546 451 2552 452
rect 2546 447 2547 451
rect 2551 447 2552 451
rect 2546 446 2552 447
rect 2538 403 2544 404
rect 2538 399 2539 403
rect 2543 399 2544 403
rect 2538 398 2544 399
rect 2374 388 2380 389
rect 2548 388 2550 446
rect 2740 404 2742 465
rect 2746 451 2752 452
rect 2746 447 2747 451
rect 2751 447 2752 451
rect 2746 446 2752 447
rect 2738 403 2744 404
rect 2738 399 2739 403
rect 2743 399 2744 403
rect 2738 398 2744 399
rect 2566 388 2572 389
rect 2748 388 2750 446
rect 2932 404 2934 465
rect 3014 455 3020 456
rect 3014 451 3015 455
rect 3019 451 3020 455
rect 3014 450 3020 451
rect 2930 403 2936 404
rect 2930 399 2931 403
rect 2935 399 2936 403
rect 2930 398 2936 399
rect 2766 388 2772 389
rect 2958 388 2964 389
rect 1974 387 1980 388
rect 1358 384 1364 385
rect 782 380 783 384
rect 787 380 788 384
rect 782 379 788 380
rect 878 383 884 384
rect 878 379 879 383
rect 883 379 884 383
rect 1070 380 1071 384
rect 1075 380 1076 384
rect 1070 379 1076 380
rect 1338 383 1344 384
rect 1338 379 1339 383
rect 1343 379 1344 383
rect 1358 380 1359 384
rect 1363 380 1364 384
rect 1358 379 1364 380
rect 1934 383 1940 384
rect 1934 379 1935 383
rect 1939 379 1940 383
rect 1974 383 1975 387
rect 1979 383 1980 387
rect 2022 384 2023 388
rect 2027 384 2028 388
rect 2022 383 2028 384
rect 2162 387 2168 388
rect 2162 383 2163 387
rect 2167 383 2168 387
rect 2182 384 2183 388
rect 2187 384 2188 388
rect 2182 383 2188 384
rect 2354 387 2360 388
rect 2354 383 2355 387
rect 2359 383 2360 387
rect 2374 384 2375 388
rect 2379 384 2380 388
rect 2374 383 2380 384
rect 2546 387 2552 388
rect 2546 383 2547 387
rect 2551 383 2552 387
rect 2566 384 2567 388
rect 2571 384 2572 388
rect 2566 383 2572 384
rect 2746 387 2752 388
rect 2746 383 2747 387
rect 2751 383 2752 387
rect 2766 384 2767 388
rect 2771 384 2772 388
rect 2766 383 2772 384
rect 2858 387 2864 388
rect 2858 383 2859 387
rect 2863 383 2864 387
rect 2958 384 2959 388
rect 2963 384 2964 388
rect 2958 383 2964 384
rect 1974 382 1980 383
rect 784 355 786 379
rect 878 378 884 379
rect 695 354 699 355
rect 695 349 699 350
rect 783 354 787 355
rect 783 349 787 350
rect 696 325 698 349
rect 694 324 700 325
rect 310 320 311 324
rect 315 320 316 324
rect 310 319 316 320
rect 430 323 436 324
rect 430 319 431 323
rect 435 319 436 323
rect 502 320 503 324
rect 507 320 508 324
rect 502 319 508 320
rect 598 323 604 324
rect 598 319 599 323
rect 603 319 604 323
rect 694 320 695 324
rect 699 320 700 324
rect 694 319 700 320
rect 430 318 436 319
rect 598 318 604 319
rect 282 309 288 310
rect 110 308 116 309
rect 110 304 111 308
rect 115 304 116 308
rect 282 305 283 309
rect 287 305 288 309
rect 282 304 288 305
rect 110 303 116 304
rect 112 207 114 303
rect 284 207 286 304
rect 432 260 434 318
rect 474 309 480 310
rect 474 305 475 309
rect 479 305 480 309
rect 474 304 480 305
rect 666 309 672 310
rect 666 305 667 309
rect 671 305 672 309
rect 666 304 672 305
rect 858 309 864 310
rect 858 305 859 309
rect 863 305 864 309
rect 858 304 864 305
rect 386 259 392 260
rect 386 255 387 259
rect 391 255 392 259
rect 386 254 392 255
rect 430 259 436 260
rect 430 255 431 259
rect 435 255 436 259
rect 430 254 436 255
rect 111 206 115 207
rect 111 201 115 202
rect 131 206 135 207
rect 131 201 135 202
rect 267 206 271 207
rect 267 201 271 202
rect 283 206 287 207
rect 283 201 287 202
rect 112 141 114 201
rect 110 140 116 141
rect 132 140 134 201
rect 268 140 270 201
rect 274 187 280 188
rect 274 183 275 187
rect 279 183 280 187
rect 274 182 280 183
rect 110 136 111 140
rect 115 136 116 140
rect 110 135 116 136
rect 130 139 136 140
rect 130 135 131 139
rect 135 135 136 139
rect 130 134 136 135
rect 266 139 272 140
rect 266 135 267 139
rect 271 135 272 139
rect 266 134 272 135
rect 158 124 164 125
rect 276 124 278 182
rect 294 124 300 125
rect 388 124 390 254
rect 476 207 478 304
rect 668 207 670 304
rect 860 207 862 304
rect 880 260 882 378
rect 1072 355 1074 379
rect 1338 378 1344 379
rect 1360 355 1362 379
rect 1934 378 1940 379
rect 1936 355 1938 378
rect 887 354 891 355
rect 887 349 891 350
rect 1071 354 1075 355
rect 1071 349 1075 350
rect 1079 354 1083 355
rect 1079 349 1083 350
rect 1359 354 1363 355
rect 1359 349 1363 350
rect 1935 354 1939 355
rect 1935 349 1939 350
rect 888 325 890 349
rect 1080 325 1082 349
rect 1936 326 1938 349
rect 1976 335 1978 382
rect 2024 335 2026 383
rect 2162 382 2168 383
rect 2184 335 2186 383
rect 2354 382 2360 383
rect 2376 335 2378 383
rect 2546 382 2552 383
rect 2568 335 2570 383
rect 2746 382 2752 383
rect 2768 335 2770 383
rect 2858 382 2864 383
rect 1975 334 1979 335
rect 1975 329 1979 330
rect 2023 334 2027 335
rect 2023 329 2027 330
rect 2159 334 2163 335
rect 2159 329 2163 330
rect 2183 334 2187 335
rect 2183 329 2187 330
rect 2295 334 2299 335
rect 2295 329 2299 330
rect 2375 334 2379 335
rect 2375 329 2379 330
rect 2431 334 2435 335
rect 2431 329 2435 330
rect 2567 334 2571 335
rect 2567 329 2571 330
rect 2703 334 2707 335
rect 2703 329 2707 330
rect 2767 334 2771 335
rect 2767 329 2771 330
rect 2839 334 2843 335
rect 2839 329 2843 330
rect 1934 325 1940 326
rect 886 324 892 325
rect 886 320 887 324
rect 891 320 892 324
rect 886 319 892 320
rect 1078 324 1084 325
rect 1078 320 1079 324
rect 1083 320 1084 324
rect 1078 319 1084 320
rect 1174 323 1180 324
rect 1174 319 1175 323
rect 1179 319 1180 323
rect 1934 321 1935 325
rect 1939 321 1940 325
rect 1934 320 1940 321
rect 1174 318 1180 319
rect 1050 309 1056 310
rect 1050 305 1051 309
rect 1055 305 1056 309
rect 1050 304 1056 305
rect 878 259 884 260
rect 878 255 879 259
rect 883 255 884 259
rect 878 254 884 255
rect 1052 207 1054 304
rect 1176 252 1178 318
rect 1934 308 1940 309
rect 1934 304 1935 308
rect 1939 304 1940 308
rect 1976 306 1978 329
rect 1934 303 1940 304
rect 1974 305 1980 306
rect 2024 305 2026 329
rect 2160 305 2162 329
rect 2296 305 2298 329
rect 2432 305 2434 329
rect 2568 305 2570 329
rect 2704 305 2706 329
rect 2840 305 2842 329
rect 1174 251 1180 252
rect 1174 247 1175 251
rect 1179 247 1180 251
rect 1174 246 1180 247
rect 1936 207 1938 303
rect 1974 301 1975 305
rect 1979 301 1980 305
rect 1974 300 1980 301
rect 2022 304 2028 305
rect 2158 304 2164 305
rect 2294 304 2300 305
rect 2430 304 2436 305
rect 2566 304 2572 305
rect 2702 304 2708 305
rect 2838 304 2844 305
rect 2022 300 2023 304
rect 2027 300 2028 304
rect 2022 299 2028 300
rect 2122 303 2128 304
rect 2122 299 2123 303
rect 2127 299 2128 303
rect 2158 300 2159 304
rect 2163 300 2164 304
rect 2158 299 2164 300
rect 2258 303 2264 304
rect 2258 299 2259 303
rect 2263 299 2264 303
rect 2294 300 2295 304
rect 2299 300 2300 304
rect 2294 299 2300 300
rect 2394 303 2400 304
rect 2394 299 2395 303
rect 2399 299 2400 303
rect 2430 300 2431 304
rect 2435 300 2436 304
rect 2430 299 2436 300
rect 2530 303 2536 304
rect 2530 299 2531 303
rect 2535 299 2536 303
rect 2566 300 2567 304
rect 2571 300 2572 304
rect 2566 299 2572 300
rect 2666 303 2672 304
rect 2666 299 2667 303
rect 2671 299 2672 303
rect 2702 300 2703 304
rect 2707 300 2708 304
rect 2702 299 2708 300
rect 2794 303 2800 304
rect 2794 299 2795 303
rect 2799 299 2800 303
rect 2838 300 2839 304
rect 2843 300 2844 304
rect 2838 299 2844 300
rect 2122 298 2128 299
rect 2258 298 2264 299
rect 2394 298 2400 299
rect 2530 298 2536 299
rect 2666 298 2672 299
rect 2794 298 2800 299
rect 1994 289 2000 290
rect 1974 288 1980 289
rect 1974 284 1975 288
rect 1979 284 1980 288
rect 1994 285 1995 289
rect 1999 285 2000 289
rect 1994 284 2000 285
rect 1974 283 1980 284
rect 403 206 407 207
rect 403 201 407 202
rect 475 206 479 207
rect 475 201 479 202
rect 539 206 543 207
rect 539 201 543 202
rect 667 206 671 207
rect 667 201 671 202
rect 675 206 679 207
rect 675 201 679 202
rect 811 206 815 207
rect 811 201 815 202
rect 859 206 863 207
rect 859 201 863 202
rect 947 206 951 207
rect 947 201 951 202
rect 1051 206 1055 207
rect 1051 201 1055 202
rect 1083 206 1087 207
rect 1083 201 1087 202
rect 1935 206 1939 207
rect 1935 201 1939 202
rect 404 140 406 201
rect 522 199 528 200
rect 522 195 523 199
rect 527 195 528 199
rect 522 194 528 195
rect 498 187 504 188
rect 498 183 499 187
rect 503 183 504 187
rect 498 182 504 183
rect 500 160 502 182
rect 498 159 504 160
rect 498 155 499 159
rect 503 155 504 159
rect 498 154 504 155
rect 402 139 408 140
rect 402 135 403 139
rect 407 135 408 139
rect 402 134 408 135
rect 430 124 436 125
rect 524 124 526 194
rect 540 140 542 201
rect 666 191 672 192
rect 666 187 667 191
rect 671 187 672 191
rect 666 186 672 187
rect 658 159 664 160
rect 658 155 659 159
rect 663 155 664 159
rect 658 154 664 155
rect 538 139 544 140
rect 538 135 539 139
rect 543 135 544 139
rect 538 134 544 135
rect 566 124 572 125
rect 110 123 116 124
rect 110 119 111 123
rect 115 119 116 123
rect 158 120 159 124
rect 163 120 164 124
rect 158 119 164 120
rect 274 123 280 124
rect 274 119 275 123
rect 279 119 280 123
rect 294 120 295 124
rect 299 120 300 124
rect 294 119 300 120
rect 386 123 392 124
rect 386 119 387 123
rect 391 119 392 123
rect 430 120 431 124
rect 435 120 436 124
rect 430 119 436 120
rect 522 123 528 124
rect 522 119 523 123
rect 527 119 528 123
rect 566 120 567 124
rect 571 120 572 124
rect 660 124 662 154
rect 668 132 670 186
rect 676 140 678 201
rect 812 140 814 201
rect 948 140 950 201
rect 954 187 960 188
rect 954 183 955 187
rect 959 183 960 187
rect 954 182 960 183
rect 674 139 680 140
rect 674 135 675 139
rect 679 135 680 139
rect 674 134 680 135
rect 810 139 816 140
rect 810 135 811 139
rect 815 135 816 139
rect 810 134 816 135
rect 946 139 952 140
rect 946 135 947 139
rect 951 135 952 139
rect 946 134 952 135
rect 666 131 672 132
rect 666 127 667 131
rect 671 127 672 131
rect 666 126 672 127
rect 702 124 708 125
rect 660 123 668 124
rect 660 121 663 123
rect 566 119 572 120
rect 662 119 663 121
rect 667 119 668 123
rect 702 120 703 124
rect 707 120 708 124
rect 702 119 708 120
rect 838 124 844 125
rect 956 124 958 182
rect 1084 140 1086 201
rect 1206 199 1212 200
rect 1206 195 1207 199
rect 1211 195 1212 199
rect 1206 194 1212 195
rect 1090 187 1096 188
rect 1090 183 1091 187
rect 1095 183 1096 187
rect 1090 182 1096 183
rect 1082 139 1088 140
rect 1082 135 1083 139
rect 1087 135 1088 139
rect 1082 134 1088 135
rect 974 124 980 125
rect 1092 124 1094 182
rect 1110 124 1116 125
rect 1208 124 1210 194
rect 1936 141 1938 201
rect 1976 191 1978 283
rect 1996 191 1998 284
rect 2090 283 2096 284
rect 2090 279 2091 283
rect 2095 279 2096 283
rect 2090 278 2096 279
rect 2092 240 2094 278
rect 2115 252 2119 253
rect 2115 247 2119 248
rect 2090 239 2096 240
rect 2090 235 2091 239
rect 2095 235 2096 239
rect 2090 234 2096 235
rect 1975 190 1979 191
rect 1975 185 1979 186
rect 1995 190 1999 191
rect 1995 185 1999 186
rect 1934 140 1940 141
rect 1934 136 1935 140
rect 1939 136 1940 140
rect 1934 135 1940 136
rect 1976 125 1978 185
rect 1974 124 1980 125
rect 1996 124 1998 185
rect 2116 176 2118 247
rect 2124 240 2126 298
rect 2130 289 2136 290
rect 2130 285 2131 289
rect 2135 285 2136 289
rect 2130 284 2136 285
rect 2122 239 2128 240
rect 2122 235 2123 239
rect 2127 235 2128 239
rect 2122 234 2128 235
rect 2132 191 2134 284
rect 2260 240 2262 298
rect 2266 289 2272 290
rect 2266 285 2267 289
rect 2271 285 2272 289
rect 2266 284 2272 285
rect 2258 239 2264 240
rect 2258 235 2259 239
rect 2263 235 2264 239
rect 2258 234 2264 235
rect 2268 191 2270 284
rect 2396 240 2398 298
rect 2402 289 2408 290
rect 2402 285 2403 289
rect 2407 285 2408 289
rect 2402 284 2408 285
rect 2394 239 2400 240
rect 2394 235 2395 239
rect 2399 235 2400 239
rect 2394 234 2400 235
rect 2404 191 2406 284
rect 2532 240 2534 298
rect 2538 289 2544 290
rect 2538 285 2539 289
rect 2543 285 2544 289
rect 2538 284 2544 285
rect 2530 239 2536 240
rect 2530 235 2531 239
rect 2535 235 2536 239
rect 2530 234 2536 235
rect 2540 191 2542 284
rect 2668 240 2670 298
rect 2674 289 2680 290
rect 2674 285 2675 289
rect 2679 285 2680 289
rect 2674 284 2680 285
rect 2666 239 2672 240
rect 2666 235 2667 239
rect 2671 235 2672 239
rect 2666 234 2672 235
rect 2676 191 2678 284
rect 2796 253 2798 298
rect 2810 289 2816 290
rect 2810 285 2811 289
rect 2815 285 2816 289
rect 2810 284 2816 285
rect 2860 284 2862 382
rect 2960 335 2962 383
rect 2959 334 2963 335
rect 2959 329 2963 330
rect 2975 334 2979 335
rect 2975 329 2979 330
rect 2976 305 2978 329
rect 3016 320 3018 450
rect 3132 404 3134 465
rect 3138 451 3144 452
rect 3138 447 3139 451
rect 3143 447 3144 451
rect 3138 446 3144 447
rect 3130 403 3136 404
rect 3130 399 3131 403
rect 3135 399 3136 403
rect 3130 398 3136 399
rect 3140 388 3142 446
rect 3332 404 3334 465
rect 3338 451 3344 452
rect 3338 447 3339 451
rect 3343 447 3344 451
rect 3338 446 3344 447
rect 3330 403 3336 404
rect 3330 399 3331 403
rect 3335 399 3336 403
rect 3330 398 3336 399
rect 3158 388 3164 389
rect 3340 388 3342 446
rect 3532 404 3534 465
rect 3538 451 3544 452
rect 3538 447 3539 451
rect 3543 447 3544 451
rect 3538 446 3544 447
rect 3530 403 3536 404
rect 3530 399 3531 403
rect 3535 399 3536 403
rect 3530 398 3536 399
rect 3358 388 3364 389
rect 3540 388 3542 446
rect 3558 388 3564 389
rect 3660 388 3662 494
rect 3800 471 3802 551
rect 3840 487 3842 563
rect 3860 487 3862 564
rect 4014 519 4020 520
rect 4014 515 4015 519
rect 4019 515 4020 519
rect 4014 514 4020 515
rect 3839 486 3843 487
rect 3839 481 3843 482
rect 3859 486 3863 487
rect 3859 481 3863 482
rect 3891 486 3895 487
rect 3891 481 3895 482
rect 3799 470 3803 471
rect 3799 465 3803 466
rect 3800 405 3802 465
rect 3840 421 3842 481
rect 3838 420 3844 421
rect 3892 420 3894 481
rect 3838 416 3839 420
rect 3843 416 3844 420
rect 3838 415 3844 416
rect 3890 419 3896 420
rect 3890 415 3891 419
rect 3895 415 3896 419
rect 3890 414 3896 415
rect 3798 404 3804 405
rect 3918 404 3924 405
rect 4016 404 4018 514
rect 4116 487 4118 564
rect 4240 512 4242 578
rect 4378 569 4384 570
rect 4378 565 4379 569
rect 4383 565 4384 569
rect 4378 564 4384 565
rect 4238 511 4244 512
rect 4238 507 4239 511
rect 4243 507 4244 511
rect 4238 506 4244 507
rect 4380 487 4382 564
rect 4448 520 4450 646
rect 4584 615 4586 647
rect 4678 646 4684 647
rect 4808 615 4810 647
rect 5010 646 5016 647
rect 5032 615 5034 647
rect 5234 646 5240 647
rect 5256 615 5258 647
rect 5346 646 5352 647
rect 4583 614 4587 615
rect 4583 609 4587 610
rect 4647 614 4651 615
rect 4647 609 4651 610
rect 4807 614 4811 615
rect 4807 609 4811 610
rect 4879 614 4883 615
rect 4879 609 4883 610
rect 5031 614 5035 615
rect 5031 609 5035 610
rect 5095 614 5099 615
rect 5095 609 5099 610
rect 5255 614 5259 615
rect 5255 609 5259 610
rect 5311 614 5315 615
rect 5311 609 5315 610
rect 4648 585 4650 609
rect 4880 585 4882 609
rect 5096 585 5098 609
rect 5312 585 5314 609
rect 4646 584 4652 585
rect 4878 584 4884 585
rect 5094 584 5100 585
rect 5310 584 5316 585
rect 4502 583 4508 584
rect 4502 579 4503 583
rect 4507 579 4508 583
rect 4646 580 4647 584
rect 4651 580 4652 584
rect 4646 579 4652 580
rect 4766 583 4772 584
rect 4766 579 4767 583
rect 4771 579 4772 583
rect 4878 580 4879 584
rect 4883 580 4884 584
rect 4878 579 4884 580
rect 4978 583 4984 584
rect 4978 579 4979 583
rect 4983 579 4984 583
rect 5094 580 5095 584
rect 5099 580 5100 584
rect 5094 579 5100 580
rect 5194 583 5200 584
rect 5194 579 5195 583
rect 5199 579 5200 583
rect 5310 580 5311 584
rect 5315 580 5316 584
rect 5310 579 5316 580
rect 4502 578 4508 579
rect 4766 578 4772 579
rect 4978 578 4984 579
rect 5194 578 5200 579
rect 4446 519 4452 520
rect 4446 515 4447 519
rect 4451 515 4452 519
rect 4446 514 4452 515
rect 4115 486 4119 487
rect 4115 481 4119 482
rect 4171 486 4175 487
rect 4171 481 4175 482
rect 4379 486 4383 487
rect 4379 481 4383 482
rect 4435 486 4439 487
rect 4435 481 4439 482
rect 4162 471 4168 472
rect 4162 467 4163 471
rect 4167 467 4168 471
rect 4162 466 4168 467
rect 4164 412 4166 466
rect 4172 420 4174 481
rect 4294 471 4300 472
rect 4294 467 4295 471
rect 4299 467 4300 471
rect 4294 466 4300 467
rect 4170 419 4176 420
rect 4170 415 4171 419
rect 4175 415 4176 419
rect 4170 414 4176 415
rect 4162 411 4168 412
rect 4162 407 4163 411
rect 4167 407 4168 411
rect 4162 406 4168 407
rect 4198 404 4204 405
rect 3798 400 3799 404
rect 3803 400 3804 404
rect 3798 399 3804 400
rect 3838 403 3844 404
rect 3838 399 3839 403
rect 3843 399 3844 403
rect 3918 400 3919 404
rect 3923 400 3924 404
rect 3918 399 3924 400
rect 4014 403 4020 404
rect 4014 399 4015 403
rect 4019 399 4020 403
rect 4198 400 4199 404
rect 4203 400 4204 404
rect 4198 399 4204 400
rect 3838 398 3844 399
rect 3138 387 3144 388
rect 3138 383 3139 387
rect 3143 383 3144 387
rect 3158 384 3159 388
rect 3163 384 3164 388
rect 3158 383 3164 384
rect 3338 387 3344 388
rect 3338 383 3339 387
rect 3343 383 3344 387
rect 3358 384 3359 388
rect 3363 384 3364 388
rect 3358 383 3364 384
rect 3538 387 3544 388
rect 3538 383 3539 387
rect 3543 383 3544 387
rect 3558 384 3559 388
rect 3563 384 3564 388
rect 3558 383 3564 384
rect 3658 387 3664 388
rect 3658 383 3659 387
rect 3663 383 3664 387
rect 3138 382 3144 383
rect 3160 335 3162 383
rect 3338 382 3344 383
rect 3360 335 3362 383
rect 3538 382 3544 383
rect 3560 335 3562 383
rect 3658 382 3664 383
rect 3798 387 3804 388
rect 3798 383 3799 387
rect 3803 383 3804 387
rect 3798 382 3804 383
rect 3800 335 3802 382
rect 3840 371 3842 398
rect 3920 371 3922 399
rect 4014 398 4020 399
rect 4200 371 4202 399
rect 3839 370 3843 371
rect 3839 365 3843 366
rect 3919 370 3923 371
rect 3919 365 3923 366
rect 4007 370 4011 371
rect 4007 365 4011 366
rect 4199 370 4203 371
rect 4199 365 4203 366
rect 3840 342 3842 365
rect 3838 341 3844 342
rect 4008 341 4010 365
rect 4200 341 4202 365
rect 3838 337 3839 341
rect 3843 337 3844 341
rect 3838 336 3844 337
rect 4006 340 4012 341
rect 4198 340 4204 341
rect 4296 340 4298 466
rect 4436 420 4438 481
rect 4504 472 4506 578
rect 4618 569 4624 570
rect 4618 565 4619 569
rect 4623 565 4624 569
rect 4618 564 4624 565
rect 4620 487 4622 564
rect 4714 555 4720 556
rect 4714 551 4715 555
rect 4719 551 4720 555
rect 4714 550 4720 551
rect 4716 520 4718 550
rect 4768 520 4770 578
rect 4850 569 4856 570
rect 4850 565 4851 569
rect 4855 565 4856 569
rect 4850 564 4856 565
rect 4778 547 4784 548
rect 4778 543 4779 547
rect 4783 543 4784 547
rect 4778 542 4784 543
rect 4714 519 4720 520
rect 4714 515 4715 519
rect 4719 515 4720 519
rect 4714 514 4720 515
rect 4766 519 4772 520
rect 4766 515 4767 519
rect 4771 515 4772 519
rect 4766 514 4772 515
rect 4619 486 4623 487
rect 4619 481 4623 482
rect 4683 486 4687 487
rect 4683 481 4687 482
rect 4502 471 4508 472
rect 4502 467 4503 471
rect 4507 467 4508 471
rect 4502 466 4508 467
rect 4684 420 4686 481
rect 4780 472 4782 542
rect 4852 487 4854 564
rect 4980 520 4982 578
rect 5066 569 5072 570
rect 5066 565 5067 569
rect 5071 565 5072 569
rect 5066 564 5072 565
rect 4978 519 4984 520
rect 4978 515 4979 519
rect 4983 515 4984 519
rect 4978 514 4984 515
rect 5068 487 5070 564
rect 5196 520 5198 578
rect 5282 569 5288 570
rect 5282 565 5283 569
rect 5287 565 5288 569
rect 5282 564 5288 565
rect 5194 519 5200 520
rect 5194 515 5195 519
rect 5199 515 5200 519
rect 5194 514 5200 515
rect 5284 487 5286 564
rect 5348 556 5350 646
rect 5488 615 5490 647
rect 5582 646 5588 647
rect 5487 614 5491 615
rect 5487 609 5491 610
rect 5527 614 5531 615
rect 5527 609 5531 610
rect 5528 585 5530 609
rect 5526 584 5532 585
rect 5402 583 5408 584
rect 5402 579 5403 583
rect 5407 579 5408 583
rect 5526 580 5527 584
rect 5531 580 5532 584
rect 5526 579 5532 580
rect 5402 578 5408 579
rect 5346 555 5352 556
rect 5346 551 5347 555
rect 5351 551 5352 555
rect 5346 550 5352 551
rect 5404 548 5406 578
rect 5498 569 5504 570
rect 5498 565 5499 569
rect 5503 565 5504 569
rect 5498 564 5504 565
rect 5402 547 5408 548
rect 5402 543 5403 547
rect 5407 543 5408 547
rect 5402 542 5408 543
rect 5500 487 5502 564
rect 5584 520 5586 646
rect 5622 583 5628 584
rect 5622 579 5623 583
rect 5627 579 5628 583
rect 5622 578 5628 579
rect 5582 519 5588 520
rect 5582 515 5583 519
rect 5587 515 5588 519
rect 5582 514 5588 515
rect 4851 486 4855 487
rect 4851 481 4855 482
rect 4907 486 4911 487
rect 4907 481 4911 482
rect 5067 486 5071 487
rect 5067 481 5071 482
rect 5123 486 5127 487
rect 5123 481 5127 482
rect 5283 486 5287 487
rect 5283 481 5287 482
rect 5331 486 5335 487
rect 5331 481 5335 482
rect 5499 486 5503 487
rect 5499 481 5503 482
rect 5515 486 5519 487
rect 5515 481 5519 482
rect 4778 471 4784 472
rect 4778 467 4779 471
rect 4783 467 4784 471
rect 4778 466 4784 467
rect 4908 420 4910 481
rect 4914 467 4920 468
rect 4914 463 4915 467
rect 4919 463 4920 467
rect 4914 462 4920 463
rect 4434 419 4440 420
rect 4434 415 4435 419
rect 4439 415 4440 419
rect 4434 414 4440 415
rect 4682 419 4688 420
rect 4682 415 4683 419
rect 4687 415 4688 419
rect 4682 414 4688 415
rect 4906 419 4912 420
rect 4906 415 4907 419
rect 4911 415 4912 419
rect 4906 414 4912 415
rect 4462 404 4468 405
rect 4710 404 4716 405
rect 4916 404 4918 462
rect 5124 420 5126 481
rect 5130 467 5136 468
rect 5130 463 5131 467
rect 5135 463 5136 467
rect 5130 462 5136 463
rect 5122 419 5128 420
rect 5122 415 5123 419
rect 5127 415 5128 419
rect 5122 414 5128 415
rect 4934 404 4940 405
rect 5132 404 5134 462
rect 5332 420 5334 481
rect 5338 467 5344 468
rect 5338 463 5339 467
rect 5343 463 5344 467
rect 5338 462 5344 463
rect 5330 419 5336 420
rect 5330 415 5331 419
rect 5335 415 5336 419
rect 5330 414 5336 415
rect 5150 404 5156 405
rect 5340 404 5342 462
rect 5516 420 5518 481
rect 5522 467 5528 468
rect 5522 463 5523 467
rect 5527 463 5528 467
rect 5522 462 5528 463
rect 5514 419 5520 420
rect 5514 415 5515 419
rect 5519 415 5520 419
rect 5514 414 5520 415
rect 5358 404 5364 405
rect 5524 404 5526 462
rect 5542 404 5548 405
rect 4462 400 4463 404
rect 4467 400 4468 404
rect 4462 399 4468 400
rect 4554 403 4560 404
rect 4554 399 4555 403
rect 4559 399 4560 403
rect 4710 400 4711 404
rect 4715 400 4716 404
rect 4710 399 4716 400
rect 4914 403 4920 404
rect 4914 399 4915 403
rect 4919 399 4920 403
rect 4934 400 4935 404
rect 4939 400 4940 404
rect 4934 399 4940 400
rect 5130 403 5136 404
rect 5130 399 5131 403
rect 5135 399 5136 403
rect 5150 400 5151 404
rect 5155 400 5156 404
rect 5150 399 5156 400
rect 5338 403 5344 404
rect 5338 399 5339 403
rect 5343 399 5344 403
rect 5358 400 5359 404
rect 5363 400 5364 404
rect 5358 399 5364 400
rect 5522 403 5528 404
rect 5522 399 5523 403
rect 5527 399 5528 403
rect 5542 400 5543 404
rect 5547 400 5548 404
rect 5542 399 5548 400
rect 4464 371 4466 399
rect 4554 398 4560 399
rect 4423 370 4427 371
rect 4423 365 4427 366
rect 4463 370 4467 371
rect 4463 365 4467 366
rect 4424 341 4426 365
rect 4556 347 4558 398
rect 4712 371 4714 399
rect 4914 398 4920 399
rect 4936 371 4938 399
rect 5130 398 5136 399
rect 5152 371 5154 399
rect 5338 398 5344 399
rect 5360 371 5362 399
rect 5522 398 5528 399
rect 5544 371 5546 399
rect 4679 370 4683 371
rect 4679 365 4683 366
rect 4711 370 4715 371
rect 4711 365 4715 366
rect 4935 370 4939 371
rect 4935 365 4939 366
rect 4967 370 4971 371
rect 4967 365 4971 366
rect 5151 370 5155 371
rect 5151 365 5155 366
rect 5263 370 5267 371
rect 5263 365 5267 366
rect 5359 370 5363 371
rect 5359 365 5363 366
rect 5543 370 5547 371
rect 5543 365 5547 366
rect 4552 345 4558 347
rect 4422 340 4428 341
rect 4006 336 4007 340
rect 4011 336 4012 340
rect 4006 335 4012 336
rect 4134 339 4140 340
rect 4134 335 4135 339
rect 4139 335 4140 339
rect 4198 336 4199 340
rect 4203 336 4204 340
rect 4198 335 4204 336
rect 4294 339 4300 340
rect 4294 335 4295 339
rect 4299 335 4300 339
rect 4422 336 4423 340
rect 4427 336 4428 340
rect 4422 335 4428 336
rect 3111 334 3115 335
rect 3111 329 3115 330
rect 3159 334 3163 335
rect 3159 329 3163 330
rect 3247 334 3251 335
rect 3247 329 3251 330
rect 3359 334 3363 335
rect 3359 329 3363 330
rect 3383 334 3387 335
rect 3383 329 3387 330
rect 3519 334 3523 335
rect 3519 329 3523 330
rect 3559 334 3563 335
rect 3559 329 3563 330
rect 3799 334 3803 335
rect 4134 334 4140 335
rect 4294 334 4300 335
rect 3799 329 3803 330
rect 3014 319 3020 320
rect 3014 315 3015 319
rect 3019 315 3020 319
rect 3014 314 3020 315
rect 3112 305 3114 329
rect 3248 305 3250 329
rect 3384 305 3386 329
rect 3520 305 3522 329
rect 3800 306 3802 329
rect 3978 325 3984 326
rect 3838 324 3844 325
rect 3838 320 3839 324
rect 3843 320 3844 324
rect 3978 321 3979 325
rect 3983 321 3984 325
rect 3978 320 3984 321
rect 3838 319 3844 320
rect 3798 305 3804 306
rect 2974 304 2980 305
rect 3110 304 3116 305
rect 3246 304 3252 305
rect 3382 304 3388 305
rect 3518 304 3524 305
rect 2938 303 2944 304
rect 2938 299 2939 303
rect 2943 299 2944 303
rect 2974 300 2975 304
rect 2979 300 2980 304
rect 2974 299 2980 300
rect 3074 303 3080 304
rect 3074 299 3075 303
rect 3079 299 3080 303
rect 3110 300 3111 304
rect 3115 300 3116 304
rect 3110 299 3116 300
rect 3210 303 3216 304
rect 3210 299 3211 303
rect 3215 299 3216 303
rect 3246 300 3247 304
rect 3251 300 3252 304
rect 3246 299 3252 300
rect 3346 303 3352 304
rect 3346 299 3347 303
rect 3351 299 3352 303
rect 3382 300 3383 304
rect 3387 300 3388 304
rect 3382 299 3388 300
rect 3482 303 3488 304
rect 3482 299 3483 303
rect 3487 299 3488 303
rect 3518 300 3519 304
rect 3523 300 3524 304
rect 3798 301 3799 305
rect 3803 301 3804 305
rect 3798 300 3804 301
rect 3518 299 3524 300
rect 2938 298 2944 299
rect 3074 298 3080 299
rect 3210 298 3216 299
rect 3346 298 3352 299
rect 3482 298 3488 299
rect 2795 252 2799 253
rect 2795 247 2799 248
rect 2812 191 2814 284
rect 2858 283 2864 284
rect 2858 279 2859 283
rect 2863 279 2864 283
rect 2858 278 2864 279
rect 2940 240 2942 298
rect 2946 289 2952 290
rect 2946 285 2947 289
rect 2951 285 2952 289
rect 2946 284 2952 285
rect 2906 239 2912 240
rect 2906 235 2907 239
rect 2911 235 2912 239
rect 2906 234 2912 235
rect 2938 239 2944 240
rect 2938 235 2939 239
rect 2943 235 2944 239
rect 2938 234 2944 235
rect 2131 190 2135 191
rect 2131 185 2135 186
rect 2267 190 2271 191
rect 2267 185 2271 186
rect 2403 190 2407 191
rect 2403 185 2407 186
rect 2539 190 2543 191
rect 2539 185 2543 186
rect 2675 190 2679 191
rect 2675 185 2679 186
rect 2811 190 2815 191
rect 2811 185 2815 186
rect 2114 175 2120 176
rect 2114 171 2115 175
rect 2119 171 2120 175
rect 2114 170 2120 171
rect 2132 124 2134 185
rect 2138 171 2144 172
rect 2138 167 2139 171
rect 2143 167 2144 171
rect 2138 166 2144 167
rect 838 120 839 124
rect 843 120 844 124
rect 838 119 844 120
rect 954 123 960 124
rect 954 119 955 123
rect 959 119 960 123
rect 974 120 975 124
rect 979 120 980 124
rect 974 119 980 120
rect 1090 123 1096 124
rect 1090 119 1091 123
rect 1095 119 1096 123
rect 1110 120 1111 124
rect 1115 120 1116 124
rect 1110 119 1116 120
rect 1206 123 1212 124
rect 1206 119 1207 123
rect 1211 119 1212 123
rect 110 118 116 119
rect 112 95 114 118
rect 160 95 162 119
rect 274 118 280 119
rect 296 95 298 119
rect 386 118 392 119
rect 432 95 434 119
rect 522 118 528 119
rect 568 95 570 119
rect 662 118 668 119
rect 704 95 706 119
rect 840 95 842 119
rect 954 118 960 119
rect 976 95 978 119
rect 1090 118 1096 119
rect 1112 95 1114 119
rect 1206 118 1212 119
rect 1934 123 1940 124
rect 1934 119 1935 123
rect 1939 119 1940 123
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 1994 123 2000 124
rect 1994 119 1995 123
rect 1999 119 2000 123
rect 1934 118 1940 119
rect 1994 118 2000 119
rect 2130 123 2136 124
rect 2130 119 2131 123
rect 2135 119 2136 123
rect 2130 118 2136 119
rect 1936 95 1938 118
rect 2022 108 2028 109
rect 2140 108 2142 166
rect 2268 124 2270 185
rect 2274 171 2280 172
rect 2274 167 2275 171
rect 2279 167 2280 171
rect 2274 166 2280 167
rect 2266 123 2272 124
rect 2266 119 2267 123
rect 2271 119 2272 123
rect 2266 118 2272 119
rect 2158 108 2164 109
rect 2276 108 2278 166
rect 2404 124 2406 185
rect 2410 171 2416 172
rect 2410 167 2411 171
rect 2415 167 2416 171
rect 2410 166 2416 167
rect 2402 123 2408 124
rect 2402 119 2403 123
rect 2407 119 2408 123
rect 2402 118 2408 119
rect 2294 108 2300 109
rect 2412 108 2414 166
rect 2540 124 2542 185
rect 2546 171 2552 172
rect 2546 167 2547 171
rect 2551 167 2552 171
rect 2546 166 2552 167
rect 2538 123 2544 124
rect 2538 119 2539 123
rect 2543 119 2544 123
rect 2538 118 2544 119
rect 2430 108 2436 109
rect 2548 108 2550 166
rect 2676 124 2678 185
rect 2682 171 2688 172
rect 2682 167 2683 171
rect 2687 167 2688 171
rect 2682 166 2688 167
rect 2674 123 2680 124
rect 2674 119 2675 123
rect 2679 119 2680 123
rect 2674 118 2680 119
rect 2566 108 2572 109
rect 2684 108 2686 166
rect 2812 124 2814 185
rect 2908 181 2910 234
rect 2948 191 2950 284
rect 3076 240 3078 298
rect 3082 289 3088 290
rect 3082 285 3083 289
rect 3087 285 3088 289
rect 3082 284 3088 285
rect 3074 239 3080 240
rect 3074 235 3075 239
rect 3079 235 3080 239
rect 3074 234 3080 235
rect 3084 191 3086 284
rect 3212 240 3214 298
rect 3218 289 3224 290
rect 3218 285 3219 289
rect 3223 285 3224 289
rect 3218 284 3224 285
rect 3210 239 3216 240
rect 3210 235 3211 239
rect 3215 235 3216 239
rect 3210 234 3216 235
rect 3220 191 3222 284
rect 3348 240 3350 298
rect 3354 289 3360 290
rect 3354 285 3355 289
rect 3359 285 3360 289
rect 3354 284 3360 285
rect 3346 239 3352 240
rect 3346 235 3347 239
rect 3351 235 3352 239
rect 3346 234 3352 235
rect 3356 191 3358 284
rect 3484 240 3486 298
rect 3490 289 3496 290
rect 3490 285 3491 289
rect 3495 285 3496 289
rect 3490 284 3496 285
rect 3798 288 3804 289
rect 3798 284 3799 288
rect 3803 284 3804 288
rect 3482 239 3488 240
rect 3482 235 3483 239
rect 3487 235 3488 239
rect 3482 234 3488 235
rect 3492 191 3494 284
rect 3798 283 3804 284
rect 3800 191 3802 283
rect 3840 207 3842 319
rect 3980 207 3982 320
rect 4136 276 4138 334
rect 4170 325 4176 326
rect 4170 321 4171 325
rect 4175 321 4176 325
rect 4170 320 4176 321
rect 4394 325 4400 326
rect 4394 321 4395 325
rect 4399 321 4400 325
rect 4394 320 4400 321
rect 4114 275 4120 276
rect 4114 271 4115 275
rect 4119 271 4120 275
rect 4114 270 4120 271
rect 4134 275 4140 276
rect 4134 271 4135 275
rect 4139 271 4140 275
rect 4134 270 4140 271
rect 3839 206 3843 207
rect 3839 201 3843 202
rect 3859 206 3863 207
rect 3859 201 3863 202
rect 3979 206 3983 207
rect 3979 201 3983 202
rect 3995 206 3999 207
rect 3995 201 3999 202
rect 2947 190 2951 191
rect 2947 185 2951 186
rect 3083 190 3087 191
rect 3083 185 3087 186
rect 3219 190 3223 191
rect 3219 185 3223 186
rect 3355 190 3359 191
rect 3355 185 3359 186
rect 3491 190 3495 191
rect 3491 185 3495 186
rect 3627 190 3631 191
rect 3627 185 3631 186
rect 3799 190 3803 191
rect 3799 185 3803 186
rect 2907 180 2911 181
rect 2907 175 2911 176
rect 2818 171 2824 172
rect 2818 167 2819 171
rect 2823 167 2824 171
rect 2818 166 2824 167
rect 2810 123 2816 124
rect 2810 119 2811 123
rect 2815 119 2816 123
rect 2810 118 2816 119
rect 2702 108 2708 109
rect 2820 108 2822 166
rect 2948 124 2950 185
rect 2954 171 2960 172
rect 2954 167 2955 171
rect 2959 167 2960 171
rect 2954 166 2960 167
rect 2946 123 2952 124
rect 2946 119 2947 123
rect 2951 119 2952 123
rect 2946 118 2952 119
rect 2838 108 2844 109
rect 2956 108 2958 166
rect 3084 124 3086 185
rect 3090 171 3096 172
rect 3090 167 3091 171
rect 3095 167 3096 171
rect 3090 166 3096 167
rect 3082 123 3088 124
rect 3082 119 3083 123
rect 3087 119 3088 123
rect 3082 118 3088 119
rect 2974 108 2980 109
rect 3092 108 3094 166
rect 3220 124 3222 185
rect 3226 171 3232 172
rect 3226 167 3227 171
rect 3231 167 3232 171
rect 3226 166 3232 167
rect 3218 123 3224 124
rect 3218 119 3219 123
rect 3223 119 3224 123
rect 3218 118 3224 119
rect 3110 108 3116 109
rect 3228 108 3230 166
rect 3356 124 3358 185
rect 3362 171 3368 172
rect 3362 167 3363 171
rect 3367 167 3368 171
rect 3362 166 3368 167
rect 3354 123 3360 124
rect 3354 119 3355 123
rect 3359 119 3360 123
rect 3354 118 3360 119
rect 3246 108 3252 109
rect 3364 108 3366 166
rect 3492 124 3494 185
rect 3498 171 3504 172
rect 3498 167 3499 171
rect 3503 167 3504 171
rect 3498 166 3504 167
rect 3490 123 3496 124
rect 3490 119 3491 123
rect 3495 119 3496 123
rect 3490 118 3496 119
rect 3382 108 3388 109
rect 3500 108 3502 166
rect 3628 124 3630 185
rect 3751 180 3755 181
rect 3751 175 3755 176
rect 3634 171 3640 172
rect 3634 167 3635 171
rect 3639 167 3640 171
rect 3634 166 3640 167
rect 3626 123 3632 124
rect 3626 119 3627 123
rect 3631 119 3632 123
rect 3626 118 3632 119
rect 3518 108 3524 109
rect 3636 108 3638 166
rect 3654 108 3660 109
rect 3752 108 3754 175
rect 3800 125 3802 185
rect 3840 141 3842 201
rect 3838 140 3844 141
rect 3860 140 3862 201
rect 3996 140 3998 201
rect 4002 187 4008 188
rect 4002 183 4003 187
rect 4007 183 4008 187
rect 4002 182 4008 183
rect 3838 136 3839 140
rect 3843 136 3844 140
rect 3838 135 3844 136
rect 3858 139 3864 140
rect 3858 135 3859 139
rect 3863 135 3864 139
rect 3858 134 3864 135
rect 3994 139 4000 140
rect 3994 135 3995 139
rect 3999 135 4000 139
rect 3994 134 4000 135
rect 3798 124 3804 125
rect 3886 124 3892 125
rect 4004 124 4006 182
rect 4022 124 4028 125
rect 4116 124 4118 270
rect 4172 207 4174 320
rect 4396 207 4398 320
rect 4552 276 4554 345
rect 4680 341 4682 365
rect 4968 341 4970 365
rect 5264 341 5266 365
rect 5544 341 5546 365
rect 4678 340 4684 341
rect 4966 340 4972 341
rect 5262 340 5268 341
rect 5542 340 5548 341
rect 4558 339 4564 340
rect 4558 335 4559 339
rect 4563 335 4564 339
rect 4678 336 4679 340
rect 4683 336 4684 340
rect 4678 335 4684 336
rect 4778 339 4784 340
rect 4778 335 4779 339
rect 4783 335 4784 339
rect 4966 336 4967 340
rect 4971 336 4972 340
rect 4966 335 4972 336
rect 5066 339 5072 340
rect 5066 335 5067 339
rect 5071 335 5072 339
rect 5262 336 5263 340
rect 5267 336 5268 340
rect 5262 335 5268 336
rect 5354 339 5360 340
rect 5354 335 5355 339
rect 5359 335 5360 339
rect 5542 336 5543 340
rect 5547 336 5548 340
rect 5542 335 5548 336
rect 4558 334 4564 335
rect 4778 334 4784 335
rect 5066 334 5072 335
rect 5354 334 5360 335
rect 4560 276 4562 334
rect 4650 325 4656 326
rect 4650 321 4651 325
rect 4655 321 4656 325
rect 4650 320 4656 321
rect 4550 275 4556 276
rect 4550 271 4551 275
rect 4555 271 4556 275
rect 4550 270 4556 271
rect 4558 275 4564 276
rect 4558 271 4559 275
rect 4563 271 4564 275
rect 4558 270 4564 271
rect 4652 207 4654 320
rect 4780 276 4782 334
rect 4938 325 4944 326
rect 4938 321 4939 325
rect 4943 321 4944 325
rect 4938 320 4944 321
rect 4778 275 4784 276
rect 4778 271 4779 275
rect 4783 271 4784 275
rect 4778 270 4784 271
rect 4722 255 4728 256
rect 4722 251 4723 255
rect 4727 251 4728 255
rect 4722 250 4728 251
rect 4131 206 4135 207
rect 4131 201 4135 202
rect 4171 206 4175 207
rect 4171 201 4175 202
rect 4267 206 4271 207
rect 4267 201 4271 202
rect 4395 206 4399 207
rect 4395 201 4399 202
rect 4435 206 4439 207
rect 4435 201 4439 202
rect 4627 206 4631 207
rect 4627 201 4631 202
rect 4651 206 4655 207
rect 4651 201 4655 202
rect 4132 140 4134 201
rect 4250 199 4256 200
rect 4250 195 4251 199
rect 4255 195 4256 199
rect 4250 194 4256 195
rect 4226 187 4232 188
rect 4226 183 4227 187
rect 4231 183 4232 187
rect 4226 182 4232 183
rect 4228 160 4230 182
rect 4226 159 4232 160
rect 4226 155 4227 159
rect 4231 155 4232 159
rect 4226 154 4232 155
rect 4130 139 4136 140
rect 4130 135 4131 139
rect 4135 135 4136 139
rect 4130 134 4136 135
rect 4158 124 4164 125
rect 4252 124 4254 194
rect 4268 140 4270 201
rect 4394 191 4400 192
rect 4394 187 4395 191
rect 4399 187 4400 191
rect 4394 186 4400 187
rect 4386 159 4392 160
rect 4386 155 4387 159
rect 4391 155 4392 159
rect 4386 154 4392 155
rect 4266 139 4272 140
rect 4266 135 4267 139
rect 4271 135 4272 139
rect 4266 134 4272 135
rect 4294 124 4300 125
rect 3798 120 3799 124
rect 3803 120 3804 124
rect 3798 119 3804 120
rect 3838 123 3844 124
rect 3838 119 3839 123
rect 3843 119 3844 123
rect 3886 120 3887 124
rect 3891 120 3892 124
rect 3886 119 3892 120
rect 4002 123 4008 124
rect 4002 119 4003 123
rect 4007 119 4008 123
rect 4022 120 4023 124
rect 4027 120 4028 124
rect 4022 119 4028 120
rect 4114 123 4120 124
rect 4114 119 4115 123
rect 4119 119 4120 123
rect 4158 120 4159 124
rect 4163 120 4164 124
rect 4158 119 4164 120
rect 4250 123 4256 124
rect 4250 119 4251 123
rect 4255 119 4256 123
rect 4294 120 4295 124
rect 4299 120 4300 124
rect 4388 124 4390 154
rect 4396 132 4398 186
rect 4436 140 4438 201
rect 4530 187 4536 188
rect 4530 183 4531 187
rect 4535 183 4536 187
rect 4530 182 4536 183
rect 4532 156 4534 182
rect 4530 155 4536 156
rect 4530 151 4531 155
rect 4535 151 4536 155
rect 4530 150 4536 151
rect 4628 140 4630 201
rect 4724 192 4726 250
rect 4940 207 4942 320
rect 5068 276 5070 334
rect 5234 325 5240 326
rect 5234 321 5235 325
rect 5239 321 5240 325
rect 5234 320 5240 321
rect 5066 275 5072 276
rect 5066 271 5067 275
rect 5071 271 5072 275
rect 5066 270 5072 271
rect 5236 207 5238 320
rect 5356 256 5358 334
rect 5514 325 5520 326
rect 5514 321 5515 325
rect 5519 321 5520 325
rect 5514 320 5520 321
rect 5354 255 5360 256
rect 5354 251 5355 255
rect 5359 251 5360 255
rect 5354 250 5360 251
rect 5516 207 5518 320
rect 5624 276 5626 578
rect 5640 404 5642 714
rect 5664 669 5666 729
rect 5662 668 5668 669
rect 5662 664 5663 668
rect 5667 664 5668 668
rect 5662 663 5668 664
rect 5662 651 5668 652
rect 5662 647 5663 651
rect 5667 647 5668 651
rect 5662 646 5668 647
rect 5664 615 5666 646
rect 5663 614 5667 615
rect 5663 609 5667 610
rect 5664 586 5666 609
rect 5662 585 5668 586
rect 5662 581 5663 585
rect 5667 581 5668 585
rect 5662 580 5668 581
rect 5662 568 5668 569
rect 5662 564 5663 568
rect 5667 564 5668 568
rect 5662 563 5668 564
rect 5664 487 5666 563
rect 5663 486 5667 487
rect 5663 481 5667 482
rect 5664 421 5666 481
rect 5662 420 5668 421
rect 5662 416 5663 420
rect 5667 416 5668 420
rect 5662 415 5668 416
rect 5638 403 5644 404
rect 5638 399 5639 403
rect 5643 399 5644 403
rect 5638 398 5644 399
rect 5662 403 5668 404
rect 5662 399 5663 403
rect 5667 399 5668 403
rect 5662 398 5668 399
rect 5664 371 5666 398
rect 5663 370 5667 371
rect 5663 365 5667 366
rect 5664 342 5666 365
rect 5662 341 5668 342
rect 5634 339 5640 340
rect 5634 335 5635 339
rect 5639 335 5640 339
rect 5662 337 5663 341
rect 5667 337 5668 341
rect 5662 336 5668 337
rect 5634 334 5640 335
rect 5622 275 5628 276
rect 5622 271 5623 275
rect 5627 271 5628 275
rect 5622 270 5628 271
rect 4843 206 4847 207
rect 4843 201 4847 202
rect 4939 206 4943 207
rect 4939 201 4943 202
rect 5067 206 5071 207
rect 5067 201 5071 202
rect 5235 206 5239 207
rect 5235 201 5239 202
rect 5299 206 5303 207
rect 5299 201 5303 202
rect 5515 206 5519 207
rect 5515 201 5519 202
rect 4722 191 4728 192
rect 4722 187 4723 191
rect 4727 187 4728 191
rect 4722 186 4728 187
rect 4844 140 4846 201
rect 4850 187 4856 188
rect 4850 183 4851 187
rect 4855 183 4856 187
rect 4850 182 4856 183
rect 4434 139 4440 140
rect 4434 135 4435 139
rect 4439 135 4440 139
rect 4434 134 4440 135
rect 4626 139 4632 140
rect 4626 135 4627 139
rect 4631 135 4632 139
rect 4626 134 4632 135
rect 4842 139 4848 140
rect 4842 135 4843 139
rect 4847 135 4848 139
rect 4842 134 4848 135
rect 4394 131 4400 132
rect 4394 127 4395 131
rect 4399 127 4400 131
rect 4394 126 4400 127
rect 4462 124 4468 125
rect 4388 123 4396 124
rect 4388 121 4391 123
rect 4294 119 4300 120
rect 4390 119 4391 121
rect 4395 119 4396 123
rect 4462 120 4463 124
rect 4467 120 4468 124
rect 4462 119 4468 120
rect 4654 124 4660 125
rect 4852 124 4854 182
rect 5068 140 5070 201
rect 5074 187 5080 188
rect 5074 183 5075 187
rect 5079 183 5080 187
rect 5074 182 5080 183
rect 5066 139 5072 140
rect 5066 135 5067 139
rect 5071 135 5072 139
rect 5066 134 5072 135
rect 4870 124 4876 125
rect 5076 124 5078 182
rect 5186 155 5192 156
rect 5186 151 5187 155
rect 5191 151 5192 155
rect 5186 150 5192 151
rect 5094 124 5100 125
rect 5188 124 5190 150
rect 5300 140 5302 201
rect 5502 191 5508 192
rect 5502 187 5503 191
rect 5507 187 5508 191
rect 5502 186 5508 187
rect 5298 139 5304 140
rect 5298 135 5299 139
rect 5303 135 5304 139
rect 5298 134 5304 135
rect 5504 132 5506 186
rect 5516 140 5518 201
rect 5636 192 5638 334
rect 5662 324 5668 325
rect 5662 320 5663 324
rect 5667 320 5668 324
rect 5662 319 5668 320
rect 5664 207 5666 319
rect 5663 206 5667 207
rect 5663 201 5667 202
rect 5634 191 5640 192
rect 5634 187 5635 191
rect 5639 187 5640 191
rect 5634 186 5640 187
rect 5664 141 5666 201
rect 5662 140 5668 141
rect 5514 139 5520 140
rect 5514 135 5515 139
rect 5519 135 5520 139
rect 5662 136 5663 140
rect 5667 136 5668 140
rect 5662 135 5668 136
rect 5514 134 5520 135
rect 5502 131 5508 132
rect 5502 127 5503 131
rect 5507 127 5508 131
rect 5502 126 5508 127
rect 5326 124 5332 125
rect 4654 120 4655 124
rect 4659 120 4660 124
rect 4654 119 4660 120
rect 4850 123 4856 124
rect 4850 119 4851 123
rect 4855 119 4856 123
rect 4870 120 4871 124
rect 4875 120 4876 124
rect 4870 119 4876 120
rect 5074 123 5080 124
rect 5074 119 5075 123
rect 5079 119 5080 123
rect 5094 120 5095 124
rect 5099 120 5100 124
rect 5094 119 5100 120
rect 5186 123 5192 124
rect 5186 119 5187 123
rect 5191 119 5192 123
rect 5326 120 5327 124
rect 5331 120 5332 124
rect 5326 119 5332 120
rect 5542 124 5548 125
rect 5542 120 5543 124
rect 5547 120 5548 124
rect 5542 119 5548 120
rect 5662 123 5668 124
rect 5662 119 5663 123
rect 5667 119 5668 123
rect 3838 118 3844 119
rect 1974 107 1980 108
rect 1974 103 1975 107
rect 1979 103 1980 107
rect 2022 104 2023 108
rect 2027 104 2028 108
rect 2022 103 2028 104
rect 2138 107 2144 108
rect 2138 103 2139 107
rect 2143 103 2144 107
rect 2158 104 2159 108
rect 2163 104 2164 108
rect 2158 103 2164 104
rect 2274 107 2280 108
rect 2274 103 2275 107
rect 2279 103 2280 107
rect 2294 104 2295 108
rect 2299 104 2300 108
rect 2294 103 2300 104
rect 2410 107 2416 108
rect 2410 103 2411 107
rect 2415 103 2416 107
rect 2430 104 2431 108
rect 2435 104 2436 108
rect 2430 103 2436 104
rect 2546 107 2552 108
rect 2546 103 2547 107
rect 2551 103 2552 107
rect 2566 104 2567 108
rect 2571 104 2572 108
rect 2566 103 2572 104
rect 2682 107 2688 108
rect 2682 103 2683 107
rect 2687 103 2688 107
rect 2702 104 2703 108
rect 2707 104 2708 108
rect 2702 103 2708 104
rect 2818 107 2824 108
rect 2818 103 2819 107
rect 2823 103 2824 107
rect 2838 104 2839 108
rect 2843 104 2844 108
rect 2838 103 2844 104
rect 2954 107 2960 108
rect 2954 103 2955 107
rect 2959 103 2960 107
rect 2974 104 2975 108
rect 2979 104 2980 108
rect 2974 103 2980 104
rect 3090 107 3096 108
rect 3090 103 3091 107
rect 3095 103 3096 107
rect 3110 104 3111 108
rect 3115 104 3116 108
rect 3110 103 3116 104
rect 3226 107 3232 108
rect 3226 103 3227 107
rect 3231 103 3232 107
rect 3246 104 3247 108
rect 3251 104 3252 108
rect 3246 103 3252 104
rect 3362 107 3368 108
rect 3362 103 3363 107
rect 3367 103 3368 107
rect 3382 104 3383 108
rect 3387 104 3388 108
rect 3382 103 3388 104
rect 3498 107 3504 108
rect 3498 103 3499 107
rect 3503 103 3504 107
rect 3518 104 3519 108
rect 3523 104 3524 108
rect 3518 103 3524 104
rect 3634 107 3640 108
rect 3634 103 3635 107
rect 3639 103 3640 107
rect 3654 104 3655 108
rect 3659 104 3660 108
rect 3654 103 3660 104
rect 3750 107 3756 108
rect 3750 103 3751 107
rect 3755 103 3756 107
rect 1974 102 1980 103
rect 111 94 115 95
rect 111 89 115 90
rect 159 94 163 95
rect 159 89 163 90
rect 295 94 299 95
rect 295 89 299 90
rect 431 94 435 95
rect 431 89 435 90
rect 567 94 571 95
rect 567 89 571 90
rect 703 94 707 95
rect 703 89 707 90
rect 839 94 843 95
rect 839 89 843 90
rect 975 94 979 95
rect 975 89 979 90
rect 1111 94 1115 95
rect 1111 89 1115 90
rect 1935 94 1939 95
rect 1935 89 1939 90
rect 1976 79 1978 102
rect 2024 79 2026 103
rect 2138 102 2144 103
rect 2160 79 2162 103
rect 2274 102 2280 103
rect 2296 79 2298 103
rect 2410 102 2416 103
rect 2432 79 2434 103
rect 2546 102 2552 103
rect 2568 79 2570 103
rect 2682 102 2688 103
rect 2704 79 2706 103
rect 2818 102 2824 103
rect 2840 79 2842 103
rect 2954 102 2960 103
rect 2976 79 2978 103
rect 3090 102 3096 103
rect 3112 79 3114 103
rect 3226 102 3232 103
rect 3248 79 3250 103
rect 3362 102 3368 103
rect 3384 79 3386 103
rect 3498 102 3504 103
rect 3520 79 3522 103
rect 3634 102 3640 103
rect 3656 79 3658 103
rect 3750 102 3756 103
rect 3798 107 3804 108
rect 3798 103 3799 107
rect 3803 103 3804 107
rect 3798 102 3804 103
rect 3800 79 3802 102
rect 3840 95 3842 118
rect 3888 95 3890 119
rect 4002 118 4008 119
rect 4024 95 4026 119
rect 4114 118 4120 119
rect 4160 95 4162 119
rect 4250 118 4256 119
rect 4296 95 4298 119
rect 4390 118 4396 119
rect 4464 95 4466 119
rect 4656 95 4658 119
rect 4850 118 4856 119
rect 4872 95 4874 119
rect 5074 118 5080 119
rect 5096 95 5098 119
rect 5186 118 5192 119
rect 5328 95 5330 119
rect 5544 95 5546 119
rect 5662 118 5668 119
rect 5664 95 5666 118
rect 3839 94 3843 95
rect 3839 89 3843 90
rect 3887 94 3891 95
rect 3887 89 3891 90
rect 4023 94 4027 95
rect 4023 89 4027 90
rect 4159 94 4163 95
rect 4159 89 4163 90
rect 4295 94 4299 95
rect 4295 89 4299 90
rect 4463 94 4467 95
rect 4463 89 4467 90
rect 4655 94 4659 95
rect 4655 89 4659 90
rect 4871 94 4875 95
rect 4871 89 4875 90
rect 5095 94 5099 95
rect 5095 89 5099 90
rect 5327 94 5331 95
rect 5327 89 5331 90
rect 5543 94 5547 95
rect 5543 89 5547 90
rect 5663 94 5667 95
rect 5663 89 5667 90
rect 1975 78 1979 79
rect 1975 73 1979 74
rect 2023 78 2027 79
rect 2023 73 2027 74
rect 2159 78 2163 79
rect 2159 73 2163 74
rect 2295 78 2299 79
rect 2295 73 2299 74
rect 2431 78 2435 79
rect 2431 73 2435 74
rect 2567 78 2571 79
rect 2567 73 2571 74
rect 2703 78 2707 79
rect 2703 73 2707 74
rect 2839 78 2843 79
rect 2839 73 2843 74
rect 2975 78 2979 79
rect 2975 73 2979 74
rect 3111 78 3115 79
rect 3111 73 3115 74
rect 3247 78 3251 79
rect 3247 73 3251 74
rect 3383 78 3387 79
rect 3383 73 3387 74
rect 3519 78 3523 79
rect 3519 73 3523 74
rect 3655 78 3659 79
rect 3655 73 3659 74
rect 3799 78 3803 79
rect 3799 73 3803 74
<< m4c >>
rect 111 5754 115 5758
rect 131 5754 135 5758
rect 371 5754 375 5758
rect 635 5754 639 5758
rect 907 5754 911 5758
rect 1179 5754 1183 5758
rect 1451 5754 1455 5758
rect 1723 5754 1727 5758
rect 1935 5754 1939 5758
rect 111 5642 115 5646
rect 159 5642 163 5646
rect 399 5642 403 5646
rect 455 5642 459 5646
rect 647 5642 651 5646
rect 663 5642 667 5646
rect 855 5642 859 5646
rect 935 5642 939 5646
rect 883 5560 887 5564
rect 111 5530 115 5534
rect 427 5530 431 5534
rect 619 5530 623 5534
rect 787 5530 791 5534
rect 827 5530 831 5534
rect 1087 5642 1091 5646
rect 1207 5642 1211 5646
rect 1327 5642 1331 5646
rect 1479 5642 1483 5646
rect 1583 5642 1587 5646
rect 1975 5718 1979 5722
rect 2511 5718 2515 5722
rect 2663 5718 2667 5722
rect 2815 5718 2819 5722
rect 2975 5718 2979 5722
rect 3143 5718 3147 5722
rect 3319 5718 3323 5722
rect 3495 5718 3499 5722
rect 3799 5718 3803 5722
rect 1751 5642 1755 5646
rect 1815 5642 1819 5646
rect 1179 5560 1183 5564
rect 923 5530 927 5534
rect 1059 5530 1063 5534
rect 1195 5530 1199 5534
rect 1299 5530 1303 5534
rect 1935 5642 1939 5646
rect 1975 5598 1979 5602
rect 1995 5598 1999 5602
rect 2203 5598 2207 5602
rect 2435 5598 2439 5602
rect 2483 5598 2487 5602
rect 2635 5598 2639 5602
rect 2659 5598 2663 5602
rect 1331 5530 1335 5534
rect 1555 5530 1559 5534
rect 1787 5530 1791 5534
rect 1935 5530 1939 5534
rect 111 5398 115 5402
rect 815 5398 819 5402
rect 903 5398 907 5402
rect 951 5398 955 5402
rect 1039 5398 1043 5402
rect 1087 5398 1091 5402
rect 1183 5398 1187 5402
rect 1223 5398 1227 5402
rect 111 5282 115 5286
rect 587 5282 591 5286
rect 739 5282 743 5286
rect 875 5282 879 5286
rect 899 5282 903 5286
rect 1011 5282 1015 5286
rect 1067 5282 1071 5286
rect 1335 5398 1339 5402
rect 1359 5398 1363 5402
rect 2787 5598 2791 5602
rect 2867 5598 2871 5602
rect 2947 5598 2951 5602
rect 3075 5598 3079 5602
rect 3115 5598 3119 5602
rect 3275 5598 3279 5602
rect 3291 5598 3295 5602
rect 3467 5598 3471 5602
rect 3475 5598 3479 5602
rect 3651 5598 3655 5602
rect 3839 5670 3843 5674
rect 4107 5670 4111 5674
rect 4243 5670 4247 5674
rect 4379 5670 4383 5674
rect 4515 5670 4519 5674
rect 4651 5670 4655 5674
rect 4787 5670 4791 5674
rect 4923 5670 4927 5674
rect 5059 5670 5063 5674
rect 5195 5670 5199 5674
rect 5663 5670 5667 5674
rect 3799 5598 3803 5602
rect 3839 5526 3843 5530
rect 4135 5526 4139 5530
rect 4271 5526 4275 5530
rect 4303 5526 4307 5530
rect 1975 5486 1979 5490
rect 2023 5486 2027 5490
rect 1495 5398 1499 5402
rect 1663 5398 1667 5402
rect 1815 5398 1819 5402
rect 1935 5398 1939 5402
rect 1155 5282 1159 5286
rect 1243 5282 1247 5286
rect 1307 5282 1311 5286
rect 1427 5282 1431 5286
rect 1467 5282 1471 5286
rect 111 5158 115 5162
rect 367 5158 371 5162
rect 535 5158 539 5162
rect 615 5158 619 5162
rect 111 5042 115 5046
rect 131 5042 135 5046
rect 323 5042 327 5046
rect 339 5042 343 5046
rect 507 5042 511 5046
rect 555 5042 559 5046
rect 711 5158 715 5162
rect 767 5158 771 5162
rect 895 5158 899 5162
rect 927 5158 931 5162
rect 1079 5158 1083 5162
rect 1095 5158 1099 5162
rect 1263 5158 1267 5162
rect 1271 5158 1275 5162
rect 1447 5158 1451 5162
rect 1455 5158 1459 5162
rect 1619 5282 1623 5286
rect 1635 5282 1639 5286
rect 1787 5282 1791 5286
rect 1975 5350 1979 5354
rect 1995 5350 1999 5354
rect 2051 5350 2055 5354
rect 2167 5486 2171 5490
rect 2231 5486 2235 5490
rect 2343 5486 2347 5490
rect 2463 5486 2467 5490
rect 2527 5486 2531 5490
rect 2139 5350 2143 5354
rect 2315 5350 2319 5354
rect 4407 5526 4411 5530
rect 4511 5526 4515 5530
rect 4543 5526 4547 5530
rect 4679 5526 4683 5530
rect 4719 5526 4723 5530
rect 4815 5526 4819 5530
rect 4927 5526 4931 5530
rect 4951 5526 4955 5530
rect 5087 5526 5091 5530
rect 5135 5526 5139 5530
rect 5223 5526 5227 5530
rect 2687 5486 2691 5490
rect 2719 5486 2723 5490
rect 2895 5486 2899 5490
rect 2911 5486 2915 5490
rect 3103 5486 3107 5490
rect 3111 5486 3115 5490
rect 3303 5486 3307 5490
rect 3311 5486 3315 5490
rect 3503 5486 3507 5490
rect 3679 5486 3683 5490
rect 3799 5486 3803 5490
rect 2459 5350 2463 5354
rect 2499 5350 2503 5354
rect 2691 5350 2695 5354
rect 2859 5350 2863 5354
rect 2883 5350 2887 5354
rect 1935 5282 1939 5286
rect 1975 5238 1979 5242
rect 2079 5238 2083 5242
rect 1631 5158 1635 5162
rect 1647 5158 1651 5162
rect 683 5042 687 5046
rect 811 5042 815 5046
rect 867 5042 871 5046
rect 1051 5042 1055 5046
rect 1083 5042 1087 5046
rect 1235 5042 1239 5046
rect 1371 5042 1375 5046
rect 1419 5042 1423 5046
rect 1603 5042 1607 5046
rect 1659 5042 1663 5046
rect 1815 5158 1819 5162
rect 1935 5158 1939 5162
rect 2239 5238 2243 5242
rect 2487 5238 2491 5242
rect 2591 5238 2595 5242
rect 3083 5350 3087 5354
rect 3267 5350 3271 5354
rect 3283 5350 3287 5354
rect 3651 5350 3655 5354
rect 2887 5238 2891 5242
rect 2943 5238 2947 5242
rect 3295 5238 3299 5242
rect 3303 5238 3307 5242
rect 3663 5238 3667 5242
rect 3679 5238 3683 5242
rect 3839 5390 3843 5394
rect 3859 5390 3863 5394
rect 3995 5390 3999 5394
rect 4131 5390 4135 5394
rect 4275 5390 4279 5394
rect 4435 5390 4439 5394
rect 4483 5390 4487 5394
rect 3799 5350 3803 5354
rect 4603 5390 4607 5394
rect 4691 5390 4695 5394
rect 4779 5390 4783 5394
rect 4899 5390 4903 5394
rect 4963 5390 4967 5394
rect 3839 5274 3843 5278
rect 3887 5274 3891 5278
rect 3999 5274 4003 5278
rect 4023 5274 4027 5278
rect 4159 5274 4163 5278
rect 3799 5238 3803 5242
rect 1975 5126 1979 5130
rect 2211 5126 2215 5130
rect 2267 5126 2271 5130
rect 2515 5126 2519 5130
rect 2563 5126 2567 5130
rect 2755 5126 2759 5130
rect 2915 5126 2919 5130
rect 2995 5126 2999 5130
rect 1787 5042 1791 5046
rect 1935 5042 1939 5046
rect 1975 4982 1979 4986
rect 2183 4982 2187 4986
rect 2295 4982 2299 4986
rect 2319 4982 2323 4986
rect 111 4906 115 4910
rect 159 4906 163 4910
rect 295 4906 299 4910
rect 351 4906 355 4910
rect 431 4906 435 4910
rect 111 4782 115 4786
rect 131 4782 135 4786
rect 567 4906 571 4910
rect 583 4906 587 4910
rect 703 4906 707 4910
rect 839 4906 843 4910
rect 1111 4906 1115 4910
rect 1399 4906 1403 4910
rect 1687 4906 1691 4910
rect 1935 4906 1939 4910
rect 2455 4982 2459 4986
rect 2543 4982 2547 4986
rect 2599 4982 2603 4986
rect 2743 4982 2747 4986
rect 2783 4982 2787 4986
rect 4199 5274 4203 5278
rect 4303 5274 4307 5278
rect 4399 5274 4403 5278
rect 4463 5274 4467 5278
rect 4607 5274 4611 5278
rect 4631 5274 4635 5278
rect 5663 5526 5667 5530
rect 5107 5390 5111 5394
rect 5663 5390 5667 5394
rect 4807 5274 4811 5278
rect 4823 5274 4827 5278
rect 3839 5142 3843 5146
rect 3971 5142 3975 5146
rect 4099 5142 4103 5146
rect 4171 5142 4175 5146
rect 4347 5142 4351 5146
rect 4371 5142 4375 5146
rect 3235 5126 3239 5130
rect 3275 5126 3279 5130
rect 3475 5126 3479 5130
rect 3635 5126 3639 5130
rect 3799 5126 3803 5130
rect 2895 4982 2899 4986
rect 3023 4982 3027 4986
rect 3047 4982 3051 4986
rect 3199 4982 3203 4986
rect 3263 4982 3267 4986
rect 3351 4982 3355 4986
rect 4579 5142 4583 5146
rect 4595 5142 4599 5146
rect 3839 5014 3843 5018
rect 3983 5014 3987 5018
rect 4127 5014 4131 5018
rect 3503 4982 3507 4986
rect 3799 4982 3803 4986
rect 1975 4862 1979 4866
rect 2155 4862 2159 4866
rect 2291 4862 2295 4866
rect 2427 4862 2431 4866
rect 2571 4862 2575 4866
rect 2715 4862 2719 4866
rect 2723 4862 2727 4866
rect 267 4782 271 4786
rect 403 4782 407 4786
rect 539 4782 543 4786
rect 675 4782 679 4786
rect 1935 4782 1939 4786
rect 2867 4862 2871 4866
rect 2875 4862 2879 4866
rect 3839 4878 3843 4882
rect 3859 4878 3863 4882
rect 3955 4878 3959 4882
rect 4075 4878 4079 4882
rect 3019 4862 3023 4866
rect 3027 4862 3031 4866
rect 3171 4862 3175 4866
rect 3179 4862 3183 4866
rect 3323 4862 3327 4866
rect 3799 4862 3803 4866
rect 1975 4746 1979 4750
rect 2023 4746 2027 4750
rect 2159 4746 2163 4750
rect 2295 4746 2299 4750
rect 2431 4746 2435 4750
rect 2455 4746 2459 4750
rect 2567 4746 2571 4750
rect 2599 4746 2603 4750
rect 2703 4746 2707 4750
rect 2751 4746 2755 4750
rect 2839 4746 2843 4750
rect 2903 4746 2907 4750
rect 2975 4746 2979 4750
rect 3055 4746 3059 4750
rect 3111 4746 3115 4750
rect 3207 4746 3211 4750
rect 3247 4746 3251 4750
rect 4223 5014 4227 5018
rect 4375 5014 4379 5018
rect 4447 5014 4451 5018
rect 4991 5274 4995 5278
rect 5039 5274 5043 5278
rect 5663 5274 5667 5278
rect 4795 5142 4799 5146
rect 4843 5142 4847 5146
rect 5011 5142 5015 5146
rect 5099 5142 5103 5146
rect 5663 5142 5667 5146
rect 4623 5014 4627 5018
rect 4655 5014 4659 5018
rect 4855 5014 4859 5018
rect 4871 5014 4875 5018
rect 4195 4878 4199 4882
rect 4299 4878 4303 4882
rect 4419 4878 4423 4882
rect 4507 4878 4511 4882
rect 4627 4878 4631 4882
rect 4699 4878 4703 4882
rect 3839 4766 3843 4770
rect 3887 4766 3891 4770
rect 3399 4746 3403 4750
rect 3543 4746 3547 4750
rect 3679 4746 3683 4750
rect 3799 4746 3803 4750
rect 111 4662 115 4666
rect 159 4662 163 4666
rect 295 4662 299 4666
rect 431 4662 435 4666
rect 567 4662 571 4666
rect 703 4662 707 4666
rect 111 4542 115 4546
rect 131 4542 135 4546
rect 267 4542 271 4546
rect 339 4542 343 4546
rect 403 4542 407 4546
rect 515 4542 519 4546
rect 539 4542 543 4546
rect 675 4542 679 4546
rect 691 4542 695 4546
rect 1935 4662 1939 4666
rect 1975 4602 1979 4606
rect 1995 4602 1999 4606
rect 2131 4602 2135 4606
rect 2267 4602 2271 4606
rect 2323 4602 2327 4606
rect 2403 4602 2407 4606
rect 875 4542 879 4546
rect 1059 4542 1063 4546
rect 1243 4542 1247 4546
rect 1427 4542 1431 4546
rect 1619 4542 1623 4546
rect 1787 4542 1791 4546
rect 1935 4542 1939 4546
rect 111 4430 115 4434
rect 367 4430 371 4434
rect 543 4430 547 4434
rect 567 4430 571 4434
rect 711 4430 715 4434
rect 719 4430 723 4434
rect 863 4430 867 4434
rect 903 4430 907 4434
rect 1023 4430 1027 4434
rect 1087 4430 1091 4434
rect 1183 4430 1187 4434
rect 1271 4430 1275 4434
rect 1343 4430 1347 4434
rect 2539 4602 2543 4606
rect 2579 4602 2583 4606
rect 2675 4602 2679 4606
rect 2811 4602 2815 4606
rect 2827 4602 2831 4606
rect 2947 4602 2951 4606
rect 3075 4602 3079 4606
rect 3083 4602 3087 4606
rect 3219 4602 3223 4606
rect 3315 4602 3319 4606
rect 3371 4602 3375 4606
rect 3515 4602 3519 4606
rect 3563 4602 3567 4606
rect 1975 4482 1979 4486
rect 2351 4482 2355 4486
rect 2543 4482 2547 4486
rect 2607 4482 2611 4486
rect 1455 4430 1459 4434
rect 1503 4430 1507 4434
rect 1647 4430 1651 4434
rect 1671 4430 1675 4434
rect 1815 4430 1819 4434
rect 111 4298 115 4302
rect 539 4298 543 4302
rect 627 4298 631 4302
rect 683 4298 687 4302
rect 771 4298 775 4302
rect 835 4298 839 4302
rect 923 4298 927 4302
rect 995 4298 999 4302
rect 1083 4298 1087 4302
rect 1155 4298 1159 4302
rect 1251 4298 1255 4302
rect 1315 4298 1319 4302
rect 1419 4298 1423 4302
rect 1475 4298 1479 4302
rect 4103 4766 4107 4770
rect 4327 4766 4331 4770
rect 4535 4766 4539 4770
rect 5039 5014 5043 5018
rect 5127 5014 5131 5018
rect 5215 5014 5219 5018
rect 5391 5014 5395 5018
rect 5543 5014 5547 5018
rect 5663 5014 5667 5018
rect 4827 4878 4831 4882
rect 4875 4878 4879 4882
rect 5011 4878 5015 4882
rect 5043 4878 5047 4882
rect 5187 4878 5191 4882
rect 5211 4878 5215 4882
rect 5363 4878 5367 4882
rect 5371 4878 5375 4882
rect 4727 4766 4731 4770
rect 4903 4766 4907 4770
rect 4943 4766 4947 4770
rect 5071 4766 5075 4770
rect 5087 4766 5091 4770
rect 5239 4766 5243 4770
rect 5515 4878 5519 4882
rect 5663 4878 5667 4882
rect 5399 4766 5403 4770
rect 5543 4766 5547 4770
rect 3839 4630 3843 4634
rect 4771 4630 4775 4634
rect 4915 4630 4919 4634
rect 4955 4630 4959 4634
rect 5059 4630 5063 4634
rect 5147 4630 5151 4634
rect 5211 4630 5215 4634
rect 5339 4630 5343 4634
rect 5371 4630 5375 4634
rect 3651 4602 3655 4606
rect 3799 4602 3803 4606
rect 4867 4568 4871 4572
rect 5423 4568 5427 4572
rect 2783 4482 2787 4486
rect 2855 4482 2859 4486
rect 1935 4430 1939 4434
rect 3839 4506 3843 4510
rect 4487 4506 4491 4510
rect 4671 4506 4675 4510
rect 4799 4506 4803 4510
rect 4879 4506 4883 4510
rect 4983 4506 4987 4510
rect 5095 4506 5099 4510
rect 5175 4506 5179 4510
rect 5327 4506 5331 4510
rect 5367 4506 5371 4510
rect 3015 4482 3019 4486
rect 3103 4482 3107 4486
rect 3247 4482 3251 4486
rect 3343 4482 3347 4486
rect 3471 4482 3475 4486
rect 3591 4482 3595 4486
rect 3679 4482 3683 4486
rect 3799 4482 3803 4486
rect 5663 4766 5667 4770
rect 5515 4630 5519 4634
rect 5663 4630 5667 4634
rect 5543 4506 5547 4510
rect 1975 4358 1979 4362
rect 1995 4358 1999 4362
rect 2379 4358 2383 4362
rect 2515 4358 2519 4362
rect 2755 4358 2759 4362
rect 2803 4358 2807 4362
rect 1595 4298 1599 4302
rect 1643 4298 1647 4302
rect 1787 4298 1791 4302
rect 1935 4298 1939 4302
rect 111 4182 115 4186
rect 519 4182 523 4186
rect 655 4182 659 4186
rect 703 4182 707 4186
rect 799 4182 803 4186
rect 111 4070 115 4074
rect 131 4070 135 4074
rect 339 4070 343 4074
rect 491 4070 495 4074
rect 595 4070 599 4074
rect 675 4070 679 4074
rect 895 4182 899 4186
rect 951 4182 955 4186
rect 1103 4182 1107 4186
rect 1111 4182 1115 4186
rect 1279 4182 1283 4186
rect 1327 4182 1331 4186
rect 1447 4182 1451 4186
rect 1551 4182 1555 4186
rect 1623 4182 1627 4186
rect 1783 4182 1787 4186
rect 2987 4358 2991 4362
rect 3219 4358 3223 4362
rect 3235 4358 3239 4362
rect 3443 4358 3447 4362
rect 3651 4358 3655 4362
rect 1975 4218 1979 4222
rect 2023 4218 2027 4222
rect 2191 4218 2195 4222
rect 2383 4218 2387 4222
rect 2407 4218 2411 4222
rect 1935 4182 1939 4186
rect 867 4070 871 4074
rect 875 4070 879 4074
rect 1075 4070 1079 4074
rect 1179 4070 1183 4074
rect 1299 4070 1303 4074
rect 1491 4070 1495 4074
rect 1523 4070 1527 4074
rect 1975 4106 1979 4110
rect 1995 4106 1999 4110
rect 2075 4106 2079 4110
rect 2163 4106 2167 4110
rect 2259 4106 2263 4110
rect 1755 4070 1759 4074
rect 1787 4070 1791 4074
rect 1935 4070 1939 4074
rect 111 3954 115 3958
rect 159 3954 163 3958
rect 343 3954 347 3958
rect 367 3954 371 3958
rect 567 3954 571 3958
rect 623 3954 627 3958
rect 807 3954 811 3958
rect 903 3954 907 3958
rect 1055 3954 1059 3958
rect 1207 3954 1211 3958
rect 1311 3954 1315 3958
rect 1519 3954 1523 3958
rect 1575 3954 1579 3958
rect 1815 3954 1819 3958
rect 111 3834 115 3838
rect 131 3834 135 3838
rect 267 3834 271 3838
rect 315 3834 319 3838
rect 2583 4218 2587 4222
rect 2783 4218 2787 4222
rect 2831 4218 2835 4222
rect 2983 4218 2987 4222
rect 3839 4370 3843 4374
rect 3859 4370 3863 4374
rect 3995 4370 3999 4374
rect 4131 4370 4135 4374
rect 4283 4370 4287 4374
rect 4459 4370 4463 4374
rect 4483 4370 4487 4374
rect 3799 4358 3803 4362
rect 3839 4258 3843 4262
rect 3887 4258 3891 4262
rect 4023 4258 4027 4262
rect 4159 4258 4163 4262
rect 3263 4218 3267 4222
rect 3679 4218 3683 4222
rect 3799 4218 3803 4222
rect 2355 4106 2359 4110
rect 2443 4106 2447 4110
rect 2555 4106 2559 4110
rect 4379 4272 4383 4276
rect 4643 4370 4647 4374
rect 4715 4370 4719 4374
rect 4851 4370 4855 4374
rect 4979 4370 4983 4374
rect 5067 4370 5071 4374
rect 5251 4370 5255 4374
rect 5299 4370 5303 4374
rect 5515 4370 5519 4374
rect 5663 4506 5667 4510
rect 5663 4370 5667 4374
rect 5367 4272 5371 4276
rect 4303 4258 4307 4262
rect 4311 4258 4315 4262
rect 4503 4258 4507 4262
rect 4511 4258 4515 4262
rect 4735 4258 4739 4262
rect 4743 4258 4747 4262
rect 4999 4258 5003 4262
rect 5007 4258 5011 4262
rect 5271 4258 5275 4262
rect 5279 4258 5283 4262
rect 5543 4258 5547 4262
rect 5663 4258 5667 4262
rect 2619 4106 2623 4110
rect 2755 4106 2759 4110
rect 2787 4106 2791 4110
rect 2955 4106 2959 4110
rect 3131 4106 3135 4110
rect 3799 4106 3803 4110
rect 3839 4106 3843 4110
rect 3859 4106 3863 4110
rect 3995 4106 3999 4110
rect 4131 4106 4135 4110
rect 4275 4106 4279 4110
rect 4475 4106 4479 4110
rect 4563 4106 4567 4110
rect 4699 4106 4703 4110
rect 4707 4106 4711 4110
rect 4835 4106 4839 4110
rect 4971 4106 4975 4110
rect 5107 4106 5111 4110
rect 5243 4106 5247 4110
rect 5379 4106 5383 4110
rect 5515 4106 5519 4110
rect 5663 4106 5667 4110
rect 1975 3986 1979 3990
rect 2103 3986 2107 3990
rect 2127 3986 2131 3990
rect 1935 3954 1939 3958
rect 475 3834 479 3838
rect 539 3834 543 3838
rect 707 3834 711 3838
rect 779 3834 783 3838
rect 963 3834 967 3838
rect 1027 3834 1031 3838
rect 1235 3834 1239 3838
rect 1283 3834 1287 3838
rect 2287 3986 2291 3990
rect 2311 3986 2315 3990
rect 2471 3986 2475 3990
rect 2487 3986 2491 3990
rect 2647 3986 2651 3990
rect 2663 3986 2667 3990
rect 2815 3986 2819 3990
rect 2831 3986 2835 3990
rect 2983 3986 2987 3990
rect 2999 3986 3003 3990
rect 3159 3986 3163 3990
rect 3175 3986 3179 3990
rect 3351 3986 3355 3990
rect 3799 3986 3803 3990
rect 3839 3974 3843 3978
rect 4359 3974 4363 3978
rect 4543 3974 4547 3978
rect 4591 3974 4595 3978
rect 4727 3974 4731 3978
rect 4735 3974 4739 3978
rect 4863 3974 4867 3978
rect 4927 3974 4931 3978
rect 1975 3866 1979 3870
rect 2099 3866 2103 3870
rect 2283 3866 2287 3870
rect 2291 3866 2295 3870
rect 2459 3866 2463 3870
rect 2523 3866 2527 3870
rect 1515 3834 1519 3838
rect 1547 3834 1551 3838
rect 1787 3834 1791 3838
rect 1935 3834 1939 3838
rect 111 3718 115 3722
rect 295 3718 299 3722
rect 503 3718 507 3722
rect 631 3718 635 3722
rect 735 3718 739 3722
rect 775 3718 779 3722
rect 927 3718 931 3722
rect 991 3718 995 3722
rect 1087 3718 1091 3722
rect 1255 3718 1259 3722
rect 1263 3718 1267 3722
rect 1423 3718 1427 3722
rect 1543 3718 1547 3722
rect 1591 3718 1595 3722
rect 1759 3718 1763 3722
rect 1815 3718 1819 3722
rect 2635 3866 2639 3870
rect 2739 3866 2743 3870
rect 2803 3866 2807 3870
rect 2947 3866 2951 3870
rect 2971 3866 2975 3870
rect 3147 3866 3151 3870
rect 3155 3866 3159 3870
rect 3323 3866 3327 3870
rect 3355 3866 3359 3870
rect 3563 3866 3567 3870
rect 3799 3866 3803 3870
rect 1975 3750 1979 3754
rect 2319 3750 2323 3754
rect 2407 3750 2411 3754
rect 2551 3750 2555 3754
rect 1935 3718 1939 3722
rect 111 3594 115 3598
rect 603 3594 607 3598
rect 747 3594 751 3598
rect 779 3594 783 3598
rect 899 3594 903 3598
rect 915 3594 919 3598
rect 1051 3594 1055 3598
rect 1059 3594 1063 3598
rect 1187 3594 1191 3598
rect 1227 3594 1231 3598
rect 1323 3594 1327 3598
rect 1395 3594 1399 3598
rect 1459 3594 1463 3598
rect 1563 3594 1567 3598
rect 1595 3594 1599 3598
rect 1731 3594 1735 3598
rect 111 3458 115 3462
rect 727 3458 731 3462
rect 807 3458 811 3462
rect 863 3458 867 3462
rect 943 3458 947 3462
rect 999 3458 1003 3462
rect 1079 3458 1083 3462
rect 1135 3458 1139 3462
rect 1215 3458 1219 3462
rect 1271 3458 1275 3462
rect 1351 3458 1355 3462
rect 1975 3630 1979 3634
rect 2379 3630 2383 3634
rect 2411 3630 2415 3634
rect 1935 3594 1939 3598
rect 2647 3750 2651 3754
rect 2767 3750 2771 3754
rect 2871 3750 2875 3754
rect 2975 3750 2979 3754
rect 3087 3750 3091 3754
rect 3183 3750 3187 3754
rect 3295 3750 3299 3754
rect 3383 3750 3387 3754
rect 3839 3854 3843 3858
rect 4051 3854 4055 3858
rect 4267 3854 4271 3858
rect 4331 3854 4335 3858
rect 4483 3854 4487 3858
rect 4515 3854 4519 3858
rect 4999 3974 5003 3978
rect 5127 3974 5131 3978
rect 5135 3974 5139 3978
rect 5271 3974 5275 3978
rect 5327 3974 5331 3978
rect 5407 3974 5411 3978
rect 5527 3974 5531 3978
rect 5543 3974 5547 3978
rect 4699 3854 4703 3858
rect 4707 3854 4711 3858
rect 4899 3854 4903 3858
rect 4907 3854 4911 3858
rect 5099 3854 5103 3858
rect 5115 3854 5119 3858
rect 5299 3854 5303 3858
rect 5323 3854 5327 3858
rect 5499 3854 5503 3858
rect 5515 3854 5519 3858
rect 5663 3974 5667 3978
rect 5663 3854 5667 3858
rect 3495 3750 3499 3754
rect 3591 3750 3595 3754
rect 3679 3750 3683 3754
rect 3799 3750 3803 3754
rect 3839 3714 3843 3718
rect 3887 3714 3891 3718
rect 4055 3714 4059 3718
rect 4079 3714 4083 3718
rect 2547 3630 2551 3634
rect 2619 3630 2623 3634
rect 2683 3630 2687 3634
rect 2843 3630 2847 3634
rect 3059 3630 3063 3634
rect 3267 3630 3271 3634
rect 3467 3630 3471 3634
rect 3651 3630 3655 3634
rect 3799 3630 3803 3634
rect 1407 3458 1411 3462
rect 111 3342 115 3346
rect 699 3342 703 3346
rect 755 3342 759 3346
rect 835 3342 839 3346
rect 1975 3478 1979 3482
rect 2439 3478 2443 3482
rect 2575 3478 2579 3482
rect 2599 3478 2603 3482
rect 2711 3478 2715 3482
rect 1487 3458 1491 3462
rect 1543 3458 1547 3462
rect 1623 3458 1627 3462
rect 1679 3458 1683 3462
rect 1759 3458 1763 3462
rect 1815 3458 1819 3462
rect 1935 3458 1939 3462
rect 891 3342 895 3346
rect 971 3342 975 3346
rect 1035 3342 1039 3346
rect 1107 3342 1111 3346
rect 1187 3342 1191 3346
rect 1243 3342 1247 3346
rect 1339 3342 1343 3346
rect 1379 3342 1383 3346
rect 1491 3342 1495 3346
rect 1515 3342 1519 3346
rect 1651 3342 1655 3346
rect 1787 3342 1791 3346
rect 111 3230 115 3234
rect 391 3230 395 3234
rect 647 3230 651 3234
rect 783 3230 787 3234
rect 919 3230 923 3234
rect 927 3230 931 3234
rect 111 3106 115 3110
rect 131 3106 135 3110
rect 307 3106 311 3110
rect 363 3106 367 3110
rect 1063 3230 1067 3234
rect 1215 3230 1219 3234
rect 1223 3230 1227 3234
rect 1367 3230 1371 3234
rect 1975 3358 1979 3362
rect 2531 3358 2535 3362
rect 2571 3358 2575 3362
rect 1935 3342 1939 3346
rect 2823 3478 2827 3482
rect 3047 3478 3051 3482
rect 3263 3478 3267 3482
rect 3479 3478 3483 3482
rect 3679 3478 3683 3482
rect 3839 3602 3843 3606
rect 3859 3602 3863 3606
rect 4247 3714 4251 3718
rect 4295 3714 4299 3718
rect 4439 3714 4443 3718
rect 4511 3714 4515 3718
rect 4631 3714 4635 3718
rect 4727 3714 4731 3718
rect 4935 3714 4939 3718
rect 5143 3714 5147 3718
rect 5351 3714 5355 3718
rect 5543 3714 5547 3718
rect 5663 3714 5667 3718
rect 3995 3602 3999 3606
rect 4027 3602 4031 3606
rect 4131 3602 4135 3606
rect 4219 3602 4223 3606
rect 4267 3602 4271 3606
rect 4403 3602 4407 3606
rect 4411 3602 4415 3606
rect 4539 3602 4543 3606
rect 4603 3602 4607 3606
rect 4675 3602 4679 3606
rect 3955 3592 3959 3596
rect 4527 3592 4531 3596
rect 4811 3602 4815 3606
rect 4947 3602 4951 3606
rect 5083 3602 5087 3606
rect 5663 3602 5667 3606
rect 3799 3478 3803 3482
rect 3839 3482 3843 3486
rect 3887 3482 3891 3486
rect 4023 3482 4027 3486
rect 4159 3482 4163 3486
rect 4295 3482 4299 3486
rect 4431 3482 4435 3486
rect 4567 3482 4571 3486
rect 4703 3482 4707 3486
rect 4831 3482 4835 3486
rect 4839 3482 4843 3486
rect 4967 3482 4971 3486
rect 2715 3358 2719 3362
rect 2795 3358 2799 3362
rect 2899 3358 2903 3362
rect 3019 3358 3023 3362
rect 3083 3358 3087 3362
rect 1519 3230 1523 3234
rect 1527 3230 1531 3234
rect 1679 3230 1683 3234
rect 1815 3230 1819 3234
rect 507 3106 511 3110
rect 619 3106 623 3110
rect 707 3106 711 3110
rect 899 3106 903 3110
rect 111 2990 115 2994
rect 159 2990 163 2994
rect 295 2990 299 2994
rect 335 2990 339 2994
rect 431 2990 435 2994
rect 535 2990 539 2994
rect 567 2990 571 2994
rect 703 2990 707 2994
rect 735 2990 739 2994
rect 1091 3106 1095 3110
rect 1195 3106 1199 3110
rect 1275 3106 1279 3110
rect 1451 3106 1455 3110
rect 1499 3106 1503 3110
rect 1975 3246 1979 3250
rect 2023 3246 2027 3250
rect 2255 3246 2259 3250
rect 2503 3246 2507 3250
rect 2559 3246 2563 3250
rect 1935 3230 1939 3234
rect 1975 3134 1979 3138
rect 1995 3134 1999 3138
rect 2227 3134 2231 3138
rect 1627 3106 1631 3110
rect 1787 3106 1791 3110
rect 1935 3106 1939 3110
rect 2475 3134 2479 3138
rect 2483 3134 2487 3138
rect 2743 3246 2747 3250
rect 2927 3246 2931 3250
rect 2975 3246 2979 3250
rect 4975 3482 4979 3486
rect 5103 3482 5107 3486
rect 5111 3482 5115 3486
rect 5239 3482 5243 3486
rect 5375 3482 5379 3486
rect 5663 3482 5667 3486
rect 3839 3370 3843 3374
rect 3859 3370 3863 3374
rect 4139 3370 4143 3374
rect 4427 3370 4431 3374
rect 4691 3370 4695 3374
rect 4803 3370 4807 3374
rect 4939 3370 4943 3374
rect 5075 3370 5079 3374
rect 5179 3370 5183 3374
rect 5211 3370 5215 3374
rect 5347 3370 5351 3374
rect 5427 3370 5431 3374
rect 3235 3358 3239 3362
rect 3267 3358 3271 3362
rect 3451 3358 3455 3362
rect 3651 3358 3655 3362
rect 3799 3358 3803 3362
rect 3111 3246 3115 3250
rect 3207 3246 3211 3250
rect 3295 3246 3299 3250
rect 2715 3134 2719 3138
rect 2779 3134 2783 3138
rect 2947 3134 2951 3138
rect 3075 3134 3079 3138
rect 3179 3134 3183 3138
rect 3447 3246 3451 3250
rect 3799 3246 3803 3250
rect 3839 3234 3843 3238
rect 3887 3234 3891 3238
rect 3911 3234 3915 3238
rect 4523 3320 4527 3324
rect 5059 3320 5063 3324
rect 5663 3370 5667 3374
rect 4167 3234 4171 3238
rect 4183 3234 4187 3238
rect 4439 3234 4443 3238
rect 4455 3234 4459 3238
rect 4687 3234 4691 3238
rect 4719 3234 4723 3238
rect 3371 3134 3375 3138
rect 3419 3134 3423 3138
rect 3651 3134 3655 3138
rect 3799 3134 3803 3138
rect 1975 3014 1979 3018
rect 2191 3014 2195 3018
rect 2351 3014 2355 3018
rect 2511 3014 2515 3018
rect 2519 3014 2523 3018
rect 927 2990 931 2994
rect 1119 2990 1123 2994
rect 1303 2990 1307 2994
rect 1479 2990 1483 2994
rect 1655 2990 1659 2994
rect 1815 2990 1819 2994
rect 1935 2990 1939 2994
rect 111 2874 115 2878
rect 131 2874 135 2878
rect 227 2874 231 2878
rect 267 2874 271 2878
rect 363 2874 367 2878
rect 403 2874 407 2878
rect 499 2874 503 2878
rect 539 2874 543 2878
rect 635 2874 639 2878
rect 675 2874 679 2878
rect 1975 2898 1979 2902
rect 1995 2898 1999 2902
rect 2131 2898 2135 2902
rect 2163 2898 2167 2902
rect 2267 2898 2271 2902
rect 771 2874 775 2878
rect 1935 2874 1939 2878
rect 111 2758 115 2762
rect 255 2758 259 2762
rect 375 2758 379 2762
rect 391 2758 395 2762
rect 527 2758 531 2762
rect 575 2758 579 2762
rect 663 2758 667 2762
rect 799 2758 803 2762
rect 2703 3014 2707 3018
rect 2807 3014 2811 3018
rect 2903 3014 2907 3018
rect 3103 3014 3107 3018
rect 3119 3014 3123 3018
rect 3839 3118 3843 3122
rect 3883 3118 3887 3122
rect 3931 3118 3935 3122
rect 3335 3014 3339 3018
rect 3399 3014 3403 3018
rect 3559 3014 3563 3018
rect 3679 3014 3683 3018
rect 2323 2898 2327 2902
rect 2403 2898 2407 2902
rect 2491 2898 2495 2902
rect 2539 2898 2543 2902
rect 2675 2898 2679 2902
rect 2683 2898 2687 2902
rect 2835 2898 2839 2902
rect 2875 2898 2879 2902
rect 111 2646 115 2650
rect 347 2646 351 2650
rect 387 2646 391 2650
rect 1975 2782 1979 2786
rect 2023 2782 2027 2786
rect 2159 2782 2163 2786
rect 1039 2758 1043 2762
rect 1295 2758 1299 2762
rect 1567 2758 1571 2762
rect 1815 2758 1819 2762
rect 1935 2758 1939 2762
rect 539 2646 543 2650
rect 547 2646 551 2650
rect 699 2646 703 2650
rect 771 2646 775 2650
rect 867 2646 871 2650
rect 1011 2646 1015 2650
rect 1035 2646 1039 2650
rect 1203 2646 1207 2650
rect 1267 2646 1271 2650
rect 1371 2646 1375 2650
rect 111 2534 115 2538
rect 327 2534 331 2538
rect 415 2534 419 2538
rect 535 2534 539 2538
rect 567 2534 571 2538
rect 1539 2646 1543 2650
rect 2295 2782 2299 2786
rect 2303 2782 2307 2786
rect 2431 2782 2435 2786
rect 2463 2782 2467 2786
rect 2567 2782 2571 2786
rect 2623 2782 2627 2786
rect 2711 2782 2715 2786
rect 2995 2898 2999 2902
rect 3091 2898 3095 2902
rect 3155 2898 3159 2902
rect 3307 2898 3311 2902
rect 3315 2898 3319 2902
rect 4131 3118 4135 3122
rect 4155 3118 4159 3122
rect 4331 3118 4335 3122
rect 4411 3118 4415 3122
rect 4523 3118 4527 3122
rect 3799 3014 3803 3018
rect 3839 2982 3843 2986
rect 3959 2982 3963 2986
rect 3999 2982 4003 2986
rect 4227 3099 4231 3100
rect 4227 3096 4231 3099
rect 4935 3234 4939 3238
rect 4967 3234 4971 3238
rect 5191 3234 5195 3238
rect 5207 3234 5211 3238
rect 5455 3234 5459 3238
rect 5663 3234 5667 3238
rect 4659 3118 4663 3122
rect 4715 3118 4719 3122
rect 4907 3118 4911 3122
rect 4915 3118 4919 3122
rect 5163 3118 5167 3122
rect 5663 3118 5667 3122
rect 5039 3096 5043 3100
rect 4159 2982 4163 2986
rect 4335 2982 4339 2986
rect 4359 2982 4363 2986
rect 3531 2898 3535 2902
rect 3799 2898 3803 2902
rect 3839 2854 3843 2858
rect 3859 2854 3863 2858
rect 3971 2854 3975 2858
rect 2783 2782 2787 2786
rect 2863 2782 2867 2786
rect 2943 2782 2947 2786
rect 3023 2782 3027 2786
rect 3103 2782 3107 2786
rect 1975 2662 1979 2666
rect 1995 2662 1999 2666
rect 2131 2662 2135 2666
rect 2275 2662 2279 2666
rect 2435 2662 2439 2666
rect 2595 2662 2599 2666
rect 2699 2662 2703 2666
rect 2755 2662 2759 2666
rect 1715 2646 1719 2650
rect 1787 2646 1791 2650
rect 1935 2646 1939 2650
rect 727 2534 731 2538
rect 735 2534 739 2538
rect 895 2534 899 2538
rect 919 2534 923 2538
rect 1063 2534 1067 2538
rect 1095 2534 1099 2538
rect 1231 2534 1235 2538
rect 1271 2534 1275 2538
rect 111 2418 115 2422
rect 131 2418 135 2422
rect 299 2418 303 2422
rect 403 2418 407 2422
rect 507 2418 511 2422
rect 691 2418 695 2422
rect 707 2418 711 2422
rect 891 2418 895 2422
rect 971 2418 975 2422
rect 1067 2418 1071 2422
rect 111 2290 115 2294
rect 159 2290 163 2294
rect 423 2290 427 2294
rect 431 2290 435 2294
rect 1975 2550 1979 2554
rect 2607 2550 2611 2554
rect 2727 2550 2731 2554
rect 2759 2550 2763 2554
rect 1399 2534 1403 2538
rect 1439 2534 1443 2538
rect 1567 2534 1571 2538
rect 1607 2534 1611 2538
rect 1743 2534 1747 2538
rect 1775 2534 1779 2538
rect 1935 2534 1939 2538
rect 2835 2662 2839 2666
rect 2915 2662 2919 2666
rect 2971 2662 2975 2666
rect 3183 2782 3187 2786
rect 3343 2782 3347 2786
rect 3799 2782 3803 2786
rect 4011 2854 4015 2858
rect 4131 2854 4135 2858
rect 4211 2854 4215 2858
rect 4307 2854 4311 2858
rect 4435 2854 4439 2858
rect 4519 2982 4523 2986
rect 4551 2982 4555 2986
rect 4719 2982 4723 2986
rect 4743 2982 4747 2986
rect 4927 2982 4931 2986
rect 4943 2982 4947 2986
rect 5135 2982 5139 2986
rect 5351 2982 5355 2986
rect 5543 2982 5547 2986
rect 5663 2982 5667 2986
rect 4491 2854 4495 2858
rect 4691 2854 4695 2858
rect 4899 2854 4903 2858
rect 4963 2854 4967 2858
rect 5107 2854 5111 2858
rect 5251 2854 5255 2858
rect 5323 2854 5327 2858
rect 5515 2854 5519 2858
rect 3839 2730 3843 2734
rect 3887 2730 3891 2734
rect 3967 2730 3971 2734
rect 4039 2730 4043 2734
rect 4223 2730 4227 2734
rect 4239 2730 4243 2734
rect 4463 2730 4467 2734
rect 4527 2730 4531 2734
rect 4719 2730 4723 2734
rect 4863 2730 4867 2734
rect 4991 2730 4995 2734
rect 5215 2730 5219 2734
rect 5279 2730 5283 2734
rect 3075 2662 3079 2666
rect 3799 2662 3803 2666
rect 3839 2618 3843 2622
rect 3891 2618 3895 2622
rect 3939 2618 3943 2622
rect 4067 2618 4071 2622
rect 2863 2550 2867 2554
rect 2911 2550 2915 2554
rect 2999 2550 3003 2554
rect 3063 2550 3067 2554
rect 1243 2418 1247 2422
rect 1251 2418 1255 2422
rect 1411 2418 1415 2422
rect 1531 2418 1535 2422
rect 1579 2418 1583 2422
rect 1747 2418 1751 2422
rect 1787 2418 1791 2422
rect 1935 2418 1939 2422
rect 1975 2422 1979 2426
rect 1995 2422 1999 2426
rect 2275 2422 2279 2426
rect 2571 2422 2575 2426
rect 2579 2422 2583 2426
rect 2731 2422 2735 2426
rect 2859 2422 2863 2426
rect 2883 2422 2887 2426
rect 711 2290 715 2294
rect 719 2290 723 2294
rect 999 2290 1003 2294
rect 1279 2290 1283 2294
rect 1295 2290 1299 2294
rect 111 2166 115 2170
rect 131 2166 135 2170
rect 395 2166 399 2170
rect 403 2166 407 2170
rect 683 2166 687 2170
rect 731 2166 735 2170
rect 971 2166 975 2170
rect 1083 2166 1087 2170
rect 111 2050 115 2054
rect 159 2050 163 2054
rect 223 2050 227 2054
rect 383 2050 387 2054
rect 431 2050 435 2054
rect 559 2050 563 2054
rect 1975 2298 1979 2302
rect 2023 2298 2027 2302
rect 1559 2290 1563 2294
rect 1815 2290 1819 2294
rect 1935 2290 1939 2294
rect 2159 2298 2163 2302
rect 2295 2298 2299 2302
rect 2303 2298 2307 2302
rect 2447 2298 2451 2302
rect 2599 2298 2603 2302
rect 2607 2298 2611 2302
rect 3223 2550 3227 2554
rect 3799 2550 3803 2554
rect 3839 2502 3843 2506
rect 3887 2502 3891 2506
rect 3919 2502 3923 2506
rect 4195 2618 4199 2622
rect 4267 2618 4271 2622
rect 4491 2618 4495 2622
rect 4499 2618 4503 2622
rect 4731 2618 4735 2622
rect 4835 2618 4839 2622
rect 4995 2618 4999 2622
rect 5187 2618 5191 2622
rect 5267 2618 5271 2622
rect 5663 2854 5667 2858
rect 5543 2730 5547 2734
rect 5515 2618 5519 2622
rect 4087 2502 4091 2506
rect 4095 2502 4099 2506
rect 4295 2502 4299 2506
rect 4319 2502 4323 2506
rect 4519 2502 4523 2506
rect 4567 2502 4571 2506
rect 4759 2502 4763 2506
rect 4823 2502 4827 2506
rect 5023 2502 5027 2506
rect 5087 2502 5091 2506
rect 3035 2422 3039 2426
rect 3147 2422 3151 2426
rect 3195 2422 3199 2426
rect 3435 2422 3439 2426
rect 3799 2422 3803 2426
rect 2767 2298 2771 2302
rect 2887 2298 2891 2302
rect 2927 2298 2931 2302
rect 3079 2298 3083 2302
rect 3175 2298 3179 2302
rect 3231 2298 3235 2302
rect 3383 2298 3387 2302
rect 3463 2298 3467 2302
rect 3543 2298 3547 2302
rect 1975 2178 1979 2182
rect 1995 2178 1999 2182
rect 2131 2178 2135 2182
rect 2267 2178 2271 2182
rect 2331 2178 2335 2182
rect 2419 2178 2423 2182
rect 2531 2178 2535 2182
rect 1267 2166 1271 2170
rect 1443 2166 1447 2170
rect 1787 2166 1791 2170
rect 1935 2166 1939 2170
rect 751 2050 755 2054
rect 759 2050 763 2054
rect 959 2050 963 2054
rect 1111 2050 1115 2054
rect 1167 2050 1171 2054
rect 1383 2050 1387 2054
rect 1471 2050 1475 2054
rect 111 1930 115 1934
rect 195 1930 199 1934
rect 355 1930 359 1934
rect 387 1930 391 1934
rect 531 1930 535 1934
rect 595 1930 599 1934
rect 723 1930 727 1934
rect 819 1930 823 1934
rect 111 1802 115 1806
rect 159 1802 163 1806
rect 223 1802 227 1806
rect 303 1802 307 1806
rect 415 1802 419 1806
rect 479 1802 483 1806
rect 931 1930 935 1934
rect 1051 1930 1055 1934
rect 1139 1930 1143 1934
rect 1283 1930 1287 1934
rect 1355 1930 1359 1934
rect 1607 2050 1611 2054
rect 1815 2050 1819 2054
rect 1975 2058 1979 2062
rect 2023 2058 2027 2062
rect 1935 2050 1939 2054
rect 2579 2178 2583 2182
rect 2731 2178 2735 2182
rect 2739 2178 2743 2182
rect 2899 2178 2903 2182
rect 2923 2178 2927 2182
rect 3051 2178 3055 2182
rect 3115 2178 3119 2182
rect 3203 2178 3207 2182
rect 3299 2178 3303 2182
rect 3355 2178 3359 2182
rect 3679 2298 3683 2302
rect 4387 2464 4391 2468
rect 3839 2390 3843 2394
rect 3859 2390 3863 2394
rect 4059 2390 4063 2394
rect 4091 2390 4095 2394
rect 5295 2502 5299 2506
rect 5351 2502 5355 2506
rect 5663 2730 5667 2734
rect 5663 2618 5667 2622
rect 5543 2502 5547 2506
rect 5115 2464 5119 2468
rect 4291 2390 4295 2394
rect 4339 2390 4343 2394
rect 4539 2390 4543 2394
rect 4579 2390 4583 2394
rect 4795 2390 4799 2394
rect 4811 2390 4815 2394
rect 5043 2390 5047 2394
rect 5059 2390 5063 2394
rect 5283 2390 5287 2394
rect 5323 2390 5327 2394
rect 5515 2390 5519 2394
rect 3799 2298 3803 2302
rect 3839 2254 3843 2258
rect 3887 2254 3891 2258
rect 4119 2254 4123 2258
rect 4367 2254 4371 2258
rect 4591 2254 4595 2258
rect 4607 2254 4611 2258
rect 4727 2254 4731 2258
rect 4839 2254 4843 2258
rect 4863 2254 4867 2258
rect 4999 2254 5003 2258
rect 5071 2254 5075 2258
rect 5135 2254 5139 2258
rect 3483 2178 3487 2182
rect 3515 2178 3519 2182
rect 3651 2178 3655 2182
rect 3799 2178 3803 2182
rect 2159 2058 2163 2062
rect 2279 2058 2283 2062
rect 2359 2058 2363 2062
rect 2551 2058 2555 2062
rect 2559 2058 2563 2062
rect 2759 2058 2763 2062
rect 2799 2058 2803 2062
rect 2951 2058 2955 2062
rect 3031 2058 3035 2062
rect 3143 2058 3147 2062
rect 1523 1930 1527 1934
rect 1579 1930 1583 1934
rect 1771 1930 1775 1934
rect 1787 1930 1791 1934
rect 1935 1930 1939 1934
rect 1975 1934 1979 1938
rect 1995 1934 1999 1938
rect 2251 1934 2255 1938
rect 2315 1934 2319 1938
rect 623 1802 627 1806
rect 655 1802 659 1806
rect 831 1802 835 1806
rect 847 1802 851 1806
rect 1007 1802 1011 1806
rect 1079 1802 1083 1806
rect 111 1686 115 1690
rect 131 1686 135 1690
rect 111 1554 115 1558
rect 159 1554 163 1558
rect 275 1686 279 1690
rect 451 1686 455 1690
rect 627 1686 631 1690
rect 803 1686 807 1690
rect 875 1686 879 1690
rect 1183 1802 1187 1806
rect 1311 1802 1315 1806
rect 1359 1802 1363 1806
rect 979 1686 983 1690
rect 1011 1686 1015 1690
rect 1147 1686 1151 1690
rect 1155 1686 1159 1690
rect 1283 1686 1287 1690
rect 1975 1818 1979 1822
rect 2023 1818 2027 1822
rect 2111 1818 2115 1822
rect 1535 1802 1539 1806
rect 1551 1802 1555 1806
rect 1711 1802 1715 1806
rect 1799 1802 1803 1806
rect 1935 1802 1939 1806
rect 2523 1934 2527 1938
rect 2619 1934 2623 1938
rect 2771 1934 2775 1938
rect 3255 2058 3259 2062
rect 3327 2058 3331 2062
rect 3479 2058 3483 2062
rect 3511 2058 3515 2062
rect 5271 2254 5275 2258
rect 5311 2254 5315 2258
rect 5407 2254 5411 2258
rect 5663 2502 5667 2506
rect 5663 2390 5667 2394
rect 5543 2254 5547 2258
rect 5663 2254 5667 2258
rect 3839 2126 3843 2130
rect 4563 2126 4567 2130
rect 4699 2126 4703 2130
rect 4835 2126 4839 2130
rect 4955 2126 4959 2130
rect 4971 2126 4975 2130
rect 5091 2126 5095 2130
rect 5107 2126 5111 2130
rect 5227 2126 5231 2130
rect 5243 2126 5247 2130
rect 5379 2126 5383 2130
rect 5515 2126 5519 2130
rect 3679 2058 3683 2062
rect 3799 2058 3803 2062
rect 3839 2014 3843 2018
rect 4727 2014 4731 2018
rect 4863 2014 4867 2018
rect 4983 2014 4987 2018
rect 5007 2014 5011 2018
rect 2899 1934 2903 1938
rect 3003 1934 3007 1938
rect 3163 1934 3167 1938
rect 3227 1934 3231 1938
rect 3419 1934 3423 1938
rect 3451 1934 3455 1938
rect 3651 1934 3655 1938
rect 2343 1818 2347 1822
rect 2391 1818 2395 1822
rect 2647 1818 2651 1822
rect 2663 1818 2667 1822
rect 2927 1818 2931 1822
rect 3183 1818 3187 1822
rect 3191 1818 3195 1822
rect 1331 1686 1335 1690
rect 1419 1686 1423 1690
rect 1507 1686 1511 1690
rect 1555 1686 1559 1690
rect 1683 1686 1687 1690
rect 1935 1686 1939 1690
rect 1975 1674 1979 1678
rect 2083 1674 2087 1678
rect 2219 1674 2223 1678
rect 2355 1674 2359 1678
rect 2363 1674 2367 1678
rect 2491 1674 2495 1678
rect 391 1554 395 1558
rect 631 1554 635 1558
rect 871 1554 875 1558
rect 903 1554 907 1558
rect 111 1430 115 1434
rect 131 1430 135 1434
rect 331 1430 335 1434
rect 363 1430 367 1434
rect 111 1318 115 1322
rect 159 1318 163 1322
rect 555 1430 559 1434
rect 603 1430 607 1434
rect 779 1430 783 1434
rect 843 1430 847 1434
rect 1039 1554 1043 1558
rect 1111 1554 1115 1558
rect 1175 1554 1179 1558
rect 1311 1554 1315 1558
rect 1351 1554 1355 1558
rect 1447 1554 1451 1558
rect 1583 1554 1587 1558
rect 1935 1554 1939 1558
rect 1975 1558 1979 1562
rect 2111 1558 2115 1562
rect 2143 1558 2147 1562
rect 2627 1674 2631 1678
rect 2635 1674 2639 1678
rect 3439 1818 3443 1822
rect 3447 1818 3451 1822
rect 3799 1934 3803 1938
rect 3839 1902 3843 1906
rect 4275 1902 4279 1906
rect 4499 1902 4503 1906
rect 4699 1902 4703 1906
rect 4731 1902 4735 1906
rect 4835 1902 4839 1906
rect 5119 2014 5123 2018
rect 5159 2014 5163 2018
rect 5255 2014 5259 2018
rect 5319 2014 5323 2018
rect 5487 2014 5491 2018
rect 4979 1902 4983 1906
rect 5131 1902 5135 1906
rect 5235 1902 5239 1906
rect 5291 1902 5295 1906
rect 3679 1818 3683 1822
rect 3799 1818 3803 1822
rect 3839 1782 3843 1786
rect 3887 1782 3891 1786
rect 4087 1782 4091 1786
rect 4303 1782 4307 1786
rect 4343 1782 4347 1786
rect 4527 1782 4531 1786
rect 4623 1782 4627 1786
rect 4759 1782 4763 1786
rect 2771 1674 2775 1678
rect 2899 1674 2903 1678
rect 2915 1674 2919 1678
rect 3155 1674 3159 1678
rect 3411 1674 3415 1678
rect 3651 1674 3655 1678
rect 3799 1674 3803 1678
rect 3839 1666 3843 1670
rect 3859 1666 3863 1670
rect 2247 1558 2251 1562
rect 2279 1558 2283 1562
rect 2383 1558 2387 1562
rect 2415 1558 2419 1562
rect 2519 1558 2523 1562
rect 2551 1558 2555 1562
rect 2655 1558 2659 1562
rect 2687 1558 2691 1562
rect 2799 1558 2803 1562
rect 2823 1558 2827 1562
rect 2943 1558 2947 1562
rect 2959 1558 2963 1562
rect 1003 1430 1007 1434
rect 1083 1430 1087 1434
rect 1323 1430 1327 1434
rect 1935 1430 1939 1434
rect 1975 1430 1979 1434
rect 2099 1430 2103 1434
rect 2115 1430 2119 1434
rect 2243 1430 2247 1434
rect 2251 1430 2255 1434
rect 2387 1430 2391 1434
rect 2523 1430 2527 1434
rect 2539 1430 2543 1434
rect 2659 1430 2663 1434
rect 2691 1430 2695 1434
rect 2795 1430 2799 1434
rect 359 1318 363 1322
rect 367 1318 371 1322
rect 583 1318 587 1322
rect 607 1318 611 1322
rect 111 1194 115 1198
rect 131 1194 135 1198
rect 275 1194 279 1198
rect 339 1194 343 1198
rect 443 1194 447 1198
rect 111 1074 115 1078
rect 159 1074 163 1078
rect 175 1074 179 1078
rect 807 1318 811 1322
rect 847 1318 851 1322
rect 1031 1318 1035 1322
rect 1087 1318 1091 1322
rect 1935 1318 1939 1322
rect 3995 1666 3999 1670
rect 4059 1666 4063 1670
rect 4139 1666 4143 1670
rect 4315 1666 4319 1670
rect 4323 1666 4327 1670
rect 3095 1558 3099 1562
rect 3231 1558 3235 1562
rect 3799 1558 3803 1562
rect 3839 1550 3843 1554
rect 3887 1550 3891 1554
rect 2851 1430 2855 1434
rect 2931 1430 2935 1434
rect 3011 1430 3015 1434
rect 3067 1430 3071 1434
rect 3171 1430 3175 1434
rect 3203 1430 3207 1434
rect 4927 1782 4931 1786
rect 5007 1782 5011 1786
rect 5247 1782 5251 1786
rect 5263 1782 5267 1786
rect 5459 1902 5463 1906
rect 5499 1902 5503 1906
rect 5663 2126 5667 2130
rect 5663 2014 5667 2018
rect 5663 1902 5667 1906
rect 5527 1782 5531 1786
rect 5543 1782 5547 1786
rect 4531 1666 4535 1670
rect 4595 1666 4599 1670
rect 4763 1666 4767 1670
rect 4899 1666 4903 1670
rect 5011 1666 5015 1670
rect 5219 1666 5223 1670
rect 5275 1666 5279 1670
rect 5663 1782 5667 1786
rect 5515 1666 5519 1670
rect 4023 1550 4027 1554
rect 4111 1550 4115 1554
rect 4167 1550 4171 1554
rect 4343 1550 4347 1554
rect 4351 1550 4355 1554
rect 4559 1550 4563 1554
rect 4575 1550 4579 1554
rect 4791 1550 4795 1554
rect 4815 1550 4819 1554
rect 5039 1550 5043 1554
rect 5063 1550 5067 1554
rect 3839 1438 3843 1442
rect 3859 1438 3863 1442
rect 4083 1438 4087 1442
rect 3799 1430 3803 1434
rect 3839 1326 3843 1330
rect 3887 1326 3891 1330
rect 1975 1314 1979 1318
rect 2023 1314 2027 1318
rect 2127 1314 2131 1318
rect 2175 1314 2179 1318
rect 2271 1314 2275 1318
rect 2367 1314 2371 1318
rect 2415 1314 2419 1318
rect 2567 1314 2571 1318
rect 2575 1314 2579 1318
rect 2719 1314 2723 1318
rect 2791 1314 2795 1318
rect 2879 1314 2883 1318
rect 3015 1314 3019 1318
rect 579 1194 583 1198
rect 603 1194 607 1198
rect 763 1194 767 1198
rect 819 1194 823 1198
rect 923 1194 927 1198
rect 1059 1194 1063 1198
rect 1075 1194 1079 1198
rect 3039 1314 3043 1318
rect 3199 1314 3203 1318
rect 3239 1314 3243 1318
rect 3471 1314 3475 1318
rect 3679 1314 3683 1318
rect 3799 1314 3803 1318
rect 4315 1438 4319 1442
rect 4323 1438 4327 1442
rect 5303 1550 5307 1554
rect 5311 1550 5315 1554
rect 5663 1666 5667 1670
rect 5543 1550 5547 1554
rect 5663 1550 5667 1554
rect 4547 1438 4551 1442
rect 4771 1438 4775 1442
rect 4787 1438 4791 1442
rect 4987 1438 4991 1442
rect 5035 1438 5039 1442
rect 5203 1438 5207 1442
rect 5283 1438 5287 1442
rect 5419 1438 5423 1442
rect 5515 1438 5519 1442
rect 4111 1326 4115 1330
rect 4119 1326 4123 1330
rect 4351 1326 4355 1330
rect 4391 1326 4395 1330
rect 4575 1326 4579 1330
rect 4671 1326 4675 1330
rect 4799 1326 4803 1330
rect 4967 1326 4971 1330
rect 5015 1326 5019 1330
rect 5231 1326 5235 1330
rect 5263 1326 5267 1330
rect 1219 1194 1223 1198
rect 1363 1194 1367 1198
rect 1507 1194 1511 1198
rect 1651 1194 1655 1198
rect 1787 1194 1791 1198
rect 303 1074 307 1078
rect 111 954 115 958
rect 147 954 151 958
rect 195 954 199 958
rect 415 1074 419 1078
rect 471 1074 475 1078
rect 631 1074 635 1078
rect 639 1074 643 1078
rect 791 1074 795 1078
rect 855 1074 859 1078
rect 387 954 391 958
rect 419 954 423 958
rect 611 954 615 958
rect 667 954 671 958
rect 111 818 115 822
rect 223 818 227 822
rect 951 1074 955 1078
rect 1055 1074 1059 1078
rect 1103 1074 1107 1078
rect 1239 1074 1243 1078
rect 1247 1074 1251 1078
rect 1935 1194 1939 1198
rect 1975 1194 1979 1198
rect 1995 1194 1999 1198
rect 2147 1194 2151 1198
rect 2339 1194 2343 1198
rect 2547 1194 2551 1198
rect 2723 1194 2727 1198
rect 2763 1194 2767 1198
rect 2899 1194 2903 1198
rect 2987 1194 2991 1198
rect 3083 1194 3087 1198
rect 3211 1194 3215 1198
rect 3275 1194 3279 1198
rect 3443 1194 3447 1198
rect 3467 1194 3471 1198
rect 3651 1194 3655 1198
rect 3799 1194 3803 1198
rect 3839 1194 3843 1198
rect 3859 1194 3863 1198
rect 4011 1194 4015 1198
rect 4091 1194 4095 1198
rect 1391 1074 1395 1078
rect 1423 1074 1427 1078
rect 1535 1074 1539 1078
rect 1607 1074 1611 1078
rect 1679 1074 1683 1078
rect 1791 1074 1795 1078
rect 1815 1074 1819 1078
rect 1935 1074 1939 1078
rect 1975 1070 1979 1074
rect 2559 1070 2563 1074
rect 2751 1070 2755 1074
rect 2927 1070 2931 1074
rect 2951 1070 2955 1074
rect 827 954 831 958
rect 931 954 935 958
rect 1027 954 1031 958
rect 1211 954 1215 958
rect 1219 954 1223 958
rect 1395 954 1399 958
rect 1515 954 1519 958
rect 1579 954 1583 958
rect 1763 954 1767 958
rect 1787 954 1791 958
rect 1935 954 1939 958
rect 1975 958 1979 962
rect 1995 958 1999 962
rect 2219 958 2223 962
rect 2467 958 2471 962
rect 2531 958 2535 962
rect 447 818 451 822
rect 663 818 667 822
rect 695 818 699 822
rect 879 818 883 822
rect 959 818 963 822
rect 1087 818 1091 822
rect 1247 818 1251 822
rect 1295 818 1299 822
rect 1511 818 1515 822
rect 1543 818 1547 822
rect 111 698 115 702
rect 131 698 135 702
rect 195 698 199 702
rect 275 698 279 702
rect 419 698 423 702
rect 443 698 447 702
rect 111 574 115 578
rect 159 574 163 578
rect 611 698 615 702
rect 635 698 639 702
rect 771 698 775 702
rect 851 698 855 702
rect 923 698 927 702
rect 1059 698 1063 702
rect 1075 698 1079 702
rect 1975 846 1979 850
rect 2023 846 2027 850
rect 2223 846 2227 850
rect 2247 846 2251 850
rect 1815 818 1819 822
rect 1935 818 1939 822
rect 3111 1070 3115 1074
rect 3151 1070 3155 1074
rect 3303 1070 3307 1074
rect 3359 1070 3363 1074
rect 3495 1070 3499 1074
rect 3575 1070 3579 1074
rect 4211 1194 4215 1198
rect 4363 1194 4367 1198
rect 4435 1194 4439 1198
rect 4643 1194 4647 1198
rect 4691 1194 4695 1198
rect 3679 1070 3683 1074
rect 3799 1070 3803 1074
rect 3839 1070 3843 1074
rect 4039 1070 4043 1074
rect 4095 1070 4099 1074
rect 5447 1326 5451 1330
rect 4939 1194 4943 1198
rect 4963 1194 4967 1198
rect 5235 1194 5239 1198
rect 5251 1194 5255 1198
rect 5515 1194 5519 1198
rect 4239 1070 4243 1074
rect 4391 1070 4395 1074
rect 4463 1070 4467 1074
rect 2707 958 2711 962
rect 2723 958 2727 962
rect 2923 958 2927 962
rect 2939 958 2943 962
rect 3123 958 3127 962
rect 3171 958 3175 962
rect 3331 958 3335 962
rect 3411 958 3415 962
rect 2439 846 2443 850
rect 2495 846 2499 850
rect 2663 846 2667 850
rect 2735 846 2739 850
rect 2887 846 2891 850
rect 2967 846 2971 850
rect 3111 846 3115 850
rect 3199 846 3203 850
rect 3547 958 3551 962
rect 3799 958 3803 962
rect 3839 954 3843 958
rect 3931 954 3935 958
rect 4067 954 4071 958
rect 4155 954 4159 958
rect 3335 846 3339 850
rect 3439 846 3443 850
rect 3559 846 3563 850
rect 3799 846 3803 850
rect 3839 842 3843 846
rect 3887 842 3891 846
rect 3959 842 3963 846
rect 1975 718 1979 722
rect 2195 718 2199 722
rect 2411 718 2415 722
rect 2635 718 2639 722
rect 2859 718 2863 722
rect 3083 718 3087 722
rect 3307 718 3311 722
rect 3379 718 3383 722
rect 1219 698 1223 702
rect 1267 698 1271 702
rect 1363 698 1367 702
rect 1483 698 1487 702
rect 1507 698 1511 702
rect 1651 698 1655 702
rect 1787 698 1791 702
rect 1935 698 1939 702
rect 4363 954 4367 958
rect 4379 954 4383 958
rect 4687 1070 4691 1074
rect 4719 1070 4723 1074
rect 4975 1070 4979 1074
rect 4991 1070 4995 1074
rect 5263 1070 5267 1074
rect 5279 1070 5283 1074
rect 4595 954 4599 958
rect 4659 954 4663 958
rect 4811 954 4815 958
rect 4947 954 4951 958
rect 5027 954 5031 958
rect 5235 954 5239 958
rect 5243 954 5247 958
rect 5467 954 5471 958
rect 5515 954 5519 958
rect 5663 1438 5667 1442
rect 5543 1326 5547 1330
rect 5663 1326 5667 1330
rect 5663 1194 5667 1198
rect 5543 1070 5547 1074
rect 5663 1070 5667 1074
rect 4111 842 4115 846
rect 4183 842 4187 846
rect 4343 842 4347 846
rect 4407 842 4411 846
rect 4575 842 4579 846
rect 4623 842 4627 846
rect 4799 842 4803 846
rect 4839 842 4843 846
rect 3839 730 3843 734
rect 3859 730 3863 734
rect 4083 730 4087 734
rect 3515 718 3519 722
rect 3531 718 3535 722
rect 3651 718 3655 722
rect 3799 718 3803 722
rect 303 574 307 578
rect 375 574 379 578
rect 471 574 475 578
rect 599 574 603 578
rect 639 574 643 578
rect 799 574 803 578
rect 807 574 811 578
rect 951 574 955 578
rect 999 574 1003 578
rect 1103 574 1107 578
rect 1175 574 1179 578
rect 1247 574 1251 578
rect 1343 574 1347 578
rect 1391 574 1395 578
rect 1511 574 1515 578
rect 1535 574 1539 578
rect 1671 574 1675 578
rect 1679 574 1683 578
rect 1815 574 1819 578
rect 111 462 115 466
rect 131 462 135 466
rect 195 462 199 466
rect 347 462 351 466
rect 475 462 479 466
rect 571 462 575 466
rect 755 462 759 466
rect 779 462 783 466
rect 971 462 975 466
rect 1043 462 1047 466
rect 111 350 115 354
rect 223 350 227 354
rect 311 350 315 354
rect 503 350 507 354
rect 1975 598 1979 602
rect 3271 598 3275 602
rect 3407 598 3411 602
rect 3543 598 3547 602
rect 3679 598 3683 602
rect 1935 574 1939 578
rect 3839 610 3843 614
rect 3887 610 3891 614
rect 3799 598 3803 602
rect 4315 730 4319 734
rect 4323 730 4327 734
rect 4547 730 4551 734
rect 4555 730 4559 734
rect 4771 730 4775 734
rect 4779 730 4783 734
rect 5031 842 5035 846
rect 5055 842 5059 846
rect 5263 842 5267 846
rect 5271 842 5275 846
rect 5495 842 5499 846
rect 5663 954 5667 958
rect 5663 842 5667 846
rect 5003 730 5007 734
rect 5227 730 5231 734
rect 5235 730 5239 734
rect 5459 730 5463 734
rect 5467 730 5471 734
rect 5663 730 5667 734
rect 4111 610 4115 614
rect 4143 610 4147 614
rect 4351 610 4355 614
rect 4407 610 4411 614
rect 1147 462 1151 466
rect 1315 462 1319 466
rect 1331 462 1335 466
rect 1483 462 1487 466
rect 1643 462 1647 466
rect 1787 462 1791 466
rect 1935 462 1939 466
rect 1975 466 1979 470
rect 1995 466 1999 470
rect 2155 466 2159 470
rect 2347 466 2351 470
rect 2539 466 2543 470
rect 2739 466 2743 470
rect 2931 466 2935 470
rect 3131 466 3135 470
rect 3243 466 3247 470
rect 3331 466 3335 470
rect 3379 466 3383 470
rect 3515 466 3519 470
rect 3531 466 3535 470
rect 3651 466 3655 470
rect 695 350 699 354
rect 783 350 787 354
rect 111 202 115 206
rect 131 202 135 206
rect 267 202 271 206
rect 283 202 287 206
rect 887 350 891 354
rect 1071 350 1075 354
rect 1079 350 1083 354
rect 1359 350 1363 354
rect 1935 350 1939 354
rect 1975 330 1979 334
rect 2023 330 2027 334
rect 2159 330 2163 334
rect 2183 330 2187 334
rect 2295 330 2299 334
rect 2375 330 2379 334
rect 2431 330 2435 334
rect 2567 330 2571 334
rect 2703 330 2707 334
rect 2767 330 2771 334
rect 2839 330 2843 334
rect 403 202 407 206
rect 475 202 479 206
rect 539 202 543 206
rect 667 202 671 206
rect 675 202 679 206
rect 811 202 815 206
rect 859 202 863 206
rect 947 202 951 206
rect 1051 202 1055 206
rect 1083 202 1087 206
rect 1935 202 1939 206
rect 2115 248 2119 252
rect 1975 186 1979 190
rect 1995 186 1999 190
rect 2959 330 2963 334
rect 2975 330 2979 334
rect 3839 482 3843 486
rect 3859 482 3863 486
rect 3891 482 3895 486
rect 3799 466 3803 470
rect 4583 610 4587 614
rect 4647 610 4651 614
rect 4807 610 4811 614
rect 4879 610 4883 614
rect 5031 610 5035 614
rect 5095 610 5099 614
rect 5255 610 5259 614
rect 5311 610 5315 614
rect 4115 482 4119 486
rect 4171 482 4175 486
rect 4379 482 4383 486
rect 4435 482 4439 486
rect 3839 366 3843 370
rect 3919 366 3923 370
rect 4007 366 4011 370
rect 4199 366 4203 370
rect 4619 482 4623 486
rect 4683 482 4687 486
rect 5487 610 5491 614
rect 5527 610 5531 614
rect 4851 482 4855 486
rect 4907 482 4911 486
rect 5067 482 5071 486
rect 5123 482 5127 486
rect 5283 482 5287 486
rect 5331 482 5335 486
rect 5499 482 5503 486
rect 5515 482 5519 486
rect 4423 366 4427 370
rect 4463 366 4467 370
rect 4679 366 4683 370
rect 4711 366 4715 370
rect 4935 366 4939 370
rect 4967 366 4971 370
rect 5151 366 5155 370
rect 5263 366 5267 370
rect 5359 366 5363 370
rect 5543 366 5547 370
rect 3111 330 3115 334
rect 3159 330 3163 334
rect 3247 330 3251 334
rect 3359 330 3363 334
rect 3383 330 3387 334
rect 3519 330 3523 334
rect 3559 330 3563 334
rect 3799 330 3803 334
rect 2795 248 2799 252
rect 2131 186 2135 190
rect 2267 186 2271 190
rect 2403 186 2407 190
rect 2539 186 2543 190
rect 2675 186 2679 190
rect 2811 186 2815 190
rect 3839 202 3843 206
rect 3859 202 3863 206
rect 3979 202 3983 206
rect 3995 202 3999 206
rect 2947 186 2951 190
rect 3083 186 3087 190
rect 3219 186 3223 190
rect 3355 186 3359 190
rect 3491 186 3495 190
rect 3627 186 3631 190
rect 3799 186 3803 190
rect 2907 176 2911 180
rect 3751 176 3755 180
rect 4131 202 4135 206
rect 4171 202 4175 206
rect 4267 202 4271 206
rect 4395 202 4399 206
rect 4435 202 4439 206
rect 4627 202 4631 206
rect 4651 202 4655 206
rect 5663 610 5667 614
rect 5663 482 5667 486
rect 5663 366 5667 370
rect 4843 202 4847 206
rect 4939 202 4943 206
rect 5067 202 5071 206
rect 5235 202 5239 206
rect 5299 202 5303 206
rect 5515 202 5519 206
rect 5663 202 5667 206
rect 111 90 115 94
rect 159 90 163 94
rect 295 90 299 94
rect 431 90 435 94
rect 567 90 571 94
rect 703 90 707 94
rect 839 90 843 94
rect 975 90 979 94
rect 1111 90 1115 94
rect 1935 90 1939 94
rect 3839 90 3843 94
rect 3887 90 3891 94
rect 4023 90 4027 94
rect 4159 90 4163 94
rect 4295 90 4299 94
rect 4463 90 4467 94
rect 4655 90 4659 94
rect 4871 90 4875 94
rect 5095 90 5099 94
rect 5327 90 5331 94
rect 5543 90 5547 94
rect 5663 90 5667 94
rect 1975 74 1979 78
rect 2023 74 2027 78
rect 2159 74 2163 78
rect 2295 74 2299 78
rect 2431 74 2435 78
rect 2567 74 2571 78
rect 2703 74 2707 78
rect 2839 74 2843 78
rect 2975 74 2979 78
rect 3111 74 3115 78
rect 3247 74 3251 78
rect 3383 74 3387 78
rect 3519 74 3523 78
rect 3655 74 3659 78
rect 3799 74 3803 78
<< m4 >>
rect 96 5753 97 5759
rect 103 5758 1959 5759
rect 103 5754 111 5758
rect 115 5754 131 5758
rect 135 5754 371 5758
rect 375 5754 635 5758
rect 639 5754 907 5758
rect 911 5754 1179 5758
rect 1183 5754 1451 5758
rect 1455 5754 1723 5758
rect 1727 5754 1935 5758
rect 1939 5754 1959 5758
rect 103 5753 1959 5754
rect 1965 5753 1966 5759
rect 1946 5717 1947 5723
rect 1953 5722 3811 5723
rect 1953 5718 1975 5722
rect 1979 5718 2511 5722
rect 2515 5718 2663 5722
rect 2667 5718 2815 5722
rect 2819 5718 2975 5722
rect 2979 5718 3143 5722
rect 3147 5718 3319 5722
rect 3323 5718 3495 5722
rect 3499 5718 3799 5722
rect 3803 5718 3811 5722
rect 1953 5717 3811 5718
rect 3817 5717 3818 5723
rect 3822 5669 3823 5675
rect 3829 5674 5707 5675
rect 3829 5670 3839 5674
rect 3843 5670 4107 5674
rect 4111 5670 4243 5674
rect 4247 5670 4379 5674
rect 4383 5670 4515 5674
rect 4519 5670 4651 5674
rect 4655 5670 4787 5674
rect 4791 5670 4923 5674
rect 4927 5670 5059 5674
rect 5063 5670 5195 5674
rect 5199 5670 5663 5674
rect 5667 5670 5707 5674
rect 3829 5669 5707 5670
rect 5713 5669 5714 5675
rect 84 5641 85 5647
rect 91 5646 1947 5647
rect 91 5642 111 5646
rect 115 5642 159 5646
rect 163 5642 399 5646
rect 403 5642 455 5646
rect 459 5642 647 5646
rect 651 5642 663 5646
rect 667 5642 855 5646
rect 859 5642 935 5646
rect 939 5642 1087 5646
rect 1091 5642 1207 5646
rect 1211 5642 1327 5646
rect 1331 5642 1479 5646
rect 1483 5642 1583 5646
rect 1587 5642 1751 5646
rect 1755 5642 1815 5646
rect 1819 5642 1935 5646
rect 1939 5642 1947 5646
rect 91 5641 1947 5642
rect 1953 5641 1954 5647
rect 1958 5597 1959 5603
rect 1965 5602 3823 5603
rect 1965 5598 1975 5602
rect 1979 5598 1995 5602
rect 1999 5598 2203 5602
rect 2207 5598 2435 5602
rect 2439 5598 2483 5602
rect 2487 5598 2635 5602
rect 2639 5598 2659 5602
rect 2663 5598 2787 5602
rect 2791 5598 2867 5602
rect 2871 5598 2947 5602
rect 2951 5598 3075 5602
rect 3079 5598 3115 5602
rect 3119 5598 3275 5602
rect 3279 5598 3291 5602
rect 3295 5598 3467 5602
rect 3471 5598 3475 5602
rect 3479 5598 3651 5602
rect 3655 5598 3799 5602
rect 3803 5598 3823 5602
rect 1965 5597 3823 5598
rect 3829 5597 3830 5603
rect 882 5564 888 5565
rect 1178 5564 1184 5565
rect 882 5560 883 5564
rect 887 5560 1179 5564
rect 1183 5560 1184 5564
rect 882 5559 888 5560
rect 1178 5559 1184 5560
rect 96 5529 97 5535
rect 103 5534 1959 5535
rect 103 5530 111 5534
rect 115 5530 427 5534
rect 431 5530 619 5534
rect 623 5530 787 5534
rect 791 5530 827 5534
rect 831 5530 923 5534
rect 927 5530 1059 5534
rect 1063 5530 1195 5534
rect 1199 5530 1299 5534
rect 1303 5530 1331 5534
rect 1335 5530 1555 5534
rect 1559 5530 1787 5534
rect 1791 5530 1935 5534
rect 1939 5530 1959 5534
rect 103 5529 1959 5530
rect 1965 5529 1966 5535
rect 3810 5525 3811 5531
rect 3817 5530 5695 5531
rect 3817 5526 3839 5530
rect 3843 5526 4135 5530
rect 4139 5526 4271 5530
rect 4275 5526 4303 5530
rect 4307 5526 4407 5530
rect 4411 5526 4511 5530
rect 4515 5526 4543 5530
rect 4547 5526 4679 5530
rect 4683 5526 4719 5530
rect 4723 5526 4815 5530
rect 4819 5526 4927 5530
rect 4931 5526 4951 5530
rect 4955 5526 5087 5530
rect 5091 5526 5135 5530
rect 5139 5526 5223 5530
rect 5227 5526 5663 5530
rect 5667 5526 5695 5530
rect 3817 5525 5695 5526
rect 5701 5525 5702 5531
rect 1946 5485 1947 5491
rect 1953 5490 3811 5491
rect 1953 5486 1975 5490
rect 1979 5486 2023 5490
rect 2027 5486 2167 5490
rect 2171 5486 2231 5490
rect 2235 5486 2343 5490
rect 2347 5486 2463 5490
rect 2467 5486 2527 5490
rect 2531 5486 2687 5490
rect 2691 5486 2719 5490
rect 2723 5486 2895 5490
rect 2899 5486 2911 5490
rect 2915 5486 3103 5490
rect 3107 5486 3111 5490
rect 3115 5486 3303 5490
rect 3307 5486 3311 5490
rect 3315 5486 3503 5490
rect 3507 5486 3679 5490
rect 3683 5486 3799 5490
rect 3803 5486 3811 5490
rect 1953 5485 3811 5486
rect 3817 5485 3818 5491
rect 84 5397 85 5403
rect 91 5402 1947 5403
rect 91 5398 111 5402
rect 115 5398 815 5402
rect 819 5398 903 5402
rect 907 5398 951 5402
rect 955 5398 1039 5402
rect 1043 5398 1087 5402
rect 1091 5398 1183 5402
rect 1187 5398 1223 5402
rect 1227 5398 1335 5402
rect 1339 5398 1359 5402
rect 1363 5398 1495 5402
rect 1499 5398 1663 5402
rect 1667 5398 1815 5402
rect 1819 5398 1935 5402
rect 1939 5398 1947 5402
rect 91 5397 1947 5398
rect 1953 5397 1954 5403
rect 3822 5389 3823 5395
rect 3829 5394 5707 5395
rect 3829 5390 3839 5394
rect 3843 5390 3859 5394
rect 3863 5390 3995 5394
rect 3999 5390 4131 5394
rect 4135 5390 4275 5394
rect 4279 5390 4435 5394
rect 4439 5390 4483 5394
rect 4487 5390 4603 5394
rect 4607 5390 4691 5394
rect 4695 5390 4779 5394
rect 4783 5390 4899 5394
rect 4903 5390 4963 5394
rect 4967 5390 5107 5394
rect 5111 5390 5663 5394
rect 5667 5390 5707 5394
rect 3829 5389 5707 5390
rect 5713 5389 5714 5395
rect 1958 5349 1959 5355
rect 1965 5354 3823 5355
rect 1965 5350 1975 5354
rect 1979 5350 1995 5354
rect 1999 5350 2051 5354
rect 2055 5350 2139 5354
rect 2143 5350 2315 5354
rect 2319 5350 2459 5354
rect 2463 5350 2499 5354
rect 2503 5350 2691 5354
rect 2695 5350 2859 5354
rect 2863 5350 2883 5354
rect 2887 5350 3083 5354
rect 3087 5350 3267 5354
rect 3271 5350 3283 5354
rect 3287 5350 3651 5354
rect 3655 5350 3799 5354
rect 3803 5350 3823 5354
rect 1965 5349 3823 5350
rect 3829 5349 3830 5355
rect 96 5281 97 5287
rect 103 5286 1959 5287
rect 103 5282 111 5286
rect 115 5282 587 5286
rect 591 5282 739 5286
rect 743 5282 875 5286
rect 879 5282 899 5286
rect 903 5282 1011 5286
rect 1015 5282 1067 5286
rect 1071 5282 1155 5286
rect 1159 5282 1243 5286
rect 1247 5282 1307 5286
rect 1311 5282 1427 5286
rect 1431 5282 1467 5286
rect 1471 5282 1619 5286
rect 1623 5282 1635 5286
rect 1639 5282 1787 5286
rect 1791 5282 1935 5286
rect 1939 5282 1959 5286
rect 103 5281 1959 5282
rect 1965 5281 1966 5287
rect 3810 5273 3811 5279
rect 3817 5278 5695 5279
rect 3817 5274 3839 5278
rect 3843 5274 3887 5278
rect 3891 5274 3999 5278
rect 4003 5274 4023 5278
rect 4027 5274 4159 5278
rect 4163 5274 4199 5278
rect 4203 5274 4303 5278
rect 4307 5274 4399 5278
rect 4403 5274 4463 5278
rect 4467 5274 4607 5278
rect 4611 5274 4631 5278
rect 4635 5274 4807 5278
rect 4811 5274 4823 5278
rect 4827 5274 4991 5278
rect 4995 5274 5039 5278
rect 5043 5274 5663 5278
rect 5667 5274 5695 5278
rect 3817 5273 5695 5274
rect 5701 5273 5702 5279
rect 1946 5237 1947 5243
rect 1953 5242 3811 5243
rect 1953 5238 1975 5242
rect 1979 5238 2079 5242
rect 2083 5238 2239 5242
rect 2243 5238 2487 5242
rect 2491 5238 2591 5242
rect 2595 5238 2887 5242
rect 2891 5238 2943 5242
rect 2947 5238 3295 5242
rect 3299 5238 3303 5242
rect 3307 5238 3663 5242
rect 3667 5238 3679 5242
rect 3683 5238 3799 5242
rect 3803 5238 3811 5242
rect 1953 5237 3811 5238
rect 3817 5237 3818 5243
rect 84 5157 85 5163
rect 91 5162 1947 5163
rect 91 5158 111 5162
rect 115 5158 367 5162
rect 371 5158 535 5162
rect 539 5158 615 5162
rect 619 5158 711 5162
rect 715 5158 767 5162
rect 771 5158 895 5162
rect 899 5158 927 5162
rect 931 5158 1079 5162
rect 1083 5158 1095 5162
rect 1099 5158 1263 5162
rect 1267 5158 1271 5162
rect 1275 5158 1447 5162
rect 1451 5158 1455 5162
rect 1459 5158 1631 5162
rect 1635 5158 1647 5162
rect 1651 5158 1815 5162
rect 1819 5158 1935 5162
rect 1939 5158 1947 5162
rect 91 5157 1947 5158
rect 1953 5157 1954 5163
rect 3822 5141 3823 5147
rect 3829 5146 5707 5147
rect 3829 5142 3839 5146
rect 3843 5142 3971 5146
rect 3975 5142 4099 5146
rect 4103 5142 4171 5146
rect 4175 5142 4347 5146
rect 4351 5142 4371 5146
rect 4375 5142 4579 5146
rect 4583 5142 4595 5146
rect 4599 5142 4795 5146
rect 4799 5142 4843 5146
rect 4847 5142 5011 5146
rect 5015 5142 5099 5146
rect 5103 5142 5663 5146
rect 5667 5142 5707 5146
rect 3829 5141 5707 5142
rect 5713 5141 5714 5147
rect 1958 5125 1959 5131
rect 1965 5130 3823 5131
rect 1965 5126 1975 5130
rect 1979 5126 2211 5130
rect 2215 5126 2267 5130
rect 2271 5126 2515 5130
rect 2519 5126 2563 5130
rect 2567 5126 2755 5130
rect 2759 5126 2915 5130
rect 2919 5126 2995 5130
rect 2999 5126 3235 5130
rect 3239 5126 3275 5130
rect 3279 5126 3475 5130
rect 3479 5126 3635 5130
rect 3639 5126 3799 5130
rect 3803 5126 3823 5130
rect 1965 5125 3823 5126
rect 3829 5125 3830 5131
rect 96 5041 97 5047
rect 103 5046 1959 5047
rect 103 5042 111 5046
rect 115 5042 131 5046
rect 135 5042 323 5046
rect 327 5042 339 5046
rect 343 5042 507 5046
rect 511 5042 555 5046
rect 559 5042 683 5046
rect 687 5042 811 5046
rect 815 5042 867 5046
rect 871 5042 1051 5046
rect 1055 5042 1083 5046
rect 1087 5042 1235 5046
rect 1239 5042 1371 5046
rect 1375 5042 1419 5046
rect 1423 5042 1603 5046
rect 1607 5042 1659 5046
rect 1663 5042 1787 5046
rect 1791 5042 1935 5046
rect 1939 5042 1959 5046
rect 103 5041 1959 5042
rect 1965 5041 1966 5047
rect 3810 5013 3811 5019
rect 3817 5018 5695 5019
rect 3817 5014 3839 5018
rect 3843 5014 3983 5018
rect 3987 5014 4127 5018
rect 4131 5014 4223 5018
rect 4227 5014 4375 5018
rect 4379 5014 4447 5018
rect 4451 5014 4623 5018
rect 4627 5014 4655 5018
rect 4659 5014 4855 5018
rect 4859 5014 4871 5018
rect 4875 5014 5039 5018
rect 5043 5014 5127 5018
rect 5131 5014 5215 5018
rect 5219 5014 5391 5018
rect 5395 5014 5543 5018
rect 5547 5014 5663 5018
rect 5667 5014 5695 5018
rect 3817 5013 5695 5014
rect 5701 5013 5702 5019
rect 1946 4981 1947 4987
rect 1953 4986 3811 4987
rect 1953 4982 1975 4986
rect 1979 4982 2183 4986
rect 2187 4982 2295 4986
rect 2299 4982 2319 4986
rect 2323 4982 2455 4986
rect 2459 4982 2543 4986
rect 2547 4982 2599 4986
rect 2603 4982 2743 4986
rect 2747 4982 2783 4986
rect 2787 4982 2895 4986
rect 2899 4982 3023 4986
rect 3027 4982 3047 4986
rect 3051 4982 3199 4986
rect 3203 4982 3263 4986
rect 3267 4982 3351 4986
rect 3355 4982 3503 4986
rect 3507 4982 3799 4986
rect 3803 4982 3811 4986
rect 1953 4981 3811 4982
rect 3817 4981 3818 4987
rect 84 4905 85 4911
rect 91 4910 1947 4911
rect 91 4906 111 4910
rect 115 4906 159 4910
rect 163 4906 295 4910
rect 299 4906 351 4910
rect 355 4906 431 4910
rect 435 4906 567 4910
rect 571 4906 583 4910
rect 587 4906 703 4910
rect 707 4906 839 4910
rect 843 4906 1111 4910
rect 1115 4906 1399 4910
rect 1403 4906 1687 4910
rect 1691 4906 1935 4910
rect 1939 4906 1947 4910
rect 91 4905 1947 4906
rect 1953 4905 1954 4911
rect 3822 4877 3823 4883
rect 3829 4882 5707 4883
rect 3829 4878 3839 4882
rect 3843 4878 3859 4882
rect 3863 4878 3955 4882
rect 3959 4878 4075 4882
rect 4079 4878 4195 4882
rect 4199 4878 4299 4882
rect 4303 4878 4419 4882
rect 4423 4878 4507 4882
rect 4511 4878 4627 4882
rect 4631 4878 4699 4882
rect 4703 4878 4827 4882
rect 4831 4878 4875 4882
rect 4879 4878 5011 4882
rect 5015 4878 5043 4882
rect 5047 4878 5187 4882
rect 5191 4878 5211 4882
rect 5215 4878 5363 4882
rect 5367 4878 5371 4882
rect 5375 4878 5515 4882
rect 5519 4878 5663 4882
rect 5667 4878 5707 4882
rect 3829 4877 5707 4878
rect 5713 4877 5714 4883
rect 1958 4861 1959 4867
rect 1965 4866 3823 4867
rect 1965 4862 1975 4866
rect 1979 4862 2155 4866
rect 2159 4862 2291 4866
rect 2295 4862 2427 4866
rect 2431 4862 2571 4866
rect 2575 4862 2715 4866
rect 2719 4862 2723 4866
rect 2727 4862 2867 4866
rect 2871 4862 2875 4866
rect 2879 4862 3019 4866
rect 3023 4862 3027 4866
rect 3031 4862 3171 4866
rect 3175 4862 3179 4866
rect 3183 4862 3323 4866
rect 3327 4862 3799 4866
rect 3803 4862 3823 4866
rect 1965 4861 3823 4862
rect 3829 4861 3830 4867
rect 96 4781 97 4787
rect 103 4786 1959 4787
rect 103 4782 111 4786
rect 115 4782 131 4786
rect 135 4782 267 4786
rect 271 4782 403 4786
rect 407 4782 539 4786
rect 543 4782 675 4786
rect 679 4782 1935 4786
rect 1939 4782 1959 4786
rect 103 4781 1959 4782
rect 1965 4781 1966 4787
rect 3810 4765 3811 4771
rect 3817 4770 5695 4771
rect 3817 4766 3839 4770
rect 3843 4766 3887 4770
rect 3891 4766 4103 4770
rect 4107 4766 4327 4770
rect 4331 4766 4535 4770
rect 4539 4766 4727 4770
rect 4731 4766 4903 4770
rect 4907 4766 4943 4770
rect 4947 4766 5071 4770
rect 5075 4766 5087 4770
rect 5091 4766 5239 4770
rect 5243 4766 5399 4770
rect 5403 4766 5543 4770
rect 5547 4766 5663 4770
rect 5667 4766 5695 4770
rect 3817 4765 5695 4766
rect 5701 4765 5702 4771
rect 1946 4745 1947 4751
rect 1953 4750 3811 4751
rect 1953 4746 1975 4750
rect 1979 4746 2023 4750
rect 2027 4746 2159 4750
rect 2163 4746 2295 4750
rect 2299 4746 2431 4750
rect 2435 4746 2455 4750
rect 2459 4746 2567 4750
rect 2571 4746 2599 4750
rect 2603 4746 2703 4750
rect 2707 4746 2751 4750
rect 2755 4746 2839 4750
rect 2843 4746 2903 4750
rect 2907 4746 2975 4750
rect 2979 4746 3055 4750
rect 3059 4746 3111 4750
rect 3115 4746 3207 4750
rect 3211 4746 3247 4750
rect 3251 4746 3399 4750
rect 3403 4746 3543 4750
rect 3547 4746 3679 4750
rect 3683 4746 3799 4750
rect 3803 4746 3811 4750
rect 1953 4745 3811 4746
rect 3817 4745 3818 4751
rect 84 4661 85 4667
rect 91 4666 1947 4667
rect 91 4662 111 4666
rect 115 4662 159 4666
rect 163 4662 295 4666
rect 299 4662 431 4666
rect 435 4662 567 4666
rect 571 4662 703 4666
rect 707 4662 1935 4666
rect 1939 4662 1947 4666
rect 91 4661 1947 4662
rect 1953 4661 1954 4667
rect 3822 4629 3823 4635
rect 3829 4634 5707 4635
rect 3829 4630 3839 4634
rect 3843 4630 4771 4634
rect 4775 4630 4915 4634
rect 4919 4630 4955 4634
rect 4959 4630 5059 4634
rect 5063 4630 5147 4634
rect 5151 4630 5211 4634
rect 5215 4630 5339 4634
rect 5343 4630 5371 4634
rect 5375 4630 5515 4634
rect 5519 4630 5663 4634
rect 5667 4630 5707 4634
rect 3829 4629 5707 4630
rect 5713 4629 5714 4635
rect 1958 4601 1959 4607
rect 1965 4606 3823 4607
rect 1965 4602 1975 4606
rect 1979 4602 1995 4606
rect 1999 4602 2131 4606
rect 2135 4602 2267 4606
rect 2271 4602 2323 4606
rect 2327 4602 2403 4606
rect 2407 4602 2539 4606
rect 2543 4602 2579 4606
rect 2583 4602 2675 4606
rect 2679 4602 2811 4606
rect 2815 4602 2827 4606
rect 2831 4602 2947 4606
rect 2951 4602 3075 4606
rect 3079 4602 3083 4606
rect 3087 4602 3219 4606
rect 3223 4602 3315 4606
rect 3319 4602 3371 4606
rect 3375 4602 3515 4606
rect 3519 4602 3563 4606
rect 3567 4602 3651 4606
rect 3655 4602 3799 4606
rect 3803 4602 3823 4606
rect 1965 4601 3823 4602
rect 3829 4601 3830 4607
rect 4866 4572 4872 4573
rect 5422 4572 5428 4573
rect 4866 4568 4867 4572
rect 4871 4568 5423 4572
rect 5427 4568 5428 4572
rect 4866 4567 4872 4568
rect 5422 4567 5428 4568
rect 96 4541 97 4547
rect 103 4546 1959 4547
rect 103 4542 111 4546
rect 115 4542 131 4546
rect 135 4542 267 4546
rect 271 4542 339 4546
rect 343 4542 403 4546
rect 407 4542 515 4546
rect 519 4542 539 4546
rect 543 4542 675 4546
rect 679 4542 691 4546
rect 695 4542 875 4546
rect 879 4542 1059 4546
rect 1063 4542 1243 4546
rect 1247 4542 1427 4546
rect 1431 4542 1619 4546
rect 1623 4542 1787 4546
rect 1791 4542 1935 4546
rect 1939 4542 1959 4546
rect 103 4541 1959 4542
rect 1965 4541 1966 4547
rect 3810 4505 3811 4511
rect 3817 4510 5695 4511
rect 3817 4506 3839 4510
rect 3843 4506 4487 4510
rect 4491 4506 4671 4510
rect 4675 4506 4799 4510
rect 4803 4506 4879 4510
rect 4883 4506 4983 4510
rect 4987 4506 5095 4510
rect 5099 4506 5175 4510
rect 5179 4506 5327 4510
rect 5331 4506 5367 4510
rect 5371 4506 5543 4510
rect 5547 4506 5663 4510
rect 5667 4506 5695 4510
rect 3817 4505 5695 4506
rect 5701 4505 5702 4511
rect 1946 4481 1947 4487
rect 1953 4486 3811 4487
rect 1953 4482 1975 4486
rect 1979 4482 2351 4486
rect 2355 4482 2543 4486
rect 2547 4482 2607 4486
rect 2611 4482 2783 4486
rect 2787 4482 2855 4486
rect 2859 4482 3015 4486
rect 3019 4482 3103 4486
rect 3107 4482 3247 4486
rect 3251 4482 3343 4486
rect 3347 4482 3471 4486
rect 3475 4482 3591 4486
rect 3595 4482 3679 4486
rect 3683 4482 3799 4486
rect 3803 4482 3811 4486
rect 1953 4481 3811 4482
rect 3817 4481 3818 4487
rect 84 4429 85 4435
rect 91 4434 1947 4435
rect 91 4430 111 4434
rect 115 4430 367 4434
rect 371 4430 543 4434
rect 547 4430 567 4434
rect 571 4430 711 4434
rect 715 4430 719 4434
rect 723 4430 863 4434
rect 867 4430 903 4434
rect 907 4430 1023 4434
rect 1027 4430 1087 4434
rect 1091 4430 1183 4434
rect 1187 4430 1271 4434
rect 1275 4430 1343 4434
rect 1347 4430 1455 4434
rect 1459 4430 1503 4434
rect 1507 4430 1647 4434
rect 1651 4430 1671 4434
rect 1675 4430 1815 4434
rect 1819 4430 1935 4434
rect 1939 4430 1947 4434
rect 91 4429 1947 4430
rect 1953 4429 1954 4435
rect 3822 4369 3823 4375
rect 3829 4374 5707 4375
rect 3829 4370 3839 4374
rect 3843 4370 3859 4374
rect 3863 4370 3995 4374
rect 3999 4370 4131 4374
rect 4135 4370 4283 4374
rect 4287 4370 4459 4374
rect 4463 4370 4483 4374
rect 4487 4370 4643 4374
rect 4647 4370 4715 4374
rect 4719 4370 4851 4374
rect 4855 4370 4979 4374
rect 4983 4370 5067 4374
rect 5071 4370 5251 4374
rect 5255 4370 5299 4374
rect 5303 4370 5515 4374
rect 5519 4370 5663 4374
rect 5667 4370 5707 4374
rect 3829 4369 5707 4370
rect 5713 4369 5714 4375
rect 1958 4357 1959 4363
rect 1965 4362 3823 4363
rect 1965 4358 1975 4362
rect 1979 4358 1995 4362
rect 1999 4358 2379 4362
rect 2383 4358 2515 4362
rect 2519 4358 2755 4362
rect 2759 4358 2803 4362
rect 2807 4358 2987 4362
rect 2991 4358 3219 4362
rect 3223 4358 3235 4362
rect 3239 4358 3443 4362
rect 3447 4358 3651 4362
rect 3655 4358 3799 4362
rect 3803 4358 3823 4362
rect 1965 4357 3823 4358
rect 3829 4357 3830 4363
rect 96 4297 97 4303
rect 103 4302 1959 4303
rect 103 4298 111 4302
rect 115 4298 539 4302
rect 543 4298 627 4302
rect 631 4298 683 4302
rect 687 4298 771 4302
rect 775 4298 835 4302
rect 839 4298 923 4302
rect 927 4298 995 4302
rect 999 4298 1083 4302
rect 1087 4298 1155 4302
rect 1159 4298 1251 4302
rect 1255 4298 1315 4302
rect 1319 4298 1419 4302
rect 1423 4298 1475 4302
rect 1479 4298 1595 4302
rect 1599 4298 1643 4302
rect 1647 4298 1787 4302
rect 1791 4298 1935 4302
rect 1939 4298 1959 4302
rect 103 4297 1959 4298
rect 1965 4297 1966 4303
rect 4378 4276 4384 4277
rect 5366 4276 5372 4277
rect 4378 4272 4379 4276
rect 4383 4272 5367 4276
rect 5371 4272 5372 4276
rect 4378 4271 4384 4272
rect 5366 4271 5372 4272
rect 3810 4257 3811 4263
rect 3817 4262 5695 4263
rect 3817 4258 3839 4262
rect 3843 4258 3887 4262
rect 3891 4258 4023 4262
rect 4027 4258 4159 4262
rect 4163 4258 4303 4262
rect 4307 4258 4311 4262
rect 4315 4258 4503 4262
rect 4507 4258 4511 4262
rect 4515 4258 4735 4262
rect 4739 4258 4743 4262
rect 4747 4258 4999 4262
rect 5003 4258 5007 4262
rect 5011 4258 5271 4262
rect 5275 4258 5279 4262
rect 5283 4258 5543 4262
rect 5547 4258 5663 4262
rect 5667 4258 5695 4262
rect 3817 4257 5695 4258
rect 5701 4257 5702 4263
rect 1946 4217 1947 4223
rect 1953 4222 3811 4223
rect 1953 4218 1975 4222
rect 1979 4218 2023 4222
rect 2027 4218 2191 4222
rect 2195 4218 2383 4222
rect 2387 4218 2407 4222
rect 2411 4218 2583 4222
rect 2587 4218 2783 4222
rect 2787 4218 2831 4222
rect 2835 4218 2983 4222
rect 2987 4218 3263 4222
rect 3267 4218 3679 4222
rect 3683 4218 3799 4222
rect 3803 4218 3811 4222
rect 1953 4217 3811 4218
rect 3817 4217 3818 4223
rect 84 4181 85 4187
rect 91 4186 1947 4187
rect 91 4182 111 4186
rect 115 4182 519 4186
rect 523 4182 655 4186
rect 659 4182 703 4186
rect 707 4182 799 4186
rect 803 4182 895 4186
rect 899 4182 951 4186
rect 955 4182 1103 4186
rect 1107 4182 1111 4186
rect 1115 4182 1279 4186
rect 1283 4182 1327 4186
rect 1331 4182 1447 4186
rect 1451 4182 1551 4186
rect 1555 4182 1623 4186
rect 1627 4182 1783 4186
rect 1787 4182 1935 4186
rect 1939 4182 1947 4186
rect 91 4181 1947 4182
rect 1953 4181 1954 4187
rect 1958 4105 1959 4111
rect 1965 4110 3823 4111
rect 1965 4106 1975 4110
rect 1979 4106 1995 4110
rect 1999 4106 2075 4110
rect 2079 4106 2163 4110
rect 2167 4106 2259 4110
rect 2263 4106 2355 4110
rect 2359 4106 2443 4110
rect 2447 4106 2555 4110
rect 2559 4106 2619 4110
rect 2623 4106 2755 4110
rect 2759 4106 2787 4110
rect 2791 4106 2955 4110
rect 2959 4106 3131 4110
rect 3135 4106 3799 4110
rect 3803 4106 3823 4110
rect 1965 4105 3823 4106
rect 3829 4110 5714 4111
rect 3829 4106 3839 4110
rect 3843 4106 3859 4110
rect 3863 4106 3995 4110
rect 3999 4106 4131 4110
rect 4135 4106 4275 4110
rect 4279 4106 4475 4110
rect 4479 4106 4563 4110
rect 4567 4106 4699 4110
rect 4703 4106 4707 4110
rect 4711 4106 4835 4110
rect 4839 4106 4971 4110
rect 4975 4106 5107 4110
rect 5111 4106 5243 4110
rect 5247 4106 5379 4110
rect 5383 4106 5515 4110
rect 5519 4106 5663 4110
rect 5667 4106 5714 4110
rect 3829 4105 5714 4106
rect 96 4069 97 4075
rect 103 4074 1959 4075
rect 103 4070 111 4074
rect 115 4070 131 4074
rect 135 4070 339 4074
rect 343 4070 491 4074
rect 495 4070 595 4074
rect 599 4070 675 4074
rect 679 4070 867 4074
rect 871 4070 875 4074
rect 879 4070 1075 4074
rect 1079 4070 1179 4074
rect 1183 4070 1299 4074
rect 1303 4070 1491 4074
rect 1495 4070 1523 4074
rect 1527 4070 1755 4074
rect 1759 4070 1787 4074
rect 1791 4070 1935 4074
rect 1939 4070 1959 4074
rect 103 4069 1959 4070
rect 1965 4069 1966 4075
rect 1946 3985 1947 3991
rect 1953 3990 3811 3991
rect 1953 3986 1975 3990
rect 1979 3986 2103 3990
rect 2107 3986 2127 3990
rect 2131 3986 2287 3990
rect 2291 3986 2311 3990
rect 2315 3986 2471 3990
rect 2475 3986 2487 3990
rect 2491 3986 2647 3990
rect 2651 3986 2663 3990
rect 2667 3986 2815 3990
rect 2819 3986 2831 3990
rect 2835 3986 2983 3990
rect 2987 3986 2999 3990
rect 3003 3986 3159 3990
rect 3163 3986 3175 3990
rect 3179 3986 3351 3990
rect 3355 3986 3799 3990
rect 3803 3986 3811 3990
rect 1953 3985 3811 3986
rect 3817 3985 3818 3991
rect 3810 3973 3811 3979
rect 3817 3978 5695 3979
rect 3817 3974 3839 3978
rect 3843 3974 4359 3978
rect 4363 3974 4543 3978
rect 4547 3974 4591 3978
rect 4595 3974 4727 3978
rect 4731 3974 4735 3978
rect 4739 3974 4863 3978
rect 4867 3974 4927 3978
rect 4931 3974 4999 3978
rect 5003 3974 5127 3978
rect 5131 3974 5135 3978
rect 5139 3974 5271 3978
rect 5275 3974 5327 3978
rect 5331 3974 5407 3978
rect 5411 3974 5527 3978
rect 5531 3974 5543 3978
rect 5547 3974 5663 3978
rect 5667 3974 5695 3978
rect 3817 3973 5695 3974
rect 5701 3973 5702 3979
rect 84 3953 85 3959
rect 91 3958 1947 3959
rect 91 3954 111 3958
rect 115 3954 159 3958
rect 163 3954 343 3958
rect 347 3954 367 3958
rect 371 3954 567 3958
rect 571 3954 623 3958
rect 627 3954 807 3958
rect 811 3954 903 3958
rect 907 3954 1055 3958
rect 1059 3954 1207 3958
rect 1211 3954 1311 3958
rect 1315 3954 1519 3958
rect 1523 3954 1575 3958
rect 1579 3954 1815 3958
rect 1819 3954 1935 3958
rect 1939 3954 1947 3958
rect 91 3953 1947 3954
rect 1953 3953 1954 3959
rect 1958 3865 1959 3871
rect 1965 3870 3823 3871
rect 1965 3866 1975 3870
rect 1979 3866 2099 3870
rect 2103 3866 2283 3870
rect 2287 3866 2291 3870
rect 2295 3866 2459 3870
rect 2463 3866 2523 3870
rect 2527 3866 2635 3870
rect 2639 3866 2739 3870
rect 2743 3866 2803 3870
rect 2807 3866 2947 3870
rect 2951 3866 2971 3870
rect 2975 3866 3147 3870
rect 3151 3866 3155 3870
rect 3159 3866 3323 3870
rect 3327 3866 3355 3870
rect 3359 3866 3563 3870
rect 3567 3866 3799 3870
rect 3803 3866 3823 3870
rect 1965 3865 3823 3866
rect 3829 3865 3830 3871
rect 3822 3853 3823 3859
rect 3829 3858 5707 3859
rect 3829 3854 3839 3858
rect 3843 3854 4051 3858
rect 4055 3854 4267 3858
rect 4271 3854 4331 3858
rect 4335 3854 4483 3858
rect 4487 3854 4515 3858
rect 4519 3854 4699 3858
rect 4703 3854 4707 3858
rect 4711 3854 4899 3858
rect 4903 3854 4907 3858
rect 4911 3854 5099 3858
rect 5103 3854 5115 3858
rect 5119 3854 5299 3858
rect 5303 3854 5323 3858
rect 5327 3854 5499 3858
rect 5503 3854 5515 3858
rect 5519 3854 5663 3858
rect 5667 3854 5707 3858
rect 3829 3853 5707 3854
rect 5713 3853 5714 3859
rect 96 3833 97 3839
rect 103 3838 1959 3839
rect 103 3834 111 3838
rect 115 3834 131 3838
rect 135 3834 267 3838
rect 271 3834 315 3838
rect 319 3834 475 3838
rect 479 3834 539 3838
rect 543 3834 707 3838
rect 711 3834 779 3838
rect 783 3834 963 3838
rect 967 3834 1027 3838
rect 1031 3834 1235 3838
rect 1239 3834 1283 3838
rect 1287 3834 1515 3838
rect 1519 3834 1547 3838
rect 1551 3834 1787 3838
rect 1791 3834 1935 3838
rect 1939 3834 1959 3838
rect 103 3833 1959 3834
rect 1965 3833 1966 3839
rect 1946 3749 1947 3755
rect 1953 3754 3811 3755
rect 1953 3750 1975 3754
rect 1979 3750 2319 3754
rect 2323 3750 2407 3754
rect 2411 3750 2551 3754
rect 2555 3750 2647 3754
rect 2651 3750 2767 3754
rect 2771 3750 2871 3754
rect 2875 3750 2975 3754
rect 2979 3750 3087 3754
rect 3091 3750 3183 3754
rect 3187 3750 3295 3754
rect 3299 3750 3383 3754
rect 3387 3750 3495 3754
rect 3499 3750 3591 3754
rect 3595 3750 3679 3754
rect 3683 3750 3799 3754
rect 3803 3750 3811 3754
rect 1953 3749 3811 3750
rect 3817 3749 3818 3755
rect 84 3717 85 3723
rect 91 3722 1947 3723
rect 91 3718 111 3722
rect 115 3718 295 3722
rect 299 3718 503 3722
rect 507 3718 631 3722
rect 635 3718 735 3722
rect 739 3718 775 3722
rect 779 3718 927 3722
rect 931 3718 991 3722
rect 995 3718 1087 3722
rect 1091 3718 1255 3722
rect 1259 3718 1263 3722
rect 1267 3718 1423 3722
rect 1427 3718 1543 3722
rect 1547 3718 1591 3722
rect 1595 3718 1759 3722
rect 1763 3718 1815 3722
rect 1819 3718 1935 3722
rect 1939 3718 1947 3722
rect 91 3717 1947 3718
rect 1953 3717 1954 3723
rect 3810 3713 3811 3719
rect 3817 3718 5695 3719
rect 3817 3714 3839 3718
rect 3843 3714 3887 3718
rect 3891 3714 4055 3718
rect 4059 3714 4079 3718
rect 4083 3714 4247 3718
rect 4251 3714 4295 3718
rect 4299 3714 4439 3718
rect 4443 3714 4511 3718
rect 4515 3714 4631 3718
rect 4635 3714 4727 3718
rect 4731 3714 4935 3718
rect 4939 3714 5143 3718
rect 5147 3714 5351 3718
rect 5355 3714 5543 3718
rect 5547 3714 5663 3718
rect 5667 3714 5695 3718
rect 3817 3713 5695 3714
rect 5701 3713 5702 3719
rect 1958 3629 1959 3635
rect 1965 3634 3823 3635
rect 1965 3630 1975 3634
rect 1979 3630 2379 3634
rect 2383 3630 2411 3634
rect 2415 3630 2547 3634
rect 2551 3630 2619 3634
rect 2623 3630 2683 3634
rect 2687 3630 2843 3634
rect 2847 3630 3059 3634
rect 3063 3630 3267 3634
rect 3271 3630 3467 3634
rect 3471 3630 3651 3634
rect 3655 3630 3799 3634
rect 3803 3630 3823 3634
rect 1965 3629 3823 3630
rect 3829 3629 3830 3635
rect 3822 3601 3823 3607
rect 3829 3606 5707 3607
rect 3829 3602 3839 3606
rect 3843 3602 3859 3606
rect 3863 3602 3995 3606
rect 3999 3602 4027 3606
rect 4031 3602 4131 3606
rect 4135 3602 4219 3606
rect 4223 3602 4267 3606
rect 4271 3602 4403 3606
rect 4407 3602 4411 3606
rect 4415 3602 4539 3606
rect 4543 3602 4603 3606
rect 4607 3602 4675 3606
rect 4679 3602 4811 3606
rect 4815 3602 4947 3606
rect 4951 3602 5083 3606
rect 5087 3602 5663 3606
rect 5667 3602 5707 3606
rect 3829 3601 5707 3602
rect 5713 3601 5714 3607
rect 96 3593 97 3599
rect 103 3598 1959 3599
rect 103 3594 111 3598
rect 115 3594 603 3598
rect 607 3594 747 3598
rect 751 3594 779 3598
rect 783 3594 899 3598
rect 903 3594 915 3598
rect 919 3594 1051 3598
rect 1055 3594 1059 3598
rect 1063 3594 1187 3598
rect 1191 3594 1227 3598
rect 1231 3594 1323 3598
rect 1327 3594 1395 3598
rect 1399 3594 1459 3598
rect 1463 3594 1563 3598
rect 1567 3594 1595 3598
rect 1599 3594 1731 3598
rect 1735 3594 1935 3598
rect 1939 3594 1959 3598
rect 103 3593 1959 3594
rect 1965 3593 1966 3599
rect 3954 3596 3960 3597
rect 4526 3596 4532 3597
rect 3954 3592 3955 3596
rect 3959 3592 4527 3596
rect 4531 3592 4532 3596
rect 3954 3591 3960 3592
rect 4526 3591 4532 3592
rect 3810 3486 5702 3487
rect 3810 3483 3839 3486
rect 1946 3477 1947 3483
rect 1953 3482 3811 3483
rect 1953 3478 1975 3482
rect 1979 3478 2439 3482
rect 2443 3478 2575 3482
rect 2579 3478 2599 3482
rect 2603 3478 2711 3482
rect 2715 3478 2823 3482
rect 2827 3478 3047 3482
rect 3051 3478 3263 3482
rect 3267 3478 3479 3482
rect 3483 3478 3679 3482
rect 3683 3478 3799 3482
rect 3803 3478 3811 3482
rect 1953 3477 3811 3478
rect 3817 3482 3839 3483
rect 3843 3482 3887 3486
rect 3891 3482 4023 3486
rect 4027 3482 4159 3486
rect 4163 3482 4295 3486
rect 4299 3482 4431 3486
rect 4435 3482 4567 3486
rect 4571 3482 4703 3486
rect 4707 3482 4831 3486
rect 4835 3482 4839 3486
rect 4843 3482 4967 3486
rect 4971 3482 4975 3486
rect 4979 3482 5103 3486
rect 5107 3482 5111 3486
rect 5115 3482 5239 3486
rect 5243 3482 5375 3486
rect 5379 3482 5663 3486
rect 5667 3482 5702 3486
rect 3817 3481 5702 3482
rect 3817 3477 3818 3481
rect 84 3457 85 3463
rect 91 3462 1947 3463
rect 91 3458 111 3462
rect 115 3458 727 3462
rect 731 3458 807 3462
rect 811 3458 863 3462
rect 867 3458 943 3462
rect 947 3458 999 3462
rect 1003 3458 1079 3462
rect 1083 3458 1135 3462
rect 1139 3458 1215 3462
rect 1219 3458 1271 3462
rect 1275 3458 1351 3462
rect 1355 3458 1407 3462
rect 1411 3458 1487 3462
rect 1491 3458 1543 3462
rect 1547 3458 1623 3462
rect 1627 3458 1679 3462
rect 1683 3458 1759 3462
rect 1763 3458 1815 3462
rect 1819 3458 1935 3462
rect 1939 3458 1947 3462
rect 91 3457 1947 3458
rect 1953 3457 1954 3463
rect 3822 3369 3823 3375
rect 3829 3374 5707 3375
rect 3829 3370 3839 3374
rect 3843 3370 3859 3374
rect 3863 3370 4139 3374
rect 4143 3370 4427 3374
rect 4431 3370 4691 3374
rect 4695 3370 4803 3374
rect 4807 3370 4939 3374
rect 4943 3370 5075 3374
rect 5079 3370 5179 3374
rect 5183 3370 5211 3374
rect 5215 3370 5347 3374
rect 5351 3370 5427 3374
rect 5431 3370 5663 3374
rect 5667 3370 5707 3374
rect 3829 3369 5707 3370
rect 5713 3369 5714 3375
rect 1958 3357 1959 3363
rect 1965 3362 3823 3363
rect 1965 3358 1975 3362
rect 1979 3358 2531 3362
rect 2535 3358 2571 3362
rect 2575 3358 2715 3362
rect 2719 3358 2795 3362
rect 2799 3358 2899 3362
rect 2903 3358 3019 3362
rect 3023 3358 3083 3362
rect 3087 3358 3235 3362
rect 3239 3358 3267 3362
rect 3271 3358 3451 3362
rect 3455 3358 3651 3362
rect 3655 3358 3799 3362
rect 3803 3358 3823 3362
rect 1965 3357 3823 3358
rect 3829 3357 3830 3363
rect 96 3341 97 3347
rect 103 3346 1959 3347
rect 103 3342 111 3346
rect 115 3342 699 3346
rect 703 3342 755 3346
rect 759 3342 835 3346
rect 839 3342 891 3346
rect 895 3342 971 3346
rect 975 3342 1035 3346
rect 1039 3342 1107 3346
rect 1111 3342 1187 3346
rect 1191 3342 1243 3346
rect 1247 3342 1339 3346
rect 1343 3342 1379 3346
rect 1383 3342 1491 3346
rect 1495 3342 1515 3346
rect 1519 3342 1651 3346
rect 1655 3342 1787 3346
rect 1791 3342 1935 3346
rect 1939 3342 1959 3346
rect 103 3341 1959 3342
rect 1965 3341 1966 3347
rect 4522 3324 4528 3325
rect 5058 3324 5064 3325
rect 4522 3320 4523 3324
rect 4527 3320 5059 3324
rect 5063 3320 5064 3324
rect 4522 3319 4528 3320
rect 5058 3319 5064 3320
rect 1946 3245 1947 3251
rect 1953 3250 3811 3251
rect 1953 3246 1975 3250
rect 1979 3246 2023 3250
rect 2027 3246 2255 3250
rect 2259 3246 2503 3250
rect 2507 3246 2559 3250
rect 2563 3246 2743 3250
rect 2747 3246 2927 3250
rect 2931 3246 2975 3250
rect 2979 3246 3111 3250
rect 3115 3246 3207 3250
rect 3211 3246 3295 3250
rect 3299 3246 3447 3250
rect 3451 3246 3799 3250
rect 3803 3246 3811 3250
rect 1953 3245 3811 3246
rect 3817 3245 3818 3251
rect 84 3229 85 3235
rect 91 3234 1947 3235
rect 91 3230 111 3234
rect 115 3230 391 3234
rect 395 3230 647 3234
rect 651 3230 783 3234
rect 787 3230 919 3234
rect 923 3230 927 3234
rect 931 3230 1063 3234
rect 1067 3230 1215 3234
rect 1219 3230 1223 3234
rect 1227 3230 1367 3234
rect 1371 3230 1519 3234
rect 1523 3230 1527 3234
rect 1531 3230 1679 3234
rect 1683 3230 1815 3234
rect 1819 3230 1935 3234
rect 1939 3230 1947 3234
rect 91 3229 1947 3230
rect 1953 3229 1954 3235
rect 3810 3233 3811 3239
rect 3817 3238 5695 3239
rect 3817 3234 3839 3238
rect 3843 3234 3887 3238
rect 3891 3234 3911 3238
rect 3915 3234 4167 3238
rect 4171 3234 4183 3238
rect 4187 3234 4439 3238
rect 4443 3234 4455 3238
rect 4459 3234 4687 3238
rect 4691 3234 4719 3238
rect 4723 3234 4935 3238
rect 4939 3234 4967 3238
rect 4971 3234 5191 3238
rect 5195 3234 5207 3238
rect 5211 3234 5455 3238
rect 5459 3234 5663 3238
rect 5667 3234 5695 3238
rect 3817 3233 5695 3234
rect 5701 3233 5702 3239
rect 1958 3133 1959 3139
rect 1965 3138 3823 3139
rect 1965 3134 1975 3138
rect 1979 3134 1995 3138
rect 1999 3134 2227 3138
rect 2231 3134 2475 3138
rect 2479 3134 2483 3138
rect 2487 3134 2715 3138
rect 2719 3134 2779 3138
rect 2783 3134 2947 3138
rect 2951 3134 3075 3138
rect 3079 3134 3179 3138
rect 3183 3134 3371 3138
rect 3375 3134 3419 3138
rect 3423 3134 3651 3138
rect 3655 3134 3799 3138
rect 3803 3134 3823 3138
rect 1965 3133 3823 3134
rect 3829 3133 3830 3139
rect 3822 3117 3823 3123
rect 3829 3122 5707 3123
rect 3829 3118 3839 3122
rect 3843 3118 3883 3122
rect 3887 3118 3931 3122
rect 3935 3118 4131 3122
rect 4135 3118 4155 3122
rect 4159 3118 4331 3122
rect 4335 3118 4411 3122
rect 4415 3118 4523 3122
rect 4527 3118 4659 3122
rect 4663 3118 4715 3122
rect 4719 3118 4907 3122
rect 4911 3118 4915 3122
rect 4919 3118 5163 3122
rect 5167 3118 5663 3122
rect 5667 3118 5707 3122
rect 3829 3117 5707 3118
rect 5713 3117 5714 3123
rect 96 3105 97 3111
rect 103 3110 1959 3111
rect 103 3106 111 3110
rect 115 3106 131 3110
rect 135 3106 307 3110
rect 311 3106 363 3110
rect 367 3106 507 3110
rect 511 3106 619 3110
rect 623 3106 707 3110
rect 711 3106 899 3110
rect 903 3106 1091 3110
rect 1095 3106 1195 3110
rect 1199 3106 1275 3110
rect 1279 3106 1451 3110
rect 1455 3106 1499 3110
rect 1503 3106 1627 3110
rect 1631 3106 1787 3110
rect 1791 3106 1935 3110
rect 1939 3106 1959 3110
rect 103 3105 1959 3106
rect 1965 3105 1966 3111
rect 4226 3100 4232 3101
rect 5038 3100 5044 3101
rect 4226 3096 4227 3100
rect 4231 3096 5039 3100
rect 5043 3096 5044 3100
rect 4226 3095 4232 3096
rect 5038 3095 5044 3096
rect 1946 3013 1947 3019
rect 1953 3018 3811 3019
rect 1953 3014 1975 3018
rect 1979 3014 2191 3018
rect 2195 3014 2351 3018
rect 2355 3014 2511 3018
rect 2515 3014 2519 3018
rect 2523 3014 2703 3018
rect 2707 3014 2807 3018
rect 2811 3014 2903 3018
rect 2907 3014 3103 3018
rect 3107 3014 3119 3018
rect 3123 3014 3335 3018
rect 3339 3014 3399 3018
rect 3403 3014 3559 3018
rect 3563 3014 3679 3018
rect 3683 3014 3799 3018
rect 3803 3014 3811 3018
rect 1953 3013 3811 3014
rect 3817 3013 3818 3019
rect 84 2989 85 2995
rect 91 2994 1947 2995
rect 91 2990 111 2994
rect 115 2990 159 2994
rect 163 2990 295 2994
rect 299 2990 335 2994
rect 339 2990 431 2994
rect 435 2990 535 2994
rect 539 2990 567 2994
rect 571 2990 703 2994
rect 707 2990 735 2994
rect 739 2990 927 2994
rect 931 2990 1119 2994
rect 1123 2990 1303 2994
rect 1307 2990 1479 2994
rect 1483 2990 1655 2994
rect 1659 2990 1815 2994
rect 1819 2990 1935 2994
rect 1939 2990 1947 2994
rect 91 2989 1947 2990
rect 1953 2989 1954 2995
rect 3810 2981 3811 2987
rect 3817 2986 5695 2987
rect 3817 2982 3839 2986
rect 3843 2982 3959 2986
rect 3963 2982 3999 2986
rect 4003 2982 4159 2986
rect 4163 2982 4335 2986
rect 4339 2982 4359 2986
rect 4363 2982 4519 2986
rect 4523 2982 4551 2986
rect 4555 2982 4719 2986
rect 4723 2982 4743 2986
rect 4747 2982 4927 2986
rect 4931 2982 4943 2986
rect 4947 2982 5135 2986
rect 5139 2982 5351 2986
rect 5355 2982 5543 2986
rect 5547 2982 5663 2986
rect 5667 2982 5695 2986
rect 3817 2981 5695 2982
rect 5701 2981 5702 2987
rect 1958 2897 1959 2903
rect 1965 2902 3823 2903
rect 1965 2898 1975 2902
rect 1979 2898 1995 2902
rect 1999 2898 2131 2902
rect 2135 2898 2163 2902
rect 2167 2898 2267 2902
rect 2271 2898 2323 2902
rect 2327 2898 2403 2902
rect 2407 2898 2491 2902
rect 2495 2898 2539 2902
rect 2543 2898 2675 2902
rect 2679 2898 2683 2902
rect 2687 2898 2835 2902
rect 2839 2898 2875 2902
rect 2879 2898 2995 2902
rect 2999 2898 3091 2902
rect 3095 2898 3155 2902
rect 3159 2898 3307 2902
rect 3311 2898 3315 2902
rect 3319 2898 3531 2902
rect 3535 2898 3799 2902
rect 3803 2898 3823 2902
rect 1965 2897 3823 2898
rect 3829 2897 3830 2903
rect 96 2873 97 2879
rect 103 2878 1959 2879
rect 103 2874 111 2878
rect 115 2874 131 2878
rect 135 2874 227 2878
rect 231 2874 267 2878
rect 271 2874 363 2878
rect 367 2874 403 2878
rect 407 2874 499 2878
rect 503 2874 539 2878
rect 543 2874 635 2878
rect 639 2874 675 2878
rect 679 2874 771 2878
rect 775 2874 1935 2878
rect 1939 2874 1959 2878
rect 103 2873 1959 2874
rect 1965 2873 1966 2879
rect 3822 2853 3823 2859
rect 3829 2858 5707 2859
rect 3829 2854 3839 2858
rect 3843 2854 3859 2858
rect 3863 2854 3971 2858
rect 3975 2854 4011 2858
rect 4015 2854 4131 2858
rect 4135 2854 4211 2858
rect 4215 2854 4307 2858
rect 4311 2854 4435 2858
rect 4439 2854 4491 2858
rect 4495 2854 4691 2858
rect 4695 2854 4899 2858
rect 4903 2854 4963 2858
rect 4967 2854 5107 2858
rect 5111 2854 5251 2858
rect 5255 2854 5323 2858
rect 5327 2854 5515 2858
rect 5519 2854 5663 2858
rect 5667 2854 5707 2858
rect 3829 2853 5707 2854
rect 5713 2853 5714 2859
rect 1946 2781 1947 2787
rect 1953 2786 3811 2787
rect 1953 2782 1975 2786
rect 1979 2782 2023 2786
rect 2027 2782 2159 2786
rect 2163 2782 2295 2786
rect 2299 2782 2303 2786
rect 2307 2782 2431 2786
rect 2435 2782 2463 2786
rect 2467 2782 2567 2786
rect 2571 2782 2623 2786
rect 2627 2782 2711 2786
rect 2715 2782 2783 2786
rect 2787 2782 2863 2786
rect 2867 2782 2943 2786
rect 2947 2782 3023 2786
rect 3027 2782 3103 2786
rect 3107 2782 3183 2786
rect 3187 2782 3343 2786
rect 3347 2782 3799 2786
rect 3803 2782 3811 2786
rect 1953 2781 3811 2782
rect 3817 2781 3818 2787
rect 84 2757 85 2763
rect 91 2762 1947 2763
rect 91 2758 111 2762
rect 115 2758 255 2762
rect 259 2758 375 2762
rect 379 2758 391 2762
rect 395 2758 527 2762
rect 531 2758 575 2762
rect 579 2758 663 2762
rect 667 2758 799 2762
rect 803 2758 1039 2762
rect 1043 2758 1295 2762
rect 1299 2758 1567 2762
rect 1571 2758 1815 2762
rect 1819 2758 1935 2762
rect 1939 2758 1947 2762
rect 91 2757 1947 2758
rect 1953 2757 1954 2763
rect 3810 2729 3811 2735
rect 3817 2734 5695 2735
rect 3817 2730 3839 2734
rect 3843 2730 3887 2734
rect 3891 2730 3967 2734
rect 3971 2730 4039 2734
rect 4043 2730 4223 2734
rect 4227 2730 4239 2734
rect 4243 2730 4463 2734
rect 4467 2730 4527 2734
rect 4531 2730 4719 2734
rect 4723 2730 4863 2734
rect 4867 2730 4991 2734
rect 4995 2730 5215 2734
rect 5219 2730 5279 2734
rect 5283 2730 5543 2734
rect 5547 2730 5663 2734
rect 5667 2730 5695 2734
rect 3817 2729 5695 2730
rect 5701 2729 5702 2735
rect 1958 2661 1959 2667
rect 1965 2666 3823 2667
rect 1965 2662 1975 2666
rect 1979 2662 1995 2666
rect 1999 2662 2131 2666
rect 2135 2662 2275 2666
rect 2279 2662 2435 2666
rect 2439 2662 2595 2666
rect 2599 2662 2699 2666
rect 2703 2662 2755 2666
rect 2759 2662 2835 2666
rect 2839 2662 2915 2666
rect 2919 2662 2971 2666
rect 2975 2662 3075 2666
rect 3079 2662 3799 2666
rect 3803 2662 3823 2666
rect 1965 2661 3823 2662
rect 3829 2661 3830 2667
rect 96 2645 97 2651
rect 103 2650 1959 2651
rect 103 2646 111 2650
rect 115 2646 347 2650
rect 351 2646 387 2650
rect 391 2646 539 2650
rect 543 2646 547 2650
rect 551 2646 699 2650
rect 703 2646 771 2650
rect 775 2646 867 2650
rect 871 2646 1011 2650
rect 1015 2646 1035 2650
rect 1039 2646 1203 2650
rect 1207 2646 1267 2650
rect 1271 2646 1371 2650
rect 1375 2646 1539 2650
rect 1543 2646 1715 2650
rect 1719 2646 1787 2650
rect 1791 2646 1935 2650
rect 1939 2646 1959 2650
rect 103 2645 1959 2646
rect 1965 2645 1966 2651
rect 3822 2617 3823 2623
rect 3829 2622 5707 2623
rect 3829 2618 3839 2622
rect 3843 2618 3891 2622
rect 3895 2618 3939 2622
rect 3943 2618 4067 2622
rect 4071 2618 4195 2622
rect 4199 2618 4267 2622
rect 4271 2618 4491 2622
rect 4495 2618 4499 2622
rect 4503 2618 4731 2622
rect 4735 2618 4835 2622
rect 4839 2618 4995 2622
rect 4999 2618 5187 2622
rect 5191 2618 5267 2622
rect 5271 2618 5515 2622
rect 5519 2618 5663 2622
rect 5667 2618 5707 2622
rect 3829 2617 5707 2618
rect 5713 2617 5714 2623
rect 1946 2549 1947 2555
rect 1953 2554 3811 2555
rect 1953 2550 1975 2554
rect 1979 2550 2607 2554
rect 2611 2550 2727 2554
rect 2731 2550 2759 2554
rect 2763 2550 2863 2554
rect 2867 2550 2911 2554
rect 2915 2550 2999 2554
rect 3003 2550 3063 2554
rect 3067 2550 3223 2554
rect 3227 2550 3799 2554
rect 3803 2550 3811 2554
rect 1953 2549 3811 2550
rect 3817 2549 3818 2555
rect 84 2533 85 2539
rect 91 2538 1947 2539
rect 91 2534 111 2538
rect 115 2534 327 2538
rect 331 2534 415 2538
rect 419 2534 535 2538
rect 539 2534 567 2538
rect 571 2534 727 2538
rect 731 2534 735 2538
rect 739 2534 895 2538
rect 899 2534 919 2538
rect 923 2534 1063 2538
rect 1067 2534 1095 2538
rect 1099 2534 1231 2538
rect 1235 2534 1271 2538
rect 1275 2534 1399 2538
rect 1403 2534 1439 2538
rect 1443 2534 1567 2538
rect 1571 2534 1607 2538
rect 1611 2534 1743 2538
rect 1747 2534 1775 2538
rect 1779 2534 1935 2538
rect 1939 2534 1947 2538
rect 91 2533 1947 2534
rect 1953 2533 1954 2539
rect 3810 2501 3811 2507
rect 3817 2506 5695 2507
rect 3817 2502 3839 2506
rect 3843 2502 3887 2506
rect 3891 2502 3919 2506
rect 3923 2502 4087 2506
rect 4091 2502 4095 2506
rect 4099 2502 4295 2506
rect 4299 2502 4319 2506
rect 4323 2502 4519 2506
rect 4523 2502 4567 2506
rect 4571 2502 4759 2506
rect 4763 2502 4823 2506
rect 4827 2502 5023 2506
rect 5027 2502 5087 2506
rect 5091 2502 5295 2506
rect 5299 2502 5351 2506
rect 5355 2502 5543 2506
rect 5547 2502 5663 2506
rect 5667 2502 5695 2506
rect 3817 2501 5695 2502
rect 5701 2501 5702 2507
rect 4386 2468 4392 2469
rect 5114 2468 5120 2469
rect 4386 2464 4387 2468
rect 4391 2464 5115 2468
rect 5119 2464 5120 2468
rect 4386 2463 4392 2464
rect 5114 2463 5120 2464
rect 1958 2426 3830 2427
rect 1958 2423 1975 2426
rect 96 2417 97 2423
rect 103 2422 1959 2423
rect 103 2418 111 2422
rect 115 2418 131 2422
rect 135 2418 299 2422
rect 303 2418 403 2422
rect 407 2418 507 2422
rect 511 2418 691 2422
rect 695 2418 707 2422
rect 711 2418 891 2422
rect 895 2418 971 2422
rect 975 2418 1067 2422
rect 1071 2418 1243 2422
rect 1247 2418 1251 2422
rect 1255 2418 1411 2422
rect 1415 2418 1531 2422
rect 1535 2418 1579 2422
rect 1583 2418 1747 2422
rect 1751 2418 1787 2422
rect 1791 2418 1935 2422
rect 1939 2418 1959 2422
rect 103 2417 1959 2418
rect 1965 2422 1975 2423
rect 1979 2422 1995 2426
rect 1999 2422 2275 2426
rect 2279 2422 2571 2426
rect 2575 2422 2579 2426
rect 2583 2422 2731 2426
rect 2735 2422 2859 2426
rect 2863 2422 2883 2426
rect 2887 2422 3035 2426
rect 3039 2422 3147 2426
rect 3151 2422 3195 2426
rect 3199 2422 3435 2426
rect 3439 2422 3799 2426
rect 3803 2422 3830 2426
rect 1965 2421 3830 2422
rect 1965 2417 1966 2421
rect 3822 2389 3823 2395
rect 3829 2394 5707 2395
rect 3829 2390 3839 2394
rect 3843 2390 3859 2394
rect 3863 2390 4059 2394
rect 4063 2390 4091 2394
rect 4095 2390 4291 2394
rect 4295 2390 4339 2394
rect 4343 2390 4539 2394
rect 4543 2390 4579 2394
rect 4583 2390 4795 2394
rect 4799 2390 4811 2394
rect 4815 2390 5043 2394
rect 5047 2390 5059 2394
rect 5063 2390 5283 2394
rect 5287 2390 5323 2394
rect 5327 2390 5515 2394
rect 5519 2390 5663 2394
rect 5667 2390 5707 2394
rect 3829 2389 5707 2390
rect 5713 2389 5714 2395
rect 1946 2297 1947 2303
rect 1953 2302 3811 2303
rect 1953 2298 1975 2302
rect 1979 2298 2023 2302
rect 2027 2298 2159 2302
rect 2163 2298 2295 2302
rect 2299 2298 2303 2302
rect 2307 2298 2447 2302
rect 2451 2298 2599 2302
rect 2603 2298 2607 2302
rect 2611 2298 2767 2302
rect 2771 2298 2887 2302
rect 2891 2298 2927 2302
rect 2931 2298 3079 2302
rect 3083 2298 3175 2302
rect 3179 2298 3231 2302
rect 3235 2298 3383 2302
rect 3387 2298 3463 2302
rect 3467 2298 3543 2302
rect 3547 2298 3679 2302
rect 3683 2298 3799 2302
rect 3803 2298 3811 2302
rect 1953 2297 3811 2298
rect 3817 2297 3818 2303
rect 1946 2295 1954 2297
rect 84 2289 85 2295
rect 91 2294 1947 2295
rect 91 2290 111 2294
rect 115 2290 159 2294
rect 163 2290 423 2294
rect 427 2290 431 2294
rect 435 2290 711 2294
rect 715 2290 719 2294
rect 723 2290 999 2294
rect 1003 2290 1279 2294
rect 1283 2290 1295 2294
rect 1299 2290 1559 2294
rect 1563 2290 1815 2294
rect 1819 2290 1935 2294
rect 1939 2290 1947 2294
rect 91 2289 1947 2290
rect 1953 2289 1954 2295
rect 3810 2253 3811 2259
rect 3817 2258 5695 2259
rect 3817 2254 3839 2258
rect 3843 2254 3887 2258
rect 3891 2254 4119 2258
rect 4123 2254 4367 2258
rect 4371 2254 4591 2258
rect 4595 2254 4607 2258
rect 4611 2254 4727 2258
rect 4731 2254 4839 2258
rect 4843 2254 4863 2258
rect 4867 2254 4999 2258
rect 5003 2254 5071 2258
rect 5075 2254 5135 2258
rect 5139 2254 5271 2258
rect 5275 2254 5311 2258
rect 5315 2254 5407 2258
rect 5411 2254 5543 2258
rect 5547 2254 5663 2258
rect 5667 2254 5695 2258
rect 3817 2253 5695 2254
rect 5701 2253 5702 2259
rect 1958 2177 1959 2183
rect 1965 2182 3823 2183
rect 1965 2178 1975 2182
rect 1979 2178 1995 2182
rect 1999 2178 2131 2182
rect 2135 2178 2267 2182
rect 2271 2178 2331 2182
rect 2335 2178 2419 2182
rect 2423 2178 2531 2182
rect 2535 2178 2579 2182
rect 2583 2178 2731 2182
rect 2735 2178 2739 2182
rect 2743 2178 2899 2182
rect 2903 2178 2923 2182
rect 2927 2178 3051 2182
rect 3055 2178 3115 2182
rect 3119 2178 3203 2182
rect 3207 2178 3299 2182
rect 3303 2178 3355 2182
rect 3359 2178 3483 2182
rect 3487 2178 3515 2182
rect 3519 2178 3651 2182
rect 3655 2178 3799 2182
rect 3803 2178 3823 2182
rect 1965 2177 3823 2178
rect 3829 2177 3830 2183
rect 96 2165 97 2171
rect 103 2170 1959 2171
rect 103 2166 111 2170
rect 115 2166 131 2170
rect 135 2166 395 2170
rect 399 2166 403 2170
rect 407 2166 683 2170
rect 687 2166 731 2170
rect 735 2166 971 2170
rect 975 2166 1083 2170
rect 1087 2166 1267 2170
rect 1271 2166 1443 2170
rect 1447 2166 1787 2170
rect 1791 2166 1935 2170
rect 1939 2166 1959 2170
rect 103 2165 1959 2166
rect 1965 2165 1966 2171
rect 3822 2125 3823 2131
rect 3829 2130 5707 2131
rect 3829 2126 3839 2130
rect 3843 2126 4563 2130
rect 4567 2126 4699 2130
rect 4703 2126 4835 2130
rect 4839 2126 4955 2130
rect 4959 2126 4971 2130
rect 4975 2126 5091 2130
rect 5095 2126 5107 2130
rect 5111 2126 5227 2130
rect 5231 2126 5243 2130
rect 5247 2126 5379 2130
rect 5383 2126 5515 2130
rect 5519 2126 5663 2130
rect 5667 2126 5707 2130
rect 3829 2125 5707 2126
rect 5713 2125 5714 2131
rect 1946 2057 1947 2063
rect 1953 2062 3811 2063
rect 1953 2058 1975 2062
rect 1979 2058 2023 2062
rect 2027 2058 2159 2062
rect 2163 2058 2279 2062
rect 2283 2058 2359 2062
rect 2363 2058 2551 2062
rect 2555 2058 2559 2062
rect 2563 2058 2759 2062
rect 2763 2058 2799 2062
rect 2803 2058 2951 2062
rect 2955 2058 3031 2062
rect 3035 2058 3143 2062
rect 3147 2058 3255 2062
rect 3259 2058 3327 2062
rect 3331 2058 3479 2062
rect 3483 2058 3511 2062
rect 3515 2058 3679 2062
rect 3683 2058 3799 2062
rect 3803 2058 3811 2062
rect 1953 2057 3811 2058
rect 3817 2057 3818 2063
rect 1946 2055 1954 2057
rect 84 2049 85 2055
rect 91 2054 1947 2055
rect 91 2050 111 2054
rect 115 2050 159 2054
rect 163 2050 223 2054
rect 227 2050 383 2054
rect 387 2050 431 2054
rect 435 2050 559 2054
rect 563 2050 751 2054
rect 755 2050 759 2054
rect 763 2050 959 2054
rect 963 2050 1111 2054
rect 1115 2050 1167 2054
rect 1171 2050 1383 2054
rect 1387 2050 1471 2054
rect 1475 2050 1607 2054
rect 1611 2050 1815 2054
rect 1819 2050 1935 2054
rect 1939 2050 1947 2054
rect 91 2049 1947 2050
rect 1953 2049 1954 2055
rect 3810 2013 3811 2019
rect 3817 2018 5695 2019
rect 3817 2014 3839 2018
rect 3843 2014 4727 2018
rect 4731 2014 4863 2018
rect 4867 2014 4983 2018
rect 4987 2014 5007 2018
rect 5011 2014 5119 2018
rect 5123 2014 5159 2018
rect 5163 2014 5255 2018
rect 5259 2014 5319 2018
rect 5323 2014 5487 2018
rect 5491 2014 5663 2018
rect 5667 2014 5695 2018
rect 3817 2013 5695 2014
rect 5701 2013 5702 2019
rect 1958 1938 3830 1939
rect 1958 1935 1975 1938
rect 96 1929 97 1935
rect 103 1934 1959 1935
rect 103 1930 111 1934
rect 115 1930 195 1934
rect 199 1930 355 1934
rect 359 1930 387 1934
rect 391 1930 531 1934
rect 535 1930 595 1934
rect 599 1930 723 1934
rect 727 1930 819 1934
rect 823 1930 931 1934
rect 935 1930 1051 1934
rect 1055 1930 1139 1934
rect 1143 1930 1283 1934
rect 1287 1930 1355 1934
rect 1359 1930 1523 1934
rect 1527 1930 1579 1934
rect 1583 1930 1771 1934
rect 1775 1930 1787 1934
rect 1791 1930 1935 1934
rect 1939 1930 1959 1934
rect 103 1929 1959 1930
rect 1965 1934 1975 1935
rect 1979 1934 1995 1938
rect 1999 1934 2251 1938
rect 2255 1934 2315 1938
rect 2319 1934 2523 1938
rect 2527 1934 2619 1938
rect 2623 1934 2771 1938
rect 2775 1934 2899 1938
rect 2903 1934 3003 1938
rect 3007 1934 3163 1938
rect 3167 1934 3227 1938
rect 3231 1934 3419 1938
rect 3423 1934 3451 1938
rect 3455 1934 3651 1938
rect 3655 1934 3799 1938
rect 3803 1934 3830 1938
rect 1965 1933 3830 1934
rect 1965 1929 1966 1933
rect 3822 1901 3823 1907
rect 3829 1906 5707 1907
rect 3829 1902 3839 1906
rect 3843 1902 4275 1906
rect 4279 1902 4499 1906
rect 4503 1902 4699 1906
rect 4703 1902 4731 1906
rect 4735 1902 4835 1906
rect 4839 1902 4979 1906
rect 4983 1902 5131 1906
rect 5135 1902 5235 1906
rect 5239 1902 5291 1906
rect 5295 1902 5459 1906
rect 5463 1902 5499 1906
rect 5503 1902 5663 1906
rect 5667 1902 5707 1906
rect 3829 1901 5707 1902
rect 5713 1901 5714 1907
rect 1946 1817 1947 1823
rect 1953 1822 3811 1823
rect 1953 1818 1975 1822
rect 1979 1818 2023 1822
rect 2027 1818 2111 1822
rect 2115 1818 2343 1822
rect 2347 1818 2391 1822
rect 2395 1818 2647 1822
rect 2651 1818 2663 1822
rect 2667 1818 2927 1822
rect 2931 1818 3183 1822
rect 3187 1818 3191 1822
rect 3195 1818 3439 1822
rect 3443 1818 3447 1822
rect 3451 1818 3679 1822
rect 3683 1818 3799 1822
rect 3803 1818 3811 1822
rect 1953 1817 3811 1818
rect 3817 1817 3818 1823
rect 84 1801 85 1807
rect 91 1806 1947 1807
rect 91 1802 111 1806
rect 115 1802 159 1806
rect 163 1802 223 1806
rect 227 1802 303 1806
rect 307 1802 415 1806
rect 419 1802 479 1806
rect 483 1802 623 1806
rect 627 1802 655 1806
rect 659 1802 831 1806
rect 835 1802 847 1806
rect 851 1802 1007 1806
rect 1011 1802 1079 1806
rect 1083 1802 1183 1806
rect 1187 1802 1311 1806
rect 1315 1802 1359 1806
rect 1363 1802 1535 1806
rect 1539 1802 1551 1806
rect 1555 1802 1711 1806
rect 1715 1802 1799 1806
rect 1803 1802 1935 1806
rect 1939 1802 1947 1806
rect 91 1801 1947 1802
rect 1953 1801 1954 1807
rect 3810 1781 3811 1787
rect 3817 1786 5695 1787
rect 3817 1782 3839 1786
rect 3843 1782 3887 1786
rect 3891 1782 4087 1786
rect 4091 1782 4303 1786
rect 4307 1782 4343 1786
rect 4347 1782 4527 1786
rect 4531 1782 4623 1786
rect 4627 1782 4759 1786
rect 4763 1782 4927 1786
rect 4931 1782 5007 1786
rect 5011 1782 5247 1786
rect 5251 1782 5263 1786
rect 5267 1782 5527 1786
rect 5531 1782 5543 1786
rect 5547 1782 5663 1786
rect 5667 1782 5695 1786
rect 3817 1781 5695 1782
rect 5701 1781 5702 1787
rect 96 1685 97 1691
rect 103 1690 1959 1691
rect 103 1686 111 1690
rect 115 1686 131 1690
rect 135 1686 275 1690
rect 279 1686 451 1690
rect 455 1686 627 1690
rect 631 1686 803 1690
rect 807 1686 875 1690
rect 879 1686 979 1690
rect 983 1686 1011 1690
rect 1015 1686 1147 1690
rect 1151 1686 1155 1690
rect 1159 1686 1283 1690
rect 1287 1686 1331 1690
rect 1335 1686 1419 1690
rect 1423 1686 1507 1690
rect 1511 1686 1555 1690
rect 1559 1686 1683 1690
rect 1687 1686 1935 1690
rect 1939 1686 1959 1690
rect 103 1685 1959 1686
rect 1965 1685 1966 1691
rect 1958 1673 1959 1679
rect 1965 1678 3823 1679
rect 1965 1674 1975 1678
rect 1979 1674 2083 1678
rect 2087 1674 2219 1678
rect 2223 1674 2355 1678
rect 2359 1674 2363 1678
rect 2367 1674 2491 1678
rect 2495 1674 2627 1678
rect 2631 1674 2635 1678
rect 2639 1674 2771 1678
rect 2775 1674 2899 1678
rect 2903 1674 2915 1678
rect 2919 1674 3155 1678
rect 3159 1674 3411 1678
rect 3415 1674 3651 1678
rect 3655 1674 3799 1678
rect 3803 1674 3823 1678
rect 1965 1673 3823 1674
rect 3829 1673 3830 1679
rect 3822 1671 3830 1673
rect 3822 1665 3823 1671
rect 3829 1670 5707 1671
rect 3829 1666 3839 1670
rect 3843 1666 3859 1670
rect 3863 1666 3995 1670
rect 3999 1666 4059 1670
rect 4063 1666 4139 1670
rect 4143 1666 4315 1670
rect 4319 1666 4323 1670
rect 4327 1666 4531 1670
rect 4535 1666 4595 1670
rect 4599 1666 4763 1670
rect 4767 1666 4899 1670
rect 4903 1666 5011 1670
rect 5015 1666 5219 1670
rect 5223 1666 5275 1670
rect 5279 1666 5515 1670
rect 5519 1666 5663 1670
rect 5667 1666 5707 1670
rect 3829 1665 5707 1666
rect 5713 1665 5714 1671
rect 1946 1562 3818 1563
rect 1946 1559 1975 1562
rect 84 1553 85 1559
rect 91 1558 1947 1559
rect 91 1554 111 1558
rect 115 1554 159 1558
rect 163 1554 391 1558
rect 395 1554 631 1558
rect 635 1554 871 1558
rect 875 1554 903 1558
rect 907 1554 1039 1558
rect 1043 1554 1111 1558
rect 1115 1554 1175 1558
rect 1179 1554 1311 1558
rect 1315 1554 1351 1558
rect 1355 1554 1447 1558
rect 1451 1554 1583 1558
rect 1587 1554 1935 1558
rect 1939 1554 1947 1558
rect 91 1553 1947 1554
rect 1953 1558 1975 1559
rect 1979 1558 2111 1562
rect 2115 1558 2143 1562
rect 2147 1558 2247 1562
rect 2251 1558 2279 1562
rect 2283 1558 2383 1562
rect 2387 1558 2415 1562
rect 2419 1558 2519 1562
rect 2523 1558 2551 1562
rect 2555 1558 2655 1562
rect 2659 1558 2687 1562
rect 2691 1558 2799 1562
rect 2803 1558 2823 1562
rect 2827 1558 2943 1562
rect 2947 1558 2959 1562
rect 2963 1558 3095 1562
rect 3099 1558 3231 1562
rect 3235 1558 3799 1562
rect 3803 1558 3818 1562
rect 1953 1557 3818 1558
rect 1953 1553 1954 1557
rect 3810 1555 3818 1557
rect 3810 1549 3811 1555
rect 3817 1554 5695 1555
rect 3817 1550 3839 1554
rect 3843 1550 3887 1554
rect 3891 1550 4023 1554
rect 4027 1550 4111 1554
rect 4115 1550 4167 1554
rect 4171 1550 4343 1554
rect 4347 1550 4351 1554
rect 4355 1550 4559 1554
rect 4563 1550 4575 1554
rect 4579 1550 4791 1554
rect 4795 1550 4815 1554
rect 4819 1550 5039 1554
rect 5043 1550 5063 1554
rect 5067 1550 5303 1554
rect 5307 1550 5311 1554
rect 5315 1550 5543 1554
rect 5547 1550 5663 1554
rect 5667 1550 5695 1554
rect 3817 1549 5695 1550
rect 5701 1549 5702 1555
rect 3822 1437 3823 1443
rect 3829 1442 5707 1443
rect 3829 1438 3839 1442
rect 3843 1438 3859 1442
rect 3863 1438 4083 1442
rect 4087 1438 4315 1442
rect 4319 1438 4323 1442
rect 4327 1438 4547 1442
rect 4551 1438 4771 1442
rect 4775 1438 4787 1442
rect 4791 1438 4987 1442
rect 4991 1438 5035 1442
rect 5039 1438 5203 1442
rect 5207 1438 5283 1442
rect 5287 1438 5419 1442
rect 5423 1438 5515 1442
rect 5519 1438 5663 1442
rect 5667 1438 5707 1442
rect 3829 1437 5707 1438
rect 5713 1437 5714 1443
rect 3822 1435 3830 1437
rect 96 1429 97 1435
rect 103 1434 1959 1435
rect 103 1430 111 1434
rect 115 1430 131 1434
rect 135 1430 331 1434
rect 335 1430 363 1434
rect 367 1430 555 1434
rect 559 1430 603 1434
rect 607 1430 779 1434
rect 783 1430 843 1434
rect 847 1430 1003 1434
rect 1007 1430 1083 1434
rect 1087 1430 1323 1434
rect 1327 1430 1935 1434
rect 1939 1430 1959 1434
rect 103 1429 1959 1430
rect 1965 1434 3830 1435
rect 1965 1430 1975 1434
rect 1979 1430 2099 1434
rect 2103 1430 2115 1434
rect 2119 1430 2243 1434
rect 2247 1430 2251 1434
rect 2255 1430 2387 1434
rect 2391 1430 2523 1434
rect 2527 1430 2539 1434
rect 2543 1430 2659 1434
rect 2663 1430 2691 1434
rect 2695 1430 2795 1434
rect 2799 1430 2851 1434
rect 2855 1430 2931 1434
rect 2935 1430 3011 1434
rect 3015 1430 3067 1434
rect 3071 1430 3171 1434
rect 3175 1430 3203 1434
rect 3207 1430 3799 1434
rect 3803 1430 3830 1434
rect 1965 1429 3830 1430
rect 3810 1325 3811 1331
rect 3817 1330 5695 1331
rect 3817 1326 3839 1330
rect 3843 1326 3887 1330
rect 3891 1326 4111 1330
rect 4115 1326 4119 1330
rect 4123 1326 4351 1330
rect 4355 1326 4391 1330
rect 4395 1326 4575 1330
rect 4579 1326 4671 1330
rect 4675 1326 4799 1330
rect 4803 1326 4967 1330
rect 4971 1326 5015 1330
rect 5019 1326 5231 1330
rect 5235 1326 5263 1330
rect 5267 1326 5447 1330
rect 5451 1326 5543 1330
rect 5547 1326 5663 1330
rect 5667 1326 5695 1330
rect 3817 1325 5695 1326
rect 5701 1325 5702 1331
rect 84 1317 85 1323
rect 91 1322 1947 1323
rect 91 1318 111 1322
rect 115 1318 159 1322
rect 163 1318 359 1322
rect 363 1318 367 1322
rect 371 1318 583 1322
rect 587 1318 607 1322
rect 611 1318 807 1322
rect 811 1318 847 1322
rect 851 1318 1031 1322
rect 1035 1318 1087 1322
rect 1091 1318 1935 1322
rect 1939 1318 1947 1322
rect 91 1317 1947 1318
rect 1953 1319 1954 1323
rect 1953 1318 3818 1319
rect 1953 1317 1975 1318
rect 1946 1314 1975 1317
rect 1979 1314 2023 1318
rect 2027 1314 2127 1318
rect 2131 1314 2175 1318
rect 2179 1314 2271 1318
rect 2275 1314 2367 1318
rect 2371 1314 2415 1318
rect 2419 1314 2567 1318
rect 2571 1314 2575 1318
rect 2579 1314 2719 1318
rect 2723 1314 2791 1318
rect 2795 1314 2879 1318
rect 2883 1314 3015 1318
rect 3019 1314 3039 1318
rect 3043 1314 3199 1318
rect 3203 1314 3239 1318
rect 3243 1314 3471 1318
rect 3475 1314 3679 1318
rect 3683 1314 3799 1318
rect 3803 1314 3818 1318
rect 1946 1313 3818 1314
rect 96 1193 97 1199
rect 103 1198 1959 1199
rect 103 1194 111 1198
rect 115 1194 131 1198
rect 135 1194 275 1198
rect 279 1194 339 1198
rect 343 1194 443 1198
rect 447 1194 579 1198
rect 583 1194 603 1198
rect 607 1194 763 1198
rect 767 1194 819 1198
rect 823 1194 923 1198
rect 927 1194 1059 1198
rect 1063 1194 1075 1198
rect 1079 1194 1219 1198
rect 1223 1194 1363 1198
rect 1367 1194 1507 1198
rect 1511 1194 1651 1198
rect 1655 1194 1787 1198
rect 1791 1194 1935 1198
rect 1939 1194 1959 1198
rect 103 1193 1959 1194
rect 1965 1198 5714 1199
rect 1965 1194 1975 1198
rect 1979 1194 1995 1198
rect 1999 1194 2147 1198
rect 2151 1194 2339 1198
rect 2343 1194 2547 1198
rect 2551 1194 2723 1198
rect 2727 1194 2763 1198
rect 2767 1194 2899 1198
rect 2903 1194 2987 1198
rect 2991 1194 3083 1198
rect 3087 1194 3211 1198
rect 3215 1194 3275 1198
rect 3279 1194 3443 1198
rect 3447 1194 3467 1198
rect 3471 1194 3651 1198
rect 3655 1194 3799 1198
rect 3803 1194 3839 1198
rect 3843 1194 3859 1198
rect 3863 1194 4011 1198
rect 4015 1194 4091 1198
rect 4095 1194 4211 1198
rect 4215 1194 4363 1198
rect 4367 1194 4435 1198
rect 4439 1194 4643 1198
rect 4647 1194 4691 1198
rect 4695 1194 4939 1198
rect 4943 1194 4963 1198
rect 4967 1194 5235 1198
rect 5239 1194 5251 1198
rect 5255 1194 5515 1198
rect 5519 1194 5663 1198
rect 5667 1194 5714 1198
rect 1965 1193 5714 1194
rect 84 1073 85 1079
rect 91 1078 1947 1079
rect 91 1074 111 1078
rect 115 1074 159 1078
rect 163 1074 175 1078
rect 179 1074 303 1078
rect 307 1074 415 1078
rect 419 1074 471 1078
rect 475 1074 631 1078
rect 635 1074 639 1078
rect 643 1074 791 1078
rect 795 1074 855 1078
rect 859 1074 951 1078
rect 955 1074 1055 1078
rect 1059 1074 1103 1078
rect 1107 1074 1239 1078
rect 1243 1074 1247 1078
rect 1251 1074 1391 1078
rect 1395 1074 1423 1078
rect 1427 1074 1535 1078
rect 1539 1074 1607 1078
rect 1611 1074 1679 1078
rect 1683 1074 1791 1078
rect 1795 1074 1815 1078
rect 1819 1074 1935 1078
rect 1939 1074 1947 1078
rect 91 1073 1947 1074
rect 1953 1075 1954 1079
rect 1953 1074 5702 1075
rect 1953 1073 1975 1074
rect 1946 1070 1975 1073
rect 1979 1070 2559 1074
rect 2563 1070 2751 1074
rect 2755 1070 2927 1074
rect 2931 1070 2951 1074
rect 2955 1070 3111 1074
rect 3115 1070 3151 1074
rect 3155 1070 3303 1074
rect 3307 1070 3359 1074
rect 3363 1070 3495 1074
rect 3499 1070 3575 1074
rect 3579 1070 3679 1074
rect 3683 1070 3799 1074
rect 3803 1070 3839 1074
rect 3843 1070 4039 1074
rect 4043 1070 4095 1074
rect 4099 1070 4239 1074
rect 4243 1070 4391 1074
rect 4395 1070 4463 1074
rect 4467 1070 4687 1074
rect 4691 1070 4719 1074
rect 4723 1070 4975 1074
rect 4979 1070 4991 1074
rect 4995 1070 5263 1074
rect 5267 1070 5279 1074
rect 5283 1070 5543 1074
rect 5547 1070 5663 1074
rect 5667 1070 5702 1074
rect 1946 1069 5702 1070
rect 1958 962 3830 963
rect 1958 959 1975 962
rect 96 953 97 959
rect 103 958 1959 959
rect 103 954 111 958
rect 115 954 147 958
rect 151 954 195 958
rect 199 954 387 958
rect 391 954 419 958
rect 423 954 611 958
rect 615 954 667 958
rect 671 954 827 958
rect 831 954 931 958
rect 935 954 1027 958
rect 1031 954 1211 958
rect 1215 954 1219 958
rect 1223 954 1395 958
rect 1399 954 1515 958
rect 1519 954 1579 958
rect 1583 954 1763 958
rect 1767 954 1787 958
rect 1791 954 1935 958
rect 1939 954 1959 958
rect 103 953 1959 954
rect 1965 958 1975 959
rect 1979 958 1995 962
rect 1999 958 2219 962
rect 2223 958 2467 962
rect 2471 958 2531 962
rect 2535 958 2707 962
rect 2711 958 2723 962
rect 2727 958 2923 962
rect 2927 958 2939 962
rect 2943 958 3123 962
rect 3127 958 3171 962
rect 3175 958 3331 962
rect 3335 958 3411 962
rect 3415 958 3547 962
rect 3551 958 3799 962
rect 3803 959 3830 962
rect 3803 958 5714 959
rect 1965 957 3839 958
rect 1965 953 1966 957
rect 3822 954 3839 957
rect 3843 954 3931 958
rect 3935 954 4067 958
rect 4071 954 4155 958
rect 4159 954 4363 958
rect 4367 954 4379 958
rect 4383 954 4595 958
rect 4599 954 4659 958
rect 4663 954 4811 958
rect 4815 954 4947 958
rect 4951 954 5027 958
rect 5031 954 5235 958
rect 5239 954 5243 958
rect 5247 954 5467 958
rect 5471 954 5515 958
rect 5519 954 5663 958
rect 5667 954 5714 958
rect 3822 953 5714 954
rect 1946 845 1947 851
rect 1953 850 3811 851
rect 1953 846 1975 850
rect 1979 846 2023 850
rect 2027 846 2223 850
rect 2227 846 2247 850
rect 2251 846 2439 850
rect 2443 846 2495 850
rect 2499 846 2663 850
rect 2667 846 2735 850
rect 2739 846 2887 850
rect 2891 846 2967 850
rect 2971 846 3111 850
rect 3115 846 3199 850
rect 3203 846 3335 850
rect 3339 846 3439 850
rect 3443 846 3559 850
rect 3563 846 3799 850
rect 3803 846 3811 850
rect 1953 845 3811 846
rect 3817 847 3818 851
rect 3817 846 5702 847
rect 3817 845 3839 846
rect 3810 842 3839 845
rect 3843 842 3887 846
rect 3891 842 3959 846
rect 3963 842 4111 846
rect 4115 842 4183 846
rect 4187 842 4343 846
rect 4347 842 4407 846
rect 4411 842 4575 846
rect 4579 842 4623 846
rect 4627 842 4799 846
rect 4803 842 4839 846
rect 4843 842 5031 846
rect 5035 842 5055 846
rect 5059 842 5263 846
rect 5267 842 5271 846
rect 5275 842 5495 846
rect 5499 842 5663 846
rect 5667 842 5702 846
rect 3810 841 5702 842
rect 84 817 85 823
rect 91 822 1947 823
rect 91 818 111 822
rect 115 818 223 822
rect 227 818 447 822
rect 451 818 663 822
rect 667 818 695 822
rect 699 818 879 822
rect 883 818 959 822
rect 963 818 1087 822
rect 1091 818 1247 822
rect 1251 818 1295 822
rect 1299 818 1511 822
rect 1515 818 1543 822
rect 1547 818 1815 822
rect 1819 818 1935 822
rect 1939 818 1947 822
rect 91 817 1947 818
rect 1953 817 1954 823
rect 3822 729 3823 735
rect 3829 734 5707 735
rect 3829 730 3839 734
rect 3843 730 3859 734
rect 3863 730 4083 734
rect 4087 730 4315 734
rect 4319 730 4323 734
rect 4327 730 4547 734
rect 4551 730 4555 734
rect 4559 730 4771 734
rect 4775 730 4779 734
rect 4783 730 5003 734
rect 5007 730 5227 734
rect 5231 730 5235 734
rect 5239 730 5459 734
rect 5463 730 5467 734
rect 5471 730 5663 734
rect 5667 730 5707 734
rect 3829 729 5707 730
rect 5713 729 5714 735
rect 1958 717 1959 723
rect 1965 722 3823 723
rect 1965 718 1975 722
rect 1979 718 2195 722
rect 2199 718 2411 722
rect 2415 718 2635 722
rect 2639 718 2859 722
rect 2863 718 3083 722
rect 3087 718 3307 722
rect 3311 718 3379 722
rect 3383 718 3515 722
rect 3519 718 3531 722
rect 3535 718 3651 722
rect 3655 718 3799 722
rect 3803 718 3823 722
rect 1965 717 3823 718
rect 3829 717 3830 723
rect 96 697 97 703
rect 103 702 1959 703
rect 103 698 111 702
rect 115 698 131 702
rect 135 698 195 702
rect 199 698 275 702
rect 279 698 419 702
rect 423 698 443 702
rect 447 698 611 702
rect 615 698 635 702
rect 639 698 771 702
rect 775 698 851 702
rect 855 698 923 702
rect 927 698 1059 702
rect 1063 698 1075 702
rect 1079 698 1219 702
rect 1223 698 1267 702
rect 1271 698 1363 702
rect 1367 698 1483 702
rect 1487 698 1507 702
rect 1511 698 1651 702
rect 1655 698 1787 702
rect 1791 698 1935 702
rect 1939 698 1959 702
rect 103 697 1959 698
rect 1965 697 1966 703
rect 3810 609 3811 615
rect 3817 614 5695 615
rect 3817 610 3839 614
rect 3843 610 3887 614
rect 3891 610 4111 614
rect 4115 610 4143 614
rect 4147 610 4351 614
rect 4355 610 4407 614
rect 4411 610 4583 614
rect 4587 610 4647 614
rect 4651 610 4807 614
rect 4811 610 4879 614
rect 4883 610 5031 614
rect 5035 610 5095 614
rect 5099 610 5255 614
rect 5259 610 5311 614
rect 5315 610 5487 614
rect 5491 610 5527 614
rect 5531 610 5663 614
rect 5667 610 5695 614
rect 3817 609 5695 610
rect 5701 609 5702 615
rect 1946 597 1947 603
rect 1953 602 3811 603
rect 1953 598 1975 602
rect 1979 598 3271 602
rect 3275 598 3407 602
rect 3411 598 3543 602
rect 3547 598 3679 602
rect 3683 598 3799 602
rect 3803 598 3811 602
rect 1953 597 3811 598
rect 3817 597 3818 603
rect 84 573 85 579
rect 91 578 1947 579
rect 91 574 111 578
rect 115 574 159 578
rect 163 574 303 578
rect 307 574 375 578
rect 379 574 471 578
rect 475 574 599 578
rect 603 574 639 578
rect 643 574 799 578
rect 803 574 807 578
rect 811 574 951 578
rect 955 574 999 578
rect 1003 574 1103 578
rect 1107 574 1175 578
rect 1179 574 1247 578
rect 1251 574 1343 578
rect 1347 574 1391 578
rect 1395 574 1511 578
rect 1515 574 1535 578
rect 1539 574 1671 578
rect 1675 574 1679 578
rect 1683 574 1815 578
rect 1819 574 1935 578
rect 1939 574 1947 578
rect 91 573 1947 574
rect 1953 573 1954 579
rect 3822 481 3823 487
rect 3829 486 5707 487
rect 3829 482 3839 486
rect 3843 482 3859 486
rect 3863 482 3891 486
rect 3895 482 4115 486
rect 4119 482 4171 486
rect 4175 482 4379 486
rect 4383 482 4435 486
rect 4439 482 4619 486
rect 4623 482 4683 486
rect 4687 482 4851 486
rect 4855 482 4907 486
rect 4911 482 5067 486
rect 5071 482 5123 486
rect 5127 482 5283 486
rect 5287 482 5331 486
rect 5335 482 5499 486
rect 5503 482 5515 486
rect 5519 482 5663 486
rect 5667 482 5707 486
rect 3829 481 5707 482
rect 5713 481 5714 487
rect 1958 470 3830 471
rect 1958 467 1975 470
rect 96 461 97 467
rect 103 466 1959 467
rect 103 462 111 466
rect 115 462 131 466
rect 135 462 195 466
rect 199 462 347 466
rect 351 462 475 466
rect 479 462 571 466
rect 575 462 755 466
rect 759 462 779 466
rect 783 462 971 466
rect 975 462 1043 466
rect 1047 462 1147 466
rect 1151 462 1315 466
rect 1319 462 1331 466
rect 1335 462 1483 466
rect 1487 462 1643 466
rect 1647 462 1787 466
rect 1791 462 1935 466
rect 1939 462 1959 466
rect 103 461 1959 462
rect 1965 466 1975 467
rect 1979 466 1995 470
rect 1999 466 2155 470
rect 2159 466 2347 470
rect 2351 466 2539 470
rect 2543 466 2739 470
rect 2743 466 2931 470
rect 2935 466 3131 470
rect 3135 466 3243 470
rect 3247 466 3331 470
rect 3335 466 3379 470
rect 3383 466 3515 470
rect 3519 466 3531 470
rect 3535 466 3651 470
rect 3655 466 3799 470
rect 3803 466 3830 470
rect 1965 465 3830 466
rect 1965 461 1966 465
rect 3810 365 3811 371
rect 3817 370 5695 371
rect 3817 366 3839 370
rect 3843 366 3919 370
rect 3923 366 4007 370
rect 4011 366 4199 370
rect 4203 366 4423 370
rect 4427 366 4463 370
rect 4467 366 4679 370
rect 4683 366 4711 370
rect 4715 366 4935 370
rect 4939 366 4967 370
rect 4971 366 5151 370
rect 5155 366 5263 370
rect 5267 366 5359 370
rect 5363 366 5543 370
rect 5547 366 5663 370
rect 5667 366 5695 370
rect 3817 365 5695 366
rect 5701 365 5702 371
rect 84 349 85 355
rect 91 354 1947 355
rect 91 350 111 354
rect 115 350 223 354
rect 227 350 311 354
rect 315 350 503 354
rect 507 350 695 354
rect 699 350 783 354
rect 787 350 887 354
rect 891 350 1071 354
rect 1075 350 1079 354
rect 1083 350 1359 354
rect 1363 350 1935 354
rect 1939 350 1947 354
rect 91 349 1947 350
rect 1953 349 1954 355
rect 1946 329 1947 335
rect 1953 334 3811 335
rect 1953 330 1975 334
rect 1979 330 2023 334
rect 2027 330 2159 334
rect 2163 330 2183 334
rect 2187 330 2295 334
rect 2299 330 2375 334
rect 2379 330 2431 334
rect 2435 330 2567 334
rect 2571 330 2703 334
rect 2707 330 2767 334
rect 2771 330 2839 334
rect 2843 330 2959 334
rect 2963 330 2975 334
rect 2979 330 3111 334
rect 3115 330 3159 334
rect 3163 330 3247 334
rect 3251 330 3359 334
rect 3363 330 3383 334
rect 3387 330 3519 334
rect 3523 330 3559 334
rect 3563 330 3799 334
rect 3803 330 3811 334
rect 1953 329 3811 330
rect 3817 329 3818 335
rect 2114 252 2120 253
rect 2794 252 2800 253
rect 2114 248 2115 252
rect 2119 248 2795 252
rect 2799 248 2800 252
rect 2114 247 2120 248
rect 2794 247 2800 248
rect 96 201 97 207
rect 103 206 1959 207
rect 103 202 111 206
rect 115 202 131 206
rect 135 202 267 206
rect 271 202 283 206
rect 287 202 403 206
rect 407 202 475 206
rect 479 202 539 206
rect 543 202 667 206
rect 671 202 675 206
rect 679 202 811 206
rect 815 202 859 206
rect 863 202 947 206
rect 951 202 1051 206
rect 1055 202 1083 206
rect 1087 202 1935 206
rect 1939 202 1959 206
rect 103 201 1959 202
rect 1965 201 1966 207
rect 3822 201 3823 207
rect 3829 206 5707 207
rect 3829 202 3839 206
rect 3843 202 3859 206
rect 3863 202 3979 206
rect 3983 202 3995 206
rect 3999 202 4131 206
rect 4135 202 4171 206
rect 4175 202 4267 206
rect 4271 202 4395 206
rect 4399 202 4435 206
rect 4439 202 4627 206
rect 4631 202 4651 206
rect 4655 202 4843 206
rect 4847 202 4939 206
rect 4943 202 5067 206
rect 5071 202 5235 206
rect 5239 202 5299 206
rect 5303 202 5515 206
rect 5519 202 5663 206
rect 5667 202 5707 206
rect 3829 201 5707 202
rect 5713 201 5714 207
rect 1958 185 1959 191
rect 1965 190 3823 191
rect 1965 186 1975 190
rect 1979 186 1995 190
rect 1999 186 2131 190
rect 2135 186 2267 190
rect 2271 186 2403 190
rect 2407 186 2539 190
rect 2543 186 2675 190
rect 2679 186 2811 190
rect 2815 186 2947 190
rect 2951 186 3083 190
rect 3087 186 3219 190
rect 3223 186 3355 190
rect 3359 186 3491 190
rect 3495 186 3627 190
rect 3631 186 3799 190
rect 3803 186 3823 190
rect 1965 185 3823 186
rect 3829 185 3830 191
rect 2906 180 2912 181
rect 3750 180 3756 181
rect 2906 176 2907 180
rect 2911 176 3751 180
rect 3755 176 3756 180
rect 2906 175 2912 176
rect 3750 175 3756 176
rect 84 89 85 95
rect 91 94 1947 95
rect 91 90 111 94
rect 115 90 159 94
rect 163 90 295 94
rect 299 90 431 94
rect 435 90 567 94
rect 571 90 703 94
rect 707 90 839 94
rect 843 90 975 94
rect 979 90 1111 94
rect 1115 90 1935 94
rect 1939 90 1947 94
rect 91 89 1947 90
rect 1953 89 1954 95
rect 3810 89 3811 95
rect 3817 94 5695 95
rect 3817 90 3839 94
rect 3843 90 3887 94
rect 3891 90 4023 94
rect 4027 90 4159 94
rect 4163 90 4295 94
rect 4299 90 4463 94
rect 4467 90 4655 94
rect 4659 90 4871 94
rect 4875 90 5095 94
rect 5099 90 5327 94
rect 5331 90 5543 94
rect 5547 90 5663 94
rect 5667 90 5695 94
rect 3817 89 5695 90
rect 5701 89 5702 95
rect 1946 73 1947 79
rect 1953 78 3811 79
rect 1953 74 1975 78
rect 1979 74 2023 78
rect 2027 74 2159 78
rect 2163 74 2295 78
rect 2299 74 2431 78
rect 2435 74 2567 78
rect 2571 74 2703 78
rect 2707 74 2839 78
rect 2843 74 2975 78
rect 2979 74 3111 78
rect 3115 74 3247 78
rect 3251 74 3383 78
rect 3387 74 3519 78
rect 3523 74 3655 78
rect 3659 74 3799 78
rect 3803 74 3811 78
rect 1953 73 3811 74
rect 3817 73 3818 79
<< m5c >>
rect 97 5753 103 5759
rect 1959 5753 1965 5759
rect 1947 5717 1953 5723
rect 3811 5717 3817 5723
rect 3823 5669 3829 5675
rect 5707 5669 5713 5675
rect 85 5641 91 5647
rect 1947 5641 1953 5647
rect 1959 5597 1965 5603
rect 3823 5597 3829 5603
rect 97 5529 103 5535
rect 1959 5529 1965 5535
rect 3811 5525 3817 5531
rect 5695 5525 5701 5531
rect 1947 5485 1953 5491
rect 3811 5485 3817 5491
rect 85 5397 91 5403
rect 1947 5397 1953 5403
rect 3823 5389 3829 5395
rect 5707 5389 5713 5395
rect 1959 5349 1965 5355
rect 3823 5349 3829 5355
rect 97 5281 103 5287
rect 1959 5281 1965 5287
rect 3811 5273 3817 5279
rect 5695 5273 5701 5279
rect 1947 5237 1953 5243
rect 3811 5237 3817 5243
rect 85 5157 91 5163
rect 1947 5157 1953 5163
rect 3823 5141 3829 5147
rect 5707 5141 5713 5147
rect 1959 5125 1965 5131
rect 3823 5125 3829 5131
rect 97 5041 103 5047
rect 1959 5041 1965 5047
rect 3811 5013 3817 5019
rect 5695 5013 5701 5019
rect 1947 4981 1953 4987
rect 3811 4981 3817 4987
rect 85 4905 91 4911
rect 1947 4905 1953 4911
rect 3823 4877 3829 4883
rect 5707 4877 5713 4883
rect 1959 4861 1965 4867
rect 3823 4861 3829 4867
rect 97 4781 103 4787
rect 1959 4781 1965 4787
rect 3811 4765 3817 4771
rect 5695 4765 5701 4771
rect 1947 4745 1953 4751
rect 3811 4745 3817 4751
rect 85 4661 91 4667
rect 1947 4661 1953 4667
rect 3823 4629 3829 4635
rect 5707 4629 5713 4635
rect 1959 4601 1965 4607
rect 3823 4601 3829 4607
rect 97 4541 103 4547
rect 1959 4541 1965 4547
rect 3811 4505 3817 4511
rect 5695 4505 5701 4511
rect 1947 4481 1953 4487
rect 3811 4481 3817 4487
rect 85 4429 91 4435
rect 1947 4429 1953 4435
rect 3823 4369 3829 4375
rect 5707 4369 5713 4375
rect 1959 4357 1965 4363
rect 3823 4357 3829 4363
rect 97 4297 103 4303
rect 1959 4297 1965 4303
rect 3811 4257 3817 4263
rect 5695 4257 5701 4263
rect 1947 4217 1953 4223
rect 3811 4217 3817 4223
rect 85 4181 91 4187
rect 1947 4181 1953 4187
rect 1959 4105 1965 4111
rect 3823 4105 3829 4111
rect 97 4069 103 4075
rect 1959 4069 1965 4075
rect 1947 3985 1953 3991
rect 3811 3985 3817 3991
rect 3811 3973 3817 3979
rect 5695 3973 5701 3979
rect 85 3953 91 3959
rect 1947 3953 1953 3959
rect 1959 3865 1965 3871
rect 3823 3865 3829 3871
rect 3823 3853 3829 3859
rect 5707 3853 5713 3859
rect 97 3833 103 3839
rect 1959 3833 1965 3839
rect 1947 3749 1953 3755
rect 3811 3749 3817 3755
rect 85 3717 91 3723
rect 1947 3717 1953 3723
rect 3811 3713 3817 3719
rect 5695 3713 5701 3719
rect 1959 3629 1965 3635
rect 3823 3629 3829 3635
rect 3823 3601 3829 3607
rect 5707 3601 5713 3607
rect 97 3593 103 3599
rect 1959 3593 1965 3599
rect 1947 3477 1953 3483
rect 3811 3477 3817 3483
rect 85 3457 91 3463
rect 1947 3457 1953 3463
rect 3823 3369 3829 3375
rect 5707 3369 5713 3375
rect 1959 3357 1965 3363
rect 3823 3357 3829 3363
rect 97 3341 103 3347
rect 1959 3341 1965 3347
rect 1947 3245 1953 3251
rect 3811 3245 3817 3251
rect 85 3229 91 3235
rect 1947 3229 1953 3235
rect 3811 3233 3817 3239
rect 5695 3233 5701 3239
rect 1959 3133 1965 3139
rect 3823 3133 3829 3139
rect 3823 3117 3829 3123
rect 5707 3117 5713 3123
rect 97 3105 103 3111
rect 1959 3105 1965 3111
rect 1947 3013 1953 3019
rect 3811 3013 3817 3019
rect 85 2989 91 2995
rect 1947 2989 1953 2995
rect 3811 2981 3817 2987
rect 5695 2981 5701 2987
rect 1959 2897 1965 2903
rect 3823 2897 3829 2903
rect 97 2873 103 2879
rect 1959 2873 1965 2879
rect 3823 2853 3829 2859
rect 5707 2853 5713 2859
rect 1947 2781 1953 2787
rect 3811 2781 3817 2787
rect 85 2757 91 2763
rect 1947 2757 1953 2763
rect 3811 2729 3817 2735
rect 5695 2729 5701 2735
rect 1959 2661 1965 2667
rect 3823 2661 3829 2667
rect 97 2645 103 2651
rect 1959 2645 1965 2651
rect 3823 2617 3829 2623
rect 5707 2617 5713 2623
rect 1947 2549 1953 2555
rect 3811 2549 3817 2555
rect 85 2533 91 2539
rect 1947 2533 1953 2539
rect 3811 2501 3817 2507
rect 5695 2501 5701 2507
rect 97 2417 103 2423
rect 1959 2417 1965 2423
rect 3823 2389 3829 2395
rect 5707 2389 5713 2395
rect 1947 2297 1953 2303
rect 3811 2297 3817 2303
rect 85 2289 91 2295
rect 1947 2289 1953 2295
rect 3811 2253 3817 2259
rect 5695 2253 5701 2259
rect 1959 2177 1965 2183
rect 3823 2177 3829 2183
rect 97 2165 103 2171
rect 1959 2165 1965 2171
rect 3823 2125 3829 2131
rect 5707 2125 5713 2131
rect 1947 2057 1953 2063
rect 3811 2057 3817 2063
rect 85 2049 91 2055
rect 1947 2049 1953 2055
rect 3811 2013 3817 2019
rect 5695 2013 5701 2019
rect 97 1929 103 1935
rect 1959 1929 1965 1935
rect 3823 1901 3829 1907
rect 5707 1901 5713 1907
rect 1947 1817 1953 1823
rect 3811 1817 3817 1823
rect 85 1801 91 1807
rect 1947 1801 1953 1807
rect 3811 1781 3817 1787
rect 5695 1781 5701 1787
rect 97 1685 103 1691
rect 1959 1685 1965 1691
rect 1959 1673 1965 1679
rect 3823 1673 3829 1679
rect 3823 1665 3829 1671
rect 5707 1665 5713 1671
rect 85 1553 91 1559
rect 1947 1553 1953 1559
rect 3811 1549 3817 1555
rect 5695 1549 5701 1555
rect 3823 1437 3829 1443
rect 5707 1437 5713 1443
rect 97 1429 103 1435
rect 1959 1429 1965 1435
rect 3811 1325 3817 1331
rect 5695 1325 5701 1331
rect 85 1317 91 1323
rect 1947 1317 1953 1323
rect 97 1193 103 1199
rect 1959 1193 1965 1199
rect 85 1073 91 1079
rect 1947 1073 1953 1079
rect 97 953 103 959
rect 1959 953 1965 959
rect 1947 845 1953 851
rect 3811 845 3817 851
rect 85 817 91 823
rect 1947 817 1953 823
rect 3823 729 3829 735
rect 5707 729 5713 735
rect 1959 717 1965 723
rect 3823 717 3829 723
rect 97 697 103 703
rect 1959 697 1965 703
rect 3811 609 3817 615
rect 5695 609 5701 615
rect 1947 597 1953 603
rect 3811 597 3817 603
rect 85 573 91 579
rect 1947 573 1953 579
rect 3823 481 3829 487
rect 5707 481 5713 487
rect 97 461 103 467
rect 1959 461 1965 467
rect 3811 365 3817 371
rect 5695 365 5701 371
rect 85 349 91 355
rect 1947 349 1953 355
rect 1947 329 1953 335
rect 3811 329 3817 335
rect 97 201 103 207
rect 1959 201 1965 207
rect 3823 201 3829 207
rect 5707 201 5713 207
rect 1959 185 1965 191
rect 3823 185 3829 191
rect 85 89 91 95
rect 1947 89 1953 95
rect 3811 89 3817 95
rect 5695 89 5701 95
rect 1947 73 1953 79
rect 3811 73 3817 79
<< m5 >>
rect 84 5647 92 5760
rect 84 5641 85 5647
rect 91 5641 92 5647
rect 84 5403 92 5641
rect 84 5397 85 5403
rect 91 5397 92 5403
rect 84 5163 92 5397
rect 84 5157 85 5163
rect 91 5157 92 5163
rect 84 4911 92 5157
rect 84 4905 85 4911
rect 91 4905 92 4911
rect 84 4667 92 4905
rect 84 4661 85 4667
rect 91 4661 92 4667
rect 84 4435 92 4661
rect 84 4429 85 4435
rect 91 4429 92 4435
rect 84 4187 92 4429
rect 84 4181 85 4187
rect 91 4181 92 4187
rect 84 3959 92 4181
rect 84 3953 85 3959
rect 91 3953 92 3959
rect 84 3723 92 3953
rect 84 3717 85 3723
rect 91 3717 92 3723
rect 84 3463 92 3717
rect 84 3457 85 3463
rect 91 3457 92 3463
rect 84 3235 92 3457
rect 84 3229 85 3235
rect 91 3229 92 3235
rect 84 2995 92 3229
rect 84 2989 85 2995
rect 91 2989 92 2995
rect 84 2763 92 2989
rect 84 2757 85 2763
rect 91 2757 92 2763
rect 84 2539 92 2757
rect 84 2533 85 2539
rect 91 2533 92 2539
rect 84 2295 92 2533
rect 84 2289 85 2295
rect 91 2289 92 2295
rect 84 2055 92 2289
rect 84 2049 85 2055
rect 91 2049 92 2055
rect 84 1807 92 2049
rect 84 1801 85 1807
rect 91 1801 92 1807
rect 84 1559 92 1801
rect 84 1553 85 1559
rect 91 1553 92 1559
rect 84 1323 92 1553
rect 84 1317 85 1323
rect 91 1317 92 1323
rect 84 1079 92 1317
rect 84 1073 85 1079
rect 91 1073 92 1079
rect 84 823 92 1073
rect 84 817 85 823
rect 91 817 92 823
rect 84 579 92 817
rect 84 573 85 579
rect 91 573 92 579
rect 84 355 92 573
rect 84 349 85 355
rect 91 349 92 355
rect 84 95 92 349
rect 84 89 85 95
rect 91 89 92 95
rect 84 72 92 89
rect 96 5759 104 5760
rect 96 5753 97 5759
rect 103 5753 104 5759
rect 96 5535 104 5753
rect 96 5529 97 5535
rect 103 5529 104 5535
rect 96 5287 104 5529
rect 96 5281 97 5287
rect 103 5281 104 5287
rect 96 5047 104 5281
rect 96 5041 97 5047
rect 103 5041 104 5047
rect 96 4787 104 5041
rect 96 4781 97 4787
rect 103 4781 104 4787
rect 96 4547 104 4781
rect 96 4541 97 4547
rect 103 4541 104 4547
rect 96 4303 104 4541
rect 96 4297 97 4303
rect 103 4297 104 4303
rect 96 4075 104 4297
rect 96 4069 97 4075
rect 103 4069 104 4075
rect 96 3839 104 4069
rect 96 3833 97 3839
rect 103 3833 104 3839
rect 96 3599 104 3833
rect 96 3593 97 3599
rect 103 3593 104 3599
rect 96 3347 104 3593
rect 96 3341 97 3347
rect 103 3341 104 3347
rect 96 3111 104 3341
rect 96 3105 97 3111
rect 103 3105 104 3111
rect 96 2879 104 3105
rect 96 2873 97 2879
rect 103 2873 104 2879
rect 96 2651 104 2873
rect 96 2645 97 2651
rect 103 2645 104 2651
rect 96 2423 104 2645
rect 96 2417 97 2423
rect 103 2417 104 2423
rect 96 2171 104 2417
rect 96 2165 97 2171
rect 103 2165 104 2171
rect 96 1935 104 2165
rect 96 1929 97 1935
rect 103 1929 104 1935
rect 96 1691 104 1929
rect 96 1685 97 1691
rect 103 1685 104 1691
rect 96 1435 104 1685
rect 96 1429 97 1435
rect 103 1429 104 1435
rect 96 1199 104 1429
rect 96 1193 97 1199
rect 103 1193 104 1199
rect 96 959 104 1193
rect 96 953 97 959
rect 103 953 104 959
rect 96 703 104 953
rect 96 697 97 703
rect 103 697 104 703
rect 96 467 104 697
rect 96 461 97 467
rect 103 461 104 467
rect 96 207 104 461
rect 96 201 97 207
rect 103 201 104 207
rect 96 72 104 201
rect 1946 5723 1954 5760
rect 1946 5717 1947 5723
rect 1953 5717 1954 5723
rect 1946 5647 1954 5717
rect 1946 5641 1947 5647
rect 1953 5641 1954 5647
rect 1946 5491 1954 5641
rect 1946 5485 1947 5491
rect 1953 5485 1954 5491
rect 1946 5403 1954 5485
rect 1946 5397 1947 5403
rect 1953 5397 1954 5403
rect 1946 5243 1954 5397
rect 1946 5237 1947 5243
rect 1953 5237 1954 5243
rect 1946 5163 1954 5237
rect 1946 5157 1947 5163
rect 1953 5157 1954 5163
rect 1946 4987 1954 5157
rect 1946 4981 1947 4987
rect 1953 4981 1954 4987
rect 1946 4911 1954 4981
rect 1946 4905 1947 4911
rect 1953 4905 1954 4911
rect 1946 4751 1954 4905
rect 1946 4745 1947 4751
rect 1953 4745 1954 4751
rect 1946 4667 1954 4745
rect 1946 4661 1947 4667
rect 1953 4661 1954 4667
rect 1946 4487 1954 4661
rect 1946 4481 1947 4487
rect 1953 4481 1954 4487
rect 1946 4435 1954 4481
rect 1946 4429 1947 4435
rect 1953 4429 1954 4435
rect 1946 4223 1954 4429
rect 1946 4217 1947 4223
rect 1953 4217 1954 4223
rect 1946 4187 1954 4217
rect 1946 4181 1947 4187
rect 1953 4181 1954 4187
rect 1946 3991 1954 4181
rect 1946 3985 1947 3991
rect 1953 3985 1954 3991
rect 1946 3959 1954 3985
rect 1946 3953 1947 3959
rect 1953 3953 1954 3959
rect 1946 3755 1954 3953
rect 1946 3749 1947 3755
rect 1953 3749 1954 3755
rect 1946 3723 1954 3749
rect 1946 3717 1947 3723
rect 1953 3717 1954 3723
rect 1946 3483 1954 3717
rect 1946 3477 1947 3483
rect 1953 3477 1954 3483
rect 1946 3463 1954 3477
rect 1946 3457 1947 3463
rect 1953 3457 1954 3463
rect 1946 3251 1954 3457
rect 1946 3245 1947 3251
rect 1953 3245 1954 3251
rect 1946 3235 1954 3245
rect 1946 3229 1947 3235
rect 1953 3229 1954 3235
rect 1946 3019 1954 3229
rect 1946 3013 1947 3019
rect 1953 3013 1954 3019
rect 1946 2995 1954 3013
rect 1946 2989 1947 2995
rect 1953 2989 1954 2995
rect 1946 2787 1954 2989
rect 1946 2781 1947 2787
rect 1953 2781 1954 2787
rect 1946 2763 1954 2781
rect 1946 2757 1947 2763
rect 1953 2757 1954 2763
rect 1946 2555 1954 2757
rect 1946 2549 1947 2555
rect 1953 2549 1954 2555
rect 1946 2539 1954 2549
rect 1946 2533 1947 2539
rect 1953 2533 1954 2539
rect 1946 2303 1954 2533
rect 1946 2297 1947 2303
rect 1953 2297 1954 2303
rect 1946 2295 1954 2297
rect 1946 2289 1947 2295
rect 1953 2289 1954 2295
rect 1946 2063 1954 2289
rect 1946 2057 1947 2063
rect 1953 2057 1954 2063
rect 1946 2055 1954 2057
rect 1946 2049 1947 2055
rect 1953 2049 1954 2055
rect 1946 1823 1954 2049
rect 1946 1817 1947 1823
rect 1953 1817 1954 1823
rect 1946 1807 1954 1817
rect 1946 1801 1947 1807
rect 1953 1801 1954 1807
rect 1946 1559 1954 1801
rect 1946 1553 1947 1559
rect 1953 1553 1954 1559
rect 1946 1323 1954 1553
rect 1946 1317 1947 1323
rect 1953 1317 1954 1323
rect 1946 1079 1954 1317
rect 1946 1073 1947 1079
rect 1953 1073 1954 1079
rect 1946 851 1954 1073
rect 1946 845 1947 851
rect 1953 845 1954 851
rect 1946 823 1954 845
rect 1946 817 1947 823
rect 1953 817 1954 823
rect 1946 603 1954 817
rect 1946 597 1947 603
rect 1953 597 1954 603
rect 1946 579 1954 597
rect 1946 573 1947 579
rect 1953 573 1954 579
rect 1946 355 1954 573
rect 1946 349 1947 355
rect 1953 349 1954 355
rect 1946 335 1954 349
rect 1946 329 1947 335
rect 1953 329 1954 335
rect 1946 95 1954 329
rect 1946 89 1947 95
rect 1953 89 1954 95
rect 1946 79 1954 89
rect 1946 73 1947 79
rect 1953 73 1954 79
rect 1946 72 1954 73
rect 1958 5759 1966 5760
rect 1958 5753 1959 5759
rect 1965 5753 1966 5759
rect 1958 5603 1966 5753
rect 1958 5597 1959 5603
rect 1965 5597 1966 5603
rect 1958 5535 1966 5597
rect 1958 5529 1959 5535
rect 1965 5529 1966 5535
rect 1958 5355 1966 5529
rect 1958 5349 1959 5355
rect 1965 5349 1966 5355
rect 1958 5287 1966 5349
rect 1958 5281 1959 5287
rect 1965 5281 1966 5287
rect 1958 5131 1966 5281
rect 1958 5125 1959 5131
rect 1965 5125 1966 5131
rect 1958 5047 1966 5125
rect 1958 5041 1959 5047
rect 1965 5041 1966 5047
rect 1958 4867 1966 5041
rect 1958 4861 1959 4867
rect 1965 4861 1966 4867
rect 1958 4787 1966 4861
rect 1958 4781 1959 4787
rect 1965 4781 1966 4787
rect 1958 4607 1966 4781
rect 1958 4601 1959 4607
rect 1965 4601 1966 4607
rect 1958 4547 1966 4601
rect 1958 4541 1959 4547
rect 1965 4541 1966 4547
rect 1958 4363 1966 4541
rect 1958 4357 1959 4363
rect 1965 4357 1966 4363
rect 1958 4303 1966 4357
rect 1958 4297 1959 4303
rect 1965 4297 1966 4303
rect 1958 4111 1966 4297
rect 1958 4105 1959 4111
rect 1965 4105 1966 4111
rect 1958 4075 1966 4105
rect 1958 4069 1959 4075
rect 1965 4069 1966 4075
rect 1958 3871 1966 4069
rect 1958 3865 1959 3871
rect 1965 3865 1966 3871
rect 1958 3839 1966 3865
rect 1958 3833 1959 3839
rect 1965 3833 1966 3839
rect 1958 3635 1966 3833
rect 1958 3629 1959 3635
rect 1965 3629 1966 3635
rect 1958 3599 1966 3629
rect 1958 3593 1959 3599
rect 1965 3593 1966 3599
rect 1958 3363 1966 3593
rect 1958 3357 1959 3363
rect 1965 3357 1966 3363
rect 1958 3347 1966 3357
rect 1958 3341 1959 3347
rect 1965 3341 1966 3347
rect 1958 3139 1966 3341
rect 1958 3133 1959 3139
rect 1965 3133 1966 3139
rect 1958 3111 1966 3133
rect 1958 3105 1959 3111
rect 1965 3105 1966 3111
rect 1958 2903 1966 3105
rect 1958 2897 1959 2903
rect 1965 2897 1966 2903
rect 1958 2879 1966 2897
rect 1958 2873 1959 2879
rect 1965 2873 1966 2879
rect 1958 2667 1966 2873
rect 1958 2661 1959 2667
rect 1965 2661 1966 2667
rect 1958 2651 1966 2661
rect 1958 2645 1959 2651
rect 1965 2645 1966 2651
rect 1958 2423 1966 2645
rect 1958 2417 1959 2423
rect 1965 2417 1966 2423
rect 1958 2183 1966 2417
rect 1958 2177 1959 2183
rect 1965 2177 1966 2183
rect 1958 2171 1966 2177
rect 1958 2165 1959 2171
rect 1965 2165 1966 2171
rect 1958 1935 1966 2165
rect 1958 1929 1959 1935
rect 1965 1929 1966 1935
rect 1958 1691 1966 1929
rect 1958 1685 1959 1691
rect 1965 1685 1966 1691
rect 1958 1679 1966 1685
rect 1958 1673 1959 1679
rect 1965 1673 1966 1679
rect 1958 1435 1966 1673
rect 1958 1429 1959 1435
rect 1965 1429 1966 1435
rect 1958 1199 1966 1429
rect 1958 1193 1959 1199
rect 1965 1193 1966 1199
rect 1958 959 1966 1193
rect 1958 953 1959 959
rect 1965 953 1966 959
rect 1958 723 1966 953
rect 1958 717 1959 723
rect 1965 717 1966 723
rect 1958 703 1966 717
rect 1958 697 1959 703
rect 1965 697 1966 703
rect 1958 467 1966 697
rect 1958 461 1959 467
rect 1965 461 1966 467
rect 1958 207 1966 461
rect 1958 201 1959 207
rect 1965 201 1966 207
rect 1958 191 1966 201
rect 1958 185 1959 191
rect 1965 185 1966 191
rect 1958 72 1966 185
rect 3810 5723 3818 5760
rect 3810 5717 3811 5723
rect 3817 5717 3818 5723
rect 3810 5531 3818 5717
rect 3810 5525 3811 5531
rect 3817 5525 3818 5531
rect 3810 5491 3818 5525
rect 3810 5485 3811 5491
rect 3817 5485 3818 5491
rect 3810 5279 3818 5485
rect 3810 5273 3811 5279
rect 3817 5273 3818 5279
rect 3810 5243 3818 5273
rect 3810 5237 3811 5243
rect 3817 5237 3818 5243
rect 3810 5019 3818 5237
rect 3810 5013 3811 5019
rect 3817 5013 3818 5019
rect 3810 4987 3818 5013
rect 3810 4981 3811 4987
rect 3817 4981 3818 4987
rect 3810 4771 3818 4981
rect 3810 4765 3811 4771
rect 3817 4765 3818 4771
rect 3810 4751 3818 4765
rect 3810 4745 3811 4751
rect 3817 4745 3818 4751
rect 3810 4511 3818 4745
rect 3810 4505 3811 4511
rect 3817 4505 3818 4511
rect 3810 4487 3818 4505
rect 3810 4481 3811 4487
rect 3817 4481 3818 4487
rect 3810 4263 3818 4481
rect 3810 4257 3811 4263
rect 3817 4257 3818 4263
rect 3810 4223 3818 4257
rect 3810 4217 3811 4223
rect 3817 4217 3818 4223
rect 3810 3991 3818 4217
rect 3810 3985 3811 3991
rect 3817 3985 3818 3991
rect 3810 3979 3818 3985
rect 3810 3973 3811 3979
rect 3817 3973 3818 3979
rect 3810 3755 3818 3973
rect 3810 3749 3811 3755
rect 3817 3749 3818 3755
rect 3810 3719 3818 3749
rect 3810 3713 3811 3719
rect 3817 3713 3818 3719
rect 3810 3483 3818 3713
rect 3810 3477 3811 3483
rect 3817 3477 3818 3483
rect 3810 3251 3818 3477
rect 3810 3245 3811 3251
rect 3817 3245 3818 3251
rect 3810 3239 3818 3245
rect 3810 3233 3811 3239
rect 3817 3233 3818 3239
rect 3810 3019 3818 3233
rect 3810 3013 3811 3019
rect 3817 3013 3818 3019
rect 3810 2987 3818 3013
rect 3810 2981 3811 2987
rect 3817 2981 3818 2987
rect 3810 2787 3818 2981
rect 3810 2781 3811 2787
rect 3817 2781 3818 2787
rect 3810 2735 3818 2781
rect 3810 2729 3811 2735
rect 3817 2729 3818 2735
rect 3810 2555 3818 2729
rect 3810 2549 3811 2555
rect 3817 2549 3818 2555
rect 3810 2507 3818 2549
rect 3810 2501 3811 2507
rect 3817 2501 3818 2507
rect 3810 2303 3818 2501
rect 3810 2297 3811 2303
rect 3817 2297 3818 2303
rect 3810 2259 3818 2297
rect 3810 2253 3811 2259
rect 3817 2253 3818 2259
rect 3810 2063 3818 2253
rect 3810 2057 3811 2063
rect 3817 2057 3818 2063
rect 3810 2019 3818 2057
rect 3810 2013 3811 2019
rect 3817 2013 3818 2019
rect 3810 1823 3818 2013
rect 3810 1817 3811 1823
rect 3817 1817 3818 1823
rect 3810 1787 3818 1817
rect 3810 1781 3811 1787
rect 3817 1781 3818 1787
rect 3810 1555 3818 1781
rect 3810 1549 3811 1555
rect 3817 1549 3818 1555
rect 3810 1331 3818 1549
rect 3810 1325 3811 1331
rect 3817 1325 3818 1331
rect 3810 851 3818 1325
rect 3810 845 3811 851
rect 3817 845 3818 851
rect 3810 615 3818 845
rect 3810 609 3811 615
rect 3817 609 3818 615
rect 3810 603 3818 609
rect 3810 597 3811 603
rect 3817 597 3818 603
rect 3810 371 3818 597
rect 3810 365 3811 371
rect 3817 365 3818 371
rect 3810 335 3818 365
rect 3810 329 3811 335
rect 3817 329 3818 335
rect 3810 95 3818 329
rect 3810 89 3811 95
rect 3817 89 3818 95
rect 3810 79 3818 89
rect 3810 73 3811 79
rect 3817 73 3818 79
rect 3810 72 3818 73
rect 3822 5675 3830 5760
rect 3822 5669 3823 5675
rect 3829 5669 3830 5675
rect 3822 5603 3830 5669
rect 3822 5597 3823 5603
rect 3829 5597 3830 5603
rect 3822 5395 3830 5597
rect 3822 5389 3823 5395
rect 3829 5389 3830 5395
rect 3822 5355 3830 5389
rect 3822 5349 3823 5355
rect 3829 5349 3830 5355
rect 3822 5147 3830 5349
rect 3822 5141 3823 5147
rect 3829 5141 3830 5147
rect 3822 5131 3830 5141
rect 3822 5125 3823 5131
rect 3829 5125 3830 5131
rect 3822 4883 3830 5125
rect 3822 4877 3823 4883
rect 3829 4877 3830 4883
rect 3822 4867 3830 4877
rect 3822 4861 3823 4867
rect 3829 4861 3830 4867
rect 3822 4635 3830 4861
rect 3822 4629 3823 4635
rect 3829 4629 3830 4635
rect 3822 4607 3830 4629
rect 3822 4601 3823 4607
rect 3829 4601 3830 4607
rect 3822 4375 3830 4601
rect 3822 4369 3823 4375
rect 3829 4369 3830 4375
rect 3822 4363 3830 4369
rect 3822 4357 3823 4363
rect 3829 4357 3830 4363
rect 3822 4111 3830 4357
rect 3822 4105 3823 4111
rect 3829 4105 3830 4111
rect 3822 3871 3830 4105
rect 3822 3865 3823 3871
rect 3829 3865 3830 3871
rect 3822 3859 3830 3865
rect 3822 3853 3823 3859
rect 3829 3853 3830 3859
rect 3822 3635 3830 3853
rect 3822 3629 3823 3635
rect 3829 3629 3830 3635
rect 3822 3607 3830 3629
rect 3822 3601 3823 3607
rect 3829 3601 3830 3607
rect 3822 3375 3830 3601
rect 3822 3369 3823 3375
rect 3829 3369 3830 3375
rect 3822 3363 3830 3369
rect 3822 3357 3823 3363
rect 3829 3357 3830 3363
rect 3822 3139 3830 3357
rect 3822 3133 3823 3139
rect 3829 3133 3830 3139
rect 3822 3123 3830 3133
rect 3822 3117 3823 3123
rect 3829 3117 3830 3123
rect 3822 2903 3830 3117
rect 3822 2897 3823 2903
rect 3829 2897 3830 2903
rect 3822 2859 3830 2897
rect 3822 2853 3823 2859
rect 3829 2853 3830 2859
rect 3822 2667 3830 2853
rect 3822 2661 3823 2667
rect 3829 2661 3830 2667
rect 3822 2623 3830 2661
rect 3822 2617 3823 2623
rect 3829 2617 3830 2623
rect 3822 2395 3830 2617
rect 3822 2389 3823 2395
rect 3829 2389 3830 2395
rect 3822 2183 3830 2389
rect 3822 2177 3823 2183
rect 3829 2177 3830 2183
rect 3822 2131 3830 2177
rect 3822 2125 3823 2131
rect 3829 2125 3830 2131
rect 3822 1907 3830 2125
rect 3822 1901 3823 1907
rect 3829 1901 3830 1907
rect 3822 1679 3830 1901
rect 3822 1673 3823 1679
rect 3829 1673 3830 1679
rect 3822 1671 3830 1673
rect 3822 1665 3823 1671
rect 3829 1665 3830 1671
rect 3822 1443 3830 1665
rect 3822 1437 3823 1443
rect 3829 1437 3830 1443
rect 3822 735 3830 1437
rect 3822 729 3823 735
rect 3829 729 3830 735
rect 3822 723 3830 729
rect 3822 717 3823 723
rect 3829 717 3830 723
rect 3822 487 3830 717
rect 3822 481 3823 487
rect 3829 481 3830 487
rect 3822 207 3830 481
rect 3822 201 3823 207
rect 3829 201 3830 207
rect 3822 191 3830 201
rect 3822 185 3823 191
rect 3829 185 3830 191
rect 3822 72 3830 185
rect 5694 5531 5702 5760
rect 5694 5525 5695 5531
rect 5701 5525 5702 5531
rect 5694 5279 5702 5525
rect 5694 5273 5695 5279
rect 5701 5273 5702 5279
rect 5694 5019 5702 5273
rect 5694 5013 5695 5019
rect 5701 5013 5702 5019
rect 5694 4771 5702 5013
rect 5694 4765 5695 4771
rect 5701 4765 5702 4771
rect 5694 4511 5702 4765
rect 5694 4505 5695 4511
rect 5701 4505 5702 4511
rect 5694 4263 5702 4505
rect 5694 4257 5695 4263
rect 5701 4257 5702 4263
rect 5694 3979 5702 4257
rect 5694 3973 5695 3979
rect 5701 3973 5702 3979
rect 5694 3719 5702 3973
rect 5694 3713 5695 3719
rect 5701 3713 5702 3719
rect 5694 3239 5702 3713
rect 5694 3233 5695 3239
rect 5701 3233 5702 3239
rect 5694 2987 5702 3233
rect 5694 2981 5695 2987
rect 5701 2981 5702 2987
rect 5694 2735 5702 2981
rect 5694 2729 5695 2735
rect 5701 2729 5702 2735
rect 5694 2507 5702 2729
rect 5694 2501 5695 2507
rect 5701 2501 5702 2507
rect 5694 2259 5702 2501
rect 5694 2253 5695 2259
rect 5701 2253 5702 2259
rect 5694 2019 5702 2253
rect 5694 2013 5695 2019
rect 5701 2013 5702 2019
rect 5694 1787 5702 2013
rect 5694 1781 5695 1787
rect 5701 1781 5702 1787
rect 5694 1555 5702 1781
rect 5694 1549 5695 1555
rect 5701 1549 5702 1555
rect 5694 1331 5702 1549
rect 5694 1325 5695 1331
rect 5701 1325 5702 1331
rect 5694 615 5702 1325
rect 5694 609 5695 615
rect 5701 609 5702 615
rect 5694 371 5702 609
rect 5694 365 5695 371
rect 5701 365 5702 371
rect 5694 95 5702 365
rect 5694 89 5695 95
rect 5701 89 5702 95
rect 5694 72 5702 89
rect 5706 5675 5714 5760
rect 5706 5669 5707 5675
rect 5713 5669 5714 5675
rect 5706 5395 5714 5669
rect 5706 5389 5707 5395
rect 5713 5389 5714 5395
rect 5706 5147 5714 5389
rect 5706 5141 5707 5147
rect 5713 5141 5714 5147
rect 5706 4883 5714 5141
rect 5706 4877 5707 4883
rect 5713 4877 5714 4883
rect 5706 4635 5714 4877
rect 5706 4629 5707 4635
rect 5713 4629 5714 4635
rect 5706 4375 5714 4629
rect 5706 4369 5707 4375
rect 5713 4369 5714 4375
rect 5706 3859 5714 4369
rect 5706 3853 5707 3859
rect 5713 3853 5714 3859
rect 5706 3607 5714 3853
rect 5706 3601 5707 3607
rect 5713 3601 5714 3607
rect 5706 3375 5714 3601
rect 5706 3369 5707 3375
rect 5713 3369 5714 3375
rect 5706 3123 5714 3369
rect 5706 3117 5707 3123
rect 5713 3117 5714 3123
rect 5706 2859 5714 3117
rect 5706 2853 5707 2859
rect 5713 2853 5714 2859
rect 5706 2623 5714 2853
rect 5706 2617 5707 2623
rect 5713 2617 5714 2623
rect 5706 2395 5714 2617
rect 5706 2389 5707 2395
rect 5713 2389 5714 2395
rect 5706 2131 5714 2389
rect 5706 2125 5707 2131
rect 5713 2125 5714 2131
rect 5706 1907 5714 2125
rect 5706 1901 5707 1907
rect 5713 1901 5714 1907
rect 5706 1671 5714 1901
rect 5706 1665 5707 1671
rect 5713 1665 5714 1671
rect 5706 1443 5714 1665
rect 5706 1437 5707 1443
rect 5713 1437 5714 1443
rect 5706 735 5714 1437
rect 5706 729 5707 735
rect 5713 729 5714 735
rect 5706 487 5714 729
rect 5706 481 5707 487
rect 5713 481 5714 487
rect 5706 207 5714 481
rect 5706 201 5707 207
rect 5713 201 5714 207
rect 5706 72 5714 201
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__275
timestamp 1731220505
transform 1 0 5656 0 1 5584
box 7 3 12 24
use welltap_svt  __well_tap__274
timestamp 1731220505
transform 1 0 3832 0 1 5584
box 7 3 12 24
use welltap_svt  __well_tap__273
timestamp 1731220505
transform 1 0 5656 0 -1 5504
box 7 3 12 24
use welltap_svt  __well_tap__272
timestamp 1731220505
transform 1 0 3832 0 -1 5504
box 7 3 12 24
use welltap_svt  __well_tap__271
timestamp 1731220505
transform 1 0 5656 0 1 5304
box 7 3 12 24
use welltap_svt  __well_tap__270
timestamp 1731220505
transform 1 0 3832 0 1 5304
box 7 3 12 24
use welltap_svt  __well_tap__269
timestamp 1731220505
transform 1 0 5656 0 -1 5252
box 7 3 12 24
use welltap_svt  __well_tap__268
timestamp 1731220505
transform 1 0 3832 0 -1 5252
box 7 3 12 24
use welltap_svt  __well_tap__267
timestamp 1731220505
transform 1 0 5656 0 1 5056
box 7 3 12 24
use welltap_svt  __well_tap__266
timestamp 1731220505
transform 1 0 3832 0 1 5056
box 7 3 12 24
use welltap_svt  __well_tap__265
timestamp 1731220505
transform 1 0 5656 0 -1 4992
box 7 3 12 24
use welltap_svt  __well_tap__264
timestamp 1731220505
transform 1 0 3832 0 -1 4992
box 7 3 12 24
use welltap_svt  __well_tap__263
timestamp 1731220505
transform 1 0 5656 0 1 4792
box 7 3 12 24
use welltap_svt  __well_tap__262
timestamp 1731220505
transform 1 0 3832 0 1 4792
box 7 3 12 24
use welltap_svt  __well_tap__261
timestamp 1731220505
transform 1 0 5656 0 -1 4744
box 7 3 12 24
use welltap_svt  __well_tap__260
timestamp 1731220505
transform 1 0 3832 0 -1 4744
box 7 3 12 24
use welltap_svt  __well_tap__259
timestamp 1731220505
transform 1 0 5656 0 1 4544
box 7 3 12 24
use welltap_svt  __well_tap__258
timestamp 1731220505
transform 1 0 3832 0 1 4544
box 7 3 12 24
use welltap_svt  __well_tap__257
timestamp 1731220505
transform 1 0 5656 0 -1 4484
box 7 3 12 24
use welltap_svt  __well_tap__256
timestamp 1731220505
transform 1 0 3832 0 -1 4484
box 7 3 12 24
use welltap_svt  __well_tap__255
timestamp 1731220505
transform 1 0 5656 0 1 4284
box 7 3 12 24
use welltap_svt  __well_tap__254
timestamp 1731220505
transform 1 0 3832 0 1 4284
box 7 3 12 24
use welltap_svt  __well_tap__253
timestamp 1731220505
transform 1 0 5656 0 -1 4236
box 7 3 12 24
use welltap_svt  __well_tap__252
timestamp 1731220505
transform 1 0 3832 0 -1 4236
box 7 3 12 24
use welltap_svt  __well_tap__251
timestamp 1731220505
transform 1 0 5656 0 1 4020
box 7 3 12 24
use welltap_svt  __well_tap__250
timestamp 1731220505
transform 1 0 3832 0 1 4020
box 7 3 12 24
use welltap_svt  __well_tap__249
timestamp 1731220505
transform 1 0 5656 0 -1 3952
box 7 3 12 24
use welltap_svt  __well_tap__248
timestamp 1731220505
transform 1 0 3832 0 -1 3952
box 7 3 12 24
use welltap_svt  __well_tap__247
timestamp 1731220505
transform 1 0 5656 0 1 3768
box 7 3 12 24
use welltap_svt  __well_tap__246
timestamp 1731220505
transform 1 0 3832 0 1 3768
box 7 3 12 24
use welltap_svt  __well_tap__245
timestamp 1731220505
transform 1 0 5656 0 -1 3692
box 7 3 12 24
use welltap_svt  __well_tap__244
timestamp 1731220505
transform 1 0 3832 0 -1 3692
box 7 3 12 24
use welltap_svt  __well_tap__243
timestamp 1731220505
transform 1 0 5656 0 1 3516
box 7 3 12 24
use welltap_svt  __well_tap__242
timestamp 1731220505
transform 1 0 3832 0 1 3516
box 7 3 12 24
use welltap_svt  __well_tap__241
timestamp 1731220505
transform 1 0 5656 0 -1 3460
box 7 3 12 24
use welltap_svt  __well_tap__240
timestamp 1731220505
transform 1 0 3832 0 -1 3460
box 7 3 12 24
use welltap_svt  __well_tap__239
timestamp 1731220505
transform 1 0 5656 0 1 3284
box 7 3 12 24
use welltap_svt  __well_tap__238
timestamp 1731220505
transform 1 0 3832 0 1 3284
box 7 3 12 24
use welltap_svt  __well_tap__237
timestamp 1731220505
transform 1 0 5656 0 -1 3212
box 7 3 12 24
use welltap_svt  __well_tap__236
timestamp 1731220505
transform 1 0 3832 0 -1 3212
box 7 3 12 24
use welltap_svt  __well_tap__235
timestamp 1731220505
transform 1 0 5656 0 1 3032
box 7 3 12 24
use welltap_svt  __well_tap__234
timestamp 1731220505
transform 1 0 3832 0 1 3032
box 7 3 12 24
use welltap_svt  __well_tap__233
timestamp 1731220505
transform 1 0 5656 0 -1 2960
box 7 3 12 24
use welltap_svt  __well_tap__232
timestamp 1731220505
transform 1 0 3832 0 -1 2960
box 7 3 12 24
use welltap_svt  __well_tap__231
timestamp 1731220505
transform 1 0 5656 0 1 2768
box 7 3 12 24
use welltap_svt  __well_tap__230
timestamp 1731220505
transform 1 0 3832 0 1 2768
box 7 3 12 24
use welltap_svt  __well_tap__229
timestamp 1731220505
transform 1 0 5656 0 -1 2708
box 7 3 12 24
use welltap_svt  __well_tap__228
timestamp 1731220505
transform 1 0 3832 0 -1 2708
box 7 3 12 24
use welltap_svt  __well_tap__227
timestamp 1731220505
transform 1 0 5656 0 1 2532
box 7 3 12 24
use welltap_svt  __well_tap__226
timestamp 1731220505
transform 1 0 3832 0 1 2532
box 7 3 12 24
use welltap_svt  __well_tap__225
timestamp 1731220505
transform 1 0 5656 0 -1 2480
box 7 3 12 24
use welltap_svt  __well_tap__224
timestamp 1731220505
transform 1 0 3832 0 -1 2480
box 7 3 12 24
use welltap_svt  __well_tap__223
timestamp 1731220505
transform 1 0 5656 0 1 2304
box 7 3 12 24
use welltap_svt  __well_tap__222
timestamp 1731220505
transform 1 0 3832 0 1 2304
box 7 3 12 24
use welltap_svt  __well_tap__221
timestamp 1731220505
transform 1 0 5656 0 -1 2232
box 7 3 12 24
use welltap_svt  __well_tap__220
timestamp 1731220505
transform 1 0 3832 0 -1 2232
box 7 3 12 24
use welltap_svt  __well_tap__219
timestamp 1731220505
transform 1 0 5656 0 1 2040
box 7 3 12 24
use welltap_svt  __well_tap__218
timestamp 1731220505
transform 1 0 3832 0 1 2040
box 7 3 12 24
use welltap_svt  __well_tap__217
timestamp 1731220505
transform 1 0 5656 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__216
timestamp 1731220505
transform 1 0 3832 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__215
timestamp 1731220505
transform 1 0 5656 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__214
timestamp 1731220505
transform 1 0 3832 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__213
timestamp 1731220505
transform 1 0 5656 0 -1 1760
box 7 3 12 24
use welltap_svt  __well_tap__212
timestamp 1731220505
transform 1 0 3832 0 -1 1760
box 7 3 12 24
use welltap_svt  __well_tap__211
timestamp 1731220505
transform 1 0 5656 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__210
timestamp 1731220505
transform 1 0 3832 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__209
timestamp 1731220505
transform 1 0 5656 0 -1 1528
box 7 3 12 24
use welltap_svt  __well_tap__208
timestamp 1731220505
transform 1 0 3832 0 -1 1528
box 7 3 12 24
use welltap_svt  __well_tap__207
timestamp 1731220505
transform 1 0 5656 0 1 1352
box 7 3 12 24
use welltap_svt  __well_tap__206
timestamp 1731220505
transform 1 0 3832 0 1 1352
box 7 3 12 24
use welltap_svt  __well_tap__205
timestamp 1731220505
transform 1 0 5656 0 -1 1304
box 7 3 12 24
use welltap_svt  __well_tap__204
timestamp 1731220505
transform 1 0 3832 0 -1 1304
box 7 3 12 24
use welltap_svt  __well_tap__203
timestamp 1731220505
transform 1 0 5656 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__202
timestamp 1731220505
transform 1 0 3832 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__201
timestamp 1731220505
transform 1 0 5656 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__200
timestamp 1731220505
transform 1 0 3832 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__199
timestamp 1731220505
transform 1 0 5656 0 1 868
box 7 3 12 24
use welltap_svt  __well_tap__198
timestamp 1731220505
transform 1 0 3832 0 1 868
box 7 3 12 24
use welltap_svt  __well_tap__197
timestamp 1731220505
transform 1 0 5656 0 -1 820
box 7 3 12 24
use welltap_svt  __well_tap__196
timestamp 1731220505
transform 1 0 3832 0 -1 820
box 7 3 12 24
use welltap_svt  __well_tap__195
timestamp 1731220505
transform 1 0 5656 0 1 644
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220505
transform 1 0 3832 0 1 644
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220505
transform 1 0 5656 0 -1 588
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220505
transform 1 0 3832 0 -1 588
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220505
transform 1 0 5656 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220505
transform 1 0 3832 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220505
transform 1 0 5656 0 -1 344
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220505
transform 1 0 3832 0 -1 344
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220505
transform 1 0 5656 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220505
transform 1 0 3832 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220505
transform 1 0 3792 0 -1 5696
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220505
transform 1 0 1968 0 -1 5696
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220505
transform 1 0 3792 0 1 5512
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220505
transform 1 0 1968 0 1 5512
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220505
transform 1 0 3792 0 -1 5464
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220505
transform 1 0 1968 0 -1 5464
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220505
transform 1 0 3792 0 1 5264
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220505
transform 1 0 1968 0 1 5264
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220505
transform 1 0 3792 0 -1 5216
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220505
transform 1 0 1968 0 -1 5216
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220505
transform 1 0 3792 0 1 5040
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220505
transform 1 0 1968 0 1 5040
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220505
transform 1 0 3792 0 -1 4960
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220505
transform 1 0 1968 0 -1 4960
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220505
transform 1 0 3792 0 1 4776
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220505
transform 1 0 1968 0 1 4776
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220505
transform 1 0 3792 0 -1 4724
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220505
transform 1 0 1968 0 -1 4724
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220505
transform 1 0 3792 0 1 4516
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220505
transform 1 0 1968 0 1 4516
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220505
transform 1 0 3792 0 -1 4460
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220505
transform 1 0 1968 0 -1 4460
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220505
transform 1 0 3792 0 1 4272
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220505
transform 1 0 1968 0 1 4272
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220505
transform 1 0 3792 0 -1 4196
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220505
transform 1 0 1968 0 -1 4196
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220505
transform 1 0 3792 0 1 4020
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220505
transform 1 0 1968 0 1 4020
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220505
transform 1 0 3792 0 -1 3964
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220505
transform 1 0 1968 0 -1 3964
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220505
transform 1 0 3792 0 1 3780
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220505
transform 1 0 1968 0 1 3780
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220505
transform 1 0 3792 0 -1 3728
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220505
transform 1 0 1968 0 -1 3728
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220505
transform 1 0 3792 0 1 3544
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220505
transform 1 0 1968 0 1 3544
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220505
transform 1 0 3792 0 -1 3456
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220505
transform 1 0 1968 0 -1 3456
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220505
transform 1 0 3792 0 1 3272
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220505
transform 1 0 1968 0 1 3272
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220505
transform 1 0 3792 0 -1 3224
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220505
transform 1 0 1968 0 -1 3224
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220505
transform 1 0 3792 0 1 3048
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220505
transform 1 0 1968 0 1 3048
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220505
transform 1 0 3792 0 -1 2992
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220505
transform 1 0 1968 0 -1 2992
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220505
transform 1 0 3792 0 1 2812
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220505
transform 1 0 1968 0 1 2812
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220505
transform 1 0 3792 0 -1 2760
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220505
transform 1 0 1968 0 -1 2760
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220505
transform 1 0 3792 0 1 2576
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220505
transform 1 0 1968 0 1 2576
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220505
transform 1 0 3792 0 -1 2528
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220505
transform 1 0 1968 0 -1 2528
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220505
transform 1 0 3792 0 1 2336
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220505
transform 1 0 1968 0 1 2336
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220505
transform 1 0 3792 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220505
transform 1 0 1968 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220505
transform 1 0 3792 0 1 2092
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220505
transform 1 0 1968 0 1 2092
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220505
transform 1 0 3792 0 -1 2036
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220505
transform 1 0 1968 0 -1 2036
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220505
transform 1 0 3792 0 1 1848
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220505
transform 1 0 1968 0 1 1848
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220505
transform 1 0 3792 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220505
transform 1 0 1968 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220505
transform 1 0 3792 0 1 1588
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220505
transform 1 0 1968 0 1 1588
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220505
transform 1 0 3792 0 -1 1536
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220505
transform 1 0 1968 0 -1 1536
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220505
transform 1 0 3792 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220505
transform 1 0 1968 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220505
transform 1 0 3792 0 -1 1292
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220505
transform 1 0 1968 0 -1 1292
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220505
transform 1 0 3792 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220505
transform 1 0 1968 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220505
transform 1 0 3792 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220505
transform 1 0 1968 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220505
transform 1 0 3792 0 1 872
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220505
transform 1 0 1968 0 1 872
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220505
transform 1 0 3792 0 -1 824
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220505
transform 1 0 1968 0 -1 824
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220505
transform 1 0 3792 0 1 632
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220505
transform 1 0 1968 0 1 632
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220505
transform 1 0 3792 0 -1 576
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220505
transform 1 0 1968 0 -1 576
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220505
transform 1 0 3792 0 1 380
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220505
transform 1 0 1968 0 1 380
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220505
transform 1 0 3792 0 -1 308
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220505
transform 1 0 1968 0 -1 308
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220505
transform 1 0 3792 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220505
transform 1 0 1968 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220505
transform 1 0 1928 0 1 5668
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220505
transform 1 0 104 0 1 5668
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220505
transform 1 0 1928 0 -1 5620
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220505
transform 1 0 104 0 -1 5620
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220505
transform 1 0 1928 0 1 5444
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220505
transform 1 0 104 0 1 5444
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220505
transform 1 0 1928 0 -1 5376
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220505
transform 1 0 104 0 -1 5376
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220505
transform 1 0 1928 0 1 5196
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220505
transform 1 0 104 0 1 5196
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220505
transform 1 0 1928 0 -1 5136
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220505
transform 1 0 104 0 -1 5136
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220505
transform 1 0 1928 0 1 4956
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220505
transform 1 0 104 0 1 4956
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220505
transform 1 0 1928 0 -1 4884
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220505
transform 1 0 104 0 -1 4884
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220505
transform 1 0 1928 0 1 4696
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220505
transform 1 0 104 0 1 4696
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220505
transform 1 0 1928 0 -1 4640
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220505
transform 1 0 104 0 -1 4640
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220505
transform 1 0 1928 0 1 4456
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220505
transform 1 0 104 0 1 4456
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220505
transform 1 0 1928 0 -1 4408
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220505
transform 1 0 104 0 -1 4408
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220505
transform 1 0 1928 0 1 4212
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220505
transform 1 0 104 0 1 4212
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220505
transform 1 0 1928 0 -1 4160
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220505
transform 1 0 104 0 -1 4160
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220505
transform 1 0 1928 0 1 3984
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220505
transform 1 0 104 0 1 3984
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220505
transform 1 0 1928 0 -1 3932
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220505
transform 1 0 104 0 -1 3932
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220505
transform 1 0 1928 0 1 3748
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220505
transform 1 0 104 0 1 3748
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220505
transform 1 0 1928 0 -1 3696
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220505
transform 1 0 104 0 -1 3696
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220505
transform 1 0 1928 0 1 3508
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220505
transform 1 0 104 0 1 3508
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220505
transform 1 0 1928 0 -1 3436
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220505
transform 1 0 104 0 -1 3436
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220505
transform 1 0 1928 0 1 3256
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220505
transform 1 0 104 0 1 3256
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220505
transform 1 0 1928 0 -1 3208
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220505
transform 1 0 104 0 -1 3208
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220505
transform 1 0 1928 0 1 3020
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220505
transform 1 0 104 0 1 3020
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220505
transform 1 0 1928 0 -1 2968
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220505
transform 1 0 104 0 -1 2968
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220505
transform 1 0 1928 0 1 2788
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220505
transform 1 0 104 0 1 2788
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220505
transform 1 0 1928 0 -1 2736
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220505
transform 1 0 104 0 -1 2736
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220505
transform 1 0 1928 0 1 2560
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220505
transform 1 0 104 0 1 2560
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220505
transform 1 0 1928 0 -1 2512
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220505
transform 1 0 104 0 -1 2512
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220505
transform 1 0 1928 0 1 2332
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220505
transform 1 0 104 0 1 2332
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220505
transform 1 0 1928 0 -1 2268
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220505
transform 1 0 104 0 -1 2268
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220505
transform 1 0 1928 0 1 2080
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220505
transform 1 0 104 0 1 2080
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220505
transform 1 0 1928 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220505
transform 1 0 104 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220505
transform 1 0 1928 0 1 1844
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220505
transform 1 0 104 0 1 1844
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220505
transform 1 0 1928 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220505
transform 1 0 104 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220505
transform 1 0 1928 0 1 1600
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220505
transform 1 0 104 0 1 1600
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220505
transform 1 0 1928 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220505
transform 1 0 104 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220505
transform 1 0 1928 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220505
transform 1 0 104 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220505
transform 1 0 1928 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220505
transform 1 0 104 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220505
transform 1 0 1928 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220505
transform 1 0 104 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220505
transform 1 0 1928 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220505
transform 1 0 104 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220505
transform 1 0 1928 0 1 868
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220505
transform 1 0 104 0 1 868
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220505
transform 1 0 1928 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220505
transform 1 0 104 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220505
transform 1 0 1928 0 1 612
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220505
transform 1 0 104 0 1 612
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220505
transform 1 0 1928 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220505
transform 1 0 104 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220505
transform 1 0 1928 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220505
transform 1 0 104 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220505
transform 1 0 1928 0 -1 328
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220505
transform 1 0 104 0 -1 328
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220505
transform 1 0 1928 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220505
transform 1 0 104 0 1 116
box 7 3 12 24
use _0_0std_0_0cells_0_0FAX1  tst_5999_6
timestamp 1731220505
transform 1 0 5296 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5998_6
timestamp 1731220505
transform 1 0 5512 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5997_6
timestamp 1731220505
transform 1 0 5512 0 -1 368
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5996_6
timestamp 1731220505
transform 1 0 5496 0 -1 612
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5995_6
timestamp 1731220505
transform 1 0 5456 0 1 620
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5994_6
timestamp 1731220505
transform 1 0 5512 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5993_6
timestamp 1731220505
transform 1 0 5328 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5992_6
timestamp 1731220505
transform 1 0 5120 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5991_6
timestamp 1731220505
transform 1 0 4904 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5990_6
timestamp 1731220505
transform 1 0 4680 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5989_6
timestamp 1731220505
transform 1 0 5280 0 -1 612
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5988_6
timestamp 1731220505
transform 1 0 5064 0 -1 612
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5987_6
timestamp 1731220505
transform 1 0 4848 0 -1 612
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5986_6
timestamp 1731220505
transform 1 0 4616 0 -1 612
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5985_6
timestamp 1731220505
transform 1 0 5224 0 1 620
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5984_6
timestamp 1731220505
transform 1 0 5000 0 1 620
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5983_6
timestamp 1731220505
transform 1 0 4776 0 1 620
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5982_6
timestamp 1731220505
transform 1 0 4768 0 -1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5981_6
timestamp 1731220505
transform 1 0 4544 0 -1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5980_6
timestamp 1731220505
transform 1 0 4312 0 -1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5979_6
timestamp 1731220505
transform 1 0 4808 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5978_6
timestamp 1731220505
transform 1 0 4592 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5977_6
timestamp 1731220505
transform 1 0 4376 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5976_6
timestamp 1731220505
transform 1 0 4360 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5975_6
timestamp 1731220505
transform 1 0 4656 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5974_6
timestamp 1731220505
transform 1 0 4432 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5973_6
timestamp 1731220505
transform 1 0 4960 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5972_6
timestamp 1731220505
transform 1 0 4688 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5971_6
timestamp 1731220505
transform 1 0 4640 0 -1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5970_6
timestamp 1731220505
transform 1 0 4360 0 -1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5969_6
timestamp 1731220505
transform 1 0 4088 0 -1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5968_6
timestamp 1731220505
transform 1 0 4008 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5967_6
timestamp 1731220505
transform 1 0 4208 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5966_6
timestamp 1731220505
transform 1 0 4064 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5965_6
timestamp 1731220505
transform 1 0 4152 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5964_6
timestamp 1731220505
transform 1 0 3928 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5963_6
timestamp 1731220505
transform 1 0 3856 0 -1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5962_6
timestamp 1731220505
transform 1 0 4080 0 -1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5961_6
timestamp 1731220505
transform 1 0 4080 0 1 620
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5960_6
timestamp 1731220505
transform 1 0 3856 0 1 620
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5959_6
timestamp 1731220505
transform 1 0 3856 0 -1 612
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5958_6
timestamp 1731220505
transform 1 0 4112 0 -1 612
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5957_6
timestamp 1731220505
transform 1 0 3888 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5956_6
timestamp 1731220505
transform 1 0 4168 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5955_6
timestamp 1731220505
transform 1 0 4168 0 -1 368
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5954_6
timestamp 1731220505
transform 1 0 3976 0 -1 368
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5953_6
timestamp 1731220505
transform 1 0 3992 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5952_6
timestamp 1731220505
transform 1 0 3856 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5951_6
timestamp 1731220505
transform 1 0 4128 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5950_6
timestamp 1731220505
transform 1 0 4264 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5949_6
timestamp 1731220505
transform 1 0 4432 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5948_6
timestamp 1731220505
transform 1 0 5064 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5947_6
timestamp 1731220505
transform 1 0 4840 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5946_6
timestamp 1731220505
transform 1 0 4624 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5945_6
timestamp 1731220505
transform 1 0 5232 0 -1 368
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5944_6
timestamp 1731220505
transform 1 0 4936 0 -1 368
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5943_6
timestamp 1731220505
transform 1 0 4648 0 -1 368
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5942_6
timestamp 1731220505
transform 1 0 4392 0 -1 368
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5941_6
timestamp 1731220505
transform 1 0 4432 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5940_6
timestamp 1731220505
transform 1 0 4376 0 -1 612
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5939_6
timestamp 1731220505
transform 1 0 4320 0 1 620
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5938_6
timestamp 1731220505
transform 1 0 4552 0 1 620
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5937_6
timestamp 1731220505
transform 1 0 5000 0 -1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5936_6
timestamp 1731220505
transform 1 0 5232 0 -1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5935_6
timestamp 1731220505
transform 1 0 5024 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5934_6
timestamp 1731220505
transform 1 0 5240 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5933_6
timestamp 1731220505
transform 1 0 5232 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5932_6
timestamp 1731220505
transform 1 0 4944 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5931_6
timestamp 1731220505
transform 1 0 5248 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5930_6
timestamp 1731220505
transform 1 0 5232 0 -1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5929_6
timestamp 1731220505
transform 1 0 4936 0 -1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5928_6
timestamp 1731220505
transform 1 0 5200 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5927_6
timestamp 1731220505
transform 1 0 4984 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5926_6
timestamp 1731220505
transform 1 0 4768 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5925_6
timestamp 1731220505
transform 1 0 4544 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5924_6
timestamp 1731220505
transform 1 0 4320 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5923_6
timestamp 1731220505
transform 1 0 5032 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5922_6
timestamp 1731220505
transform 1 0 4784 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5921_6
timestamp 1731220505
transform 1 0 4544 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5920_6
timestamp 1731220505
transform 1 0 4312 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5919_6
timestamp 1731220505
transform 1 0 5008 0 1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5918_6
timestamp 1731220505
transform 1 0 4760 0 1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5917_6
timestamp 1731220505
transform 1 0 4528 0 1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5916_6
timestamp 1731220505
transform 1 0 4320 0 1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5915_6
timestamp 1731220505
transform 1 0 4312 0 -1 1784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5914_6
timestamp 1731220505
transform 1 0 4056 0 -1 1784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5913_6
timestamp 1731220505
transform 1 0 4592 0 -1 1784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5912_6
timestamp 1731220505
transform 1 0 4896 0 -1 1784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5911_6
timestamp 1731220505
transform 1 0 4728 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5910_6
timestamp 1731220505
transform 1 0 4496 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5909_6
timestamp 1731220505
transform 1 0 4272 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5908_6
timestamp 1731220505
transform 1 0 4976 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5907_6
timestamp 1731220505
transform 1 0 4832 0 -1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5906_6
timestamp 1731220505
transform 1 0 4696 0 -1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5905_6
timestamp 1731220505
transform 1 0 5128 0 -1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5904_6
timestamp 1731220505
transform 1 0 4976 0 -1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5903_6
timestamp 1731220505
transform 1 0 4952 0 1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5902_6
timestamp 1731220505
transform 1 0 5088 0 1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5901_6
timestamp 1731220505
transform 1 0 5224 0 1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5900_6
timestamp 1731220505
transform 1 0 5288 0 -1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5899_6
timestamp 1731220505
transform 1 0 5232 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5898_6
timestamp 1731220505
transform 1 0 5216 0 -1 1784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5897_6
timestamp 1731220505
transform 1 0 5272 0 1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5896_6
timestamp 1731220505
transform 1 0 5280 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5895_6
timestamp 1731220505
transform 1 0 5416 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5894_6
timestamp 1731220505
transform 1 0 5464 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5893_6
timestamp 1731220505
transform 1 0 5464 0 -1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5892_6
timestamp 1731220505
transform 1 0 5512 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5891_6
timestamp 1731220505
transform 1 0 5512 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5890_6
timestamp 1731220505
transform 1 0 5512 0 -1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5889_6
timestamp 1731220505
transform 1 0 5512 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5888_6
timestamp 1731220505
transform 1 0 5512 0 1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5887_6
timestamp 1731220505
transform 1 0 5512 0 -1 1784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5886_6
timestamp 1731220505
transform 1 0 5496 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5885_6
timestamp 1731220505
transform 1 0 5456 0 -1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5884_6
timestamp 1731220505
transform 1 0 5512 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5883_6
timestamp 1731220505
transform 1 0 5512 0 1 2280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5882_6
timestamp 1731220505
transform 1 0 5512 0 1 2508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5881_6
timestamp 1731220505
transform 1 0 5512 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5880_6
timestamp 1731220505
transform 1 0 5512 0 1 2744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5879_6
timestamp 1731220505
transform 1 0 5512 0 -1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5878_6
timestamp 1731220505
transform 1 0 5320 0 -1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5877_6
timestamp 1731220505
transform 1 0 5104 0 -1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5876_6
timestamp 1731220505
transform 1 0 5248 0 1 2744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5875_6
timestamp 1731220505
transform 1 0 5264 0 1 2508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5874_6
timestamp 1731220505
transform 1 0 5320 0 -1 2504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5873_6
timestamp 1731220505
transform 1 0 5280 0 1 2280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5872_6
timestamp 1731220505
transform 1 0 5376 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5871_6
timestamp 1731220505
transform 1 0 5240 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5870_6
timestamp 1731220505
transform 1 0 5104 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5869_6
timestamp 1731220505
transform 1 0 4968 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5868_6
timestamp 1731220505
transform 1 0 4832 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5867_6
timestamp 1731220505
transform 1 0 4696 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5866_6
timestamp 1731220505
transform 1 0 4560 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5865_6
timestamp 1731220505
transform 1 0 5040 0 1 2280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5864_6
timestamp 1731220505
transform 1 0 4808 0 1 2280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5863_6
timestamp 1731220505
transform 1 0 4576 0 1 2280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5862_6
timestamp 1731220505
transform 1 0 4336 0 1 2280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5861_6
timestamp 1731220505
transform 1 0 5056 0 -1 2504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5860_6
timestamp 1731220505
transform 1 0 4792 0 -1 2504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5859_6
timestamp 1731220505
transform 1 0 4536 0 -1 2504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5858_6
timestamp 1731220505
transform 1 0 4288 0 -1 2504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5857_6
timestamp 1731220505
transform 1 0 4992 0 1 2508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5856_6
timestamp 1731220505
transform 1 0 4728 0 1 2508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5855_6
timestamp 1731220505
transform 1 0 4488 0 1 2508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5854_6
timestamp 1731220505
transform 1 0 4264 0 1 2508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5853_6
timestamp 1731220505
transform 1 0 5184 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5852_6
timestamp 1731220505
transform 1 0 4832 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5851_6
timestamp 1731220505
transform 1 0 4496 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5850_6
timestamp 1731220505
transform 1 0 4192 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5849_6
timestamp 1731220505
transform 1 0 4008 0 1 2744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5848_6
timestamp 1731220505
transform 1 0 4208 0 1 2744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5847_6
timestamp 1731220505
transform 1 0 4960 0 1 2744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5846_6
timestamp 1731220505
transform 1 0 4688 0 1 2744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5845_6
timestamp 1731220505
transform 1 0 4432 0 1 2744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5844_6
timestamp 1731220505
transform 1 0 4304 0 -1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5843_6
timestamp 1731220505
transform 1 0 4128 0 -1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5842_6
timestamp 1731220505
transform 1 0 4896 0 -1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5841_6
timestamp 1731220505
transform 1 0 4688 0 -1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5840_6
timestamp 1731220505
transform 1 0 4488 0 -1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5839_6
timestamp 1731220505
transform 1 0 4328 0 1 3008
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5838_6
timestamp 1731220505
transform 1 0 4128 0 1 3008
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5837_6
timestamp 1731220505
transform 1 0 4912 0 1 3008
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5836_6
timestamp 1731220505
transform 1 0 4712 0 1 3008
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5835_6
timestamp 1731220505
transform 1 0 4520 0 1 3008
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5834_6
timestamp 1731220505
transform 1 0 4408 0 -1 3236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5833_6
timestamp 1731220505
transform 1 0 4152 0 -1 3236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5832_6
timestamp 1731220505
transform 1 0 4656 0 -1 3236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5831_6
timestamp 1731220505
transform 1 0 5160 0 -1 3236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5830_6
timestamp 1731220505
transform 1 0 4904 0 -1 3236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5829_6
timestamp 1731220505
transform 1 0 4688 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5828_6
timestamp 1731220505
transform 1 0 4424 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5827_6
timestamp 1731220505
transform 1 0 4936 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5826_6
timestamp 1731220505
transform 1 0 5176 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5825_6
timestamp 1731220505
transform 1 0 5424 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5824_6
timestamp 1731220505
transform 1 0 5344 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5823_6
timestamp 1731220505
transform 1 0 5208 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5822_6
timestamp 1731220505
transform 1 0 5072 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5821_6
timestamp 1731220505
transform 1 0 4936 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5820_6
timestamp 1731220505
transform 1 0 4800 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5819_6
timestamp 1731220505
transform 1 0 5080 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5818_6
timestamp 1731220505
transform 1 0 4944 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5817_6
timestamp 1731220505
transform 1 0 4808 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5816_6
timestamp 1731220505
transform 1 0 4672 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5815_6
timestamp 1731220505
transform 1 0 4536 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5814_6
timestamp 1731220505
transform 1 0 4600 0 -1 3716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5813_6
timestamp 1731220505
transform 1 0 4408 0 -1 3716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5812_6
timestamp 1731220505
transform 1 0 4216 0 -1 3716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5811_6
timestamp 1731220505
transform 1 0 4024 0 -1 3716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5810_6
timestamp 1731220505
transform 1 0 4048 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5809_6
timestamp 1731220505
transform 1 0 4264 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5808_6
timestamp 1731220505
transform 1 0 4480 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5807_6
timestamp 1731220505
transform 1 0 4696 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5806_6
timestamp 1731220505
transform 1 0 4512 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5805_6
timestamp 1731220505
transform 1 0 4328 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5804_6
timestamp 1731220505
transform 1 0 4704 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5803_6
timestamp 1731220505
transform 1 0 4896 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5802_6
timestamp 1731220505
transform 1 0 4832 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5801_6
timestamp 1731220505
transform 1 0 4696 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5800_6
timestamp 1731220505
transform 1 0 4560 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5799_6
timestamp 1731220505
transform 1 0 4968 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5798_6
timestamp 1731220505
transform 1 0 5104 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5797_6
timestamp 1731220505
transform 1 0 5240 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5796_6
timestamp 1731220505
transform 1 0 5376 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5795_6
timestamp 1731220505
transform 1 0 5296 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5794_6
timestamp 1731220505
transform 1 0 5096 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5793_6
timestamp 1731220505
transform 1 0 4904 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5792_6
timestamp 1731220505
transform 1 0 5112 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5791_6
timestamp 1731220505
transform 1 0 5320 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5790_6
timestamp 1731220505
transform 1 0 5512 0 1 3744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5789_6
timestamp 1731220505
transform 1 0 5496 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5788_6
timestamp 1731220505
transform 1 0 5512 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5787_6
timestamp 1731220505
transform 1 0 5512 0 -1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5786_6
timestamp 1731220505
transform 1 0 5512 0 1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5785_6
timestamp 1731220505
transform 1 0 5512 0 -1 4508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5784_6
timestamp 1731220505
transform 1 0 5512 0 1 4520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5783_6
timestamp 1731220505
transform 1 0 5512 0 -1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5782_6
timestamp 1731220505
transform 1 0 5512 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5781_6
timestamp 1731220505
transform 1 0 5512 0 -1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5780_6
timestamp 1731220505
transform 1 0 5360 0 -1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5779_6
timestamp 1731220505
transform 1 0 5184 0 -1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5778_6
timestamp 1731220505
transform 1 0 5008 0 -1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5777_6
timestamp 1731220505
transform 1 0 5368 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5776_6
timestamp 1731220505
transform 1 0 5208 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5775_6
timestamp 1731220505
transform 1 0 5208 0 -1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5774_6
timestamp 1731220505
transform 1 0 5056 0 -1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5773_6
timestamp 1731220505
transform 1 0 5040 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5772_6
timestamp 1731220505
transform 1 0 4872 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5771_6
timestamp 1731220505
transform 1 0 4696 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5770_6
timestamp 1731220505
transform 1 0 4624 0 -1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5769_6
timestamp 1731220505
transform 1 0 4824 0 -1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5768_6
timestamp 1731220505
transform 1 0 4840 0 1 5032
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5767_6
timestamp 1731220505
transform 1 0 5096 0 1 5032
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5766_6
timestamp 1731220505
transform 1 0 5008 0 -1 5276
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5765_6
timestamp 1731220505
transform 1 0 4792 0 -1 5276
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5764_6
timestamp 1731220505
transform 1 0 4776 0 1 5280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5763_6
timestamp 1731220505
transform 1 0 4960 0 1 5280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5762_6
timestamp 1731220505
transform 1 0 4896 0 -1 5528
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5761_6
timestamp 1731220505
transform 1 0 4688 0 -1 5528
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5760_6
timestamp 1731220505
transform 1 0 5104 0 -1 5528
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5759_6
timestamp 1731220505
transform 1 0 5192 0 1 5560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5758_6
timestamp 1731220505
transform 1 0 5056 0 1 5560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5757_6
timestamp 1731220505
transform 1 0 4920 0 1 5560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5756_6
timestamp 1731220505
transform 1 0 4784 0 1 5560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5755_6
timestamp 1731220505
transform 1 0 4648 0 1 5560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5754_6
timestamp 1731220505
transform 1 0 4512 0 1 5560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5753_6
timestamp 1731220505
transform 1 0 4376 0 1 5560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5752_6
timestamp 1731220505
transform 1 0 4240 0 1 5560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5751_6
timestamp 1731220505
transform 1 0 4104 0 1 5560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5750_6
timestamp 1731220505
transform 1 0 4272 0 -1 5528
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5749_6
timestamp 1731220505
transform 1 0 4480 0 -1 5528
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5748_6
timestamp 1731220505
transform 1 0 4432 0 1 5280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5747_6
timestamp 1731220505
transform 1 0 4600 0 1 5280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5746_6
timestamp 1731220505
transform 1 0 4576 0 -1 5276
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5745_6
timestamp 1731220505
transform 1 0 4592 0 1 5032
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5744_6
timestamp 1731220505
transform 1 0 4416 0 -1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5743_6
timestamp 1731220505
transform 1 0 4296 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5742_6
timestamp 1731220505
transform 1 0 4504 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5741_6
timestamp 1731220505
transform 1 0 4912 0 -1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5740_6
timestamp 1731220505
transform 1 0 5368 0 -1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5739_6
timestamp 1731220505
transform 1 0 5336 0 1 4520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5738_6
timestamp 1731220505
transform 1 0 5144 0 1 4520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5737_6
timestamp 1731220505
transform 1 0 4952 0 1 4520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5736_6
timestamp 1731220505
transform 1 0 4768 0 1 4520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5735_6
timestamp 1731220505
transform 1 0 5296 0 -1 4508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5734_6
timestamp 1731220505
transform 1 0 5064 0 -1 4508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5733_6
timestamp 1731220505
transform 1 0 4848 0 -1 4508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5732_6
timestamp 1731220505
transform 1 0 4640 0 -1 4508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5731_6
timestamp 1731220505
transform 1 0 4456 0 -1 4508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5730_6
timestamp 1731220505
transform 1 0 5248 0 1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5729_6
timestamp 1731220505
transform 1 0 4976 0 1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5728_6
timestamp 1731220505
transform 1 0 4712 0 1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5727_6
timestamp 1731220505
transform 1 0 4480 0 1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5726_6
timestamp 1731220505
transform 1 0 4280 0 1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5725_6
timestamp 1731220505
transform 1 0 5240 0 -1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5724_6
timestamp 1731220505
transform 1 0 4968 0 -1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5723_6
timestamp 1731220505
transform 1 0 4704 0 -1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5722_6
timestamp 1731220505
transform 1 0 4472 0 -1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5721_6
timestamp 1731220505
transform 1 0 4272 0 -1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5720_6
timestamp 1731220505
transform 1 0 4128 0 -1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5719_6
timestamp 1731220505
transform 1 0 3992 0 -1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5718_6
timestamp 1731220505
transform 1 0 3856 0 -1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5717_6
timestamp 1731220505
transform 1 0 4128 0 1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5716_6
timestamp 1731220505
transform 1 0 3992 0 1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5715_6
timestamp 1731220505
transform 1 0 3856 0 1 4260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5714_6
timestamp 1731220505
transform 1 0 3648 0 1 4248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5713_6
timestamp 1731220505
transform 1 0 3648 0 -1 4484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5712_6
timestamp 1731220505
transform 1 0 3440 0 -1 4484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5711_6
timestamp 1731220505
transform 1 0 3216 0 -1 4484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5710_6
timestamp 1731220505
transform 1 0 2984 0 -1 4484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5709_6
timestamp 1731220505
transform 1 0 2752 0 -1 4484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5708_6
timestamp 1731220505
transform 1 0 2824 0 1 4492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5707_6
timestamp 1731220505
transform 1 0 3072 0 1 4492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5706_6
timestamp 1731220505
transform 1 0 3312 0 1 4492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5705_6
timestamp 1731220505
transform 1 0 3560 0 1 4492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5704_6
timestamp 1731220505
transform 1 0 3512 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5703_6
timestamp 1731220505
transform 1 0 3368 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5702_6
timestamp 1731220505
transform 1 0 3648 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5701_6
timestamp 1731220505
transform 1 0 3856 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5700_6
timestamp 1731220505
transform 1 0 4072 0 1 4768
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5699_6
timestamp 1731220505
transform 1 0 3952 0 -1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5698_6
timestamp 1731220505
transform 1 0 4192 0 -1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5697_6
timestamp 1731220505
transform 1 0 4096 0 1 5032
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5696_6
timestamp 1731220505
transform 1 0 4344 0 1 5032
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5695_6
timestamp 1731220505
transform 1 0 4368 0 -1 5276
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5694_6
timestamp 1731220505
transform 1 0 4168 0 -1 5276
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5693_6
timestamp 1731220505
transform 1 0 3968 0 -1 5276
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5692_6
timestamp 1731220505
transform 1 0 4272 0 1 5280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5691_6
timestamp 1731220505
transform 1 0 4128 0 1 5280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5690_6
timestamp 1731220505
transform 1 0 3992 0 1 5280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5689_6
timestamp 1731220505
transform 1 0 3856 0 1 5280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5688_6
timestamp 1731220505
transform 1 0 3648 0 1 5240
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5687_6
timestamp 1731220505
transform 1 0 3264 0 1 5240
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5686_6
timestamp 1731220505
transform 1 0 3632 0 -1 5240
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5685_6
timestamp 1731220505
transform 1 0 3272 0 -1 5240
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5684_6
timestamp 1731220505
transform 1 0 2912 0 -1 5240
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5683_6
timestamp 1731220505
transform 1 0 2992 0 1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5682_6
timestamp 1731220505
transform 1 0 3232 0 1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5681_6
timestamp 1731220505
transform 1 0 3472 0 1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5680_6
timestamp 1731220505
transform 1 0 3320 0 -1 4984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5679_6
timestamp 1731220505
transform 1 0 3168 0 -1 4984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5678_6
timestamp 1731220505
transform 1 0 3016 0 -1 4984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5677_6
timestamp 1731220505
transform 1 0 2872 0 1 4752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5676_6
timestamp 1731220505
transform 1 0 3024 0 1 4752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5675_6
timestamp 1731220505
transform 1 0 3176 0 1 4752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5674_6
timestamp 1731220505
transform 1 0 3216 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5673_6
timestamp 1731220505
transform 1 0 3080 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5672_6
timestamp 1731220505
transform 1 0 2944 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5671_6
timestamp 1731220505
transform 1 0 2808 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5670_6
timestamp 1731220505
transform 1 0 2672 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5669_6
timestamp 1731220505
transform 1 0 2536 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5668_6
timestamp 1731220505
transform 1 0 2400 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5667_6
timestamp 1731220505
transform 1 0 2264 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5666_6
timestamp 1731220505
transform 1 0 2128 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5665_6
timestamp 1731220505
transform 1 0 1992 0 -1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5664_6
timestamp 1731220505
transform 1 0 2320 0 1 4492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5663_6
timestamp 1731220505
transform 1 0 2576 0 1 4492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5662_6
timestamp 1731220505
transform 1 0 2512 0 -1 4484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5661_6
timestamp 1731220505
transform 1 0 2800 0 1 4248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5660_6
timestamp 1731220505
transform 1 0 3232 0 1 4248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5659_6
timestamp 1731220505
transform 1 0 2952 0 -1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5658_6
timestamp 1731220505
transform 1 0 2752 0 -1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5657_6
timestamp 1731220505
transform 1 0 2552 0 -1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5656_6
timestamp 1731220505
transform 1 0 2440 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5655_6
timestamp 1731220505
transform 1 0 2616 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5654_6
timestamp 1731220505
transform 1 0 2784 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5653_6
timestamp 1731220505
transform 1 0 2952 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5652_6
timestamp 1731220505
transform 1 0 3128 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5651_6
timestamp 1731220505
transform 1 0 2968 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5650_6
timestamp 1731220505
transform 1 0 2800 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5649_6
timestamp 1731220505
transform 1 0 2632 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5648_6
timestamp 1731220505
transform 1 0 3144 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5647_6
timestamp 1731220505
transform 1 0 3320 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5646_6
timestamp 1731220505
transform 1 0 3152 0 1 3756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5645_6
timestamp 1731220505
transform 1 0 2944 0 1 3756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5644_6
timestamp 1731220505
transform 1 0 2736 0 1 3756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5643_6
timestamp 1731220505
transform 1 0 3560 0 1 3756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5642_6
timestamp 1731220505
transform 1 0 3352 0 1 3756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5641_6
timestamp 1731220505
transform 1 0 3264 0 -1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5640_6
timestamp 1731220505
transform 1 0 3056 0 -1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5639_6
timestamp 1731220505
transform 1 0 2840 0 -1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5638_6
timestamp 1731220505
transform 1 0 3464 0 -1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5637_6
timestamp 1731220505
transform 1 0 3648 0 -1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5636_6
timestamp 1731220505
transform 1 0 3856 0 -1 3716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5635_6
timestamp 1731220505
transform 1 0 4400 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5634_6
timestamp 1731220505
transform 1 0 4264 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5633_6
timestamp 1731220505
transform 1 0 4128 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5632_6
timestamp 1731220505
transform 1 0 3992 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5631_6
timestamp 1731220505
transform 1 0 3856 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5630_6
timestamp 1731220505
transform 1 0 3648 0 -1 3480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5629_6
timestamp 1731220505
transform 1 0 3448 0 -1 3480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5628_6
timestamp 1731220505
transform 1 0 3232 0 -1 3480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5627_6
timestamp 1731220505
transform 1 0 3016 0 -1 3480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5626_6
timestamp 1731220505
transform 1 0 3856 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5625_6
timestamp 1731220505
transform 1 0 4136 0 1 3260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5624_6
timestamp 1731220505
transform 1 0 3880 0 -1 3236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5623_6
timestamp 1731220505
transform 1 0 3928 0 1 3008
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5622_6
timestamp 1731220505
transform 1 0 3968 0 -1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5621_6
timestamp 1731220505
transform 1 0 3856 0 1 2744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5620_6
timestamp 1731220505
transform 1 0 3936 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5619_6
timestamp 1731220505
transform 1 0 4064 0 1 2508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5618_6
timestamp 1731220505
transform 1 0 3888 0 1 2508
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5617_6
timestamp 1731220505
transform 1 0 3856 0 -1 2504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5616_6
timestamp 1731220505
transform 1 0 4056 0 -1 2504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5615_6
timestamp 1731220505
transform 1 0 4088 0 1 2280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5614_6
timestamp 1731220505
transform 1 0 3856 0 1 2280
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5613_6
timestamp 1731220505
transform 1 0 3648 0 -1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5612_6
timestamp 1731220505
transform 1 0 3512 0 -1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5611_6
timestamp 1731220505
transform 1 0 3432 0 1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5610_6
timestamp 1731220505
transform 1 0 3144 0 1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5609_6
timestamp 1731220505
transform 1 0 2856 0 1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5608_6
timestamp 1731220505
transform 1 0 2880 0 -1 2552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5607_6
timestamp 1731220505
transform 1 0 3192 0 -1 2552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5606_6
timestamp 1731220505
transform 1 0 3032 0 -1 2552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5605_6
timestamp 1731220505
transform 1 0 2968 0 1 2552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5604_6
timestamp 1731220505
transform 1 0 2832 0 1 2552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5603_6
timestamp 1731220505
transform 1 0 2912 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5602_6
timestamp 1731220505
transform 1 0 3072 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5601_6
timestamp 1731220505
transform 1 0 2992 0 1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5600_6
timestamp 1731220505
transform 1 0 3152 0 1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5599_6
timestamp 1731220505
transform 1 0 3312 0 1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5598_6
timestamp 1731220505
transform 1 0 3304 0 -1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5597_6
timestamp 1731220505
transform 1 0 3528 0 -1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5596_6
timestamp 1731220505
transform 1 0 3648 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5595_6
timestamp 1731220505
transform 1 0 3368 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5594_6
timestamp 1731220505
transform 1 0 3072 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5593_6
timestamp 1731220505
transform 1 0 3176 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5592_6
timestamp 1731220505
transform 1 0 3416 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5591_6
timestamp 1731220505
transform 1 0 3264 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5590_6
timestamp 1731220505
transform 1 0 3080 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5589_6
timestamp 1731220505
transform 1 0 2896 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5588_6
timestamp 1731220505
transform 1 0 2944 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5587_6
timestamp 1731220505
transform 1 0 2712 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5586_6
timestamp 1731220505
transform 1 0 2776 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5585_6
timestamp 1731220505
transform 1 0 3088 0 -1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5584_6
timestamp 1731220505
transform 1 0 2872 0 -1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5583_6
timestamp 1731220505
transform 1 0 2832 0 1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5582_6
timestamp 1731220505
transform 1 0 2680 0 1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5581_6
timestamp 1731220505
transform 1 0 2592 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5580_6
timestamp 1731220505
transform 1 0 2752 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5579_6
timestamp 1731220505
transform 1 0 2696 0 1 2552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5578_6
timestamp 1731220505
transform 1 0 2728 0 -1 2552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5577_6
timestamp 1731220505
transform 1 0 2576 0 -1 2552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5576_6
timestamp 1731220505
transform 1 0 2568 0 1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5575_6
timestamp 1731220505
transform 1 0 2272 0 1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5574_6
timestamp 1731220505
transform 1 0 2576 0 -1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5573_6
timestamp 1731220505
transform 1 0 2736 0 -1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5572_6
timestamp 1731220505
transform 1 0 2728 0 1 2068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5571_6
timestamp 1731220505
transform 1 0 2528 0 1 2068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5570_6
timestamp 1731220505
transform 1 0 2328 0 1 2068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5569_6
timestamp 1731220505
transform 1 0 2128 0 1 2068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5568_6
timestamp 1731220505
transform 1 0 2416 0 -1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5567_6
timestamp 1731220505
transform 1 0 2264 0 -1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5566_6
timestamp 1731220505
transform 1 0 2128 0 -1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5565_6
timestamp 1731220505
transform 1 0 1992 0 -1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5564_6
timestamp 1731220505
transform 1 0 1992 0 1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5563_6
timestamp 1731220505
transform 1 0 1784 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5562_6
timestamp 1731220505
transform 1 0 1528 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5561_6
timestamp 1731220505
transform 1 0 1744 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5560_6
timestamp 1731220505
transform 1 0 1576 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5559_6
timestamp 1731220505
transform 1 0 1408 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5558_6
timestamp 1731220505
transform 1 0 1240 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5557_6
timestamp 1731220505
transform 1 0 1200 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5556_6
timestamp 1731220505
transform 1 0 1368 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5555_6
timestamp 1731220505
transform 1 0 1712 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5554_6
timestamp 1731220505
transform 1 0 1536 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5553_6
timestamp 1731220505
transform 1 0 1536 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5552_6
timestamp 1731220505
transform 1 0 1784 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5551_6
timestamp 1731220505
transform 1 0 1992 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5550_6
timestamp 1731220505
transform 1 0 2432 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5549_6
timestamp 1731220505
transform 1 0 2272 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5548_6
timestamp 1731220505
transform 1 0 2128 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5547_6
timestamp 1731220505
transform 1 0 2128 0 1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5546_6
timestamp 1731220505
transform 1 0 1992 0 1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5545_6
timestamp 1731220505
transform 1 0 2536 0 1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5544_6
timestamp 1731220505
transform 1 0 2400 0 1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5543_6
timestamp 1731220505
transform 1 0 2264 0 1 2788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5542_6
timestamp 1731220505
transform 1 0 2160 0 -1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5541_6
timestamp 1731220505
transform 1 0 2320 0 -1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5540_6
timestamp 1731220505
transform 1 0 2672 0 -1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5539_6
timestamp 1731220505
transform 1 0 2488 0 -1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5538_6
timestamp 1731220505
transform 1 0 2480 0 1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5537_6
timestamp 1731220505
transform 1 0 2472 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5536_6
timestamp 1731220505
transform 1 0 2528 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5535_6
timestamp 1731220505
transform 1 0 2712 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5534_6
timestamp 1731220505
transform 1 0 2568 0 -1 3480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5533_6
timestamp 1731220505
transform 1 0 2792 0 -1 3480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5532_6
timestamp 1731220505
transform 1 0 2680 0 1 3520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5531_6
timestamp 1731220505
transform 1 0 2544 0 1 3520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5530_6
timestamp 1731220505
transform 1 0 2408 0 1 3520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5529_6
timestamp 1731220505
transform 1 0 2376 0 -1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5528_6
timestamp 1731220505
transform 1 0 2616 0 -1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5527_6
timestamp 1731220505
transform 1 0 2520 0 1 3756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5526_6
timestamp 1731220505
transform 1 0 2288 0 1 3756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5525_6
timestamp 1731220505
transform 1 0 2456 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5524_6
timestamp 1731220505
transform 1 0 2280 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5523_6
timestamp 1731220505
transform 1 0 2096 0 -1 3988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5522_6
timestamp 1731220505
transform 1 0 2072 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5521_6
timestamp 1731220505
transform 1 0 2256 0 1 3996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5520_6
timestamp 1731220505
transform 1 0 2160 0 -1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5519_6
timestamp 1731220505
transform 1 0 1992 0 -1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5518_6
timestamp 1731220505
transform 1 0 2352 0 -1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5517_6
timestamp 1731220505
transform 1 0 2376 0 1 4248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5516_6
timestamp 1731220505
transform 1 0 1992 0 1 4248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5515_6
timestamp 1731220505
transform 1 0 1784 0 -1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5514_6
timestamp 1731220505
transform 1 0 1640 0 -1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5513_6
timestamp 1731220505
transform 1 0 1784 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5512_6
timestamp 1731220505
transform 1 0 1616 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5511_6
timestamp 1731220505
transform 1 0 1424 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5510_6
timestamp 1731220505
transform 1 0 1240 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5509_6
timestamp 1731220505
transform 1 0 1312 0 -1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5508_6
timestamp 1731220505
transform 1 0 1472 0 -1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5507_6
timestamp 1731220505
transform 1 0 1416 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5506_6
timestamp 1731220505
transform 1 0 1592 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5505_6
timestamp 1731220505
transform 1 0 1752 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5504_6
timestamp 1731220505
transform 1 0 1520 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5503_6
timestamp 1731220505
transform 1 0 1488 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5502_6
timestamp 1731220505
transform 1 0 1784 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5501_6
timestamp 1731220505
transform 1 0 1784 0 -1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5500_6
timestamp 1731220505
transform 1 0 1544 0 -1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5499_6
timestamp 1731220505
transform 1 0 1280 0 -1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5498_6
timestamp 1731220505
transform 1 0 1512 0 1 3724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5497_6
timestamp 1731220505
transform 1 0 1784 0 1 3724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5496_6
timestamp 1731220505
transform 1 0 1728 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5495_6
timestamp 1731220505
transform 1 0 1560 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5494_6
timestamp 1731220505
transform 1 0 1392 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5493_6
timestamp 1731220505
transform 1 0 1728 0 1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5492_6
timestamp 1731220505
transform 1 0 1592 0 1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5491_6
timestamp 1731220505
transform 1 0 1456 0 1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5490_6
timestamp 1731220505
transform 1 0 1240 0 -1 3460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5489_6
timestamp 1731220505
transform 1 0 1104 0 -1 3460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5488_6
timestamp 1731220505
transform 1 0 968 0 -1 3460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5487_6
timestamp 1731220505
transform 1 0 832 0 -1 3460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5486_6
timestamp 1731220505
transform 1 0 696 0 -1 3460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5485_6
timestamp 1731220505
transform 1 0 752 0 1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5484_6
timestamp 1731220505
transform 1 0 1032 0 1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5483_6
timestamp 1731220505
transform 1 0 1192 0 -1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5482_6
timestamp 1731220505
transform 1 0 896 0 1 2996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5481_6
timestamp 1731220505
transform 1 0 704 0 1 2996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5480_6
timestamp 1731220505
transform 1 0 672 0 -1 2992
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5479_6
timestamp 1731220505
transform 1 0 632 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5478_6
timestamp 1731220505
transform 1 0 768 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5477_6
timestamp 1731220505
transform 1 0 768 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5476_6
timestamp 1731220505
transform 1 0 544 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5475_6
timestamp 1731220505
transform 1 0 344 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5474_6
timestamp 1731220505
transform 1 0 384 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5473_6
timestamp 1731220505
transform 1 0 536 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5472_6
timestamp 1731220505
transform 1 0 504 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5471_6
timestamp 1731220505
transform 1 0 296 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5470_6
timestamp 1731220505
transform 1 0 128 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5469_6
timestamp 1731220505
transform 1 0 688 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5468_6
timestamp 1731220505
transform 1 0 400 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5467_6
timestamp 1731220505
transform 1 0 392 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5466_6
timestamp 1731220505
transform 1 0 128 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5465_6
timestamp 1731220505
transform 1 0 128 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5464_6
timestamp 1731220505
transform 1 0 400 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5463_6
timestamp 1731220505
transform 1 0 728 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5462_6
timestamp 1731220505
transform 1 0 528 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5461_6
timestamp 1731220505
transform 1 0 352 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5460_6
timestamp 1731220505
transform 1 0 192 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5459_6
timestamp 1731220505
transform 1 0 192 0 1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5458_6
timestamp 1731220505
transform 1 0 384 0 1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5457_6
timestamp 1731220505
transform 1 0 448 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5456_6
timestamp 1731220505
transform 1 0 272 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5455_6
timestamp 1731220505
transform 1 0 128 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5454_6
timestamp 1731220505
transform 1 0 128 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5453_6
timestamp 1731220505
transform 1 0 328 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5452_6
timestamp 1731220505
transform 1 0 128 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5451_6
timestamp 1731220505
transform 1 0 128 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5450_6
timestamp 1731220505
transform 1 0 128 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5449_6
timestamp 1731220505
transform 1 0 144 0 -1 1076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5448_6
timestamp 1731220505
transform 1 0 192 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5447_6
timestamp 1731220505
transform 1 0 416 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5446_6
timestamp 1731220505
transform 1 0 192 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5445_6
timestamp 1731220505
transform 1 0 440 0 1 588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5444_6
timestamp 1731220505
transform 1 0 272 0 1 588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5443_6
timestamp 1731220505
transform 1 0 128 0 1 588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5442_6
timestamp 1731220505
transform 1 0 128 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5441_6
timestamp 1731220505
transform 1 0 344 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5440_6
timestamp 1731220505
transform 1 0 192 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5439_6
timestamp 1731220505
transform 1 0 472 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5438_6
timestamp 1731220505
transform 1 0 472 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5437_6
timestamp 1731220505
transform 1 0 280 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5436_6
timestamp 1731220505
transform 1 0 264 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5435_6
timestamp 1731220505
transform 1 0 128 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5434_6
timestamp 1731220505
transform 1 0 400 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5433_6
timestamp 1731220505
transform 1 0 536 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5432_6
timestamp 1731220505
transform 1 0 672 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5431_6
timestamp 1731220505
transform 1 0 1080 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5430_6
timestamp 1731220505
transform 1 0 944 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5429_6
timestamp 1731220505
transform 1 0 808 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5428_6
timestamp 1731220505
transform 1 0 664 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5427_6
timestamp 1731220505
transform 1 0 1048 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5426_6
timestamp 1731220505
transform 1 0 856 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5425_6
timestamp 1731220505
transform 1 0 752 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5424_6
timestamp 1731220505
transform 1 0 1328 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5423_6
timestamp 1731220505
transform 1 0 1040 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5422_6
timestamp 1731220505
transform 1 0 968 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5421_6
timestamp 1731220505
transform 1 0 776 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5420_6
timestamp 1731220505
transform 1 0 568 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5419_6
timestamp 1731220505
transform 1 0 608 0 1 588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5418_6
timestamp 1731220505
transform 1 0 768 0 1 588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5417_6
timestamp 1731220505
transform 1 0 920 0 1 588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5416_6
timestamp 1731220505
transform 1 0 848 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5415_6
timestamp 1731220505
transform 1 0 632 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5414_6
timestamp 1731220505
transform 1 0 416 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5413_6
timestamp 1731220505
transform 1 0 928 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5412_6
timestamp 1731220505
transform 1 0 664 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5411_6
timestamp 1731220505
transform 1 0 608 0 -1 1076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5410_6
timestamp 1731220505
transform 1 0 384 0 -1 1076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5409_6
timestamp 1731220505
transform 1 0 272 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5408_6
timestamp 1731220505
transform 1 0 600 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5407_6
timestamp 1731220505
transform 1 0 440 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5406_6
timestamp 1731220505
transform 1 0 336 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5405_6
timestamp 1731220505
transform 1 0 576 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5404_6
timestamp 1731220505
transform 1 0 552 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5403_6
timestamp 1731220505
transform 1 0 1000 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5402_6
timestamp 1731220505
transform 1 0 840 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5401_6
timestamp 1731220505
transform 1 0 1320 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5400_6
timestamp 1731220505
transform 1 0 1080 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5399_6
timestamp 1731220505
transform 1 0 1008 0 1 1576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5398_6
timestamp 1731220505
transform 1 0 1144 0 1 1576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5397_6
timestamp 1731220505
transform 1 0 1552 0 1 1576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5396_6
timestamp 1731220505
transform 1 0 1416 0 1 1576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5395_6
timestamp 1731220505
transform 1 0 1280 0 1 1576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5394_6
timestamp 1731220505
transform 1 0 1152 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5393_6
timestamp 1731220505
transform 1 0 1680 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5392_6
timestamp 1731220505
transform 1 0 1504 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5391_6
timestamp 1731220505
transform 1 0 1328 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5390_6
timestamp 1731220505
transform 1 0 1280 0 1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5389_6
timestamp 1731220505
transform 1 0 1768 0 1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5388_6
timestamp 1731220505
transform 1 0 1520 0 1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5387_6
timestamp 1731220505
transform 1 0 1352 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5386_6
timestamp 1731220505
transform 1 0 1576 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5385_6
timestamp 1731220505
transform 1 0 1784 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5384_6
timestamp 1731220505
transform 1 0 1784 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5383_6
timestamp 1731220505
transform 1 0 1992 0 -1 2060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5382_6
timestamp 1731220505
transform 1 0 2248 0 -1 2060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5381_6
timestamp 1731220505
transform 1 0 2520 0 -1 2060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5380_6
timestamp 1731220505
transform 1 0 2312 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5379_6
timestamp 1731220505
transform 1 0 1992 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5378_6
timestamp 1731220505
transform 1 0 2080 0 -1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5377_6
timestamp 1731220505
transform 1 0 2360 0 -1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5376_6
timestamp 1731220505
transform 1 0 2488 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5375_6
timestamp 1731220505
transform 1 0 2352 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5374_6
timestamp 1731220505
transform 1 0 2216 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5373_6
timestamp 1731220505
transform 1 0 2080 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5372_6
timestamp 1731220505
transform 1 0 2112 0 -1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5371_6
timestamp 1731220505
transform 1 0 2248 0 -1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5370_6
timestamp 1731220505
transform 1 0 2792 0 -1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5369_6
timestamp 1731220505
transform 1 0 2656 0 -1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5368_6
timestamp 1731220505
transform 1 0 2520 0 -1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5367_6
timestamp 1731220505
transform 1 0 2384 0 -1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5366_6
timestamp 1731220505
transform 1 0 2688 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5365_6
timestamp 1731220505
transform 1 0 2536 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5364_6
timestamp 1731220505
transform 1 0 2384 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5363_6
timestamp 1731220505
transform 1 0 2240 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5362_6
timestamp 1731220505
transform 1 0 2096 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5361_6
timestamp 1731220505
transform 1 0 2760 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5360_6
timestamp 1731220505
transform 1 0 2544 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5359_6
timestamp 1731220505
transform 1 0 2336 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5358_6
timestamp 1731220505
transform 1 0 2144 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5357_6
timestamp 1731220505
transform 1 0 1992 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5356_6
timestamp 1731220505
transform 1 0 1784 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5355_6
timestamp 1731220505
transform 1 0 1648 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5354_6
timestamp 1731220505
transform 1 0 1504 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5353_6
timestamp 1731220505
transform 1 0 1360 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5352_6
timestamp 1731220505
transform 1 0 1216 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5351_6
timestamp 1731220505
transform 1 0 1072 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5350_6
timestamp 1731220505
transform 1 0 1208 0 -1 1076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5349_6
timestamp 1731220505
transform 1 0 1392 0 -1 1076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5348_6
timestamp 1731220505
transform 1 0 1576 0 -1 1076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5347_6
timestamp 1731220505
transform 1 0 1760 0 -1 1076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5346_6
timestamp 1731220505
transform 1 0 1784 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5345_6
timestamp 1731220505
transform 1 0 1992 0 1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5344_6
timestamp 1731220505
transform 1 0 2216 0 1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5343_6
timestamp 1731220505
transform 1 0 2192 0 -1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5342_6
timestamp 1731220505
transform 1 0 2408 0 -1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5341_6
timestamp 1731220505
transform 1 0 2632 0 -1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5340_6
timestamp 1731220505
transform 1 0 2856 0 -1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5339_6
timestamp 1731220505
transform 1 0 2704 0 1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5338_6
timestamp 1731220505
transform 1 0 2464 0 1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5337_6
timestamp 1731220505
transform 1 0 2528 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5336_6
timestamp 1731220505
transform 1 0 2720 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5335_6
timestamp 1731220505
transform 1 0 3120 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5334_6
timestamp 1731220505
transform 1 0 2920 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5333_6
timestamp 1731220505
transform 1 0 2896 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5332_6
timestamp 1731220505
transform 1 0 2720 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5331_6
timestamp 1731220505
transform 1 0 3080 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5330_6
timestamp 1731220505
transform 1 0 3272 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5329_6
timestamp 1731220505
transform 1 0 3208 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5328_6
timestamp 1731220505
transform 1 0 2984 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5327_6
timestamp 1731220505
transform 1 0 2848 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5326_6
timestamp 1731220505
transform 1 0 3008 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5325_6
timestamp 1731220505
transform 1 0 3168 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5324_6
timestamp 1731220505
transform 1 0 3200 0 -1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5323_6
timestamp 1731220505
transform 1 0 3064 0 -1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5322_6
timestamp 1731220505
transform 1 0 2928 0 -1 1560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5321_6
timestamp 1731220505
transform 1 0 2912 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5320_6
timestamp 1731220505
transform 1 0 2768 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5319_6
timestamp 1731220505
transform 1 0 2624 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5318_6
timestamp 1731220505
transform 1 0 2632 0 -1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5317_6
timestamp 1731220505
transform 1 0 2896 0 -1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5316_6
timestamp 1731220505
transform 1 0 3152 0 -1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5315_6
timestamp 1731220505
transform 1 0 3160 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5314_6
timestamp 1731220505
transform 1 0 2896 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5313_6
timestamp 1731220505
transform 1 0 2616 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5312_6
timestamp 1731220505
transform 1 0 2768 0 -1 2060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5311_6
timestamp 1731220505
transform 1 0 3000 0 -1 2060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5310_6
timestamp 1731220505
transform 1 0 3224 0 -1 2060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5309_6
timestamp 1731220505
transform 1 0 3112 0 1 2068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5308_6
timestamp 1731220505
transform 1 0 2920 0 1 2068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5307_6
timestamp 1731220505
transform 1 0 2896 0 -1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5306_6
timestamp 1731220505
transform 1 0 3048 0 -1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5305_6
timestamp 1731220505
transform 1 0 3200 0 -1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5304_6
timestamp 1731220505
transform 1 0 3352 0 -1 2300
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5303_6
timestamp 1731220505
transform 1 0 3296 0 1 2068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5302_6
timestamp 1731220505
transform 1 0 3648 0 1 2068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5301_6
timestamp 1731220505
transform 1 0 3480 0 1 2068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5300_6
timestamp 1731220505
transform 1 0 3448 0 -1 2060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5299_6
timestamp 1731220505
transform 1 0 3648 0 -1 2060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5298_6
timestamp 1731220505
transform 1 0 3648 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5297_6
timestamp 1731220505
transform 1 0 3416 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5296_6
timestamp 1731220505
transform 1 0 3408 0 -1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5295_6
timestamp 1731220505
transform 1 0 3648 0 -1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5294_6
timestamp 1731220505
transform 1 0 3856 0 -1 1784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5293_6
timestamp 1731220505
transform 1 0 3856 0 1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5292_6
timestamp 1731220505
transform 1 0 4136 0 1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5291_6
timestamp 1731220505
transform 1 0 3992 0 1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5290_6
timestamp 1731220505
transform 1 0 3856 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5289_6
timestamp 1731220505
transform 1 0 4080 0 -1 1552
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5288_6
timestamp 1731220505
transform 1 0 4080 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5287_6
timestamp 1731220505
transform 1 0 3856 0 1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5286_6
timestamp 1731220505
transform 1 0 3856 0 -1 1328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5285_6
timestamp 1731220505
transform 1 0 3648 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5284_6
timestamp 1731220505
transform 1 0 3440 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5283_6
timestamp 1731220505
transform 1 0 3464 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5282_6
timestamp 1731220505
transform 1 0 3648 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5281_6
timestamp 1731220505
transform 1 0 3544 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5280_6
timestamp 1731220505
transform 1 0 3328 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5279_6
timestamp 1731220505
transform 1 0 3408 0 1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5278_6
timestamp 1731220505
transform 1 0 3168 0 1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5277_6
timestamp 1731220505
transform 1 0 2936 0 1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5276_6
timestamp 1731220505
transform 1 0 3080 0 -1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5275_6
timestamp 1731220505
transform 1 0 3304 0 -1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5274_6
timestamp 1731220505
transform 1 0 3528 0 -1 848
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5273_6
timestamp 1731220505
transform 1 0 3376 0 1 608
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5272_6
timestamp 1731220505
transform 1 0 3512 0 1 608
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5271_6
timestamp 1731220505
transform 1 0 3648 0 1 608
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5270_6
timestamp 1731220505
transform 1 0 3648 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5269_6
timestamp 1731220505
transform 1 0 3512 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5268_6
timestamp 1731220505
transform 1 0 3376 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5267_6
timestamp 1731220505
transform 1 0 3240 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5266_6
timestamp 1731220505
transform 1 0 3528 0 1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5265_6
timestamp 1731220505
transform 1 0 3328 0 1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5264_6
timestamp 1731220505
transform 1 0 3128 0 1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5263_6
timestamp 1731220505
transform 1 0 2928 0 1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5262_6
timestamp 1731220505
transform 1 0 3488 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5261_6
timestamp 1731220505
transform 1 0 3352 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5260_6
timestamp 1731220505
transform 1 0 3216 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5259_6
timestamp 1731220505
transform 1 0 3080 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5258_6
timestamp 1731220505
transform 1 0 2944 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5257_6
timestamp 1731220505
transform 1 0 2808 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5256_6
timestamp 1731220505
transform 1 0 3624 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5255_6
timestamp 1731220505
transform 1 0 3488 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5254_6
timestamp 1731220505
transform 1 0 3352 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5253_6
timestamp 1731220505
transform 1 0 3216 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5252_6
timestamp 1731220505
transform 1 0 3080 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5251_6
timestamp 1731220505
transform 1 0 2944 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5250_6
timestamp 1731220505
transform 1 0 2808 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5249_6
timestamp 1731220505
transform 1 0 2672 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5248_6
timestamp 1731220505
transform 1 0 2536 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5247_6
timestamp 1731220505
transform 1 0 2400 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5246_6
timestamp 1731220505
transform 1 0 2264 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5245_6
timestamp 1731220505
transform 1 0 2128 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5244_6
timestamp 1731220505
transform 1 0 1992 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5243_6
timestamp 1731220505
transform 1 0 2672 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5242_6
timestamp 1731220505
transform 1 0 2536 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5241_6
timestamp 1731220505
transform 1 0 2400 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5240_6
timestamp 1731220505
transform 1 0 2264 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5239_6
timestamp 1731220505
transform 1 0 2128 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5238_6
timestamp 1731220505
transform 1 0 1992 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5237_6
timestamp 1731220505
transform 1 0 2736 0 1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5236_6
timestamp 1731220505
transform 1 0 2536 0 1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5235_6
timestamp 1731220505
transform 1 0 2344 0 1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5234_6
timestamp 1731220505
transform 1 0 2152 0 1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5233_6
timestamp 1731220505
transform 1 0 1992 0 1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5232_6
timestamp 1731220505
transform 1 0 1784 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5231_6
timestamp 1731220505
transform 1 0 1640 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5230_6
timestamp 1731220505
transform 1 0 1480 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5229_6
timestamp 1731220505
transform 1 0 1312 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5228_6
timestamp 1731220505
transform 1 0 1144 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5227_6
timestamp 1731220505
transform 1 0 1784 0 1 588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5226_6
timestamp 1731220505
transform 1 0 1648 0 1 588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5225_6
timestamp 1731220505
transform 1 0 1504 0 1 588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5224_6
timestamp 1731220505
transform 1 0 1360 0 1 588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5223_6
timestamp 1731220505
transform 1 0 1216 0 1 588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5222_6
timestamp 1731220505
transform 1 0 1072 0 1 588
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5221_6
timestamp 1731220505
transform 1 0 1056 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5220_6
timestamp 1731220505
transform 1 0 1264 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5219_6
timestamp 1731220505
transform 1 0 1480 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5218_6
timestamp 1731220505
transform 1 0 1512 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5217_6
timestamp 1731220505
transform 1 0 1216 0 1 844
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5216_6
timestamp 1731220505
transform 1 0 1024 0 -1 1076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5215_6
timestamp 1731220505
transform 1 0 824 0 -1 1076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5214_6
timestamp 1731220505
transform 1 0 760 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5213_6
timestamp 1731220505
transform 1 0 920 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5212_6
timestamp 1731220505
transform 1 0 1056 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5211_6
timestamp 1731220505
transform 1 0 816 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5210_6
timestamp 1731220505
transform 1 0 776 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5209_6
timestamp 1731220505
transform 1 0 600 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5208_6
timestamp 1731220505
transform 1 0 360 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5207_6
timestamp 1731220505
transform 1 0 872 0 1 1576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5206_6
timestamp 1731220505
transform 1 0 800 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5205_6
timestamp 1731220505
transform 1 0 624 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5204_6
timestamp 1731220505
transform 1 0 976 0 -1 1804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5203_6
timestamp 1731220505
transform 1 0 1048 0 1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5202_6
timestamp 1731220505
transform 1 0 816 0 1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5201_6
timestamp 1731220505
transform 1 0 592 0 1 1820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5200_6
timestamp 1731220505
transform 1 0 720 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5199_6
timestamp 1731220505
transform 1 0 928 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5198_6
timestamp 1731220505
transform 1 0 1136 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5197_6
timestamp 1731220505
transform 1 0 1440 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5196_6
timestamp 1731220505
transform 1 0 1080 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5195_6
timestamp 1731220505
transform 1 0 968 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5194_6
timestamp 1731220505
transform 1 0 680 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5193_6
timestamp 1731220505
transform 1 0 1264 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5192_6
timestamp 1731220505
transform 1 0 1248 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5191_6
timestamp 1731220505
transform 1 0 968 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5190_6
timestamp 1731220505
transform 1 0 1064 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5189_6
timestamp 1731220505
transform 1 0 888 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5188_6
timestamp 1731220505
transform 1 0 704 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5187_6
timestamp 1731220505
transform 1 0 696 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5186_6
timestamp 1731220505
transform 1 0 864 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5185_6
timestamp 1731220505
transform 1 0 1032 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5184_6
timestamp 1731220505
transform 1 0 1264 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5183_6
timestamp 1731220505
transform 1 0 1008 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5182_6
timestamp 1731220505
transform 1 0 496 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5181_6
timestamp 1731220505
transform 1 0 360 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5180_6
timestamp 1731220505
transform 1 0 224 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5179_6
timestamp 1731220505
transform 1 0 536 0 -1 2992
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5178_6
timestamp 1731220505
transform 1 0 400 0 -1 2992
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5177_6
timestamp 1731220505
transform 1 0 264 0 -1 2992
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5176_6
timestamp 1731220505
transform 1 0 128 0 -1 2992
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5175_6
timestamp 1731220505
transform 1 0 128 0 1 2996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5174_6
timestamp 1731220505
transform 1 0 304 0 1 2996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5173_6
timestamp 1731220505
transform 1 0 504 0 1 2996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5172_6
timestamp 1731220505
transform 1 0 360 0 -1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5171_6
timestamp 1731220505
transform 1 0 616 0 -1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5170_6
timestamp 1731220505
transform 1 0 896 0 -1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5169_6
timestamp 1731220505
transform 1 0 888 0 1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5168_6
timestamp 1731220505
transform 1 0 1184 0 1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5167_6
timestamp 1731220505
transform 1 0 1336 0 1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5166_6
timestamp 1731220505
transform 1 0 1496 0 -1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5165_6
timestamp 1731220505
transform 1 0 1448 0 1 2996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5164_6
timestamp 1731220505
transform 1 0 1272 0 1 2996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5163_6
timestamp 1731220505
transform 1 0 1088 0 1 2996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5162_6
timestamp 1731220505
transform 1 0 1624 0 1 2996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5161_6
timestamp 1731220505
transform 1 0 1784 0 1 2996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5160_6
timestamp 1731220505
transform 1 0 2224 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5159_6
timestamp 1731220505
transform 1 0 1992 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5158_6
timestamp 1731220505
transform 1 0 1784 0 -1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5157_6
timestamp 1731220505
transform 1 0 1784 0 1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5156_6
timestamp 1731220505
transform 1 0 1648 0 1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5155_6
timestamp 1731220505
transform 1 0 1488 0 1 3232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5154_6
timestamp 1731220505
transform 1 0 1784 0 -1 3460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5153_6
timestamp 1731220505
transform 1 0 1648 0 -1 3460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5152_6
timestamp 1731220505
transform 1 0 1512 0 -1 3460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5151_6
timestamp 1731220505
transform 1 0 1376 0 -1 3460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5150_6
timestamp 1731220505
transform 1 0 1320 0 1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5149_6
timestamp 1731220505
transform 1 0 1184 0 1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5148_6
timestamp 1731220505
transform 1 0 1048 0 1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5147_6
timestamp 1731220505
transform 1 0 912 0 1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5146_6
timestamp 1731220505
transform 1 0 776 0 1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5145_6
timestamp 1731220505
transform 1 0 1224 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5144_6
timestamp 1731220505
transform 1 0 1056 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5143_6
timestamp 1731220505
transform 1 0 896 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5142_6
timestamp 1731220505
transform 1 0 744 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5141_6
timestamp 1731220505
transform 1 0 600 0 -1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5140_6
timestamp 1731220505
transform 1 0 1232 0 1 3724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5139_6
timestamp 1731220505
transform 1 0 960 0 1 3724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5138_6
timestamp 1731220505
transform 1 0 704 0 1 3724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5137_6
timestamp 1731220505
transform 1 0 472 0 1 3724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5136_6
timestamp 1731220505
transform 1 0 264 0 1 3724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5135_6
timestamp 1731220505
transform 1 0 1024 0 -1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5134_6
timestamp 1731220505
transform 1 0 776 0 -1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5133_6
timestamp 1731220505
transform 1 0 536 0 -1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5132_6
timestamp 1731220505
transform 1 0 312 0 -1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5131_6
timestamp 1731220505
transform 1 0 128 0 -1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5130_6
timestamp 1731220505
transform 1 0 128 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5129_6
timestamp 1731220505
transform 1 0 336 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5128_6
timestamp 1731220505
transform 1 0 592 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5127_6
timestamp 1731220505
transform 1 0 1176 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5126_6
timestamp 1731220505
transform 1 0 872 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5125_6
timestamp 1731220505
transform 1 0 672 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5124_6
timestamp 1731220505
transform 1 0 488 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5123_6
timestamp 1731220505
transform 1 0 1296 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5122_6
timestamp 1731220505
transform 1 0 1072 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5121_6
timestamp 1731220505
transform 1 0 864 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5120_6
timestamp 1731220505
transform 1 0 768 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5119_6
timestamp 1731220505
transform 1 0 624 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5118_6
timestamp 1731220505
transform 1 0 920 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5117_6
timestamp 1731220505
transform 1 0 1080 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5116_6
timestamp 1731220505
transform 1 0 1248 0 1 4188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5115_6
timestamp 1731220505
transform 1 0 1152 0 -1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5114_6
timestamp 1731220505
transform 1 0 992 0 -1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5113_6
timestamp 1731220505
transform 1 0 832 0 -1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5112_6
timestamp 1731220505
transform 1 0 680 0 -1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5111_6
timestamp 1731220505
transform 1 0 536 0 -1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5110_6
timestamp 1731220505
transform 1 0 1056 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5109_6
timestamp 1731220505
transform 1 0 872 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5108_6
timestamp 1731220505
transform 1 0 688 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5107_6
timestamp 1731220505
transform 1 0 512 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5106_6
timestamp 1731220505
transform 1 0 336 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5105_6
timestamp 1731220505
transform 1 0 672 0 -1 4664
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5104_6
timestamp 1731220505
transform 1 0 536 0 -1 4664
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5103_6
timestamp 1731220505
transform 1 0 400 0 -1 4664
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5102_6
timestamp 1731220505
transform 1 0 264 0 -1 4664
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5101_6
timestamp 1731220505
transform 1 0 128 0 -1 4664
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5100_6
timestamp 1731220505
transform 1 0 672 0 1 4672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_599_6
timestamp 1731220505
transform 1 0 536 0 1 4672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_598_6
timestamp 1731220505
transform 1 0 400 0 1 4672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_597_6
timestamp 1731220505
transform 1 0 264 0 1 4672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_596_6
timestamp 1731220505
transform 1 0 128 0 1 4672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_595_6
timestamp 1731220505
transform 1 0 128 0 -1 4908
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_594_6
timestamp 1731220505
transform 1 0 264 0 -1 4908
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_593_6
timestamp 1731220505
transform 1 0 672 0 -1 4908
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_592_6
timestamp 1731220505
transform 1 0 536 0 -1 4908
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_591_6
timestamp 1731220505
transform 1 0 400 0 -1 4908
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_590_6
timestamp 1731220505
transform 1 0 320 0 1 4932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_589_6
timestamp 1731220505
transform 1 0 128 0 1 4932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_588_6
timestamp 1731220505
transform 1 0 1080 0 1 4932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_587_6
timestamp 1731220505
transform 1 0 808 0 1 4932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_586_6
timestamp 1731220505
transform 1 0 552 0 1 4932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_585_6
timestamp 1731220505
transform 1 0 504 0 -1 5160
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_584_6
timestamp 1731220505
transform 1 0 336 0 -1 5160
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_583_6
timestamp 1731220505
transform 1 0 1048 0 -1 5160
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_582_6
timestamp 1731220505
transform 1 0 864 0 -1 5160
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_581_6
timestamp 1731220505
transform 1 0 680 0 -1 5160
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_580_6
timestamp 1731220505
transform 1 0 584 0 1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_579_6
timestamp 1731220505
transform 1 0 736 0 1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_578_6
timestamp 1731220505
transform 1 0 896 0 1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_577_6
timestamp 1731220505
transform 1 0 1240 0 1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_576_6
timestamp 1731220505
transform 1 0 1064 0 1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_575_6
timestamp 1731220505
transform 1 0 1008 0 -1 5400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_574_6
timestamp 1731220505
transform 1 0 872 0 -1 5400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_573_6
timestamp 1731220505
transform 1 0 1152 0 -1 5400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_572_6
timestamp 1731220505
transform 1 0 1328 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_571_6
timestamp 1731220505
transform 1 0 1304 0 -1 5400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_570_6
timestamp 1731220505
transform 1 0 1632 0 -1 5400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_569_6
timestamp 1731220505
transform 1 0 1464 0 -1 5400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_568_6
timestamp 1731220505
transform 1 0 1424 0 1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_567_6
timestamp 1731220505
transform 1 0 1416 0 -1 5160
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_566_6
timestamp 1731220505
transform 1 0 1232 0 -1 5160
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_565_6
timestamp 1731220505
transform 1 0 1368 0 1 4932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_564_6
timestamp 1731220505
transform 1 0 1656 0 1 4932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_563_6
timestamp 1731220505
transform 1 0 1600 0 -1 5160
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_562_6
timestamp 1731220505
transform 1 0 1784 0 -1 5160
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_561_6
timestamp 1731220505
transform 1 0 1616 0 1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_560_6
timestamp 1731220505
transform 1 0 1784 0 1 5172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_559_6
timestamp 1731220505
transform 1 0 1784 0 -1 5400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_558_6
timestamp 1731220505
transform 1 0 1992 0 -1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_557_6
timestamp 1731220505
transform 1 0 2688 0 -1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_556_6
timestamp 1731220505
transform 1 0 2496 0 -1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_555_6
timestamp 1731220505
transform 1 0 2432 0 1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_554_6
timestamp 1731220505
transform 1 0 2200 0 1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_553_6
timestamp 1731220505
transform 1 0 2656 0 1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_552_6
timestamp 1731220505
transform 1 0 2632 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_551_6
timestamp 1731220505
transform 1 0 2480 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_550_6
timestamp 1731220505
transform 1 0 2784 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_549_6
timestamp 1731220505
transform 1 0 2944 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_548_6
timestamp 1731220505
transform 1 0 3112 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_547_6
timestamp 1731220505
transform 1 0 3288 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_546_6
timestamp 1731220505
transform 1 0 3464 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_545_6
timestamp 1731220505
transform 1 0 3648 0 1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_544_6
timestamp 1731220505
transform 1 0 3472 0 1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_543_6
timestamp 1731220505
transform 1 0 3272 0 1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_542_6
timestamp 1731220505
transform 1 0 3072 0 1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_541_6
timestamp 1731220505
transform 1 0 2864 0 1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_540_6
timestamp 1731220505
transform 1 0 3280 0 -1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_539_6
timestamp 1731220505
transform 1 0 3080 0 -1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_538_6
timestamp 1731220505
transform 1 0 2880 0 -1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_537_6
timestamp 1731220505
transform 1 0 2856 0 1 5240
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_536_6
timestamp 1731220505
transform 1 0 2560 0 -1 5240
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_535_6
timestamp 1731220505
transform 1 0 2512 0 1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_534_6
timestamp 1731220505
transform 1 0 2752 0 1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_533_6
timestamp 1731220505
transform 1 0 2712 0 -1 4984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_532_6
timestamp 1731220505
transform 1 0 2864 0 -1 4984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_531_6
timestamp 1731220505
transform 1 0 2720 0 1 4752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_530_6
timestamp 1731220505
transform 1 0 2568 0 1 4752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_529_6
timestamp 1731220505
transform 1 0 2424 0 1 4752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_528_6
timestamp 1731220505
transform 1 0 2568 0 -1 4984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_527_6
timestamp 1731220505
transform 1 0 2424 0 -1 4984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_526_6
timestamp 1731220505
transform 1 0 2288 0 -1 4984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_525_6
timestamp 1731220505
transform 1 0 2152 0 -1 4984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_524_6
timestamp 1731220505
transform 1 0 2264 0 1 5016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_523_6
timestamp 1731220505
transform 1 0 2208 0 -1 5240
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_522_6
timestamp 1731220505
transform 1 0 2048 0 1 5240
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_521_6
timestamp 1731220505
transform 1 0 2456 0 1 5240
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_520_6
timestamp 1731220505
transform 1 0 2312 0 -1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_519_6
timestamp 1731220505
transform 1 0 2136 0 -1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_518_6
timestamp 1731220505
transform 1 0 1992 0 1 5488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_517_6
timestamp 1731220505
transform 1 0 1784 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_516_6
timestamp 1731220505
transform 1 0 1720 0 1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_515_6
timestamp 1731220505
transform 1 0 1448 0 1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_514_6
timestamp 1731220505
transform 1 0 1176 0 1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_513_6
timestamp 1731220505
transform 1 0 1552 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_512_6
timestamp 1731220505
transform 1 0 1296 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_511_6
timestamp 1731220505
transform 1 0 1192 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_510_6
timestamp 1731220505
transform 1 0 1056 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_59_6
timestamp 1731220505
transform 1 0 920 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_58_6
timestamp 1731220505
transform 1 0 784 0 1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_57_6
timestamp 1731220505
transform 1 0 1056 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_56_6
timestamp 1731220505
transform 1 0 824 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_55_6
timestamp 1731220505
transform 1 0 616 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_54_6
timestamp 1731220505
transform 1 0 424 0 -1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_53_6
timestamp 1731220505
transform 1 0 904 0 1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_52_6
timestamp 1731220505
transform 1 0 632 0 1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_51_6
timestamp 1731220505
transform 1 0 368 0 1 5644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_50_6
timestamp 1731220505
transform 1 0 128 0 1 5644
box 3 5 132 108
<< end >>
