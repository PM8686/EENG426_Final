magic
tech sky130l
timestamp 1731220588
<< m2 >>
rect 238 3633 244 3634
rect 238 3629 239 3633
rect 243 3629 244 3633
rect 238 3628 244 3629
rect 326 3633 332 3634
rect 326 3629 327 3633
rect 331 3629 332 3633
rect 326 3628 332 3629
rect 414 3633 420 3634
rect 414 3629 415 3633
rect 419 3629 420 3633
rect 414 3628 420 3629
rect 502 3633 508 3634
rect 502 3629 503 3633
rect 507 3629 508 3633
rect 502 3628 508 3629
rect 590 3633 596 3634
rect 590 3629 591 3633
rect 595 3629 596 3633
rect 590 3628 596 3629
rect 678 3633 684 3634
rect 678 3629 679 3633
rect 683 3629 684 3633
rect 678 3628 684 3629
rect 110 3620 116 3621
rect 110 3616 111 3620
rect 115 3616 116 3620
rect 110 3615 116 3616
rect 1822 3620 1828 3621
rect 1822 3616 1823 3620
rect 1827 3616 1828 3620
rect 1822 3615 1828 3616
rect 110 3603 116 3604
rect 110 3599 111 3603
rect 115 3599 116 3603
rect 110 3598 116 3599
rect 1822 3603 1828 3604
rect 1822 3599 1823 3603
rect 1827 3599 1828 3603
rect 1822 3598 1828 3599
rect 230 3593 236 3594
rect 230 3589 231 3593
rect 235 3589 236 3593
rect 230 3588 236 3589
rect 318 3593 324 3594
rect 318 3589 319 3593
rect 323 3589 324 3593
rect 318 3588 324 3589
rect 406 3593 412 3594
rect 406 3589 407 3593
rect 411 3589 412 3593
rect 406 3588 412 3589
rect 494 3593 500 3594
rect 494 3589 495 3593
rect 499 3589 500 3593
rect 494 3588 500 3589
rect 582 3593 588 3594
rect 582 3589 583 3593
rect 587 3589 588 3593
rect 582 3588 588 3589
rect 670 3593 676 3594
rect 670 3589 671 3593
rect 675 3589 676 3593
rect 670 3588 676 3589
rect 1886 3575 1892 3576
rect 1886 3571 1887 3575
rect 1891 3571 1892 3575
rect 1886 3570 1892 3571
rect 1974 3575 1980 3576
rect 1974 3571 1975 3575
rect 1979 3571 1980 3575
rect 1974 3570 1980 3571
rect 2062 3575 2068 3576
rect 2062 3571 2063 3575
rect 2067 3571 2068 3575
rect 2062 3570 2068 3571
rect 2150 3575 2156 3576
rect 2150 3571 2151 3575
rect 2155 3571 2156 3575
rect 2150 3570 2156 3571
rect 2238 3575 2244 3576
rect 2238 3571 2239 3575
rect 2243 3571 2244 3575
rect 2238 3570 2244 3571
rect 2326 3575 2332 3576
rect 2326 3571 2327 3575
rect 2331 3571 2332 3575
rect 2326 3570 2332 3571
rect 2414 3575 2420 3576
rect 2414 3571 2415 3575
rect 2419 3571 2420 3575
rect 2414 3570 2420 3571
rect 2502 3575 2508 3576
rect 2502 3571 2503 3575
rect 2507 3571 2508 3575
rect 2502 3570 2508 3571
rect 2590 3575 2596 3576
rect 2590 3571 2591 3575
rect 2595 3571 2596 3575
rect 2590 3570 2596 3571
rect 2678 3575 2684 3576
rect 2678 3571 2679 3575
rect 2683 3571 2684 3575
rect 2678 3570 2684 3571
rect 2766 3575 2772 3576
rect 2766 3571 2767 3575
rect 2771 3571 2772 3575
rect 2766 3570 2772 3571
rect 2854 3575 2860 3576
rect 2854 3571 2855 3575
rect 2859 3571 2860 3575
rect 2854 3570 2860 3571
rect 2942 3575 2948 3576
rect 2942 3571 2943 3575
rect 2947 3571 2948 3575
rect 2942 3570 2948 3571
rect 3030 3575 3036 3576
rect 3030 3571 3031 3575
rect 3035 3571 3036 3575
rect 3030 3570 3036 3571
rect 3118 3575 3124 3576
rect 3118 3571 3119 3575
rect 3123 3571 3124 3575
rect 3118 3570 3124 3571
rect 3206 3575 3212 3576
rect 3206 3571 3207 3575
rect 3211 3571 3212 3575
rect 3206 3570 3212 3571
rect 3294 3575 3300 3576
rect 3294 3571 3295 3575
rect 3299 3571 3300 3575
rect 3294 3570 3300 3571
rect 1862 3565 1868 3566
rect 246 3563 252 3564
rect 246 3559 247 3563
rect 251 3559 252 3563
rect 246 3558 252 3559
rect 398 3563 404 3564
rect 398 3559 399 3563
rect 403 3559 404 3563
rect 398 3558 404 3559
rect 542 3563 548 3564
rect 542 3559 543 3563
rect 547 3559 548 3563
rect 542 3558 548 3559
rect 686 3563 692 3564
rect 686 3559 687 3563
rect 691 3559 692 3563
rect 686 3558 692 3559
rect 822 3563 828 3564
rect 822 3559 823 3563
rect 827 3559 828 3563
rect 822 3558 828 3559
rect 950 3563 956 3564
rect 950 3559 951 3563
rect 955 3559 956 3563
rect 950 3558 956 3559
rect 1078 3563 1084 3564
rect 1078 3559 1079 3563
rect 1083 3559 1084 3563
rect 1078 3558 1084 3559
rect 1198 3563 1204 3564
rect 1198 3559 1199 3563
rect 1203 3559 1204 3563
rect 1198 3558 1204 3559
rect 1310 3563 1316 3564
rect 1310 3559 1311 3563
rect 1315 3559 1316 3563
rect 1310 3558 1316 3559
rect 1422 3563 1428 3564
rect 1422 3559 1423 3563
rect 1427 3559 1428 3563
rect 1422 3558 1428 3559
rect 1542 3563 1548 3564
rect 1542 3559 1543 3563
rect 1547 3559 1548 3563
rect 1862 3561 1863 3565
rect 1867 3561 1868 3565
rect 1862 3560 1868 3561
rect 3574 3565 3580 3566
rect 3574 3561 3575 3565
rect 3579 3561 3580 3565
rect 3574 3560 3580 3561
rect 1542 3558 1548 3559
rect 110 3553 116 3554
rect 110 3549 111 3553
rect 115 3549 116 3553
rect 110 3548 116 3549
rect 1822 3553 1828 3554
rect 1822 3549 1823 3553
rect 1827 3549 1828 3553
rect 1822 3548 1828 3549
rect 1862 3548 1868 3549
rect 1862 3544 1863 3548
rect 1867 3544 1868 3548
rect 1862 3543 1868 3544
rect 3574 3548 3580 3549
rect 3574 3544 3575 3548
rect 3579 3544 3580 3548
rect 3574 3543 3580 3544
rect 110 3536 116 3537
rect 110 3532 111 3536
rect 115 3532 116 3536
rect 110 3531 116 3532
rect 1822 3536 1828 3537
rect 1822 3532 1823 3536
rect 1827 3532 1828 3536
rect 1822 3531 1828 3532
rect 1894 3535 1900 3536
rect 1894 3531 1895 3535
rect 1899 3531 1900 3535
rect 1894 3530 1900 3531
rect 1982 3535 1988 3536
rect 1982 3531 1983 3535
rect 1987 3531 1988 3535
rect 1982 3530 1988 3531
rect 2070 3535 2076 3536
rect 2070 3531 2071 3535
rect 2075 3531 2076 3535
rect 2070 3530 2076 3531
rect 2158 3535 2164 3536
rect 2158 3531 2159 3535
rect 2163 3531 2164 3535
rect 2158 3530 2164 3531
rect 2246 3535 2252 3536
rect 2246 3531 2247 3535
rect 2251 3531 2252 3535
rect 2246 3530 2252 3531
rect 2334 3535 2340 3536
rect 2334 3531 2335 3535
rect 2339 3531 2340 3535
rect 2334 3530 2340 3531
rect 2422 3535 2428 3536
rect 2422 3531 2423 3535
rect 2427 3531 2428 3535
rect 2422 3530 2428 3531
rect 2510 3535 2516 3536
rect 2510 3531 2511 3535
rect 2515 3531 2516 3535
rect 2510 3530 2516 3531
rect 2598 3535 2604 3536
rect 2598 3531 2599 3535
rect 2603 3531 2604 3535
rect 2598 3530 2604 3531
rect 2686 3535 2692 3536
rect 2686 3531 2687 3535
rect 2691 3531 2692 3535
rect 2686 3530 2692 3531
rect 2774 3535 2780 3536
rect 2774 3531 2775 3535
rect 2779 3531 2780 3535
rect 2774 3530 2780 3531
rect 2862 3535 2868 3536
rect 2862 3531 2863 3535
rect 2867 3531 2868 3535
rect 2862 3530 2868 3531
rect 2950 3535 2956 3536
rect 2950 3531 2951 3535
rect 2955 3531 2956 3535
rect 2950 3530 2956 3531
rect 3038 3535 3044 3536
rect 3038 3531 3039 3535
rect 3043 3531 3044 3535
rect 3038 3530 3044 3531
rect 3126 3535 3132 3536
rect 3126 3531 3127 3535
rect 3131 3531 3132 3535
rect 3126 3530 3132 3531
rect 3214 3535 3220 3536
rect 3214 3531 3215 3535
rect 3219 3531 3220 3535
rect 3214 3530 3220 3531
rect 3302 3535 3308 3536
rect 3302 3531 3303 3535
rect 3307 3531 3308 3535
rect 3302 3530 3308 3531
rect 254 3523 260 3524
rect 254 3519 255 3523
rect 259 3519 260 3523
rect 254 3518 260 3519
rect 406 3523 412 3524
rect 406 3519 407 3523
rect 411 3519 412 3523
rect 406 3518 412 3519
rect 550 3523 556 3524
rect 550 3519 551 3523
rect 555 3519 556 3523
rect 550 3518 556 3519
rect 694 3523 700 3524
rect 694 3519 695 3523
rect 699 3519 700 3523
rect 694 3518 700 3519
rect 830 3523 836 3524
rect 830 3519 831 3523
rect 835 3519 836 3523
rect 830 3518 836 3519
rect 958 3523 964 3524
rect 958 3519 959 3523
rect 963 3519 964 3523
rect 958 3518 964 3519
rect 1086 3523 1092 3524
rect 1086 3519 1087 3523
rect 1091 3519 1092 3523
rect 1086 3518 1092 3519
rect 1206 3523 1212 3524
rect 1206 3519 1207 3523
rect 1211 3519 1212 3523
rect 1206 3518 1212 3519
rect 1318 3523 1324 3524
rect 1318 3519 1319 3523
rect 1323 3519 1324 3523
rect 1318 3518 1324 3519
rect 1430 3523 1436 3524
rect 1430 3519 1431 3523
rect 1435 3519 1436 3523
rect 1430 3518 1436 3519
rect 1550 3523 1556 3524
rect 1550 3519 1551 3523
rect 1555 3519 1556 3523
rect 1550 3518 1556 3519
rect 1910 3493 1916 3494
rect 182 3489 188 3490
rect 182 3485 183 3489
rect 187 3485 188 3489
rect 182 3484 188 3485
rect 350 3489 356 3490
rect 350 3485 351 3489
rect 355 3485 356 3489
rect 350 3484 356 3485
rect 518 3489 524 3490
rect 518 3485 519 3489
rect 523 3485 524 3489
rect 518 3484 524 3485
rect 678 3489 684 3490
rect 678 3485 679 3489
rect 683 3485 684 3489
rect 678 3484 684 3485
rect 830 3489 836 3490
rect 830 3485 831 3489
rect 835 3485 836 3489
rect 830 3484 836 3485
rect 966 3489 972 3490
rect 966 3485 967 3489
rect 971 3485 972 3489
rect 966 3484 972 3485
rect 1094 3489 1100 3490
rect 1094 3485 1095 3489
rect 1099 3485 1100 3489
rect 1094 3484 1100 3485
rect 1214 3489 1220 3490
rect 1214 3485 1215 3489
rect 1219 3485 1220 3489
rect 1214 3484 1220 3485
rect 1334 3489 1340 3490
rect 1334 3485 1335 3489
rect 1339 3485 1340 3489
rect 1334 3484 1340 3485
rect 1454 3489 1460 3490
rect 1454 3485 1455 3489
rect 1459 3485 1460 3489
rect 1454 3484 1460 3485
rect 1574 3489 1580 3490
rect 1574 3485 1575 3489
rect 1579 3485 1580 3489
rect 1910 3489 1911 3493
rect 1915 3489 1916 3493
rect 1910 3488 1916 3489
rect 2014 3493 2020 3494
rect 2014 3489 2015 3493
rect 2019 3489 2020 3493
rect 2014 3488 2020 3489
rect 2134 3493 2140 3494
rect 2134 3489 2135 3493
rect 2139 3489 2140 3493
rect 2134 3488 2140 3489
rect 2262 3493 2268 3494
rect 2262 3489 2263 3493
rect 2267 3489 2268 3493
rect 2262 3488 2268 3489
rect 2390 3493 2396 3494
rect 2390 3489 2391 3493
rect 2395 3489 2396 3493
rect 2390 3488 2396 3489
rect 2526 3493 2532 3494
rect 2526 3489 2527 3493
rect 2531 3489 2532 3493
rect 2526 3488 2532 3489
rect 2662 3493 2668 3494
rect 2662 3489 2663 3493
rect 2667 3489 2668 3493
rect 2662 3488 2668 3489
rect 2798 3493 2804 3494
rect 2798 3489 2799 3493
rect 2803 3489 2804 3493
rect 2798 3488 2804 3489
rect 2942 3493 2948 3494
rect 2942 3489 2943 3493
rect 2947 3489 2948 3493
rect 2942 3488 2948 3489
rect 3086 3493 3092 3494
rect 3086 3489 3087 3493
rect 3091 3489 3092 3493
rect 3086 3488 3092 3489
rect 1574 3484 1580 3485
rect 1862 3480 1868 3481
rect 110 3476 116 3477
rect 110 3472 111 3476
rect 115 3472 116 3476
rect 110 3471 116 3472
rect 1822 3476 1828 3477
rect 1822 3472 1823 3476
rect 1827 3472 1828 3476
rect 1862 3476 1863 3480
rect 1867 3476 1868 3480
rect 1862 3475 1868 3476
rect 3574 3480 3580 3481
rect 3574 3476 3575 3480
rect 3579 3476 3580 3480
rect 3574 3475 3580 3476
rect 1822 3471 1828 3472
rect 1862 3463 1868 3464
rect 110 3459 116 3460
rect 110 3455 111 3459
rect 115 3455 116 3459
rect 110 3454 116 3455
rect 1822 3459 1828 3460
rect 1822 3455 1823 3459
rect 1827 3455 1828 3459
rect 1862 3459 1863 3463
rect 1867 3459 1868 3463
rect 1862 3458 1868 3459
rect 3574 3463 3580 3464
rect 3574 3459 3575 3463
rect 3579 3459 3580 3463
rect 3574 3458 3580 3459
rect 1822 3454 1828 3455
rect 1902 3453 1908 3454
rect 174 3449 180 3450
rect 174 3445 175 3449
rect 179 3445 180 3449
rect 174 3444 180 3445
rect 342 3449 348 3450
rect 342 3445 343 3449
rect 347 3445 348 3449
rect 342 3444 348 3445
rect 510 3449 516 3450
rect 510 3445 511 3449
rect 515 3445 516 3449
rect 510 3444 516 3445
rect 670 3449 676 3450
rect 670 3445 671 3449
rect 675 3445 676 3449
rect 670 3444 676 3445
rect 822 3449 828 3450
rect 822 3445 823 3449
rect 827 3445 828 3449
rect 822 3444 828 3445
rect 958 3449 964 3450
rect 958 3445 959 3449
rect 963 3445 964 3449
rect 958 3444 964 3445
rect 1086 3449 1092 3450
rect 1086 3445 1087 3449
rect 1091 3445 1092 3449
rect 1086 3444 1092 3445
rect 1206 3449 1212 3450
rect 1206 3445 1207 3449
rect 1211 3445 1212 3449
rect 1206 3444 1212 3445
rect 1326 3449 1332 3450
rect 1326 3445 1327 3449
rect 1331 3445 1332 3449
rect 1326 3444 1332 3445
rect 1446 3449 1452 3450
rect 1446 3445 1447 3449
rect 1451 3445 1452 3449
rect 1446 3444 1452 3445
rect 1566 3449 1572 3450
rect 1566 3445 1567 3449
rect 1571 3445 1572 3449
rect 1902 3449 1903 3453
rect 1907 3449 1908 3453
rect 1902 3448 1908 3449
rect 2006 3453 2012 3454
rect 2006 3449 2007 3453
rect 2011 3449 2012 3453
rect 2006 3448 2012 3449
rect 2126 3453 2132 3454
rect 2126 3449 2127 3453
rect 2131 3449 2132 3453
rect 2126 3448 2132 3449
rect 2254 3453 2260 3454
rect 2254 3449 2255 3453
rect 2259 3449 2260 3453
rect 2254 3448 2260 3449
rect 2382 3453 2388 3454
rect 2382 3449 2383 3453
rect 2387 3449 2388 3453
rect 2382 3448 2388 3449
rect 2518 3453 2524 3454
rect 2518 3449 2519 3453
rect 2523 3449 2524 3453
rect 2518 3448 2524 3449
rect 2654 3453 2660 3454
rect 2654 3449 2655 3453
rect 2659 3449 2660 3453
rect 2654 3448 2660 3449
rect 2790 3453 2796 3454
rect 2790 3449 2791 3453
rect 2795 3449 2796 3453
rect 2790 3448 2796 3449
rect 2934 3453 2940 3454
rect 2934 3449 2935 3453
rect 2939 3449 2940 3453
rect 2934 3448 2940 3449
rect 3078 3453 3084 3454
rect 3078 3449 3079 3453
rect 3083 3449 3084 3453
rect 3078 3448 3084 3449
rect 1566 3444 1572 3445
rect 134 3427 140 3428
rect 134 3423 135 3427
rect 139 3423 140 3427
rect 134 3422 140 3423
rect 254 3427 260 3428
rect 254 3423 255 3427
rect 259 3423 260 3427
rect 254 3422 260 3423
rect 414 3427 420 3428
rect 414 3423 415 3427
rect 419 3423 420 3427
rect 414 3422 420 3423
rect 582 3427 588 3428
rect 582 3423 583 3427
rect 587 3423 588 3427
rect 582 3422 588 3423
rect 758 3427 764 3428
rect 758 3423 759 3427
rect 763 3423 764 3427
rect 758 3422 764 3423
rect 934 3427 940 3428
rect 934 3423 935 3427
rect 939 3423 940 3427
rect 934 3422 940 3423
rect 1110 3427 1116 3428
rect 1110 3423 1111 3427
rect 1115 3423 1116 3427
rect 1110 3422 1116 3423
rect 1294 3427 1300 3428
rect 1294 3423 1295 3427
rect 1299 3423 1300 3427
rect 1294 3422 1300 3423
rect 1478 3427 1484 3428
rect 1478 3423 1479 3427
rect 1483 3423 1484 3427
rect 1478 3422 1484 3423
rect 1910 3423 1916 3424
rect 1910 3419 1911 3423
rect 1915 3419 1916 3423
rect 1910 3418 1916 3419
rect 2070 3423 2076 3424
rect 2070 3419 2071 3423
rect 2075 3419 2076 3423
rect 2070 3418 2076 3419
rect 2222 3423 2228 3424
rect 2222 3419 2223 3423
rect 2227 3419 2228 3423
rect 2222 3418 2228 3419
rect 2366 3423 2372 3424
rect 2366 3419 2367 3423
rect 2371 3419 2372 3423
rect 2366 3418 2372 3419
rect 2502 3423 2508 3424
rect 2502 3419 2503 3423
rect 2507 3419 2508 3423
rect 2502 3418 2508 3419
rect 2630 3423 2636 3424
rect 2630 3419 2631 3423
rect 2635 3419 2636 3423
rect 2630 3418 2636 3419
rect 2758 3423 2764 3424
rect 2758 3419 2759 3423
rect 2763 3419 2764 3423
rect 2758 3418 2764 3419
rect 2886 3423 2892 3424
rect 2886 3419 2887 3423
rect 2891 3419 2892 3423
rect 2886 3418 2892 3419
rect 3022 3423 3028 3424
rect 3022 3419 3023 3423
rect 3027 3419 3028 3423
rect 3022 3418 3028 3419
rect 110 3417 116 3418
rect 110 3413 111 3417
rect 115 3413 116 3417
rect 110 3412 116 3413
rect 1822 3417 1828 3418
rect 1822 3413 1823 3417
rect 1827 3413 1828 3417
rect 1822 3412 1828 3413
rect 1862 3413 1868 3414
rect 1862 3409 1863 3413
rect 1867 3409 1868 3413
rect 1862 3408 1868 3409
rect 3574 3413 3580 3414
rect 3574 3409 3575 3413
rect 3579 3409 3580 3413
rect 3574 3408 3580 3409
rect 110 3400 116 3401
rect 110 3396 111 3400
rect 115 3396 116 3400
rect 110 3395 116 3396
rect 1822 3400 1828 3401
rect 1822 3396 1823 3400
rect 1827 3396 1828 3400
rect 1822 3395 1828 3396
rect 1862 3396 1868 3397
rect 1862 3392 1863 3396
rect 1867 3392 1868 3396
rect 1862 3391 1868 3392
rect 3574 3396 3580 3397
rect 3574 3392 3575 3396
rect 3579 3392 3580 3396
rect 3574 3391 3580 3392
rect 142 3387 148 3388
rect 142 3383 143 3387
rect 147 3383 148 3387
rect 142 3382 148 3383
rect 262 3387 268 3388
rect 262 3383 263 3387
rect 267 3383 268 3387
rect 262 3382 268 3383
rect 422 3387 428 3388
rect 422 3383 423 3387
rect 427 3383 428 3387
rect 422 3382 428 3383
rect 590 3387 596 3388
rect 590 3383 591 3387
rect 595 3383 596 3387
rect 590 3382 596 3383
rect 766 3387 772 3388
rect 766 3383 767 3387
rect 771 3383 772 3387
rect 766 3382 772 3383
rect 942 3387 948 3388
rect 942 3383 943 3387
rect 947 3383 948 3387
rect 942 3382 948 3383
rect 1118 3387 1124 3388
rect 1118 3383 1119 3387
rect 1123 3383 1124 3387
rect 1118 3382 1124 3383
rect 1302 3387 1308 3388
rect 1302 3383 1303 3387
rect 1307 3383 1308 3387
rect 1302 3382 1308 3383
rect 1486 3387 1492 3388
rect 1486 3383 1487 3387
rect 1491 3383 1492 3387
rect 1486 3382 1492 3383
rect 1918 3383 1924 3384
rect 1918 3379 1919 3383
rect 1923 3379 1924 3383
rect 1918 3378 1924 3379
rect 2078 3383 2084 3384
rect 2078 3379 2079 3383
rect 2083 3379 2084 3383
rect 2078 3378 2084 3379
rect 2230 3383 2236 3384
rect 2230 3379 2231 3383
rect 2235 3379 2236 3383
rect 2230 3378 2236 3379
rect 2374 3383 2380 3384
rect 2374 3379 2375 3383
rect 2379 3379 2380 3383
rect 2374 3378 2380 3379
rect 2510 3383 2516 3384
rect 2510 3379 2511 3383
rect 2515 3379 2516 3383
rect 2510 3378 2516 3379
rect 2638 3383 2644 3384
rect 2638 3379 2639 3383
rect 2643 3379 2644 3383
rect 2638 3378 2644 3379
rect 2766 3383 2772 3384
rect 2766 3379 2767 3383
rect 2771 3379 2772 3383
rect 2766 3378 2772 3379
rect 2894 3383 2900 3384
rect 2894 3379 2895 3383
rect 2899 3379 2900 3383
rect 2894 3378 2900 3379
rect 3030 3383 3036 3384
rect 3030 3379 3031 3383
rect 3035 3379 3036 3383
rect 3030 3378 3036 3379
rect 206 3345 212 3346
rect 206 3341 207 3345
rect 211 3341 212 3345
rect 206 3340 212 3341
rect 366 3345 372 3346
rect 366 3341 367 3345
rect 371 3341 372 3345
rect 366 3340 372 3341
rect 534 3345 540 3346
rect 534 3341 535 3345
rect 539 3341 540 3345
rect 534 3340 540 3341
rect 694 3345 700 3346
rect 694 3341 695 3345
rect 699 3341 700 3345
rect 694 3340 700 3341
rect 854 3345 860 3346
rect 854 3341 855 3345
rect 859 3341 860 3345
rect 854 3340 860 3341
rect 998 3345 1004 3346
rect 998 3341 999 3345
rect 1003 3341 1004 3345
rect 998 3340 1004 3341
rect 1142 3345 1148 3346
rect 1142 3341 1143 3345
rect 1147 3341 1148 3345
rect 1142 3340 1148 3341
rect 1278 3345 1284 3346
rect 1278 3341 1279 3345
rect 1283 3341 1284 3345
rect 1278 3340 1284 3341
rect 1414 3345 1420 3346
rect 1414 3341 1415 3345
rect 1419 3341 1420 3345
rect 1414 3340 1420 3341
rect 1558 3345 1564 3346
rect 1558 3341 1559 3345
rect 1563 3341 1564 3345
rect 1558 3340 1564 3341
rect 1894 3345 1900 3346
rect 1894 3341 1895 3345
rect 1899 3341 1900 3345
rect 1894 3340 1900 3341
rect 2046 3345 2052 3346
rect 2046 3341 2047 3345
rect 2051 3341 2052 3345
rect 2046 3340 2052 3341
rect 2206 3345 2212 3346
rect 2206 3341 2207 3345
rect 2211 3341 2212 3345
rect 2206 3340 2212 3341
rect 2366 3345 2372 3346
rect 2366 3341 2367 3345
rect 2371 3341 2372 3345
rect 2366 3340 2372 3341
rect 2534 3345 2540 3346
rect 2534 3341 2535 3345
rect 2539 3341 2540 3345
rect 2534 3340 2540 3341
rect 2702 3345 2708 3346
rect 2702 3341 2703 3345
rect 2707 3341 2708 3345
rect 2702 3340 2708 3341
rect 2878 3345 2884 3346
rect 2878 3341 2879 3345
rect 2883 3341 2884 3345
rect 2878 3340 2884 3341
rect 3054 3345 3060 3346
rect 3054 3341 3055 3345
rect 3059 3341 3060 3345
rect 3054 3340 3060 3341
rect 110 3332 116 3333
rect 110 3328 111 3332
rect 115 3328 116 3332
rect 110 3327 116 3328
rect 1822 3332 1828 3333
rect 1822 3328 1823 3332
rect 1827 3328 1828 3332
rect 1822 3327 1828 3328
rect 1862 3332 1868 3333
rect 1862 3328 1863 3332
rect 1867 3328 1868 3332
rect 1862 3327 1868 3328
rect 3574 3332 3580 3333
rect 3574 3328 3575 3332
rect 3579 3328 3580 3332
rect 3574 3327 3580 3328
rect 110 3315 116 3316
rect 110 3311 111 3315
rect 115 3311 116 3315
rect 110 3310 116 3311
rect 1822 3315 1828 3316
rect 1822 3311 1823 3315
rect 1827 3311 1828 3315
rect 1822 3310 1828 3311
rect 1862 3315 1868 3316
rect 1862 3311 1863 3315
rect 1867 3311 1868 3315
rect 1862 3310 1868 3311
rect 3574 3315 3580 3316
rect 3574 3311 3575 3315
rect 3579 3311 3580 3315
rect 3574 3310 3580 3311
rect 198 3305 204 3306
rect 198 3301 199 3305
rect 203 3301 204 3305
rect 198 3300 204 3301
rect 358 3305 364 3306
rect 358 3301 359 3305
rect 363 3301 364 3305
rect 358 3300 364 3301
rect 526 3305 532 3306
rect 526 3301 527 3305
rect 531 3301 532 3305
rect 526 3300 532 3301
rect 686 3305 692 3306
rect 686 3301 687 3305
rect 691 3301 692 3305
rect 686 3300 692 3301
rect 846 3305 852 3306
rect 846 3301 847 3305
rect 851 3301 852 3305
rect 846 3300 852 3301
rect 990 3305 996 3306
rect 990 3301 991 3305
rect 995 3301 996 3305
rect 990 3300 996 3301
rect 1134 3305 1140 3306
rect 1134 3301 1135 3305
rect 1139 3301 1140 3305
rect 1134 3300 1140 3301
rect 1270 3305 1276 3306
rect 1270 3301 1271 3305
rect 1275 3301 1276 3305
rect 1270 3300 1276 3301
rect 1406 3305 1412 3306
rect 1406 3301 1407 3305
rect 1411 3301 1412 3305
rect 1406 3300 1412 3301
rect 1550 3305 1556 3306
rect 1550 3301 1551 3305
rect 1555 3301 1556 3305
rect 1550 3300 1556 3301
rect 1886 3305 1892 3306
rect 1886 3301 1887 3305
rect 1891 3301 1892 3305
rect 1886 3300 1892 3301
rect 2038 3305 2044 3306
rect 2038 3301 2039 3305
rect 2043 3301 2044 3305
rect 2038 3300 2044 3301
rect 2198 3305 2204 3306
rect 2198 3301 2199 3305
rect 2203 3301 2204 3305
rect 2198 3300 2204 3301
rect 2358 3305 2364 3306
rect 2358 3301 2359 3305
rect 2363 3301 2364 3305
rect 2358 3300 2364 3301
rect 2526 3305 2532 3306
rect 2526 3301 2527 3305
rect 2531 3301 2532 3305
rect 2526 3300 2532 3301
rect 2694 3305 2700 3306
rect 2694 3301 2695 3305
rect 2699 3301 2700 3305
rect 2694 3300 2700 3301
rect 2870 3305 2876 3306
rect 2870 3301 2871 3305
rect 2875 3301 2876 3305
rect 2870 3300 2876 3301
rect 3046 3305 3052 3306
rect 3046 3301 3047 3305
rect 3051 3301 3052 3305
rect 3046 3300 3052 3301
rect 254 3279 260 3280
rect 254 3275 255 3279
rect 259 3275 260 3279
rect 254 3274 260 3275
rect 374 3279 380 3280
rect 374 3275 375 3279
rect 379 3275 380 3279
rect 374 3274 380 3275
rect 510 3279 516 3280
rect 510 3275 511 3279
rect 515 3275 516 3279
rect 510 3274 516 3275
rect 662 3279 668 3280
rect 662 3275 663 3279
rect 667 3275 668 3279
rect 662 3274 668 3275
rect 822 3279 828 3280
rect 822 3275 823 3279
rect 827 3275 828 3279
rect 822 3274 828 3275
rect 990 3279 996 3280
rect 990 3275 991 3279
rect 995 3275 996 3279
rect 990 3274 996 3275
rect 1166 3279 1172 3280
rect 1166 3275 1167 3279
rect 1171 3275 1172 3279
rect 1166 3274 1172 3275
rect 1342 3279 1348 3280
rect 1342 3275 1343 3279
rect 1347 3275 1348 3279
rect 1342 3274 1348 3275
rect 1518 3279 1524 3280
rect 1518 3275 1519 3279
rect 1523 3275 1524 3279
rect 1518 3274 1524 3275
rect 1886 3279 1892 3280
rect 1886 3275 1887 3279
rect 1891 3275 1892 3279
rect 1886 3274 1892 3275
rect 2062 3279 2068 3280
rect 2062 3275 2063 3279
rect 2067 3275 2068 3279
rect 2062 3274 2068 3275
rect 2262 3279 2268 3280
rect 2262 3275 2263 3279
rect 2267 3275 2268 3279
rect 2262 3274 2268 3275
rect 2454 3279 2460 3280
rect 2454 3275 2455 3279
rect 2459 3275 2460 3279
rect 2454 3274 2460 3275
rect 2638 3279 2644 3280
rect 2638 3275 2639 3279
rect 2643 3275 2644 3279
rect 2638 3274 2644 3275
rect 2814 3279 2820 3280
rect 2814 3275 2815 3279
rect 2819 3275 2820 3279
rect 2814 3274 2820 3275
rect 2982 3279 2988 3280
rect 2982 3275 2983 3279
rect 2987 3275 2988 3279
rect 2982 3274 2988 3275
rect 3150 3279 3156 3280
rect 3150 3275 3151 3279
rect 3155 3275 3156 3279
rect 3150 3274 3156 3275
rect 3318 3279 3324 3280
rect 3318 3275 3319 3279
rect 3323 3275 3324 3279
rect 3318 3274 3324 3275
rect 3478 3279 3484 3280
rect 3478 3275 3479 3279
rect 3483 3275 3484 3279
rect 3478 3274 3484 3275
rect 110 3269 116 3270
rect 110 3265 111 3269
rect 115 3265 116 3269
rect 110 3264 116 3265
rect 1822 3269 1828 3270
rect 1822 3265 1823 3269
rect 1827 3265 1828 3269
rect 1822 3264 1828 3265
rect 1862 3269 1868 3270
rect 1862 3265 1863 3269
rect 1867 3265 1868 3269
rect 1862 3264 1868 3265
rect 3574 3269 3580 3270
rect 3574 3265 3575 3269
rect 3579 3265 3580 3269
rect 3574 3264 3580 3265
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 110 3247 116 3248
rect 1822 3252 1828 3253
rect 1822 3248 1823 3252
rect 1827 3248 1828 3252
rect 1822 3247 1828 3248
rect 1862 3252 1868 3253
rect 1862 3248 1863 3252
rect 1867 3248 1868 3252
rect 1862 3247 1868 3248
rect 3574 3252 3580 3253
rect 3574 3248 3575 3252
rect 3579 3248 3580 3252
rect 3574 3247 3580 3248
rect 262 3239 268 3240
rect 262 3235 263 3239
rect 267 3235 268 3239
rect 262 3234 268 3235
rect 382 3239 388 3240
rect 382 3235 383 3239
rect 387 3235 388 3239
rect 382 3234 388 3235
rect 518 3239 524 3240
rect 518 3235 519 3239
rect 523 3235 524 3239
rect 518 3234 524 3235
rect 670 3239 676 3240
rect 670 3235 671 3239
rect 675 3235 676 3239
rect 670 3234 676 3235
rect 830 3239 836 3240
rect 830 3235 831 3239
rect 835 3235 836 3239
rect 830 3234 836 3235
rect 998 3239 1004 3240
rect 998 3235 999 3239
rect 1003 3235 1004 3239
rect 998 3234 1004 3235
rect 1174 3239 1180 3240
rect 1174 3235 1175 3239
rect 1179 3235 1180 3239
rect 1174 3234 1180 3235
rect 1350 3239 1356 3240
rect 1350 3235 1351 3239
rect 1355 3235 1356 3239
rect 1350 3234 1356 3235
rect 1526 3239 1532 3240
rect 1526 3235 1527 3239
rect 1531 3235 1532 3239
rect 1526 3234 1532 3235
rect 1894 3239 1900 3240
rect 1894 3235 1895 3239
rect 1899 3235 1900 3239
rect 1894 3234 1900 3235
rect 2070 3239 2076 3240
rect 2070 3235 2071 3239
rect 2075 3235 2076 3239
rect 2070 3234 2076 3235
rect 2270 3239 2276 3240
rect 2270 3235 2271 3239
rect 2275 3235 2276 3239
rect 2270 3234 2276 3235
rect 2462 3239 2468 3240
rect 2462 3235 2463 3239
rect 2467 3235 2468 3239
rect 2462 3234 2468 3235
rect 2646 3239 2652 3240
rect 2646 3235 2647 3239
rect 2651 3235 2652 3239
rect 2646 3234 2652 3235
rect 2822 3239 2828 3240
rect 2822 3235 2823 3239
rect 2827 3235 2828 3239
rect 2822 3234 2828 3235
rect 2990 3239 2996 3240
rect 2990 3235 2991 3239
rect 2995 3235 2996 3239
rect 2990 3234 2996 3235
rect 3158 3239 3164 3240
rect 3158 3235 3159 3239
rect 3163 3235 3164 3239
rect 3158 3234 3164 3235
rect 3326 3239 3332 3240
rect 3326 3235 3327 3239
rect 3331 3235 3332 3239
rect 3326 3234 3332 3235
rect 3486 3239 3492 3240
rect 3486 3235 3487 3239
rect 3491 3235 3492 3239
rect 3486 3234 3492 3235
rect 1894 3205 1900 3206
rect 430 3201 436 3202
rect 430 3197 431 3201
rect 435 3197 436 3201
rect 430 3196 436 3197
rect 550 3201 556 3202
rect 550 3197 551 3201
rect 555 3197 556 3201
rect 550 3196 556 3197
rect 670 3201 676 3202
rect 670 3197 671 3201
rect 675 3197 676 3201
rect 670 3196 676 3197
rect 798 3201 804 3202
rect 798 3197 799 3201
rect 803 3197 804 3201
rect 798 3196 804 3197
rect 934 3201 940 3202
rect 934 3197 935 3201
rect 939 3197 940 3201
rect 934 3196 940 3197
rect 1078 3201 1084 3202
rect 1078 3197 1079 3201
rect 1083 3197 1084 3201
rect 1078 3196 1084 3197
rect 1230 3201 1236 3202
rect 1230 3197 1231 3201
rect 1235 3197 1236 3201
rect 1230 3196 1236 3197
rect 1382 3201 1388 3202
rect 1382 3197 1383 3201
rect 1387 3197 1388 3201
rect 1382 3196 1388 3197
rect 1534 3201 1540 3202
rect 1534 3197 1535 3201
rect 1539 3197 1540 3201
rect 1894 3201 1895 3205
rect 1899 3201 1900 3205
rect 1894 3200 1900 3201
rect 2086 3205 2092 3206
rect 2086 3201 2087 3205
rect 2091 3201 2092 3205
rect 2086 3200 2092 3201
rect 2302 3205 2308 3206
rect 2302 3201 2303 3205
rect 2307 3201 2308 3205
rect 2302 3200 2308 3201
rect 2510 3205 2516 3206
rect 2510 3201 2511 3205
rect 2515 3201 2516 3205
rect 2510 3200 2516 3201
rect 2702 3205 2708 3206
rect 2702 3201 2703 3205
rect 2707 3201 2708 3205
rect 2702 3200 2708 3201
rect 2878 3205 2884 3206
rect 2878 3201 2879 3205
rect 2883 3201 2884 3205
rect 2878 3200 2884 3201
rect 3038 3205 3044 3206
rect 3038 3201 3039 3205
rect 3043 3201 3044 3205
rect 3038 3200 3044 3201
rect 3198 3205 3204 3206
rect 3198 3201 3199 3205
rect 3203 3201 3204 3205
rect 3198 3200 3204 3201
rect 3350 3205 3356 3206
rect 3350 3201 3351 3205
rect 3355 3201 3356 3205
rect 3350 3200 3356 3201
rect 3486 3205 3492 3206
rect 3486 3201 3487 3205
rect 3491 3201 3492 3205
rect 3486 3200 3492 3201
rect 1534 3196 1540 3197
rect 1862 3192 1868 3193
rect 110 3188 116 3189
rect 110 3184 111 3188
rect 115 3184 116 3188
rect 110 3183 116 3184
rect 1822 3188 1828 3189
rect 1822 3184 1823 3188
rect 1827 3184 1828 3188
rect 1862 3188 1863 3192
rect 1867 3188 1868 3192
rect 1862 3187 1868 3188
rect 3574 3192 3580 3193
rect 3574 3188 3575 3192
rect 3579 3188 3580 3192
rect 3574 3187 3580 3188
rect 1822 3183 1828 3184
rect 1862 3175 1868 3176
rect 110 3171 116 3172
rect 110 3167 111 3171
rect 115 3167 116 3171
rect 110 3166 116 3167
rect 1822 3171 1828 3172
rect 1822 3167 1823 3171
rect 1827 3167 1828 3171
rect 1862 3171 1863 3175
rect 1867 3171 1868 3175
rect 1862 3170 1868 3171
rect 3574 3175 3580 3176
rect 3574 3171 3575 3175
rect 3579 3171 3580 3175
rect 3574 3170 3580 3171
rect 1822 3166 1828 3167
rect 1886 3165 1892 3166
rect 422 3161 428 3162
rect 422 3157 423 3161
rect 427 3157 428 3161
rect 422 3156 428 3157
rect 542 3161 548 3162
rect 542 3157 543 3161
rect 547 3157 548 3161
rect 542 3156 548 3157
rect 662 3161 668 3162
rect 662 3157 663 3161
rect 667 3157 668 3161
rect 662 3156 668 3157
rect 790 3161 796 3162
rect 790 3157 791 3161
rect 795 3157 796 3161
rect 790 3156 796 3157
rect 926 3161 932 3162
rect 926 3157 927 3161
rect 931 3157 932 3161
rect 926 3156 932 3157
rect 1070 3161 1076 3162
rect 1070 3157 1071 3161
rect 1075 3157 1076 3161
rect 1070 3156 1076 3157
rect 1222 3161 1228 3162
rect 1222 3157 1223 3161
rect 1227 3157 1228 3161
rect 1222 3156 1228 3157
rect 1374 3161 1380 3162
rect 1374 3157 1375 3161
rect 1379 3157 1380 3161
rect 1374 3156 1380 3157
rect 1526 3161 1532 3162
rect 1526 3157 1527 3161
rect 1531 3157 1532 3161
rect 1886 3161 1887 3165
rect 1891 3161 1892 3165
rect 1886 3160 1892 3161
rect 2078 3165 2084 3166
rect 2078 3161 2079 3165
rect 2083 3161 2084 3165
rect 2078 3160 2084 3161
rect 2294 3165 2300 3166
rect 2294 3161 2295 3165
rect 2299 3161 2300 3165
rect 2294 3160 2300 3161
rect 2502 3165 2508 3166
rect 2502 3161 2503 3165
rect 2507 3161 2508 3165
rect 2502 3160 2508 3161
rect 2694 3165 2700 3166
rect 2694 3161 2695 3165
rect 2699 3161 2700 3165
rect 2694 3160 2700 3161
rect 2870 3165 2876 3166
rect 2870 3161 2871 3165
rect 2875 3161 2876 3165
rect 2870 3160 2876 3161
rect 3030 3165 3036 3166
rect 3030 3161 3031 3165
rect 3035 3161 3036 3165
rect 3030 3160 3036 3161
rect 3190 3165 3196 3166
rect 3190 3161 3191 3165
rect 3195 3161 3196 3165
rect 3190 3160 3196 3161
rect 3342 3165 3348 3166
rect 3342 3161 3343 3165
rect 3347 3161 3348 3165
rect 3342 3160 3348 3161
rect 3478 3165 3484 3166
rect 3478 3161 3479 3165
rect 3483 3161 3484 3165
rect 3478 3160 3484 3161
rect 1526 3156 1532 3157
rect 1886 3139 1892 3140
rect 462 3135 468 3136
rect 462 3131 463 3135
rect 467 3131 468 3135
rect 462 3130 468 3131
rect 550 3135 556 3136
rect 550 3131 551 3135
rect 555 3131 556 3135
rect 550 3130 556 3131
rect 638 3135 644 3136
rect 638 3131 639 3135
rect 643 3131 644 3135
rect 638 3130 644 3131
rect 734 3135 740 3136
rect 734 3131 735 3135
rect 739 3131 740 3135
rect 734 3130 740 3131
rect 846 3135 852 3136
rect 846 3131 847 3135
rect 851 3131 852 3135
rect 846 3130 852 3131
rect 966 3135 972 3136
rect 966 3131 967 3135
rect 971 3131 972 3135
rect 966 3130 972 3131
rect 1094 3135 1100 3136
rect 1094 3131 1095 3135
rect 1099 3131 1100 3135
rect 1094 3130 1100 3131
rect 1230 3135 1236 3136
rect 1230 3131 1231 3135
rect 1235 3131 1236 3135
rect 1230 3130 1236 3131
rect 1374 3135 1380 3136
rect 1374 3131 1375 3135
rect 1379 3131 1380 3135
rect 1374 3130 1380 3131
rect 1518 3135 1524 3136
rect 1518 3131 1519 3135
rect 1523 3131 1524 3135
rect 1886 3135 1887 3139
rect 1891 3135 1892 3139
rect 1886 3134 1892 3135
rect 2078 3139 2084 3140
rect 2078 3135 2079 3139
rect 2083 3135 2084 3139
rect 2078 3134 2084 3135
rect 2294 3139 2300 3140
rect 2294 3135 2295 3139
rect 2299 3135 2300 3139
rect 2294 3134 2300 3135
rect 2502 3139 2508 3140
rect 2502 3135 2503 3139
rect 2507 3135 2508 3139
rect 2502 3134 2508 3135
rect 2694 3139 2700 3140
rect 2694 3135 2695 3139
rect 2699 3135 2700 3139
rect 2694 3134 2700 3135
rect 2870 3139 2876 3140
rect 2870 3135 2871 3139
rect 2875 3135 2876 3139
rect 2870 3134 2876 3135
rect 3038 3139 3044 3140
rect 3038 3135 3039 3139
rect 3043 3135 3044 3139
rect 3038 3134 3044 3135
rect 3190 3139 3196 3140
rect 3190 3135 3191 3139
rect 3195 3135 3196 3139
rect 3190 3134 3196 3135
rect 3342 3139 3348 3140
rect 3342 3135 3343 3139
rect 3347 3135 3348 3139
rect 3342 3134 3348 3135
rect 3478 3139 3484 3140
rect 3478 3135 3479 3139
rect 3483 3135 3484 3139
rect 3478 3134 3484 3135
rect 1518 3130 1524 3131
rect 1862 3129 1868 3130
rect 110 3125 116 3126
rect 110 3121 111 3125
rect 115 3121 116 3125
rect 110 3120 116 3121
rect 1822 3125 1828 3126
rect 1822 3121 1823 3125
rect 1827 3121 1828 3125
rect 1862 3125 1863 3129
rect 1867 3125 1868 3129
rect 1862 3124 1868 3125
rect 3574 3129 3580 3130
rect 3574 3125 3575 3129
rect 3579 3125 3580 3129
rect 3574 3124 3580 3125
rect 1822 3120 1828 3121
rect 1862 3112 1868 3113
rect 110 3108 116 3109
rect 110 3104 111 3108
rect 115 3104 116 3108
rect 110 3103 116 3104
rect 1822 3108 1828 3109
rect 1822 3104 1823 3108
rect 1827 3104 1828 3108
rect 1862 3108 1863 3112
rect 1867 3108 1868 3112
rect 1862 3107 1868 3108
rect 3574 3112 3580 3113
rect 3574 3108 3575 3112
rect 3579 3108 3580 3112
rect 3574 3107 3580 3108
rect 1822 3103 1828 3104
rect 1894 3099 1900 3100
rect 470 3095 476 3096
rect 470 3091 471 3095
rect 475 3091 476 3095
rect 470 3090 476 3091
rect 558 3095 564 3096
rect 558 3091 559 3095
rect 563 3091 564 3095
rect 558 3090 564 3091
rect 646 3095 652 3096
rect 646 3091 647 3095
rect 651 3091 652 3095
rect 646 3090 652 3091
rect 742 3095 748 3096
rect 742 3091 743 3095
rect 747 3091 748 3095
rect 742 3090 748 3091
rect 854 3095 860 3096
rect 854 3091 855 3095
rect 859 3091 860 3095
rect 854 3090 860 3091
rect 974 3095 980 3096
rect 974 3091 975 3095
rect 979 3091 980 3095
rect 974 3090 980 3091
rect 1102 3095 1108 3096
rect 1102 3091 1103 3095
rect 1107 3091 1108 3095
rect 1102 3090 1108 3091
rect 1238 3095 1244 3096
rect 1238 3091 1239 3095
rect 1243 3091 1244 3095
rect 1238 3090 1244 3091
rect 1382 3095 1388 3096
rect 1382 3091 1383 3095
rect 1387 3091 1388 3095
rect 1382 3090 1388 3091
rect 1526 3095 1532 3096
rect 1526 3091 1527 3095
rect 1531 3091 1532 3095
rect 1894 3095 1895 3099
rect 1899 3095 1900 3099
rect 1894 3094 1900 3095
rect 2086 3099 2092 3100
rect 2086 3095 2087 3099
rect 2091 3095 2092 3099
rect 2086 3094 2092 3095
rect 2302 3099 2308 3100
rect 2302 3095 2303 3099
rect 2307 3095 2308 3099
rect 2302 3094 2308 3095
rect 2510 3099 2516 3100
rect 2510 3095 2511 3099
rect 2515 3095 2516 3099
rect 2510 3094 2516 3095
rect 2702 3099 2708 3100
rect 2702 3095 2703 3099
rect 2707 3095 2708 3099
rect 2702 3094 2708 3095
rect 2878 3099 2884 3100
rect 2878 3095 2879 3099
rect 2883 3095 2884 3099
rect 2878 3094 2884 3095
rect 3046 3099 3052 3100
rect 3046 3095 3047 3099
rect 3051 3095 3052 3099
rect 3046 3094 3052 3095
rect 3198 3099 3204 3100
rect 3198 3095 3199 3099
rect 3203 3095 3204 3099
rect 3198 3094 3204 3095
rect 3350 3099 3356 3100
rect 3350 3095 3351 3099
rect 3355 3095 3356 3099
rect 3350 3094 3356 3095
rect 3486 3099 3492 3100
rect 3486 3095 3487 3099
rect 3491 3095 3492 3099
rect 3486 3094 3492 3095
rect 1526 3090 1532 3091
rect 150 3053 156 3054
rect 150 3049 151 3053
rect 155 3049 156 3053
rect 150 3048 156 3049
rect 238 3053 244 3054
rect 238 3049 239 3053
rect 243 3049 244 3053
rect 238 3048 244 3049
rect 326 3053 332 3054
rect 326 3049 327 3053
rect 331 3049 332 3053
rect 326 3048 332 3049
rect 414 3053 420 3054
rect 414 3049 415 3053
rect 419 3049 420 3053
rect 414 3048 420 3049
rect 502 3053 508 3054
rect 502 3049 503 3053
rect 507 3049 508 3053
rect 502 3048 508 3049
rect 590 3053 596 3054
rect 590 3049 591 3053
rect 595 3049 596 3053
rect 590 3048 596 3049
rect 678 3053 684 3054
rect 678 3049 679 3053
rect 683 3049 684 3053
rect 678 3048 684 3049
rect 766 3053 772 3054
rect 766 3049 767 3053
rect 771 3049 772 3053
rect 766 3048 772 3049
rect 854 3053 860 3054
rect 854 3049 855 3053
rect 859 3049 860 3053
rect 854 3048 860 3049
rect 942 3053 948 3054
rect 942 3049 943 3053
rect 947 3049 948 3053
rect 942 3048 948 3049
rect 1030 3053 1036 3054
rect 1030 3049 1031 3053
rect 1035 3049 1036 3053
rect 1030 3048 1036 3049
rect 1118 3053 1124 3054
rect 1118 3049 1119 3053
rect 1123 3049 1124 3053
rect 1118 3048 1124 3049
rect 1206 3053 1212 3054
rect 1206 3049 1207 3053
rect 1211 3049 1212 3053
rect 1206 3048 1212 3049
rect 1294 3053 1300 3054
rect 1294 3049 1295 3053
rect 1299 3049 1300 3053
rect 1294 3048 1300 3049
rect 1382 3053 1388 3054
rect 1382 3049 1383 3053
rect 1387 3049 1388 3053
rect 1382 3048 1388 3049
rect 1470 3053 1476 3054
rect 1470 3049 1471 3053
rect 1475 3049 1476 3053
rect 1470 3048 1476 3049
rect 1558 3053 1564 3054
rect 1558 3049 1559 3053
rect 1563 3049 1564 3053
rect 1558 3048 1564 3049
rect 1646 3053 1652 3054
rect 1646 3049 1647 3053
rect 1651 3049 1652 3053
rect 1646 3048 1652 3049
rect 1734 3053 1740 3054
rect 1734 3049 1735 3053
rect 1739 3049 1740 3053
rect 1734 3048 1740 3049
rect 2254 3053 2260 3054
rect 2254 3049 2255 3053
rect 2259 3049 2260 3053
rect 2254 3048 2260 3049
rect 2422 3053 2428 3054
rect 2422 3049 2423 3053
rect 2427 3049 2428 3053
rect 2422 3048 2428 3049
rect 2590 3053 2596 3054
rect 2590 3049 2591 3053
rect 2595 3049 2596 3053
rect 2590 3048 2596 3049
rect 2750 3053 2756 3054
rect 2750 3049 2751 3053
rect 2755 3049 2756 3053
rect 2750 3048 2756 3049
rect 2918 3053 2924 3054
rect 2918 3049 2919 3053
rect 2923 3049 2924 3053
rect 2918 3048 2924 3049
rect 3086 3053 3092 3054
rect 3086 3049 3087 3053
rect 3091 3049 3092 3053
rect 3086 3048 3092 3049
rect 110 3040 116 3041
rect 110 3036 111 3040
rect 115 3036 116 3040
rect 110 3035 116 3036
rect 1822 3040 1828 3041
rect 1822 3036 1823 3040
rect 1827 3036 1828 3040
rect 1822 3035 1828 3036
rect 1862 3040 1868 3041
rect 1862 3036 1863 3040
rect 1867 3036 1868 3040
rect 1862 3035 1868 3036
rect 3574 3040 3580 3041
rect 3574 3036 3575 3040
rect 3579 3036 3580 3040
rect 3574 3035 3580 3036
rect 110 3023 116 3024
rect 110 3019 111 3023
rect 115 3019 116 3023
rect 110 3018 116 3019
rect 1822 3023 1828 3024
rect 1822 3019 1823 3023
rect 1827 3019 1828 3023
rect 1822 3018 1828 3019
rect 1862 3023 1868 3024
rect 1862 3019 1863 3023
rect 1867 3019 1868 3023
rect 1862 3018 1868 3019
rect 3574 3023 3580 3024
rect 3574 3019 3575 3023
rect 3579 3019 3580 3023
rect 3574 3018 3580 3019
rect 142 3013 148 3014
rect 142 3009 143 3013
rect 147 3009 148 3013
rect 142 3008 148 3009
rect 230 3013 236 3014
rect 230 3009 231 3013
rect 235 3009 236 3013
rect 230 3008 236 3009
rect 318 3013 324 3014
rect 318 3009 319 3013
rect 323 3009 324 3013
rect 318 3008 324 3009
rect 406 3013 412 3014
rect 406 3009 407 3013
rect 411 3009 412 3013
rect 406 3008 412 3009
rect 494 3013 500 3014
rect 494 3009 495 3013
rect 499 3009 500 3013
rect 494 3008 500 3009
rect 582 3013 588 3014
rect 582 3009 583 3013
rect 587 3009 588 3013
rect 582 3008 588 3009
rect 670 3013 676 3014
rect 670 3009 671 3013
rect 675 3009 676 3013
rect 670 3008 676 3009
rect 758 3013 764 3014
rect 758 3009 759 3013
rect 763 3009 764 3013
rect 758 3008 764 3009
rect 846 3013 852 3014
rect 846 3009 847 3013
rect 851 3009 852 3013
rect 846 3008 852 3009
rect 934 3013 940 3014
rect 934 3009 935 3013
rect 939 3009 940 3013
rect 934 3008 940 3009
rect 1022 3013 1028 3014
rect 1022 3009 1023 3013
rect 1027 3009 1028 3013
rect 1022 3008 1028 3009
rect 1110 3013 1116 3014
rect 1110 3009 1111 3013
rect 1115 3009 1116 3013
rect 1110 3008 1116 3009
rect 1198 3013 1204 3014
rect 1198 3009 1199 3013
rect 1203 3009 1204 3013
rect 1198 3008 1204 3009
rect 1286 3013 1292 3014
rect 1286 3009 1287 3013
rect 1291 3009 1292 3013
rect 1286 3008 1292 3009
rect 1374 3013 1380 3014
rect 1374 3009 1375 3013
rect 1379 3009 1380 3013
rect 1374 3008 1380 3009
rect 1462 3013 1468 3014
rect 1462 3009 1463 3013
rect 1467 3009 1468 3013
rect 1462 3008 1468 3009
rect 1550 3013 1556 3014
rect 1550 3009 1551 3013
rect 1555 3009 1556 3013
rect 1550 3008 1556 3009
rect 1638 3013 1644 3014
rect 1638 3009 1639 3013
rect 1643 3009 1644 3013
rect 1638 3008 1644 3009
rect 1726 3013 1732 3014
rect 1726 3009 1727 3013
rect 1731 3009 1732 3013
rect 1726 3008 1732 3009
rect 2246 3013 2252 3014
rect 2246 3009 2247 3013
rect 2251 3009 2252 3013
rect 2246 3008 2252 3009
rect 2414 3013 2420 3014
rect 2414 3009 2415 3013
rect 2419 3009 2420 3013
rect 2414 3008 2420 3009
rect 2582 3013 2588 3014
rect 2582 3009 2583 3013
rect 2587 3009 2588 3013
rect 2582 3008 2588 3009
rect 2742 3013 2748 3014
rect 2742 3009 2743 3013
rect 2747 3009 2748 3013
rect 2742 3008 2748 3009
rect 2910 3013 2916 3014
rect 2910 3009 2911 3013
rect 2915 3009 2916 3013
rect 2910 3008 2916 3009
rect 3078 3013 3084 3014
rect 3078 3009 3079 3013
rect 3083 3009 3084 3013
rect 3078 3008 3084 3009
rect 2238 2987 2244 2988
rect 1406 2983 1412 2984
rect 1406 2979 1407 2983
rect 1411 2979 1412 2983
rect 1406 2978 1412 2979
rect 1518 2983 1524 2984
rect 1518 2979 1519 2983
rect 1523 2979 1524 2983
rect 1518 2978 1524 2979
rect 1630 2983 1636 2984
rect 1630 2979 1631 2983
rect 1635 2979 1636 2983
rect 1630 2978 1636 2979
rect 1726 2983 1732 2984
rect 1726 2979 1727 2983
rect 1731 2979 1732 2983
rect 2238 2983 2239 2987
rect 2243 2983 2244 2987
rect 2238 2982 2244 2983
rect 2462 2987 2468 2988
rect 2462 2983 2463 2987
rect 2467 2983 2468 2987
rect 2462 2982 2468 2983
rect 2670 2987 2676 2988
rect 2670 2983 2671 2987
rect 2675 2983 2676 2987
rect 2670 2982 2676 2983
rect 2862 2987 2868 2988
rect 2862 2983 2863 2987
rect 2867 2983 2868 2987
rect 2862 2982 2868 2983
rect 3030 2987 3036 2988
rect 3030 2983 3031 2987
rect 3035 2983 3036 2987
rect 3030 2982 3036 2983
rect 3190 2987 3196 2988
rect 3190 2983 3191 2987
rect 3195 2983 3196 2987
rect 3190 2982 3196 2983
rect 3342 2987 3348 2988
rect 3342 2983 3343 2987
rect 3347 2983 3348 2987
rect 3342 2982 3348 2983
rect 3478 2987 3484 2988
rect 3478 2983 3479 2987
rect 3483 2983 3484 2987
rect 3478 2982 3484 2983
rect 1726 2978 1732 2979
rect 1862 2977 1868 2978
rect 110 2973 116 2974
rect 110 2969 111 2973
rect 115 2969 116 2973
rect 110 2968 116 2969
rect 1822 2973 1828 2974
rect 1822 2969 1823 2973
rect 1827 2969 1828 2973
rect 1862 2973 1863 2977
rect 1867 2973 1868 2977
rect 1862 2972 1868 2973
rect 3574 2977 3580 2978
rect 3574 2973 3575 2977
rect 3579 2973 3580 2977
rect 3574 2972 3580 2973
rect 1822 2968 1828 2969
rect 1862 2960 1868 2961
rect 110 2956 116 2957
rect 110 2952 111 2956
rect 115 2952 116 2956
rect 110 2951 116 2952
rect 1822 2956 1828 2957
rect 1822 2952 1823 2956
rect 1827 2952 1828 2956
rect 1862 2956 1863 2960
rect 1867 2956 1868 2960
rect 1862 2955 1868 2956
rect 3574 2960 3580 2961
rect 3574 2956 3575 2960
rect 3579 2956 3580 2960
rect 3574 2955 3580 2956
rect 1822 2951 1828 2952
rect 2246 2947 2252 2948
rect 1414 2943 1420 2944
rect 1414 2939 1415 2943
rect 1419 2939 1420 2943
rect 1414 2938 1420 2939
rect 1526 2943 1532 2944
rect 1526 2939 1527 2943
rect 1531 2939 1532 2943
rect 1526 2938 1532 2939
rect 1638 2943 1644 2944
rect 1638 2939 1639 2943
rect 1643 2939 1644 2943
rect 1638 2938 1644 2939
rect 1734 2943 1740 2944
rect 1734 2939 1735 2943
rect 1739 2939 1740 2943
rect 2246 2943 2247 2947
rect 2251 2943 2252 2947
rect 2246 2942 2252 2943
rect 2470 2947 2476 2948
rect 2470 2943 2471 2947
rect 2475 2943 2476 2947
rect 2470 2942 2476 2943
rect 2678 2947 2684 2948
rect 2678 2943 2679 2947
rect 2683 2943 2684 2947
rect 2678 2942 2684 2943
rect 2870 2947 2876 2948
rect 2870 2943 2871 2947
rect 2875 2943 2876 2947
rect 2870 2942 2876 2943
rect 3038 2947 3044 2948
rect 3038 2943 3039 2947
rect 3043 2943 3044 2947
rect 3038 2942 3044 2943
rect 3198 2947 3204 2948
rect 3198 2943 3199 2947
rect 3203 2943 3204 2947
rect 3198 2942 3204 2943
rect 3350 2947 3356 2948
rect 3350 2943 3351 2947
rect 3355 2943 3356 2947
rect 3350 2942 3356 2943
rect 3486 2947 3492 2948
rect 3486 2943 3487 2947
rect 3491 2943 3492 2947
rect 3486 2942 3492 2943
rect 1734 2938 1740 2939
rect 1358 2909 1364 2910
rect 1358 2905 1359 2909
rect 1363 2905 1364 2909
rect 1358 2904 1364 2905
rect 1470 2909 1476 2910
rect 1470 2905 1471 2909
rect 1475 2905 1476 2909
rect 1470 2904 1476 2905
rect 1582 2909 1588 2910
rect 1582 2905 1583 2909
rect 1587 2905 1588 2909
rect 1582 2904 1588 2905
rect 1702 2909 1708 2910
rect 1702 2905 1703 2909
rect 1707 2905 1708 2909
rect 1702 2904 1708 2905
rect 2238 2897 2244 2898
rect 110 2896 116 2897
rect 110 2892 111 2896
rect 115 2892 116 2896
rect 110 2891 116 2892
rect 1822 2896 1828 2897
rect 1822 2892 1823 2896
rect 1827 2892 1828 2896
rect 2238 2893 2239 2897
rect 2243 2893 2244 2897
rect 2238 2892 2244 2893
rect 2462 2897 2468 2898
rect 2462 2893 2463 2897
rect 2467 2893 2468 2897
rect 2462 2892 2468 2893
rect 2670 2897 2676 2898
rect 2670 2893 2671 2897
rect 2675 2893 2676 2897
rect 2670 2892 2676 2893
rect 2854 2897 2860 2898
rect 2854 2893 2855 2897
rect 2859 2893 2860 2897
rect 2854 2892 2860 2893
rect 3022 2897 3028 2898
rect 3022 2893 3023 2897
rect 3027 2893 3028 2897
rect 3022 2892 3028 2893
rect 3182 2897 3188 2898
rect 3182 2893 3183 2897
rect 3187 2893 3188 2897
rect 3182 2892 3188 2893
rect 3334 2897 3340 2898
rect 3334 2893 3335 2897
rect 3339 2893 3340 2897
rect 3334 2892 3340 2893
rect 3486 2897 3492 2898
rect 3486 2893 3487 2897
rect 3491 2893 3492 2897
rect 3486 2892 3492 2893
rect 1822 2891 1828 2892
rect 1862 2884 1868 2885
rect 1862 2880 1863 2884
rect 1867 2880 1868 2884
rect 110 2879 116 2880
rect 110 2875 111 2879
rect 115 2875 116 2879
rect 110 2874 116 2875
rect 1822 2879 1828 2880
rect 1862 2879 1868 2880
rect 3574 2884 3580 2885
rect 3574 2880 3575 2884
rect 3579 2880 3580 2884
rect 3574 2879 3580 2880
rect 1822 2875 1823 2879
rect 1827 2875 1828 2879
rect 1822 2874 1828 2875
rect 1350 2869 1356 2870
rect 1350 2865 1351 2869
rect 1355 2865 1356 2869
rect 1350 2864 1356 2865
rect 1462 2869 1468 2870
rect 1462 2865 1463 2869
rect 1467 2865 1468 2869
rect 1462 2864 1468 2865
rect 1574 2869 1580 2870
rect 1574 2865 1575 2869
rect 1579 2865 1580 2869
rect 1574 2864 1580 2865
rect 1694 2869 1700 2870
rect 1694 2865 1695 2869
rect 1699 2865 1700 2869
rect 1694 2864 1700 2865
rect 1862 2867 1868 2868
rect 1862 2863 1863 2867
rect 1867 2863 1868 2867
rect 1862 2862 1868 2863
rect 3574 2867 3580 2868
rect 3574 2863 3575 2867
rect 3579 2863 3580 2867
rect 3574 2862 3580 2863
rect 2230 2857 2236 2858
rect 2230 2853 2231 2857
rect 2235 2853 2236 2857
rect 2230 2852 2236 2853
rect 2454 2857 2460 2858
rect 2454 2853 2455 2857
rect 2459 2853 2460 2857
rect 2454 2852 2460 2853
rect 2662 2857 2668 2858
rect 2662 2853 2663 2857
rect 2667 2853 2668 2857
rect 2662 2852 2668 2853
rect 2846 2857 2852 2858
rect 2846 2853 2847 2857
rect 2851 2853 2852 2857
rect 2846 2852 2852 2853
rect 3014 2857 3020 2858
rect 3014 2853 3015 2857
rect 3019 2853 3020 2857
rect 3014 2852 3020 2853
rect 3174 2857 3180 2858
rect 3174 2853 3175 2857
rect 3179 2853 3180 2857
rect 3174 2852 3180 2853
rect 3326 2857 3332 2858
rect 3326 2853 3327 2857
rect 3331 2853 3332 2857
rect 3326 2852 3332 2853
rect 3478 2857 3484 2858
rect 3478 2853 3479 2857
rect 3483 2853 3484 2857
rect 3478 2852 3484 2853
rect 134 2843 140 2844
rect 134 2839 135 2843
rect 139 2839 140 2843
rect 134 2838 140 2839
rect 222 2843 228 2844
rect 222 2839 223 2843
rect 227 2839 228 2843
rect 222 2838 228 2839
rect 310 2843 316 2844
rect 310 2839 311 2843
rect 315 2839 316 2843
rect 310 2838 316 2839
rect 398 2843 404 2844
rect 398 2839 399 2843
rect 403 2839 404 2843
rect 398 2838 404 2839
rect 486 2843 492 2844
rect 486 2839 487 2843
rect 491 2839 492 2843
rect 486 2838 492 2839
rect 598 2843 604 2844
rect 598 2839 599 2843
rect 603 2839 604 2843
rect 598 2838 604 2839
rect 726 2843 732 2844
rect 726 2839 727 2843
rect 731 2839 732 2843
rect 726 2838 732 2839
rect 862 2843 868 2844
rect 862 2839 863 2843
rect 867 2839 868 2843
rect 862 2838 868 2839
rect 998 2843 1004 2844
rect 998 2839 999 2843
rect 1003 2839 1004 2843
rect 998 2838 1004 2839
rect 1134 2843 1140 2844
rect 1134 2839 1135 2843
rect 1139 2839 1140 2843
rect 1134 2838 1140 2839
rect 1262 2843 1268 2844
rect 1262 2839 1263 2843
rect 1267 2839 1268 2843
rect 1262 2838 1268 2839
rect 1382 2843 1388 2844
rect 1382 2839 1383 2843
rect 1387 2839 1388 2843
rect 1382 2838 1388 2839
rect 1502 2843 1508 2844
rect 1502 2839 1503 2843
rect 1507 2839 1508 2843
rect 1502 2838 1508 2839
rect 1622 2843 1628 2844
rect 1622 2839 1623 2843
rect 1627 2839 1628 2843
rect 1622 2838 1628 2839
rect 1726 2843 1732 2844
rect 1726 2839 1727 2843
rect 1731 2839 1732 2843
rect 1726 2838 1732 2839
rect 110 2833 116 2834
rect 110 2829 111 2833
rect 115 2829 116 2833
rect 110 2828 116 2829
rect 1822 2833 1828 2834
rect 1822 2829 1823 2833
rect 1827 2829 1828 2833
rect 1822 2828 1828 2829
rect 1894 2831 1900 2832
rect 1894 2827 1895 2831
rect 1899 2827 1900 2831
rect 1894 2826 1900 2827
rect 1982 2831 1988 2832
rect 1982 2827 1983 2831
rect 1987 2827 1988 2831
rect 1982 2826 1988 2827
rect 2070 2831 2076 2832
rect 2070 2827 2071 2831
rect 2075 2827 2076 2831
rect 2070 2826 2076 2827
rect 2158 2831 2164 2832
rect 2158 2827 2159 2831
rect 2163 2827 2164 2831
rect 2158 2826 2164 2827
rect 2246 2831 2252 2832
rect 2246 2827 2247 2831
rect 2251 2827 2252 2831
rect 2246 2826 2252 2827
rect 2334 2831 2340 2832
rect 2334 2827 2335 2831
rect 2339 2827 2340 2831
rect 2334 2826 2340 2827
rect 2422 2831 2428 2832
rect 2422 2827 2423 2831
rect 2427 2827 2428 2831
rect 2422 2826 2428 2827
rect 2510 2831 2516 2832
rect 2510 2827 2511 2831
rect 2515 2827 2516 2831
rect 2510 2826 2516 2827
rect 2598 2831 2604 2832
rect 2598 2827 2599 2831
rect 2603 2827 2604 2831
rect 2598 2826 2604 2827
rect 2686 2831 2692 2832
rect 2686 2827 2687 2831
rect 2691 2827 2692 2831
rect 2686 2826 2692 2827
rect 2790 2831 2796 2832
rect 2790 2827 2791 2831
rect 2795 2827 2796 2831
rect 2790 2826 2796 2827
rect 2902 2831 2908 2832
rect 2902 2827 2903 2831
rect 2907 2827 2908 2831
rect 2902 2826 2908 2827
rect 3030 2831 3036 2832
rect 3030 2827 3031 2831
rect 3035 2827 3036 2831
rect 3030 2826 3036 2827
rect 3174 2831 3180 2832
rect 3174 2827 3175 2831
rect 3179 2827 3180 2831
rect 3174 2826 3180 2827
rect 3326 2831 3332 2832
rect 3326 2827 3327 2831
rect 3331 2827 3332 2831
rect 3326 2826 3332 2827
rect 3478 2831 3484 2832
rect 3478 2827 3479 2831
rect 3483 2827 3484 2831
rect 3478 2826 3484 2827
rect 1862 2821 1868 2822
rect 1862 2817 1863 2821
rect 1867 2817 1868 2821
rect 110 2816 116 2817
rect 110 2812 111 2816
rect 115 2812 116 2816
rect 110 2811 116 2812
rect 1822 2816 1828 2817
rect 1862 2816 1868 2817
rect 3574 2821 3580 2822
rect 3574 2817 3575 2821
rect 3579 2817 3580 2821
rect 3574 2816 3580 2817
rect 1822 2812 1823 2816
rect 1827 2812 1828 2816
rect 1822 2811 1828 2812
rect 1862 2804 1868 2805
rect 142 2803 148 2804
rect 142 2799 143 2803
rect 147 2799 148 2803
rect 142 2798 148 2799
rect 230 2803 236 2804
rect 230 2799 231 2803
rect 235 2799 236 2803
rect 230 2798 236 2799
rect 318 2803 324 2804
rect 318 2799 319 2803
rect 323 2799 324 2803
rect 318 2798 324 2799
rect 406 2803 412 2804
rect 406 2799 407 2803
rect 411 2799 412 2803
rect 406 2798 412 2799
rect 494 2803 500 2804
rect 494 2799 495 2803
rect 499 2799 500 2803
rect 494 2798 500 2799
rect 606 2803 612 2804
rect 606 2799 607 2803
rect 611 2799 612 2803
rect 606 2798 612 2799
rect 734 2803 740 2804
rect 734 2799 735 2803
rect 739 2799 740 2803
rect 734 2798 740 2799
rect 870 2803 876 2804
rect 870 2799 871 2803
rect 875 2799 876 2803
rect 870 2798 876 2799
rect 1006 2803 1012 2804
rect 1006 2799 1007 2803
rect 1011 2799 1012 2803
rect 1006 2798 1012 2799
rect 1142 2803 1148 2804
rect 1142 2799 1143 2803
rect 1147 2799 1148 2803
rect 1142 2798 1148 2799
rect 1270 2803 1276 2804
rect 1270 2799 1271 2803
rect 1275 2799 1276 2803
rect 1270 2798 1276 2799
rect 1390 2803 1396 2804
rect 1390 2799 1391 2803
rect 1395 2799 1396 2803
rect 1390 2798 1396 2799
rect 1510 2803 1516 2804
rect 1510 2799 1511 2803
rect 1515 2799 1516 2803
rect 1510 2798 1516 2799
rect 1630 2803 1636 2804
rect 1630 2799 1631 2803
rect 1635 2799 1636 2803
rect 1630 2798 1636 2799
rect 1734 2803 1740 2804
rect 1734 2799 1735 2803
rect 1739 2799 1740 2803
rect 1862 2800 1863 2804
rect 1867 2800 1868 2804
rect 1862 2799 1868 2800
rect 3574 2804 3580 2805
rect 3574 2800 3575 2804
rect 3579 2800 3580 2804
rect 3574 2799 3580 2800
rect 1734 2798 1740 2799
rect 1902 2791 1908 2792
rect 1902 2787 1903 2791
rect 1907 2787 1908 2791
rect 1902 2786 1908 2787
rect 1990 2791 1996 2792
rect 1990 2787 1991 2791
rect 1995 2787 1996 2791
rect 1990 2786 1996 2787
rect 2078 2791 2084 2792
rect 2078 2787 2079 2791
rect 2083 2787 2084 2791
rect 2078 2786 2084 2787
rect 2166 2791 2172 2792
rect 2166 2787 2167 2791
rect 2171 2787 2172 2791
rect 2166 2786 2172 2787
rect 2254 2791 2260 2792
rect 2254 2787 2255 2791
rect 2259 2787 2260 2791
rect 2254 2786 2260 2787
rect 2342 2791 2348 2792
rect 2342 2787 2343 2791
rect 2347 2787 2348 2791
rect 2342 2786 2348 2787
rect 2430 2791 2436 2792
rect 2430 2787 2431 2791
rect 2435 2787 2436 2791
rect 2430 2786 2436 2787
rect 2518 2791 2524 2792
rect 2518 2787 2519 2791
rect 2523 2787 2524 2791
rect 2518 2786 2524 2787
rect 2606 2791 2612 2792
rect 2606 2787 2607 2791
rect 2611 2787 2612 2791
rect 2606 2786 2612 2787
rect 2694 2791 2700 2792
rect 2694 2787 2695 2791
rect 2699 2787 2700 2791
rect 2694 2786 2700 2787
rect 2798 2791 2804 2792
rect 2798 2787 2799 2791
rect 2803 2787 2804 2791
rect 2798 2786 2804 2787
rect 2910 2791 2916 2792
rect 2910 2787 2911 2791
rect 2915 2787 2916 2791
rect 2910 2786 2916 2787
rect 3038 2791 3044 2792
rect 3038 2787 3039 2791
rect 3043 2787 3044 2791
rect 3038 2786 3044 2787
rect 3182 2791 3188 2792
rect 3182 2787 3183 2791
rect 3187 2787 3188 2791
rect 3182 2786 3188 2787
rect 3334 2791 3340 2792
rect 3334 2787 3335 2791
rect 3339 2787 3340 2791
rect 3334 2786 3340 2787
rect 3486 2791 3492 2792
rect 3486 2787 3487 2791
rect 3491 2787 3492 2791
rect 3486 2786 3492 2787
rect 190 2769 196 2770
rect 190 2765 191 2769
rect 195 2765 196 2769
rect 190 2764 196 2765
rect 294 2769 300 2770
rect 294 2765 295 2769
rect 299 2765 300 2769
rect 294 2764 300 2765
rect 414 2769 420 2770
rect 414 2765 415 2769
rect 419 2765 420 2769
rect 414 2764 420 2765
rect 550 2769 556 2770
rect 550 2765 551 2769
rect 555 2765 556 2769
rect 550 2764 556 2765
rect 686 2769 692 2770
rect 686 2765 687 2769
rect 691 2765 692 2769
rect 686 2764 692 2765
rect 822 2769 828 2770
rect 822 2765 823 2769
rect 827 2765 828 2769
rect 822 2764 828 2765
rect 958 2769 964 2770
rect 958 2765 959 2769
rect 963 2765 964 2769
rect 958 2764 964 2765
rect 1086 2769 1092 2770
rect 1086 2765 1087 2769
rect 1091 2765 1092 2769
rect 1086 2764 1092 2765
rect 1206 2769 1212 2770
rect 1206 2765 1207 2769
rect 1211 2765 1212 2769
rect 1206 2764 1212 2765
rect 1318 2769 1324 2770
rect 1318 2765 1319 2769
rect 1323 2765 1324 2769
rect 1318 2764 1324 2765
rect 1430 2769 1436 2770
rect 1430 2765 1431 2769
rect 1435 2765 1436 2769
rect 1430 2764 1436 2765
rect 1534 2769 1540 2770
rect 1534 2765 1535 2769
rect 1539 2765 1540 2769
rect 1534 2764 1540 2765
rect 1646 2769 1652 2770
rect 1646 2765 1647 2769
rect 1651 2765 1652 2769
rect 1646 2764 1652 2765
rect 1734 2769 1740 2770
rect 1734 2765 1735 2769
rect 1739 2765 1740 2769
rect 1734 2764 1740 2765
rect 110 2756 116 2757
rect 110 2752 111 2756
rect 115 2752 116 2756
rect 110 2751 116 2752
rect 1822 2756 1828 2757
rect 1822 2752 1823 2756
rect 1827 2752 1828 2756
rect 1822 2751 1828 2752
rect 2046 2745 2052 2746
rect 2046 2741 2047 2745
rect 2051 2741 2052 2745
rect 2046 2740 2052 2741
rect 2166 2745 2172 2746
rect 2166 2741 2167 2745
rect 2171 2741 2172 2745
rect 2166 2740 2172 2741
rect 2294 2745 2300 2746
rect 2294 2741 2295 2745
rect 2299 2741 2300 2745
rect 2294 2740 2300 2741
rect 2446 2745 2452 2746
rect 2446 2741 2447 2745
rect 2451 2741 2452 2745
rect 2446 2740 2452 2741
rect 2622 2745 2628 2746
rect 2622 2741 2623 2745
rect 2627 2741 2628 2745
rect 2622 2740 2628 2741
rect 2822 2745 2828 2746
rect 2822 2741 2823 2745
rect 2827 2741 2828 2745
rect 2822 2740 2828 2741
rect 3038 2745 3044 2746
rect 3038 2741 3039 2745
rect 3043 2741 3044 2745
rect 3038 2740 3044 2741
rect 3270 2745 3276 2746
rect 3270 2741 3271 2745
rect 3275 2741 3276 2745
rect 3270 2740 3276 2741
rect 3486 2745 3492 2746
rect 3486 2741 3487 2745
rect 3491 2741 3492 2745
rect 3486 2740 3492 2741
rect 110 2739 116 2740
rect 110 2735 111 2739
rect 115 2735 116 2739
rect 110 2734 116 2735
rect 1822 2739 1828 2740
rect 1822 2735 1823 2739
rect 1827 2735 1828 2739
rect 1822 2734 1828 2735
rect 1862 2732 1868 2733
rect 182 2729 188 2730
rect 182 2725 183 2729
rect 187 2725 188 2729
rect 182 2724 188 2725
rect 286 2729 292 2730
rect 286 2725 287 2729
rect 291 2725 292 2729
rect 286 2724 292 2725
rect 406 2729 412 2730
rect 406 2725 407 2729
rect 411 2725 412 2729
rect 406 2724 412 2725
rect 542 2729 548 2730
rect 542 2725 543 2729
rect 547 2725 548 2729
rect 542 2724 548 2725
rect 678 2729 684 2730
rect 678 2725 679 2729
rect 683 2725 684 2729
rect 678 2724 684 2725
rect 814 2729 820 2730
rect 814 2725 815 2729
rect 819 2725 820 2729
rect 814 2724 820 2725
rect 950 2729 956 2730
rect 950 2725 951 2729
rect 955 2725 956 2729
rect 950 2724 956 2725
rect 1078 2729 1084 2730
rect 1078 2725 1079 2729
rect 1083 2725 1084 2729
rect 1078 2724 1084 2725
rect 1198 2729 1204 2730
rect 1198 2725 1199 2729
rect 1203 2725 1204 2729
rect 1198 2724 1204 2725
rect 1310 2729 1316 2730
rect 1310 2725 1311 2729
rect 1315 2725 1316 2729
rect 1310 2724 1316 2725
rect 1422 2729 1428 2730
rect 1422 2725 1423 2729
rect 1427 2725 1428 2729
rect 1422 2724 1428 2725
rect 1526 2729 1532 2730
rect 1526 2725 1527 2729
rect 1531 2725 1532 2729
rect 1526 2724 1532 2725
rect 1638 2729 1644 2730
rect 1638 2725 1639 2729
rect 1643 2725 1644 2729
rect 1638 2724 1644 2725
rect 1726 2729 1732 2730
rect 1726 2725 1727 2729
rect 1731 2725 1732 2729
rect 1862 2728 1863 2732
rect 1867 2728 1868 2732
rect 1862 2727 1868 2728
rect 3574 2732 3580 2733
rect 3574 2728 3575 2732
rect 3579 2728 3580 2732
rect 3574 2727 3580 2728
rect 1726 2724 1732 2725
rect 1862 2715 1868 2716
rect 1862 2711 1863 2715
rect 1867 2711 1868 2715
rect 1862 2710 1868 2711
rect 3574 2715 3580 2716
rect 3574 2711 3575 2715
rect 3579 2711 3580 2715
rect 3574 2710 3580 2711
rect 2038 2705 2044 2706
rect 2038 2701 2039 2705
rect 2043 2701 2044 2705
rect 2038 2700 2044 2701
rect 2158 2705 2164 2706
rect 2158 2701 2159 2705
rect 2163 2701 2164 2705
rect 2158 2700 2164 2701
rect 2286 2705 2292 2706
rect 2286 2701 2287 2705
rect 2291 2701 2292 2705
rect 2286 2700 2292 2701
rect 2438 2705 2444 2706
rect 2438 2701 2439 2705
rect 2443 2701 2444 2705
rect 2438 2700 2444 2701
rect 2614 2705 2620 2706
rect 2614 2701 2615 2705
rect 2619 2701 2620 2705
rect 2614 2700 2620 2701
rect 2814 2705 2820 2706
rect 2814 2701 2815 2705
rect 2819 2701 2820 2705
rect 2814 2700 2820 2701
rect 3030 2705 3036 2706
rect 3030 2701 3031 2705
rect 3035 2701 3036 2705
rect 3030 2700 3036 2701
rect 3262 2705 3268 2706
rect 3262 2701 3263 2705
rect 3267 2701 3268 2705
rect 3262 2700 3268 2701
rect 3478 2705 3484 2706
rect 3478 2701 3479 2705
rect 3483 2701 3484 2705
rect 3478 2700 3484 2701
rect 166 2699 172 2700
rect 166 2695 167 2699
rect 171 2695 172 2699
rect 166 2694 172 2695
rect 278 2699 284 2700
rect 278 2695 279 2699
rect 283 2695 284 2699
rect 278 2694 284 2695
rect 390 2699 396 2700
rect 390 2695 391 2699
rect 395 2695 396 2699
rect 390 2694 396 2695
rect 502 2699 508 2700
rect 502 2695 503 2699
rect 507 2695 508 2699
rect 502 2694 508 2695
rect 614 2699 620 2700
rect 614 2695 615 2699
rect 619 2695 620 2699
rect 614 2694 620 2695
rect 110 2689 116 2690
rect 110 2685 111 2689
rect 115 2685 116 2689
rect 110 2684 116 2685
rect 1822 2689 1828 2690
rect 1822 2685 1823 2689
rect 1827 2685 1828 2689
rect 1822 2684 1828 2685
rect 1942 2683 1948 2684
rect 1942 2679 1943 2683
rect 1947 2679 1948 2683
rect 1942 2678 1948 2679
rect 2054 2683 2060 2684
rect 2054 2679 2055 2683
rect 2059 2679 2060 2683
rect 2054 2678 2060 2679
rect 2166 2683 2172 2684
rect 2166 2679 2167 2683
rect 2171 2679 2172 2683
rect 2166 2678 2172 2679
rect 2286 2683 2292 2684
rect 2286 2679 2287 2683
rect 2291 2679 2292 2683
rect 2286 2678 2292 2679
rect 2406 2683 2412 2684
rect 2406 2679 2407 2683
rect 2411 2679 2412 2683
rect 2406 2678 2412 2679
rect 2518 2683 2524 2684
rect 2518 2679 2519 2683
rect 2523 2679 2524 2683
rect 2518 2678 2524 2679
rect 2630 2683 2636 2684
rect 2630 2679 2631 2683
rect 2635 2679 2636 2683
rect 2630 2678 2636 2679
rect 2734 2683 2740 2684
rect 2734 2679 2735 2683
rect 2739 2679 2740 2683
rect 2734 2678 2740 2679
rect 2846 2683 2852 2684
rect 2846 2679 2847 2683
rect 2851 2679 2852 2683
rect 2846 2678 2852 2679
rect 2958 2683 2964 2684
rect 2958 2679 2959 2683
rect 2963 2679 2964 2683
rect 2958 2678 2964 2679
rect 3070 2683 3076 2684
rect 3070 2679 3071 2683
rect 3075 2679 3076 2683
rect 3070 2678 3076 2679
rect 1862 2673 1868 2674
rect 110 2672 116 2673
rect 110 2668 111 2672
rect 115 2668 116 2672
rect 110 2667 116 2668
rect 1822 2672 1828 2673
rect 1822 2668 1823 2672
rect 1827 2668 1828 2672
rect 1862 2669 1863 2673
rect 1867 2669 1868 2673
rect 1862 2668 1868 2669
rect 3574 2673 3580 2674
rect 3574 2669 3575 2673
rect 3579 2669 3580 2673
rect 3574 2668 3580 2669
rect 1822 2667 1828 2668
rect 174 2659 180 2660
rect 174 2655 175 2659
rect 179 2655 180 2659
rect 174 2654 180 2655
rect 286 2659 292 2660
rect 286 2655 287 2659
rect 291 2655 292 2659
rect 286 2654 292 2655
rect 398 2659 404 2660
rect 398 2655 399 2659
rect 403 2655 404 2659
rect 398 2654 404 2655
rect 510 2659 516 2660
rect 510 2655 511 2659
rect 515 2655 516 2659
rect 510 2654 516 2655
rect 622 2659 628 2660
rect 622 2655 623 2659
rect 627 2655 628 2659
rect 622 2654 628 2655
rect 1862 2656 1868 2657
rect 1862 2652 1863 2656
rect 1867 2652 1868 2656
rect 1862 2651 1868 2652
rect 3574 2656 3580 2657
rect 3574 2652 3575 2656
rect 3579 2652 3580 2656
rect 3574 2651 3580 2652
rect 1950 2643 1956 2644
rect 1950 2639 1951 2643
rect 1955 2639 1956 2643
rect 1950 2638 1956 2639
rect 2062 2643 2068 2644
rect 2062 2639 2063 2643
rect 2067 2639 2068 2643
rect 2062 2638 2068 2639
rect 2174 2643 2180 2644
rect 2174 2639 2175 2643
rect 2179 2639 2180 2643
rect 2174 2638 2180 2639
rect 2294 2643 2300 2644
rect 2294 2639 2295 2643
rect 2299 2639 2300 2643
rect 2294 2638 2300 2639
rect 2414 2643 2420 2644
rect 2414 2639 2415 2643
rect 2419 2639 2420 2643
rect 2414 2638 2420 2639
rect 2526 2643 2532 2644
rect 2526 2639 2527 2643
rect 2531 2639 2532 2643
rect 2526 2638 2532 2639
rect 2638 2643 2644 2644
rect 2638 2639 2639 2643
rect 2643 2639 2644 2643
rect 2638 2638 2644 2639
rect 2742 2643 2748 2644
rect 2742 2639 2743 2643
rect 2747 2639 2748 2643
rect 2742 2638 2748 2639
rect 2854 2643 2860 2644
rect 2854 2639 2855 2643
rect 2859 2639 2860 2643
rect 2854 2638 2860 2639
rect 2966 2643 2972 2644
rect 2966 2639 2967 2643
rect 2971 2639 2972 2643
rect 2966 2638 2972 2639
rect 3078 2643 3084 2644
rect 3078 2639 3079 2643
rect 3083 2639 3084 2643
rect 3078 2638 3084 2639
rect 222 2609 228 2610
rect 222 2605 223 2609
rect 227 2605 228 2609
rect 222 2604 228 2605
rect 350 2609 356 2610
rect 350 2605 351 2609
rect 355 2605 356 2609
rect 350 2604 356 2605
rect 494 2609 500 2610
rect 494 2605 495 2609
rect 499 2605 500 2609
rect 494 2604 500 2605
rect 662 2609 668 2610
rect 662 2605 663 2609
rect 667 2605 668 2609
rect 662 2604 668 2605
rect 838 2609 844 2610
rect 838 2605 839 2609
rect 843 2605 844 2609
rect 838 2604 844 2605
rect 1022 2609 1028 2610
rect 1022 2605 1023 2609
rect 1027 2605 1028 2609
rect 1022 2604 1028 2605
rect 1214 2609 1220 2610
rect 1214 2605 1215 2609
rect 1219 2605 1220 2609
rect 1214 2604 1220 2605
rect 1406 2609 1412 2610
rect 1406 2605 1407 2609
rect 1411 2605 1412 2609
rect 1406 2604 1412 2605
rect 1606 2609 1612 2610
rect 1606 2605 1607 2609
rect 1611 2605 1612 2609
rect 1606 2604 1612 2605
rect 1894 2605 1900 2606
rect 1894 2601 1895 2605
rect 1899 2601 1900 2605
rect 1894 2600 1900 2601
rect 2070 2605 2076 2606
rect 2070 2601 2071 2605
rect 2075 2601 2076 2605
rect 2070 2600 2076 2601
rect 2262 2605 2268 2606
rect 2262 2601 2263 2605
rect 2267 2601 2268 2605
rect 2262 2600 2268 2601
rect 2462 2605 2468 2606
rect 2462 2601 2463 2605
rect 2467 2601 2468 2605
rect 2462 2600 2468 2601
rect 2662 2605 2668 2606
rect 2662 2601 2663 2605
rect 2667 2601 2668 2605
rect 2662 2600 2668 2601
rect 2870 2605 2876 2606
rect 2870 2601 2871 2605
rect 2875 2601 2876 2605
rect 2870 2600 2876 2601
rect 3078 2605 3084 2606
rect 3078 2601 3079 2605
rect 3083 2601 3084 2605
rect 3078 2600 3084 2601
rect 3294 2605 3300 2606
rect 3294 2601 3295 2605
rect 3299 2601 3300 2605
rect 3294 2600 3300 2601
rect 3486 2605 3492 2606
rect 3486 2601 3487 2605
rect 3491 2601 3492 2605
rect 3486 2600 3492 2601
rect 110 2596 116 2597
rect 110 2592 111 2596
rect 115 2592 116 2596
rect 110 2591 116 2592
rect 1822 2596 1828 2597
rect 1822 2592 1823 2596
rect 1827 2592 1828 2596
rect 1822 2591 1828 2592
rect 1862 2592 1868 2593
rect 1862 2588 1863 2592
rect 1867 2588 1868 2592
rect 1862 2587 1868 2588
rect 3574 2592 3580 2593
rect 3574 2588 3575 2592
rect 3579 2588 3580 2592
rect 3574 2587 3580 2588
rect 110 2579 116 2580
rect 110 2575 111 2579
rect 115 2575 116 2579
rect 110 2574 116 2575
rect 1822 2579 1828 2580
rect 1822 2575 1823 2579
rect 1827 2575 1828 2579
rect 1822 2574 1828 2575
rect 1862 2575 1868 2576
rect 1862 2571 1863 2575
rect 1867 2571 1868 2575
rect 1862 2570 1868 2571
rect 3574 2575 3580 2576
rect 3574 2571 3575 2575
rect 3579 2571 3580 2575
rect 3574 2570 3580 2571
rect 214 2569 220 2570
rect 214 2565 215 2569
rect 219 2565 220 2569
rect 214 2564 220 2565
rect 342 2569 348 2570
rect 342 2565 343 2569
rect 347 2565 348 2569
rect 342 2564 348 2565
rect 486 2569 492 2570
rect 486 2565 487 2569
rect 491 2565 492 2569
rect 486 2564 492 2565
rect 654 2569 660 2570
rect 654 2565 655 2569
rect 659 2565 660 2569
rect 654 2564 660 2565
rect 830 2569 836 2570
rect 830 2565 831 2569
rect 835 2565 836 2569
rect 830 2564 836 2565
rect 1014 2569 1020 2570
rect 1014 2565 1015 2569
rect 1019 2565 1020 2569
rect 1014 2564 1020 2565
rect 1206 2569 1212 2570
rect 1206 2565 1207 2569
rect 1211 2565 1212 2569
rect 1206 2564 1212 2565
rect 1398 2569 1404 2570
rect 1398 2565 1399 2569
rect 1403 2565 1404 2569
rect 1398 2564 1404 2565
rect 1598 2569 1604 2570
rect 1598 2565 1599 2569
rect 1603 2565 1604 2569
rect 1598 2564 1604 2565
rect 1886 2565 1892 2566
rect 1886 2561 1887 2565
rect 1891 2561 1892 2565
rect 1886 2560 1892 2561
rect 2062 2565 2068 2566
rect 2062 2561 2063 2565
rect 2067 2561 2068 2565
rect 2062 2560 2068 2561
rect 2254 2565 2260 2566
rect 2254 2561 2255 2565
rect 2259 2561 2260 2565
rect 2254 2560 2260 2561
rect 2454 2565 2460 2566
rect 2454 2561 2455 2565
rect 2459 2561 2460 2565
rect 2454 2560 2460 2561
rect 2654 2565 2660 2566
rect 2654 2561 2655 2565
rect 2659 2561 2660 2565
rect 2654 2560 2660 2561
rect 2862 2565 2868 2566
rect 2862 2561 2863 2565
rect 2867 2561 2868 2565
rect 2862 2560 2868 2561
rect 3070 2565 3076 2566
rect 3070 2561 3071 2565
rect 3075 2561 3076 2565
rect 3070 2560 3076 2561
rect 3286 2565 3292 2566
rect 3286 2561 3287 2565
rect 3291 2561 3292 2565
rect 3286 2560 3292 2561
rect 3478 2565 3484 2566
rect 3478 2561 3479 2565
rect 3483 2561 3484 2565
rect 3478 2560 3484 2561
rect 270 2547 276 2548
rect 270 2543 271 2547
rect 275 2543 276 2547
rect 270 2542 276 2543
rect 470 2547 476 2548
rect 470 2543 471 2547
rect 475 2543 476 2547
rect 470 2542 476 2543
rect 670 2547 676 2548
rect 670 2543 671 2547
rect 675 2543 676 2547
rect 670 2542 676 2543
rect 854 2547 860 2548
rect 854 2543 855 2547
rect 859 2543 860 2547
rect 854 2542 860 2543
rect 1022 2547 1028 2548
rect 1022 2543 1023 2547
rect 1027 2543 1028 2547
rect 1022 2542 1028 2543
rect 1174 2547 1180 2548
rect 1174 2543 1175 2547
rect 1179 2543 1180 2547
rect 1174 2542 1180 2543
rect 1318 2547 1324 2548
rect 1318 2543 1319 2547
rect 1323 2543 1324 2547
rect 1318 2542 1324 2543
rect 1454 2547 1460 2548
rect 1454 2543 1455 2547
rect 1459 2543 1460 2547
rect 1454 2542 1460 2543
rect 1590 2547 1596 2548
rect 1590 2543 1591 2547
rect 1595 2543 1596 2547
rect 1590 2542 1596 2543
rect 1726 2547 1732 2548
rect 1726 2543 1727 2547
rect 1731 2543 1732 2547
rect 1726 2542 1732 2543
rect 1886 2543 1892 2544
rect 1886 2539 1887 2543
rect 1891 2539 1892 2543
rect 1886 2538 1892 2539
rect 2038 2543 2044 2544
rect 2038 2539 2039 2543
rect 2043 2539 2044 2543
rect 2038 2538 2044 2539
rect 2214 2543 2220 2544
rect 2214 2539 2215 2543
rect 2219 2539 2220 2543
rect 2214 2538 2220 2539
rect 2398 2543 2404 2544
rect 2398 2539 2399 2543
rect 2403 2539 2404 2543
rect 2398 2538 2404 2539
rect 2574 2543 2580 2544
rect 2574 2539 2575 2543
rect 2579 2539 2580 2543
rect 2574 2538 2580 2539
rect 2742 2543 2748 2544
rect 2742 2539 2743 2543
rect 2747 2539 2748 2543
rect 2742 2538 2748 2539
rect 2902 2543 2908 2544
rect 2902 2539 2903 2543
rect 2907 2539 2908 2543
rect 2902 2538 2908 2539
rect 3054 2543 3060 2544
rect 3054 2539 3055 2543
rect 3059 2539 3060 2543
rect 3054 2538 3060 2539
rect 3198 2543 3204 2544
rect 3198 2539 3199 2543
rect 3203 2539 3204 2543
rect 3198 2538 3204 2539
rect 3342 2543 3348 2544
rect 3342 2539 3343 2543
rect 3347 2539 3348 2543
rect 3342 2538 3348 2539
rect 3478 2543 3484 2544
rect 3478 2539 3479 2543
rect 3483 2539 3484 2543
rect 3478 2538 3484 2539
rect 110 2537 116 2538
rect 110 2533 111 2537
rect 115 2533 116 2537
rect 110 2532 116 2533
rect 1822 2537 1828 2538
rect 1822 2533 1823 2537
rect 1827 2533 1828 2537
rect 1822 2532 1828 2533
rect 1862 2533 1868 2534
rect 1862 2529 1863 2533
rect 1867 2529 1868 2533
rect 1862 2528 1868 2529
rect 3574 2533 3580 2534
rect 3574 2529 3575 2533
rect 3579 2529 3580 2533
rect 3574 2528 3580 2529
rect 110 2520 116 2521
rect 110 2516 111 2520
rect 115 2516 116 2520
rect 110 2515 116 2516
rect 1822 2520 1828 2521
rect 1822 2516 1823 2520
rect 1827 2516 1828 2520
rect 1822 2515 1828 2516
rect 1862 2516 1868 2517
rect 1862 2512 1863 2516
rect 1867 2512 1868 2516
rect 1862 2511 1868 2512
rect 3574 2516 3580 2517
rect 3574 2512 3575 2516
rect 3579 2512 3580 2516
rect 3574 2511 3580 2512
rect 278 2507 284 2508
rect 278 2503 279 2507
rect 283 2503 284 2507
rect 278 2502 284 2503
rect 478 2507 484 2508
rect 478 2503 479 2507
rect 483 2503 484 2507
rect 478 2502 484 2503
rect 678 2507 684 2508
rect 678 2503 679 2507
rect 683 2503 684 2507
rect 678 2502 684 2503
rect 862 2507 868 2508
rect 862 2503 863 2507
rect 867 2503 868 2507
rect 862 2502 868 2503
rect 1030 2507 1036 2508
rect 1030 2503 1031 2507
rect 1035 2503 1036 2507
rect 1030 2502 1036 2503
rect 1182 2507 1188 2508
rect 1182 2503 1183 2507
rect 1187 2503 1188 2507
rect 1182 2502 1188 2503
rect 1326 2507 1332 2508
rect 1326 2503 1327 2507
rect 1331 2503 1332 2507
rect 1326 2502 1332 2503
rect 1462 2507 1468 2508
rect 1462 2503 1463 2507
rect 1467 2503 1468 2507
rect 1462 2502 1468 2503
rect 1598 2507 1604 2508
rect 1598 2503 1599 2507
rect 1603 2503 1604 2507
rect 1598 2502 1604 2503
rect 1734 2507 1740 2508
rect 1734 2503 1735 2507
rect 1739 2503 1740 2507
rect 1734 2502 1740 2503
rect 1894 2503 1900 2504
rect 1894 2499 1895 2503
rect 1899 2499 1900 2503
rect 1894 2498 1900 2499
rect 2046 2503 2052 2504
rect 2046 2499 2047 2503
rect 2051 2499 2052 2503
rect 2046 2498 2052 2499
rect 2222 2503 2228 2504
rect 2222 2499 2223 2503
rect 2227 2499 2228 2503
rect 2222 2498 2228 2499
rect 2406 2503 2412 2504
rect 2406 2499 2407 2503
rect 2411 2499 2412 2503
rect 2406 2498 2412 2499
rect 2582 2503 2588 2504
rect 2582 2499 2583 2503
rect 2587 2499 2588 2503
rect 2582 2498 2588 2499
rect 2750 2503 2756 2504
rect 2750 2499 2751 2503
rect 2755 2499 2756 2503
rect 2750 2498 2756 2499
rect 2910 2503 2916 2504
rect 2910 2499 2911 2503
rect 2915 2499 2916 2503
rect 2910 2498 2916 2499
rect 3062 2503 3068 2504
rect 3062 2499 3063 2503
rect 3067 2499 3068 2503
rect 3062 2498 3068 2499
rect 3206 2503 3212 2504
rect 3206 2499 3207 2503
rect 3211 2499 3212 2503
rect 3206 2498 3212 2499
rect 3350 2503 3356 2504
rect 3350 2499 3351 2503
rect 3355 2499 3356 2503
rect 3350 2498 3356 2499
rect 3486 2503 3492 2504
rect 3486 2499 3487 2503
rect 3491 2499 3492 2503
rect 3486 2498 3492 2499
rect 182 2469 188 2470
rect 182 2465 183 2469
rect 187 2465 188 2469
rect 182 2464 188 2465
rect 318 2469 324 2470
rect 318 2465 319 2469
rect 323 2465 324 2469
rect 318 2464 324 2465
rect 462 2469 468 2470
rect 462 2465 463 2469
rect 467 2465 468 2469
rect 462 2464 468 2465
rect 606 2469 612 2470
rect 606 2465 607 2469
rect 611 2465 612 2469
rect 606 2464 612 2465
rect 742 2469 748 2470
rect 742 2465 743 2469
rect 747 2465 748 2469
rect 742 2464 748 2465
rect 878 2469 884 2470
rect 878 2465 879 2469
rect 883 2465 884 2469
rect 878 2464 884 2465
rect 1006 2469 1012 2470
rect 1006 2465 1007 2469
rect 1011 2465 1012 2469
rect 1006 2464 1012 2465
rect 1126 2469 1132 2470
rect 1126 2465 1127 2469
rect 1131 2465 1132 2469
rect 1126 2464 1132 2465
rect 1238 2469 1244 2470
rect 1238 2465 1239 2469
rect 1243 2465 1244 2469
rect 1238 2464 1244 2465
rect 1342 2469 1348 2470
rect 1342 2465 1343 2469
rect 1347 2465 1348 2469
rect 1342 2464 1348 2465
rect 1446 2469 1452 2470
rect 1446 2465 1447 2469
rect 1451 2465 1452 2469
rect 1446 2464 1452 2465
rect 1550 2469 1556 2470
rect 1550 2465 1551 2469
rect 1555 2465 1556 2469
rect 1550 2464 1556 2465
rect 1646 2469 1652 2470
rect 1646 2465 1647 2469
rect 1651 2465 1652 2469
rect 1646 2464 1652 2465
rect 1734 2469 1740 2470
rect 1734 2465 1735 2469
rect 1739 2465 1740 2469
rect 1734 2464 1740 2465
rect 1894 2469 1900 2470
rect 1894 2465 1895 2469
rect 1899 2465 1900 2469
rect 1894 2464 1900 2465
rect 1990 2469 1996 2470
rect 1990 2465 1991 2469
rect 1995 2465 1996 2469
rect 1990 2464 1996 2465
rect 2126 2469 2132 2470
rect 2126 2465 2127 2469
rect 2131 2465 2132 2469
rect 2126 2464 2132 2465
rect 2278 2469 2284 2470
rect 2278 2465 2279 2469
rect 2283 2465 2284 2469
rect 2278 2464 2284 2465
rect 2438 2469 2444 2470
rect 2438 2465 2439 2469
rect 2443 2465 2444 2469
rect 2438 2464 2444 2465
rect 2598 2469 2604 2470
rect 2598 2465 2599 2469
rect 2603 2465 2604 2469
rect 2598 2464 2604 2465
rect 2766 2469 2772 2470
rect 2766 2465 2767 2469
rect 2771 2465 2772 2469
rect 2766 2464 2772 2465
rect 2942 2469 2948 2470
rect 2942 2465 2943 2469
rect 2947 2465 2948 2469
rect 2942 2464 2948 2465
rect 3118 2469 3124 2470
rect 3118 2465 3119 2469
rect 3123 2465 3124 2469
rect 3118 2464 3124 2465
rect 3294 2469 3300 2470
rect 3294 2465 3295 2469
rect 3299 2465 3300 2469
rect 3294 2464 3300 2465
rect 3470 2469 3476 2470
rect 3470 2465 3471 2469
rect 3475 2465 3476 2469
rect 3470 2464 3476 2465
rect 110 2456 116 2457
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 110 2451 116 2452
rect 1822 2456 1828 2457
rect 1822 2452 1823 2456
rect 1827 2452 1828 2456
rect 1822 2451 1828 2452
rect 1862 2456 1868 2457
rect 1862 2452 1863 2456
rect 1867 2452 1868 2456
rect 1862 2451 1868 2452
rect 3574 2456 3580 2457
rect 3574 2452 3575 2456
rect 3579 2452 3580 2456
rect 3574 2451 3580 2452
rect 110 2439 116 2440
rect 110 2435 111 2439
rect 115 2435 116 2439
rect 110 2434 116 2435
rect 1822 2439 1828 2440
rect 1822 2435 1823 2439
rect 1827 2435 1828 2439
rect 1822 2434 1828 2435
rect 1862 2439 1868 2440
rect 1862 2435 1863 2439
rect 1867 2435 1868 2439
rect 1862 2434 1868 2435
rect 3574 2439 3580 2440
rect 3574 2435 3575 2439
rect 3579 2435 3580 2439
rect 3574 2434 3580 2435
rect 174 2429 180 2430
rect 174 2425 175 2429
rect 179 2425 180 2429
rect 174 2424 180 2425
rect 310 2429 316 2430
rect 310 2425 311 2429
rect 315 2425 316 2429
rect 310 2424 316 2425
rect 454 2429 460 2430
rect 454 2425 455 2429
rect 459 2425 460 2429
rect 454 2424 460 2425
rect 598 2429 604 2430
rect 598 2425 599 2429
rect 603 2425 604 2429
rect 598 2424 604 2425
rect 734 2429 740 2430
rect 734 2425 735 2429
rect 739 2425 740 2429
rect 734 2424 740 2425
rect 870 2429 876 2430
rect 870 2425 871 2429
rect 875 2425 876 2429
rect 870 2424 876 2425
rect 998 2429 1004 2430
rect 998 2425 999 2429
rect 1003 2425 1004 2429
rect 998 2424 1004 2425
rect 1118 2429 1124 2430
rect 1118 2425 1119 2429
rect 1123 2425 1124 2429
rect 1118 2424 1124 2425
rect 1230 2429 1236 2430
rect 1230 2425 1231 2429
rect 1235 2425 1236 2429
rect 1230 2424 1236 2425
rect 1334 2429 1340 2430
rect 1334 2425 1335 2429
rect 1339 2425 1340 2429
rect 1334 2424 1340 2425
rect 1438 2429 1444 2430
rect 1438 2425 1439 2429
rect 1443 2425 1444 2429
rect 1438 2424 1444 2425
rect 1542 2429 1548 2430
rect 1542 2425 1543 2429
rect 1547 2425 1548 2429
rect 1542 2424 1548 2425
rect 1638 2429 1644 2430
rect 1638 2425 1639 2429
rect 1643 2425 1644 2429
rect 1638 2424 1644 2425
rect 1726 2429 1732 2430
rect 1726 2425 1727 2429
rect 1731 2425 1732 2429
rect 1726 2424 1732 2425
rect 1886 2429 1892 2430
rect 1886 2425 1887 2429
rect 1891 2425 1892 2429
rect 1886 2424 1892 2425
rect 1982 2429 1988 2430
rect 1982 2425 1983 2429
rect 1987 2425 1988 2429
rect 1982 2424 1988 2425
rect 2118 2429 2124 2430
rect 2118 2425 2119 2429
rect 2123 2425 2124 2429
rect 2118 2424 2124 2425
rect 2270 2429 2276 2430
rect 2270 2425 2271 2429
rect 2275 2425 2276 2429
rect 2270 2424 2276 2425
rect 2430 2429 2436 2430
rect 2430 2425 2431 2429
rect 2435 2425 2436 2429
rect 2430 2424 2436 2425
rect 2590 2429 2596 2430
rect 2590 2425 2591 2429
rect 2595 2425 2596 2429
rect 2590 2424 2596 2425
rect 2758 2429 2764 2430
rect 2758 2425 2759 2429
rect 2763 2425 2764 2429
rect 2758 2424 2764 2425
rect 2934 2429 2940 2430
rect 2934 2425 2935 2429
rect 2939 2425 2940 2429
rect 2934 2424 2940 2425
rect 3110 2429 3116 2430
rect 3110 2425 3111 2429
rect 3115 2425 3116 2429
rect 3110 2424 3116 2425
rect 3286 2429 3292 2430
rect 3286 2425 3287 2429
rect 3291 2425 3292 2429
rect 3286 2424 3292 2425
rect 3462 2429 3468 2430
rect 3462 2425 3463 2429
rect 3467 2425 3468 2429
rect 3462 2424 3468 2425
rect 150 2399 156 2400
rect 150 2395 151 2399
rect 155 2395 156 2399
rect 150 2394 156 2395
rect 318 2399 324 2400
rect 318 2395 319 2399
rect 323 2395 324 2399
rect 318 2394 324 2395
rect 478 2399 484 2400
rect 478 2395 479 2399
rect 483 2395 484 2399
rect 478 2394 484 2395
rect 638 2399 644 2400
rect 638 2395 639 2399
rect 643 2395 644 2399
rect 638 2394 644 2395
rect 782 2399 788 2400
rect 782 2395 783 2399
rect 787 2395 788 2399
rect 782 2394 788 2395
rect 918 2399 924 2400
rect 918 2395 919 2399
rect 923 2395 924 2399
rect 918 2394 924 2395
rect 1046 2399 1052 2400
rect 1046 2395 1047 2399
rect 1051 2395 1052 2399
rect 1046 2394 1052 2395
rect 1174 2399 1180 2400
rect 1174 2395 1175 2399
rect 1179 2395 1180 2399
rect 1174 2394 1180 2395
rect 1302 2399 1308 2400
rect 1302 2395 1303 2399
rect 1307 2395 1308 2399
rect 1302 2394 1308 2395
rect 1430 2399 1436 2400
rect 1430 2395 1431 2399
rect 1435 2395 1436 2399
rect 1430 2394 1436 2395
rect 2350 2399 2356 2400
rect 2350 2395 2351 2399
rect 2355 2395 2356 2399
rect 2350 2394 2356 2395
rect 2502 2399 2508 2400
rect 2502 2395 2503 2399
rect 2507 2395 2508 2399
rect 2502 2394 2508 2395
rect 2654 2399 2660 2400
rect 2654 2395 2655 2399
rect 2659 2395 2660 2399
rect 2654 2394 2660 2395
rect 2806 2399 2812 2400
rect 2806 2395 2807 2399
rect 2811 2395 2812 2399
rect 2806 2394 2812 2395
rect 2966 2399 2972 2400
rect 2966 2395 2967 2399
rect 2971 2395 2972 2399
rect 2966 2394 2972 2395
rect 3134 2399 3140 2400
rect 3134 2395 3135 2399
rect 3139 2395 3140 2399
rect 3134 2394 3140 2395
rect 3302 2399 3308 2400
rect 3302 2395 3303 2399
rect 3307 2395 3308 2399
rect 3302 2394 3308 2395
rect 3470 2399 3476 2400
rect 3470 2395 3471 2399
rect 3475 2395 3476 2399
rect 3470 2394 3476 2395
rect 110 2389 116 2390
rect 110 2385 111 2389
rect 115 2385 116 2389
rect 110 2384 116 2385
rect 1822 2389 1828 2390
rect 1822 2385 1823 2389
rect 1827 2385 1828 2389
rect 1822 2384 1828 2385
rect 1862 2389 1868 2390
rect 1862 2385 1863 2389
rect 1867 2385 1868 2389
rect 1862 2384 1868 2385
rect 3574 2389 3580 2390
rect 3574 2385 3575 2389
rect 3579 2385 3580 2389
rect 3574 2384 3580 2385
rect 110 2372 116 2373
rect 110 2368 111 2372
rect 115 2368 116 2372
rect 110 2367 116 2368
rect 1822 2372 1828 2373
rect 1822 2368 1823 2372
rect 1827 2368 1828 2372
rect 1822 2367 1828 2368
rect 1862 2372 1868 2373
rect 1862 2368 1863 2372
rect 1867 2368 1868 2372
rect 1862 2367 1868 2368
rect 3574 2372 3580 2373
rect 3574 2368 3575 2372
rect 3579 2368 3580 2372
rect 3574 2367 3580 2368
rect 158 2359 164 2360
rect 158 2355 159 2359
rect 163 2355 164 2359
rect 158 2354 164 2355
rect 326 2359 332 2360
rect 326 2355 327 2359
rect 331 2355 332 2359
rect 326 2354 332 2355
rect 486 2359 492 2360
rect 486 2355 487 2359
rect 491 2355 492 2359
rect 486 2354 492 2355
rect 646 2359 652 2360
rect 646 2355 647 2359
rect 651 2355 652 2359
rect 646 2354 652 2355
rect 790 2359 796 2360
rect 790 2355 791 2359
rect 795 2355 796 2359
rect 790 2354 796 2355
rect 926 2359 932 2360
rect 926 2355 927 2359
rect 931 2355 932 2359
rect 926 2354 932 2355
rect 1054 2359 1060 2360
rect 1054 2355 1055 2359
rect 1059 2355 1060 2359
rect 1054 2354 1060 2355
rect 1182 2359 1188 2360
rect 1182 2355 1183 2359
rect 1187 2355 1188 2359
rect 1182 2354 1188 2355
rect 1310 2359 1316 2360
rect 1310 2355 1311 2359
rect 1315 2355 1316 2359
rect 1310 2354 1316 2355
rect 1438 2359 1444 2360
rect 1438 2355 1439 2359
rect 1443 2355 1444 2359
rect 1438 2354 1444 2355
rect 2358 2359 2364 2360
rect 2358 2355 2359 2359
rect 2363 2355 2364 2359
rect 2358 2354 2364 2355
rect 2510 2359 2516 2360
rect 2510 2355 2511 2359
rect 2515 2355 2516 2359
rect 2510 2354 2516 2355
rect 2662 2359 2668 2360
rect 2662 2355 2663 2359
rect 2667 2355 2668 2359
rect 2662 2354 2668 2355
rect 2814 2359 2820 2360
rect 2814 2355 2815 2359
rect 2819 2355 2820 2359
rect 2814 2354 2820 2355
rect 2974 2359 2980 2360
rect 2974 2355 2975 2359
rect 2979 2355 2980 2359
rect 2974 2354 2980 2355
rect 3142 2359 3148 2360
rect 3142 2355 3143 2359
rect 3147 2355 3148 2359
rect 3142 2354 3148 2355
rect 3310 2359 3316 2360
rect 3310 2355 3311 2359
rect 3315 2355 3316 2359
rect 3310 2354 3316 2355
rect 3478 2359 3484 2360
rect 3478 2355 3479 2359
rect 3483 2355 3484 2359
rect 3478 2354 3484 2355
rect 142 2321 148 2322
rect 142 2317 143 2321
rect 147 2317 148 2321
rect 142 2316 148 2317
rect 262 2321 268 2322
rect 262 2317 263 2321
rect 267 2317 268 2321
rect 262 2316 268 2317
rect 406 2321 412 2322
rect 406 2317 407 2321
rect 411 2317 412 2321
rect 406 2316 412 2317
rect 542 2321 548 2322
rect 542 2317 543 2321
rect 547 2317 548 2321
rect 542 2316 548 2317
rect 678 2321 684 2322
rect 678 2317 679 2321
rect 683 2317 684 2321
rect 678 2316 684 2317
rect 806 2321 812 2322
rect 806 2317 807 2321
rect 811 2317 812 2321
rect 806 2316 812 2317
rect 926 2321 932 2322
rect 926 2317 927 2321
rect 931 2317 932 2321
rect 926 2316 932 2317
rect 1038 2321 1044 2322
rect 1038 2317 1039 2321
rect 1043 2317 1044 2321
rect 1038 2316 1044 2317
rect 1158 2321 1164 2322
rect 1158 2317 1159 2321
rect 1163 2317 1164 2321
rect 1158 2316 1164 2317
rect 1278 2321 1284 2322
rect 1278 2317 1279 2321
rect 1283 2317 1284 2321
rect 1278 2316 1284 2317
rect 2350 2321 2356 2322
rect 2350 2317 2351 2321
rect 2355 2317 2356 2321
rect 2350 2316 2356 2317
rect 2446 2321 2452 2322
rect 2446 2317 2447 2321
rect 2451 2317 2452 2321
rect 2446 2316 2452 2317
rect 2558 2321 2564 2322
rect 2558 2317 2559 2321
rect 2563 2317 2564 2321
rect 2558 2316 2564 2317
rect 2702 2321 2708 2322
rect 2702 2317 2703 2321
rect 2707 2317 2708 2321
rect 2702 2316 2708 2317
rect 2878 2321 2884 2322
rect 2878 2317 2879 2321
rect 2883 2317 2884 2321
rect 2878 2316 2884 2317
rect 3078 2321 3084 2322
rect 3078 2317 3079 2321
rect 3083 2317 3084 2321
rect 3078 2316 3084 2317
rect 3286 2321 3292 2322
rect 3286 2317 3287 2321
rect 3291 2317 3292 2321
rect 3286 2316 3292 2317
rect 3486 2321 3492 2322
rect 3486 2317 3487 2321
rect 3491 2317 3492 2321
rect 3486 2316 3492 2317
rect 110 2308 116 2309
rect 110 2304 111 2308
rect 115 2304 116 2308
rect 110 2303 116 2304
rect 1822 2308 1828 2309
rect 1822 2304 1823 2308
rect 1827 2304 1828 2308
rect 1822 2303 1828 2304
rect 1862 2308 1868 2309
rect 1862 2304 1863 2308
rect 1867 2304 1868 2308
rect 1862 2303 1868 2304
rect 3574 2308 3580 2309
rect 3574 2304 3575 2308
rect 3579 2304 3580 2308
rect 3574 2303 3580 2304
rect 110 2291 116 2292
rect 110 2287 111 2291
rect 115 2287 116 2291
rect 110 2286 116 2287
rect 1822 2291 1828 2292
rect 1822 2287 1823 2291
rect 1827 2287 1828 2291
rect 1822 2286 1828 2287
rect 1862 2291 1868 2292
rect 1862 2287 1863 2291
rect 1867 2287 1868 2291
rect 1862 2286 1868 2287
rect 3574 2291 3580 2292
rect 3574 2287 3575 2291
rect 3579 2287 3580 2291
rect 3574 2286 3580 2287
rect 134 2281 140 2282
rect 134 2277 135 2281
rect 139 2277 140 2281
rect 134 2276 140 2277
rect 254 2281 260 2282
rect 254 2277 255 2281
rect 259 2277 260 2281
rect 254 2276 260 2277
rect 398 2281 404 2282
rect 398 2277 399 2281
rect 403 2277 404 2281
rect 398 2276 404 2277
rect 534 2281 540 2282
rect 534 2277 535 2281
rect 539 2277 540 2281
rect 534 2276 540 2277
rect 670 2281 676 2282
rect 670 2277 671 2281
rect 675 2277 676 2281
rect 670 2276 676 2277
rect 798 2281 804 2282
rect 798 2277 799 2281
rect 803 2277 804 2281
rect 798 2276 804 2277
rect 918 2281 924 2282
rect 918 2277 919 2281
rect 923 2277 924 2281
rect 918 2276 924 2277
rect 1030 2281 1036 2282
rect 1030 2277 1031 2281
rect 1035 2277 1036 2281
rect 1030 2276 1036 2277
rect 1150 2281 1156 2282
rect 1150 2277 1151 2281
rect 1155 2277 1156 2281
rect 1150 2276 1156 2277
rect 1270 2281 1276 2282
rect 1270 2277 1271 2281
rect 1275 2277 1276 2281
rect 1270 2276 1276 2277
rect 2342 2281 2348 2282
rect 2342 2277 2343 2281
rect 2347 2277 2348 2281
rect 2342 2276 2348 2277
rect 2438 2281 2444 2282
rect 2438 2277 2439 2281
rect 2443 2277 2444 2281
rect 2438 2276 2444 2277
rect 2550 2281 2556 2282
rect 2550 2277 2551 2281
rect 2555 2277 2556 2281
rect 2550 2276 2556 2277
rect 2694 2281 2700 2282
rect 2694 2277 2695 2281
rect 2699 2277 2700 2281
rect 2694 2276 2700 2277
rect 2870 2281 2876 2282
rect 2870 2277 2871 2281
rect 2875 2277 2876 2281
rect 2870 2276 2876 2277
rect 3070 2281 3076 2282
rect 3070 2277 3071 2281
rect 3075 2277 3076 2281
rect 3070 2276 3076 2277
rect 3278 2281 3284 2282
rect 3278 2277 3279 2281
rect 3283 2277 3284 2281
rect 3278 2276 3284 2277
rect 3478 2281 3484 2282
rect 3478 2277 3479 2281
rect 3483 2277 3484 2281
rect 3478 2276 3484 2277
rect 134 2259 140 2260
rect 134 2255 135 2259
rect 139 2255 140 2259
rect 134 2254 140 2255
rect 230 2259 236 2260
rect 230 2255 231 2259
rect 235 2255 236 2259
rect 230 2254 236 2255
rect 350 2259 356 2260
rect 350 2255 351 2259
rect 355 2255 356 2259
rect 350 2254 356 2255
rect 470 2259 476 2260
rect 470 2255 471 2259
rect 475 2255 476 2259
rect 470 2254 476 2255
rect 590 2259 596 2260
rect 590 2255 591 2259
rect 595 2255 596 2259
rect 590 2254 596 2255
rect 710 2259 716 2260
rect 710 2255 711 2259
rect 715 2255 716 2259
rect 710 2254 716 2255
rect 822 2259 828 2260
rect 822 2255 823 2259
rect 827 2255 828 2259
rect 822 2254 828 2255
rect 934 2259 940 2260
rect 934 2255 935 2259
rect 939 2255 940 2259
rect 934 2254 940 2255
rect 1054 2259 1060 2260
rect 1054 2255 1055 2259
rect 1059 2255 1060 2259
rect 1054 2254 1060 2255
rect 1174 2259 1180 2260
rect 1174 2255 1175 2259
rect 1179 2255 1180 2259
rect 1174 2254 1180 2255
rect 2334 2259 2340 2260
rect 2334 2255 2335 2259
rect 2339 2255 2340 2259
rect 2334 2254 2340 2255
rect 2446 2259 2452 2260
rect 2446 2255 2447 2259
rect 2451 2255 2452 2259
rect 2446 2254 2452 2255
rect 2582 2259 2588 2260
rect 2582 2255 2583 2259
rect 2587 2255 2588 2259
rect 2582 2254 2588 2255
rect 2734 2259 2740 2260
rect 2734 2255 2735 2259
rect 2739 2255 2740 2259
rect 2734 2254 2740 2255
rect 2910 2259 2916 2260
rect 2910 2255 2911 2259
rect 2915 2255 2916 2259
rect 2910 2254 2916 2255
rect 3102 2259 3108 2260
rect 3102 2255 3103 2259
rect 3107 2255 3108 2259
rect 3102 2254 3108 2255
rect 3302 2259 3308 2260
rect 3302 2255 3303 2259
rect 3307 2255 3308 2259
rect 3302 2254 3308 2255
rect 3478 2259 3484 2260
rect 3478 2255 3479 2259
rect 3483 2255 3484 2259
rect 3478 2254 3484 2255
rect 110 2249 116 2250
rect 110 2245 111 2249
rect 115 2245 116 2249
rect 110 2244 116 2245
rect 1822 2249 1828 2250
rect 1822 2245 1823 2249
rect 1827 2245 1828 2249
rect 1822 2244 1828 2245
rect 1862 2249 1868 2250
rect 1862 2245 1863 2249
rect 1867 2245 1868 2249
rect 1862 2244 1868 2245
rect 3574 2249 3580 2250
rect 3574 2245 3575 2249
rect 3579 2245 3580 2249
rect 3574 2244 3580 2245
rect 110 2232 116 2233
rect 110 2228 111 2232
rect 115 2228 116 2232
rect 110 2227 116 2228
rect 1822 2232 1828 2233
rect 1822 2228 1823 2232
rect 1827 2228 1828 2232
rect 1822 2227 1828 2228
rect 1862 2232 1868 2233
rect 1862 2228 1863 2232
rect 1867 2228 1868 2232
rect 1862 2227 1868 2228
rect 3574 2232 3580 2233
rect 3574 2228 3575 2232
rect 3579 2228 3580 2232
rect 3574 2227 3580 2228
rect 142 2219 148 2220
rect 142 2215 143 2219
rect 147 2215 148 2219
rect 142 2214 148 2215
rect 238 2219 244 2220
rect 238 2215 239 2219
rect 243 2215 244 2219
rect 238 2214 244 2215
rect 358 2219 364 2220
rect 358 2215 359 2219
rect 363 2215 364 2219
rect 358 2214 364 2215
rect 478 2219 484 2220
rect 478 2215 479 2219
rect 483 2215 484 2219
rect 478 2214 484 2215
rect 598 2219 604 2220
rect 598 2215 599 2219
rect 603 2215 604 2219
rect 598 2214 604 2215
rect 718 2219 724 2220
rect 718 2215 719 2219
rect 723 2215 724 2219
rect 718 2214 724 2215
rect 830 2219 836 2220
rect 830 2215 831 2219
rect 835 2215 836 2219
rect 830 2214 836 2215
rect 942 2219 948 2220
rect 942 2215 943 2219
rect 947 2215 948 2219
rect 942 2214 948 2215
rect 1062 2219 1068 2220
rect 1062 2215 1063 2219
rect 1067 2215 1068 2219
rect 1062 2214 1068 2215
rect 1182 2219 1188 2220
rect 1182 2215 1183 2219
rect 1187 2215 1188 2219
rect 1182 2214 1188 2215
rect 2342 2219 2348 2220
rect 2342 2215 2343 2219
rect 2347 2215 2348 2219
rect 2342 2214 2348 2215
rect 2454 2219 2460 2220
rect 2454 2215 2455 2219
rect 2459 2215 2460 2219
rect 2454 2214 2460 2215
rect 2590 2219 2596 2220
rect 2590 2215 2591 2219
rect 2595 2215 2596 2219
rect 2590 2214 2596 2215
rect 2742 2219 2748 2220
rect 2742 2215 2743 2219
rect 2747 2215 2748 2219
rect 2742 2214 2748 2215
rect 2918 2219 2924 2220
rect 2918 2215 2919 2219
rect 2923 2215 2924 2219
rect 2918 2214 2924 2215
rect 3110 2219 3116 2220
rect 3110 2215 3111 2219
rect 3115 2215 3116 2219
rect 3110 2214 3116 2215
rect 3310 2219 3316 2220
rect 3310 2215 3311 2219
rect 3315 2215 3316 2219
rect 3310 2214 3316 2215
rect 3486 2219 3492 2220
rect 3486 2215 3487 2219
rect 3491 2215 3492 2219
rect 3486 2214 3492 2215
rect 2254 2185 2260 2186
rect 142 2181 148 2182
rect 142 2177 143 2181
rect 147 2177 148 2181
rect 142 2176 148 2177
rect 246 2181 252 2182
rect 246 2177 247 2181
rect 251 2177 252 2181
rect 246 2176 252 2177
rect 382 2181 388 2182
rect 382 2177 383 2181
rect 387 2177 388 2181
rect 382 2176 388 2177
rect 518 2181 524 2182
rect 518 2177 519 2181
rect 523 2177 524 2181
rect 518 2176 524 2177
rect 654 2181 660 2182
rect 654 2177 655 2181
rect 659 2177 660 2181
rect 654 2176 660 2177
rect 782 2181 788 2182
rect 782 2177 783 2181
rect 787 2177 788 2181
rect 782 2176 788 2177
rect 910 2181 916 2182
rect 910 2177 911 2181
rect 915 2177 916 2181
rect 910 2176 916 2177
rect 1030 2181 1036 2182
rect 1030 2177 1031 2181
rect 1035 2177 1036 2181
rect 1030 2176 1036 2177
rect 1158 2181 1164 2182
rect 1158 2177 1159 2181
rect 1163 2177 1164 2181
rect 1158 2176 1164 2177
rect 1286 2181 1292 2182
rect 1286 2177 1287 2181
rect 1291 2177 1292 2181
rect 2254 2181 2255 2185
rect 2259 2181 2260 2185
rect 2254 2180 2260 2181
rect 2342 2185 2348 2186
rect 2342 2181 2343 2185
rect 2347 2181 2348 2185
rect 2342 2180 2348 2181
rect 2438 2185 2444 2186
rect 2438 2181 2439 2185
rect 2443 2181 2444 2185
rect 2438 2180 2444 2181
rect 2550 2185 2556 2186
rect 2550 2181 2551 2185
rect 2555 2181 2556 2185
rect 2550 2180 2556 2181
rect 2694 2185 2700 2186
rect 2694 2181 2695 2185
rect 2699 2181 2700 2185
rect 2694 2180 2700 2181
rect 2870 2185 2876 2186
rect 2870 2181 2871 2185
rect 2875 2181 2876 2185
rect 2870 2180 2876 2181
rect 3070 2185 3076 2186
rect 3070 2181 3071 2185
rect 3075 2181 3076 2185
rect 3070 2180 3076 2181
rect 3286 2185 3292 2186
rect 3286 2181 3287 2185
rect 3291 2181 3292 2185
rect 3286 2180 3292 2181
rect 3486 2185 3492 2186
rect 3486 2181 3487 2185
rect 3491 2181 3492 2185
rect 3486 2180 3492 2181
rect 1286 2176 1292 2177
rect 1862 2172 1868 2173
rect 110 2168 116 2169
rect 110 2164 111 2168
rect 115 2164 116 2168
rect 110 2163 116 2164
rect 1822 2168 1828 2169
rect 1822 2164 1823 2168
rect 1827 2164 1828 2168
rect 1862 2168 1863 2172
rect 1867 2168 1868 2172
rect 1862 2167 1868 2168
rect 3574 2172 3580 2173
rect 3574 2168 3575 2172
rect 3579 2168 3580 2172
rect 3574 2167 3580 2168
rect 1822 2163 1828 2164
rect 1862 2155 1868 2156
rect 110 2151 116 2152
rect 110 2147 111 2151
rect 115 2147 116 2151
rect 110 2146 116 2147
rect 1822 2151 1828 2152
rect 1822 2147 1823 2151
rect 1827 2147 1828 2151
rect 1862 2151 1863 2155
rect 1867 2151 1868 2155
rect 1862 2150 1868 2151
rect 3574 2155 3580 2156
rect 3574 2151 3575 2155
rect 3579 2151 3580 2155
rect 3574 2150 3580 2151
rect 1822 2146 1828 2147
rect 2246 2145 2252 2146
rect 134 2141 140 2142
rect 134 2137 135 2141
rect 139 2137 140 2141
rect 134 2136 140 2137
rect 238 2141 244 2142
rect 238 2137 239 2141
rect 243 2137 244 2141
rect 238 2136 244 2137
rect 374 2141 380 2142
rect 374 2137 375 2141
rect 379 2137 380 2141
rect 374 2136 380 2137
rect 510 2141 516 2142
rect 510 2137 511 2141
rect 515 2137 516 2141
rect 510 2136 516 2137
rect 646 2141 652 2142
rect 646 2137 647 2141
rect 651 2137 652 2141
rect 646 2136 652 2137
rect 774 2141 780 2142
rect 774 2137 775 2141
rect 779 2137 780 2141
rect 774 2136 780 2137
rect 902 2141 908 2142
rect 902 2137 903 2141
rect 907 2137 908 2141
rect 902 2136 908 2137
rect 1022 2141 1028 2142
rect 1022 2137 1023 2141
rect 1027 2137 1028 2141
rect 1022 2136 1028 2137
rect 1150 2141 1156 2142
rect 1150 2137 1151 2141
rect 1155 2137 1156 2141
rect 1150 2136 1156 2137
rect 1278 2141 1284 2142
rect 1278 2137 1279 2141
rect 1283 2137 1284 2141
rect 2246 2141 2247 2145
rect 2251 2141 2252 2145
rect 2246 2140 2252 2141
rect 2334 2145 2340 2146
rect 2334 2141 2335 2145
rect 2339 2141 2340 2145
rect 2334 2140 2340 2141
rect 2430 2145 2436 2146
rect 2430 2141 2431 2145
rect 2435 2141 2436 2145
rect 2430 2140 2436 2141
rect 2542 2145 2548 2146
rect 2542 2141 2543 2145
rect 2547 2141 2548 2145
rect 2542 2140 2548 2141
rect 2686 2145 2692 2146
rect 2686 2141 2687 2145
rect 2691 2141 2692 2145
rect 2686 2140 2692 2141
rect 2862 2145 2868 2146
rect 2862 2141 2863 2145
rect 2867 2141 2868 2145
rect 2862 2140 2868 2141
rect 3062 2145 3068 2146
rect 3062 2141 3063 2145
rect 3067 2141 3068 2145
rect 3062 2140 3068 2141
rect 3278 2145 3284 2146
rect 3278 2141 3279 2145
rect 3283 2141 3284 2145
rect 3278 2140 3284 2141
rect 3478 2145 3484 2146
rect 3478 2141 3479 2145
rect 3483 2141 3484 2145
rect 3478 2140 3484 2141
rect 1278 2136 1284 2137
rect 2150 2115 2156 2116
rect 134 2111 140 2112
rect 134 2107 135 2111
rect 139 2107 140 2111
rect 134 2106 140 2107
rect 230 2111 236 2112
rect 230 2107 231 2111
rect 235 2107 236 2111
rect 230 2106 236 2107
rect 358 2111 364 2112
rect 358 2107 359 2111
rect 363 2107 364 2111
rect 358 2106 364 2107
rect 478 2111 484 2112
rect 478 2107 479 2111
rect 483 2107 484 2111
rect 478 2106 484 2107
rect 598 2111 604 2112
rect 598 2107 599 2111
rect 603 2107 604 2111
rect 598 2106 604 2107
rect 718 2111 724 2112
rect 718 2107 719 2111
rect 723 2107 724 2111
rect 718 2106 724 2107
rect 830 2111 836 2112
rect 830 2107 831 2111
rect 835 2107 836 2111
rect 830 2106 836 2107
rect 942 2111 948 2112
rect 942 2107 943 2111
rect 947 2107 948 2111
rect 942 2106 948 2107
rect 1054 2111 1060 2112
rect 1054 2107 1055 2111
rect 1059 2107 1060 2111
rect 1054 2106 1060 2107
rect 1174 2111 1180 2112
rect 1174 2107 1175 2111
rect 1179 2107 1180 2111
rect 2150 2111 2151 2115
rect 2155 2111 2156 2115
rect 2150 2110 2156 2111
rect 2238 2115 2244 2116
rect 2238 2111 2239 2115
rect 2243 2111 2244 2115
rect 2238 2110 2244 2111
rect 2326 2115 2332 2116
rect 2326 2111 2327 2115
rect 2331 2111 2332 2115
rect 2326 2110 2332 2111
rect 2414 2115 2420 2116
rect 2414 2111 2415 2115
rect 2419 2111 2420 2115
rect 2414 2110 2420 2111
rect 2502 2115 2508 2116
rect 2502 2111 2503 2115
rect 2507 2111 2508 2115
rect 2502 2110 2508 2111
rect 2614 2115 2620 2116
rect 2614 2111 2615 2115
rect 2619 2111 2620 2115
rect 2614 2110 2620 2111
rect 2750 2115 2756 2116
rect 2750 2111 2751 2115
rect 2755 2111 2756 2115
rect 2750 2110 2756 2111
rect 2918 2115 2924 2116
rect 2918 2111 2919 2115
rect 2923 2111 2924 2115
rect 2918 2110 2924 2111
rect 3102 2115 3108 2116
rect 3102 2111 3103 2115
rect 3107 2111 3108 2115
rect 3102 2110 3108 2111
rect 3302 2115 3308 2116
rect 3302 2111 3303 2115
rect 3307 2111 3308 2115
rect 3302 2110 3308 2111
rect 3478 2115 3484 2116
rect 3478 2111 3479 2115
rect 3483 2111 3484 2115
rect 3478 2110 3484 2111
rect 1174 2106 1180 2107
rect 1862 2105 1868 2106
rect 110 2101 116 2102
rect 110 2097 111 2101
rect 115 2097 116 2101
rect 110 2096 116 2097
rect 1822 2101 1828 2102
rect 1822 2097 1823 2101
rect 1827 2097 1828 2101
rect 1862 2101 1863 2105
rect 1867 2101 1868 2105
rect 1862 2100 1868 2101
rect 3574 2105 3580 2106
rect 3574 2101 3575 2105
rect 3579 2101 3580 2105
rect 3574 2100 3580 2101
rect 1822 2096 1828 2097
rect 1862 2088 1868 2089
rect 110 2084 116 2085
rect 110 2080 111 2084
rect 115 2080 116 2084
rect 110 2079 116 2080
rect 1822 2084 1828 2085
rect 1822 2080 1823 2084
rect 1827 2080 1828 2084
rect 1862 2084 1863 2088
rect 1867 2084 1868 2088
rect 1862 2083 1868 2084
rect 3574 2088 3580 2089
rect 3574 2084 3575 2088
rect 3579 2084 3580 2088
rect 3574 2083 3580 2084
rect 1822 2079 1828 2080
rect 2158 2075 2164 2076
rect 142 2071 148 2072
rect 142 2067 143 2071
rect 147 2067 148 2071
rect 142 2066 148 2067
rect 238 2071 244 2072
rect 238 2067 239 2071
rect 243 2067 244 2071
rect 238 2066 244 2067
rect 366 2071 372 2072
rect 366 2067 367 2071
rect 371 2067 372 2071
rect 366 2066 372 2067
rect 486 2071 492 2072
rect 486 2067 487 2071
rect 491 2067 492 2071
rect 486 2066 492 2067
rect 606 2071 612 2072
rect 606 2067 607 2071
rect 611 2067 612 2071
rect 606 2066 612 2067
rect 726 2071 732 2072
rect 726 2067 727 2071
rect 731 2067 732 2071
rect 726 2066 732 2067
rect 838 2071 844 2072
rect 838 2067 839 2071
rect 843 2067 844 2071
rect 838 2066 844 2067
rect 950 2071 956 2072
rect 950 2067 951 2071
rect 955 2067 956 2071
rect 950 2066 956 2067
rect 1062 2071 1068 2072
rect 1062 2067 1063 2071
rect 1067 2067 1068 2071
rect 1062 2066 1068 2067
rect 1182 2071 1188 2072
rect 1182 2067 1183 2071
rect 1187 2067 1188 2071
rect 2158 2071 2159 2075
rect 2163 2071 2164 2075
rect 2158 2070 2164 2071
rect 2246 2075 2252 2076
rect 2246 2071 2247 2075
rect 2251 2071 2252 2075
rect 2246 2070 2252 2071
rect 2334 2075 2340 2076
rect 2334 2071 2335 2075
rect 2339 2071 2340 2075
rect 2334 2070 2340 2071
rect 2422 2075 2428 2076
rect 2422 2071 2423 2075
rect 2427 2071 2428 2075
rect 2422 2070 2428 2071
rect 2510 2075 2516 2076
rect 2510 2071 2511 2075
rect 2515 2071 2516 2075
rect 2510 2070 2516 2071
rect 2622 2075 2628 2076
rect 2622 2071 2623 2075
rect 2627 2071 2628 2075
rect 2622 2070 2628 2071
rect 2758 2075 2764 2076
rect 2758 2071 2759 2075
rect 2763 2071 2764 2075
rect 2758 2070 2764 2071
rect 2926 2075 2932 2076
rect 2926 2071 2927 2075
rect 2931 2071 2932 2075
rect 2926 2070 2932 2071
rect 3110 2075 3116 2076
rect 3110 2071 3111 2075
rect 3115 2071 3116 2075
rect 3110 2070 3116 2071
rect 3310 2075 3316 2076
rect 3310 2071 3311 2075
rect 3315 2071 3316 2075
rect 3310 2070 3316 2071
rect 3486 2075 3492 2076
rect 3486 2071 3487 2075
rect 3491 2071 3492 2075
rect 3486 2070 3492 2071
rect 1182 2066 1188 2067
rect 1998 2037 2004 2038
rect 1998 2033 1999 2037
rect 2003 2033 2004 2037
rect 1998 2032 2004 2033
rect 2126 2037 2132 2038
rect 2126 2033 2127 2037
rect 2131 2033 2132 2037
rect 2126 2032 2132 2033
rect 2254 2037 2260 2038
rect 2254 2033 2255 2037
rect 2259 2033 2260 2037
rect 2254 2032 2260 2033
rect 2398 2037 2404 2038
rect 2398 2033 2399 2037
rect 2403 2033 2404 2037
rect 2398 2032 2404 2033
rect 2550 2037 2556 2038
rect 2550 2033 2551 2037
rect 2555 2033 2556 2037
rect 2550 2032 2556 2033
rect 2710 2037 2716 2038
rect 2710 2033 2711 2037
rect 2715 2033 2716 2037
rect 2710 2032 2716 2033
rect 2878 2037 2884 2038
rect 2878 2033 2879 2037
rect 2883 2033 2884 2037
rect 2878 2032 2884 2033
rect 3062 2037 3068 2038
rect 3062 2033 3063 2037
rect 3067 2033 3068 2037
rect 3062 2032 3068 2033
rect 3246 2037 3252 2038
rect 3246 2033 3247 2037
rect 3251 2033 3252 2037
rect 3246 2032 3252 2033
rect 3438 2037 3444 2038
rect 3438 2033 3439 2037
rect 3443 2033 3444 2037
rect 3438 2032 3444 2033
rect 166 2025 172 2026
rect 166 2021 167 2025
rect 171 2021 172 2025
rect 166 2020 172 2021
rect 310 2025 316 2026
rect 310 2021 311 2025
rect 315 2021 316 2025
rect 310 2020 316 2021
rect 446 2025 452 2026
rect 446 2021 447 2025
rect 451 2021 452 2025
rect 446 2020 452 2021
rect 574 2025 580 2026
rect 574 2021 575 2025
rect 579 2021 580 2025
rect 574 2020 580 2021
rect 694 2025 700 2026
rect 694 2021 695 2025
rect 699 2021 700 2025
rect 694 2020 700 2021
rect 806 2025 812 2026
rect 806 2021 807 2025
rect 811 2021 812 2025
rect 806 2020 812 2021
rect 910 2025 916 2026
rect 910 2021 911 2025
rect 915 2021 916 2025
rect 910 2020 916 2021
rect 1014 2025 1020 2026
rect 1014 2021 1015 2025
rect 1019 2021 1020 2025
rect 1014 2020 1020 2021
rect 1118 2025 1124 2026
rect 1118 2021 1119 2025
rect 1123 2021 1124 2025
rect 1118 2020 1124 2021
rect 1222 2025 1228 2026
rect 1222 2021 1223 2025
rect 1227 2021 1228 2025
rect 1222 2020 1228 2021
rect 1326 2025 1332 2026
rect 1326 2021 1327 2025
rect 1331 2021 1332 2025
rect 1326 2020 1332 2021
rect 1862 2024 1868 2025
rect 1862 2020 1863 2024
rect 1867 2020 1868 2024
rect 1862 2019 1868 2020
rect 3574 2024 3580 2025
rect 3574 2020 3575 2024
rect 3579 2020 3580 2024
rect 3574 2019 3580 2020
rect 110 2012 116 2013
rect 110 2008 111 2012
rect 115 2008 116 2012
rect 110 2007 116 2008
rect 1822 2012 1828 2013
rect 1822 2008 1823 2012
rect 1827 2008 1828 2012
rect 1822 2007 1828 2008
rect 1862 2007 1868 2008
rect 1862 2003 1863 2007
rect 1867 2003 1868 2007
rect 1862 2002 1868 2003
rect 3574 2007 3580 2008
rect 3574 2003 3575 2007
rect 3579 2003 3580 2007
rect 3574 2002 3580 2003
rect 1990 1997 1996 1998
rect 110 1995 116 1996
rect 110 1991 111 1995
rect 115 1991 116 1995
rect 110 1990 116 1991
rect 1822 1995 1828 1996
rect 1822 1991 1823 1995
rect 1827 1991 1828 1995
rect 1990 1993 1991 1997
rect 1995 1993 1996 1997
rect 1990 1992 1996 1993
rect 2118 1997 2124 1998
rect 2118 1993 2119 1997
rect 2123 1993 2124 1997
rect 2118 1992 2124 1993
rect 2246 1997 2252 1998
rect 2246 1993 2247 1997
rect 2251 1993 2252 1997
rect 2246 1992 2252 1993
rect 2390 1997 2396 1998
rect 2390 1993 2391 1997
rect 2395 1993 2396 1997
rect 2390 1992 2396 1993
rect 2542 1997 2548 1998
rect 2542 1993 2543 1997
rect 2547 1993 2548 1997
rect 2542 1992 2548 1993
rect 2702 1997 2708 1998
rect 2702 1993 2703 1997
rect 2707 1993 2708 1997
rect 2702 1992 2708 1993
rect 2870 1997 2876 1998
rect 2870 1993 2871 1997
rect 2875 1993 2876 1997
rect 2870 1992 2876 1993
rect 3054 1997 3060 1998
rect 3054 1993 3055 1997
rect 3059 1993 3060 1997
rect 3054 1992 3060 1993
rect 3238 1997 3244 1998
rect 3238 1993 3239 1997
rect 3243 1993 3244 1997
rect 3238 1992 3244 1993
rect 3430 1997 3436 1998
rect 3430 1993 3431 1997
rect 3435 1993 3436 1997
rect 3430 1992 3436 1993
rect 1822 1990 1828 1991
rect 158 1985 164 1986
rect 158 1981 159 1985
rect 163 1981 164 1985
rect 158 1980 164 1981
rect 302 1985 308 1986
rect 302 1981 303 1985
rect 307 1981 308 1985
rect 302 1980 308 1981
rect 438 1985 444 1986
rect 438 1981 439 1985
rect 443 1981 444 1985
rect 438 1980 444 1981
rect 566 1985 572 1986
rect 566 1981 567 1985
rect 571 1981 572 1985
rect 566 1980 572 1981
rect 686 1985 692 1986
rect 686 1981 687 1985
rect 691 1981 692 1985
rect 686 1980 692 1981
rect 798 1985 804 1986
rect 798 1981 799 1985
rect 803 1981 804 1985
rect 798 1980 804 1981
rect 902 1985 908 1986
rect 902 1981 903 1985
rect 907 1981 908 1985
rect 902 1980 908 1981
rect 1006 1985 1012 1986
rect 1006 1981 1007 1985
rect 1011 1981 1012 1985
rect 1006 1980 1012 1981
rect 1110 1985 1116 1986
rect 1110 1981 1111 1985
rect 1115 1981 1116 1985
rect 1110 1980 1116 1981
rect 1214 1985 1220 1986
rect 1214 1981 1215 1985
rect 1219 1981 1220 1985
rect 1214 1980 1220 1981
rect 1318 1985 1324 1986
rect 1318 1981 1319 1985
rect 1323 1981 1324 1985
rect 1318 1980 1324 1981
rect 1902 1967 1908 1968
rect 158 1963 164 1964
rect 158 1959 159 1963
rect 163 1959 164 1963
rect 158 1958 164 1959
rect 294 1963 300 1964
rect 294 1959 295 1963
rect 299 1959 300 1963
rect 294 1958 300 1959
rect 438 1963 444 1964
rect 438 1959 439 1963
rect 443 1959 444 1963
rect 438 1958 444 1959
rect 582 1963 588 1964
rect 582 1959 583 1963
rect 587 1959 588 1963
rect 582 1958 588 1959
rect 718 1963 724 1964
rect 718 1959 719 1963
rect 723 1959 724 1963
rect 718 1958 724 1959
rect 854 1963 860 1964
rect 854 1959 855 1963
rect 859 1959 860 1963
rect 854 1958 860 1959
rect 990 1963 996 1964
rect 990 1959 991 1963
rect 995 1959 996 1963
rect 990 1958 996 1959
rect 1118 1963 1124 1964
rect 1118 1959 1119 1963
rect 1123 1959 1124 1963
rect 1118 1958 1124 1959
rect 1238 1963 1244 1964
rect 1238 1959 1239 1963
rect 1243 1959 1244 1963
rect 1238 1958 1244 1959
rect 1358 1963 1364 1964
rect 1358 1959 1359 1963
rect 1363 1959 1364 1963
rect 1358 1958 1364 1959
rect 1478 1963 1484 1964
rect 1478 1959 1479 1963
rect 1483 1959 1484 1963
rect 1478 1958 1484 1959
rect 1598 1963 1604 1964
rect 1598 1959 1599 1963
rect 1603 1959 1604 1963
rect 1902 1963 1903 1967
rect 1907 1963 1908 1967
rect 1902 1962 1908 1963
rect 2158 1967 2164 1968
rect 2158 1963 2159 1967
rect 2163 1963 2164 1967
rect 2158 1962 2164 1963
rect 2398 1967 2404 1968
rect 2398 1963 2399 1967
rect 2403 1963 2404 1967
rect 2398 1962 2404 1963
rect 2614 1967 2620 1968
rect 2614 1963 2615 1967
rect 2619 1963 2620 1967
rect 2614 1962 2620 1963
rect 2814 1967 2820 1968
rect 2814 1963 2815 1967
rect 2819 1963 2820 1967
rect 2814 1962 2820 1963
rect 2998 1967 3004 1968
rect 2998 1963 2999 1967
rect 3003 1963 3004 1967
rect 2998 1962 3004 1963
rect 3166 1967 3172 1968
rect 3166 1963 3167 1967
rect 3171 1963 3172 1967
rect 3166 1962 3172 1963
rect 3334 1967 3340 1968
rect 3334 1963 3335 1967
rect 3339 1963 3340 1967
rect 3334 1962 3340 1963
rect 3478 1967 3484 1968
rect 3478 1963 3479 1967
rect 3483 1963 3484 1967
rect 3478 1962 3484 1963
rect 1598 1958 1604 1959
rect 1862 1957 1868 1958
rect 110 1953 116 1954
rect 110 1949 111 1953
rect 115 1949 116 1953
rect 110 1948 116 1949
rect 1822 1953 1828 1954
rect 1822 1949 1823 1953
rect 1827 1949 1828 1953
rect 1862 1953 1863 1957
rect 1867 1953 1868 1957
rect 1862 1952 1868 1953
rect 3574 1957 3580 1958
rect 3574 1953 3575 1957
rect 3579 1953 3580 1957
rect 3574 1952 3580 1953
rect 1822 1948 1828 1949
rect 1862 1940 1868 1941
rect 110 1936 116 1937
rect 110 1932 111 1936
rect 115 1932 116 1936
rect 110 1931 116 1932
rect 1822 1936 1828 1937
rect 1822 1932 1823 1936
rect 1827 1932 1828 1936
rect 1862 1936 1863 1940
rect 1867 1936 1868 1940
rect 1862 1935 1868 1936
rect 3574 1940 3580 1941
rect 3574 1936 3575 1940
rect 3579 1936 3580 1940
rect 3574 1935 3580 1936
rect 1822 1931 1828 1932
rect 1910 1927 1916 1928
rect 166 1923 172 1924
rect 166 1919 167 1923
rect 171 1919 172 1923
rect 166 1918 172 1919
rect 302 1923 308 1924
rect 302 1919 303 1923
rect 307 1919 308 1923
rect 302 1918 308 1919
rect 446 1923 452 1924
rect 446 1919 447 1923
rect 451 1919 452 1923
rect 446 1918 452 1919
rect 590 1923 596 1924
rect 590 1919 591 1923
rect 595 1919 596 1923
rect 590 1918 596 1919
rect 726 1923 732 1924
rect 726 1919 727 1923
rect 731 1919 732 1923
rect 726 1918 732 1919
rect 862 1923 868 1924
rect 862 1919 863 1923
rect 867 1919 868 1923
rect 862 1918 868 1919
rect 998 1923 1004 1924
rect 998 1919 999 1923
rect 1003 1919 1004 1923
rect 998 1918 1004 1919
rect 1126 1923 1132 1924
rect 1126 1919 1127 1923
rect 1131 1919 1132 1923
rect 1126 1918 1132 1919
rect 1246 1923 1252 1924
rect 1246 1919 1247 1923
rect 1251 1919 1252 1923
rect 1246 1918 1252 1919
rect 1366 1923 1372 1924
rect 1366 1919 1367 1923
rect 1371 1919 1372 1923
rect 1366 1918 1372 1919
rect 1486 1923 1492 1924
rect 1486 1919 1487 1923
rect 1491 1919 1492 1923
rect 1486 1918 1492 1919
rect 1606 1923 1612 1924
rect 1606 1919 1607 1923
rect 1611 1919 1612 1923
rect 1910 1923 1911 1927
rect 1915 1923 1916 1927
rect 1910 1922 1916 1923
rect 2166 1927 2172 1928
rect 2166 1923 2167 1927
rect 2171 1923 2172 1927
rect 2166 1922 2172 1923
rect 2406 1927 2412 1928
rect 2406 1923 2407 1927
rect 2411 1923 2412 1927
rect 2406 1922 2412 1923
rect 2622 1927 2628 1928
rect 2622 1923 2623 1927
rect 2627 1923 2628 1927
rect 2622 1922 2628 1923
rect 2822 1927 2828 1928
rect 2822 1923 2823 1927
rect 2827 1923 2828 1927
rect 2822 1922 2828 1923
rect 3006 1927 3012 1928
rect 3006 1923 3007 1927
rect 3011 1923 3012 1927
rect 3006 1922 3012 1923
rect 3174 1927 3180 1928
rect 3174 1923 3175 1927
rect 3179 1923 3180 1927
rect 3174 1922 3180 1923
rect 3342 1927 3348 1928
rect 3342 1923 3343 1927
rect 3347 1923 3348 1927
rect 3342 1922 3348 1923
rect 3486 1927 3492 1928
rect 3486 1923 3487 1927
rect 3491 1923 3492 1927
rect 3486 1922 3492 1923
rect 1606 1918 1612 1919
rect 1894 1893 1900 1894
rect 1894 1889 1895 1893
rect 1899 1889 1900 1893
rect 1894 1888 1900 1889
rect 1982 1893 1988 1894
rect 1982 1889 1983 1893
rect 1987 1889 1988 1893
rect 1982 1888 1988 1889
rect 2070 1893 2076 1894
rect 2070 1889 2071 1893
rect 2075 1889 2076 1893
rect 2070 1888 2076 1889
rect 2166 1893 2172 1894
rect 2166 1889 2167 1893
rect 2171 1889 2172 1893
rect 2166 1888 2172 1889
rect 2294 1893 2300 1894
rect 2294 1889 2295 1893
rect 2299 1889 2300 1893
rect 2294 1888 2300 1889
rect 2446 1893 2452 1894
rect 2446 1889 2447 1893
rect 2451 1889 2452 1893
rect 2446 1888 2452 1889
rect 2606 1893 2612 1894
rect 2606 1889 2607 1893
rect 2611 1889 2612 1893
rect 2606 1888 2612 1889
rect 2766 1893 2772 1894
rect 2766 1889 2767 1893
rect 2771 1889 2772 1893
rect 2766 1888 2772 1889
rect 2918 1893 2924 1894
rect 2918 1889 2919 1893
rect 2923 1889 2924 1893
rect 2918 1888 2924 1889
rect 3070 1893 3076 1894
rect 3070 1889 3071 1893
rect 3075 1889 3076 1893
rect 3070 1888 3076 1889
rect 3214 1893 3220 1894
rect 3214 1889 3215 1893
rect 3219 1889 3220 1893
rect 3214 1888 3220 1889
rect 3358 1893 3364 1894
rect 3358 1889 3359 1893
rect 3363 1889 3364 1893
rect 3358 1888 3364 1889
rect 3486 1893 3492 1894
rect 3486 1889 3487 1893
rect 3491 1889 3492 1893
rect 3486 1888 3492 1889
rect 222 1881 228 1882
rect 222 1877 223 1881
rect 227 1877 228 1881
rect 222 1876 228 1877
rect 478 1881 484 1882
rect 478 1877 479 1881
rect 483 1877 484 1881
rect 478 1876 484 1877
rect 718 1881 724 1882
rect 718 1877 719 1881
rect 723 1877 724 1881
rect 718 1876 724 1877
rect 934 1881 940 1882
rect 934 1877 935 1881
rect 939 1877 940 1881
rect 934 1876 940 1877
rect 1126 1881 1132 1882
rect 1126 1877 1127 1881
rect 1131 1877 1132 1881
rect 1126 1876 1132 1877
rect 1294 1881 1300 1882
rect 1294 1877 1295 1881
rect 1299 1877 1300 1881
rect 1294 1876 1300 1877
rect 1454 1881 1460 1882
rect 1454 1877 1455 1881
rect 1459 1877 1460 1881
rect 1454 1876 1460 1877
rect 1606 1881 1612 1882
rect 1606 1877 1607 1881
rect 1611 1877 1612 1881
rect 1606 1876 1612 1877
rect 1734 1881 1740 1882
rect 1734 1877 1735 1881
rect 1739 1877 1740 1881
rect 1734 1876 1740 1877
rect 1862 1880 1868 1881
rect 1862 1876 1863 1880
rect 1867 1876 1868 1880
rect 1862 1875 1868 1876
rect 3574 1880 3580 1881
rect 3574 1876 3575 1880
rect 3579 1876 3580 1880
rect 3574 1875 3580 1876
rect 110 1868 116 1869
rect 110 1864 111 1868
rect 115 1864 116 1868
rect 110 1863 116 1864
rect 1822 1868 1828 1869
rect 1822 1864 1823 1868
rect 1827 1864 1828 1868
rect 1822 1863 1828 1864
rect 1862 1863 1868 1864
rect 1862 1859 1863 1863
rect 1867 1859 1868 1863
rect 1862 1858 1868 1859
rect 3574 1863 3580 1864
rect 3574 1859 3575 1863
rect 3579 1859 3580 1863
rect 3574 1858 3580 1859
rect 1886 1853 1892 1854
rect 110 1851 116 1852
rect 110 1847 111 1851
rect 115 1847 116 1851
rect 110 1846 116 1847
rect 1822 1851 1828 1852
rect 1822 1847 1823 1851
rect 1827 1847 1828 1851
rect 1886 1849 1887 1853
rect 1891 1849 1892 1853
rect 1886 1848 1892 1849
rect 1974 1853 1980 1854
rect 1974 1849 1975 1853
rect 1979 1849 1980 1853
rect 1974 1848 1980 1849
rect 2062 1853 2068 1854
rect 2062 1849 2063 1853
rect 2067 1849 2068 1853
rect 2062 1848 2068 1849
rect 2158 1853 2164 1854
rect 2158 1849 2159 1853
rect 2163 1849 2164 1853
rect 2158 1848 2164 1849
rect 2286 1853 2292 1854
rect 2286 1849 2287 1853
rect 2291 1849 2292 1853
rect 2286 1848 2292 1849
rect 2438 1853 2444 1854
rect 2438 1849 2439 1853
rect 2443 1849 2444 1853
rect 2438 1848 2444 1849
rect 2598 1853 2604 1854
rect 2598 1849 2599 1853
rect 2603 1849 2604 1853
rect 2598 1848 2604 1849
rect 2758 1853 2764 1854
rect 2758 1849 2759 1853
rect 2763 1849 2764 1853
rect 2758 1848 2764 1849
rect 2910 1853 2916 1854
rect 2910 1849 2911 1853
rect 2915 1849 2916 1853
rect 2910 1848 2916 1849
rect 3062 1853 3068 1854
rect 3062 1849 3063 1853
rect 3067 1849 3068 1853
rect 3062 1848 3068 1849
rect 3206 1853 3212 1854
rect 3206 1849 3207 1853
rect 3211 1849 3212 1853
rect 3206 1848 3212 1849
rect 3350 1853 3356 1854
rect 3350 1849 3351 1853
rect 3355 1849 3356 1853
rect 3350 1848 3356 1849
rect 3478 1853 3484 1854
rect 3478 1849 3479 1853
rect 3483 1849 3484 1853
rect 3478 1848 3484 1849
rect 1822 1846 1828 1847
rect 214 1841 220 1842
rect 214 1837 215 1841
rect 219 1837 220 1841
rect 214 1836 220 1837
rect 470 1841 476 1842
rect 470 1837 471 1841
rect 475 1837 476 1841
rect 470 1836 476 1837
rect 710 1841 716 1842
rect 710 1837 711 1841
rect 715 1837 716 1841
rect 710 1836 716 1837
rect 926 1841 932 1842
rect 926 1837 927 1841
rect 931 1837 932 1841
rect 926 1836 932 1837
rect 1118 1841 1124 1842
rect 1118 1837 1119 1841
rect 1123 1837 1124 1841
rect 1118 1836 1124 1837
rect 1286 1841 1292 1842
rect 1286 1837 1287 1841
rect 1291 1837 1292 1841
rect 1286 1836 1292 1837
rect 1446 1841 1452 1842
rect 1446 1837 1447 1841
rect 1451 1837 1452 1841
rect 1446 1836 1452 1837
rect 1598 1841 1604 1842
rect 1598 1837 1599 1841
rect 1603 1837 1604 1841
rect 1598 1836 1604 1837
rect 1726 1841 1732 1842
rect 1726 1837 1727 1841
rect 1731 1837 1732 1841
rect 1726 1836 1732 1837
rect 1998 1827 2004 1828
rect 1998 1823 1999 1827
rect 2003 1823 2004 1827
rect 1998 1822 2004 1823
rect 2222 1827 2228 1828
rect 2222 1823 2223 1827
rect 2227 1823 2228 1827
rect 2222 1822 2228 1823
rect 2438 1827 2444 1828
rect 2438 1823 2439 1827
rect 2443 1823 2444 1827
rect 2438 1822 2444 1823
rect 2638 1827 2644 1828
rect 2638 1823 2639 1827
rect 2643 1823 2644 1827
rect 2638 1822 2644 1823
rect 2830 1827 2836 1828
rect 2830 1823 2831 1827
rect 2835 1823 2836 1827
rect 2830 1822 2836 1823
rect 3014 1827 3020 1828
rect 3014 1823 3015 1827
rect 3019 1823 3020 1827
rect 3014 1822 3020 1823
rect 3198 1827 3204 1828
rect 3198 1823 3199 1827
rect 3203 1823 3204 1827
rect 3198 1822 3204 1823
rect 3390 1827 3396 1828
rect 3390 1823 3391 1827
rect 3395 1823 3396 1827
rect 3390 1822 3396 1823
rect 246 1819 252 1820
rect 246 1815 247 1819
rect 251 1815 252 1819
rect 246 1814 252 1815
rect 414 1819 420 1820
rect 414 1815 415 1819
rect 419 1815 420 1819
rect 414 1814 420 1815
rect 590 1819 596 1820
rect 590 1815 591 1819
rect 595 1815 596 1819
rect 590 1814 596 1815
rect 758 1819 764 1820
rect 758 1815 759 1819
rect 763 1815 764 1819
rect 758 1814 764 1815
rect 926 1819 932 1820
rect 926 1815 927 1819
rect 931 1815 932 1819
rect 926 1814 932 1815
rect 1078 1819 1084 1820
rect 1078 1815 1079 1819
rect 1083 1815 1084 1819
rect 1078 1814 1084 1815
rect 1222 1819 1228 1820
rect 1222 1815 1223 1819
rect 1227 1815 1228 1819
rect 1222 1814 1228 1815
rect 1358 1819 1364 1820
rect 1358 1815 1359 1819
rect 1363 1815 1364 1819
rect 1358 1814 1364 1815
rect 1486 1819 1492 1820
rect 1486 1815 1487 1819
rect 1491 1815 1492 1819
rect 1486 1814 1492 1815
rect 1614 1819 1620 1820
rect 1614 1815 1615 1819
rect 1619 1815 1620 1819
rect 1614 1814 1620 1815
rect 1726 1819 1732 1820
rect 1726 1815 1727 1819
rect 1731 1815 1732 1819
rect 1726 1814 1732 1815
rect 1862 1817 1868 1818
rect 1862 1813 1863 1817
rect 1867 1813 1868 1817
rect 1862 1812 1868 1813
rect 3574 1817 3580 1818
rect 3574 1813 3575 1817
rect 3579 1813 3580 1817
rect 3574 1812 3580 1813
rect 110 1809 116 1810
rect 110 1805 111 1809
rect 115 1805 116 1809
rect 110 1804 116 1805
rect 1822 1809 1828 1810
rect 1822 1805 1823 1809
rect 1827 1805 1828 1809
rect 1822 1804 1828 1805
rect 1862 1800 1868 1801
rect 1862 1796 1863 1800
rect 1867 1796 1868 1800
rect 1862 1795 1868 1796
rect 3574 1800 3580 1801
rect 3574 1796 3575 1800
rect 3579 1796 3580 1800
rect 3574 1795 3580 1796
rect 110 1792 116 1793
rect 110 1788 111 1792
rect 115 1788 116 1792
rect 110 1787 116 1788
rect 1822 1792 1828 1793
rect 1822 1788 1823 1792
rect 1827 1788 1828 1792
rect 1822 1787 1828 1788
rect 2006 1787 2012 1788
rect 2006 1783 2007 1787
rect 2011 1783 2012 1787
rect 2006 1782 2012 1783
rect 2230 1787 2236 1788
rect 2230 1783 2231 1787
rect 2235 1783 2236 1787
rect 2230 1782 2236 1783
rect 2446 1787 2452 1788
rect 2446 1783 2447 1787
rect 2451 1783 2452 1787
rect 2446 1782 2452 1783
rect 2646 1787 2652 1788
rect 2646 1783 2647 1787
rect 2651 1783 2652 1787
rect 2646 1782 2652 1783
rect 2838 1787 2844 1788
rect 2838 1783 2839 1787
rect 2843 1783 2844 1787
rect 2838 1782 2844 1783
rect 3022 1787 3028 1788
rect 3022 1783 3023 1787
rect 3027 1783 3028 1787
rect 3022 1782 3028 1783
rect 3206 1787 3212 1788
rect 3206 1783 3207 1787
rect 3211 1783 3212 1787
rect 3206 1782 3212 1783
rect 3398 1787 3404 1788
rect 3398 1783 3399 1787
rect 3403 1783 3404 1787
rect 3398 1782 3404 1783
rect 254 1779 260 1780
rect 254 1775 255 1779
rect 259 1775 260 1779
rect 254 1774 260 1775
rect 422 1779 428 1780
rect 422 1775 423 1779
rect 427 1775 428 1779
rect 422 1774 428 1775
rect 598 1779 604 1780
rect 598 1775 599 1779
rect 603 1775 604 1779
rect 598 1774 604 1775
rect 766 1779 772 1780
rect 766 1775 767 1779
rect 771 1775 772 1779
rect 766 1774 772 1775
rect 934 1779 940 1780
rect 934 1775 935 1779
rect 939 1775 940 1779
rect 934 1774 940 1775
rect 1086 1779 1092 1780
rect 1086 1775 1087 1779
rect 1091 1775 1092 1779
rect 1086 1774 1092 1775
rect 1230 1779 1236 1780
rect 1230 1775 1231 1779
rect 1235 1775 1236 1779
rect 1230 1774 1236 1775
rect 1366 1779 1372 1780
rect 1366 1775 1367 1779
rect 1371 1775 1372 1779
rect 1366 1774 1372 1775
rect 1494 1779 1500 1780
rect 1494 1775 1495 1779
rect 1499 1775 1500 1779
rect 1494 1774 1500 1775
rect 1622 1779 1628 1780
rect 1622 1775 1623 1779
rect 1627 1775 1628 1779
rect 1622 1774 1628 1775
rect 1734 1779 1740 1780
rect 1734 1775 1735 1779
rect 1739 1775 1740 1779
rect 1734 1774 1740 1775
rect 1942 1749 1948 1750
rect 1942 1745 1943 1749
rect 1947 1745 1948 1749
rect 1942 1744 1948 1745
rect 2086 1749 2092 1750
rect 2086 1745 2087 1749
rect 2091 1745 2092 1749
rect 2086 1744 2092 1745
rect 2246 1749 2252 1750
rect 2246 1745 2247 1749
rect 2251 1745 2252 1749
rect 2246 1744 2252 1745
rect 2414 1749 2420 1750
rect 2414 1745 2415 1749
rect 2419 1745 2420 1749
rect 2414 1744 2420 1745
rect 2598 1749 2604 1750
rect 2598 1745 2599 1749
rect 2603 1745 2604 1749
rect 2598 1744 2604 1745
rect 2790 1749 2796 1750
rect 2790 1745 2791 1749
rect 2795 1745 2796 1749
rect 2790 1744 2796 1745
rect 2990 1749 2996 1750
rect 2990 1745 2991 1749
rect 2995 1745 2996 1749
rect 2990 1744 2996 1745
rect 3198 1749 3204 1750
rect 3198 1745 3199 1749
rect 3203 1745 3204 1749
rect 3198 1744 3204 1745
rect 3414 1749 3420 1750
rect 3414 1745 3415 1749
rect 3419 1745 3420 1749
rect 3414 1744 3420 1745
rect 326 1741 332 1742
rect 326 1737 327 1741
rect 331 1737 332 1741
rect 326 1736 332 1737
rect 470 1741 476 1742
rect 470 1737 471 1741
rect 475 1737 476 1741
rect 470 1736 476 1737
rect 614 1741 620 1742
rect 614 1737 615 1741
rect 619 1737 620 1741
rect 614 1736 620 1737
rect 766 1741 772 1742
rect 766 1737 767 1741
rect 771 1737 772 1741
rect 766 1736 772 1737
rect 918 1741 924 1742
rect 918 1737 919 1741
rect 923 1737 924 1741
rect 918 1736 924 1737
rect 1070 1741 1076 1742
rect 1070 1737 1071 1741
rect 1075 1737 1076 1741
rect 1070 1736 1076 1737
rect 1222 1741 1228 1742
rect 1222 1737 1223 1741
rect 1227 1737 1228 1741
rect 1222 1736 1228 1737
rect 1374 1741 1380 1742
rect 1374 1737 1375 1741
rect 1379 1737 1380 1741
rect 1374 1736 1380 1737
rect 1526 1741 1532 1742
rect 1526 1737 1527 1741
rect 1531 1737 1532 1741
rect 1526 1736 1532 1737
rect 1686 1741 1692 1742
rect 1686 1737 1687 1741
rect 1691 1737 1692 1741
rect 1686 1736 1692 1737
rect 1862 1736 1868 1737
rect 1862 1732 1863 1736
rect 1867 1732 1868 1736
rect 1862 1731 1868 1732
rect 3574 1736 3580 1737
rect 3574 1732 3575 1736
rect 3579 1732 3580 1736
rect 3574 1731 3580 1732
rect 110 1728 116 1729
rect 110 1724 111 1728
rect 115 1724 116 1728
rect 110 1723 116 1724
rect 1822 1728 1828 1729
rect 1822 1724 1823 1728
rect 1827 1724 1828 1728
rect 1822 1723 1828 1724
rect 1862 1719 1868 1720
rect 1862 1715 1863 1719
rect 1867 1715 1868 1719
rect 1862 1714 1868 1715
rect 3574 1719 3580 1720
rect 3574 1715 3575 1719
rect 3579 1715 3580 1719
rect 3574 1714 3580 1715
rect 110 1711 116 1712
rect 110 1707 111 1711
rect 115 1707 116 1711
rect 110 1706 116 1707
rect 1822 1711 1828 1712
rect 1822 1707 1823 1711
rect 1827 1707 1828 1711
rect 1822 1706 1828 1707
rect 1934 1709 1940 1710
rect 1934 1705 1935 1709
rect 1939 1705 1940 1709
rect 1934 1704 1940 1705
rect 2078 1709 2084 1710
rect 2078 1705 2079 1709
rect 2083 1705 2084 1709
rect 2078 1704 2084 1705
rect 2238 1709 2244 1710
rect 2238 1705 2239 1709
rect 2243 1705 2244 1709
rect 2238 1704 2244 1705
rect 2406 1709 2412 1710
rect 2406 1705 2407 1709
rect 2411 1705 2412 1709
rect 2406 1704 2412 1705
rect 2590 1709 2596 1710
rect 2590 1705 2591 1709
rect 2595 1705 2596 1709
rect 2590 1704 2596 1705
rect 2782 1709 2788 1710
rect 2782 1705 2783 1709
rect 2787 1705 2788 1709
rect 2782 1704 2788 1705
rect 2982 1709 2988 1710
rect 2982 1705 2983 1709
rect 2987 1705 2988 1709
rect 2982 1704 2988 1705
rect 3190 1709 3196 1710
rect 3190 1705 3191 1709
rect 3195 1705 3196 1709
rect 3190 1704 3196 1705
rect 3406 1709 3412 1710
rect 3406 1705 3407 1709
rect 3411 1705 3412 1709
rect 3406 1704 3412 1705
rect 318 1701 324 1702
rect 318 1697 319 1701
rect 323 1697 324 1701
rect 318 1696 324 1697
rect 462 1701 468 1702
rect 462 1697 463 1701
rect 467 1697 468 1701
rect 462 1696 468 1697
rect 606 1701 612 1702
rect 606 1697 607 1701
rect 611 1697 612 1701
rect 606 1696 612 1697
rect 758 1701 764 1702
rect 758 1697 759 1701
rect 763 1697 764 1701
rect 758 1696 764 1697
rect 910 1701 916 1702
rect 910 1697 911 1701
rect 915 1697 916 1701
rect 910 1696 916 1697
rect 1062 1701 1068 1702
rect 1062 1697 1063 1701
rect 1067 1697 1068 1701
rect 1062 1696 1068 1697
rect 1214 1701 1220 1702
rect 1214 1697 1215 1701
rect 1219 1697 1220 1701
rect 1214 1696 1220 1697
rect 1366 1701 1372 1702
rect 1366 1697 1367 1701
rect 1371 1697 1372 1701
rect 1366 1696 1372 1697
rect 1518 1701 1524 1702
rect 1518 1697 1519 1701
rect 1523 1697 1524 1701
rect 1518 1696 1524 1697
rect 1678 1701 1684 1702
rect 1678 1697 1679 1701
rect 1683 1697 1684 1701
rect 1678 1696 1684 1697
rect 1910 1683 1916 1684
rect 1910 1679 1911 1683
rect 1915 1679 1916 1683
rect 1910 1678 1916 1679
rect 2030 1683 2036 1684
rect 2030 1679 2031 1683
rect 2035 1679 2036 1683
rect 2030 1678 2036 1679
rect 2150 1683 2156 1684
rect 2150 1679 2151 1683
rect 2155 1679 2156 1683
rect 2150 1678 2156 1679
rect 2270 1683 2276 1684
rect 2270 1679 2271 1683
rect 2275 1679 2276 1683
rect 2270 1678 2276 1679
rect 2398 1683 2404 1684
rect 2398 1679 2399 1683
rect 2403 1679 2404 1683
rect 2398 1678 2404 1679
rect 2542 1683 2548 1684
rect 2542 1679 2543 1683
rect 2547 1679 2548 1683
rect 2542 1678 2548 1679
rect 2694 1683 2700 1684
rect 2694 1679 2695 1683
rect 2699 1679 2700 1683
rect 2694 1678 2700 1679
rect 2862 1683 2868 1684
rect 2862 1679 2863 1683
rect 2867 1679 2868 1683
rect 2862 1678 2868 1679
rect 3046 1683 3052 1684
rect 3046 1679 3047 1683
rect 3051 1679 3052 1683
rect 3046 1678 3052 1679
rect 3238 1683 3244 1684
rect 3238 1679 3239 1683
rect 3243 1679 3244 1683
rect 3238 1678 3244 1679
rect 3430 1683 3436 1684
rect 3430 1679 3431 1683
rect 3435 1679 3436 1683
rect 3430 1678 3436 1679
rect 310 1675 316 1676
rect 310 1671 311 1675
rect 315 1671 316 1675
rect 310 1670 316 1671
rect 446 1675 452 1676
rect 446 1671 447 1675
rect 451 1671 452 1675
rect 446 1670 452 1671
rect 590 1675 596 1676
rect 590 1671 591 1675
rect 595 1671 596 1675
rect 590 1670 596 1671
rect 734 1675 740 1676
rect 734 1671 735 1675
rect 739 1671 740 1675
rect 734 1670 740 1671
rect 886 1675 892 1676
rect 886 1671 887 1675
rect 891 1671 892 1675
rect 886 1670 892 1671
rect 1038 1675 1044 1676
rect 1038 1671 1039 1675
rect 1043 1671 1044 1675
rect 1038 1670 1044 1671
rect 1190 1675 1196 1676
rect 1190 1671 1191 1675
rect 1195 1671 1196 1675
rect 1190 1670 1196 1671
rect 1342 1675 1348 1676
rect 1342 1671 1343 1675
rect 1347 1671 1348 1675
rect 1342 1670 1348 1671
rect 1494 1675 1500 1676
rect 1494 1671 1495 1675
rect 1499 1671 1500 1675
rect 1494 1670 1500 1671
rect 1646 1675 1652 1676
rect 1646 1671 1647 1675
rect 1651 1671 1652 1675
rect 1646 1670 1652 1671
rect 1862 1673 1868 1674
rect 1862 1669 1863 1673
rect 1867 1669 1868 1673
rect 1862 1668 1868 1669
rect 3574 1673 3580 1674
rect 3574 1669 3575 1673
rect 3579 1669 3580 1673
rect 3574 1668 3580 1669
rect 110 1665 116 1666
rect 110 1661 111 1665
rect 115 1661 116 1665
rect 110 1660 116 1661
rect 1822 1665 1828 1666
rect 1822 1661 1823 1665
rect 1827 1661 1828 1665
rect 1822 1660 1828 1661
rect 1862 1656 1868 1657
rect 1862 1652 1863 1656
rect 1867 1652 1868 1656
rect 1862 1651 1868 1652
rect 3574 1656 3580 1657
rect 3574 1652 3575 1656
rect 3579 1652 3580 1656
rect 3574 1651 3580 1652
rect 110 1648 116 1649
rect 110 1644 111 1648
rect 115 1644 116 1648
rect 110 1643 116 1644
rect 1822 1648 1828 1649
rect 1822 1644 1823 1648
rect 1827 1644 1828 1648
rect 1822 1643 1828 1644
rect 1918 1643 1924 1644
rect 1918 1639 1919 1643
rect 1923 1639 1924 1643
rect 1918 1638 1924 1639
rect 2038 1643 2044 1644
rect 2038 1639 2039 1643
rect 2043 1639 2044 1643
rect 2038 1638 2044 1639
rect 2158 1643 2164 1644
rect 2158 1639 2159 1643
rect 2163 1639 2164 1643
rect 2158 1638 2164 1639
rect 2278 1643 2284 1644
rect 2278 1639 2279 1643
rect 2283 1639 2284 1643
rect 2278 1638 2284 1639
rect 2406 1643 2412 1644
rect 2406 1639 2407 1643
rect 2411 1639 2412 1643
rect 2406 1638 2412 1639
rect 2550 1643 2556 1644
rect 2550 1639 2551 1643
rect 2555 1639 2556 1643
rect 2550 1638 2556 1639
rect 2702 1643 2708 1644
rect 2702 1639 2703 1643
rect 2707 1639 2708 1643
rect 2702 1638 2708 1639
rect 2870 1643 2876 1644
rect 2870 1639 2871 1643
rect 2875 1639 2876 1643
rect 2870 1638 2876 1639
rect 3054 1643 3060 1644
rect 3054 1639 3055 1643
rect 3059 1639 3060 1643
rect 3054 1638 3060 1639
rect 3246 1643 3252 1644
rect 3246 1639 3247 1643
rect 3251 1639 3252 1643
rect 3246 1638 3252 1639
rect 3438 1643 3444 1644
rect 3438 1639 3439 1643
rect 3443 1639 3444 1643
rect 3438 1638 3444 1639
rect 318 1635 324 1636
rect 318 1631 319 1635
rect 323 1631 324 1635
rect 318 1630 324 1631
rect 454 1635 460 1636
rect 454 1631 455 1635
rect 459 1631 460 1635
rect 454 1630 460 1631
rect 598 1635 604 1636
rect 598 1631 599 1635
rect 603 1631 604 1635
rect 598 1630 604 1631
rect 742 1635 748 1636
rect 742 1631 743 1635
rect 747 1631 748 1635
rect 742 1630 748 1631
rect 894 1635 900 1636
rect 894 1631 895 1635
rect 899 1631 900 1635
rect 894 1630 900 1631
rect 1046 1635 1052 1636
rect 1046 1631 1047 1635
rect 1051 1631 1052 1635
rect 1046 1630 1052 1631
rect 1198 1635 1204 1636
rect 1198 1631 1199 1635
rect 1203 1631 1204 1635
rect 1198 1630 1204 1631
rect 1350 1635 1356 1636
rect 1350 1631 1351 1635
rect 1355 1631 1356 1635
rect 1350 1630 1356 1631
rect 1502 1635 1508 1636
rect 1502 1631 1503 1635
rect 1507 1631 1508 1635
rect 1502 1630 1508 1631
rect 1654 1635 1660 1636
rect 1654 1631 1655 1635
rect 1659 1631 1660 1635
rect 1654 1630 1660 1631
rect 1894 1601 1900 1602
rect 1894 1597 1895 1601
rect 1899 1597 1900 1601
rect 1894 1596 1900 1597
rect 2014 1601 2020 1602
rect 2014 1597 2015 1601
rect 2019 1597 2020 1601
rect 2014 1596 2020 1597
rect 2150 1601 2156 1602
rect 2150 1597 2151 1601
rect 2155 1597 2156 1601
rect 2150 1596 2156 1597
rect 2286 1601 2292 1602
rect 2286 1597 2287 1601
rect 2291 1597 2292 1601
rect 2286 1596 2292 1597
rect 2430 1601 2436 1602
rect 2430 1597 2431 1601
rect 2435 1597 2436 1601
rect 2430 1596 2436 1597
rect 2582 1601 2588 1602
rect 2582 1597 2583 1601
rect 2587 1597 2588 1601
rect 2582 1596 2588 1597
rect 2742 1601 2748 1602
rect 2742 1597 2743 1601
rect 2747 1597 2748 1601
rect 2742 1596 2748 1597
rect 2910 1601 2916 1602
rect 2910 1597 2911 1601
rect 2915 1597 2916 1601
rect 2910 1596 2916 1597
rect 3094 1601 3100 1602
rect 3094 1597 3095 1601
rect 3099 1597 3100 1601
rect 3094 1596 3100 1597
rect 3278 1601 3284 1602
rect 3278 1597 3279 1601
rect 3283 1597 3284 1601
rect 3278 1596 3284 1597
rect 3470 1601 3476 1602
rect 3470 1597 3471 1601
rect 3475 1597 3476 1601
rect 3470 1596 3476 1597
rect 222 1593 228 1594
rect 222 1589 223 1593
rect 227 1589 228 1593
rect 222 1588 228 1589
rect 350 1593 356 1594
rect 350 1589 351 1593
rect 355 1589 356 1593
rect 350 1588 356 1589
rect 486 1593 492 1594
rect 486 1589 487 1593
rect 491 1589 492 1593
rect 486 1588 492 1589
rect 622 1593 628 1594
rect 622 1589 623 1593
rect 627 1589 628 1593
rect 622 1588 628 1589
rect 758 1593 764 1594
rect 758 1589 759 1593
rect 763 1589 764 1593
rect 758 1588 764 1589
rect 902 1593 908 1594
rect 902 1589 903 1593
rect 907 1589 908 1593
rect 902 1588 908 1589
rect 1054 1593 1060 1594
rect 1054 1589 1055 1593
rect 1059 1589 1060 1593
rect 1054 1588 1060 1589
rect 1214 1593 1220 1594
rect 1214 1589 1215 1593
rect 1219 1589 1220 1593
rect 1214 1588 1220 1589
rect 1374 1593 1380 1594
rect 1374 1589 1375 1593
rect 1379 1589 1380 1593
rect 1374 1588 1380 1589
rect 1542 1593 1548 1594
rect 1542 1589 1543 1593
rect 1547 1589 1548 1593
rect 1542 1588 1548 1589
rect 1862 1588 1868 1589
rect 1862 1584 1863 1588
rect 1867 1584 1868 1588
rect 1862 1583 1868 1584
rect 3574 1588 3580 1589
rect 3574 1584 3575 1588
rect 3579 1584 3580 1588
rect 3574 1583 3580 1584
rect 110 1580 116 1581
rect 110 1576 111 1580
rect 115 1576 116 1580
rect 110 1575 116 1576
rect 1822 1580 1828 1581
rect 1822 1576 1823 1580
rect 1827 1576 1828 1580
rect 1822 1575 1828 1576
rect 1862 1571 1868 1572
rect 1862 1567 1863 1571
rect 1867 1567 1868 1571
rect 1862 1566 1868 1567
rect 3574 1571 3580 1572
rect 3574 1567 3575 1571
rect 3579 1567 3580 1571
rect 3574 1566 3580 1567
rect 110 1563 116 1564
rect 110 1559 111 1563
rect 115 1559 116 1563
rect 110 1558 116 1559
rect 1822 1563 1828 1564
rect 1822 1559 1823 1563
rect 1827 1559 1828 1563
rect 1822 1558 1828 1559
rect 1886 1561 1892 1562
rect 1886 1557 1887 1561
rect 1891 1557 1892 1561
rect 1886 1556 1892 1557
rect 2006 1561 2012 1562
rect 2006 1557 2007 1561
rect 2011 1557 2012 1561
rect 2006 1556 2012 1557
rect 2142 1561 2148 1562
rect 2142 1557 2143 1561
rect 2147 1557 2148 1561
rect 2142 1556 2148 1557
rect 2278 1561 2284 1562
rect 2278 1557 2279 1561
rect 2283 1557 2284 1561
rect 2278 1556 2284 1557
rect 2422 1561 2428 1562
rect 2422 1557 2423 1561
rect 2427 1557 2428 1561
rect 2422 1556 2428 1557
rect 2574 1561 2580 1562
rect 2574 1557 2575 1561
rect 2579 1557 2580 1561
rect 2574 1556 2580 1557
rect 2734 1561 2740 1562
rect 2734 1557 2735 1561
rect 2739 1557 2740 1561
rect 2734 1556 2740 1557
rect 2902 1561 2908 1562
rect 2902 1557 2903 1561
rect 2907 1557 2908 1561
rect 2902 1556 2908 1557
rect 3086 1561 3092 1562
rect 3086 1557 3087 1561
rect 3091 1557 3092 1561
rect 3086 1556 3092 1557
rect 3270 1561 3276 1562
rect 3270 1557 3271 1561
rect 3275 1557 3276 1561
rect 3270 1556 3276 1557
rect 3462 1561 3468 1562
rect 3462 1557 3463 1561
rect 3467 1557 3468 1561
rect 3462 1556 3468 1557
rect 214 1553 220 1554
rect 214 1549 215 1553
rect 219 1549 220 1553
rect 214 1548 220 1549
rect 342 1553 348 1554
rect 342 1549 343 1553
rect 347 1549 348 1553
rect 342 1548 348 1549
rect 478 1553 484 1554
rect 478 1549 479 1553
rect 483 1549 484 1553
rect 478 1548 484 1549
rect 614 1553 620 1554
rect 614 1549 615 1553
rect 619 1549 620 1553
rect 614 1548 620 1549
rect 750 1553 756 1554
rect 750 1549 751 1553
rect 755 1549 756 1553
rect 750 1548 756 1549
rect 894 1553 900 1554
rect 894 1549 895 1553
rect 899 1549 900 1553
rect 894 1548 900 1549
rect 1046 1553 1052 1554
rect 1046 1549 1047 1553
rect 1051 1549 1052 1553
rect 1046 1548 1052 1549
rect 1206 1553 1212 1554
rect 1206 1549 1207 1553
rect 1211 1549 1212 1553
rect 1206 1548 1212 1549
rect 1366 1553 1372 1554
rect 1366 1549 1367 1553
rect 1371 1549 1372 1553
rect 1366 1548 1372 1549
rect 1534 1553 1540 1554
rect 1534 1549 1535 1553
rect 1539 1549 1540 1553
rect 1534 1548 1540 1549
rect 1886 1531 1892 1532
rect 134 1527 140 1528
rect 134 1523 135 1527
rect 139 1523 140 1527
rect 134 1522 140 1523
rect 270 1527 276 1528
rect 270 1523 271 1527
rect 275 1523 276 1527
rect 270 1522 276 1523
rect 422 1527 428 1528
rect 422 1523 423 1527
rect 427 1523 428 1527
rect 422 1522 428 1523
rect 582 1527 588 1528
rect 582 1523 583 1527
rect 587 1523 588 1527
rect 582 1522 588 1523
rect 734 1527 740 1528
rect 734 1523 735 1527
rect 739 1523 740 1527
rect 734 1522 740 1523
rect 886 1527 892 1528
rect 886 1523 887 1527
rect 891 1523 892 1527
rect 886 1522 892 1523
rect 1038 1527 1044 1528
rect 1038 1523 1039 1527
rect 1043 1523 1044 1527
rect 1038 1522 1044 1523
rect 1190 1527 1196 1528
rect 1190 1523 1191 1527
rect 1195 1523 1196 1527
rect 1190 1522 1196 1523
rect 1342 1527 1348 1528
rect 1342 1523 1343 1527
rect 1347 1523 1348 1527
rect 1342 1522 1348 1523
rect 1494 1527 1500 1528
rect 1494 1523 1495 1527
rect 1499 1523 1500 1527
rect 1886 1527 1887 1531
rect 1891 1527 1892 1531
rect 1886 1526 1892 1527
rect 2022 1531 2028 1532
rect 2022 1527 2023 1531
rect 2027 1527 2028 1531
rect 2022 1526 2028 1527
rect 2182 1531 2188 1532
rect 2182 1527 2183 1531
rect 2187 1527 2188 1531
rect 2182 1526 2188 1527
rect 2342 1531 2348 1532
rect 2342 1527 2343 1531
rect 2347 1527 2348 1531
rect 2342 1526 2348 1527
rect 2502 1531 2508 1532
rect 2502 1527 2503 1531
rect 2507 1527 2508 1531
rect 2502 1526 2508 1527
rect 2662 1531 2668 1532
rect 2662 1527 2663 1531
rect 2667 1527 2668 1531
rect 2662 1526 2668 1527
rect 2822 1531 2828 1532
rect 2822 1527 2823 1531
rect 2827 1527 2828 1531
rect 2822 1526 2828 1527
rect 2982 1531 2988 1532
rect 2982 1527 2983 1531
rect 2987 1527 2988 1531
rect 2982 1526 2988 1527
rect 3150 1531 3156 1532
rect 3150 1527 3151 1531
rect 3155 1527 3156 1531
rect 3150 1526 3156 1527
rect 3318 1531 3324 1532
rect 3318 1527 3319 1531
rect 3323 1527 3324 1531
rect 3318 1526 3324 1527
rect 3478 1531 3484 1532
rect 3478 1527 3479 1531
rect 3483 1527 3484 1531
rect 3478 1526 3484 1527
rect 1494 1522 1500 1523
rect 1862 1521 1868 1522
rect 110 1517 116 1518
rect 110 1513 111 1517
rect 115 1513 116 1517
rect 110 1512 116 1513
rect 1822 1517 1828 1518
rect 1822 1513 1823 1517
rect 1827 1513 1828 1517
rect 1862 1517 1863 1521
rect 1867 1517 1868 1521
rect 1862 1516 1868 1517
rect 3574 1521 3580 1522
rect 3574 1517 3575 1521
rect 3579 1517 3580 1521
rect 3574 1516 3580 1517
rect 1822 1512 1828 1513
rect 1862 1504 1868 1505
rect 110 1500 116 1501
rect 110 1496 111 1500
rect 115 1496 116 1500
rect 110 1495 116 1496
rect 1822 1500 1828 1501
rect 1822 1496 1823 1500
rect 1827 1496 1828 1500
rect 1862 1500 1863 1504
rect 1867 1500 1868 1504
rect 1862 1499 1868 1500
rect 3574 1504 3580 1505
rect 3574 1500 3575 1504
rect 3579 1500 3580 1504
rect 3574 1499 3580 1500
rect 1822 1495 1828 1496
rect 1894 1491 1900 1492
rect 142 1487 148 1488
rect 142 1483 143 1487
rect 147 1483 148 1487
rect 142 1482 148 1483
rect 278 1487 284 1488
rect 278 1483 279 1487
rect 283 1483 284 1487
rect 278 1482 284 1483
rect 430 1487 436 1488
rect 430 1483 431 1487
rect 435 1483 436 1487
rect 430 1482 436 1483
rect 590 1487 596 1488
rect 590 1483 591 1487
rect 595 1483 596 1487
rect 590 1482 596 1483
rect 742 1487 748 1488
rect 742 1483 743 1487
rect 747 1483 748 1487
rect 742 1482 748 1483
rect 894 1487 900 1488
rect 894 1483 895 1487
rect 899 1483 900 1487
rect 894 1482 900 1483
rect 1046 1487 1052 1488
rect 1046 1483 1047 1487
rect 1051 1483 1052 1487
rect 1046 1482 1052 1483
rect 1198 1487 1204 1488
rect 1198 1483 1199 1487
rect 1203 1483 1204 1487
rect 1198 1482 1204 1483
rect 1350 1487 1356 1488
rect 1350 1483 1351 1487
rect 1355 1483 1356 1487
rect 1350 1482 1356 1483
rect 1502 1487 1508 1488
rect 1502 1483 1503 1487
rect 1507 1483 1508 1487
rect 1894 1487 1895 1491
rect 1899 1487 1900 1491
rect 1894 1486 1900 1487
rect 2030 1491 2036 1492
rect 2030 1487 2031 1491
rect 2035 1487 2036 1491
rect 2030 1486 2036 1487
rect 2190 1491 2196 1492
rect 2190 1487 2191 1491
rect 2195 1487 2196 1491
rect 2190 1486 2196 1487
rect 2350 1491 2356 1492
rect 2350 1487 2351 1491
rect 2355 1487 2356 1491
rect 2350 1486 2356 1487
rect 2510 1491 2516 1492
rect 2510 1487 2511 1491
rect 2515 1487 2516 1491
rect 2510 1486 2516 1487
rect 2670 1491 2676 1492
rect 2670 1487 2671 1491
rect 2675 1487 2676 1491
rect 2670 1486 2676 1487
rect 2830 1491 2836 1492
rect 2830 1487 2831 1491
rect 2835 1487 2836 1491
rect 2830 1486 2836 1487
rect 2990 1491 2996 1492
rect 2990 1487 2991 1491
rect 2995 1487 2996 1491
rect 2990 1486 2996 1487
rect 3158 1491 3164 1492
rect 3158 1487 3159 1491
rect 3163 1487 3164 1491
rect 3158 1486 3164 1487
rect 3326 1491 3332 1492
rect 3326 1487 3327 1491
rect 3331 1487 3332 1491
rect 3326 1486 3332 1487
rect 3486 1491 3492 1492
rect 3486 1487 3487 1491
rect 3491 1487 3492 1491
rect 3486 1486 3492 1487
rect 1502 1482 1508 1483
rect 2182 1449 2188 1450
rect 142 1445 148 1446
rect 142 1441 143 1445
rect 147 1441 148 1445
rect 142 1440 148 1441
rect 262 1445 268 1446
rect 262 1441 263 1445
rect 267 1441 268 1445
rect 262 1440 268 1441
rect 398 1445 404 1446
rect 398 1441 399 1445
rect 403 1441 404 1445
rect 398 1440 404 1441
rect 534 1445 540 1446
rect 534 1441 535 1445
rect 539 1441 540 1445
rect 534 1440 540 1441
rect 662 1445 668 1446
rect 662 1441 663 1445
rect 667 1441 668 1445
rect 662 1440 668 1441
rect 790 1445 796 1446
rect 790 1441 791 1445
rect 795 1441 796 1445
rect 790 1440 796 1441
rect 910 1445 916 1446
rect 910 1441 911 1445
rect 915 1441 916 1445
rect 910 1440 916 1441
rect 1022 1445 1028 1446
rect 1022 1441 1023 1445
rect 1027 1441 1028 1445
rect 1022 1440 1028 1441
rect 1142 1445 1148 1446
rect 1142 1441 1143 1445
rect 1147 1441 1148 1445
rect 1142 1440 1148 1441
rect 1262 1445 1268 1446
rect 1262 1441 1263 1445
rect 1267 1441 1268 1445
rect 1262 1440 1268 1441
rect 1382 1445 1388 1446
rect 1382 1441 1383 1445
rect 1387 1441 1388 1445
rect 1382 1440 1388 1441
rect 1502 1445 1508 1446
rect 1502 1441 1503 1445
rect 1507 1441 1508 1445
rect 1502 1440 1508 1441
rect 1630 1445 1636 1446
rect 1630 1441 1631 1445
rect 1635 1441 1636 1445
rect 1630 1440 1636 1441
rect 1734 1445 1740 1446
rect 1734 1441 1735 1445
rect 1739 1441 1740 1445
rect 2182 1445 2183 1449
rect 2187 1445 2188 1449
rect 2182 1444 2188 1445
rect 2358 1449 2364 1450
rect 2358 1445 2359 1449
rect 2363 1445 2364 1449
rect 2358 1444 2364 1445
rect 2526 1449 2532 1450
rect 2526 1445 2527 1449
rect 2531 1445 2532 1449
rect 2526 1444 2532 1445
rect 2686 1449 2692 1450
rect 2686 1445 2687 1449
rect 2691 1445 2692 1449
rect 2686 1444 2692 1445
rect 2846 1449 2852 1450
rect 2846 1445 2847 1449
rect 2851 1445 2852 1449
rect 2846 1444 2852 1445
rect 3006 1449 3012 1450
rect 3006 1445 3007 1449
rect 3011 1445 3012 1449
rect 3006 1444 3012 1445
rect 3174 1449 3180 1450
rect 3174 1445 3175 1449
rect 3179 1445 3180 1449
rect 3174 1444 3180 1445
rect 3342 1449 3348 1450
rect 3342 1445 3343 1449
rect 3347 1445 3348 1449
rect 3342 1444 3348 1445
rect 3486 1449 3492 1450
rect 3486 1445 3487 1449
rect 3491 1445 3492 1449
rect 3486 1444 3492 1445
rect 1734 1440 1740 1441
rect 1862 1436 1868 1437
rect 110 1432 116 1433
rect 110 1428 111 1432
rect 115 1428 116 1432
rect 110 1427 116 1428
rect 1822 1432 1828 1433
rect 1822 1428 1823 1432
rect 1827 1428 1828 1432
rect 1862 1432 1863 1436
rect 1867 1432 1868 1436
rect 1862 1431 1868 1432
rect 3574 1436 3580 1437
rect 3574 1432 3575 1436
rect 3579 1432 3580 1436
rect 3574 1431 3580 1432
rect 1822 1427 1828 1428
rect 1862 1419 1868 1420
rect 110 1415 116 1416
rect 110 1411 111 1415
rect 115 1411 116 1415
rect 110 1410 116 1411
rect 1822 1415 1828 1416
rect 1822 1411 1823 1415
rect 1827 1411 1828 1415
rect 1862 1415 1863 1419
rect 1867 1415 1868 1419
rect 1862 1414 1868 1415
rect 3574 1419 3580 1420
rect 3574 1415 3575 1419
rect 3579 1415 3580 1419
rect 3574 1414 3580 1415
rect 1822 1410 1828 1411
rect 2174 1409 2180 1410
rect 134 1405 140 1406
rect 134 1401 135 1405
rect 139 1401 140 1405
rect 134 1400 140 1401
rect 254 1405 260 1406
rect 254 1401 255 1405
rect 259 1401 260 1405
rect 254 1400 260 1401
rect 390 1405 396 1406
rect 390 1401 391 1405
rect 395 1401 396 1405
rect 390 1400 396 1401
rect 526 1405 532 1406
rect 526 1401 527 1405
rect 531 1401 532 1405
rect 526 1400 532 1401
rect 654 1405 660 1406
rect 654 1401 655 1405
rect 659 1401 660 1405
rect 654 1400 660 1401
rect 782 1405 788 1406
rect 782 1401 783 1405
rect 787 1401 788 1405
rect 782 1400 788 1401
rect 902 1405 908 1406
rect 902 1401 903 1405
rect 907 1401 908 1405
rect 902 1400 908 1401
rect 1014 1405 1020 1406
rect 1014 1401 1015 1405
rect 1019 1401 1020 1405
rect 1014 1400 1020 1401
rect 1134 1405 1140 1406
rect 1134 1401 1135 1405
rect 1139 1401 1140 1405
rect 1134 1400 1140 1401
rect 1254 1405 1260 1406
rect 1254 1401 1255 1405
rect 1259 1401 1260 1405
rect 1254 1400 1260 1401
rect 1374 1405 1380 1406
rect 1374 1401 1375 1405
rect 1379 1401 1380 1405
rect 1374 1400 1380 1401
rect 1494 1405 1500 1406
rect 1494 1401 1495 1405
rect 1499 1401 1500 1405
rect 1494 1400 1500 1401
rect 1622 1405 1628 1406
rect 1622 1401 1623 1405
rect 1627 1401 1628 1405
rect 1622 1400 1628 1401
rect 1726 1405 1732 1406
rect 1726 1401 1727 1405
rect 1731 1401 1732 1405
rect 2174 1405 2175 1409
rect 2179 1405 2180 1409
rect 2174 1404 2180 1405
rect 2350 1409 2356 1410
rect 2350 1405 2351 1409
rect 2355 1405 2356 1409
rect 2350 1404 2356 1405
rect 2518 1409 2524 1410
rect 2518 1405 2519 1409
rect 2523 1405 2524 1409
rect 2518 1404 2524 1405
rect 2678 1409 2684 1410
rect 2678 1405 2679 1409
rect 2683 1405 2684 1409
rect 2678 1404 2684 1405
rect 2838 1409 2844 1410
rect 2838 1405 2839 1409
rect 2843 1405 2844 1409
rect 2838 1404 2844 1405
rect 2998 1409 3004 1410
rect 2998 1405 2999 1409
rect 3003 1405 3004 1409
rect 2998 1404 3004 1405
rect 3166 1409 3172 1410
rect 3166 1405 3167 1409
rect 3171 1405 3172 1409
rect 3166 1404 3172 1405
rect 3334 1409 3340 1410
rect 3334 1405 3335 1409
rect 3339 1405 3340 1409
rect 3334 1404 3340 1405
rect 3478 1409 3484 1410
rect 3478 1405 3479 1409
rect 3483 1405 3484 1409
rect 3478 1404 3484 1405
rect 1726 1400 1732 1401
rect 134 1383 140 1384
rect 134 1379 135 1383
rect 139 1379 140 1383
rect 134 1378 140 1379
rect 326 1383 332 1384
rect 326 1379 327 1383
rect 331 1379 332 1383
rect 326 1378 332 1379
rect 550 1383 556 1384
rect 550 1379 551 1383
rect 555 1379 556 1383
rect 550 1378 556 1379
rect 782 1383 788 1384
rect 782 1379 783 1383
rect 787 1379 788 1383
rect 782 1378 788 1379
rect 1022 1383 1028 1384
rect 1022 1379 1023 1383
rect 1027 1379 1028 1383
rect 1022 1378 1028 1379
rect 1262 1383 1268 1384
rect 1262 1379 1263 1383
rect 1267 1379 1268 1383
rect 1262 1378 1268 1379
rect 1502 1383 1508 1384
rect 1502 1379 1503 1383
rect 1507 1379 1508 1383
rect 1502 1378 1508 1379
rect 1726 1383 1732 1384
rect 1726 1379 1727 1383
rect 1731 1379 1732 1383
rect 1726 1378 1732 1379
rect 2078 1379 2084 1380
rect 2078 1375 2079 1379
rect 2083 1375 2084 1379
rect 2078 1374 2084 1375
rect 2262 1379 2268 1380
rect 2262 1375 2263 1379
rect 2267 1375 2268 1379
rect 2262 1374 2268 1375
rect 2438 1379 2444 1380
rect 2438 1375 2439 1379
rect 2443 1375 2444 1379
rect 2438 1374 2444 1375
rect 2614 1379 2620 1380
rect 2614 1375 2615 1379
rect 2619 1375 2620 1379
rect 2614 1374 2620 1375
rect 2782 1379 2788 1380
rect 2782 1375 2783 1379
rect 2787 1375 2788 1379
rect 2782 1374 2788 1375
rect 2934 1379 2940 1380
rect 2934 1375 2935 1379
rect 2939 1375 2940 1379
rect 2934 1374 2940 1375
rect 3078 1379 3084 1380
rect 3078 1375 3079 1379
rect 3083 1375 3084 1379
rect 3078 1374 3084 1375
rect 3222 1379 3228 1380
rect 3222 1375 3223 1379
rect 3227 1375 3228 1379
rect 3222 1374 3228 1375
rect 3358 1379 3364 1380
rect 3358 1375 3359 1379
rect 3363 1375 3364 1379
rect 3358 1374 3364 1375
rect 3478 1379 3484 1380
rect 3478 1375 3479 1379
rect 3483 1375 3484 1379
rect 3478 1374 3484 1375
rect 110 1373 116 1374
rect 110 1369 111 1373
rect 115 1369 116 1373
rect 110 1368 116 1369
rect 1822 1373 1828 1374
rect 1822 1369 1823 1373
rect 1827 1369 1828 1373
rect 1822 1368 1828 1369
rect 1862 1369 1868 1370
rect 1862 1365 1863 1369
rect 1867 1365 1868 1369
rect 1862 1364 1868 1365
rect 3574 1369 3580 1370
rect 3574 1365 3575 1369
rect 3579 1365 3580 1369
rect 3574 1364 3580 1365
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 110 1351 116 1352
rect 1822 1356 1828 1357
rect 1822 1352 1823 1356
rect 1827 1352 1828 1356
rect 1822 1351 1828 1352
rect 1862 1352 1868 1353
rect 1862 1348 1863 1352
rect 1867 1348 1868 1352
rect 1862 1347 1868 1348
rect 3574 1352 3580 1353
rect 3574 1348 3575 1352
rect 3579 1348 3580 1352
rect 3574 1347 3580 1348
rect 142 1343 148 1344
rect 142 1339 143 1343
rect 147 1339 148 1343
rect 142 1338 148 1339
rect 334 1343 340 1344
rect 334 1339 335 1343
rect 339 1339 340 1343
rect 334 1338 340 1339
rect 558 1343 564 1344
rect 558 1339 559 1343
rect 563 1339 564 1343
rect 558 1338 564 1339
rect 790 1343 796 1344
rect 790 1339 791 1343
rect 795 1339 796 1343
rect 790 1338 796 1339
rect 1030 1343 1036 1344
rect 1030 1339 1031 1343
rect 1035 1339 1036 1343
rect 1030 1338 1036 1339
rect 1270 1343 1276 1344
rect 1270 1339 1271 1343
rect 1275 1339 1276 1343
rect 1270 1338 1276 1339
rect 1510 1343 1516 1344
rect 1510 1339 1511 1343
rect 1515 1339 1516 1343
rect 1510 1338 1516 1339
rect 1734 1343 1740 1344
rect 1734 1339 1735 1343
rect 1739 1339 1740 1343
rect 1734 1338 1740 1339
rect 2086 1339 2092 1340
rect 2086 1335 2087 1339
rect 2091 1335 2092 1339
rect 2086 1334 2092 1335
rect 2270 1339 2276 1340
rect 2270 1335 2271 1339
rect 2275 1335 2276 1339
rect 2270 1334 2276 1335
rect 2446 1339 2452 1340
rect 2446 1335 2447 1339
rect 2451 1335 2452 1339
rect 2446 1334 2452 1335
rect 2622 1339 2628 1340
rect 2622 1335 2623 1339
rect 2627 1335 2628 1339
rect 2622 1334 2628 1335
rect 2790 1339 2796 1340
rect 2790 1335 2791 1339
rect 2795 1335 2796 1339
rect 2790 1334 2796 1335
rect 2942 1339 2948 1340
rect 2942 1335 2943 1339
rect 2947 1335 2948 1339
rect 2942 1334 2948 1335
rect 3086 1339 3092 1340
rect 3086 1335 3087 1339
rect 3091 1335 3092 1339
rect 3086 1334 3092 1335
rect 3230 1339 3236 1340
rect 3230 1335 3231 1339
rect 3235 1335 3236 1339
rect 3230 1334 3236 1335
rect 3366 1339 3372 1340
rect 3366 1335 3367 1339
rect 3371 1335 3372 1339
rect 3366 1334 3372 1335
rect 3486 1339 3492 1340
rect 3486 1335 3487 1339
rect 3491 1335 3492 1339
rect 3486 1334 3492 1335
rect 2086 1305 2092 1306
rect 142 1301 148 1302
rect 142 1297 143 1301
rect 147 1297 148 1301
rect 142 1296 148 1297
rect 326 1301 332 1302
rect 326 1297 327 1301
rect 331 1297 332 1301
rect 326 1296 332 1297
rect 526 1301 532 1302
rect 526 1297 527 1301
rect 531 1297 532 1301
rect 526 1296 532 1297
rect 718 1301 724 1302
rect 718 1297 719 1301
rect 723 1297 724 1301
rect 718 1296 724 1297
rect 902 1301 908 1302
rect 902 1297 903 1301
rect 907 1297 908 1301
rect 902 1296 908 1297
rect 1070 1301 1076 1302
rect 1070 1297 1071 1301
rect 1075 1297 1076 1301
rect 1070 1296 1076 1297
rect 1230 1301 1236 1302
rect 1230 1297 1231 1301
rect 1235 1297 1236 1301
rect 1230 1296 1236 1297
rect 1382 1301 1388 1302
rect 1382 1297 1383 1301
rect 1387 1297 1388 1301
rect 1382 1296 1388 1297
rect 1534 1301 1540 1302
rect 1534 1297 1535 1301
rect 1539 1297 1540 1301
rect 1534 1296 1540 1297
rect 1686 1301 1692 1302
rect 1686 1297 1687 1301
rect 1691 1297 1692 1301
rect 2086 1301 2087 1305
rect 2091 1301 2092 1305
rect 2086 1300 2092 1301
rect 2310 1305 2316 1306
rect 2310 1301 2311 1305
rect 2315 1301 2316 1305
rect 2310 1300 2316 1301
rect 2518 1305 2524 1306
rect 2518 1301 2519 1305
rect 2523 1301 2524 1305
rect 2518 1300 2524 1301
rect 2710 1305 2716 1306
rect 2710 1301 2711 1305
rect 2715 1301 2716 1305
rect 2710 1300 2716 1301
rect 2886 1305 2892 1306
rect 2886 1301 2887 1305
rect 2891 1301 2892 1305
rect 2886 1300 2892 1301
rect 3046 1305 3052 1306
rect 3046 1301 3047 1305
rect 3051 1301 3052 1305
rect 3046 1300 3052 1301
rect 3198 1305 3204 1306
rect 3198 1301 3199 1305
rect 3203 1301 3204 1305
rect 3198 1300 3204 1301
rect 3350 1305 3356 1306
rect 3350 1301 3351 1305
rect 3355 1301 3356 1305
rect 3350 1300 3356 1301
rect 3486 1305 3492 1306
rect 3486 1301 3487 1305
rect 3491 1301 3492 1305
rect 3486 1300 3492 1301
rect 1686 1296 1692 1297
rect 1862 1292 1868 1293
rect 110 1288 116 1289
rect 110 1284 111 1288
rect 115 1284 116 1288
rect 110 1283 116 1284
rect 1822 1288 1828 1289
rect 1822 1284 1823 1288
rect 1827 1284 1828 1288
rect 1862 1288 1863 1292
rect 1867 1288 1868 1292
rect 1862 1287 1868 1288
rect 3574 1292 3580 1293
rect 3574 1288 3575 1292
rect 3579 1288 3580 1292
rect 3574 1287 3580 1288
rect 1822 1283 1828 1284
rect 1862 1275 1868 1276
rect 110 1271 116 1272
rect 110 1267 111 1271
rect 115 1267 116 1271
rect 110 1266 116 1267
rect 1822 1271 1828 1272
rect 1822 1267 1823 1271
rect 1827 1267 1828 1271
rect 1862 1271 1863 1275
rect 1867 1271 1868 1275
rect 1862 1270 1868 1271
rect 3574 1275 3580 1276
rect 3574 1271 3575 1275
rect 3579 1271 3580 1275
rect 3574 1270 3580 1271
rect 1822 1266 1828 1267
rect 2078 1265 2084 1266
rect 134 1261 140 1262
rect 134 1257 135 1261
rect 139 1257 140 1261
rect 134 1256 140 1257
rect 318 1261 324 1262
rect 318 1257 319 1261
rect 323 1257 324 1261
rect 318 1256 324 1257
rect 518 1261 524 1262
rect 518 1257 519 1261
rect 523 1257 524 1261
rect 518 1256 524 1257
rect 710 1261 716 1262
rect 710 1257 711 1261
rect 715 1257 716 1261
rect 710 1256 716 1257
rect 894 1261 900 1262
rect 894 1257 895 1261
rect 899 1257 900 1261
rect 894 1256 900 1257
rect 1062 1261 1068 1262
rect 1062 1257 1063 1261
rect 1067 1257 1068 1261
rect 1062 1256 1068 1257
rect 1222 1261 1228 1262
rect 1222 1257 1223 1261
rect 1227 1257 1228 1261
rect 1222 1256 1228 1257
rect 1374 1261 1380 1262
rect 1374 1257 1375 1261
rect 1379 1257 1380 1261
rect 1374 1256 1380 1257
rect 1526 1261 1532 1262
rect 1526 1257 1527 1261
rect 1531 1257 1532 1261
rect 1526 1256 1532 1257
rect 1678 1261 1684 1262
rect 1678 1257 1679 1261
rect 1683 1257 1684 1261
rect 2078 1261 2079 1265
rect 2083 1261 2084 1265
rect 2078 1260 2084 1261
rect 2302 1265 2308 1266
rect 2302 1261 2303 1265
rect 2307 1261 2308 1265
rect 2302 1260 2308 1261
rect 2510 1265 2516 1266
rect 2510 1261 2511 1265
rect 2515 1261 2516 1265
rect 2510 1260 2516 1261
rect 2702 1265 2708 1266
rect 2702 1261 2703 1265
rect 2707 1261 2708 1265
rect 2702 1260 2708 1261
rect 2878 1265 2884 1266
rect 2878 1261 2879 1265
rect 2883 1261 2884 1265
rect 2878 1260 2884 1261
rect 3038 1265 3044 1266
rect 3038 1261 3039 1265
rect 3043 1261 3044 1265
rect 3038 1260 3044 1261
rect 3190 1265 3196 1266
rect 3190 1261 3191 1265
rect 3195 1261 3196 1265
rect 3190 1260 3196 1261
rect 3342 1265 3348 1266
rect 3342 1261 3343 1265
rect 3347 1261 3348 1265
rect 3342 1260 3348 1261
rect 3478 1265 3484 1266
rect 3478 1261 3479 1265
rect 3483 1261 3484 1265
rect 3478 1260 3484 1261
rect 1678 1256 1684 1257
rect 1902 1239 1908 1240
rect 134 1235 140 1236
rect 134 1231 135 1235
rect 139 1231 140 1235
rect 134 1230 140 1231
rect 294 1235 300 1236
rect 294 1231 295 1235
rect 299 1231 300 1235
rect 294 1230 300 1231
rect 478 1235 484 1236
rect 478 1231 479 1235
rect 483 1231 484 1235
rect 478 1230 484 1231
rect 654 1235 660 1236
rect 654 1231 655 1235
rect 659 1231 660 1235
rect 654 1230 660 1231
rect 814 1235 820 1236
rect 814 1231 815 1235
rect 819 1231 820 1235
rect 814 1230 820 1231
rect 966 1235 972 1236
rect 966 1231 967 1235
rect 971 1231 972 1235
rect 966 1230 972 1231
rect 1110 1235 1116 1236
rect 1110 1231 1111 1235
rect 1115 1231 1116 1235
rect 1110 1230 1116 1231
rect 1246 1235 1252 1236
rect 1246 1231 1247 1235
rect 1251 1231 1252 1235
rect 1246 1230 1252 1231
rect 1382 1235 1388 1236
rect 1382 1231 1383 1235
rect 1387 1231 1388 1235
rect 1382 1230 1388 1231
rect 1526 1235 1532 1236
rect 1526 1231 1527 1235
rect 1531 1231 1532 1235
rect 1902 1235 1903 1239
rect 1907 1235 1908 1239
rect 1902 1234 1908 1235
rect 1990 1239 1996 1240
rect 1990 1235 1991 1239
rect 1995 1235 1996 1239
rect 1990 1234 1996 1235
rect 2094 1239 2100 1240
rect 2094 1235 2095 1239
rect 2099 1235 2100 1239
rect 2094 1234 2100 1235
rect 2214 1239 2220 1240
rect 2214 1235 2215 1239
rect 2219 1235 2220 1239
rect 2214 1234 2220 1235
rect 2350 1239 2356 1240
rect 2350 1235 2351 1239
rect 2355 1235 2356 1239
rect 2350 1234 2356 1235
rect 2486 1239 2492 1240
rect 2486 1235 2487 1239
rect 2491 1235 2492 1239
rect 2486 1234 2492 1235
rect 2630 1239 2636 1240
rect 2630 1235 2631 1239
rect 2635 1235 2636 1239
rect 2630 1234 2636 1235
rect 2774 1239 2780 1240
rect 2774 1235 2775 1239
rect 2779 1235 2780 1239
rect 2774 1234 2780 1235
rect 2918 1239 2924 1240
rect 2918 1235 2919 1239
rect 2923 1235 2924 1239
rect 2918 1234 2924 1235
rect 3062 1239 3068 1240
rect 3062 1235 3063 1239
rect 3067 1235 3068 1239
rect 3062 1234 3068 1235
rect 3206 1239 3212 1240
rect 3206 1235 3207 1239
rect 3211 1235 3212 1239
rect 3206 1234 3212 1235
rect 3350 1239 3356 1240
rect 3350 1235 3351 1239
rect 3355 1235 3356 1239
rect 3350 1234 3356 1235
rect 3478 1239 3484 1240
rect 3478 1235 3479 1239
rect 3483 1235 3484 1239
rect 3478 1234 3484 1235
rect 1526 1230 1532 1231
rect 1862 1229 1868 1230
rect 110 1225 116 1226
rect 110 1221 111 1225
rect 115 1221 116 1225
rect 110 1220 116 1221
rect 1822 1225 1828 1226
rect 1822 1221 1823 1225
rect 1827 1221 1828 1225
rect 1862 1225 1863 1229
rect 1867 1225 1868 1229
rect 1862 1224 1868 1225
rect 3574 1229 3580 1230
rect 3574 1225 3575 1229
rect 3579 1225 3580 1229
rect 3574 1224 3580 1225
rect 1822 1220 1828 1221
rect 1862 1212 1868 1213
rect 110 1208 116 1209
rect 110 1204 111 1208
rect 115 1204 116 1208
rect 110 1203 116 1204
rect 1822 1208 1828 1209
rect 1822 1204 1823 1208
rect 1827 1204 1828 1208
rect 1862 1208 1863 1212
rect 1867 1208 1868 1212
rect 1862 1207 1868 1208
rect 3574 1212 3580 1213
rect 3574 1208 3575 1212
rect 3579 1208 3580 1212
rect 3574 1207 3580 1208
rect 1822 1203 1828 1204
rect 1910 1199 1916 1200
rect 142 1195 148 1196
rect 142 1191 143 1195
rect 147 1191 148 1195
rect 142 1190 148 1191
rect 302 1195 308 1196
rect 302 1191 303 1195
rect 307 1191 308 1195
rect 302 1190 308 1191
rect 486 1195 492 1196
rect 486 1191 487 1195
rect 491 1191 492 1195
rect 486 1190 492 1191
rect 662 1195 668 1196
rect 662 1191 663 1195
rect 667 1191 668 1195
rect 662 1190 668 1191
rect 822 1195 828 1196
rect 822 1191 823 1195
rect 827 1191 828 1195
rect 822 1190 828 1191
rect 974 1195 980 1196
rect 974 1191 975 1195
rect 979 1191 980 1195
rect 974 1190 980 1191
rect 1118 1195 1124 1196
rect 1118 1191 1119 1195
rect 1123 1191 1124 1195
rect 1118 1190 1124 1191
rect 1254 1195 1260 1196
rect 1254 1191 1255 1195
rect 1259 1191 1260 1195
rect 1254 1190 1260 1191
rect 1390 1195 1396 1196
rect 1390 1191 1391 1195
rect 1395 1191 1396 1195
rect 1390 1190 1396 1191
rect 1534 1195 1540 1196
rect 1534 1191 1535 1195
rect 1539 1191 1540 1195
rect 1910 1195 1911 1199
rect 1915 1195 1916 1199
rect 1910 1194 1916 1195
rect 1998 1199 2004 1200
rect 1998 1195 1999 1199
rect 2003 1195 2004 1199
rect 1998 1194 2004 1195
rect 2102 1199 2108 1200
rect 2102 1195 2103 1199
rect 2107 1195 2108 1199
rect 2102 1194 2108 1195
rect 2222 1199 2228 1200
rect 2222 1195 2223 1199
rect 2227 1195 2228 1199
rect 2222 1194 2228 1195
rect 2358 1199 2364 1200
rect 2358 1195 2359 1199
rect 2363 1195 2364 1199
rect 2358 1194 2364 1195
rect 2494 1199 2500 1200
rect 2494 1195 2495 1199
rect 2499 1195 2500 1199
rect 2494 1194 2500 1195
rect 2638 1199 2644 1200
rect 2638 1195 2639 1199
rect 2643 1195 2644 1199
rect 2638 1194 2644 1195
rect 2782 1199 2788 1200
rect 2782 1195 2783 1199
rect 2787 1195 2788 1199
rect 2782 1194 2788 1195
rect 2926 1199 2932 1200
rect 2926 1195 2927 1199
rect 2931 1195 2932 1199
rect 2926 1194 2932 1195
rect 3070 1199 3076 1200
rect 3070 1195 3071 1199
rect 3075 1195 3076 1199
rect 3070 1194 3076 1195
rect 3214 1199 3220 1200
rect 3214 1195 3215 1199
rect 3219 1195 3220 1199
rect 3214 1194 3220 1195
rect 3358 1199 3364 1200
rect 3358 1195 3359 1199
rect 3363 1195 3364 1199
rect 3358 1194 3364 1195
rect 3486 1199 3492 1200
rect 3486 1195 3487 1199
rect 3491 1195 3492 1199
rect 3486 1194 3492 1195
rect 1534 1190 1540 1191
rect 1894 1161 1900 1162
rect 166 1157 172 1158
rect 166 1153 167 1157
rect 171 1153 172 1157
rect 166 1152 172 1153
rect 318 1157 324 1158
rect 318 1153 319 1157
rect 323 1153 324 1157
rect 318 1152 324 1153
rect 470 1157 476 1158
rect 470 1153 471 1157
rect 475 1153 476 1157
rect 470 1152 476 1153
rect 614 1157 620 1158
rect 614 1153 615 1157
rect 619 1153 620 1157
rect 614 1152 620 1153
rect 758 1157 764 1158
rect 758 1153 759 1157
rect 763 1153 764 1157
rect 758 1152 764 1153
rect 910 1157 916 1158
rect 910 1153 911 1157
rect 915 1153 916 1157
rect 910 1152 916 1153
rect 1062 1157 1068 1158
rect 1062 1153 1063 1157
rect 1067 1153 1068 1157
rect 1062 1152 1068 1153
rect 1230 1157 1236 1158
rect 1230 1153 1231 1157
rect 1235 1153 1236 1157
rect 1230 1152 1236 1153
rect 1398 1157 1404 1158
rect 1398 1153 1399 1157
rect 1403 1153 1404 1157
rect 1398 1152 1404 1153
rect 1574 1157 1580 1158
rect 1574 1153 1575 1157
rect 1579 1153 1580 1157
rect 1574 1152 1580 1153
rect 1734 1157 1740 1158
rect 1734 1153 1735 1157
rect 1739 1153 1740 1157
rect 1894 1157 1895 1161
rect 1899 1157 1900 1161
rect 1894 1156 1900 1157
rect 2062 1161 2068 1162
rect 2062 1157 2063 1161
rect 2067 1157 2068 1161
rect 2062 1156 2068 1157
rect 2254 1161 2260 1162
rect 2254 1157 2255 1161
rect 2259 1157 2260 1161
rect 2254 1156 2260 1157
rect 2438 1161 2444 1162
rect 2438 1157 2439 1161
rect 2443 1157 2444 1161
rect 2438 1156 2444 1157
rect 2614 1161 2620 1162
rect 2614 1157 2615 1161
rect 2619 1157 2620 1161
rect 2614 1156 2620 1157
rect 2790 1161 2796 1162
rect 2790 1157 2791 1161
rect 2795 1157 2796 1161
rect 2790 1156 2796 1157
rect 2966 1161 2972 1162
rect 2966 1157 2967 1161
rect 2971 1157 2972 1161
rect 2966 1156 2972 1157
rect 3142 1161 3148 1162
rect 3142 1157 3143 1161
rect 3147 1157 3148 1161
rect 3142 1156 3148 1157
rect 3326 1161 3332 1162
rect 3326 1157 3327 1161
rect 3331 1157 3332 1161
rect 3326 1156 3332 1157
rect 3486 1161 3492 1162
rect 3486 1157 3487 1161
rect 3491 1157 3492 1161
rect 3486 1156 3492 1157
rect 1734 1152 1740 1153
rect 1862 1148 1868 1149
rect 110 1144 116 1145
rect 110 1140 111 1144
rect 115 1140 116 1144
rect 110 1139 116 1140
rect 1822 1144 1828 1145
rect 1822 1140 1823 1144
rect 1827 1140 1828 1144
rect 1862 1144 1863 1148
rect 1867 1144 1868 1148
rect 1862 1143 1868 1144
rect 3574 1148 3580 1149
rect 3574 1144 3575 1148
rect 3579 1144 3580 1148
rect 3574 1143 3580 1144
rect 1822 1139 1828 1140
rect 1862 1131 1868 1132
rect 110 1127 116 1128
rect 110 1123 111 1127
rect 115 1123 116 1127
rect 110 1122 116 1123
rect 1822 1127 1828 1128
rect 1822 1123 1823 1127
rect 1827 1123 1828 1127
rect 1862 1127 1863 1131
rect 1867 1127 1868 1131
rect 1862 1126 1868 1127
rect 3574 1131 3580 1132
rect 3574 1127 3575 1131
rect 3579 1127 3580 1131
rect 3574 1126 3580 1127
rect 1822 1122 1828 1123
rect 1886 1121 1892 1122
rect 158 1117 164 1118
rect 158 1113 159 1117
rect 163 1113 164 1117
rect 158 1112 164 1113
rect 310 1117 316 1118
rect 310 1113 311 1117
rect 315 1113 316 1117
rect 310 1112 316 1113
rect 462 1117 468 1118
rect 462 1113 463 1117
rect 467 1113 468 1117
rect 462 1112 468 1113
rect 606 1117 612 1118
rect 606 1113 607 1117
rect 611 1113 612 1117
rect 606 1112 612 1113
rect 750 1117 756 1118
rect 750 1113 751 1117
rect 755 1113 756 1117
rect 750 1112 756 1113
rect 902 1117 908 1118
rect 902 1113 903 1117
rect 907 1113 908 1117
rect 902 1112 908 1113
rect 1054 1117 1060 1118
rect 1054 1113 1055 1117
rect 1059 1113 1060 1117
rect 1054 1112 1060 1113
rect 1222 1117 1228 1118
rect 1222 1113 1223 1117
rect 1227 1113 1228 1117
rect 1222 1112 1228 1113
rect 1390 1117 1396 1118
rect 1390 1113 1391 1117
rect 1395 1113 1396 1117
rect 1390 1112 1396 1113
rect 1566 1117 1572 1118
rect 1566 1113 1567 1117
rect 1571 1113 1572 1117
rect 1566 1112 1572 1113
rect 1726 1117 1732 1118
rect 1726 1113 1727 1117
rect 1731 1113 1732 1117
rect 1886 1117 1887 1121
rect 1891 1117 1892 1121
rect 1886 1116 1892 1117
rect 2054 1121 2060 1122
rect 2054 1117 2055 1121
rect 2059 1117 2060 1121
rect 2054 1116 2060 1117
rect 2246 1121 2252 1122
rect 2246 1117 2247 1121
rect 2251 1117 2252 1121
rect 2246 1116 2252 1117
rect 2430 1121 2436 1122
rect 2430 1117 2431 1121
rect 2435 1117 2436 1121
rect 2430 1116 2436 1117
rect 2606 1121 2612 1122
rect 2606 1117 2607 1121
rect 2611 1117 2612 1121
rect 2606 1116 2612 1117
rect 2782 1121 2788 1122
rect 2782 1117 2783 1121
rect 2787 1117 2788 1121
rect 2782 1116 2788 1117
rect 2958 1121 2964 1122
rect 2958 1117 2959 1121
rect 2963 1117 2964 1121
rect 2958 1116 2964 1117
rect 3134 1121 3140 1122
rect 3134 1117 3135 1121
rect 3139 1117 3140 1121
rect 3134 1116 3140 1117
rect 3318 1121 3324 1122
rect 3318 1117 3319 1121
rect 3323 1117 3324 1121
rect 3318 1116 3324 1117
rect 3478 1121 3484 1122
rect 3478 1117 3479 1121
rect 3483 1117 3484 1121
rect 3478 1116 3484 1117
rect 1726 1112 1732 1113
rect 214 1091 220 1092
rect 214 1087 215 1091
rect 219 1087 220 1091
rect 214 1086 220 1087
rect 326 1091 332 1092
rect 326 1087 327 1091
rect 331 1087 332 1091
rect 326 1086 332 1087
rect 438 1091 444 1092
rect 438 1087 439 1091
rect 443 1087 444 1091
rect 438 1086 444 1087
rect 558 1091 564 1092
rect 558 1087 559 1091
rect 563 1087 564 1091
rect 558 1086 564 1087
rect 678 1091 684 1092
rect 678 1087 679 1091
rect 683 1087 684 1091
rect 678 1086 684 1087
rect 806 1091 812 1092
rect 806 1087 807 1091
rect 811 1087 812 1091
rect 806 1086 812 1087
rect 942 1091 948 1092
rect 942 1087 943 1091
rect 947 1087 948 1091
rect 942 1086 948 1087
rect 1086 1091 1092 1092
rect 1086 1087 1087 1091
rect 1091 1087 1092 1091
rect 1086 1086 1092 1087
rect 1246 1091 1252 1092
rect 1246 1087 1247 1091
rect 1251 1087 1252 1091
rect 1246 1086 1252 1087
rect 1406 1091 1412 1092
rect 1406 1087 1407 1091
rect 1411 1087 1412 1091
rect 1406 1086 1412 1087
rect 1574 1091 1580 1092
rect 1574 1087 1575 1091
rect 1579 1087 1580 1091
rect 1574 1086 1580 1087
rect 1726 1091 1732 1092
rect 1726 1087 1727 1091
rect 1731 1087 1732 1091
rect 1726 1086 1732 1087
rect 1934 1087 1940 1088
rect 1934 1083 1935 1087
rect 1939 1083 1940 1087
rect 1934 1082 1940 1083
rect 2094 1087 2100 1088
rect 2094 1083 2095 1087
rect 2099 1083 2100 1087
rect 2094 1082 2100 1083
rect 2246 1087 2252 1088
rect 2246 1083 2247 1087
rect 2251 1083 2252 1087
rect 2246 1082 2252 1083
rect 2406 1087 2412 1088
rect 2406 1083 2407 1087
rect 2411 1083 2412 1087
rect 2406 1082 2412 1083
rect 2566 1087 2572 1088
rect 2566 1083 2567 1087
rect 2571 1083 2572 1087
rect 2566 1082 2572 1083
rect 2734 1087 2740 1088
rect 2734 1083 2735 1087
rect 2739 1083 2740 1087
rect 2734 1082 2740 1083
rect 2910 1087 2916 1088
rect 2910 1083 2911 1087
rect 2915 1083 2916 1087
rect 2910 1082 2916 1083
rect 3094 1087 3100 1088
rect 3094 1083 3095 1087
rect 3099 1083 3100 1087
rect 3094 1082 3100 1083
rect 3286 1087 3292 1088
rect 3286 1083 3287 1087
rect 3291 1083 3292 1087
rect 3286 1082 3292 1083
rect 3478 1087 3484 1088
rect 3478 1083 3479 1087
rect 3483 1083 3484 1087
rect 3478 1082 3484 1083
rect 110 1081 116 1082
rect 110 1077 111 1081
rect 115 1077 116 1081
rect 110 1076 116 1077
rect 1822 1081 1828 1082
rect 1822 1077 1823 1081
rect 1827 1077 1828 1081
rect 1822 1076 1828 1077
rect 1862 1077 1868 1078
rect 1862 1073 1863 1077
rect 1867 1073 1868 1077
rect 1862 1072 1868 1073
rect 3574 1077 3580 1078
rect 3574 1073 3575 1077
rect 3579 1073 3580 1077
rect 3574 1072 3580 1073
rect 110 1064 116 1065
rect 110 1060 111 1064
rect 115 1060 116 1064
rect 110 1059 116 1060
rect 1822 1064 1828 1065
rect 1822 1060 1823 1064
rect 1827 1060 1828 1064
rect 1822 1059 1828 1060
rect 1862 1060 1868 1061
rect 1862 1056 1863 1060
rect 1867 1056 1868 1060
rect 1862 1055 1868 1056
rect 3574 1060 3580 1061
rect 3574 1056 3575 1060
rect 3579 1056 3580 1060
rect 3574 1055 3580 1056
rect 222 1051 228 1052
rect 222 1047 223 1051
rect 227 1047 228 1051
rect 222 1046 228 1047
rect 334 1051 340 1052
rect 334 1047 335 1051
rect 339 1047 340 1051
rect 334 1046 340 1047
rect 446 1051 452 1052
rect 446 1047 447 1051
rect 451 1047 452 1051
rect 446 1046 452 1047
rect 566 1051 572 1052
rect 566 1047 567 1051
rect 571 1047 572 1051
rect 566 1046 572 1047
rect 686 1051 692 1052
rect 686 1047 687 1051
rect 691 1047 692 1051
rect 686 1046 692 1047
rect 814 1051 820 1052
rect 814 1047 815 1051
rect 819 1047 820 1051
rect 814 1046 820 1047
rect 950 1051 956 1052
rect 950 1047 951 1051
rect 955 1047 956 1051
rect 950 1046 956 1047
rect 1094 1051 1100 1052
rect 1094 1047 1095 1051
rect 1099 1047 1100 1051
rect 1094 1046 1100 1047
rect 1254 1051 1260 1052
rect 1254 1047 1255 1051
rect 1259 1047 1260 1051
rect 1254 1046 1260 1047
rect 1414 1051 1420 1052
rect 1414 1047 1415 1051
rect 1419 1047 1420 1051
rect 1414 1046 1420 1047
rect 1582 1051 1588 1052
rect 1582 1047 1583 1051
rect 1587 1047 1588 1051
rect 1582 1046 1588 1047
rect 1734 1051 1740 1052
rect 1734 1047 1735 1051
rect 1739 1047 1740 1051
rect 1734 1046 1740 1047
rect 1942 1047 1948 1048
rect 1942 1043 1943 1047
rect 1947 1043 1948 1047
rect 1942 1042 1948 1043
rect 2102 1047 2108 1048
rect 2102 1043 2103 1047
rect 2107 1043 2108 1047
rect 2102 1042 2108 1043
rect 2254 1047 2260 1048
rect 2254 1043 2255 1047
rect 2259 1043 2260 1047
rect 2254 1042 2260 1043
rect 2414 1047 2420 1048
rect 2414 1043 2415 1047
rect 2419 1043 2420 1047
rect 2414 1042 2420 1043
rect 2574 1047 2580 1048
rect 2574 1043 2575 1047
rect 2579 1043 2580 1047
rect 2574 1042 2580 1043
rect 2742 1047 2748 1048
rect 2742 1043 2743 1047
rect 2747 1043 2748 1047
rect 2742 1042 2748 1043
rect 2918 1047 2924 1048
rect 2918 1043 2919 1047
rect 2923 1043 2924 1047
rect 2918 1042 2924 1043
rect 3102 1047 3108 1048
rect 3102 1043 3103 1047
rect 3107 1043 3108 1047
rect 3102 1042 3108 1043
rect 3294 1047 3300 1048
rect 3294 1043 3295 1047
rect 3299 1043 3300 1047
rect 3294 1042 3300 1043
rect 3486 1047 3492 1048
rect 3486 1043 3487 1047
rect 3491 1043 3492 1047
rect 3486 1042 3492 1043
rect 342 1009 348 1010
rect 342 1005 343 1009
rect 347 1005 348 1009
rect 342 1004 348 1005
rect 430 1009 436 1010
rect 430 1005 431 1009
rect 435 1005 436 1009
rect 430 1004 436 1005
rect 534 1009 540 1010
rect 534 1005 535 1009
rect 539 1005 540 1009
rect 534 1004 540 1005
rect 654 1009 660 1010
rect 654 1005 655 1009
rect 659 1005 660 1009
rect 654 1004 660 1005
rect 790 1009 796 1010
rect 790 1005 791 1009
rect 795 1005 796 1009
rect 790 1004 796 1005
rect 950 1009 956 1010
rect 950 1005 951 1009
rect 955 1005 956 1009
rect 950 1004 956 1005
rect 1134 1009 1140 1010
rect 1134 1005 1135 1009
rect 1139 1005 1140 1009
rect 1134 1004 1140 1005
rect 1326 1009 1332 1010
rect 1326 1005 1327 1009
rect 1331 1005 1332 1009
rect 1326 1004 1332 1005
rect 1534 1009 1540 1010
rect 1534 1005 1535 1009
rect 1539 1005 1540 1009
rect 1534 1004 1540 1005
rect 1734 1009 1740 1010
rect 1734 1005 1735 1009
rect 1739 1005 1740 1009
rect 1734 1004 1740 1005
rect 1942 1009 1948 1010
rect 1942 1005 1943 1009
rect 1947 1005 1948 1009
rect 1942 1004 1948 1005
rect 2070 1009 2076 1010
rect 2070 1005 2071 1009
rect 2075 1005 2076 1009
rect 2070 1004 2076 1005
rect 2190 1009 2196 1010
rect 2190 1005 2191 1009
rect 2195 1005 2196 1009
rect 2190 1004 2196 1005
rect 2310 1009 2316 1010
rect 2310 1005 2311 1009
rect 2315 1005 2316 1009
rect 2310 1004 2316 1005
rect 2438 1009 2444 1010
rect 2438 1005 2439 1009
rect 2443 1005 2444 1009
rect 2438 1004 2444 1005
rect 2574 1009 2580 1010
rect 2574 1005 2575 1009
rect 2579 1005 2580 1009
rect 2574 1004 2580 1005
rect 2718 1009 2724 1010
rect 2718 1005 2719 1009
rect 2723 1005 2724 1009
rect 2718 1004 2724 1005
rect 2870 1009 2876 1010
rect 2870 1005 2871 1009
rect 2875 1005 2876 1009
rect 2870 1004 2876 1005
rect 3030 1009 3036 1010
rect 3030 1005 3031 1009
rect 3035 1005 3036 1009
rect 3030 1004 3036 1005
rect 3190 1009 3196 1010
rect 3190 1005 3191 1009
rect 3195 1005 3196 1009
rect 3190 1004 3196 1005
rect 3350 1009 3356 1010
rect 3350 1005 3351 1009
rect 3355 1005 3356 1009
rect 3350 1004 3356 1005
rect 3486 1009 3492 1010
rect 3486 1005 3487 1009
rect 3491 1005 3492 1009
rect 3486 1004 3492 1005
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 110 991 116 992
rect 1822 996 1828 997
rect 1822 992 1823 996
rect 1827 992 1828 996
rect 1822 991 1828 992
rect 1862 996 1868 997
rect 1862 992 1863 996
rect 1867 992 1868 996
rect 1862 991 1868 992
rect 3574 996 3580 997
rect 3574 992 3575 996
rect 3579 992 3580 996
rect 3574 991 3580 992
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 110 974 116 975
rect 1822 979 1828 980
rect 1822 975 1823 979
rect 1827 975 1828 979
rect 1822 974 1828 975
rect 1862 979 1868 980
rect 1862 975 1863 979
rect 1867 975 1868 979
rect 1862 974 1868 975
rect 3574 979 3580 980
rect 3574 975 3575 979
rect 3579 975 3580 979
rect 3574 974 3580 975
rect 334 969 340 970
rect 334 965 335 969
rect 339 965 340 969
rect 334 964 340 965
rect 422 969 428 970
rect 422 965 423 969
rect 427 965 428 969
rect 422 964 428 965
rect 526 969 532 970
rect 526 965 527 969
rect 531 965 532 969
rect 526 964 532 965
rect 646 969 652 970
rect 646 965 647 969
rect 651 965 652 969
rect 646 964 652 965
rect 782 969 788 970
rect 782 965 783 969
rect 787 965 788 969
rect 782 964 788 965
rect 942 969 948 970
rect 942 965 943 969
rect 947 965 948 969
rect 942 964 948 965
rect 1126 969 1132 970
rect 1126 965 1127 969
rect 1131 965 1132 969
rect 1126 964 1132 965
rect 1318 969 1324 970
rect 1318 965 1319 969
rect 1323 965 1324 969
rect 1318 964 1324 965
rect 1526 969 1532 970
rect 1526 965 1527 969
rect 1531 965 1532 969
rect 1526 964 1532 965
rect 1726 969 1732 970
rect 1726 965 1727 969
rect 1731 965 1732 969
rect 1726 964 1732 965
rect 1934 969 1940 970
rect 1934 965 1935 969
rect 1939 965 1940 969
rect 1934 964 1940 965
rect 2062 969 2068 970
rect 2062 965 2063 969
rect 2067 965 2068 969
rect 2062 964 2068 965
rect 2182 969 2188 970
rect 2182 965 2183 969
rect 2187 965 2188 969
rect 2182 964 2188 965
rect 2302 969 2308 970
rect 2302 965 2303 969
rect 2307 965 2308 969
rect 2302 964 2308 965
rect 2430 969 2436 970
rect 2430 965 2431 969
rect 2435 965 2436 969
rect 2430 964 2436 965
rect 2566 969 2572 970
rect 2566 965 2567 969
rect 2571 965 2572 969
rect 2566 964 2572 965
rect 2710 969 2716 970
rect 2710 965 2711 969
rect 2715 965 2716 969
rect 2710 964 2716 965
rect 2862 969 2868 970
rect 2862 965 2863 969
rect 2867 965 2868 969
rect 2862 964 2868 965
rect 3022 969 3028 970
rect 3022 965 3023 969
rect 3027 965 3028 969
rect 3022 964 3028 965
rect 3182 969 3188 970
rect 3182 965 3183 969
rect 3187 965 3188 969
rect 3182 964 3188 965
rect 3342 969 3348 970
rect 3342 965 3343 969
rect 3347 965 3348 969
rect 3342 964 3348 965
rect 3478 969 3484 970
rect 3478 965 3479 969
rect 3483 965 3484 969
rect 3478 964 3484 965
rect 366 943 372 944
rect 366 939 367 943
rect 371 939 372 943
rect 366 938 372 939
rect 462 943 468 944
rect 462 939 463 943
rect 467 939 468 943
rect 462 938 468 939
rect 574 943 580 944
rect 574 939 575 943
rect 579 939 580 943
rect 574 938 580 939
rect 702 943 708 944
rect 702 939 703 943
rect 707 939 708 943
rect 702 938 708 939
rect 846 943 852 944
rect 846 939 847 943
rect 851 939 852 943
rect 846 938 852 939
rect 1006 943 1012 944
rect 1006 939 1007 943
rect 1011 939 1012 943
rect 1006 938 1012 939
rect 1174 943 1180 944
rect 1174 939 1175 943
rect 1179 939 1180 943
rect 1174 938 1180 939
rect 1350 943 1356 944
rect 1350 939 1351 943
rect 1355 939 1356 943
rect 1350 938 1356 939
rect 1526 943 1532 944
rect 1526 939 1527 943
rect 1531 939 1532 943
rect 1526 938 1532 939
rect 1710 943 1716 944
rect 1710 939 1711 943
rect 1715 939 1716 943
rect 1710 938 1716 939
rect 1886 943 1892 944
rect 1886 939 1887 943
rect 1891 939 1892 943
rect 1886 938 1892 939
rect 2046 943 2052 944
rect 2046 939 2047 943
rect 2051 939 2052 943
rect 2046 938 2052 939
rect 2198 943 2204 944
rect 2198 939 2199 943
rect 2203 939 2204 943
rect 2198 938 2204 939
rect 2350 943 2356 944
rect 2350 939 2351 943
rect 2355 939 2356 943
rect 2350 938 2356 939
rect 2494 943 2500 944
rect 2494 939 2495 943
rect 2499 939 2500 943
rect 2494 938 2500 939
rect 2630 943 2636 944
rect 2630 939 2631 943
rect 2635 939 2636 943
rect 2630 938 2636 939
rect 2758 943 2764 944
rect 2758 939 2759 943
rect 2763 939 2764 943
rect 2758 938 2764 939
rect 2886 943 2892 944
rect 2886 939 2887 943
rect 2891 939 2892 943
rect 2886 938 2892 939
rect 3022 943 3028 944
rect 3022 939 3023 943
rect 3027 939 3028 943
rect 3022 938 3028 939
rect 110 933 116 934
rect 110 929 111 933
rect 115 929 116 933
rect 110 928 116 929
rect 1822 933 1828 934
rect 1822 929 1823 933
rect 1827 929 1828 933
rect 1822 928 1828 929
rect 1862 933 1868 934
rect 1862 929 1863 933
rect 1867 929 1868 933
rect 1862 928 1868 929
rect 3574 933 3580 934
rect 3574 929 3575 933
rect 3579 929 3580 933
rect 3574 928 3580 929
rect 110 916 116 917
rect 110 912 111 916
rect 115 912 116 916
rect 110 911 116 912
rect 1822 916 1828 917
rect 1822 912 1823 916
rect 1827 912 1828 916
rect 1822 911 1828 912
rect 1862 916 1868 917
rect 1862 912 1863 916
rect 1867 912 1868 916
rect 1862 911 1868 912
rect 3574 916 3580 917
rect 3574 912 3575 916
rect 3579 912 3580 916
rect 3574 911 3580 912
rect 374 903 380 904
rect 374 899 375 903
rect 379 899 380 903
rect 374 898 380 899
rect 470 903 476 904
rect 470 899 471 903
rect 475 899 476 903
rect 470 898 476 899
rect 582 903 588 904
rect 582 899 583 903
rect 587 899 588 903
rect 582 898 588 899
rect 710 903 716 904
rect 710 899 711 903
rect 715 899 716 903
rect 710 898 716 899
rect 854 903 860 904
rect 854 899 855 903
rect 859 899 860 903
rect 854 898 860 899
rect 1014 903 1020 904
rect 1014 899 1015 903
rect 1019 899 1020 903
rect 1014 898 1020 899
rect 1182 903 1188 904
rect 1182 899 1183 903
rect 1187 899 1188 903
rect 1182 898 1188 899
rect 1358 903 1364 904
rect 1358 899 1359 903
rect 1363 899 1364 903
rect 1358 898 1364 899
rect 1534 903 1540 904
rect 1534 899 1535 903
rect 1539 899 1540 903
rect 1534 898 1540 899
rect 1718 903 1724 904
rect 1718 899 1719 903
rect 1723 899 1724 903
rect 1718 898 1724 899
rect 1894 903 1900 904
rect 1894 899 1895 903
rect 1899 899 1900 903
rect 1894 898 1900 899
rect 2054 903 2060 904
rect 2054 899 2055 903
rect 2059 899 2060 903
rect 2054 898 2060 899
rect 2206 903 2212 904
rect 2206 899 2207 903
rect 2211 899 2212 903
rect 2206 898 2212 899
rect 2358 903 2364 904
rect 2358 899 2359 903
rect 2363 899 2364 903
rect 2358 898 2364 899
rect 2502 903 2508 904
rect 2502 899 2503 903
rect 2507 899 2508 903
rect 2502 898 2508 899
rect 2638 903 2644 904
rect 2638 899 2639 903
rect 2643 899 2644 903
rect 2638 898 2644 899
rect 2766 903 2772 904
rect 2766 899 2767 903
rect 2771 899 2772 903
rect 2766 898 2772 899
rect 2894 903 2900 904
rect 2894 899 2895 903
rect 2899 899 2900 903
rect 2894 898 2900 899
rect 3030 903 3036 904
rect 3030 899 3031 903
rect 3035 899 3036 903
rect 3030 898 3036 899
rect 1894 869 1900 870
rect 342 865 348 866
rect 342 861 343 865
rect 347 861 348 865
rect 342 860 348 861
rect 430 865 436 866
rect 430 861 431 865
rect 435 861 436 865
rect 430 860 436 861
rect 534 865 540 866
rect 534 861 535 865
rect 539 861 540 865
rect 534 860 540 861
rect 646 865 652 866
rect 646 861 647 865
rect 651 861 652 865
rect 646 860 652 861
rect 782 865 788 866
rect 782 861 783 865
rect 787 861 788 865
rect 782 860 788 861
rect 926 865 932 866
rect 926 861 927 865
rect 931 861 932 865
rect 926 860 932 861
rect 1086 865 1092 866
rect 1086 861 1087 865
rect 1091 861 1092 865
rect 1086 860 1092 861
rect 1262 865 1268 866
rect 1262 861 1263 865
rect 1267 861 1268 865
rect 1262 860 1268 861
rect 1446 865 1452 866
rect 1446 861 1447 865
rect 1451 861 1452 865
rect 1446 860 1452 861
rect 1630 865 1636 866
rect 1630 861 1631 865
rect 1635 861 1636 865
rect 1894 865 1895 869
rect 1899 865 1900 869
rect 1894 864 1900 865
rect 2014 869 2020 870
rect 2014 865 2015 869
rect 2019 865 2020 869
rect 2014 864 2020 865
rect 2166 869 2172 870
rect 2166 865 2167 869
rect 2171 865 2172 869
rect 2166 864 2172 865
rect 2318 869 2324 870
rect 2318 865 2319 869
rect 2323 865 2324 869
rect 2318 864 2324 865
rect 2486 869 2492 870
rect 2486 865 2487 869
rect 2491 865 2492 869
rect 2486 864 2492 865
rect 2662 869 2668 870
rect 2662 865 2663 869
rect 2667 865 2668 869
rect 2662 864 2668 865
rect 2846 869 2852 870
rect 2846 865 2847 869
rect 2851 865 2852 869
rect 2846 864 2852 865
rect 3038 869 3044 870
rect 3038 865 3039 869
rect 3043 865 3044 869
rect 3038 864 3044 865
rect 3238 869 3244 870
rect 3238 865 3239 869
rect 3243 865 3244 869
rect 3238 864 3244 865
rect 3438 869 3444 870
rect 3438 865 3439 869
rect 3443 865 3444 869
rect 3438 864 3444 865
rect 1630 860 1636 861
rect 1862 856 1868 857
rect 110 852 116 853
rect 110 848 111 852
rect 115 848 116 852
rect 110 847 116 848
rect 1822 852 1828 853
rect 1822 848 1823 852
rect 1827 848 1828 852
rect 1862 852 1863 856
rect 1867 852 1868 856
rect 1862 851 1868 852
rect 3574 856 3580 857
rect 3574 852 3575 856
rect 3579 852 3580 856
rect 3574 851 3580 852
rect 1822 847 1828 848
rect 1862 839 1868 840
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 110 830 116 831
rect 1822 835 1828 836
rect 1822 831 1823 835
rect 1827 831 1828 835
rect 1862 835 1863 839
rect 1867 835 1868 839
rect 1862 834 1868 835
rect 3574 839 3580 840
rect 3574 835 3575 839
rect 3579 835 3580 839
rect 3574 834 3580 835
rect 1822 830 1828 831
rect 1886 829 1892 830
rect 334 825 340 826
rect 334 821 335 825
rect 339 821 340 825
rect 334 820 340 821
rect 422 825 428 826
rect 422 821 423 825
rect 427 821 428 825
rect 422 820 428 821
rect 526 825 532 826
rect 526 821 527 825
rect 531 821 532 825
rect 526 820 532 821
rect 638 825 644 826
rect 638 821 639 825
rect 643 821 644 825
rect 638 820 644 821
rect 774 825 780 826
rect 774 821 775 825
rect 779 821 780 825
rect 774 820 780 821
rect 918 825 924 826
rect 918 821 919 825
rect 923 821 924 825
rect 918 820 924 821
rect 1078 825 1084 826
rect 1078 821 1079 825
rect 1083 821 1084 825
rect 1078 820 1084 821
rect 1254 825 1260 826
rect 1254 821 1255 825
rect 1259 821 1260 825
rect 1254 820 1260 821
rect 1438 825 1444 826
rect 1438 821 1439 825
rect 1443 821 1444 825
rect 1438 820 1444 821
rect 1622 825 1628 826
rect 1622 821 1623 825
rect 1627 821 1628 825
rect 1886 825 1887 829
rect 1891 825 1892 829
rect 1886 824 1892 825
rect 2006 829 2012 830
rect 2006 825 2007 829
rect 2011 825 2012 829
rect 2006 824 2012 825
rect 2158 829 2164 830
rect 2158 825 2159 829
rect 2163 825 2164 829
rect 2158 824 2164 825
rect 2310 829 2316 830
rect 2310 825 2311 829
rect 2315 825 2316 829
rect 2310 824 2316 825
rect 2478 829 2484 830
rect 2478 825 2479 829
rect 2483 825 2484 829
rect 2478 824 2484 825
rect 2654 829 2660 830
rect 2654 825 2655 829
rect 2659 825 2660 829
rect 2654 824 2660 825
rect 2838 829 2844 830
rect 2838 825 2839 829
rect 2843 825 2844 829
rect 2838 824 2844 825
rect 3030 829 3036 830
rect 3030 825 3031 829
rect 3035 825 3036 829
rect 3030 824 3036 825
rect 3230 829 3236 830
rect 3230 825 3231 829
rect 3235 825 3236 829
rect 3230 824 3236 825
rect 3430 829 3436 830
rect 3430 825 3431 829
rect 3435 825 3436 829
rect 3430 824 3436 825
rect 1622 820 1628 821
rect 1886 807 1892 808
rect 286 803 292 804
rect 286 799 287 803
rect 291 799 292 803
rect 286 798 292 799
rect 406 803 412 804
rect 406 799 407 803
rect 411 799 412 803
rect 406 798 412 799
rect 534 803 540 804
rect 534 799 535 803
rect 539 799 540 803
rect 534 798 540 799
rect 678 803 684 804
rect 678 799 679 803
rect 683 799 684 803
rect 678 798 684 799
rect 822 803 828 804
rect 822 799 823 803
rect 827 799 828 803
rect 822 798 828 799
rect 974 803 980 804
rect 974 799 975 803
rect 979 799 980 803
rect 974 798 980 799
rect 1126 803 1132 804
rect 1126 799 1127 803
rect 1131 799 1132 803
rect 1126 798 1132 799
rect 1278 803 1284 804
rect 1278 799 1279 803
rect 1283 799 1284 803
rect 1278 798 1284 799
rect 1438 803 1444 804
rect 1438 799 1439 803
rect 1443 799 1444 803
rect 1438 798 1444 799
rect 1598 803 1604 804
rect 1598 799 1599 803
rect 1603 799 1604 803
rect 1886 803 1887 807
rect 1891 803 1892 807
rect 1886 802 1892 803
rect 1990 807 1996 808
rect 1990 803 1991 807
rect 1995 803 1996 807
rect 1990 802 1996 803
rect 2134 807 2140 808
rect 2134 803 2135 807
rect 2139 803 2140 807
rect 2134 802 2140 803
rect 2286 807 2292 808
rect 2286 803 2287 807
rect 2291 803 2292 807
rect 2286 802 2292 803
rect 2454 807 2460 808
rect 2454 803 2455 807
rect 2459 803 2460 807
rect 2454 802 2460 803
rect 2622 807 2628 808
rect 2622 803 2623 807
rect 2627 803 2628 807
rect 2622 802 2628 803
rect 2798 807 2804 808
rect 2798 803 2799 807
rect 2803 803 2804 807
rect 2798 802 2804 803
rect 2966 807 2972 808
rect 2966 803 2967 807
rect 2971 803 2972 807
rect 2966 802 2972 803
rect 3142 807 3148 808
rect 3142 803 3143 807
rect 3147 803 3148 807
rect 3142 802 3148 803
rect 3318 807 3324 808
rect 3318 803 3319 807
rect 3323 803 3324 807
rect 3318 802 3324 803
rect 3478 807 3484 808
rect 3478 803 3479 807
rect 3483 803 3484 807
rect 3478 802 3484 803
rect 1598 798 1604 799
rect 1862 797 1868 798
rect 110 793 116 794
rect 110 789 111 793
rect 115 789 116 793
rect 110 788 116 789
rect 1822 793 1828 794
rect 1822 789 1823 793
rect 1827 789 1828 793
rect 1862 793 1863 797
rect 1867 793 1868 797
rect 1862 792 1868 793
rect 3574 797 3580 798
rect 3574 793 3575 797
rect 3579 793 3580 797
rect 3574 792 3580 793
rect 1822 788 1828 789
rect 1862 780 1868 781
rect 110 776 116 777
rect 110 772 111 776
rect 115 772 116 776
rect 110 771 116 772
rect 1822 776 1828 777
rect 1822 772 1823 776
rect 1827 772 1828 776
rect 1862 776 1863 780
rect 1867 776 1868 780
rect 1862 775 1868 776
rect 3574 780 3580 781
rect 3574 776 3575 780
rect 3579 776 3580 780
rect 3574 775 3580 776
rect 1822 771 1828 772
rect 1894 767 1900 768
rect 294 763 300 764
rect 294 759 295 763
rect 299 759 300 763
rect 294 758 300 759
rect 414 763 420 764
rect 414 759 415 763
rect 419 759 420 763
rect 414 758 420 759
rect 542 763 548 764
rect 542 759 543 763
rect 547 759 548 763
rect 542 758 548 759
rect 686 763 692 764
rect 686 759 687 763
rect 691 759 692 763
rect 686 758 692 759
rect 830 763 836 764
rect 830 759 831 763
rect 835 759 836 763
rect 830 758 836 759
rect 982 763 988 764
rect 982 759 983 763
rect 987 759 988 763
rect 982 758 988 759
rect 1134 763 1140 764
rect 1134 759 1135 763
rect 1139 759 1140 763
rect 1134 758 1140 759
rect 1286 763 1292 764
rect 1286 759 1287 763
rect 1291 759 1292 763
rect 1286 758 1292 759
rect 1446 763 1452 764
rect 1446 759 1447 763
rect 1451 759 1452 763
rect 1446 758 1452 759
rect 1606 763 1612 764
rect 1606 759 1607 763
rect 1611 759 1612 763
rect 1894 763 1895 767
rect 1899 763 1900 767
rect 1894 762 1900 763
rect 1998 767 2004 768
rect 1998 763 1999 767
rect 2003 763 2004 767
rect 1998 762 2004 763
rect 2142 767 2148 768
rect 2142 763 2143 767
rect 2147 763 2148 767
rect 2142 762 2148 763
rect 2294 767 2300 768
rect 2294 763 2295 767
rect 2299 763 2300 767
rect 2294 762 2300 763
rect 2462 767 2468 768
rect 2462 763 2463 767
rect 2467 763 2468 767
rect 2462 762 2468 763
rect 2630 767 2636 768
rect 2630 763 2631 767
rect 2635 763 2636 767
rect 2630 762 2636 763
rect 2806 767 2812 768
rect 2806 763 2807 767
rect 2811 763 2812 767
rect 2806 762 2812 763
rect 2974 767 2980 768
rect 2974 763 2975 767
rect 2979 763 2980 767
rect 2974 762 2980 763
rect 3150 767 3156 768
rect 3150 763 3151 767
rect 3155 763 3156 767
rect 3150 762 3156 763
rect 3326 767 3332 768
rect 3326 763 3327 767
rect 3331 763 3332 767
rect 3326 762 3332 763
rect 3486 767 3492 768
rect 3486 763 3487 767
rect 3491 763 3492 767
rect 3486 762 3492 763
rect 1606 758 1612 759
rect 1894 729 1900 730
rect 214 725 220 726
rect 214 721 215 725
rect 219 721 220 725
rect 214 720 220 721
rect 358 725 364 726
rect 358 721 359 725
rect 363 721 364 725
rect 358 720 364 721
rect 502 725 508 726
rect 502 721 503 725
rect 507 721 508 725
rect 502 720 508 721
rect 646 725 652 726
rect 646 721 647 725
rect 651 721 652 725
rect 646 720 652 721
rect 790 725 796 726
rect 790 721 791 725
rect 795 721 796 725
rect 790 720 796 721
rect 934 725 940 726
rect 934 721 935 725
rect 939 721 940 725
rect 934 720 940 721
rect 1086 725 1092 726
rect 1086 721 1087 725
rect 1091 721 1092 725
rect 1086 720 1092 721
rect 1246 725 1252 726
rect 1246 721 1247 725
rect 1251 721 1252 725
rect 1246 720 1252 721
rect 1414 725 1420 726
rect 1414 721 1415 725
rect 1419 721 1420 725
rect 1414 720 1420 721
rect 1582 725 1588 726
rect 1582 721 1583 725
rect 1587 721 1588 725
rect 1582 720 1588 721
rect 1734 725 1740 726
rect 1734 721 1735 725
rect 1739 721 1740 725
rect 1894 725 1895 729
rect 1899 725 1900 729
rect 1894 724 1900 725
rect 2062 729 2068 730
rect 2062 725 2063 729
rect 2067 725 2068 729
rect 2062 724 2068 725
rect 2254 729 2260 730
rect 2254 725 2255 729
rect 2259 725 2260 729
rect 2254 724 2260 725
rect 2446 729 2452 730
rect 2446 725 2447 729
rect 2451 725 2452 729
rect 2446 724 2452 725
rect 2638 729 2644 730
rect 2638 725 2639 729
rect 2643 725 2644 729
rect 2638 724 2644 725
rect 2822 729 2828 730
rect 2822 725 2823 729
rect 2827 725 2828 729
rect 2822 724 2828 725
rect 2998 729 3004 730
rect 2998 725 2999 729
rect 3003 725 3004 729
rect 2998 724 3004 725
rect 3166 729 3172 730
rect 3166 725 3167 729
rect 3171 725 3172 729
rect 3166 724 3172 725
rect 3334 729 3340 730
rect 3334 725 3335 729
rect 3339 725 3340 729
rect 3334 724 3340 725
rect 3486 729 3492 730
rect 3486 725 3487 729
rect 3491 725 3492 729
rect 3486 724 3492 725
rect 1734 720 1740 721
rect 1862 716 1868 717
rect 110 712 116 713
rect 110 708 111 712
rect 115 708 116 712
rect 110 707 116 708
rect 1822 712 1828 713
rect 1822 708 1823 712
rect 1827 708 1828 712
rect 1862 712 1863 716
rect 1867 712 1868 716
rect 1862 711 1868 712
rect 3574 716 3580 717
rect 3574 712 3575 716
rect 3579 712 3580 716
rect 3574 711 3580 712
rect 1822 707 1828 708
rect 1862 699 1868 700
rect 110 695 116 696
rect 110 691 111 695
rect 115 691 116 695
rect 110 690 116 691
rect 1822 695 1828 696
rect 1822 691 1823 695
rect 1827 691 1828 695
rect 1862 695 1863 699
rect 1867 695 1868 699
rect 1862 694 1868 695
rect 3574 699 3580 700
rect 3574 695 3575 699
rect 3579 695 3580 699
rect 3574 694 3580 695
rect 1822 690 1828 691
rect 1886 689 1892 690
rect 206 685 212 686
rect 206 681 207 685
rect 211 681 212 685
rect 206 680 212 681
rect 350 685 356 686
rect 350 681 351 685
rect 355 681 356 685
rect 350 680 356 681
rect 494 685 500 686
rect 494 681 495 685
rect 499 681 500 685
rect 494 680 500 681
rect 638 685 644 686
rect 638 681 639 685
rect 643 681 644 685
rect 638 680 644 681
rect 782 685 788 686
rect 782 681 783 685
rect 787 681 788 685
rect 782 680 788 681
rect 926 685 932 686
rect 926 681 927 685
rect 931 681 932 685
rect 926 680 932 681
rect 1078 685 1084 686
rect 1078 681 1079 685
rect 1083 681 1084 685
rect 1078 680 1084 681
rect 1238 685 1244 686
rect 1238 681 1239 685
rect 1243 681 1244 685
rect 1238 680 1244 681
rect 1406 685 1412 686
rect 1406 681 1407 685
rect 1411 681 1412 685
rect 1406 680 1412 681
rect 1574 685 1580 686
rect 1574 681 1575 685
rect 1579 681 1580 685
rect 1574 680 1580 681
rect 1726 685 1732 686
rect 1726 681 1727 685
rect 1731 681 1732 685
rect 1886 685 1887 689
rect 1891 685 1892 689
rect 1886 684 1892 685
rect 2054 689 2060 690
rect 2054 685 2055 689
rect 2059 685 2060 689
rect 2054 684 2060 685
rect 2246 689 2252 690
rect 2246 685 2247 689
rect 2251 685 2252 689
rect 2246 684 2252 685
rect 2438 689 2444 690
rect 2438 685 2439 689
rect 2443 685 2444 689
rect 2438 684 2444 685
rect 2630 689 2636 690
rect 2630 685 2631 689
rect 2635 685 2636 689
rect 2630 684 2636 685
rect 2814 689 2820 690
rect 2814 685 2815 689
rect 2819 685 2820 689
rect 2814 684 2820 685
rect 2990 689 2996 690
rect 2990 685 2991 689
rect 2995 685 2996 689
rect 2990 684 2996 685
rect 3158 689 3164 690
rect 3158 685 3159 689
rect 3163 685 3164 689
rect 3158 684 3164 685
rect 3326 689 3332 690
rect 3326 685 3327 689
rect 3331 685 3332 689
rect 3326 684 3332 685
rect 3478 689 3484 690
rect 3478 685 3479 689
rect 3483 685 3484 689
rect 3478 684 3484 685
rect 1726 680 1732 681
rect 134 663 140 664
rect 134 659 135 663
rect 139 659 140 663
rect 134 658 140 659
rect 294 663 300 664
rect 294 659 295 663
rect 299 659 300 663
rect 294 658 300 659
rect 462 663 468 664
rect 462 659 463 663
rect 467 659 468 663
rect 462 658 468 659
rect 622 663 628 664
rect 622 659 623 663
rect 627 659 628 663
rect 622 658 628 659
rect 774 663 780 664
rect 774 659 775 663
rect 779 659 780 663
rect 774 658 780 659
rect 926 663 932 664
rect 926 659 927 663
rect 931 659 932 663
rect 926 658 932 659
rect 1070 663 1076 664
rect 1070 659 1071 663
rect 1075 659 1076 663
rect 1070 658 1076 659
rect 1206 663 1212 664
rect 1206 659 1207 663
rect 1211 659 1212 663
rect 1206 658 1212 659
rect 1342 663 1348 664
rect 1342 659 1343 663
rect 1347 659 1348 663
rect 1342 658 1348 659
rect 1478 663 1484 664
rect 1478 659 1479 663
rect 1483 659 1484 663
rect 1478 658 1484 659
rect 1614 663 1620 664
rect 1614 659 1615 663
rect 1619 659 1620 663
rect 1614 658 1620 659
rect 1726 663 1732 664
rect 1726 659 1727 663
rect 1731 659 1732 663
rect 1726 658 1732 659
rect 2214 663 2220 664
rect 2214 659 2215 663
rect 2219 659 2220 663
rect 2214 658 2220 659
rect 2358 663 2364 664
rect 2358 659 2359 663
rect 2363 659 2364 663
rect 2358 658 2364 659
rect 2510 663 2516 664
rect 2510 659 2511 663
rect 2515 659 2516 663
rect 2510 658 2516 659
rect 2670 663 2676 664
rect 2670 659 2671 663
rect 2675 659 2676 663
rect 2670 658 2676 659
rect 2830 663 2836 664
rect 2830 659 2831 663
rect 2835 659 2836 663
rect 2830 658 2836 659
rect 2990 663 2996 664
rect 2990 659 2991 663
rect 2995 659 2996 663
rect 2990 658 2996 659
rect 3158 663 3164 664
rect 3158 659 3159 663
rect 3163 659 3164 663
rect 3158 658 3164 659
rect 3326 663 3332 664
rect 3326 659 3327 663
rect 3331 659 3332 663
rect 3326 658 3332 659
rect 3478 663 3484 664
rect 3478 659 3479 663
rect 3483 659 3484 663
rect 3478 658 3484 659
rect 110 653 116 654
rect 110 649 111 653
rect 115 649 116 653
rect 110 648 116 649
rect 1822 653 1828 654
rect 1822 649 1823 653
rect 1827 649 1828 653
rect 1822 648 1828 649
rect 1862 653 1868 654
rect 1862 649 1863 653
rect 1867 649 1868 653
rect 1862 648 1868 649
rect 3574 653 3580 654
rect 3574 649 3575 653
rect 3579 649 3580 653
rect 3574 648 3580 649
rect 110 636 116 637
rect 110 632 111 636
rect 115 632 116 636
rect 110 631 116 632
rect 1822 636 1828 637
rect 1822 632 1823 636
rect 1827 632 1828 636
rect 1822 631 1828 632
rect 1862 636 1868 637
rect 1862 632 1863 636
rect 1867 632 1868 636
rect 1862 631 1868 632
rect 3574 636 3580 637
rect 3574 632 3575 636
rect 3579 632 3580 636
rect 3574 631 3580 632
rect 142 623 148 624
rect 142 619 143 623
rect 147 619 148 623
rect 142 618 148 619
rect 302 623 308 624
rect 302 619 303 623
rect 307 619 308 623
rect 302 618 308 619
rect 470 623 476 624
rect 470 619 471 623
rect 475 619 476 623
rect 470 618 476 619
rect 630 623 636 624
rect 630 619 631 623
rect 635 619 636 623
rect 630 618 636 619
rect 782 623 788 624
rect 782 619 783 623
rect 787 619 788 623
rect 782 618 788 619
rect 934 623 940 624
rect 934 619 935 623
rect 939 619 940 623
rect 934 618 940 619
rect 1078 623 1084 624
rect 1078 619 1079 623
rect 1083 619 1084 623
rect 1078 618 1084 619
rect 1214 623 1220 624
rect 1214 619 1215 623
rect 1219 619 1220 623
rect 1214 618 1220 619
rect 1350 623 1356 624
rect 1350 619 1351 623
rect 1355 619 1356 623
rect 1350 618 1356 619
rect 1486 623 1492 624
rect 1486 619 1487 623
rect 1491 619 1492 623
rect 1486 618 1492 619
rect 1622 623 1628 624
rect 1622 619 1623 623
rect 1627 619 1628 623
rect 1622 618 1628 619
rect 1734 623 1740 624
rect 1734 619 1735 623
rect 1739 619 1740 623
rect 1734 618 1740 619
rect 2222 623 2228 624
rect 2222 619 2223 623
rect 2227 619 2228 623
rect 2222 618 2228 619
rect 2366 623 2372 624
rect 2366 619 2367 623
rect 2371 619 2372 623
rect 2366 618 2372 619
rect 2518 623 2524 624
rect 2518 619 2519 623
rect 2523 619 2524 623
rect 2518 618 2524 619
rect 2678 623 2684 624
rect 2678 619 2679 623
rect 2683 619 2684 623
rect 2678 618 2684 619
rect 2838 623 2844 624
rect 2838 619 2839 623
rect 2843 619 2844 623
rect 2838 618 2844 619
rect 2998 623 3004 624
rect 2998 619 2999 623
rect 3003 619 3004 623
rect 2998 618 3004 619
rect 3166 623 3172 624
rect 3166 619 3167 623
rect 3171 619 3172 623
rect 3166 618 3172 619
rect 3334 623 3340 624
rect 3334 619 3335 623
rect 3339 619 3340 623
rect 3334 618 3340 619
rect 3486 623 3492 624
rect 3486 619 3487 623
rect 3491 619 3492 623
rect 3486 618 3492 619
rect 142 585 148 586
rect 142 581 143 585
rect 147 581 148 585
rect 142 580 148 581
rect 302 585 308 586
rect 302 581 303 585
rect 307 581 308 585
rect 302 580 308 581
rect 486 585 492 586
rect 486 581 487 585
rect 491 581 492 585
rect 486 580 492 581
rect 670 585 676 586
rect 670 581 671 585
rect 675 581 676 585
rect 670 580 676 581
rect 846 585 852 586
rect 846 581 847 585
rect 851 581 852 585
rect 846 580 852 581
rect 1022 585 1028 586
rect 1022 581 1023 585
rect 1027 581 1028 585
rect 1022 580 1028 581
rect 1198 585 1204 586
rect 1198 581 1199 585
rect 1203 581 1204 585
rect 1198 580 1204 581
rect 1374 585 1380 586
rect 1374 581 1375 585
rect 1379 581 1380 585
rect 1374 580 1380 581
rect 1558 585 1564 586
rect 1558 581 1559 585
rect 1563 581 1564 585
rect 1558 580 1564 581
rect 1734 585 1740 586
rect 1734 581 1735 585
rect 1739 581 1740 585
rect 1734 580 1740 581
rect 2198 585 2204 586
rect 2198 581 2199 585
rect 2203 581 2204 585
rect 2198 580 2204 581
rect 2286 585 2292 586
rect 2286 581 2287 585
rect 2291 581 2292 585
rect 2286 580 2292 581
rect 2374 585 2380 586
rect 2374 581 2375 585
rect 2379 581 2380 585
rect 2374 580 2380 581
rect 2462 585 2468 586
rect 2462 581 2463 585
rect 2467 581 2468 585
rect 2462 580 2468 581
rect 2566 585 2572 586
rect 2566 581 2567 585
rect 2571 581 2572 585
rect 2566 580 2572 581
rect 2678 585 2684 586
rect 2678 581 2679 585
rect 2683 581 2684 585
rect 2678 580 2684 581
rect 2814 585 2820 586
rect 2814 581 2815 585
rect 2819 581 2820 585
rect 2814 580 2820 581
rect 2974 585 2980 586
rect 2974 581 2975 585
rect 2979 581 2980 585
rect 2974 580 2980 581
rect 3142 585 3148 586
rect 3142 581 3143 585
rect 3147 581 3148 585
rect 3142 580 3148 581
rect 3326 585 3332 586
rect 3326 581 3327 585
rect 3331 581 3332 585
rect 3326 580 3332 581
rect 3486 585 3492 586
rect 3486 581 3487 585
rect 3491 581 3492 585
rect 3486 580 3492 581
rect 110 572 116 573
rect 110 568 111 572
rect 115 568 116 572
rect 110 567 116 568
rect 1822 572 1828 573
rect 1822 568 1823 572
rect 1827 568 1828 572
rect 1822 567 1828 568
rect 1862 572 1868 573
rect 1862 568 1863 572
rect 1867 568 1868 572
rect 1862 567 1868 568
rect 3574 572 3580 573
rect 3574 568 3575 572
rect 3579 568 3580 572
rect 3574 567 3580 568
rect 110 555 116 556
rect 110 551 111 555
rect 115 551 116 555
rect 110 550 116 551
rect 1822 555 1828 556
rect 1822 551 1823 555
rect 1827 551 1828 555
rect 1822 550 1828 551
rect 1862 555 1868 556
rect 1862 551 1863 555
rect 1867 551 1868 555
rect 1862 550 1868 551
rect 3574 555 3580 556
rect 3574 551 3575 555
rect 3579 551 3580 555
rect 3574 550 3580 551
rect 134 545 140 546
rect 134 541 135 545
rect 139 541 140 545
rect 134 540 140 541
rect 294 545 300 546
rect 294 541 295 545
rect 299 541 300 545
rect 294 540 300 541
rect 478 545 484 546
rect 478 541 479 545
rect 483 541 484 545
rect 478 540 484 541
rect 662 545 668 546
rect 662 541 663 545
rect 667 541 668 545
rect 662 540 668 541
rect 838 545 844 546
rect 838 541 839 545
rect 843 541 844 545
rect 838 540 844 541
rect 1014 545 1020 546
rect 1014 541 1015 545
rect 1019 541 1020 545
rect 1014 540 1020 541
rect 1190 545 1196 546
rect 1190 541 1191 545
rect 1195 541 1196 545
rect 1190 540 1196 541
rect 1366 545 1372 546
rect 1366 541 1367 545
rect 1371 541 1372 545
rect 1366 540 1372 541
rect 1550 545 1556 546
rect 1550 541 1551 545
rect 1555 541 1556 545
rect 1550 540 1556 541
rect 1726 545 1732 546
rect 1726 541 1727 545
rect 1731 541 1732 545
rect 1726 540 1732 541
rect 2190 545 2196 546
rect 2190 541 2191 545
rect 2195 541 2196 545
rect 2190 540 2196 541
rect 2278 545 2284 546
rect 2278 541 2279 545
rect 2283 541 2284 545
rect 2278 540 2284 541
rect 2366 545 2372 546
rect 2366 541 2367 545
rect 2371 541 2372 545
rect 2366 540 2372 541
rect 2454 545 2460 546
rect 2454 541 2455 545
rect 2459 541 2460 545
rect 2454 540 2460 541
rect 2558 545 2564 546
rect 2558 541 2559 545
rect 2563 541 2564 545
rect 2558 540 2564 541
rect 2670 545 2676 546
rect 2670 541 2671 545
rect 2675 541 2676 545
rect 2670 540 2676 541
rect 2806 545 2812 546
rect 2806 541 2807 545
rect 2811 541 2812 545
rect 2806 540 2812 541
rect 2966 545 2972 546
rect 2966 541 2967 545
rect 2971 541 2972 545
rect 2966 540 2972 541
rect 3134 545 3140 546
rect 3134 541 3135 545
rect 3139 541 3140 545
rect 3134 540 3140 541
rect 3318 545 3324 546
rect 3318 541 3319 545
rect 3323 541 3324 545
rect 3318 540 3324 541
rect 3478 545 3484 546
rect 3478 541 3479 545
rect 3483 541 3484 545
rect 3478 540 3484 541
rect 134 519 140 520
rect 134 515 135 519
rect 139 515 140 519
rect 134 514 140 515
rect 302 519 308 520
rect 302 515 303 519
rect 307 515 308 519
rect 302 514 308 515
rect 494 519 500 520
rect 494 515 495 519
rect 499 515 500 519
rect 494 514 500 515
rect 678 519 684 520
rect 678 515 679 519
rect 683 515 684 519
rect 678 514 684 515
rect 862 519 868 520
rect 862 515 863 519
rect 867 515 868 519
rect 862 514 868 515
rect 1030 519 1036 520
rect 1030 515 1031 519
rect 1035 515 1036 519
rect 1030 514 1036 515
rect 1190 519 1196 520
rect 1190 515 1191 519
rect 1195 515 1196 519
rect 1190 514 1196 515
rect 1350 519 1356 520
rect 1350 515 1351 519
rect 1355 515 1356 519
rect 1350 514 1356 515
rect 1502 519 1508 520
rect 1502 515 1503 519
rect 1507 515 1508 519
rect 1502 514 1508 515
rect 1662 519 1668 520
rect 1662 515 1663 519
rect 1667 515 1668 519
rect 1662 514 1668 515
rect 2302 519 2308 520
rect 2302 515 2303 519
rect 2307 515 2308 519
rect 2302 514 2308 515
rect 2398 519 2404 520
rect 2398 515 2399 519
rect 2403 515 2404 519
rect 2398 514 2404 515
rect 2502 519 2508 520
rect 2502 515 2503 519
rect 2507 515 2508 519
rect 2502 514 2508 515
rect 2606 519 2612 520
rect 2606 515 2607 519
rect 2611 515 2612 519
rect 2606 514 2612 515
rect 2718 519 2724 520
rect 2718 515 2719 519
rect 2723 515 2724 519
rect 2718 514 2724 515
rect 2838 519 2844 520
rect 2838 515 2839 519
rect 2843 515 2844 519
rect 2838 514 2844 515
rect 2966 519 2972 520
rect 2966 515 2967 519
rect 2971 515 2972 519
rect 2966 514 2972 515
rect 3094 519 3100 520
rect 3094 515 3095 519
rect 3099 515 3100 519
rect 3094 514 3100 515
rect 3222 519 3228 520
rect 3222 515 3223 519
rect 3227 515 3228 519
rect 3222 514 3228 515
rect 3350 519 3356 520
rect 3350 515 3351 519
rect 3355 515 3356 519
rect 3350 514 3356 515
rect 3478 519 3484 520
rect 3478 515 3479 519
rect 3483 515 3484 519
rect 3478 514 3484 515
rect 110 509 116 510
rect 110 505 111 509
rect 115 505 116 509
rect 110 504 116 505
rect 1822 509 1828 510
rect 1822 505 1823 509
rect 1827 505 1828 509
rect 1822 504 1828 505
rect 1862 509 1868 510
rect 1862 505 1863 509
rect 1867 505 1868 509
rect 1862 504 1868 505
rect 3574 509 3580 510
rect 3574 505 3575 509
rect 3579 505 3580 509
rect 3574 504 3580 505
rect 110 492 116 493
rect 110 488 111 492
rect 115 488 116 492
rect 110 487 116 488
rect 1822 492 1828 493
rect 1822 488 1823 492
rect 1827 488 1828 492
rect 1822 487 1828 488
rect 1862 492 1868 493
rect 1862 488 1863 492
rect 1867 488 1868 492
rect 1862 487 1868 488
rect 3574 492 3580 493
rect 3574 488 3575 492
rect 3579 488 3580 492
rect 3574 487 3580 488
rect 142 479 148 480
rect 142 475 143 479
rect 147 475 148 479
rect 142 474 148 475
rect 310 479 316 480
rect 310 475 311 479
rect 315 475 316 479
rect 310 474 316 475
rect 502 479 508 480
rect 502 475 503 479
rect 507 475 508 479
rect 502 474 508 475
rect 686 479 692 480
rect 686 475 687 479
rect 691 475 692 479
rect 686 474 692 475
rect 870 479 876 480
rect 870 475 871 479
rect 875 475 876 479
rect 870 474 876 475
rect 1038 479 1044 480
rect 1038 475 1039 479
rect 1043 475 1044 479
rect 1038 474 1044 475
rect 1198 479 1204 480
rect 1198 475 1199 479
rect 1203 475 1204 479
rect 1198 474 1204 475
rect 1358 479 1364 480
rect 1358 475 1359 479
rect 1363 475 1364 479
rect 1358 474 1364 475
rect 1510 479 1516 480
rect 1510 475 1511 479
rect 1515 475 1516 479
rect 1510 474 1516 475
rect 1670 479 1676 480
rect 1670 475 1671 479
rect 1675 475 1676 479
rect 1670 474 1676 475
rect 2310 479 2316 480
rect 2310 475 2311 479
rect 2315 475 2316 479
rect 2310 474 2316 475
rect 2406 479 2412 480
rect 2406 475 2407 479
rect 2411 475 2412 479
rect 2406 474 2412 475
rect 2510 479 2516 480
rect 2510 475 2511 479
rect 2515 475 2516 479
rect 2510 474 2516 475
rect 2614 479 2620 480
rect 2614 475 2615 479
rect 2619 475 2620 479
rect 2614 474 2620 475
rect 2726 479 2732 480
rect 2726 475 2727 479
rect 2731 475 2732 479
rect 2726 474 2732 475
rect 2846 479 2852 480
rect 2846 475 2847 479
rect 2851 475 2852 479
rect 2846 474 2852 475
rect 2974 479 2980 480
rect 2974 475 2975 479
rect 2979 475 2980 479
rect 2974 474 2980 475
rect 3102 479 3108 480
rect 3102 475 3103 479
rect 3107 475 3108 479
rect 3102 474 3108 475
rect 3230 479 3236 480
rect 3230 475 3231 479
rect 3235 475 3236 479
rect 3230 474 3236 475
rect 3358 479 3364 480
rect 3358 475 3359 479
rect 3363 475 3364 479
rect 3358 474 3364 475
rect 3486 479 3492 480
rect 3486 475 3487 479
rect 3491 475 3492 479
rect 3486 474 3492 475
rect 2238 445 2244 446
rect 142 441 148 442
rect 142 437 143 441
rect 147 437 148 441
rect 142 436 148 437
rect 302 441 308 442
rect 302 437 303 441
rect 307 437 308 441
rect 302 436 308 437
rect 494 441 500 442
rect 494 437 495 441
rect 499 437 500 441
rect 494 436 500 437
rect 686 441 692 442
rect 686 437 687 441
rect 691 437 692 441
rect 686 436 692 437
rect 878 441 884 442
rect 878 437 879 441
rect 883 437 884 441
rect 878 436 884 437
rect 1054 441 1060 442
rect 1054 437 1055 441
rect 1059 437 1060 441
rect 1054 436 1060 437
rect 1222 441 1228 442
rect 1222 437 1223 441
rect 1227 437 1228 441
rect 1222 436 1228 437
rect 1390 441 1396 442
rect 1390 437 1391 441
rect 1395 437 1396 441
rect 1390 436 1396 437
rect 1558 441 1564 442
rect 1558 437 1559 441
rect 1563 437 1564 441
rect 1558 436 1564 437
rect 1726 441 1732 442
rect 1726 437 1727 441
rect 1731 437 1732 441
rect 2238 441 2239 445
rect 2243 441 2244 445
rect 2238 440 2244 441
rect 2326 445 2332 446
rect 2326 441 2327 445
rect 2331 441 2332 445
rect 2326 440 2332 441
rect 2430 445 2436 446
rect 2430 441 2431 445
rect 2435 441 2436 445
rect 2430 440 2436 441
rect 2558 445 2564 446
rect 2558 441 2559 445
rect 2563 441 2564 445
rect 2558 440 2564 441
rect 2694 445 2700 446
rect 2694 441 2695 445
rect 2699 441 2700 445
rect 2694 440 2700 441
rect 2846 445 2852 446
rect 2846 441 2847 445
rect 2851 441 2852 445
rect 2846 440 2852 441
rect 2998 445 3004 446
rect 2998 441 2999 445
rect 3003 441 3004 445
rect 2998 440 3004 441
rect 3158 445 3164 446
rect 3158 441 3159 445
rect 3163 441 3164 445
rect 3158 440 3164 441
rect 3326 445 3332 446
rect 3326 441 3327 445
rect 3331 441 3332 445
rect 3326 440 3332 441
rect 3486 445 3492 446
rect 3486 441 3487 445
rect 3491 441 3492 445
rect 3486 440 3492 441
rect 1726 436 1732 437
rect 1862 432 1868 433
rect 110 428 116 429
rect 110 424 111 428
rect 115 424 116 428
rect 110 423 116 424
rect 1822 428 1828 429
rect 1822 424 1823 428
rect 1827 424 1828 428
rect 1862 428 1863 432
rect 1867 428 1868 432
rect 1862 427 1868 428
rect 3574 432 3580 433
rect 3574 428 3575 432
rect 3579 428 3580 432
rect 3574 427 3580 428
rect 1822 423 1828 424
rect 1862 415 1868 416
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 110 406 116 407
rect 1822 411 1828 412
rect 1822 407 1823 411
rect 1827 407 1828 411
rect 1862 411 1863 415
rect 1867 411 1868 415
rect 1862 410 1868 411
rect 3574 415 3580 416
rect 3574 411 3575 415
rect 3579 411 3580 415
rect 3574 410 3580 411
rect 1822 406 1828 407
rect 2230 405 2236 406
rect 134 401 140 402
rect 134 397 135 401
rect 139 397 140 401
rect 134 396 140 397
rect 294 401 300 402
rect 294 397 295 401
rect 299 397 300 401
rect 294 396 300 397
rect 486 401 492 402
rect 486 397 487 401
rect 491 397 492 401
rect 486 396 492 397
rect 678 401 684 402
rect 678 397 679 401
rect 683 397 684 401
rect 678 396 684 397
rect 870 401 876 402
rect 870 397 871 401
rect 875 397 876 401
rect 870 396 876 397
rect 1046 401 1052 402
rect 1046 397 1047 401
rect 1051 397 1052 401
rect 1046 396 1052 397
rect 1214 401 1220 402
rect 1214 397 1215 401
rect 1219 397 1220 401
rect 1214 396 1220 397
rect 1382 401 1388 402
rect 1382 397 1383 401
rect 1387 397 1388 401
rect 1382 396 1388 397
rect 1550 401 1556 402
rect 1550 397 1551 401
rect 1555 397 1556 401
rect 1550 396 1556 397
rect 1718 401 1724 402
rect 1718 397 1719 401
rect 1723 397 1724 401
rect 2230 401 2231 405
rect 2235 401 2236 405
rect 2230 400 2236 401
rect 2318 405 2324 406
rect 2318 401 2319 405
rect 2323 401 2324 405
rect 2318 400 2324 401
rect 2422 405 2428 406
rect 2422 401 2423 405
rect 2427 401 2428 405
rect 2422 400 2428 401
rect 2550 405 2556 406
rect 2550 401 2551 405
rect 2555 401 2556 405
rect 2550 400 2556 401
rect 2686 405 2692 406
rect 2686 401 2687 405
rect 2691 401 2692 405
rect 2686 400 2692 401
rect 2838 405 2844 406
rect 2838 401 2839 405
rect 2843 401 2844 405
rect 2838 400 2844 401
rect 2990 405 2996 406
rect 2990 401 2991 405
rect 2995 401 2996 405
rect 2990 400 2996 401
rect 3150 405 3156 406
rect 3150 401 3151 405
rect 3155 401 3156 405
rect 3150 400 3156 401
rect 3318 405 3324 406
rect 3318 401 3319 405
rect 3323 401 3324 405
rect 3318 400 3324 401
rect 3478 405 3484 406
rect 3478 401 3479 405
rect 3483 401 3484 405
rect 3478 400 3484 401
rect 1718 396 1724 397
rect 2182 383 2188 384
rect 134 379 140 380
rect 134 375 135 379
rect 139 375 140 379
rect 134 374 140 375
rect 262 379 268 380
rect 262 375 263 379
rect 267 375 268 379
rect 262 374 268 375
rect 422 379 428 380
rect 422 375 423 379
rect 427 375 428 379
rect 422 374 428 375
rect 590 379 596 380
rect 590 375 591 379
rect 595 375 596 379
rect 590 374 596 375
rect 766 379 772 380
rect 766 375 767 379
rect 771 375 772 379
rect 766 374 772 375
rect 934 379 940 380
rect 934 375 935 379
rect 939 375 940 379
rect 934 374 940 375
rect 1102 379 1108 380
rect 1102 375 1103 379
rect 1107 375 1108 379
rect 1102 374 1108 375
rect 1262 379 1268 380
rect 1262 375 1263 379
rect 1267 375 1268 379
rect 1262 374 1268 375
rect 1422 379 1428 380
rect 1422 375 1423 379
rect 1427 375 1428 379
rect 1422 374 1428 375
rect 1582 379 1588 380
rect 1582 375 1583 379
rect 1587 375 1588 379
rect 1582 374 1588 375
rect 1726 379 1732 380
rect 1726 375 1727 379
rect 1731 375 1732 379
rect 2182 379 2183 383
rect 2187 379 2188 383
rect 2182 378 2188 379
rect 2286 383 2292 384
rect 2286 379 2287 383
rect 2291 379 2292 383
rect 2286 378 2292 379
rect 2398 383 2404 384
rect 2398 379 2399 383
rect 2403 379 2404 383
rect 2398 378 2404 379
rect 2526 383 2532 384
rect 2526 379 2527 383
rect 2531 379 2532 383
rect 2526 378 2532 379
rect 2670 383 2676 384
rect 2670 379 2671 383
rect 2675 379 2676 383
rect 2670 378 2676 379
rect 2814 383 2820 384
rect 2814 379 2815 383
rect 2819 379 2820 383
rect 2814 378 2820 379
rect 2966 383 2972 384
rect 2966 379 2967 383
rect 2971 379 2972 383
rect 2966 378 2972 379
rect 3126 383 3132 384
rect 3126 379 3127 383
rect 3131 379 3132 383
rect 3126 378 3132 379
rect 3294 383 3300 384
rect 3294 379 3295 383
rect 3299 379 3300 383
rect 3294 378 3300 379
rect 3462 383 3468 384
rect 3462 379 3463 383
rect 3467 379 3468 383
rect 3462 378 3468 379
rect 1726 374 1732 375
rect 1862 373 1868 374
rect 110 369 116 370
rect 110 365 111 369
rect 115 365 116 369
rect 110 364 116 365
rect 1822 369 1828 370
rect 1822 365 1823 369
rect 1827 365 1828 369
rect 1862 369 1863 373
rect 1867 369 1868 373
rect 1862 368 1868 369
rect 3574 373 3580 374
rect 3574 369 3575 373
rect 3579 369 3580 373
rect 3574 368 3580 369
rect 1822 364 1828 365
rect 1862 356 1868 357
rect 110 352 116 353
rect 110 348 111 352
rect 115 348 116 352
rect 110 347 116 348
rect 1822 352 1828 353
rect 1822 348 1823 352
rect 1827 348 1828 352
rect 1862 352 1863 356
rect 1867 352 1868 356
rect 1862 351 1868 352
rect 3574 356 3580 357
rect 3574 352 3575 356
rect 3579 352 3580 356
rect 3574 351 3580 352
rect 1822 347 1828 348
rect 2190 343 2196 344
rect 142 339 148 340
rect 142 335 143 339
rect 147 335 148 339
rect 142 334 148 335
rect 270 339 276 340
rect 270 335 271 339
rect 275 335 276 339
rect 270 334 276 335
rect 430 339 436 340
rect 430 335 431 339
rect 435 335 436 339
rect 430 334 436 335
rect 598 339 604 340
rect 598 335 599 339
rect 603 335 604 339
rect 598 334 604 335
rect 774 339 780 340
rect 774 335 775 339
rect 779 335 780 339
rect 774 334 780 335
rect 942 339 948 340
rect 942 335 943 339
rect 947 335 948 339
rect 942 334 948 335
rect 1110 339 1116 340
rect 1110 335 1111 339
rect 1115 335 1116 339
rect 1110 334 1116 335
rect 1270 339 1276 340
rect 1270 335 1271 339
rect 1275 335 1276 339
rect 1270 334 1276 335
rect 1430 339 1436 340
rect 1430 335 1431 339
rect 1435 335 1436 339
rect 1430 334 1436 335
rect 1590 339 1596 340
rect 1590 335 1591 339
rect 1595 335 1596 339
rect 1590 334 1596 335
rect 1734 339 1740 340
rect 1734 335 1735 339
rect 1739 335 1740 339
rect 2190 339 2191 343
rect 2195 339 2196 343
rect 2190 338 2196 339
rect 2294 343 2300 344
rect 2294 339 2295 343
rect 2299 339 2300 343
rect 2294 338 2300 339
rect 2406 343 2412 344
rect 2406 339 2407 343
rect 2411 339 2412 343
rect 2406 338 2412 339
rect 2534 343 2540 344
rect 2534 339 2535 343
rect 2539 339 2540 343
rect 2534 338 2540 339
rect 2678 343 2684 344
rect 2678 339 2679 343
rect 2683 339 2684 343
rect 2678 338 2684 339
rect 2822 343 2828 344
rect 2822 339 2823 343
rect 2827 339 2828 343
rect 2822 338 2828 339
rect 2974 343 2980 344
rect 2974 339 2975 343
rect 2979 339 2980 343
rect 2974 338 2980 339
rect 3134 343 3140 344
rect 3134 339 3135 343
rect 3139 339 3140 343
rect 3134 338 3140 339
rect 3302 343 3308 344
rect 3302 339 3303 343
rect 3307 339 3308 343
rect 3302 338 3308 339
rect 3470 343 3476 344
rect 3470 339 3471 343
rect 3475 339 3476 343
rect 3470 338 3476 339
rect 1734 334 1740 335
rect 214 305 220 306
rect 214 301 215 305
rect 219 301 220 305
rect 214 300 220 301
rect 350 305 356 306
rect 350 301 351 305
rect 355 301 356 305
rect 350 300 356 301
rect 494 305 500 306
rect 494 301 495 305
rect 499 301 500 305
rect 494 300 500 301
rect 638 305 644 306
rect 638 301 639 305
rect 643 301 644 305
rect 638 300 644 301
rect 790 305 796 306
rect 790 301 791 305
rect 795 301 796 305
rect 790 300 796 301
rect 934 305 940 306
rect 934 301 935 305
rect 939 301 940 305
rect 934 300 940 301
rect 1078 305 1084 306
rect 1078 301 1079 305
rect 1083 301 1084 305
rect 1078 300 1084 301
rect 1222 305 1228 306
rect 1222 301 1223 305
rect 1227 301 1228 305
rect 1222 300 1228 301
rect 1358 305 1364 306
rect 1358 301 1359 305
rect 1363 301 1364 305
rect 1358 300 1364 301
rect 1486 305 1492 306
rect 1486 301 1487 305
rect 1491 301 1492 305
rect 1486 300 1492 301
rect 1622 305 1628 306
rect 1622 301 1623 305
rect 1627 301 1628 305
rect 1622 300 1628 301
rect 1734 305 1740 306
rect 1734 301 1735 305
rect 1739 301 1740 305
rect 1734 300 1740 301
rect 1894 301 1900 302
rect 1894 297 1895 301
rect 1899 297 1900 301
rect 1894 296 1900 297
rect 2086 301 2092 302
rect 2086 297 2087 301
rect 2091 297 2092 301
rect 2086 296 2092 297
rect 2302 301 2308 302
rect 2302 297 2303 301
rect 2307 297 2308 301
rect 2302 296 2308 297
rect 2510 301 2516 302
rect 2510 297 2511 301
rect 2515 297 2516 301
rect 2510 296 2516 297
rect 2710 301 2716 302
rect 2710 297 2711 301
rect 2715 297 2716 301
rect 2710 296 2716 297
rect 2902 301 2908 302
rect 2902 297 2903 301
rect 2907 297 2908 301
rect 2902 296 2908 297
rect 3094 301 3100 302
rect 3094 297 3095 301
rect 3099 297 3100 301
rect 3094 296 3100 297
rect 3294 301 3300 302
rect 3294 297 3295 301
rect 3299 297 3300 301
rect 3294 296 3300 297
rect 3486 301 3492 302
rect 3486 297 3487 301
rect 3491 297 3492 301
rect 3486 296 3492 297
rect 110 292 116 293
rect 110 288 111 292
rect 115 288 116 292
rect 110 287 116 288
rect 1822 292 1828 293
rect 1822 288 1823 292
rect 1827 288 1828 292
rect 1822 287 1828 288
rect 1862 288 1868 289
rect 1862 284 1863 288
rect 1867 284 1868 288
rect 1862 283 1868 284
rect 3574 288 3580 289
rect 3574 284 3575 288
rect 3579 284 3580 288
rect 3574 283 3580 284
rect 110 275 116 276
rect 110 271 111 275
rect 115 271 116 275
rect 110 270 116 271
rect 1822 275 1828 276
rect 1822 271 1823 275
rect 1827 271 1828 275
rect 1822 270 1828 271
rect 1862 271 1868 272
rect 1862 267 1863 271
rect 1867 267 1868 271
rect 1862 266 1868 267
rect 3574 271 3580 272
rect 3574 267 3575 271
rect 3579 267 3580 271
rect 3574 266 3580 267
rect 206 265 212 266
rect 206 261 207 265
rect 211 261 212 265
rect 206 260 212 261
rect 342 265 348 266
rect 342 261 343 265
rect 347 261 348 265
rect 342 260 348 261
rect 486 265 492 266
rect 486 261 487 265
rect 491 261 492 265
rect 486 260 492 261
rect 630 265 636 266
rect 630 261 631 265
rect 635 261 636 265
rect 630 260 636 261
rect 782 265 788 266
rect 782 261 783 265
rect 787 261 788 265
rect 782 260 788 261
rect 926 265 932 266
rect 926 261 927 265
rect 931 261 932 265
rect 926 260 932 261
rect 1070 265 1076 266
rect 1070 261 1071 265
rect 1075 261 1076 265
rect 1070 260 1076 261
rect 1214 265 1220 266
rect 1214 261 1215 265
rect 1219 261 1220 265
rect 1214 260 1220 261
rect 1350 265 1356 266
rect 1350 261 1351 265
rect 1355 261 1356 265
rect 1350 260 1356 261
rect 1478 265 1484 266
rect 1478 261 1479 265
rect 1483 261 1484 265
rect 1478 260 1484 261
rect 1614 265 1620 266
rect 1614 261 1615 265
rect 1619 261 1620 265
rect 1614 260 1620 261
rect 1726 265 1732 266
rect 1726 261 1727 265
rect 1731 261 1732 265
rect 1726 260 1732 261
rect 1886 261 1892 262
rect 1886 257 1887 261
rect 1891 257 1892 261
rect 1886 256 1892 257
rect 2078 261 2084 262
rect 2078 257 2079 261
rect 2083 257 2084 261
rect 2078 256 2084 257
rect 2294 261 2300 262
rect 2294 257 2295 261
rect 2299 257 2300 261
rect 2294 256 2300 257
rect 2502 261 2508 262
rect 2502 257 2503 261
rect 2507 257 2508 261
rect 2502 256 2508 257
rect 2702 261 2708 262
rect 2702 257 2703 261
rect 2707 257 2708 261
rect 2702 256 2708 257
rect 2894 261 2900 262
rect 2894 257 2895 261
rect 2899 257 2900 261
rect 2894 256 2900 257
rect 3086 261 3092 262
rect 3086 257 3087 261
rect 3091 257 3092 261
rect 3086 256 3092 257
rect 3286 261 3292 262
rect 3286 257 3287 261
rect 3291 257 3292 261
rect 3286 256 3292 257
rect 3478 261 3484 262
rect 3478 257 3479 261
rect 3483 257 3484 261
rect 3478 256 3484 257
rect 1886 239 1892 240
rect 230 235 236 236
rect 230 231 231 235
rect 235 231 236 235
rect 230 230 236 231
rect 358 235 364 236
rect 358 231 359 235
rect 363 231 364 235
rect 358 230 364 231
rect 486 235 492 236
rect 486 231 487 235
rect 491 231 492 235
rect 486 230 492 231
rect 622 235 628 236
rect 622 231 623 235
rect 627 231 628 235
rect 622 230 628 231
rect 758 235 764 236
rect 758 231 759 235
rect 763 231 764 235
rect 758 230 764 231
rect 894 235 900 236
rect 894 231 895 235
rect 899 231 900 235
rect 894 230 900 231
rect 1030 235 1036 236
rect 1030 231 1031 235
rect 1035 231 1036 235
rect 1030 230 1036 231
rect 1158 235 1164 236
rect 1158 231 1159 235
rect 1163 231 1164 235
rect 1158 230 1164 231
rect 1294 235 1300 236
rect 1294 231 1295 235
rect 1299 231 1300 235
rect 1294 230 1300 231
rect 1430 235 1436 236
rect 1430 231 1431 235
rect 1435 231 1436 235
rect 1886 235 1887 239
rect 1891 235 1892 239
rect 1886 234 1892 235
rect 1998 239 2004 240
rect 1998 235 1999 239
rect 2003 235 2004 239
rect 1998 234 2004 235
rect 2142 239 2148 240
rect 2142 235 2143 239
rect 2147 235 2148 239
rect 2142 234 2148 235
rect 2294 239 2300 240
rect 2294 235 2295 239
rect 2299 235 2300 239
rect 2294 234 2300 235
rect 2454 239 2460 240
rect 2454 235 2455 239
rect 2459 235 2460 239
rect 2454 234 2460 235
rect 2614 239 2620 240
rect 2614 235 2615 239
rect 2619 235 2620 239
rect 2614 234 2620 235
rect 2782 239 2788 240
rect 2782 235 2783 239
rect 2787 235 2788 239
rect 2782 234 2788 235
rect 2950 239 2956 240
rect 2950 235 2951 239
rect 2955 235 2956 239
rect 2950 234 2956 235
rect 3126 239 3132 240
rect 3126 235 3127 239
rect 3131 235 3132 239
rect 3126 234 3132 235
rect 3310 239 3316 240
rect 3310 235 3311 239
rect 3315 235 3316 239
rect 3310 234 3316 235
rect 3478 239 3484 240
rect 3478 235 3479 239
rect 3483 235 3484 239
rect 3478 234 3484 235
rect 1430 230 1436 231
rect 1862 229 1868 230
rect 110 225 116 226
rect 110 221 111 225
rect 115 221 116 225
rect 110 220 116 221
rect 1822 225 1828 226
rect 1822 221 1823 225
rect 1827 221 1828 225
rect 1862 225 1863 229
rect 1867 225 1868 229
rect 1862 224 1868 225
rect 3574 229 3580 230
rect 3574 225 3575 229
rect 3579 225 3580 229
rect 3574 224 3580 225
rect 1822 220 1828 221
rect 1862 212 1868 213
rect 110 208 116 209
rect 110 204 111 208
rect 115 204 116 208
rect 110 203 116 204
rect 1822 208 1828 209
rect 1822 204 1823 208
rect 1827 204 1828 208
rect 1862 208 1863 212
rect 1867 208 1868 212
rect 1862 207 1868 208
rect 3574 212 3580 213
rect 3574 208 3575 212
rect 3579 208 3580 212
rect 3574 207 3580 208
rect 1822 203 1828 204
rect 1894 199 1900 200
rect 238 195 244 196
rect 238 191 239 195
rect 243 191 244 195
rect 238 190 244 191
rect 366 195 372 196
rect 366 191 367 195
rect 371 191 372 195
rect 366 190 372 191
rect 494 195 500 196
rect 494 191 495 195
rect 499 191 500 195
rect 494 190 500 191
rect 630 195 636 196
rect 630 191 631 195
rect 635 191 636 195
rect 630 190 636 191
rect 766 195 772 196
rect 766 191 767 195
rect 771 191 772 195
rect 766 190 772 191
rect 902 195 908 196
rect 902 191 903 195
rect 907 191 908 195
rect 902 190 908 191
rect 1038 195 1044 196
rect 1038 191 1039 195
rect 1043 191 1044 195
rect 1038 190 1044 191
rect 1166 195 1172 196
rect 1166 191 1167 195
rect 1171 191 1172 195
rect 1166 190 1172 191
rect 1302 195 1308 196
rect 1302 191 1303 195
rect 1307 191 1308 195
rect 1302 190 1308 191
rect 1438 195 1444 196
rect 1438 191 1439 195
rect 1443 191 1444 195
rect 1894 195 1895 199
rect 1899 195 1900 199
rect 1894 194 1900 195
rect 2006 199 2012 200
rect 2006 195 2007 199
rect 2011 195 2012 199
rect 2006 194 2012 195
rect 2150 199 2156 200
rect 2150 195 2151 199
rect 2155 195 2156 199
rect 2150 194 2156 195
rect 2302 199 2308 200
rect 2302 195 2303 199
rect 2307 195 2308 199
rect 2302 194 2308 195
rect 2462 199 2468 200
rect 2462 195 2463 199
rect 2467 195 2468 199
rect 2462 194 2468 195
rect 2622 199 2628 200
rect 2622 195 2623 199
rect 2627 195 2628 199
rect 2622 194 2628 195
rect 2790 199 2796 200
rect 2790 195 2791 199
rect 2795 195 2796 199
rect 2790 194 2796 195
rect 2958 199 2964 200
rect 2958 195 2959 199
rect 2963 195 2964 199
rect 2958 194 2964 195
rect 3134 199 3140 200
rect 3134 195 3135 199
rect 3139 195 3140 199
rect 3134 194 3140 195
rect 3318 199 3324 200
rect 3318 195 3319 199
rect 3323 195 3324 199
rect 3318 194 3324 195
rect 3486 199 3492 200
rect 3486 195 3487 199
rect 3491 195 3492 199
rect 3486 194 3492 195
rect 1438 190 1444 191
rect 174 137 180 138
rect 174 133 175 137
rect 179 133 180 137
rect 174 132 180 133
rect 262 137 268 138
rect 262 133 263 137
rect 267 133 268 137
rect 262 132 268 133
rect 350 137 356 138
rect 350 133 351 137
rect 355 133 356 137
rect 350 132 356 133
rect 438 137 444 138
rect 438 133 439 137
rect 443 133 444 137
rect 438 132 444 133
rect 526 137 532 138
rect 526 133 527 137
rect 531 133 532 137
rect 526 132 532 133
rect 614 137 620 138
rect 614 133 615 137
rect 619 133 620 137
rect 614 132 620 133
rect 702 137 708 138
rect 702 133 703 137
rect 707 133 708 137
rect 702 132 708 133
rect 790 137 796 138
rect 790 133 791 137
rect 795 133 796 137
rect 790 132 796 133
rect 878 137 884 138
rect 878 133 879 137
rect 883 133 884 137
rect 878 132 884 133
rect 966 137 972 138
rect 966 133 967 137
rect 971 133 972 137
rect 966 132 972 133
rect 1054 137 1060 138
rect 1054 133 1055 137
rect 1059 133 1060 137
rect 1054 132 1060 133
rect 1142 137 1148 138
rect 1142 133 1143 137
rect 1147 133 1148 137
rect 1142 132 1148 133
rect 1230 137 1236 138
rect 1230 133 1231 137
rect 1235 133 1236 137
rect 1230 132 1236 133
rect 1318 137 1324 138
rect 1318 133 1319 137
rect 1323 133 1324 137
rect 1318 132 1324 133
rect 1406 137 1412 138
rect 1406 133 1407 137
rect 1411 133 1412 137
rect 1406 132 1412 133
rect 1502 137 1508 138
rect 1502 133 1503 137
rect 1507 133 1508 137
rect 1502 132 1508 133
rect 1894 137 1900 138
rect 1894 133 1895 137
rect 1899 133 1900 137
rect 1894 132 1900 133
rect 1982 137 1988 138
rect 1982 133 1983 137
rect 1987 133 1988 137
rect 1982 132 1988 133
rect 2070 137 2076 138
rect 2070 133 2071 137
rect 2075 133 2076 137
rect 2070 132 2076 133
rect 2158 137 2164 138
rect 2158 133 2159 137
rect 2163 133 2164 137
rect 2158 132 2164 133
rect 2246 137 2252 138
rect 2246 133 2247 137
rect 2251 133 2252 137
rect 2246 132 2252 133
rect 2334 137 2340 138
rect 2334 133 2335 137
rect 2339 133 2340 137
rect 2334 132 2340 133
rect 2438 137 2444 138
rect 2438 133 2439 137
rect 2443 133 2444 137
rect 2438 132 2444 133
rect 2542 137 2548 138
rect 2542 133 2543 137
rect 2547 133 2548 137
rect 2542 132 2548 133
rect 2646 137 2652 138
rect 2646 133 2647 137
rect 2651 133 2652 137
rect 2646 132 2652 133
rect 2742 137 2748 138
rect 2742 133 2743 137
rect 2747 133 2748 137
rect 2742 132 2748 133
rect 2838 137 2844 138
rect 2838 133 2839 137
rect 2843 133 2844 137
rect 2838 132 2844 133
rect 2934 137 2940 138
rect 2934 133 2935 137
rect 2939 133 2940 137
rect 2934 132 2940 133
rect 3030 137 3036 138
rect 3030 133 3031 137
rect 3035 133 3036 137
rect 3030 132 3036 133
rect 3126 137 3132 138
rect 3126 133 3127 137
rect 3131 133 3132 137
rect 3126 132 3132 133
rect 3222 137 3228 138
rect 3222 133 3223 137
rect 3227 133 3228 137
rect 3222 132 3228 133
rect 3310 137 3316 138
rect 3310 133 3311 137
rect 3315 133 3316 137
rect 3310 132 3316 133
rect 3398 137 3404 138
rect 3398 133 3399 137
rect 3403 133 3404 137
rect 3398 132 3404 133
rect 3486 137 3492 138
rect 3486 133 3487 137
rect 3491 133 3492 137
rect 3486 132 3492 133
rect 110 124 116 125
rect 110 120 111 124
rect 115 120 116 124
rect 110 119 116 120
rect 1822 124 1828 125
rect 1822 120 1823 124
rect 1827 120 1828 124
rect 1822 119 1828 120
rect 1862 124 1868 125
rect 1862 120 1863 124
rect 1867 120 1868 124
rect 1862 119 1868 120
rect 3574 124 3580 125
rect 3574 120 3575 124
rect 3579 120 3580 124
rect 3574 119 3580 120
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 110 102 116 103
rect 1822 107 1828 108
rect 1822 103 1823 107
rect 1827 103 1828 107
rect 1822 102 1828 103
rect 1862 107 1868 108
rect 1862 103 1863 107
rect 1867 103 1868 107
rect 1862 102 1868 103
rect 3574 107 3580 108
rect 3574 103 3575 107
rect 3579 103 3580 107
rect 3574 102 3580 103
rect 166 97 172 98
rect 166 93 167 97
rect 171 93 172 97
rect 166 92 172 93
rect 254 97 260 98
rect 254 93 255 97
rect 259 93 260 97
rect 254 92 260 93
rect 342 97 348 98
rect 342 93 343 97
rect 347 93 348 97
rect 342 92 348 93
rect 430 97 436 98
rect 430 93 431 97
rect 435 93 436 97
rect 430 92 436 93
rect 518 97 524 98
rect 518 93 519 97
rect 523 93 524 97
rect 518 92 524 93
rect 606 97 612 98
rect 606 93 607 97
rect 611 93 612 97
rect 606 92 612 93
rect 694 97 700 98
rect 694 93 695 97
rect 699 93 700 97
rect 694 92 700 93
rect 782 97 788 98
rect 782 93 783 97
rect 787 93 788 97
rect 782 92 788 93
rect 870 97 876 98
rect 870 93 871 97
rect 875 93 876 97
rect 870 92 876 93
rect 958 97 964 98
rect 958 93 959 97
rect 963 93 964 97
rect 958 92 964 93
rect 1046 97 1052 98
rect 1046 93 1047 97
rect 1051 93 1052 97
rect 1046 92 1052 93
rect 1134 97 1140 98
rect 1134 93 1135 97
rect 1139 93 1140 97
rect 1134 92 1140 93
rect 1222 97 1228 98
rect 1222 93 1223 97
rect 1227 93 1228 97
rect 1222 92 1228 93
rect 1310 97 1316 98
rect 1310 93 1311 97
rect 1315 93 1316 97
rect 1310 92 1316 93
rect 1398 97 1404 98
rect 1398 93 1399 97
rect 1403 93 1404 97
rect 1398 92 1404 93
rect 1494 97 1500 98
rect 1494 93 1495 97
rect 1499 93 1500 97
rect 1494 92 1500 93
rect 1886 97 1892 98
rect 1886 93 1887 97
rect 1891 93 1892 97
rect 1886 92 1892 93
rect 1974 97 1980 98
rect 1974 93 1975 97
rect 1979 93 1980 97
rect 1974 92 1980 93
rect 2062 97 2068 98
rect 2062 93 2063 97
rect 2067 93 2068 97
rect 2062 92 2068 93
rect 2150 97 2156 98
rect 2150 93 2151 97
rect 2155 93 2156 97
rect 2150 92 2156 93
rect 2238 97 2244 98
rect 2238 93 2239 97
rect 2243 93 2244 97
rect 2238 92 2244 93
rect 2326 97 2332 98
rect 2326 93 2327 97
rect 2331 93 2332 97
rect 2326 92 2332 93
rect 2430 97 2436 98
rect 2430 93 2431 97
rect 2435 93 2436 97
rect 2430 92 2436 93
rect 2534 97 2540 98
rect 2534 93 2535 97
rect 2539 93 2540 97
rect 2534 92 2540 93
rect 2638 97 2644 98
rect 2638 93 2639 97
rect 2643 93 2644 97
rect 2638 92 2644 93
rect 2734 97 2740 98
rect 2734 93 2735 97
rect 2739 93 2740 97
rect 2734 92 2740 93
rect 2830 97 2836 98
rect 2830 93 2831 97
rect 2835 93 2836 97
rect 2830 92 2836 93
rect 2926 97 2932 98
rect 2926 93 2927 97
rect 2931 93 2932 97
rect 2926 92 2932 93
rect 3022 97 3028 98
rect 3022 93 3023 97
rect 3027 93 3028 97
rect 3022 92 3028 93
rect 3118 97 3124 98
rect 3118 93 3119 97
rect 3123 93 3124 97
rect 3118 92 3124 93
rect 3214 97 3220 98
rect 3214 93 3215 97
rect 3219 93 3220 97
rect 3214 92 3220 93
rect 3302 97 3308 98
rect 3302 93 3303 97
rect 3307 93 3308 97
rect 3302 92 3308 93
rect 3390 97 3396 98
rect 3390 93 3391 97
rect 3395 93 3396 97
rect 3390 92 3396 93
rect 3478 97 3484 98
rect 3478 93 3479 97
rect 3483 93 3484 97
rect 3478 92 3484 93
<< m3c >>
rect 239 3629 243 3633
rect 327 3629 331 3633
rect 415 3629 419 3633
rect 503 3629 507 3633
rect 591 3629 595 3633
rect 679 3629 683 3633
rect 111 3616 115 3620
rect 1823 3616 1827 3620
rect 111 3599 115 3603
rect 1823 3599 1827 3603
rect 231 3589 235 3593
rect 319 3589 323 3593
rect 407 3589 411 3593
rect 495 3589 499 3593
rect 583 3589 587 3593
rect 671 3589 675 3593
rect 1887 3571 1891 3575
rect 1975 3571 1979 3575
rect 2063 3571 2067 3575
rect 2151 3571 2155 3575
rect 2239 3571 2243 3575
rect 2327 3571 2331 3575
rect 2415 3571 2419 3575
rect 2503 3571 2507 3575
rect 2591 3571 2595 3575
rect 2679 3571 2683 3575
rect 2767 3571 2771 3575
rect 2855 3571 2859 3575
rect 2943 3571 2947 3575
rect 3031 3571 3035 3575
rect 3119 3571 3123 3575
rect 3207 3571 3211 3575
rect 3295 3571 3299 3575
rect 247 3559 251 3563
rect 399 3559 403 3563
rect 543 3559 547 3563
rect 687 3559 691 3563
rect 823 3559 827 3563
rect 951 3559 955 3563
rect 1079 3559 1083 3563
rect 1199 3559 1203 3563
rect 1311 3559 1315 3563
rect 1423 3559 1427 3563
rect 1543 3559 1547 3563
rect 1863 3561 1867 3565
rect 3575 3561 3579 3565
rect 111 3549 115 3553
rect 1823 3549 1827 3553
rect 1863 3544 1867 3548
rect 3575 3544 3579 3548
rect 111 3532 115 3536
rect 1823 3532 1827 3536
rect 1895 3531 1899 3535
rect 1983 3531 1987 3535
rect 2071 3531 2075 3535
rect 2159 3531 2163 3535
rect 2247 3531 2251 3535
rect 2335 3531 2339 3535
rect 2423 3531 2427 3535
rect 2511 3531 2515 3535
rect 2599 3531 2603 3535
rect 2687 3531 2691 3535
rect 2775 3531 2779 3535
rect 2863 3531 2867 3535
rect 2951 3531 2955 3535
rect 3039 3531 3043 3535
rect 3127 3531 3131 3535
rect 3215 3531 3219 3535
rect 3303 3531 3307 3535
rect 255 3519 259 3523
rect 407 3519 411 3523
rect 551 3519 555 3523
rect 695 3519 699 3523
rect 831 3519 835 3523
rect 959 3519 963 3523
rect 1087 3519 1091 3523
rect 1207 3519 1211 3523
rect 1319 3519 1323 3523
rect 1431 3519 1435 3523
rect 1551 3519 1555 3523
rect 183 3485 187 3489
rect 351 3485 355 3489
rect 519 3485 523 3489
rect 679 3485 683 3489
rect 831 3485 835 3489
rect 967 3485 971 3489
rect 1095 3485 1099 3489
rect 1215 3485 1219 3489
rect 1335 3485 1339 3489
rect 1455 3485 1459 3489
rect 1575 3485 1579 3489
rect 1911 3489 1915 3493
rect 2015 3489 2019 3493
rect 2135 3489 2139 3493
rect 2263 3489 2267 3493
rect 2391 3489 2395 3493
rect 2527 3489 2531 3493
rect 2663 3489 2667 3493
rect 2799 3489 2803 3493
rect 2943 3489 2947 3493
rect 3087 3489 3091 3493
rect 111 3472 115 3476
rect 1823 3472 1827 3476
rect 1863 3476 1867 3480
rect 3575 3476 3579 3480
rect 111 3455 115 3459
rect 1823 3455 1827 3459
rect 1863 3459 1867 3463
rect 3575 3459 3579 3463
rect 175 3445 179 3449
rect 343 3445 347 3449
rect 511 3445 515 3449
rect 671 3445 675 3449
rect 823 3445 827 3449
rect 959 3445 963 3449
rect 1087 3445 1091 3449
rect 1207 3445 1211 3449
rect 1327 3445 1331 3449
rect 1447 3445 1451 3449
rect 1567 3445 1571 3449
rect 1903 3449 1907 3453
rect 2007 3449 2011 3453
rect 2127 3449 2131 3453
rect 2255 3449 2259 3453
rect 2383 3449 2387 3453
rect 2519 3449 2523 3453
rect 2655 3449 2659 3453
rect 2791 3449 2795 3453
rect 2935 3449 2939 3453
rect 3079 3449 3083 3453
rect 135 3423 139 3427
rect 255 3423 259 3427
rect 415 3423 419 3427
rect 583 3423 587 3427
rect 759 3423 763 3427
rect 935 3423 939 3427
rect 1111 3423 1115 3427
rect 1295 3423 1299 3427
rect 1479 3423 1483 3427
rect 1911 3419 1915 3423
rect 2071 3419 2075 3423
rect 2223 3419 2227 3423
rect 2367 3419 2371 3423
rect 2503 3419 2507 3423
rect 2631 3419 2635 3423
rect 2759 3419 2763 3423
rect 2887 3419 2891 3423
rect 3023 3419 3027 3423
rect 111 3413 115 3417
rect 1823 3413 1827 3417
rect 1863 3409 1867 3413
rect 3575 3409 3579 3413
rect 111 3396 115 3400
rect 1823 3396 1827 3400
rect 1863 3392 1867 3396
rect 3575 3392 3579 3396
rect 143 3383 147 3387
rect 263 3383 267 3387
rect 423 3383 427 3387
rect 591 3383 595 3387
rect 767 3383 771 3387
rect 943 3383 947 3387
rect 1119 3383 1123 3387
rect 1303 3383 1307 3387
rect 1487 3383 1491 3387
rect 1919 3379 1923 3383
rect 2079 3379 2083 3383
rect 2231 3379 2235 3383
rect 2375 3379 2379 3383
rect 2511 3379 2515 3383
rect 2639 3379 2643 3383
rect 2767 3379 2771 3383
rect 2895 3379 2899 3383
rect 3031 3379 3035 3383
rect 207 3341 211 3345
rect 367 3341 371 3345
rect 535 3341 539 3345
rect 695 3341 699 3345
rect 855 3341 859 3345
rect 999 3341 1003 3345
rect 1143 3341 1147 3345
rect 1279 3341 1283 3345
rect 1415 3341 1419 3345
rect 1559 3341 1563 3345
rect 1895 3341 1899 3345
rect 2047 3341 2051 3345
rect 2207 3341 2211 3345
rect 2367 3341 2371 3345
rect 2535 3341 2539 3345
rect 2703 3341 2707 3345
rect 2879 3341 2883 3345
rect 3055 3341 3059 3345
rect 111 3328 115 3332
rect 1823 3328 1827 3332
rect 1863 3328 1867 3332
rect 3575 3328 3579 3332
rect 111 3311 115 3315
rect 1823 3311 1827 3315
rect 1863 3311 1867 3315
rect 3575 3311 3579 3315
rect 199 3301 203 3305
rect 359 3301 363 3305
rect 527 3301 531 3305
rect 687 3301 691 3305
rect 847 3301 851 3305
rect 991 3301 995 3305
rect 1135 3301 1139 3305
rect 1271 3301 1275 3305
rect 1407 3301 1411 3305
rect 1551 3301 1555 3305
rect 1887 3301 1891 3305
rect 2039 3301 2043 3305
rect 2199 3301 2203 3305
rect 2359 3301 2363 3305
rect 2527 3301 2531 3305
rect 2695 3301 2699 3305
rect 2871 3301 2875 3305
rect 3047 3301 3051 3305
rect 255 3275 259 3279
rect 375 3275 379 3279
rect 511 3275 515 3279
rect 663 3275 667 3279
rect 823 3275 827 3279
rect 991 3275 995 3279
rect 1167 3275 1171 3279
rect 1343 3275 1347 3279
rect 1519 3275 1523 3279
rect 1887 3275 1891 3279
rect 2063 3275 2067 3279
rect 2263 3275 2267 3279
rect 2455 3275 2459 3279
rect 2639 3275 2643 3279
rect 2815 3275 2819 3279
rect 2983 3275 2987 3279
rect 3151 3275 3155 3279
rect 3319 3275 3323 3279
rect 3479 3275 3483 3279
rect 111 3265 115 3269
rect 1823 3265 1827 3269
rect 1863 3265 1867 3269
rect 3575 3265 3579 3269
rect 111 3248 115 3252
rect 1823 3248 1827 3252
rect 1863 3248 1867 3252
rect 3575 3248 3579 3252
rect 263 3235 267 3239
rect 383 3235 387 3239
rect 519 3235 523 3239
rect 671 3235 675 3239
rect 831 3235 835 3239
rect 999 3235 1003 3239
rect 1175 3235 1179 3239
rect 1351 3235 1355 3239
rect 1527 3235 1531 3239
rect 1895 3235 1899 3239
rect 2071 3235 2075 3239
rect 2271 3235 2275 3239
rect 2463 3235 2467 3239
rect 2647 3235 2651 3239
rect 2823 3235 2827 3239
rect 2991 3235 2995 3239
rect 3159 3235 3163 3239
rect 3327 3235 3331 3239
rect 3487 3235 3491 3239
rect 431 3197 435 3201
rect 551 3197 555 3201
rect 671 3197 675 3201
rect 799 3197 803 3201
rect 935 3197 939 3201
rect 1079 3197 1083 3201
rect 1231 3197 1235 3201
rect 1383 3197 1387 3201
rect 1535 3197 1539 3201
rect 1895 3201 1899 3205
rect 2087 3201 2091 3205
rect 2303 3201 2307 3205
rect 2511 3201 2515 3205
rect 2703 3201 2707 3205
rect 2879 3201 2883 3205
rect 3039 3201 3043 3205
rect 3199 3201 3203 3205
rect 3351 3201 3355 3205
rect 3487 3201 3491 3205
rect 111 3184 115 3188
rect 1823 3184 1827 3188
rect 1863 3188 1867 3192
rect 3575 3188 3579 3192
rect 111 3167 115 3171
rect 1823 3167 1827 3171
rect 1863 3171 1867 3175
rect 3575 3171 3579 3175
rect 423 3157 427 3161
rect 543 3157 547 3161
rect 663 3157 667 3161
rect 791 3157 795 3161
rect 927 3157 931 3161
rect 1071 3157 1075 3161
rect 1223 3157 1227 3161
rect 1375 3157 1379 3161
rect 1527 3157 1531 3161
rect 1887 3161 1891 3165
rect 2079 3161 2083 3165
rect 2295 3161 2299 3165
rect 2503 3161 2507 3165
rect 2695 3161 2699 3165
rect 2871 3161 2875 3165
rect 3031 3161 3035 3165
rect 3191 3161 3195 3165
rect 3343 3161 3347 3165
rect 3479 3161 3483 3165
rect 463 3131 467 3135
rect 551 3131 555 3135
rect 639 3131 643 3135
rect 735 3131 739 3135
rect 847 3131 851 3135
rect 967 3131 971 3135
rect 1095 3131 1099 3135
rect 1231 3131 1235 3135
rect 1375 3131 1379 3135
rect 1519 3131 1523 3135
rect 1887 3135 1891 3139
rect 2079 3135 2083 3139
rect 2295 3135 2299 3139
rect 2503 3135 2507 3139
rect 2695 3135 2699 3139
rect 2871 3135 2875 3139
rect 3039 3135 3043 3139
rect 3191 3135 3195 3139
rect 3343 3135 3347 3139
rect 3479 3135 3483 3139
rect 111 3121 115 3125
rect 1823 3121 1827 3125
rect 1863 3125 1867 3129
rect 3575 3125 3579 3129
rect 111 3104 115 3108
rect 1823 3104 1827 3108
rect 1863 3108 1867 3112
rect 3575 3108 3579 3112
rect 471 3091 475 3095
rect 559 3091 563 3095
rect 647 3091 651 3095
rect 743 3091 747 3095
rect 855 3091 859 3095
rect 975 3091 979 3095
rect 1103 3091 1107 3095
rect 1239 3091 1243 3095
rect 1383 3091 1387 3095
rect 1527 3091 1531 3095
rect 1895 3095 1899 3099
rect 2087 3095 2091 3099
rect 2303 3095 2307 3099
rect 2511 3095 2515 3099
rect 2703 3095 2707 3099
rect 2879 3095 2883 3099
rect 3047 3095 3051 3099
rect 3199 3095 3203 3099
rect 3351 3095 3355 3099
rect 3487 3095 3491 3099
rect 151 3049 155 3053
rect 239 3049 243 3053
rect 327 3049 331 3053
rect 415 3049 419 3053
rect 503 3049 507 3053
rect 591 3049 595 3053
rect 679 3049 683 3053
rect 767 3049 771 3053
rect 855 3049 859 3053
rect 943 3049 947 3053
rect 1031 3049 1035 3053
rect 1119 3049 1123 3053
rect 1207 3049 1211 3053
rect 1295 3049 1299 3053
rect 1383 3049 1387 3053
rect 1471 3049 1475 3053
rect 1559 3049 1563 3053
rect 1647 3049 1651 3053
rect 1735 3049 1739 3053
rect 2255 3049 2259 3053
rect 2423 3049 2427 3053
rect 2591 3049 2595 3053
rect 2751 3049 2755 3053
rect 2919 3049 2923 3053
rect 3087 3049 3091 3053
rect 111 3036 115 3040
rect 1823 3036 1827 3040
rect 1863 3036 1867 3040
rect 3575 3036 3579 3040
rect 111 3019 115 3023
rect 1823 3019 1827 3023
rect 1863 3019 1867 3023
rect 3575 3019 3579 3023
rect 143 3009 147 3013
rect 231 3009 235 3013
rect 319 3009 323 3013
rect 407 3009 411 3013
rect 495 3009 499 3013
rect 583 3009 587 3013
rect 671 3009 675 3013
rect 759 3009 763 3013
rect 847 3009 851 3013
rect 935 3009 939 3013
rect 1023 3009 1027 3013
rect 1111 3009 1115 3013
rect 1199 3009 1203 3013
rect 1287 3009 1291 3013
rect 1375 3009 1379 3013
rect 1463 3009 1467 3013
rect 1551 3009 1555 3013
rect 1639 3009 1643 3013
rect 1727 3009 1731 3013
rect 2247 3009 2251 3013
rect 2415 3009 2419 3013
rect 2583 3009 2587 3013
rect 2743 3009 2747 3013
rect 2911 3009 2915 3013
rect 3079 3009 3083 3013
rect 1407 2979 1411 2983
rect 1519 2979 1523 2983
rect 1631 2979 1635 2983
rect 1727 2979 1731 2983
rect 2239 2983 2243 2987
rect 2463 2983 2467 2987
rect 2671 2983 2675 2987
rect 2863 2983 2867 2987
rect 3031 2983 3035 2987
rect 3191 2983 3195 2987
rect 3343 2983 3347 2987
rect 3479 2983 3483 2987
rect 111 2969 115 2973
rect 1823 2969 1827 2973
rect 1863 2973 1867 2977
rect 3575 2973 3579 2977
rect 111 2952 115 2956
rect 1823 2952 1827 2956
rect 1863 2956 1867 2960
rect 3575 2956 3579 2960
rect 1415 2939 1419 2943
rect 1527 2939 1531 2943
rect 1639 2939 1643 2943
rect 1735 2939 1739 2943
rect 2247 2943 2251 2947
rect 2471 2943 2475 2947
rect 2679 2943 2683 2947
rect 2871 2943 2875 2947
rect 3039 2943 3043 2947
rect 3199 2943 3203 2947
rect 3351 2943 3355 2947
rect 3487 2943 3491 2947
rect 1359 2905 1363 2909
rect 1471 2905 1475 2909
rect 1583 2905 1587 2909
rect 1703 2905 1707 2909
rect 111 2892 115 2896
rect 1823 2892 1827 2896
rect 2239 2893 2243 2897
rect 2463 2893 2467 2897
rect 2671 2893 2675 2897
rect 2855 2893 2859 2897
rect 3023 2893 3027 2897
rect 3183 2893 3187 2897
rect 3335 2893 3339 2897
rect 3487 2893 3491 2897
rect 1863 2880 1867 2884
rect 111 2875 115 2879
rect 3575 2880 3579 2884
rect 1823 2875 1827 2879
rect 1351 2865 1355 2869
rect 1463 2865 1467 2869
rect 1575 2865 1579 2869
rect 1695 2865 1699 2869
rect 1863 2863 1867 2867
rect 3575 2863 3579 2867
rect 2231 2853 2235 2857
rect 2455 2853 2459 2857
rect 2663 2853 2667 2857
rect 2847 2853 2851 2857
rect 3015 2853 3019 2857
rect 3175 2853 3179 2857
rect 3327 2853 3331 2857
rect 3479 2853 3483 2857
rect 135 2839 139 2843
rect 223 2839 227 2843
rect 311 2839 315 2843
rect 399 2839 403 2843
rect 487 2839 491 2843
rect 599 2839 603 2843
rect 727 2839 731 2843
rect 863 2839 867 2843
rect 999 2839 1003 2843
rect 1135 2839 1139 2843
rect 1263 2839 1267 2843
rect 1383 2839 1387 2843
rect 1503 2839 1507 2843
rect 1623 2839 1627 2843
rect 1727 2839 1731 2843
rect 111 2829 115 2833
rect 1823 2829 1827 2833
rect 1895 2827 1899 2831
rect 1983 2827 1987 2831
rect 2071 2827 2075 2831
rect 2159 2827 2163 2831
rect 2247 2827 2251 2831
rect 2335 2827 2339 2831
rect 2423 2827 2427 2831
rect 2511 2827 2515 2831
rect 2599 2827 2603 2831
rect 2687 2827 2691 2831
rect 2791 2827 2795 2831
rect 2903 2827 2907 2831
rect 3031 2827 3035 2831
rect 3175 2827 3179 2831
rect 3327 2827 3331 2831
rect 3479 2827 3483 2831
rect 1863 2817 1867 2821
rect 111 2812 115 2816
rect 3575 2817 3579 2821
rect 1823 2812 1827 2816
rect 143 2799 147 2803
rect 231 2799 235 2803
rect 319 2799 323 2803
rect 407 2799 411 2803
rect 495 2799 499 2803
rect 607 2799 611 2803
rect 735 2799 739 2803
rect 871 2799 875 2803
rect 1007 2799 1011 2803
rect 1143 2799 1147 2803
rect 1271 2799 1275 2803
rect 1391 2799 1395 2803
rect 1511 2799 1515 2803
rect 1631 2799 1635 2803
rect 1735 2799 1739 2803
rect 1863 2800 1867 2804
rect 3575 2800 3579 2804
rect 1903 2787 1907 2791
rect 1991 2787 1995 2791
rect 2079 2787 2083 2791
rect 2167 2787 2171 2791
rect 2255 2787 2259 2791
rect 2343 2787 2347 2791
rect 2431 2787 2435 2791
rect 2519 2787 2523 2791
rect 2607 2787 2611 2791
rect 2695 2787 2699 2791
rect 2799 2787 2803 2791
rect 2911 2787 2915 2791
rect 3039 2787 3043 2791
rect 3183 2787 3187 2791
rect 3335 2787 3339 2791
rect 3487 2787 3491 2791
rect 191 2765 195 2769
rect 295 2765 299 2769
rect 415 2765 419 2769
rect 551 2765 555 2769
rect 687 2765 691 2769
rect 823 2765 827 2769
rect 959 2765 963 2769
rect 1087 2765 1091 2769
rect 1207 2765 1211 2769
rect 1319 2765 1323 2769
rect 1431 2765 1435 2769
rect 1535 2765 1539 2769
rect 1647 2765 1651 2769
rect 1735 2765 1739 2769
rect 111 2752 115 2756
rect 1823 2752 1827 2756
rect 2047 2741 2051 2745
rect 2167 2741 2171 2745
rect 2295 2741 2299 2745
rect 2447 2741 2451 2745
rect 2623 2741 2627 2745
rect 2823 2741 2827 2745
rect 3039 2741 3043 2745
rect 3271 2741 3275 2745
rect 3487 2741 3491 2745
rect 111 2735 115 2739
rect 1823 2735 1827 2739
rect 183 2725 187 2729
rect 287 2725 291 2729
rect 407 2725 411 2729
rect 543 2725 547 2729
rect 679 2725 683 2729
rect 815 2725 819 2729
rect 951 2725 955 2729
rect 1079 2725 1083 2729
rect 1199 2725 1203 2729
rect 1311 2725 1315 2729
rect 1423 2725 1427 2729
rect 1527 2725 1531 2729
rect 1639 2725 1643 2729
rect 1727 2725 1731 2729
rect 1863 2728 1867 2732
rect 3575 2728 3579 2732
rect 1863 2711 1867 2715
rect 3575 2711 3579 2715
rect 2039 2701 2043 2705
rect 2159 2701 2163 2705
rect 2287 2701 2291 2705
rect 2439 2701 2443 2705
rect 2615 2701 2619 2705
rect 2815 2701 2819 2705
rect 3031 2701 3035 2705
rect 3263 2701 3267 2705
rect 3479 2701 3483 2705
rect 167 2695 171 2699
rect 279 2695 283 2699
rect 391 2695 395 2699
rect 503 2695 507 2699
rect 615 2695 619 2699
rect 111 2685 115 2689
rect 1823 2685 1827 2689
rect 1943 2679 1947 2683
rect 2055 2679 2059 2683
rect 2167 2679 2171 2683
rect 2287 2679 2291 2683
rect 2407 2679 2411 2683
rect 2519 2679 2523 2683
rect 2631 2679 2635 2683
rect 2735 2679 2739 2683
rect 2847 2679 2851 2683
rect 2959 2679 2963 2683
rect 3071 2679 3075 2683
rect 111 2668 115 2672
rect 1823 2668 1827 2672
rect 1863 2669 1867 2673
rect 3575 2669 3579 2673
rect 175 2655 179 2659
rect 287 2655 291 2659
rect 399 2655 403 2659
rect 511 2655 515 2659
rect 623 2655 627 2659
rect 1863 2652 1867 2656
rect 3575 2652 3579 2656
rect 1951 2639 1955 2643
rect 2063 2639 2067 2643
rect 2175 2639 2179 2643
rect 2295 2639 2299 2643
rect 2415 2639 2419 2643
rect 2527 2639 2531 2643
rect 2639 2639 2643 2643
rect 2743 2639 2747 2643
rect 2855 2639 2859 2643
rect 2967 2639 2971 2643
rect 3079 2639 3083 2643
rect 223 2605 227 2609
rect 351 2605 355 2609
rect 495 2605 499 2609
rect 663 2605 667 2609
rect 839 2605 843 2609
rect 1023 2605 1027 2609
rect 1215 2605 1219 2609
rect 1407 2605 1411 2609
rect 1607 2605 1611 2609
rect 1895 2601 1899 2605
rect 2071 2601 2075 2605
rect 2263 2601 2267 2605
rect 2463 2601 2467 2605
rect 2663 2601 2667 2605
rect 2871 2601 2875 2605
rect 3079 2601 3083 2605
rect 3295 2601 3299 2605
rect 3487 2601 3491 2605
rect 111 2592 115 2596
rect 1823 2592 1827 2596
rect 1863 2588 1867 2592
rect 3575 2588 3579 2592
rect 111 2575 115 2579
rect 1823 2575 1827 2579
rect 1863 2571 1867 2575
rect 3575 2571 3579 2575
rect 215 2565 219 2569
rect 343 2565 347 2569
rect 487 2565 491 2569
rect 655 2565 659 2569
rect 831 2565 835 2569
rect 1015 2565 1019 2569
rect 1207 2565 1211 2569
rect 1399 2565 1403 2569
rect 1599 2565 1603 2569
rect 1887 2561 1891 2565
rect 2063 2561 2067 2565
rect 2255 2561 2259 2565
rect 2455 2561 2459 2565
rect 2655 2561 2659 2565
rect 2863 2561 2867 2565
rect 3071 2561 3075 2565
rect 3287 2561 3291 2565
rect 3479 2561 3483 2565
rect 271 2543 275 2547
rect 471 2543 475 2547
rect 671 2543 675 2547
rect 855 2543 859 2547
rect 1023 2543 1027 2547
rect 1175 2543 1179 2547
rect 1319 2543 1323 2547
rect 1455 2543 1459 2547
rect 1591 2543 1595 2547
rect 1727 2543 1731 2547
rect 1887 2539 1891 2543
rect 2039 2539 2043 2543
rect 2215 2539 2219 2543
rect 2399 2539 2403 2543
rect 2575 2539 2579 2543
rect 2743 2539 2747 2543
rect 2903 2539 2907 2543
rect 3055 2539 3059 2543
rect 3199 2539 3203 2543
rect 3343 2539 3347 2543
rect 3479 2539 3483 2543
rect 111 2533 115 2537
rect 1823 2533 1827 2537
rect 1863 2529 1867 2533
rect 3575 2529 3579 2533
rect 111 2516 115 2520
rect 1823 2516 1827 2520
rect 1863 2512 1867 2516
rect 3575 2512 3579 2516
rect 279 2503 283 2507
rect 479 2503 483 2507
rect 679 2503 683 2507
rect 863 2503 867 2507
rect 1031 2503 1035 2507
rect 1183 2503 1187 2507
rect 1327 2503 1331 2507
rect 1463 2503 1467 2507
rect 1599 2503 1603 2507
rect 1735 2503 1739 2507
rect 1895 2499 1899 2503
rect 2047 2499 2051 2503
rect 2223 2499 2227 2503
rect 2407 2499 2411 2503
rect 2583 2499 2587 2503
rect 2751 2499 2755 2503
rect 2911 2499 2915 2503
rect 3063 2499 3067 2503
rect 3207 2499 3211 2503
rect 3351 2499 3355 2503
rect 3487 2499 3491 2503
rect 183 2465 187 2469
rect 319 2465 323 2469
rect 463 2465 467 2469
rect 607 2465 611 2469
rect 743 2465 747 2469
rect 879 2465 883 2469
rect 1007 2465 1011 2469
rect 1127 2465 1131 2469
rect 1239 2465 1243 2469
rect 1343 2465 1347 2469
rect 1447 2465 1451 2469
rect 1551 2465 1555 2469
rect 1647 2465 1651 2469
rect 1735 2465 1739 2469
rect 1895 2465 1899 2469
rect 1991 2465 1995 2469
rect 2127 2465 2131 2469
rect 2279 2465 2283 2469
rect 2439 2465 2443 2469
rect 2599 2465 2603 2469
rect 2767 2465 2771 2469
rect 2943 2465 2947 2469
rect 3119 2465 3123 2469
rect 3295 2465 3299 2469
rect 3471 2465 3475 2469
rect 111 2452 115 2456
rect 1823 2452 1827 2456
rect 1863 2452 1867 2456
rect 3575 2452 3579 2456
rect 111 2435 115 2439
rect 1823 2435 1827 2439
rect 1863 2435 1867 2439
rect 3575 2435 3579 2439
rect 175 2425 179 2429
rect 311 2425 315 2429
rect 455 2425 459 2429
rect 599 2425 603 2429
rect 735 2425 739 2429
rect 871 2425 875 2429
rect 999 2425 1003 2429
rect 1119 2425 1123 2429
rect 1231 2425 1235 2429
rect 1335 2425 1339 2429
rect 1439 2425 1443 2429
rect 1543 2425 1547 2429
rect 1639 2425 1643 2429
rect 1727 2425 1731 2429
rect 1887 2425 1891 2429
rect 1983 2425 1987 2429
rect 2119 2425 2123 2429
rect 2271 2425 2275 2429
rect 2431 2425 2435 2429
rect 2591 2425 2595 2429
rect 2759 2425 2763 2429
rect 2935 2425 2939 2429
rect 3111 2425 3115 2429
rect 3287 2425 3291 2429
rect 3463 2425 3467 2429
rect 151 2395 155 2399
rect 319 2395 323 2399
rect 479 2395 483 2399
rect 639 2395 643 2399
rect 783 2395 787 2399
rect 919 2395 923 2399
rect 1047 2395 1051 2399
rect 1175 2395 1179 2399
rect 1303 2395 1307 2399
rect 1431 2395 1435 2399
rect 2351 2395 2355 2399
rect 2503 2395 2507 2399
rect 2655 2395 2659 2399
rect 2807 2395 2811 2399
rect 2967 2395 2971 2399
rect 3135 2395 3139 2399
rect 3303 2395 3307 2399
rect 3471 2395 3475 2399
rect 111 2385 115 2389
rect 1823 2385 1827 2389
rect 1863 2385 1867 2389
rect 3575 2385 3579 2389
rect 111 2368 115 2372
rect 1823 2368 1827 2372
rect 1863 2368 1867 2372
rect 3575 2368 3579 2372
rect 159 2355 163 2359
rect 327 2355 331 2359
rect 487 2355 491 2359
rect 647 2355 651 2359
rect 791 2355 795 2359
rect 927 2355 931 2359
rect 1055 2355 1059 2359
rect 1183 2355 1187 2359
rect 1311 2355 1315 2359
rect 1439 2355 1443 2359
rect 2359 2355 2363 2359
rect 2511 2355 2515 2359
rect 2663 2355 2667 2359
rect 2815 2355 2819 2359
rect 2975 2355 2979 2359
rect 3143 2355 3147 2359
rect 3311 2355 3315 2359
rect 3479 2355 3483 2359
rect 143 2317 147 2321
rect 263 2317 267 2321
rect 407 2317 411 2321
rect 543 2317 547 2321
rect 679 2317 683 2321
rect 807 2317 811 2321
rect 927 2317 931 2321
rect 1039 2317 1043 2321
rect 1159 2317 1163 2321
rect 1279 2317 1283 2321
rect 2351 2317 2355 2321
rect 2447 2317 2451 2321
rect 2559 2317 2563 2321
rect 2703 2317 2707 2321
rect 2879 2317 2883 2321
rect 3079 2317 3083 2321
rect 3287 2317 3291 2321
rect 3487 2317 3491 2321
rect 111 2304 115 2308
rect 1823 2304 1827 2308
rect 1863 2304 1867 2308
rect 3575 2304 3579 2308
rect 111 2287 115 2291
rect 1823 2287 1827 2291
rect 1863 2287 1867 2291
rect 3575 2287 3579 2291
rect 135 2277 139 2281
rect 255 2277 259 2281
rect 399 2277 403 2281
rect 535 2277 539 2281
rect 671 2277 675 2281
rect 799 2277 803 2281
rect 919 2277 923 2281
rect 1031 2277 1035 2281
rect 1151 2277 1155 2281
rect 1271 2277 1275 2281
rect 2343 2277 2347 2281
rect 2439 2277 2443 2281
rect 2551 2277 2555 2281
rect 2695 2277 2699 2281
rect 2871 2277 2875 2281
rect 3071 2277 3075 2281
rect 3279 2277 3283 2281
rect 3479 2277 3483 2281
rect 135 2255 139 2259
rect 231 2255 235 2259
rect 351 2255 355 2259
rect 471 2255 475 2259
rect 591 2255 595 2259
rect 711 2255 715 2259
rect 823 2255 827 2259
rect 935 2255 939 2259
rect 1055 2255 1059 2259
rect 1175 2255 1179 2259
rect 2335 2255 2339 2259
rect 2447 2255 2451 2259
rect 2583 2255 2587 2259
rect 2735 2255 2739 2259
rect 2911 2255 2915 2259
rect 3103 2255 3107 2259
rect 3303 2255 3307 2259
rect 3479 2255 3483 2259
rect 111 2245 115 2249
rect 1823 2245 1827 2249
rect 1863 2245 1867 2249
rect 3575 2245 3579 2249
rect 111 2228 115 2232
rect 1823 2228 1827 2232
rect 1863 2228 1867 2232
rect 3575 2228 3579 2232
rect 143 2215 147 2219
rect 239 2215 243 2219
rect 359 2215 363 2219
rect 479 2215 483 2219
rect 599 2215 603 2219
rect 719 2215 723 2219
rect 831 2215 835 2219
rect 943 2215 947 2219
rect 1063 2215 1067 2219
rect 1183 2215 1187 2219
rect 2343 2215 2347 2219
rect 2455 2215 2459 2219
rect 2591 2215 2595 2219
rect 2743 2215 2747 2219
rect 2919 2215 2923 2219
rect 3111 2215 3115 2219
rect 3311 2215 3315 2219
rect 3487 2215 3491 2219
rect 143 2177 147 2181
rect 247 2177 251 2181
rect 383 2177 387 2181
rect 519 2177 523 2181
rect 655 2177 659 2181
rect 783 2177 787 2181
rect 911 2177 915 2181
rect 1031 2177 1035 2181
rect 1159 2177 1163 2181
rect 1287 2177 1291 2181
rect 2255 2181 2259 2185
rect 2343 2181 2347 2185
rect 2439 2181 2443 2185
rect 2551 2181 2555 2185
rect 2695 2181 2699 2185
rect 2871 2181 2875 2185
rect 3071 2181 3075 2185
rect 3287 2181 3291 2185
rect 3487 2181 3491 2185
rect 111 2164 115 2168
rect 1823 2164 1827 2168
rect 1863 2168 1867 2172
rect 3575 2168 3579 2172
rect 111 2147 115 2151
rect 1823 2147 1827 2151
rect 1863 2151 1867 2155
rect 3575 2151 3579 2155
rect 135 2137 139 2141
rect 239 2137 243 2141
rect 375 2137 379 2141
rect 511 2137 515 2141
rect 647 2137 651 2141
rect 775 2137 779 2141
rect 903 2137 907 2141
rect 1023 2137 1027 2141
rect 1151 2137 1155 2141
rect 1279 2137 1283 2141
rect 2247 2141 2251 2145
rect 2335 2141 2339 2145
rect 2431 2141 2435 2145
rect 2543 2141 2547 2145
rect 2687 2141 2691 2145
rect 2863 2141 2867 2145
rect 3063 2141 3067 2145
rect 3279 2141 3283 2145
rect 3479 2141 3483 2145
rect 135 2107 139 2111
rect 231 2107 235 2111
rect 359 2107 363 2111
rect 479 2107 483 2111
rect 599 2107 603 2111
rect 719 2107 723 2111
rect 831 2107 835 2111
rect 943 2107 947 2111
rect 1055 2107 1059 2111
rect 1175 2107 1179 2111
rect 2151 2111 2155 2115
rect 2239 2111 2243 2115
rect 2327 2111 2331 2115
rect 2415 2111 2419 2115
rect 2503 2111 2507 2115
rect 2615 2111 2619 2115
rect 2751 2111 2755 2115
rect 2919 2111 2923 2115
rect 3103 2111 3107 2115
rect 3303 2111 3307 2115
rect 3479 2111 3483 2115
rect 111 2097 115 2101
rect 1823 2097 1827 2101
rect 1863 2101 1867 2105
rect 3575 2101 3579 2105
rect 111 2080 115 2084
rect 1823 2080 1827 2084
rect 1863 2084 1867 2088
rect 3575 2084 3579 2088
rect 143 2067 147 2071
rect 239 2067 243 2071
rect 367 2067 371 2071
rect 487 2067 491 2071
rect 607 2067 611 2071
rect 727 2067 731 2071
rect 839 2067 843 2071
rect 951 2067 955 2071
rect 1063 2067 1067 2071
rect 1183 2067 1187 2071
rect 2159 2071 2163 2075
rect 2247 2071 2251 2075
rect 2335 2071 2339 2075
rect 2423 2071 2427 2075
rect 2511 2071 2515 2075
rect 2623 2071 2627 2075
rect 2759 2071 2763 2075
rect 2927 2071 2931 2075
rect 3111 2071 3115 2075
rect 3311 2071 3315 2075
rect 3487 2071 3491 2075
rect 1999 2033 2003 2037
rect 2127 2033 2131 2037
rect 2255 2033 2259 2037
rect 2399 2033 2403 2037
rect 2551 2033 2555 2037
rect 2711 2033 2715 2037
rect 2879 2033 2883 2037
rect 3063 2033 3067 2037
rect 3247 2033 3251 2037
rect 3439 2033 3443 2037
rect 167 2021 171 2025
rect 311 2021 315 2025
rect 447 2021 451 2025
rect 575 2021 579 2025
rect 695 2021 699 2025
rect 807 2021 811 2025
rect 911 2021 915 2025
rect 1015 2021 1019 2025
rect 1119 2021 1123 2025
rect 1223 2021 1227 2025
rect 1327 2021 1331 2025
rect 1863 2020 1867 2024
rect 3575 2020 3579 2024
rect 111 2008 115 2012
rect 1823 2008 1827 2012
rect 1863 2003 1867 2007
rect 3575 2003 3579 2007
rect 111 1991 115 1995
rect 1823 1991 1827 1995
rect 1991 1993 1995 1997
rect 2119 1993 2123 1997
rect 2247 1993 2251 1997
rect 2391 1993 2395 1997
rect 2543 1993 2547 1997
rect 2703 1993 2707 1997
rect 2871 1993 2875 1997
rect 3055 1993 3059 1997
rect 3239 1993 3243 1997
rect 3431 1993 3435 1997
rect 159 1981 163 1985
rect 303 1981 307 1985
rect 439 1981 443 1985
rect 567 1981 571 1985
rect 687 1981 691 1985
rect 799 1981 803 1985
rect 903 1981 907 1985
rect 1007 1981 1011 1985
rect 1111 1981 1115 1985
rect 1215 1981 1219 1985
rect 1319 1981 1323 1985
rect 159 1959 163 1963
rect 295 1959 299 1963
rect 439 1959 443 1963
rect 583 1959 587 1963
rect 719 1959 723 1963
rect 855 1959 859 1963
rect 991 1959 995 1963
rect 1119 1959 1123 1963
rect 1239 1959 1243 1963
rect 1359 1959 1363 1963
rect 1479 1959 1483 1963
rect 1599 1959 1603 1963
rect 1903 1963 1907 1967
rect 2159 1963 2163 1967
rect 2399 1963 2403 1967
rect 2615 1963 2619 1967
rect 2815 1963 2819 1967
rect 2999 1963 3003 1967
rect 3167 1963 3171 1967
rect 3335 1963 3339 1967
rect 3479 1963 3483 1967
rect 111 1949 115 1953
rect 1823 1949 1827 1953
rect 1863 1953 1867 1957
rect 3575 1953 3579 1957
rect 111 1932 115 1936
rect 1823 1932 1827 1936
rect 1863 1936 1867 1940
rect 3575 1936 3579 1940
rect 167 1919 171 1923
rect 303 1919 307 1923
rect 447 1919 451 1923
rect 591 1919 595 1923
rect 727 1919 731 1923
rect 863 1919 867 1923
rect 999 1919 1003 1923
rect 1127 1919 1131 1923
rect 1247 1919 1251 1923
rect 1367 1919 1371 1923
rect 1487 1919 1491 1923
rect 1607 1919 1611 1923
rect 1911 1923 1915 1927
rect 2167 1923 2171 1927
rect 2407 1923 2411 1927
rect 2623 1923 2627 1927
rect 2823 1923 2827 1927
rect 3007 1923 3011 1927
rect 3175 1923 3179 1927
rect 3343 1923 3347 1927
rect 3487 1923 3491 1927
rect 1895 1889 1899 1893
rect 1983 1889 1987 1893
rect 2071 1889 2075 1893
rect 2167 1889 2171 1893
rect 2295 1889 2299 1893
rect 2447 1889 2451 1893
rect 2607 1889 2611 1893
rect 2767 1889 2771 1893
rect 2919 1889 2923 1893
rect 3071 1889 3075 1893
rect 3215 1889 3219 1893
rect 3359 1889 3363 1893
rect 3487 1889 3491 1893
rect 223 1877 227 1881
rect 479 1877 483 1881
rect 719 1877 723 1881
rect 935 1877 939 1881
rect 1127 1877 1131 1881
rect 1295 1877 1299 1881
rect 1455 1877 1459 1881
rect 1607 1877 1611 1881
rect 1735 1877 1739 1881
rect 1863 1876 1867 1880
rect 3575 1876 3579 1880
rect 111 1864 115 1868
rect 1823 1864 1827 1868
rect 1863 1859 1867 1863
rect 3575 1859 3579 1863
rect 111 1847 115 1851
rect 1823 1847 1827 1851
rect 1887 1849 1891 1853
rect 1975 1849 1979 1853
rect 2063 1849 2067 1853
rect 2159 1849 2163 1853
rect 2287 1849 2291 1853
rect 2439 1849 2443 1853
rect 2599 1849 2603 1853
rect 2759 1849 2763 1853
rect 2911 1849 2915 1853
rect 3063 1849 3067 1853
rect 3207 1849 3211 1853
rect 3351 1849 3355 1853
rect 3479 1849 3483 1853
rect 215 1837 219 1841
rect 471 1837 475 1841
rect 711 1837 715 1841
rect 927 1837 931 1841
rect 1119 1837 1123 1841
rect 1287 1837 1291 1841
rect 1447 1837 1451 1841
rect 1599 1837 1603 1841
rect 1727 1837 1731 1841
rect 1999 1823 2003 1827
rect 2223 1823 2227 1827
rect 2439 1823 2443 1827
rect 2639 1823 2643 1827
rect 2831 1823 2835 1827
rect 3015 1823 3019 1827
rect 3199 1823 3203 1827
rect 3391 1823 3395 1827
rect 247 1815 251 1819
rect 415 1815 419 1819
rect 591 1815 595 1819
rect 759 1815 763 1819
rect 927 1815 931 1819
rect 1079 1815 1083 1819
rect 1223 1815 1227 1819
rect 1359 1815 1363 1819
rect 1487 1815 1491 1819
rect 1615 1815 1619 1819
rect 1727 1815 1731 1819
rect 1863 1813 1867 1817
rect 3575 1813 3579 1817
rect 111 1805 115 1809
rect 1823 1805 1827 1809
rect 1863 1796 1867 1800
rect 3575 1796 3579 1800
rect 111 1788 115 1792
rect 1823 1788 1827 1792
rect 2007 1783 2011 1787
rect 2231 1783 2235 1787
rect 2447 1783 2451 1787
rect 2647 1783 2651 1787
rect 2839 1783 2843 1787
rect 3023 1783 3027 1787
rect 3207 1783 3211 1787
rect 3399 1783 3403 1787
rect 255 1775 259 1779
rect 423 1775 427 1779
rect 599 1775 603 1779
rect 767 1775 771 1779
rect 935 1775 939 1779
rect 1087 1775 1091 1779
rect 1231 1775 1235 1779
rect 1367 1775 1371 1779
rect 1495 1775 1499 1779
rect 1623 1775 1627 1779
rect 1735 1775 1739 1779
rect 1943 1745 1947 1749
rect 2087 1745 2091 1749
rect 2247 1745 2251 1749
rect 2415 1745 2419 1749
rect 2599 1745 2603 1749
rect 2791 1745 2795 1749
rect 2991 1745 2995 1749
rect 3199 1745 3203 1749
rect 3415 1745 3419 1749
rect 327 1737 331 1741
rect 471 1737 475 1741
rect 615 1737 619 1741
rect 767 1737 771 1741
rect 919 1737 923 1741
rect 1071 1737 1075 1741
rect 1223 1737 1227 1741
rect 1375 1737 1379 1741
rect 1527 1737 1531 1741
rect 1687 1737 1691 1741
rect 1863 1732 1867 1736
rect 3575 1732 3579 1736
rect 111 1724 115 1728
rect 1823 1724 1827 1728
rect 1863 1715 1867 1719
rect 3575 1715 3579 1719
rect 111 1707 115 1711
rect 1823 1707 1827 1711
rect 1935 1705 1939 1709
rect 2079 1705 2083 1709
rect 2239 1705 2243 1709
rect 2407 1705 2411 1709
rect 2591 1705 2595 1709
rect 2783 1705 2787 1709
rect 2983 1705 2987 1709
rect 3191 1705 3195 1709
rect 3407 1705 3411 1709
rect 319 1697 323 1701
rect 463 1697 467 1701
rect 607 1697 611 1701
rect 759 1697 763 1701
rect 911 1697 915 1701
rect 1063 1697 1067 1701
rect 1215 1697 1219 1701
rect 1367 1697 1371 1701
rect 1519 1697 1523 1701
rect 1679 1697 1683 1701
rect 1911 1679 1915 1683
rect 2031 1679 2035 1683
rect 2151 1679 2155 1683
rect 2271 1679 2275 1683
rect 2399 1679 2403 1683
rect 2543 1679 2547 1683
rect 2695 1679 2699 1683
rect 2863 1679 2867 1683
rect 3047 1679 3051 1683
rect 3239 1679 3243 1683
rect 3431 1679 3435 1683
rect 311 1671 315 1675
rect 447 1671 451 1675
rect 591 1671 595 1675
rect 735 1671 739 1675
rect 887 1671 891 1675
rect 1039 1671 1043 1675
rect 1191 1671 1195 1675
rect 1343 1671 1347 1675
rect 1495 1671 1499 1675
rect 1647 1671 1651 1675
rect 1863 1669 1867 1673
rect 3575 1669 3579 1673
rect 111 1661 115 1665
rect 1823 1661 1827 1665
rect 1863 1652 1867 1656
rect 3575 1652 3579 1656
rect 111 1644 115 1648
rect 1823 1644 1827 1648
rect 1919 1639 1923 1643
rect 2039 1639 2043 1643
rect 2159 1639 2163 1643
rect 2279 1639 2283 1643
rect 2407 1639 2411 1643
rect 2551 1639 2555 1643
rect 2703 1639 2707 1643
rect 2871 1639 2875 1643
rect 3055 1639 3059 1643
rect 3247 1639 3251 1643
rect 3439 1639 3443 1643
rect 319 1631 323 1635
rect 455 1631 459 1635
rect 599 1631 603 1635
rect 743 1631 747 1635
rect 895 1631 899 1635
rect 1047 1631 1051 1635
rect 1199 1631 1203 1635
rect 1351 1631 1355 1635
rect 1503 1631 1507 1635
rect 1655 1631 1659 1635
rect 1895 1597 1899 1601
rect 2015 1597 2019 1601
rect 2151 1597 2155 1601
rect 2287 1597 2291 1601
rect 2431 1597 2435 1601
rect 2583 1597 2587 1601
rect 2743 1597 2747 1601
rect 2911 1597 2915 1601
rect 3095 1597 3099 1601
rect 3279 1597 3283 1601
rect 3471 1597 3475 1601
rect 223 1589 227 1593
rect 351 1589 355 1593
rect 487 1589 491 1593
rect 623 1589 627 1593
rect 759 1589 763 1593
rect 903 1589 907 1593
rect 1055 1589 1059 1593
rect 1215 1589 1219 1593
rect 1375 1589 1379 1593
rect 1543 1589 1547 1593
rect 1863 1584 1867 1588
rect 3575 1584 3579 1588
rect 111 1576 115 1580
rect 1823 1576 1827 1580
rect 1863 1567 1867 1571
rect 3575 1567 3579 1571
rect 111 1559 115 1563
rect 1823 1559 1827 1563
rect 1887 1557 1891 1561
rect 2007 1557 2011 1561
rect 2143 1557 2147 1561
rect 2279 1557 2283 1561
rect 2423 1557 2427 1561
rect 2575 1557 2579 1561
rect 2735 1557 2739 1561
rect 2903 1557 2907 1561
rect 3087 1557 3091 1561
rect 3271 1557 3275 1561
rect 3463 1557 3467 1561
rect 215 1549 219 1553
rect 343 1549 347 1553
rect 479 1549 483 1553
rect 615 1549 619 1553
rect 751 1549 755 1553
rect 895 1549 899 1553
rect 1047 1549 1051 1553
rect 1207 1549 1211 1553
rect 1367 1549 1371 1553
rect 1535 1549 1539 1553
rect 135 1523 139 1527
rect 271 1523 275 1527
rect 423 1523 427 1527
rect 583 1523 587 1527
rect 735 1523 739 1527
rect 887 1523 891 1527
rect 1039 1523 1043 1527
rect 1191 1523 1195 1527
rect 1343 1523 1347 1527
rect 1495 1523 1499 1527
rect 1887 1527 1891 1531
rect 2023 1527 2027 1531
rect 2183 1527 2187 1531
rect 2343 1527 2347 1531
rect 2503 1527 2507 1531
rect 2663 1527 2667 1531
rect 2823 1527 2827 1531
rect 2983 1527 2987 1531
rect 3151 1527 3155 1531
rect 3319 1527 3323 1531
rect 3479 1527 3483 1531
rect 111 1513 115 1517
rect 1823 1513 1827 1517
rect 1863 1517 1867 1521
rect 3575 1517 3579 1521
rect 111 1496 115 1500
rect 1823 1496 1827 1500
rect 1863 1500 1867 1504
rect 3575 1500 3579 1504
rect 143 1483 147 1487
rect 279 1483 283 1487
rect 431 1483 435 1487
rect 591 1483 595 1487
rect 743 1483 747 1487
rect 895 1483 899 1487
rect 1047 1483 1051 1487
rect 1199 1483 1203 1487
rect 1351 1483 1355 1487
rect 1503 1483 1507 1487
rect 1895 1487 1899 1491
rect 2031 1487 2035 1491
rect 2191 1487 2195 1491
rect 2351 1487 2355 1491
rect 2511 1487 2515 1491
rect 2671 1487 2675 1491
rect 2831 1487 2835 1491
rect 2991 1487 2995 1491
rect 3159 1487 3163 1491
rect 3327 1487 3331 1491
rect 3487 1487 3491 1491
rect 143 1441 147 1445
rect 263 1441 267 1445
rect 399 1441 403 1445
rect 535 1441 539 1445
rect 663 1441 667 1445
rect 791 1441 795 1445
rect 911 1441 915 1445
rect 1023 1441 1027 1445
rect 1143 1441 1147 1445
rect 1263 1441 1267 1445
rect 1383 1441 1387 1445
rect 1503 1441 1507 1445
rect 1631 1441 1635 1445
rect 1735 1441 1739 1445
rect 2183 1445 2187 1449
rect 2359 1445 2363 1449
rect 2527 1445 2531 1449
rect 2687 1445 2691 1449
rect 2847 1445 2851 1449
rect 3007 1445 3011 1449
rect 3175 1445 3179 1449
rect 3343 1445 3347 1449
rect 3487 1445 3491 1449
rect 111 1428 115 1432
rect 1823 1428 1827 1432
rect 1863 1432 1867 1436
rect 3575 1432 3579 1436
rect 111 1411 115 1415
rect 1823 1411 1827 1415
rect 1863 1415 1867 1419
rect 3575 1415 3579 1419
rect 135 1401 139 1405
rect 255 1401 259 1405
rect 391 1401 395 1405
rect 527 1401 531 1405
rect 655 1401 659 1405
rect 783 1401 787 1405
rect 903 1401 907 1405
rect 1015 1401 1019 1405
rect 1135 1401 1139 1405
rect 1255 1401 1259 1405
rect 1375 1401 1379 1405
rect 1495 1401 1499 1405
rect 1623 1401 1627 1405
rect 1727 1401 1731 1405
rect 2175 1405 2179 1409
rect 2351 1405 2355 1409
rect 2519 1405 2523 1409
rect 2679 1405 2683 1409
rect 2839 1405 2843 1409
rect 2999 1405 3003 1409
rect 3167 1405 3171 1409
rect 3335 1405 3339 1409
rect 3479 1405 3483 1409
rect 135 1379 139 1383
rect 327 1379 331 1383
rect 551 1379 555 1383
rect 783 1379 787 1383
rect 1023 1379 1027 1383
rect 1263 1379 1267 1383
rect 1503 1379 1507 1383
rect 1727 1379 1731 1383
rect 2079 1375 2083 1379
rect 2263 1375 2267 1379
rect 2439 1375 2443 1379
rect 2615 1375 2619 1379
rect 2783 1375 2787 1379
rect 2935 1375 2939 1379
rect 3079 1375 3083 1379
rect 3223 1375 3227 1379
rect 3359 1375 3363 1379
rect 3479 1375 3483 1379
rect 111 1369 115 1373
rect 1823 1369 1827 1373
rect 1863 1365 1867 1369
rect 3575 1365 3579 1369
rect 111 1352 115 1356
rect 1823 1352 1827 1356
rect 1863 1348 1867 1352
rect 3575 1348 3579 1352
rect 143 1339 147 1343
rect 335 1339 339 1343
rect 559 1339 563 1343
rect 791 1339 795 1343
rect 1031 1339 1035 1343
rect 1271 1339 1275 1343
rect 1511 1339 1515 1343
rect 1735 1339 1739 1343
rect 2087 1335 2091 1339
rect 2271 1335 2275 1339
rect 2447 1335 2451 1339
rect 2623 1335 2627 1339
rect 2791 1335 2795 1339
rect 2943 1335 2947 1339
rect 3087 1335 3091 1339
rect 3231 1335 3235 1339
rect 3367 1335 3371 1339
rect 3487 1335 3491 1339
rect 143 1297 147 1301
rect 327 1297 331 1301
rect 527 1297 531 1301
rect 719 1297 723 1301
rect 903 1297 907 1301
rect 1071 1297 1075 1301
rect 1231 1297 1235 1301
rect 1383 1297 1387 1301
rect 1535 1297 1539 1301
rect 1687 1297 1691 1301
rect 2087 1301 2091 1305
rect 2311 1301 2315 1305
rect 2519 1301 2523 1305
rect 2711 1301 2715 1305
rect 2887 1301 2891 1305
rect 3047 1301 3051 1305
rect 3199 1301 3203 1305
rect 3351 1301 3355 1305
rect 3487 1301 3491 1305
rect 111 1284 115 1288
rect 1823 1284 1827 1288
rect 1863 1288 1867 1292
rect 3575 1288 3579 1292
rect 111 1267 115 1271
rect 1823 1267 1827 1271
rect 1863 1271 1867 1275
rect 3575 1271 3579 1275
rect 135 1257 139 1261
rect 319 1257 323 1261
rect 519 1257 523 1261
rect 711 1257 715 1261
rect 895 1257 899 1261
rect 1063 1257 1067 1261
rect 1223 1257 1227 1261
rect 1375 1257 1379 1261
rect 1527 1257 1531 1261
rect 1679 1257 1683 1261
rect 2079 1261 2083 1265
rect 2303 1261 2307 1265
rect 2511 1261 2515 1265
rect 2703 1261 2707 1265
rect 2879 1261 2883 1265
rect 3039 1261 3043 1265
rect 3191 1261 3195 1265
rect 3343 1261 3347 1265
rect 3479 1261 3483 1265
rect 135 1231 139 1235
rect 295 1231 299 1235
rect 479 1231 483 1235
rect 655 1231 659 1235
rect 815 1231 819 1235
rect 967 1231 971 1235
rect 1111 1231 1115 1235
rect 1247 1231 1251 1235
rect 1383 1231 1387 1235
rect 1527 1231 1531 1235
rect 1903 1235 1907 1239
rect 1991 1235 1995 1239
rect 2095 1235 2099 1239
rect 2215 1235 2219 1239
rect 2351 1235 2355 1239
rect 2487 1235 2491 1239
rect 2631 1235 2635 1239
rect 2775 1235 2779 1239
rect 2919 1235 2923 1239
rect 3063 1235 3067 1239
rect 3207 1235 3211 1239
rect 3351 1235 3355 1239
rect 3479 1235 3483 1239
rect 111 1221 115 1225
rect 1823 1221 1827 1225
rect 1863 1225 1867 1229
rect 3575 1225 3579 1229
rect 111 1204 115 1208
rect 1823 1204 1827 1208
rect 1863 1208 1867 1212
rect 3575 1208 3579 1212
rect 143 1191 147 1195
rect 303 1191 307 1195
rect 487 1191 491 1195
rect 663 1191 667 1195
rect 823 1191 827 1195
rect 975 1191 979 1195
rect 1119 1191 1123 1195
rect 1255 1191 1259 1195
rect 1391 1191 1395 1195
rect 1535 1191 1539 1195
rect 1911 1195 1915 1199
rect 1999 1195 2003 1199
rect 2103 1195 2107 1199
rect 2223 1195 2227 1199
rect 2359 1195 2363 1199
rect 2495 1195 2499 1199
rect 2639 1195 2643 1199
rect 2783 1195 2787 1199
rect 2927 1195 2931 1199
rect 3071 1195 3075 1199
rect 3215 1195 3219 1199
rect 3359 1195 3363 1199
rect 3487 1195 3491 1199
rect 167 1153 171 1157
rect 319 1153 323 1157
rect 471 1153 475 1157
rect 615 1153 619 1157
rect 759 1153 763 1157
rect 911 1153 915 1157
rect 1063 1153 1067 1157
rect 1231 1153 1235 1157
rect 1399 1153 1403 1157
rect 1575 1153 1579 1157
rect 1735 1153 1739 1157
rect 1895 1157 1899 1161
rect 2063 1157 2067 1161
rect 2255 1157 2259 1161
rect 2439 1157 2443 1161
rect 2615 1157 2619 1161
rect 2791 1157 2795 1161
rect 2967 1157 2971 1161
rect 3143 1157 3147 1161
rect 3327 1157 3331 1161
rect 3487 1157 3491 1161
rect 111 1140 115 1144
rect 1823 1140 1827 1144
rect 1863 1144 1867 1148
rect 3575 1144 3579 1148
rect 111 1123 115 1127
rect 1823 1123 1827 1127
rect 1863 1127 1867 1131
rect 3575 1127 3579 1131
rect 159 1113 163 1117
rect 311 1113 315 1117
rect 463 1113 467 1117
rect 607 1113 611 1117
rect 751 1113 755 1117
rect 903 1113 907 1117
rect 1055 1113 1059 1117
rect 1223 1113 1227 1117
rect 1391 1113 1395 1117
rect 1567 1113 1571 1117
rect 1727 1113 1731 1117
rect 1887 1117 1891 1121
rect 2055 1117 2059 1121
rect 2247 1117 2251 1121
rect 2431 1117 2435 1121
rect 2607 1117 2611 1121
rect 2783 1117 2787 1121
rect 2959 1117 2963 1121
rect 3135 1117 3139 1121
rect 3319 1117 3323 1121
rect 3479 1117 3483 1121
rect 215 1087 219 1091
rect 327 1087 331 1091
rect 439 1087 443 1091
rect 559 1087 563 1091
rect 679 1087 683 1091
rect 807 1087 811 1091
rect 943 1087 947 1091
rect 1087 1087 1091 1091
rect 1247 1087 1251 1091
rect 1407 1087 1411 1091
rect 1575 1087 1579 1091
rect 1727 1087 1731 1091
rect 1935 1083 1939 1087
rect 2095 1083 2099 1087
rect 2247 1083 2251 1087
rect 2407 1083 2411 1087
rect 2567 1083 2571 1087
rect 2735 1083 2739 1087
rect 2911 1083 2915 1087
rect 3095 1083 3099 1087
rect 3287 1083 3291 1087
rect 3479 1083 3483 1087
rect 111 1077 115 1081
rect 1823 1077 1827 1081
rect 1863 1073 1867 1077
rect 3575 1073 3579 1077
rect 111 1060 115 1064
rect 1823 1060 1827 1064
rect 1863 1056 1867 1060
rect 3575 1056 3579 1060
rect 223 1047 227 1051
rect 335 1047 339 1051
rect 447 1047 451 1051
rect 567 1047 571 1051
rect 687 1047 691 1051
rect 815 1047 819 1051
rect 951 1047 955 1051
rect 1095 1047 1099 1051
rect 1255 1047 1259 1051
rect 1415 1047 1419 1051
rect 1583 1047 1587 1051
rect 1735 1047 1739 1051
rect 1943 1043 1947 1047
rect 2103 1043 2107 1047
rect 2255 1043 2259 1047
rect 2415 1043 2419 1047
rect 2575 1043 2579 1047
rect 2743 1043 2747 1047
rect 2919 1043 2923 1047
rect 3103 1043 3107 1047
rect 3295 1043 3299 1047
rect 3487 1043 3491 1047
rect 343 1005 347 1009
rect 431 1005 435 1009
rect 535 1005 539 1009
rect 655 1005 659 1009
rect 791 1005 795 1009
rect 951 1005 955 1009
rect 1135 1005 1139 1009
rect 1327 1005 1331 1009
rect 1535 1005 1539 1009
rect 1735 1005 1739 1009
rect 1943 1005 1947 1009
rect 2071 1005 2075 1009
rect 2191 1005 2195 1009
rect 2311 1005 2315 1009
rect 2439 1005 2443 1009
rect 2575 1005 2579 1009
rect 2719 1005 2723 1009
rect 2871 1005 2875 1009
rect 3031 1005 3035 1009
rect 3191 1005 3195 1009
rect 3351 1005 3355 1009
rect 3487 1005 3491 1009
rect 111 992 115 996
rect 1823 992 1827 996
rect 1863 992 1867 996
rect 3575 992 3579 996
rect 111 975 115 979
rect 1823 975 1827 979
rect 1863 975 1867 979
rect 3575 975 3579 979
rect 335 965 339 969
rect 423 965 427 969
rect 527 965 531 969
rect 647 965 651 969
rect 783 965 787 969
rect 943 965 947 969
rect 1127 965 1131 969
rect 1319 965 1323 969
rect 1527 965 1531 969
rect 1727 965 1731 969
rect 1935 965 1939 969
rect 2063 965 2067 969
rect 2183 965 2187 969
rect 2303 965 2307 969
rect 2431 965 2435 969
rect 2567 965 2571 969
rect 2711 965 2715 969
rect 2863 965 2867 969
rect 3023 965 3027 969
rect 3183 965 3187 969
rect 3343 965 3347 969
rect 3479 965 3483 969
rect 367 939 371 943
rect 463 939 467 943
rect 575 939 579 943
rect 703 939 707 943
rect 847 939 851 943
rect 1007 939 1011 943
rect 1175 939 1179 943
rect 1351 939 1355 943
rect 1527 939 1531 943
rect 1711 939 1715 943
rect 1887 939 1891 943
rect 2047 939 2051 943
rect 2199 939 2203 943
rect 2351 939 2355 943
rect 2495 939 2499 943
rect 2631 939 2635 943
rect 2759 939 2763 943
rect 2887 939 2891 943
rect 3023 939 3027 943
rect 111 929 115 933
rect 1823 929 1827 933
rect 1863 929 1867 933
rect 3575 929 3579 933
rect 111 912 115 916
rect 1823 912 1827 916
rect 1863 912 1867 916
rect 3575 912 3579 916
rect 375 899 379 903
rect 471 899 475 903
rect 583 899 587 903
rect 711 899 715 903
rect 855 899 859 903
rect 1015 899 1019 903
rect 1183 899 1187 903
rect 1359 899 1363 903
rect 1535 899 1539 903
rect 1719 899 1723 903
rect 1895 899 1899 903
rect 2055 899 2059 903
rect 2207 899 2211 903
rect 2359 899 2363 903
rect 2503 899 2507 903
rect 2639 899 2643 903
rect 2767 899 2771 903
rect 2895 899 2899 903
rect 3031 899 3035 903
rect 343 861 347 865
rect 431 861 435 865
rect 535 861 539 865
rect 647 861 651 865
rect 783 861 787 865
rect 927 861 931 865
rect 1087 861 1091 865
rect 1263 861 1267 865
rect 1447 861 1451 865
rect 1631 861 1635 865
rect 1895 865 1899 869
rect 2015 865 2019 869
rect 2167 865 2171 869
rect 2319 865 2323 869
rect 2487 865 2491 869
rect 2663 865 2667 869
rect 2847 865 2851 869
rect 3039 865 3043 869
rect 3239 865 3243 869
rect 3439 865 3443 869
rect 111 848 115 852
rect 1823 848 1827 852
rect 1863 852 1867 856
rect 3575 852 3579 856
rect 111 831 115 835
rect 1823 831 1827 835
rect 1863 835 1867 839
rect 3575 835 3579 839
rect 335 821 339 825
rect 423 821 427 825
rect 527 821 531 825
rect 639 821 643 825
rect 775 821 779 825
rect 919 821 923 825
rect 1079 821 1083 825
rect 1255 821 1259 825
rect 1439 821 1443 825
rect 1623 821 1627 825
rect 1887 825 1891 829
rect 2007 825 2011 829
rect 2159 825 2163 829
rect 2311 825 2315 829
rect 2479 825 2483 829
rect 2655 825 2659 829
rect 2839 825 2843 829
rect 3031 825 3035 829
rect 3231 825 3235 829
rect 3431 825 3435 829
rect 287 799 291 803
rect 407 799 411 803
rect 535 799 539 803
rect 679 799 683 803
rect 823 799 827 803
rect 975 799 979 803
rect 1127 799 1131 803
rect 1279 799 1283 803
rect 1439 799 1443 803
rect 1599 799 1603 803
rect 1887 803 1891 807
rect 1991 803 1995 807
rect 2135 803 2139 807
rect 2287 803 2291 807
rect 2455 803 2459 807
rect 2623 803 2627 807
rect 2799 803 2803 807
rect 2967 803 2971 807
rect 3143 803 3147 807
rect 3319 803 3323 807
rect 3479 803 3483 807
rect 111 789 115 793
rect 1823 789 1827 793
rect 1863 793 1867 797
rect 3575 793 3579 797
rect 111 772 115 776
rect 1823 772 1827 776
rect 1863 776 1867 780
rect 3575 776 3579 780
rect 295 759 299 763
rect 415 759 419 763
rect 543 759 547 763
rect 687 759 691 763
rect 831 759 835 763
rect 983 759 987 763
rect 1135 759 1139 763
rect 1287 759 1291 763
rect 1447 759 1451 763
rect 1607 759 1611 763
rect 1895 763 1899 767
rect 1999 763 2003 767
rect 2143 763 2147 767
rect 2295 763 2299 767
rect 2463 763 2467 767
rect 2631 763 2635 767
rect 2807 763 2811 767
rect 2975 763 2979 767
rect 3151 763 3155 767
rect 3327 763 3331 767
rect 3487 763 3491 767
rect 215 721 219 725
rect 359 721 363 725
rect 503 721 507 725
rect 647 721 651 725
rect 791 721 795 725
rect 935 721 939 725
rect 1087 721 1091 725
rect 1247 721 1251 725
rect 1415 721 1419 725
rect 1583 721 1587 725
rect 1735 721 1739 725
rect 1895 725 1899 729
rect 2063 725 2067 729
rect 2255 725 2259 729
rect 2447 725 2451 729
rect 2639 725 2643 729
rect 2823 725 2827 729
rect 2999 725 3003 729
rect 3167 725 3171 729
rect 3335 725 3339 729
rect 3487 725 3491 729
rect 111 708 115 712
rect 1823 708 1827 712
rect 1863 712 1867 716
rect 3575 712 3579 716
rect 111 691 115 695
rect 1823 691 1827 695
rect 1863 695 1867 699
rect 3575 695 3579 699
rect 207 681 211 685
rect 351 681 355 685
rect 495 681 499 685
rect 639 681 643 685
rect 783 681 787 685
rect 927 681 931 685
rect 1079 681 1083 685
rect 1239 681 1243 685
rect 1407 681 1411 685
rect 1575 681 1579 685
rect 1727 681 1731 685
rect 1887 685 1891 689
rect 2055 685 2059 689
rect 2247 685 2251 689
rect 2439 685 2443 689
rect 2631 685 2635 689
rect 2815 685 2819 689
rect 2991 685 2995 689
rect 3159 685 3163 689
rect 3327 685 3331 689
rect 3479 685 3483 689
rect 135 659 139 663
rect 295 659 299 663
rect 463 659 467 663
rect 623 659 627 663
rect 775 659 779 663
rect 927 659 931 663
rect 1071 659 1075 663
rect 1207 659 1211 663
rect 1343 659 1347 663
rect 1479 659 1483 663
rect 1615 659 1619 663
rect 1727 659 1731 663
rect 2215 659 2219 663
rect 2359 659 2363 663
rect 2511 659 2515 663
rect 2671 659 2675 663
rect 2831 659 2835 663
rect 2991 659 2995 663
rect 3159 659 3163 663
rect 3327 659 3331 663
rect 3479 659 3483 663
rect 111 649 115 653
rect 1823 649 1827 653
rect 1863 649 1867 653
rect 3575 649 3579 653
rect 111 632 115 636
rect 1823 632 1827 636
rect 1863 632 1867 636
rect 3575 632 3579 636
rect 143 619 147 623
rect 303 619 307 623
rect 471 619 475 623
rect 631 619 635 623
rect 783 619 787 623
rect 935 619 939 623
rect 1079 619 1083 623
rect 1215 619 1219 623
rect 1351 619 1355 623
rect 1487 619 1491 623
rect 1623 619 1627 623
rect 1735 619 1739 623
rect 2223 619 2227 623
rect 2367 619 2371 623
rect 2519 619 2523 623
rect 2679 619 2683 623
rect 2839 619 2843 623
rect 2999 619 3003 623
rect 3167 619 3171 623
rect 3335 619 3339 623
rect 3487 619 3491 623
rect 143 581 147 585
rect 303 581 307 585
rect 487 581 491 585
rect 671 581 675 585
rect 847 581 851 585
rect 1023 581 1027 585
rect 1199 581 1203 585
rect 1375 581 1379 585
rect 1559 581 1563 585
rect 1735 581 1739 585
rect 2199 581 2203 585
rect 2287 581 2291 585
rect 2375 581 2379 585
rect 2463 581 2467 585
rect 2567 581 2571 585
rect 2679 581 2683 585
rect 2815 581 2819 585
rect 2975 581 2979 585
rect 3143 581 3147 585
rect 3327 581 3331 585
rect 3487 581 3491 585
rect 111 568 115 572
rect 1823 568 1827 572
rect 1863 568 1867 572
rect 3575 568 3579 572
rect 111 551 115 555
rect 1823 551 1827 555
rect 1863 551 1867 555
rect 3575 551 3579 555
rect 135 541 139 545
rect 295 541 299 545
rect 479 541 483 545
rect 663 541 667 545
rect 839 541 843 545
rect 1015 541 1019 545
rect 1191 541 1195 545
rect 1367 541 1371 545
rect 1551 541 1555 545
rect 1727 541 1731 545
rect 2191 541 2195 545
rect 2279 541 2283 545
rect 2367 541 2371 545
rect 2455 541 2459 545
rect 2559 541 2563 545
rect 2671 541 2675 545
rect 2807 541 2811 545
rect 2967 541 2971 545
rect 3135 541 3139 545
rect 3319 541 3323 545
rect 3479 541 3483 545
rect 135 515 139 519
rect 303 515 307 519
rect 495 515 499 519
rect 679 515 683 519
rect 863 515 867 519
rect 1031 515 1035 519
rect 1191 515 1195 519
rect 1351 515 1355 519
rect 1503 515 1507 519
rect 1663 515 1667 519
rect 2303 515 2307 519
rect 2399 515 2403 519
rect 2503 515 2507 519
rect 2607 515 2611 519
rect 2719 515 2723 519
rect 2839 515 2843 519
rect 2967 515 2971 519
rect 3095 515 3099 519
rect 3223 515 3227 519
rect 3351 515 3355 519
rect 3479 515 3483 519
rect 111 505 115 509
rect 1823 505 1827 509
rect 1863 505 1867 509
rect 3575 505 3579 509
rect 111 488 115 492
rect 1823 488 1827 492
rect 1863 488 1867 492
rect 3575 488 3579 492
rect 143 475 147 479
rect 311 475 315 479
rect 503 475 507 479
rect 687 475 691 479
rect 871 475 875 479
rect 1039 475 1043 479
rect 1199 475 1203 479
rect 1359 475 1363 479
rect 1511 475 1515 479
rect 1671 475 1675 479
rect 2311 475 2315 479
rect 2407 475 2411 479
rect 2511 475 2515 479
rect 2615 475 2619 479
rect 2727 475 2731 479
rect 2847 475 2851 479
rect 2975 475 2979 479
rect 3103 475 3107 479
rect 3231 475 3235 479
rect 3359 475 3363 479
rect 3487 475 3491 479
rect 143 437 147 441
rect 303 437 307 441
rect 495 437 499 441
rect 687 437 691 441
rect 879 437 883 441
rect 1055 437 1059 441
rect 1223 437 1227 441
rect 1391 437 1395 441
rect 1559 437 1563 441
rect 1727 437 1731 441
rect 2239 441 2243 445
rect 2327 441 2331 445
rect 2431 441 2435 445
rect 2559 441 2563 445
rect 2695 441 2699 445
rect 2847 441 2851 445
rect 2999 441 3003 445
rect 3159 441 3163 445
rect 3327 441 3331 445
rect 3487 441 3491 445
rect 111 424 115 428
rect 1823 424 1827 428
rect 1863 428 1867 432
rect 3575 428 3579 432
rect 111 407 115 411
rect 1823 407 1827 411
rect 1863 411 1867 415
rect 3575 411 3579 415
rect 135 397 139 401
rect 295 397 299 401
rect 487 397 491 401
rect 679 397 683 401
rect 871 397 875 401
rect 1047 397 1051 401
rect 1215 397 1219 401
rect 1383 397 1387 401
rect 1551 397 1555 401
rect 1719 397 1723 401
rect 2231 401 2235 405
rect 2319 401 2323 405
rect 2423 401 2427 405
rect 2551 401 2555 405
rect 2687 401 2691 405
rect 2839 401 2843 405
rect 2991 401 2995 405
rect 3151 401 3155 405
rect 3319 401 3323 405
rect 3479 401 3483 405
rect 135 375 139 379
rect 263 375 267 379
rect 423 375 427 379
rect 591 375 595 379
rect 767 375 771 379
rect 935 375 939 379
rect 1103 375 1107 379
rect 1263 375 1267 379
rect 1423 375 1427 379
rect 1583 375 1587 379
rect 1727 375 1731 379
rect 2183 379 2187 383
rect 2287 379 2291 383
rect 2399 379 2403 383
rect 2527 379 2531 383
rect 2671 379 2675 383
rect 2815 379 2819 383
rect 2967 379 2971 383
rect 3127 379 3131 383
rect 3295 379 3299 383
rect 3463 379 3467 383
rect 111 365 115 369
rect 1823 365 1827 369
rect 1863 369 1867 373
rect 3575 369 3579 373
rect 111 348 115 352
rect 1823 348 1827 352
rect 1863 352 1867 356
rect 3575 352 3579 356
rect 143 335 147 339
rect 271 335 275 339
rect 431 335 435 339
rect 599 335 603 339
rect 775 335 779 339
rect 943 335 947 339
rect 1111 335 1115 339
rect 1271 335 1275 339
rect 1431 335 1435 339
rect 1591 335 1595 339
rect 1735 335 1739 339
rect 2191 339 2195 343
rect 2295 339 2299 343
rect 2407 339 2411 343
rect 2535 339 2539 343
rect 2679 339 2683 343
rect 2823 339 2827 343
rect 2975 339 2979 343
rect 3135 339 3139 343
rect 3303 339 3307 343
rect 3471 339 3475 343
rect 215 301 219 305
rect 351 301 355 305
rect 495 301 499 305
rect 639 301 643 305
rect 791 301 795 305
rect 935 301 939 305
rect 1079 301 1083 305
rect 1223 301 1227 305
rect 1359 301 1363 305
rect 1487 301 1491 305
rect 1623 301 1627 305
rect 1735 301 1739 305
rect 1895 297 1899 301
rect 2087 297 2091 301
rect 2303 297 2307 301
rect 2511 297 2515 301
rect 2711 297 2715 301
rect 2903 297 2907 301
rect 3095 297 3099 301
rect 3295 297 3299 301
rect 3487 297 3491 301
rect 111 288 115 292
rect 1823 288 1827 292
rect 1863 284 1867 288
rect 3575 284 3579 288
rect 111 271 115 275
rect 1823 271 1827 275
rect 1863 267 1867 271
rect 3575 267 3579 271
rect 207 261 211 265
rect 343 261 347 265
rect 487 261 491 265
rect 631 261 635 265
rect 783 261 787 265
rect 927 261 931 265
rect 1071 261 1075 265
rect 1215 261 1219 265
rect 1351 261 1355 265
rect 1479 261 1483 265
rect 1615 261 1619 265
rect 1727 261 1731 265
rect 1887 257 1891 261
rect 2079 257 2083 261
rect 2295 257 2299 261
rect 2503 257 2507 261
rect 2703 257 2707 261
rect 2895 257 2899 261
rect 3087 257 3091 261
rect 3287 257 3291 261
rect 3479 257 3483 261
rect 231 231 235 235
rect 359 231 363 235
rect 487 231 491 235
rect 623 231 627 235
rect 759 231 763 235
rect 895 231 899 235
rect 1031 231 1035 235
rect 1159 231 1163 235
rect 1295 231 1299 235
rect 1431 231 1435 235
rect 1887 235 1891 239
rect 1999 235 2003 239
rect 2143 235 2147 239
rect 2295 235 2299 239
rect 2455 235 2459 239
rect 2615 235 2619 239
rect 2783 235 2787 239
rect 2951 235 2955 239
rect 3127 235 3131 239
rect 3311 235 3315 239
rect 3479 235 3483 239
rect 111 221 115 225
rect 1823 221 1827 225
rect 1863 225 1867 229
rect 3575 225 3579 229
rect 111 204 115 208
rect 1823 204 1827 208
rect 1863 208 1867 212
rect 3575 208 3579 212
rect 239 191 243 195
rect 367 191 371 195
rect 495 191 499 195
rect 631 191 635 195
rect 767 191 771 195
rect 903 191 907 195
rect 1039 191 1043 195
rect 1167 191 1171 195
rect 1303 191 1307 195
rect 1439 191 1443 195
rect 1895 195 1899 199
rect 2007 195 2011 199
rect 2151 195 2155 199
rect 2303 195 2307 199
rect 2463 195 2467 199
rect 2623 195 2627 199
rect 2791 195 2795 199
rect 2959 195 2963 199
rect 3135 195 3139 199
rect 3319 195 3323 199
rect 3487 195 3491 199
rect 175 133 179 137
rect 263 133 267 137
rect 351 133 355 137
rect 439 133 443 137
rect 527 133 531 137
rect 615 133 619 137
rect 703 133 707 137
rect 791 133 795 137
rect 879 133 883 137
rect 967 133 971 137
rect 1055 133 1059 137
rect 1143 133 1147 137
rect 1231 133 1235 137
rect 1319 133 1323 137
rect 1407 133 1411 137
rect 1503 133 1507 137
rect 1895 133 1899 137
rect 1983 133 1987 137
rect 2071 133 2075 137
rect 2159 133 2163 137
rect 2247 133 2251 137
rect 2335 133 2339 137
rect 2439 133 2443 137
rect 2543 133 2547 137
rect 2647 133 2651 137
rect 2743 133 2747 137
rect 2839 133 2843 137
rect 2935 133 2939 137
rect 3031 133 3035 137
rect 3127 133 3131 137
rect 3223 133 3227 137
rect 3311 133 3315 137
rect 3399 133 3403 137
rect 3487 133 3491 137
rect 111 120 115 124
rect 1823 120 1827 124
rect 1863 120 1867 124
rect 3575 120 3579 124
rect 111 103 115 107
rect 1823 103 1827 107
rect 1863 103 1867 107
rect 3575 103 3579 107
rect 167 93 171 97
rect 255 93 259 97
rect 343 93 347 97
rect 431 93 435 97
rect 519 93 523 97
rect 607 93 611 97
rect 695 93 699 97
rect 783 93 787 97
rect 871 93 875 97
rect 959 93 963 97
rect 1047 93 1051 97
rect 1135 93 1139 97
rect 1223 93 1227 97
rect 1311 93 1315 97
rect 1399 93 1403 97
rect 1495 93 1499 97
rect 1887 93 1891 97
rect 1975 93 1979 97
rect 2063 93 2067 97
rect 2151 93 2155 97
rect 2239 93 2243 97
rect 2327 93 2331 97
rect 2431 93 2435 97
rect 2535 93 2539 97
rect 2639 93 2643 97
rect 2735 93 2739 97
rect 2831 93 2835 97
rect 2927 93 2931 97
rect 3023 93 3027 97
rect 3119 93 3123 97
rect 3215 93 3219 97
rect 3303 93 3307 97
rect 3391 93 3395 97
rect 3479 93 3483 97
<< m3 >>
rect 111 3650 115 3651
rect 111 3645 115 3646
rect 239 3650 243 3651
rect 239 3645 243 3646
rect 327 3650 331 3651
rect 327 3645 331 3646
rect 415 3650 419 3651
rect 415 3645 419 3646
rect 503 3650 507 3651
rect 503 3645 507 3646
rect 591 3650 595 3651
rect 591 3645 595 3646
rect 679 3650 683 3651
rect 679 3645 683 3646
rect 1823 3650 1827 3651
rect 1823 3645 1827 3646
rect 112 3621 114 3645
rect 240 3634 242 3645
rect 328 3634 330 3645
rect 416 3634 418 3645
rect 504 3634 506 3645
rect 592 3634 594 3645
rect 680 3634 682 3645
rect 238 3633 244 3634
rect 238 3629 239 3633
rect 243 3629 244 3633
rect 238 3628 244 3629
rect 326 3633 332 3634
rect 326 3629 327 3633
rect 331 3629 332 3633
rect 326 3628 332 3629
rect 414 3633 420 3634
rect 414 3629 415 3633
rect 419 3629 420 3633
rect 414 3628 420 3629
rect 502 3633 508 3634
rect 502 3629 503 3633
rect 507 3629 508 3633
rect 502 3628 508 3629
rect 590 3633 596 3634
rect 590 3629 591 3633
rect 595 3629 596 3633
rect 590 3628 596 3629
rect 678 3633 684 3634
rect 678 3629 679 3633
rect 683 3629 684 3633
rect 678 3628 684 3629
rect 1824 3621 1826 3645
rect 110 3620 116 3621
rect 110 3616 111 3620
rect 115 3616 116 3620
rect 110 3615 116 3616
rect 1822 3620 1828 3621
rect 1822 3616 1823 3620
rect 1827 3616 1828 3620
rect 1822 3615 1828 3616
rect 110 3603 116 3604
rect 110 3599 111 3603
rect 115 3599 116 3603
rect 110 3598 116 3599
rect 1822 3603 1828 3604
rect 1822 3599 1823 3603
rect 1827 3599 1828 3603
rect 1822 3598 1828 3599
rect 112 3575 114 3598
rect 230 3593 236 3594
rect 230 3589 231 3593
rect 235 3589 236 3593
rect 230 3588 236 3589
rect 318 3593 324 3594
rect 318 3589 319 3593
rect 323 3589 324 3593
rect 318 3588 324 3589
rect 406 3593 412 3594
rect 406 3589 407 3593
rect 411 3589 412 3593
rect 406 3588 412 3589
rect 494 3593 500 3594
rect 494 3589 495 3593
rect 499 3589 500 3593
rect 494 3588 500 3589
rect 582 3593 588 3594
rect 582 3589 583 3593
rect 587 3589 588 3593
rect 582 3588 588 3589
rect 670 3593 676 3594
rect 670 3589 671 3593
rect 675 3589 676 3593
rect 670 3588 676 3589
rect 232 3575 234 3588
rect 320 3575 322 3588
rect 408 3575 410 3588
rect 496 3575 498 3588
rect 584 3575 586 3588
rect 672 3575 674 3588
rect 1824 3575 1826 3598
rect 1863 3586 1867 3587
rect 1863 3581 1867 3582
rect 1887 3586 1891 3587
rect 1887 3581 1891 3582
rect 1975 3586 1979 3587
rect 1975 3581 1979 3582
rect 2063 3586 2067 3587
rect 2063 3581 2067 3582
rect 2151 3586 2155 3587
rect 2151 3581 2155 3582
rect 2239 3586 2243 3587
rect 2239 3581 2243 3582
rect 2327 3586 2331 3587
rect 2327 3581 2331 3582
rect 2415 3586 2419 3587
rect 2415 3581 2419 3582
rect 2503 3586 2507 3587
rect 2503 3581 2507 3582
rect 2591 3586 2595 3587
rect 2591 3581 2595 3582
rect 2679 3586 2683 3587
rect 2679 3581 2683 3582
rect 2767 3586 2771 3587
rect 2767 3581 2771 3582
rect 2855 3586 2859 3587
rect 2855 3581 2859 3582
rect 2943 3586 2947 3587
rect 2943 3581 2947 3582
rect 3031 3586 3035 3587
rect 3031 3581 3035 3582
rect 3119 3586 3123 3587
rect 3119 3581 3123 3582
rect 3207 3586 3211 3587
rect 3207 3581 3211 3582
rect 3295 3586 3299 3587
rect 3295 3581 3299 3582
rect 3575 3586 3579 3587
rect 3575 3581 3579 3582
rect 111 3574 115 3575
rect 111 3569 115 3570
rect 231 3574 235 3575
rect 231 3569 235 3570
rect 247 3574 251 3575
rect 247 3569 251 3570
rect 319 3574 323 3575
rect 319 3569 323 3570
rect 399 3574 403 3575
rect 399 3569 403 3570
rect 407 3574 411 3575
rect 407 3569 411 3570
rect 495 3574 499 3575
rect 495 3569 499 3570
rect 543 3574 547 3575
rect 543 3569 547 3570
rect 583 3574 587 3575
rect 583 3569 587 3570
rect 671 3574 675 3575
rect 671 3569 675 3570
rect 687 3574 691 3575
rect 687 3569 691 3570
rect 823 3574 827 3575
rect 823 3569 827 3570
rect 951 3574 955 3575
rect 951 3569 955 3570
rect 1079 3574 1083 3575
rect 1079 3569 1083 3570
rect 1199 3574 1203 3575
rect 1199 3569 1203 3570
rect 1311 3574 1315 3575
rect 1311 3569 1315 3570
rect 1423 3574 1427 3575
rect 1423 3569 1427 3570
rect 1543 3574 1547 3575
rect 1543 3569 1547 3570
rect 1823 3574 1827 3575
rect 1823 3569 1827 3570
rect 112 3554 114 3569
rect 248 3564 250 3569
rect 400 3564 402 3569
rect 544 3564 546 3569
rect 688 3564 690 3569
rect 824 3564 826 3569
rect 952 3564 954 3569
rect 1080 3564 1082 3569
rect 1200 3564 1202 3569
rect 1312 3564 1314 3569
rect 1424 3564 1426 3569
rect 1544 3564 1546 3569
rect 246 3563 252 3564
rect 246 3559 247 3563
rect 251 3559 252 3563
rect 246 3558 252 3559
rect 398 3563 404 3564
rect 398 3559 399 3563
rect 403 3559 404 3563
rect 398 3558 404 3559
rect 542 3563 548 3564
rect 542 3559 543 3563
rect 547 3559 548 3563
rect 542 3558 548 3559
rect 686 3563 692 3564
rect 686 3559 687 3563
rect 691 3559 692 3563
rect 686 3558 692 3559
rect 822 3563 828 3564
rect 822 3559 823 3563
rect 827 3559 828 3563
rect 822 3558 828 3559
rect 950 3563 956 3564
rect 950 3559 951 3563
rect 955 3559 956 3563
rect 950 3558 956 3559
rect 1078 3563 1084 3564
rect 1078 3559 1079 3563
rect 1083 3559 1084 3563
rect 1078 3558 1084 3559
rect 1198 3563 1204 3564
rect 1198 3559 1199 3563
rect 1203 3559 1204 3563
rect 1198 3558 1204 3559
rect 1310 3563 1316 3564
rect 1310 3559 1311 3563
rect 1315 3559 1316 3563
rect 1310 3558 1316 3559
rect 1422 3563 1428 3564
rect 1422 3559 1423 3563
rect 1427 3559 1428 3563
rect 1422 3558 1428 3559
rect 1542 3563 1548 3564
rect 1542 3559 1543 3563
rect 1547 3559 1548 3563
rect 1542 3558 1548 3559
rect 1824 3554 1826 3569
rect 1864 3566 1866 3581
rect 1888 3576 1890 3581
rect 1976 3576 1978 3581
rect 2064 3576 2066 3581
rect 2152 3576 2154 3581
rect 2240 3576 2242 3581
rect 2328 3576 2330 3581
rect 2416 3576 2418 3581
rect 2504 3576 2506 3581
rect 2592 3576 2594 3581
rect 2680 3576 2682 3581
rect 2768 3576 2770 3581
rect 2856 3576 2858 3581
rect 2944 3576 2946 3581
rect 3032 3576 3034 3581
rect 3120 3576 3122 3581
rect 3208 3576 3210 3581
rect 3296 3576 3298 3581
rect 1886 3575 1892 3576
rect 1886 3571 1887 3575
rect 1891 3571 1892 3575
rect 1886 3570 1892 3571
rect 1974 3575 1980 3576
rect 1974 3571 1975 3575
rect 1979 3571 1980 3575
rect 1974 3570 1980 3571
rect 2062 3575 2068 3576
rect 2062 3571 2063 3575
rect 2067 3571 2068 3575
rect 2062 3570 2068 3571
rect 2150 3575 2156 3576
rect 2150 3571 2151 3575
rect 2155 3571 2156 3575
rect 2150 3570 2156 3571
rect 2238 3575 2244 3576
rect 2238 3571 2239 3575
rect 2243 3571 2244 3575
rect 2238 3570 2244 3571
rect 2326 3575 2332 3576
rect 2326 3571 2327 3575
rect 2331 3571 2332 3575
rect 2326 3570 2332 3571
rect 2414 3575 2420 3576
rect 2414 3571 2415 3575
rect 2419 3571 2420 3575
rect 2414 3570 2420 3571
rect 2502 3575 2508 3576
rect 2502 3571 2503 3575
rect 2507 3571 2508 3575
rect 2502 3570 2508 3571
rect 2590 3575 2596 3576
rect 2590 3571 2591 3575
rect 2595 3571 2596 3575
rect 2590 3570 2596 3571
rect 2678 3575 2684 3576
rect 2678 3571 2679 3575
rect 2683 3571 2684 3575
rect 2678 3570 2684 3571
rect 2766 3575 2772 3576
rect 2766 3571 2767 3575
rect 2771 3571 2772 3575
rect 2766 3570 2772 3571
rect 2854 3575 2860 3576
rect 2854 3571 2855 3575
rect 2859 3571 2860 3575
rect 2854 3570 2860 3571
rect 2942 3575 2948 3576
rect 2942 3571 2943 3575
rect 2947 3571 2948 3575
rect 2942 3570 2948 3571
rect 3030 3575 3036 3576
rect 3030 3571 3031 3575
rect 3035 3571 3036 3575
rect 3030 3570 3036 3571
rect 3118 3575 3124 3576
rect 3118 3571 3119 3575
rect 3123 3571 3124 3575
rect 3118 3570 3124 3571
rect 3206 3575 3212 3576
rect 3206 3571 3207 3575
rect 3211 3571 3212 3575
rect 3206 3570 3212 3571
rect 3294 3575 3300 3576
rect 3294 3571 3295 3575
rect 3299 3571 3300 3575
rect 3294 3570 3300 3571
rect 3576 3566 3578 3581
rect 1862 3565 1868 3566
rect 1862 3561 1863 3565
rect 1867 3561 1868 3565
rect 1862 3560 1868 3561
rect 3574 3565 3580 3566
rect 3574 3561 3575 3565
rect 3579 3561 3580 3565
rect 3574 3560 3580 3561
rect 110 3553 116 3554
rect 110 3549 111 3553
rect 115 3549 116 3553
rect 110 3548 116 3549
rect 1822 3553 1828 3554
rect 1822 3549 1823 3553
rect 1827 3549 1828 3553
rect 1822 3548 1828 3549
rect 1862 3548 1868 3549
rect 1862 3544 1863 3548
rect 1867 3544 1868 3548
rect 1862 3543 1868 3544
rect 3574 3548 3580 3549
rect 3574 3544 3575 3548
rect 3579 3544 3580 3548
rect 3574 3543 3580 3544
rect 110 3536 116 3537
rect 110 3532 111 3536
rect 115 3532 116 3536
rect 110 3531 116 3532
rect 1822 3536 1828 3537
rect 1822 3532 1823 3536
rect 1827 3532 1828 3536
rect 1822 3531 1828 3532
rect 112 3507 114 3531
rect 254 3523 260 3524
rect 254 3519 255 3523
rect 259 3519 260 3523
rect 254 3518 260 3519
rect 406 3523 412 3524
rect 406 3519 407 3523
rect 411 3519 412 3523
rect 406 3518 412 3519
rect 550 3523 556 3524
rect 550 3519 551 3523
rect 555 3519 556 3523
rect 550 3518 556 3519
rect 694 3523 700 3524
rect 694 3519 695 3523
rect 699 3519 700 3523
rect 694 3518 700 3519
rect 830 3523 836 3524
rect 830 3519 831 3523
rect 835 3519 836 3523
rect 830 3518 836 3519
rect 958 3523 964 3524
rect 958 3519 959 3523
rect 963 3519 964 3523
rect 958 3518 964 3519
rect 1086 3523 1092 3524
rect 1086 3519 1087 3523
rect 1091 3519 1092 3523
rect 1086 3518 1092 3519
rect 1206 3523 1212 3524
rect 1206 3519 1207 3523
rect 1211 3519 1212 3523
rect 1206 3518 1212 3519
rect 1318 3523 1324 3524
rect 1318 3519 1319 3523
rect 1323 3519 1324 3523
rect 1318 3518 1324 3519
rect 1430 3523 1436 3524
rect 1430 3519 1431 3523
rect 1435 3519 1436 3523
rect 1430 3518 1436 3519
rect 1550 3523 1556 3524
rect 1550 3519 1551 3523
rect 1555 3519 1556 3523
rect 1550 3518 1556 3519
rect 256 3507 258 3518
rect 408 3507 410 3518
rect 552 3507 554 3518
rect 696 3507 698 3518
rect 832 3507 834 3518
rect 960 3507 962 3518
rect 1088 3507 1090 3518
rect 1208 3507 1210 3518
rect 1320 3507 1322 3518
rect 1432 3507 1434 3518
rect 1552 3507 1554 3518
rect 1824 3507 1826 3531
rect 1864 3511 1866 3543
rect 1894 3535 1900 3536
rect 1894 3531 1895 3535
rect 1899 3531 1900 3535
rect 1894 3530 1900 3531
rect 1982 3535 1988 3536
rect 1982 3531 1983 3535
rect 1987 3531 1988 3535
rect 1982 3530 1988 3531
rect 2070 3535 2076 3536
rect 2070 3531 2071 3535
rect 2075 3531 2076 3535
rect 2070 3530 2076 3531
rect 2158 3535 2164 3536
rect 2158 3531 2159 3535
rect 2163 3531 2164 3535
rect 2158 3530 2164 3531
rect 2246 3535 2252 3536
rect 2246 3531 2247 3535
rect 2251 3531 2252 3535
rect 2246 3530 2252 3531
rect 2334 3535 2340 3536
rect 2334 3531 2335 3535
rect 2339 3531 2340 3535
rect 2334 3530 2340 3531
rect 2422 3535 2428 3536
rect 2422 3531 2423 3535
rect 2427 3531 2428 3535
rect 2422 3530 2428 3531
rect 2510 3535 2516 3536
rect 2510 3531 2511 3535
rect 2515 3531 2516 3535
rect 2510 3530 2516 3531
rect 2598 3535 2604 3536
rect 2598 3531 2599 3535
rect 2603 3531 2604 3535
rect 2598 3530 2604 3531
rect 2686 3535 2692 3536
rect 2686 3531 2687 3535
rect 2691 3531 2692 3535
rect 2686 3530 2692 3531
rect 2774 3535 2780 3536
rect 2774 3531 2775 3535
rect 2779 3531 2780 3535
rect 2774 3530 2780 3531
rect 2862 3535 2868 3536
rect 2862 3531 2863 3535
rect 2867 3531 2868 3535
rect 2862 3530 2868 3531
rect 2950 3535 2956 3536
rect 2950 3531 2951 3535
rect 2955 3531 2956 3535
rect 2950 3530 2956 3531
rect 3038 3535 3044 3536
rect 3038 3531 3039 3535
rect 3043 3531 3044 3535
rect 3038 3530 3044 3531
rect 3126 3535 3132 3536
rect 3126 3531 3127 3535
rect 3131 3531 3132 3535
rect 3126 3530 3132 3531
rect 3214 3535 3220 3536
rect 3214 3531 3215 3535
rect 3219 3531 3220 3535
rect 3214 3530 3220 3531
rect 3302 3535 3308 3536
rect 3302 3531 3303 3535
rect 3307 3531 3308 3535
rect 3302 3530 3308 3531
rect 1896 3511 1898 3530
rect 1984 3511 1986 3530
rect 2072 3511 2074 3530
rect 2160 3511 2162 3530
rect 2248 3511 2250 3530
rect 2336 3511 2338 3530
rect 2424 3511 2426 3530
rect 2512 3511 2514 3530
rect 2600 3511 2602 3530
rect 2688 3511 2690 3530
rect 2776 3511 2778 3530
rect 2864 3511 2866 3530
rect 2952 3511 2954 3530
rect 3040 3511 3042 3530
rect 3128 3511 3130 3530
rect 3216 3511 3218 3530
rect 3304 3511 3306 3530
rect 3576 3511 3578 3543
rect 1863 3510 1867 3511
rect 111 3506 115 3507
rect 111 3501 115 3502
rect 183 3506 187 3507
rect 183 3501 187 3502
rect 255 3506 259 3507
rect 255 3501 259 3502
rect 351 3506 355 3507
rect 351 3501 355 3502
rect 407 3506 411 3507
rect 407 3501 411 3502
rect 519 3506 523 3507
rect 519 3501 523 3502
rect 551 3506 555 3507
rect 551 3501 555 3502
rect 679 3506 683 3507
rect 679 3501 683 3502
rect 695 3506 699 3507
rect 695 3501 699 3502
rect 831 3506 835 3507
rect 831 3501 835 3502
rect 959 3506 963 3507
rect 959 3501 963 3502
rect 967 3506 971 3507
rect 967 3501 971 3502
rect 1087 3506 1091 3507
rect 1087 3501 1091 3502
rect 1095 3506 1099 3507
rect 1095 3501 1099 3502
rect 1207 3506 1211 3507
rect 1207 3501 1211 3502
rect 1215 3506 1219 3507
rect 1215 3501 1219 3502
rect 1319 3506 1323 3507
rect 1319 3501 1323 3502
rect 1335 3506 1339 3507
rect 1335 3501 1339 3502
rect 1431 3506 1435 3507
rect 1431 3501 1435 3502
rect 1455 3506 1459 3507
rect 1455 3501 1459 3502
rect 1551 3506 1555 3507
rect 1551 3501 1555 3502
rect 1575 3506 1579 3507
rect 1575 3501 1579 3502
rect 1823 3506 1827 3507
rect 1863 3505 1867 3506
rect 1895 3510 1899 3511
rect 1895 3505 1899 3506
rect 1911 3510 1915 3511
rect 1911 3505 1915 3506
rect 1983 3510 1987 3511
rect 1983 3505 1987 3506
rect 2015 3510 2019 3511
rect 2015 3505 2019 3506
rect 2071 3510 2075 3511
rect 2071 3505 2075 3506
rect 2135 3510 2139 3511
rect 2135 3505 2139 3506
rect 2159 3510 2163 3511
rect 2159 3505 2163 3506
rect 2247 3510 2251 3511
rect 2247 3505 2251 3506
rect 2263 3510 2267 3511
rect 2263 3505 2267 3506
rect 2335 3510 2339 3511
rect 2335 3505 2339 3506
rect 2391 3510 2395 3511
rect 2391 3505 2395 3506
rect 2423 3510 2427 3511
rect 2423 3505 2427 3506
rect 2511 3510 2515 3511
rect 2511 3505 2515 3506
rect 2527 3510 2531 3511
rect 2527 3505 2531 3506
rect 2599 3510 2603 3511
rect 2599 3505 2603 3506
rect 2663 3510 2667 3511
rect 2663 3505 2667 3506
rect 2687 3510 2691 3511
rect 2687 3505 2691 3506
rect 2775 3510 2779 3511
rect 2775 3505 2779 3506
rect 2799 3510 2803 3511
rect 2799 3505 2803 3506
rect 2863 3510 2867 3511
rect 2863 3505 2867 3506
rect 2943 3510 2947 3511
rect 2943 3505 2947 3506
rect 2951 3510 2955 3511
rect 2951 3505 2955 3506
rect 3039 3510 3043 3511
rect 3039 3505 3043 3506
rect 3087 3510 3091 3511
rect 3087 3505 3091 3506
rect 3127 3510 3131 3511
rect 3127 3505 3131 3506
rect 3215 3510 3219 3511
rect 3215 3505 3219 3506
rect 3303 3510 3307 3511
rect 3303 3505 3307 3506
rect 3575 3510 3579 3511
rect 3575 3505 3579 3506
rect 1823 3501 1827 3502
rect 112 3477 114 3501
rect 184 3490 186 3501
rect 352 3490 354 3501
rect 520 3490 522 3501
rect 680 3490 682 3501
rect 832 3490 834 3501
rect 968 3490 970 3501
rect 1096 3490 1098 3501
rect 1216 3490 1218 3501
rect 1336 3490 1338 3501
rect 1456 3490 1458 3501
rect 1576 3490 1578 3501
rect 182 3489 188 3490
rect 182 3485 183 3489
rect 187 3485 188 3489
rect 182 3484 188 3485
rect 350 3489 356 3490
rect 350 3485 351 3489
rect 355 3485 356 3489
rect 350 3484 356 3485
rect 518 3489 524 3490
rect 518 3485 519 3489
rect 523 3485 524 3489
rect 518 3484 524 3485
rect 678 3489 684 3490
rect 678 3485 679 3489
rect 683 3485 684 3489
rect 678 3484 684 3485
rect 830 3489 836 3490
rect 830 3485 831 3489
rect 835 3485 836 3489
rect 830 3484 836 3485
rect 966 3489 972 3490
rect 966 3485 967 3489
rect 971 3485 972 3489
rect 966 3484 972 3485
rect 1094 3489 1100 3490
rect 1094 3485 1095 3489
rect 1099 3485 1100 3489
rect 1094 3484 1100 3485
rect 1214 3489 1220 3490
rect 1214 3485 1215 3489
rect 1219 3485 1220 3489
rect 1214 3484 1220 3485
rect 1334 3489 1340 3490
rect 1334 3485 1335 3489
rect 1339 3485 1340 3489
rect 1334 3484 1340 3485
rect 1454 3489 1460 3490
rect 1454 3485 1455 3489
rect 1459 3485 1460 3489
rect 1454 3484 1460 3485
rect 1574 3489 1580 3490
rect 1574 3485 1575 3489
rect 1579 3485 1580 3489
rect 1574 3484 1580 3485
rect 1824 3477 1826 3501
rect 1864 3481 1866 3505
rect 1912 3494 1914 3505
rect 2016 3494 2018 3505
rect 2136 3494 2138 3505
rect 2264 3494 2266 3505
rect 2392 3494 2394 3505
rect 2528 3494 2530 3505
rect 2664 3494 2666 3505
rect 2800 3494 2802 3505
rect 2944 3494 2946 3505
rect 3088 3494 3090 3505
rect 1910 3493 1916 3494
rect 1910 3489 1911 3493
rect 1915 3489 1916 3493
rect 1910 3488 1916 3489
rect 2014 3493 2020 3494
rect 2014 3489 2015 3493
rect 2019 3489 2020 3493
rect 2014 3488 2020 3489
rect 2134 3493 2140 3494
rect 2134 3489 2135 3493
rect 2139 3489 2140 3493
rect 2134 3488 2140 3489
rect 2262 3493 2268 3494
rect 2262 3489 2263 3493
rect 2267 3489 2268 3493
rect 2262 3488 2268 3489
rect 2390 3493 2396 3494
rect 2390 3489 2391 3493
rect 2395 3489 2396 3493
rect 2390 3488 2396 3489
rect 2526 3493 2532 3494
rect 2526 3489 2527 3493
rect 2531 3489 2532 3493
rect 2526 3488 2532 3489
rect 2662 3493 2668 3494
rect 2662 3489 2663 3493
rect 2667 3489 2668 3493
rect 2662 3488 2668 3489
rect 2798 3493 2804 3494
rect 2798 3489 2799 3493
rect 2803 3489 2804 3493
rect 2798 3488 2804 3489
rect 2942 3493 2948 3494
rect 2942 3489 2943 3493
rect 2947 3489 2948 3493
rect 2942 3488 2948 3489
rect 3086 3493 3092 3494
rect 3086 3489 3087 3493
rect 3091 3489 3092 3493
rect 3086 3488 3092 3489
rect 3576 3481 3578 3505
rect 1862 3480 1868 3481
rect 110 3476 116 3477
rect 110 3472 111 3476
rect 115 3472 116 3476
rect 110 3471 116 3472
rect 1822 3476 1828 3477
rect 1822 3472 1823 3476
rect 1827 3472 1828 3476
rect 1862 3476 1863 3480
rect 1867 3476 1868 3480
rect 1862 3475 1868 3476
rect 3574 3480 3580 3481
rect 3574 3476 3575 3480
rect 3579 3476 3580 3480
rect 3574 3475 3580 3476
rect 1822 3471 1828 3472
rect 1862 3463 1868 3464
rect 110 3459 116 3460
rect 110 3455 111 3459
rect 115 3455 116 3459
rect 110 3454 116 3455
rect 1822 3459 1828 3460
rect 1822 3455 1823 3459
rect 1827 3455 1828 3459
rect 1862 3459 1863 3463
rect 1867 3459 1868 3463
rect 1862 3458 1868 3459
rect 3574 3463 3580 3464
rect 3574 3459 3575 3463
rect 3579 3459 3580 3463
rect 3574 3458 3580 3459
rect 1822 3454 1828 3455
rect 112 3439 114 3454
rect 174 3449 180 3450
rect 174 3445 175 3449
rect 179 3445 180 3449
rect 174 3444 180 3445
rect 342 3449 348 3450
rect 342 3445 343 3449
rect 347 3445 348 3449
rect 342 3444 348 3445
rect 510 3449 516 3450
rect 510 3445 511 3449
rect 515 3445 516 3449
rect 510 3444 516 3445
rect 670 3449 676 3450
rect 670 3445 671 3449
rect 675 3445 676 3449
rect 670 3444 676 3445
rect 822 3449 828 3450
rect 822 3445 823 3449
rect 827 3445 828 3449
rect 822 3444 828 3445
rect 958 3449 964 3450
rect 958 3445 959 3449
rect 963 3445 964 3449
rect 958 3444 964 3445
rect 1086 3449 1092 3450
rect 1086 3445 1087 3449
rect 1091 3445 1092 3449
rect 1086 3444 1092 3445
rect 1206 3449 1212 3450
rect 1206 3445 1207 3449
rect 1211 3445 1212 3449
rect 1206 3444 1212 3445
rect 1326 3449 1332 3450
rect 1326 3445 1327 3449
rect 1331 3445 1332 3449
rect 1326 3444 1332 3445
rect 1446 3449 1452 3450
rect 1446 3445 1447 3449
rect 1451 3445 1452 3449
rect 1446 3444 1452 3445
rect 1566 3449 1572 3450
rect 1566 3445 1567 3449
rect 1571 3445 1572 3449
rect 1566 3444 1572 3445
rect 176 3439 178 3444
rect 344 3439 346 3444
rect 512 3439 514 3444
rect 672 3439 674 3444
rect 824 3439 826 3444
rect 960 3439 962 3444
rect 1088 3439 1090 3444
rect 1208 3439 1210 3444
rect 1328 3439 1330 3444
rect 1448 3439 1450 3444
rect 1568 3439 1570 3444
rect 1824 3439 1826 3454
rect 111 3438 115 3439
rect 111 3433 115 3434
rect 135 3438 139 3439
rect 135 3433 139 3434
rect 175 3438 179 3439
rect 175 3433 179 3434
rect 255 3438 259 3439
rect 255 3433 259 3434
rect 343 3438 347 3439
rect 343 3433 347 3434
rect 415 3438 419 3439
rect 415 3433 419 3434
rect 511 3438 515 3439
rect 511 3433 515 3434
rect 583 3438 587 3439
rect 583 3433 587 3434
rect 671 3438 675 3439
rect 671 3433 675 3434
rect 759 3438 763 3439
rect 759 3433 763 3434
rect 823 3438 827 3439
rect 823 3433 827 3434
rect 935 3438 939 3439
rect 935 3433 939 3434
rect 959 3438 963 3439
rect 959 3433 963 3434
rect 1087 3438 1091 3439
rect 1087 3433 1091 3434
rect 1111 3438 1115 3439
rect 1111 3433 1115 3434
rect 1207 3438 1211 3439
rect 1207 3433 1211 3434
rect 1295 3438 1299 3439
rect 1295 3433 1299 3434
rect 1327 3438 1331 3439
rect 1327 3433 1331 3434
rect 1447 3438 1451 3439
rect 1447 3433 1451 3434
rect 1479 3438 1483 3439
rect 1479 3433 1483 3434
rect 1567 3438 1571 3439
rect 1567 3433 1571 3434
rect 1823 3438 1827 3439
rect 1864 3435 1866 3458
rect 1902 3453 1908 3454
rect 1902 3449 1903 3453
rect 1907 3449 1908 3453
rect 1902 3448 1908 3449
rect 2006 3453 2012 3454
rect 2006 3449 2007 3453
rect 2011 3449 2012 3453
rect 2006 3448 2012 3449
rect 2126 3453 2132 3454
rect 2126 3449 2127 3453
rect 2131 3449 2132 3453
rect 2126 3448 2132 3449
rect 2254 3453 2260 3454
rect 2254 3449 2255 3453
rect 2259 3449 2260 3453
rect 2254 3448 2260 3449
rect 2382 3453 2388 3454
rect 2382 3449 2383 3453
rect 2387 3449 2388 3453
rect 2382 3448 2388 3449
rect 2518 3453 2524 3454
rect 2518 3449 2519 3453
rect 2523 3449 2524 3453
rect 2518 3448 2524 3449
rect 2654 3453 2660 3454
rect 2654 3449 2655 3453
rect 2659 3449 2660 3453
rect 2654 3448 2660 3449
rect 2790 3453 2796 3454
rect 2790 3449 2791 3453
rect 2795 3449 2796 3453
rect 2790 3448 2796 3449
rect 2934 3453 2940 3454
rect 2934 3449 2935 3453
rect 2939 3449 2940 3453
rect 2934 3448 2940 3449
rect 3078 3453 3084 3454
rect 3078 3449 3079 3453
rect 3083 3449 3084 3453
rect 3078 3448 3084 3449
rect 1904 3435 1906 3448
rect 2008 3435 2010 3448
rect 2128 3435 2130 3448
rect 2256 3435 2258 3448
rect 2384 3435 2386 3448
rect 2520 3435 2522 3448
rect 2656 3435 2658 3448
rect 2792 3435 2794 3448
rect 2936 3435 2938 3448
rect 3080 3435 3082 3448
rect 3576 3435 3578 3458
rect 1823 3433 1827 3434
rect 1863 3434 1867 3435
rect 112 3418 114 3433
rect 136 3428 138 3433
rect 256 3428 258 3433
rect 416 3428 418 3433
rect 584 3428 586 3433
rect 760 3428 762 3433
rect 936 3428 938 3433
rect 1112 3428 1114 3433
rect 1296 3428 1298 3433
rect 1480 3428 1482 3433
rect 134 3427 140 3428
rect 134 3423 135 3427
rect 139 3423 140 3427
rect 134 3422 140 3423
rect 254 3427 260 3428
rect 254 3423 255 3427
rect 259 3423 260 3427
rect 254 3422 260 3423
rect 414 3427 420 3428
rect 414 3423 415 3427
rect 419 3423 420 3427
rect 414 3422 420 3423
rect 582 3427 588 3428
rect 582 3423 583 3427
rect 587 3423 588 3427
rect 582 3422 588 3423
rect 758 3427 764 3428
rect 758 3423 759 3427
rect 763 3423 764 3427
rect 758 3422 764 3423
rect 934 3427 940 3428
rect 934 3423 935 3427
rect 939 3423 940 3427
rect 934 3422 940 3423
rect 1110 3427 1116 3428
rect 1110 3423 1111 3427
rect 1115 3423 1116 3427
rect 1110 3422 1116 3423
rect 1294 3427 1300 3428
rect 1294 3423 1295 3427
rect 1299 3423 1300 3427
rect 1294 3422 1300 3423
rect 1478 3427 1484 3428
rect 1478 3423 1479 3427
rect 1483 3423 1484 3427
rect 1478 3422 1484 3423
rect 1824 3418 1826 3433
rect 1863 3429 1867 3430
rect 1903 3434 1907 3435
rect 1903 3429 1907 3430
rect 1911 3434 1915 3435
rect 1911 3429 1915 3430
rect 2007 3434 2011 3435
rect 2007 3429 2011 3430
rect 2071 3434 2075 3435
rect 2071 3429 2075 3430
rect 2127 3434 2131 3435
rect 2127 3429 2131 3430
rect 2223 3434 2227 3435
rect 2223 3429 2227 3430
rect 2255 3434 2259 3435
rect 2255 3429 2259 3430
rect 2367 3434 2371 3435
rect 2367 3429 2371 3430
rect 2383 3434 2387 3435
rect 2383 3429 2387 3430
rect 2503 3434 2507 3435
rect 2503 3429 2507 3430
rect 2519 3434 2523 3435
rect 2519 3429 2523 3430
rect 2631 3434 2635 3435
rect 2631 3429 2635 3430
rect 2655 3434 2659 3435
rect 2655 3429 2659 3430
rect 2759 3434 2763 3435
rect 2759 3429 2763 3430
rect 2791 3434 2795 3435
rect 2791 3429 2795 3430
rect 2887 3434 2891 3435
rect 2887 3429 2891 3430
rect 2935 3434 2939 3435
rect 2935 3429 2939 3430
rect 3023 3434 3027 3435
rect 3023 3429 3027 3430
rect 3079 3434 3083 3435
rect 3079 3429 3083 3430
rect 3575 3434 3579 3435
rect 3575 3429 3579 3430
rect 110 3417 116 3418
rect 110 3413 111 3417
rect 115 3413 116 3417
rect 110 3412 116 3413
rect 1822 3417 1828 3418
rect 1822 3413 1823 3417
rect 1827 3413 1828 3417
rect 1864 3414 1866 3429
rect 1912 3424 1914 3429
rect 2072 3424 2074 3429
rect 2224 3424 2226 3429
rect 2368 3424 2370 3429
rect 2504 3424 2506 3429
rect 2632 3424 2634 3429
rect 2760 3424 2762 3429
rect 2888 3424 2890 3429
rect 3024 3424 3026 3429
rect 1910 3423 1916 3424
rect 1910 3419 1911 3423
rect 1915 3419 1916 3423
rect 1910 3418 1916 3419
rect 2070 3423 2076 3424
rect 2070 3419 2071 3423
rect 2075 3419 2076 3423
rect 2070 3418 2076 3419
rect 2222 3423 2228 3424
rect 2222 3419 2223 3423
rect 2227 3419 2228 3423
rect 2222 3418 2228 3419
rect 2366 3423 2372 3424
rect 2366 3419 2367 3423
rect 2371 3419 2372 3423
rect 2366 3418 2372 3419
rect 2502 3423 2508 3424
rect 2502 3419 2503 3423
rect 2507 3419 2508 3423
rect 2502 3418 2508 3419
rect 2630 3423 2636 3424
rect 2630 3419 2631 3423
rect 2635 3419 2636 3423
rect 2630 3418 2636 3419
rect 2758 3423 2764 3424
rect 2758 3419 2759 3423
rect 2763 3419 2764 3423
rect 2758 3418 2764 3419
rect 2886 3423 2892 3424
rect 2886 3419 2887 3423
rect 2891 3419 2892 3423
rect 2886 3418 2892 3419
rect 3022 3423 3028 3424
rect 3022 3419 3023 3423
rect 3027 3419 3028 3423
rect 3022 3418 3028 3419
rect 3576 3414 3578 3429
rect 1822 3412 1828 3413
rect 1862 3413 1868 3414
rect 1862 3409 1863 3413
rect 1867 3409 1868 3413
rect 1862 3408 1868 3409
rect 3574 3413 3580 3414
rect 3574 3409 3575 3413
rect 3579 3409 3580 3413
rect 3574 3408 3580 3409
rect 110 3400 116 3401
rect 110 3396 111 3400
rect 115 3396 116 3400
rect 110 3395 116 3396
rect 1822 3400 1828 3401
rect 1822 3396 1823 3400
rect 1827 3396 1828 3400
rect 1822 3395 1828 3396
rect 1862 3396 1868 3397
rect 112 3363 114 3395
rect 142 3387 148 3388
rect 142 3383 143 3387
rect 147 3383 148 3387
rect 142 3382 148 3383
rect 262 3387 268 3388
rect 262 3383 263 3387
rect 267 3383 268 3387
rect 262 3382 268 3383
rect 422 3387 428 3388
rect 422 3383 423 3387
rect 427 3383 428 3387
rect 422 3382 428 3383
rect 590 3387 596 3388
rect 590 3383 591 3387
rect 595 3383 596 3387
rect 590 3382 596 3383
rect 766 3387 772 3388
rect 766 3383 767 3387
rect 771 3383 772 3387
rect 766 3382 772 3383
rect 942 3387 948 3388
rect 942 3383 943 3387
rect 947 3383 948 3387
rect 942 3382 948 3383
rect 1118 3387 1124 3388
rect 1118 3383 1119 3387
rect 1123 3383 1124 3387
rect 1118 3382 1124 3383
rect 1302 3387 1308 3388
rect 1302 3383 1303 3387
rect 1307 3383 1308 3387
rect 1302 3382 1308 3383
rect 1486 3387 1492 3388
rect 1486 3383 1487 3387
rect 1491 3383 1492 3387
rect 1486 3382 1492 3383
rect 144 3363 146 3382
rect 264 3363 266 3382
rect 424 3363 426 3382
rect 592 3363 594 3382
rect 768 3363 770 3382
rect 944 3363 946 3382
rect 1120 3363 1122 3382
rect 1304 3363 1306 3382
rect 1488 3363 1490 3382
rect 1824 3363 1826 3395
rect 1862 3392 1863 3396
rect 1867 3392 1868 3396
rect 1862 3391 1868 3392
rect 3574 3396 3580 3397
rect 3574 3392 3575 3396
rect 3579 3392 3580 3396
rect 3574 3391 3580 3392
rect 1864 3363 1866 3391
rect 1918 3383 1924 3384
rect 1918 3379 1919 3383
rect 1923 3379 1924 3383
rect 1918 3378 1924 3379
rect 2078 3383 2084 3384
rect 2078 3379 2079 3383
rect 2083 3379 2084 3383
rect 2078 3378 2084 3379
rect 2230 3383 2236 3384
rect 2230 3379 2231 3383
rect 2235 3379 2236 3383
rect 2230 3378 2236 3379
rect 2374 3383 2380 3384
rect 2374 3379 2375 3383
rect 2379 3379 2380 3383
rect 2374 3378 2380 3379
rect 2510 3383 2516 3384
rect 2510 3379 2511 3383
rect 2515 3379 2516 3383
rect 2510 3378 2516 3379
rect 2638 3383 2644 3384
rect 2638 3379 2639 3383
rect 2643 3379 2644 3383
rect 2638 3378 2644 3379
rect 2766 3383 2772 3384
rect 2766 3379 2767 3383
rect 2771 3379 2772 3383
rect 2766 3378 2772 3379
rect 2894 3383 2900 3384
rect 2894 3379 2895 3383
rect 2899 3379 2900 3383
rect 2894 3378 2900 3379
rect 3030 3383 3036 3384
rect 3030 3379 3031 3383
rect 3035 3379 3036 3383
rect 3030 3378 3036 3379
rect 1920 3363 1922 3378
rect 2080 3363 2082 3378
rect 2232 3363 2234 3378
rect 2376 3363 2378 3378
rect 2512 3363 2514 3378
rect 2640 3363 2642 3378
rect 2768 3363 2770 3378
rect 2896 3363 2898 3378
rect 3032 3363 3034 3378
rect 3576 3363 3578 3391
rect 111 3362 115 3363
rect 111 3357 115 3358
rect 143 3362 147 3363
rect 143 3357 147 3358
rect 207 3362 211 3363
rect 207 3357 211 3358
rect 263 3362 267 3363
rect 263 3357 267 3358
rect 367 3362 371 3363
rect 367 3357 371 3358
rect 423 3362 427 3363
rect 423 3357 427 3358
rect 535 3362 539 3363
rect 535 3357 539 3358
rect 591 3362 595 3363
rect 591 3357 595 3358
rect 695 3362 699 3363
rect 695 3357 699 3358
rect 767 3362 771 3363
rect 767 3357 771 3358
rect 855 3362 859 3363
rect 855 3357 859 3358
rect 943 3362 947 3363
rect 943 3357 947 3358
rect 999 3362 1003 3363
rect 999 3357 1003 3358
rect 1119 3362 1123 3363
rect 1119 3357 1123 3358
rect 1143 3362 1147 3363
rect 1143 3357 1147 3358
rect 1279 3362 1283 3363
rect 1279 3357 1283 3358
rect 1303 3362 1307 3363
rect 1303 3357 1307 3358
rect 1415 3362 1419 3363
rect 1415 3357 1419 3358
rect 1487 3362 1491 3363
rect 1487 3357 1491 3358
rect 1559 3362 1563 3363
rect 1559 3357 1563 3358
rect 1823 3362 1827 3363
rect 1823 3357 1827 3358
rect 1863 3362 1867 3363
rect 1863 3357 1867 3358
rect 1895 3362 1899 3363
rect 1895 3357 1899 3358
rect 1919 3362 1923 3363
rect 1919 3357 1923 3358
rect 2047 3362 2051 3363
rect 2047 3357 2051 3358
rect 2079 3362 2083 3363
rect 2079 3357 2083 3358
rect 2207 3362 2211 3363
rect 2207 3357 2211 3358
rect 2231 3362 2235 3363
rect 2231 3357 2235 3358
rect 2367 3362 2371 3363
rect 2367 3357 2371 3358
rect 2375 3362 2379 3363
rect 2375 3357 2379 3358
rect 2511 3362 2515 3363
rect 2511 3357 2515 3358
rect 2535 3362 2539 3363
rect 2535 3357 2539 3358
rect 2639 3362 2643 3363
rect 2639 3357 2643 3358
rect 2703 3362 2707 3363
rect 2703 3357 2707 3358
rect 2767 3362 2771 3363
rect 2767 3357 2771 3358
rect 2879 3362 2883 3363
rect 2879 3357 2883 3358
rect 2895 3362 2899 3363
rect 2895 3357 2899 3358
rect 3031 3362 3035 3363
rect 3031 3357 3035 3358
rect 3055 3362 3059 3363
rect 3055 3357 3059 3358
rect 3575 3362 3579 3363
rect 3575 3357 3579 3358
rect 112 3333 114 3357
rect 208 3346 210 3357
rect 368 3346 370 3357
rect 536 3346 538 3357
rect 696 3346 698 3357
rect 856 3346 858 3357
rect 1000 3346 1002 3357
rect 1144 3346 1146 3357
rect 1280 3346 1282 3357
rect 1416 3346 1418 3357
rect 1560 3346 1562 3357
rect 206 3345 212 3346
rect 206 3341 207 3345
rect 211 3341 212 3345
rect 206 3340 212 3341
rect 366 3345 372 3346
rect 366 3341 367 3345
rect 371 3341 372 3345
rect 366 3340 372 3341
rect 534 3345 540 3346
rect 534 3341 535 3345
rect 539 3341 540 3345
rect 534 3340 540 3341
rect 694 3345 700 3346
rect 694 3341 695 3345
rect 699 3341 700 3345
rect 694 3340 700 3341
rect 854 3345 860 3346
rect 854 3341 855 3345
rect 859 3341 860 3345
rect 854 3340 860 3341
rect 998 3345 1004 3346
rect 998 3341 999 3345
rect 1003 3341 1004 3345
rect 998 3340 1004 3341
rect 1142 3345 1148 3346
rect 1142 3341 1143 3345
rect 1147 3341 1148 3345
rect 1142 3340 1148 3341
rect 1278 3345 1284 3346
rect 1278 3341 1279 3345
rect 1283 3341 1284 3345
rect 1278 3340 1284 3341
rect 1414 3345 1420 3346
rect 1414 3341 1415 3345
rect 1419 3341 1420 3345
rect 1414 3340 1420 3341
rect 1558 3345 1564 3346
rect 1558 3341 1559 3345
rect 1563 3341 1564 3345
rect 1558 3340 1564 3341
rect 1824 3333 1826 3357
rect 1864 3333 1866 3357
rect 1896 3346 1898 3357
rect 2048 3346 2050 3357
rect 2208 3346 2210 3357
rect 2368 3346 2370 3357
rect 2536 3346 2538 3357
rect 2704 3346 2706 3357
rect 2880 3346 2882 3357
rect 3056 3346 3058 3357
rect 1894 3345 1900 3346
rect 1894 3341 1895 3345
rect 1899 3341 1900 3345
rect 1894 3340 1900 3341
rect 2046 3345 2052 3346
rect 2046 3341 2047 3345
rect 2051 3341 2052 3345
rect 2046 3340 2052 3341
rect 2206 3345 2212 3346
rect 2206 3341 2207 3345
rect 2211 3341 2212 3345
rect 2206 3340 2212 3341
rect 2366 3345 2372 3346
rect 2366 3341 2367 3345
rect 2371 3341 2372 3345
rect 2366 3340 2372 3341
rect 2534 3345 2540 3346
rect 2534 3341 2535 3345
rect 2539 3341 2540 3345
rect 2534 3340 2540 3341
rect 2702 3345 2708 3346
rect 2702 3341 2703 3345
rect 2707 3341 2708 3345
rect 2702 3340 2708 3341
rect 2878 3345 2884 3346
rect 2878 3341 2879 3345
rect 2883 3341 2884 3345
rect 2878 3340 2884 3341
rect 3054 3345 3060 3346
rect 3054 3341 3055 3345
rect 3059 3341 3060 3345
rect 3054 3340 3060 3341
rect 3576 3333 3578 3357
rect 110 3332 116 3333
rect 110 3328 111 3332
rect 115 3328 116 3332
rect 110 3327 116 3328
rect 1822 3332 1828 3333
rect 1822 3328 1823 3332
rect 1827 3328 1828 3332
rect 1822 3327 1828 3328
rect 1862 3332 1868 3333
rect 1862 3328 1863 3332
rect 1867 3328 1868 3332
rect 1862 3327 1868 3328
rect 3574 3332 3580 3333
rect 3574 3328 3575 3332
rect 3579 3328 3580 3332
rect 3574 3327 3580 3328
rect 110 3315 116 3316
rect 110 3311 111 3315
rect 115 3311 116 3315
rect 110 3310 116 3311
rect 1822 3315 1828 3316
rect 1822 3311 1823 3315
rect 1827 3311 1828 3315
rect 1822 3310 1828 3311
rect 1862 3315 1868 3316
rect 1862 3311 1863 3315
rect 1867 3311 1868 3315
rect 1862 3310 1868 3311
rect 3574 3315 3580 3316
rect 3574 3311 3575 3315
rect 3579 3311 3580 3315
rect 3574 3310 3580 3311
rect 112 3291 114 3310
rect 198 3305 204 3306
rect 198 3301 199 3305
rect 203 3301 204 3305
rect 198 3300 204 3301
rect 358 3305 364 3306
rect 358 3301 359 3305
rect 363 3301 364 3305
rect 358 3300 364 3301
rect 526 3305 532 3306
rect 526 3301 527 3305
rect 531 3301 532 3305
rect 526 3300 532 3301
rect 686 3305 692 3306
rect 686 3301 687 3305
rect 691 3301 692 3305
rect 686 3300 692 3301
rect 846 3305 852 3306
rect 846 3301 847 3305
rect 851 3301 852 3305
rect 846 3300 852 3301
rect 990 3305 996 3306
rect 990 3301 991 3305
rect 995 3301 996 3305
rect 990 3300 996 3301
rect 1134 3305 1140 3306
rect 1134 3301 1135 3305
rect 1139 3301 1140 3305
rect 1134 3300 1140 3301
rect 1270 3305 1276 3306
rect 1270 3301 1271 3305
rect 1275 3301 1276 3305
rect 1270 3300 1276 3301
rect 1406 3305 1412 3306
rect 1406 3301 1407 3305
rect 1411 3301 1412 3305
rect 1406 3300 1412 3301
rect 1550 3305 1556 3306
rect 1550 3301 1551 3305
rect 1555 3301 1556 3305
rect 1550 3300 1556 3301
rect 200 3291 202 3300
rect 360 3291 362 3300
rect 528 3291 530 3300
rect 688 3291 690 3300
rect 848 3291 850 3300
rect 992 3291 994 3300
rect 1136 3291 1138 3300
rect 1272 3291 1274 3300
rect 1408 3291 1410 3300
rect 1552 3291 1554 3300
rect 1824 3291 1826 3310
rect 1864 3291 1866 3310
rect 1886 3305 1892 3306
rect 1886 3301 1887 3305
rect 1891 3301 1892 3305
rect 1886 3300 1892 3301
rect 2038 3305 2044 3306
rect 2038 3301 2039 3305
rect 2043 3301 2044 3305
rect 2038 3300 2044 3301
rect 2198 3305 2204 3306
rect 2198 3301 2199 3305
rect 2203 3301 2204 3305
rect 2198 3300 2204 3301
rect 2358 3305 2364 3306
rect 2358 3301 2359 3305
rect 2363 3301 2364 3305
rect 2358 3300 2364 3301
rect 2526 3305 2532 3306
rect 2526 3301 2527 3305
rect 2531 3301 2532 3305
rect 2526 3300 2532 3301
rect 2694 3305 2700 3306
rect 2694 3301 2695 3305
rect 2699 3301 2700 3305
rect 2694 3300 2700 3301
rect 2870 3305 2876 3306
rect 2870 3301 2871 3305
rect 2875 3301 2876 3305
rect 2870 3300 2876 3301
rect 3046 3305 3052 3306
rect 3046 3301 3047 3305
rect 3051 3301 3052 3305
rect 3046 3300 3052 3301
rect 1888 3291 1890 3300
rect 2040 3291 2042 3300
rect 2200 3291 2202 3300
rect 2360 3291 2362 3300
rect 2528 3291 2530 3300
rect 2696 3291 2698 3300
rect 2872 3291 2874 3300
rect 3048 3291 3050 3300
rect 3576 3291 3578 3310
rect 111 3290 115 3291
rect 111 3285 115 3286
rect 199 3290 203 3291
rect 199 3285 203 3286
rect 255 3290 259 3291
rect 255 3285 259 3286
rect 359 3290 363 3291
rect 359 3285 363 3286
rect 375 3290 379 3291
rect 375 3285 379 3286
rect 511 3290 515 3291
rect 511 3285 515 3286
rect 527 3290 531 3291
rect 527 3285 531 3286
rect 663 3290 667 3291
rect 663 3285 667 3286
rect 687 3290 691 3291
rect 687 3285 691 3286
rect 823 3290 827 3291
rect 823 3285 827 3286
rect 847 3290 851 3291
rect 847 3285 851 3286
rect 991 3290 995 3291
rect 991 3285 995 3286
rect 1135 3290 1139 3291
rect 1135 3285 1139 3286
rect 1167 3290 1171 3291
rect 1167 3285 1171 3286
rect 1271 3290 1275 3291
rect 1271 3285 1275 3286
rect 1343 3290 1347 3291
rect 1343 3285 1347 3286
rect 1407 3290 1411 3291
rect 1407 3285 1411 3286
rect 1519 3290 1523 3291
rect 1519 3285 1523 3286
rect 1551 3290 1555 3291
rect 1551 3285 1555 3286
rect 1823 3290 1827 3291
rect 1823 3285 1827 3286
rect 1863 3290 1867 3291
rect 1863 3285 1867 3286
rect 1887 3290 1891 3291
rect 1887 3285 1891 3286
rect 2039 3290 2043 3291
rect 2039 3285 2043 3286
rect 2063 3290 2067 3291
rect 2063 3285 2067 3286
rect 2199 3290 2203 3291
rect 2199 3285 2203 3286
rect 2263 3290 2267 3291
rect 2263 3285 2267 3286
rect 2359 3290 2363 3291
rect 2359 3285 2363 3286
rect 2455 3290 2459 3291
rect 2455 3285 2459 3286
rect 2527 3290 2531 3291
rect 2527 3285 2531 3286
rect 2639 3290 2643 3291
rect 2639 3285 2643 3286
rect 2695 3290 2699 3291
rect 2695 3285 2699 3286
rect 2815 3290 2819 3291
rect 2815 3285 2819 3286
rect 2871 3290 2875 3291
rect 2871 3285 2875 3286
rect 2983 3290 2987 3291
rect 2983 3285 2987 3286
rect 3047 3290 3051 3291
rect 3047 3285 3051 3286
rect 3151 3290 3155 3291
rect 3151 3285 3155 3286
rect 3319 3290 3323 3291
rect 3319 3285 3323 3286
rect 3479 3290 3483 3291
rect 3479 3285 3483 3286
rect 3575 3290 3579 3291
rect 3575 3285 3579 3286
rect 112 3270 114 3285
rect 256 3280 258 3285
rect 376 3280 378 3285
rect 512 3280 514 3285
rect 664 3280 666 3285
rect 824 3280 826 3285
rect 992 3280 994 3285
rect 1168 3280 1170 3285
rect 1344 3280 1346 3285
rect 1520 3280 1522 3285
rect 254 3279 260 3280
rect 254 3275 255 3279
rect 259 3275 260 3279
rect 254 3274 260 3275
rect 374 3279 380 3280
rect 374 3275 375 3279
rect 379 3275 380 3279
rect 374 3274 380 3275
rect 510 3279 516 3280
rect 510 3275 511 3279
rect 515 3275 516 3279
rect 510 3274 516 3275
rect 662 3279 668 3280
rect 662 3275 663 3279
rect 667 3275 668 3279
rect 662 3274 668 3275
rect 822 3279 828 3280
rect 822 3275 823 3279
rect 827 3275 828 3279
rect 822 3274 828 3275
rect 990 3279 996 3280
rect 990 3275 991 3279
rect 995 3275 996 3279
rect 990 3274 996 3275
rect 1166 3279 1172 3280
rect 1166 3275 1167 3279
rect 1171 3275 1172 3279
rect 1166 3274 1172 3275
rect 1342 3279 1348 3280
rect 1342 3275 1343 3279
rect 1347 3275 1348 3279
rect 1342 3274 1348 3275
rect 1518 3279 1524 3280
rect 1518 3275 1519 3279
rect 1523 3275 1524 3279
rect 1518 3274 1524 3275
rect 1824 3270 1826 3285
rect 1864 3270 1866 3285
rect 1888 3280 1890 3285
rect 2064 3280 2066 3285
rect 2264 3280 2266 3285
rect 2456 3280 2458 3285
rect 2640 3280 2642 3285
rect 2816 3280 2818 3285
rect 2984 3280 2986 3285
rect 3152 3280 3154 3285
rect 3320 3280 3322 3285
rect 3480 3280 3482 3285
rect 1886 3279 1892 3280
rect 1886 3275 1887 3279
rect 1891 3275 1892 3279
rect 1886 3274 1892 3275
rect 2062 3279 2068 3280
rect 2062 3275 2063 3279
rect 2067 3275 2068 3279
rect 2062 3274 2068 3275
rect 2262 3279 2268 3280
rect 2262 3275 2263 3279
rect 2267 3275 2268 3279
rect 2262 3274 2268 3275
rect 2454 3279 2460 3280
rect 2454 3275 2455 3279
rect 2459 3275 2460 3279
rect 2454 3274 2460 3275
rect 2638 3279 2644 3280
rect 2638 3275 2639 3279
rect 2643 3275 2644 3279
rect 2638 3274 2644 3275
rect 2814 3279 2820 3280
rect 2814 3275 2815 3279
rect 2819 3275 2820 3279
rect 2814 3274 2820 3275
rect 2982 3279 2988 3280
rect 2982 3275 2983 3279
rect 2987 3275 2988 3279
rect 2982 3274 2988 3275
rect 3150 3279 3156 3280
rect 3150 3275 3151 3279
rect 3155 3275 3156 3279
rect 3150 3274 3156 3275
rect 3318 3279 3324 3280
rect 3318 3275 3319 3279
rect 3323 3275 3324 3279
rect 3318 3274 3324 3275
rect 3478 3279 3484 3280
rect 3478 3275 3479 3279
rect 3483 3275 3484 3279
rect 3478 3274 3484 3275
rect 3576 3270 3578 3285
rect 110 3269 116 3270
rect 110 3265 111 3269
rect 115 3265 116 3269
rect 110 3264 116 3265
rect 1822 3269 1828 3270
rect 1822 3265 1823 3269
rect 1827 3265 1828 3269
rect 1822 3264 1828 3265
rect 1862 3269 1868 3270
rect 1862 3265 1863 3269
rect 1867 3265 1868 3269
rect 1862 3264 1868 3265
rect 3574 3269 3580 3270
rect 3574 3265 3575 3269
rect 3579 3265 3580 3269
rect 3574 3264 3580 3265
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 110 3247 116 3248
rect 1822 3252 1828 3253
rect 1822 3248 1823 3252
rect 1827 3248 1828 3252
rect 1822 3247 1828 3248
rect 1862 3252 1868 3253
rect 1862 3248 1863 3252
rect 1867 3248 1868 3252
rect 1862 3247 1868 3248
rect 3574 3252 3580 3253
rect 3574 3248 3575 3252
rect 3579 3248 3580 3252
rect 3574 3247 3580 3248
rect 112 3219 114 3247
rect 262 3239 268 3240
rect 262 3235 263 3239
rect 267 3235 268 3239
rect 262 3234 268 3235
rect 382 3239 388 3240
rect 382 3235 383 3239
rect 387 3235 388 3239
rect 382 3234 388 3235
rect 518 3239 524 3240
rect 518 3235 519 3239
rect 523 3235 524 3239
rect 518 3234 524 3235
rect 670 3239 676 3240
rect 670 3235 671 3239
rect 675 3235 676 3239
rect 670 3234 676 3235
rect 830 3239 836 3240
rect 830 3235 831 3239
rect 835 3235 836 3239
rect 830 3234 836 3235
rect 998 3239 1004 3240
rect 998 3235 999 3239
rect 1003 3235 1004 3239
rect 998 3234 1004 3235
rect 1174 3239 1180 3240
rect 1174 3235 1175 3239
rect 1179 3235 1180 3239
rect 1174 3234 1180 3235
rect 1350 3239 1356 3240
rect 1350 3235 1351 3239
rect 1355 3235 1356 3239
rect 1350 3234 1356 3235
rect 1526 3239 1532 3240
rect 1526 3235 1527 3239
rect 1531 3235 1532 3239
rect 1526 3234 1532 3235
rect 264 3219 266 3234
rect 384 3219 386 3234
rect 520 3219 522 3234
rect 672 3219 674 3234
rect 832 3219 834 3234
rect 1000 3219 1002 3234
rect 1176 3219 1178 3234
rect 1352 3219 1354 3234
rect 1528 3219 1530 3234
rect 1824 3219 1826 3247
rect 1864 3223 1866 3247
rect 1894 3239 1900 3240
rect 1894 3235 1895 3239
rect 1899 3235 1900 3239
rect 1894 3234 1900 3235
rect 2070 3239 2076 3240
rect 2070 3235 2071 3239
rect 2075 3235 2076 3239
rect 2070 3234 2076 3235
rect 2270 3239 2276 3240
rect 2270 3235 2271 3239
rect 2275 3235 2276 3239
rect 2270 3234 2276 3235
rect 2462 3239 2468 3240
rect 2462 3235 2463 3239
rect 2467 3235 2468 3239
rect 2462 3234 2468 3235
rect 2646 3239 2652 3240
rect 2646 3235 2647 3239
rect 2651 3235 2652 3239
rect 2646 3234 2652 3235
rect 2822 3239 2828 3240
rect 2822 3235 2823 3239
rect 2827 3235 2828 3239
rect 2822 3234 2828 3235
rect 2990 3239 2996 3240
rect 2990 3235 2991 3239
rect 2995 3235 2996 3239
rect 2990 3234 2996 3235
rect 3158 3239 3164 3240
rect 3158 3235 3159 3239
rect 3163 3235 3164 3239
rect 3158 3234 3164 3235
rect 3326 3239 3332 3240
rect 3326 3235 3327 3239
rect 3331 3235 3332 3239
rect 3326 3234 3332 3235
rect 3486 3239 3492 3240
rect 3486 3235 3487 3239
rect 3491 3235 3492 3239
rect 3486 3234 3492 3235
rect 1896 3223 1898 3234
rect 2072 3223 2074 3234
rect 2272 3223 2274 3234
rect 2464 3223 2466 3234
rect 2648 3223 2650 3234
rect 2824 3223 2826 3234
rect 2992 3223 2994 3234
rect 3160 3223 3162 3234
rect 3328 3223 3330 3234
rect 3488 3223 3490 3234
rect 3576 3223 3578 3247
rect 1863 3222 1867 3223
rect 111 3218 115 3219
rect 111 3213 115 3214
rect 263 3218 267 3219
rect 263 3213 267 3214
rect 383 3218 387 3219
rect 383 3213 387 3214
rect 431 3218 435 3219
rect 431 3213 435 3214
rect 519 3218 523 3219
rect 519 3213 523 3214
rect 551 3218 555 3219
rect 551 3213 555 3214
rect 671 3218 675 3219
rect 671 3213 675 3214
rect 799 3218 803 3219
rect 799 3213 803 3214
rect 831 3218 835 3219
rect 831 3213 835 3214
rect 935 3218 939 3219
rect 935 3213 939 3214
rect 999 3218 1003 3219
rect 999 3213 1003 3214
rect 1079 3218 1083 3219
rect 1079 3213 1083 3214
rect 1175 3218 1179 3219
rect 1175 3213 1179 3214
rect 1231 3218 1235 3219
rect 1231 3213 1235 3214
rect 1351 3218 1355 3219
rect 1351 3213 1355 3214
rect 1383 3218 1387 3219
rect 1383 3213 1387 3214
rect 1527 3218 1531 3219
rect 1527 3213 1531 3214
rect 1535 3218 1539 3219
rect 1535 3213 1539 3214
rect 1823 3218 1827 3219
rect 1863 3217 1867 3218
rect 1895 3222 1899 3223
rect 1895 3217 1899 3218
rect 2071 3222 2075 3223
rect 2071 3217 2075 3218
rect 2087 3222 2091 3223
rect 2087 3217 2091 3218
rect 2271 3222 2275 3223
rect 2271 3217 2275 3218
rect 2303 3222 2307 3223
rect 2303 3217 2307 3218
rect 2463 3222 2467 3223
rect 2463 3217 2467 3218
rect 2511 3222 2515 3223
rect 2511 3217 2515 3218
rect 2647 3222 2651 3223
rect 2647 3217 2651 3218
rect 2703 3222 2707 3223
rect 2703 3217 2707 3218
rect 2823 3222 2827 3223
rect 2823 3217 2827 3218
rect 2879 3222 2883 3223
rect 2879 3217 2883 3218
rect 2991 3222 2995 3223
rect 2991 3217 2995 3218
rect 3039 3222 3043 3223
rect 3039 3217 3043 3218
rect 3159 3222 3163 3223
rect 3159 3217 3163 3218
rect 3199 3222 3203 3223
rect 3199 3217 3203 3218
rect 3327 3222 3331 3223
rect 3327 3217 3331 3218
rect 3351 3222 3355 3223
rect 3351 3217 3355 3218
rect 3487 3222 3491 3223
rect 3487 3217 3491 3218
rect 3575 3222 3579 3223
rect 3575 3217 3579 3218
rect 1823 3213 1827 3214
rect 112 3189 114 3213
rect 432 3202 434 3213
rect 552 3202 554 3213
rect 672 3202 674 3213
rect 800 3202 802 3213
rect 936 3202 938 3213
rect 1080 3202 1082 3213
rect 1232 3202 1234 3213
rect 1384 3202 1386 3213
rect 1536 3202 1538 3213
rect 430 3201 436 3202
rect 430 3197 431 3201
rect 435 3197 436 3201
rect 430 3196 436 3197
rect 550 3201 556 3202
rect 550 3197 551 3201
rect 555 3197 556 3201
rect 550 3196 556 3197
rect 670 3201 676 3202
rect 670 3197 671 3201
rect 675 3197 676 3201
rect 670 3196 676 3197
rect 798 3201 804 3202
rect 798 3197 799 3201
rect 803 3197 804 3201
rect 798 3196 804 3197
rect 934 3201 940 3202
rect 934 3197 935 3201
rect 939 3197 940 3201
rect 934 3196 940 3197
rect 1078 3201 1084 3202
rect 1078 3197 1079 3201
rect 1083 3197 1084 3201
rect 1078 3196 1084 3197
rect 1230 3201 1236 3202
rect 1230 3197 1231 3201
rect 1235 3197 1236 3201
rect 1230 3196 1236 3197
rect 1382 3201 1388 3202
rect 1382 3197 1383 3201
rect 1387 3197 1388 3201
rect 1382 3196 1388 3197
rect 1534 3201 1540 3202
rect 1534 3197 1535 3201
rect 1539 3197 1540 3201
rect 1534 3196 1540 3197
rect 1824 3189 1826 3213
rect 1864 3193 1866 3217
rect 1896 3206 1898 3217
rect 2088 3206 2090 3217
rect 2304 3206 2306 3217
rect 2512 3206 2514 3217
rect 2704 3206 2706 3217
rect 2880 3206 2882 3217
rect 3040 3206 3042 3217
rect 3200 3206 3202 3217
rect 3352 3206 3354 3217
rect 3488 3206 3490 3217
rect 1894 3205 1900 3206
rect 1894 3201 1895 3205
rect 1899 3201 1900 3205
rect 1894 3200 1900 3201
rect 2086 3205 2092 3206
rect 2086 3201 2087 3205
rect 2091 3201 2092 3205
rect 2086 3200 2092 3201
rect 2302 3205 2308 3206
rect 2302 3201 2303 3205
rect 2307 3201 2308 3205
rect 2302 3200 2308 3201
rect 2510 3205 2516 3206
rect 2510 3201 2511 3205
rect 2515 3201 2516 3205
rect 2510 3200 2516 3201
rect 2702 3205 2708 3206
rect 2702 3201 2703 3205
rect 2707 3201 2708 3205
rect 2702 3200 2708 3201
rect 2878 3205 2884 3206
rect 2878 3201 2879 3205
rect 2883 3201 2884 3205
rect 2878 3200 2884 3201
rect 3038 3205 3044 3206
rect 3038 3201 3039 3205
rect 3043 3201 3044 3205
rect 3038 3200 3044 3201
rect 3198 3205 3204 3206
rect 3198 3201 3199 3205
rect 3203 3201 3204 3205
rect 3198 3200 3204 3201
rect 3350 3205 3356 3206
rect 3350 3201 3351 3205
rect 3355 3201 3356 3205
rect 3350 3200 3356 3201
rect 3486 3205 3492 3206
rect 3486 3201 3487 3205
rect 3491 3201 3492 3205
rect 3486 3200 3492 3201
rect 3576 3193 3578 3217
rect 1862 3192 1868 3193
rect 110 3188 116 3189
rect 110 3184 111 3188
rect 115 3184 116 3188
rect 110 3183 116 3184
rect 1822 3188 1828 3189
rect 1822 3184 1823 3188
rect 1827 3184 1828 3188
rect 1862 3188 1863 3192
rect 1867 3188 1868 3192
rect 1862 3187 1868 3188
rect 3574 3192 3580 3193
rect 3574 3188 3575 3192
rect 3579 3188 3580 3192
rect 3574 3187 3580 3188
rect 1822 3183 1828 3184
rect 1862 3175 1868 3176
rect 110 3171 116 3172
rect 110 3167 111 3171
rect 115 3167 116 3171
rect 110 3166 116 3167
rect 1822 3171 1828 3172
rect 1822 3167 1823 3171
rect 1827 3167 1828 3171
rect 1862 3171 1863 3175
rect 1867 3171 1868 3175
rect 1862 3170 1868 3171
rect 3574 3175 3580 3176
rect 3574 3171 3575 3175
rect 3579 3171 3580 3175
rect 3574 3170 3580 3171
rect 1822 3166 1828 3167
rect 112 3147 114 3166
rect 422 3161 428 3162
rect 422 3157 423 3161
rect 427 3157 428 3161
rect 422 3156 428 3157
rect 542 3161 548 3162
rect 542 3157 543 3161
rect 547 3157 548 3161
rect 542 3156 548 3157
rect 662 3161 668 3162
rect 662 3157 663 3161
rect 667 3157 668 3161
rect 662 3156 668 3157
rect 790 3161 796 3162
rect 790 3157 791 3161
rect 795 3157 796 3161
rect 790 3156 796 3157
rect 926 3161 932 3162
rect 926 3157 927 3161
rect 931 3157 932 3161
rect 926 3156 932 3157
rect 1070 3161 1076 3162
rect 1070 3157 1071 3161
rect 1075 3157 1076 3161
rect 1070 3156 1076 3157
rect 1222 3161 1228 3162
rect 1222 3157 1223 3161
rect 1227 3157 1228 3161
rect 1222 3156 1228 3157
rect 1374 3161 1380 3162
rect 1374 3157 1375 3161
rect 1379 3157 1380 3161
rect 1374 3156 1380 3157
rect 1526 3161 1532 3162
rect 1526 3157 1527 3161
rect 1531 3157 1532 3161
rect 1526 3156 1532 3157
rect 424 3147 426 3156
rect 544 3147 546 3156
rect 664 3147 666 3156
rect 792 3147 794 3156
rect 928 3147 930 3156
rect 1072 3147 1074 3156
rect 1224 3147 1226 3156
rect 1376 3147 1378 3156
rect 1528 3147 1530 3156
rect 1824 3147 1826 3166
rect 1864 3151 1866 3170
rect 1886 3165 1892 3166
rect 1886 3161 1887 3165
rect 1891 3161 1892 3165
rect 1886 3160 1892 3161
rect 2078 3165 2084 3166
rect 2078 3161 2079 3165
rect 2083 3161 2084 3165
rect 2078 3160 2084 3161
rect 2294 3165 2300 3166
rect 2294 3161 2295 3165
rect 2299 3161 2300 3165
rect 2294 3160 2300 3161
rect 2502 3165 2508 3166
rect 2502 3161 2503 3165
rect 2507 3161 2508 3165
rect 2502 3160 2508 3161
rect 2694 3165 2700 3166
rect 2694 3161 2695 3165
rect 2699 3161 2700 3165
rect 2694 3160 2700 3161
rect 2870 3165 2876 3166
rect 2870 3161 2871 3165
rect 2875 3161 2876 3165
rect 2870 3160 2876 3161
rect 3030 3165 3036 3166
rect 3030 3161 3031 3165
rect 3035 3161 3036 3165
rect 3030 3160 3036 3161
rect 3190 3165 3196 3166
rect 3190 3161 3191 3165
rect 3195 3161 3196 3165
rect 3190 3160 3196 3161
rect 3342 3165 3348 3166
rect 3342 3161 3343 3165
rect 3347 3161 3348 3165
rect 3342 3160 3348 3161
rect 3478 3165 3484 3166
rect 3478 3161 3479 3165
rect 3483 3161 3484 3165
rect 3478 3160 3484 3161
rect 1888 3151 1890 3160
rect 2080 3151 2082 3160
rect 2296 3151 2298 3160
rect 2504 3151 2506 3160
rect 2696 3151 2698 3160
rect 2872 3151 2874 3160
rect 3032 3151 3034 3160
rect 3192 3151 3194 3160
rect 3344 3151 3346 3160
rect 3480 3151 3482 3160
rect 3576 3151 3578 3170
rect 1863 3150 1867 3151
rect 111 3146 115 3147
rect 111 3141 115 3142
rect 423 3146 427 3147
rect 423 3141 427 3142
rect 463 3146 467 3147
rect 463 3141 467 3142
rect 543 3146 547 3147
rect 543 3141 547 3142
rect 551 3146 555 3147
rect 551 3141 555 3142
rect 639 3146 643 3147
rect 639 3141 643 3142
rect 663 3146 667 3147
rect 663 3141 667 3142
rect 735 3146 739 3147
rect 735 3141 739 3142
rect 791 3146 795 3147
rect 791 3141 795 3142
rect 847 3146 851 3147
rect 847 3141 851 3142
rect 927 3146 931 3147
rect 927 3141 931 3142
rect 967 3146 971 3147
rect 967 3141 971 3142
rect 1071 3146 1075 3147
rect 1071 3141 1075 3142
rect 1095 3146 1099 3147
rect 1095 3141 1099 3142
rect 1223 3146 1227 3147
rect 1223 3141 1227 3142
rect 1231 3146 1235 3147
rect 1231 3141 1235 3142
rect 1375 3146 1379 3147
rect 1375 3141 1379 3142
rect 1519 3146 1523 3147
rect 1519 3141 1523 3142
rect 1527 3146 1531 3147
rect 1527 3141 1531 3142
rect 1823 3146 1827 3147
rect 1863 3145 1867 3146
rect 1887 3150 1891 3151
rect 1887 3145 1891 3146
rect 2079 3150 2083 3151
rect 2079 3145 2083 3146
rect 2295 3150 2299 3151
rect 2295 3145 2299 3146
rect 2503 3150 2507 3151
rect 2503 3145 2507 3146
rect 2695 3150 2699 3151
rect 2695 3145 2699 3146
rect 2871 3150 2875 3151
rect 2871 3145 2875 3146
rect 3031 3150 3035 3151
rect 3031 3145 3035 3146
rect 3039 3150 3043 3151
rect 3039 3145 3043 3146
rect 3191 3150 3195 3151
rect 3191 3145 3195 3146
rect 3343 3150 3347 3151
rect 3343 3145 3347 3146
rect 3479 3150 3483 3151
rect 3479 3145 3483 3146
rect 3575 3150 3579 3151
rect 3575 3145 3579 3146
rect 1823 3141 1827 3142
rect 112 3126 114 3141
rect 464 3136 466 3141
rect 552 3136 554 3141
rect 640 3136 642 3141
rect 736 3136 738 3141
rect 848 3136 850 3141
rect 968 3136 970 3141
rect 1096 3136 1098 3141
rect 1232 3136 1234 3141
rect 1376 3136 1378 3141
rect 1520 3136 1522 3141
rect 462 3135 468 3136
rect 462 3131 463 3135
rect 467 3131 468 3135
rect 462 3130 468 3131
rect 550 3135 556 3136
rect 550 3131 551 3135
rect 555 3131 556 3135
rect 550 3130 556 3131
rect 638 3135 644 3136
rect 638 3131 639 3135
rect 643 3131 644 3135
rect 638 3130 644 3131
rect 734 3135 740 3136
rect 734 3131 735 3135
rect 739 3131 740 3135
rect 734 3130 740 3131
rect 846 3135 852 3136
rect 846 3131 847 3135
rect 851 3131 852 3135
rect 846 3130 852 3131
rect 966 3135 972 3136
rect 966 3131 967 3135
rect 971 3131 972 3135
rect 966 3130 972 3131
rect 1094 3135 1100 3136
rect 1094 3131 1095 3135
rect 1099 3131 1100 3135
rect 1094 3130 1100 3131
rect 1230 3135 1236 3136
rect 1230 3131 1231 3135
rect 1235 3131 1236 3135
rect 1230 3130 1236 3131
rect 1374 3135 1380 3136
rect 1374 3131 1375 3135
rect 1379 3131 1380 3135
rect 1374 3130 1380 3131
rect 1518 3135 1524 3136
rect 1518 3131 1519 3135
rect 1523 3131 1524 3135
rect 1518 3130 1524 3131
rect 1824 3126 1826 3141
rect 1864 3130 1866 3145
rect 1888 3140 1890 3145
rect 2080 3140 2082 3145
rect 2296 3140 2298 3145
rect 2504 3140 2506 3145
rect 2696 3140 2698 3145
rect 2872 3140 2874 3145
rect 3040 3140 3042 3145
rect 3192 3140 3194 3145
rect 3344 3140 3346 3145
rect 3480 3140 3482 3145
rect 1886 3139 1892 3140
rect 1886 3135 1887 3139
rect 1891 3135 1892 3139
rect 1886 3134 1892 3135
rect 2078 3139 2084 3140
rect 2078 3135 2079 3139
rect 2083 3135 2084 3139
rect 2078 3134 2084 3135
rect 2294 3139 2300 3140
rect 2294 3135 2295 3139
rect 2299 3135 2300 3139
rect 2294 3134 2300 3135
rect 2502 3139 2508 3140
rect 2502 3135 2503 3139
rect 2507 3135 2508 3139
rect 2502 3134 2508 3135
rect 2694 3139 2700 3140
rect 2694 3135 2695 3139
rect 2699 3135 2700 3139
rect 2694 3134 2700 3135
rect 2870 3139 2876 3140
rect 2870 3135 2871 3139
rect 2875 3135 2876 3139
rect 2870 3134 2876 3135
rect 3038 3139 3044 3140
rect 3038 3135 3039 3139
rect 3043 3135 3044 3139
rect 3038 3134 3044 3135
rect 3190 3139 3196 3140
rect 3190 3135 3191 3139
rect 3195 3135 3196 3139
rect 3190 3134 3196 3135
rect 3342 3139 3348 3140
rect 3342 3135 3343 3139
rect 3347 3135 3348 3139
rect 3342 3134 3348 3135
rect 3478 3139 3484 3140
rect 3478 3135 3479 3139
rect 3483 3135 3484 3139
rect 3478 3134 3484 3135
rect 3576 3130 3578 3145
rect 1862 3129 1868 3130
rect 110 3125 116 3126
rect 110 3121 111 3125
rect 115 3121 116 3125
rect 110 3120 116 3121
rect 1822 3125 1828 3126
rect 1822 3121 1823 3125
rect 1827 3121 1828 3125
rect 1862 3125 1863 3129
rect 1867 3125 1868 3129
rect 1862 3124 1868 3125
rect 3574 3129 3580 3130
rect 3574 3125 3575 3129
rect 3579 3125 3580 3129
rect 3574 3124 3580 3125
rect 1822 3120 1828 3121
rect 1862 3112 1868 3113
rect 110 3108 116 3109
rect 110 3104 111 3108
rect 115 3104 116 3108
rect 110 3103 116 3104
rect 1822 3108 1828 3109
rect 1822 3104 1823 3108
rect 1827 3104 1828 3108
rect 1862 3108 1863 3112
rect 1867 3108 1868 3112
rect 1862 3107 1868 3108
rect 3574 3112 3580 3113
rect 3574 3108 3575 3112
rect 3579 3108 3580 3112
rect 3574 3107 3580 3108
rect 1822 3103 1828 3104
rect 112 3071 114 3103
rect 470 3095 476 3096
rect 470 3091 471 3095
rect 475 3091 476 3095
rect 470 3090 476 3091
rect 558 3095 564 3096
rect 558 3091 559 3095
rect 563 3091 564 3095
rect 558 3090 564 3091
rect 646 3095 652 3096
rect 646 3091 647 3095
rect 651 3091 652 3095
rect 646 3090 652 3091
rect 742 3095 748 3096
rect 742 3091 743 3095
rect 747 3091 748 3095
rect 742 3090 748 3091
rect 854 3095 860 3096
rect 854 3091 855 3095
rect 859 3091 860 3095
rect 854 3090 860 3091
rect 974 3095 980 3096
rect 974 3091 975 3095
rect 979 3091 980 3095
rect 974 3090 980 3091
rect 1102 3095 1108 3096
rect 1102 3091 1103 3095
rect 1107 3091 1108 3095
rect 1102 3090 1108 3091
rect 1238 3095 1244 3096
rect 1238 3091 1239 3095
rect 1243 3091 1244 3095
rect 1238 3090 1244 3091
rect 1382 3095 1388 3096
rect 1382 3091 1383 3095
rect 1387 3091 1388 3095
rect 1382 3090 1388 3091
rect 1526 3095 1532 3096
rect 1526 3091 1527 3095
rect 1531 3091 1532 3095
rect 1526 3090 1532 3091
rect 472 3071 474 3090
rect 560 3071 562 3090
rect 648 3071 650 3090
rect 744 3071 746 3090
rect 856 3071 858 3090
rect 976 3071 978 3090
rect 1104 3071 1106 3090
rect 1240 3071 1242 3090
rect 1384 3071 1386 3090
rect 1528 3071 1530 3090
rect 1824 3071 1826 3103
rect 1864 3071 1866 3107
rect 1894 3099 1900 3100
rect 1894 3095 1895 3099
rect 1899 3095 1900 3099
rect 1894 3094 1900 3095
rect 2086 3099 2092 3100
rect 2086 3095 2087 3099
rect 2091 3095 2092 3099
rect 2086 3094 2092 3095
rect 2302 3099 2308 3100
rect 2302 3095 2303 3099
rect 2307 3095 2308 3099
rect 2302 3094 2308 3095
rect 2510 3099 2516 3100
rect 2510 3095 2511 3099
rect 2515 3095 2516 3099
rect 2510 3094 2516 3095
rect 2702 3099 2708 3100
rect 2702 3095 2703 3099
rect 2707 3095 2708 3099
rect 2702 3094 2708 3095
rect 2878 3099 2884 3100
rect 2878 3095 2879 3099
rect 2883 3095 2884 3099
rect 2878 3094 2884 3095
rect 3046 3099 3052 3100
rect 3046 3095 3047 3099
rect 3051 3095 3052 3099
rect 3046 3094 3052 3095
rect 3198 3099 3204 3100
rect 3198 3095 3199 3099
rect 3203 3095 3204 3099
rect 3198 3094 3204 3095
rect 3350 3099 3356 3100
rect 3350 3095 3351 3099
rect 3355 3095 3356 3099
rect 3350 3094 3356 3095
rect 3486 3099 3492 3100
rect 3486 3095 3487 3099
rect 3491 3095 3492 3099
rect 3486 3094 3492 3095
rect 1896 3071 1898 3094
rect 2088 3071 2090 3094
rect 2304 3071 2306 3094
rect 2512 3071 2514 3094
rect 2704 3071 2706 3094
rect 2880 3071 2882 3094
rect 3048 3071 3050 3094
rect 3200 3071 3202 3094
rect 3352 3071 3354 3094
rect 3488 3071 3490 3094
rect 3576 3071 3578 3107
rect 111 3070 115 3071
rect 111 3065 115 3066
rect 151 3070 155 3071
rect 151 3065 155 3066
rect 239 3070 243 3071
rect 239 3065 243 3066
rect 327 3070 331 3071
rect 327 3065 331 3066
rect 415 3070 419 3071
rect 415 3065 419 3066
rect 471 3070 475 3071
rect 471 3065 475 3066
rect 503 3070 507 3071
rect 503 3065 507 3066
rect 559 3070 563 3071
rect 559 3065 563 3066
rect 591 3070 595 3071
rect 591 3065 595 3066
rect 647 3070 651 3071
rect 647 3065 651 3066
rect 679 3070 683 3071
rect 679 3065 683 3066
rect 743 3070 747 3071
rect 743 3065 747 3066
rect 767 3070 771 3071
rect 767 3065 771 3066
rect 855 3070 859 3071
rect 855 3065 859 3066
rect 943 3070 947 3071
rect 943 3065 947 3066
rect 975 3070 979 3071
rect 975 3065 979 3066
rect 1031 3070 1035 3071
rect 1031 3065 1035 3066
rect 1103 3070 1107 3071
rect 1103 3065 1107 3066
rect 1119 3070 1123 3071
rect 1119 3065 1123 3066
rect 1207 3070 1211 3071
rect 1207 3065 1211 3066
rect 1239 3070 1243 3071
rect 1239 3065 1243 3066
rect 1295 3070 1299 3071
rect 1295 3065 1299 3066
rect 1383 3070 1387 3071
rect 1383 3065 1387 3066
rect 1471 3070 1475 3071
rect 1471 3065 1475 3066
rect 1527 3070 1531 3071
rect 1527 3065 1531 3066
rect 1559 3070 1563 3071
rect 1559 3065 1563 3066
rect 1647 3070 1651 3071
rect 1647 3065 1651 3066
rect 1735 3070 1739 3071
rect 1735 3065 1739 3066
rect 1823 3070 1827 3071
rect 1823 3065 1827 3066
rect 1863 3070 1867 3071
rect 1863 3065 1867 3066
rect 1895 3070 1899 3071
rect 1895 3065 1899 3066
rect 2087 3070 2091 3071
rect 2087 3065 2091 3066
rect 2255 3070 2259 3071
rect 2255 3065 2259 3066
rect 2303 3070 2307 3071
rect 2303 3065 2307 3066
rect 2423 3070 2427 3071
rect 2423 3065 2427 3066
rect 2511 3070 2515 3071
rect 2511 3065 2515 3066
rect 2591 3070 2595 3071
rect 2591 3065 2595 3066
rect 2703 3070 2707 3071
rect 2703 3065 2707 3066
rect 2751 3070 2755 3071
rect 2751 3065 2755 3066
rect 2879 3070 2883 3071
rect 2879 3065 2883 3066
rect 2919 3070 2923 3071
rect 2919 3065 2923 3066
rect 3047 3070 3051 3071
rect 3047 3065 3051 3066
rect 3087 3070 3091 3071
rect 3087 3065 3091 3066
rect 3199 3070 3203 3071
rect 3199 3065 3203 3066
rect 3351 3070 3355 3071
rect 3351 3065 3355 3066
rect 3487 3070 3491 3071
rect 3487 3065 3491 3066
rect 3575 3070 3579 3071
rect 3575 3065 3579 3066
rect 112 3041 114 3065
rect 152 3054 154 3065
rect 240 3054 242 3065
rect 328 3054 330 3065
rect 416 3054 418 3065
rect 504 3054 506 3065
rect 592 3054 594 3065
rect 680 3054 682 3065
rect 768 3054 770 3065
rect 856 3054 858 3065
rect 944 3054 946 3065
rect 1032 3054 1034 3065
rect 1120 3054 1122 3065
rect 1208 3054 1210 3065
rect 1296 3054 1298 3065
rect 1384 3054 1386 3065
rect 1472 3054 1474 3065
rect 1560 3054 1562 3065
rect 1648 3054 1650 3065
rect 1736 3054 1738 3065
rect 150 3053 156 3054
rect 150 3049 151 3053
rect 155 3049 156 3053
rect 150 3048 156 3049
rect 238 3053 244 3054
rect 238 3049 239 3053
rect 243 3049 244 3053
rect 238 3048 244 3049
rect 326 3053 332 3054
rect 326 3049 327 3053
rect 331 3049 332 3053
rect 326 3048 332 3049
rect 414 3053 420 3054
rect 414 3049 415 3053
rect 419 3049 420 3053
rect 414 3048 420 3049
rect 502 3053 508 3054
rect 502 3049 503 3053
rect 507 3049 508 3053
rect 502 3048 508 3049
rect 590 3053 596 3054
rect 590 3049 591 3053
rect 595 3049 596 3053
rect 590 3048 596 3049
rect 678 3053 684 3054
rect 678 3049 679 3053
rect 683 3049 684 3053
rect 678 3048 684 3049
rect 766 3053 772 3054
rect 766 3049 767 3053
rect 771 3049 772 3053
rect 766 3048 772 3049
rect 854 3053 860 3054
rect 854 3049 855 3053
rect 859 3049 860 3053
rect 854 3048 860 3049
rect 942 3053 948 3054
rect 942 3049 943 3053
rect 947 3049 948 3053
rect 942 3048 948 3049
rect 1030 3053 1036 3054
rect 1030 3049 1031 3053
rect 1035 3049 1036 3053
rect 1030 3048 1036 3049
rect 1118 3053 1124 3054
rect 1118 3049 1119 3053
rect 1123 3049 1124 3053
rect 1118 3048 1124 3049
rect 1206 3053 1212 3054
rect 1206 3049 1207 3053
rect 1211 3049 1212 3053
rect 1206 3048 1212 3049
rect 1294 3053 1300 3054
rect 1294 3049 1295 3053
rect 1299 3049 1300 3053
rect 1294 3048 1300 3049
rect 1382 3053 1388 3054
rect 1382 3049 1383 3053
rect 1387 3049 1388 3053
rect 1382 3048 1388 3049
rect 1470 3053 1476 3054
rect 1470 3049 1471 3053
rect 1475 3049 1476 3053
rect 1470 3048 1476 3049
rect 1558 3053 1564 3054
rect 1558 3049 1559 3053
rect 1563 3049 1564 3053
rect 1558 3048 1564 3049
rect 1646 3053 1652 3054
rect 1646 3049 1647 3053
rect 1651 3049 1652 3053
rect 1646 3048 1652 3049
rect 1734 3053 1740 3054
rect 1734 3049 1735 3053
rect 1739 3049 1740 3053
rect 1734 3048 1740 3049
rect 1824 3041 1826 3065
rect 1864 3041 1866 3065
rect 2256 3054 2258 3065
rect 2424 3054 2426 3065
rect 2592 3054 2594 3065
rect 2752 3054 2754 3065
rect 2920 3054 2922 3065
rect 3088 3054 3090 3065
rect 2254 3053 2260 3054
rect 2254 3049 2255 3053
rect 2259 3049 2260 3053
rect 2254 3048 2260 3049
rect 2422 3053 2428 3054
rect 2422 3049 2423 3053
rect 2427 3049 2428 3053
rect 2422 3048 2428 3049
rect 2590 3053 2596 3054
rect 2590 3049 2591 3053
rect 2595 3049 2596 3053
rect 2590 3048 2596 3049
rect 2750 3053 2756 3054
rect 2750 3049 2751 3053
rect 2755 3049 2756 3053
rect 2750 3048 2756 3049
rect 2918 3053 2924 3054
rect 2918 3049 2919 3053
rect 2923 3049 2924 3053
rect 2918 3048 2924 3049
rect 3086 3053 3092 3054
rect 3086 3049 3087 3053
rect 3091 3049 3092 3053
rect 3086 3048 3092 3049
rect 3576 3041 3578 3065
rect 110 3040 116 3041
rect 110 3036 111 3040
rect 115 3036 116 3040
rect 110 3035 116 3036
rect 1822 3040 1828 3041
rect 1822 3036 1823 3040
rect 1827 3036 1828 3040
rect 1822 3035 1828 3036
rect 1862 3040 1868 3041
rect 1862 3036 1863 3040
rect 1867 3036 1868 3040
rect 1862 3035 1868 3036
rect 3574 3040 3580 3041
rect 3574 3036 3575 3040
rect 3579 3036 3580 3040
rect 3574 3035 3580 3036
rect 110 3023 116 3024
rect 110 3019 111 3023
rect 115 3019 116 3023
rect 110 3018 116 3019
rect 1822 3023 1828 3024
rect 1822 3019 1823 3023
rect 1827 3019 1828 3023
rect 1822 3018 1828 3019
rect 1862 3023 1868 3024
rect 1862 3019 1863 3023
rect 1867 3019 1868 3023
rect 1862 3018 1868 3019
rect 3574 3023 3580 3024
rect 3574 3019 3575 3023
rect 3579 3019 3580 3023
rect 3574 3018 3580 3019
rect 112 2995 114 3018
rect 142 3013 148 3014
rect 142 3009 143 3013
rect 147 3009 148 3013
rect 142 3008 148 3009
rect 230 3013 236 3014
rect 230 3009 231 3013
rect 235 3009 236 3013
rect 230 3008 236 3009
rect 318 3013 324 3014
rect 318 3009 319 3013
rect 323 3009 324 3013
rect 318 3008 324 3009
rect 406 3013 412 3014
rect 406 3009 407 3013
rect 411 3009 412 3013
rect 406 3008 412 3009
rect 494 3013 500 3014
rect 494 3009 495 3013
rect 499 3009 500 3013
rect 494 3008 500 3009
rect 582 3013 588 3014
rect 582 3009 583 3013
rect 587 3009 588 3013
rect 582 3008 588 3009
rect 670 3013 676 3014
rect 670 3009 671 3013
rect 675 3009 676 3013
rect 670 3008 676 3009
rect 758 3013 764 3014
rect 758 3009 759 3013
rect 763 3009 764 3013
rect 758 3008 764 3009
rect 846 3013 852 3014
rect 846 3009 847 3013
rect 851 3009 852 3013
rect 846 3008 852 3009
rect 934 3013 940 3014
rect 934 3009 935 3013
rect 939 3009 940 3013
rect 934 3008 940 3009
rect 1022 3013 1028 3014
rect 1022 3009 1023 3013
rect 1027 3009 1028 3013
rect 1022 3008 1028 3009
rect 1110 3013 1116 3014
rect 1110 3009 1111 3013
rect 1115 3009 1116 3013
rect 1110 3008 1116 3009
rect 1198 3013 1204 3014
rect 1198 3009 1199 3013
rect 1203 3009 1204 3013
rect 1198 3008 1204 3009
rect 1286 3013 1292 3014
rect 1286 3009 1287 3013
rect 1291 3009 1292 3013
rect 1286 3008 1292 3009
rect 1374 3013 1380 3014
rect 1374 3009 1375 3013
rect 1379 3009 1380 3013
rect 1374 3008 1380 3009
rect 1462 3013 1468 3014
rect 1462 3009 1463 3013
rect 1467 3009 1468 3013
rect 1462 3008 1468 3009
rect 1550 3013 1556 3014
rect 1550 3009 1551 3013
rect 1555 3009 1556 3013
rect 1550 3008 1556 3009
rect 1638 3013 1644 3014
rect 1638 3009 1639 3013
rect 1643 3009 1644 3013
rect 1638 3008 1644 3009
rect 1726 3013 1732 3014
rect 1726 3009 1727 3013
rect 1731 3009 1732 3013
rect 1726 3008 1732 3009
rect 144 2995 146 3008
rect 232 2995 234 3008
rect 320 2995 322 3008
rect 408 2995 410 3008
rect 496 2995 498 3008
rect 584 2995 586 3008
rect 672 2995 674 3008
rect 760 2995 762 3008
rect 848 2995 850 3008
rect 936 2995 938 3008
rect 1024 2995 1026 3008
rect 1112 2995 1114 3008
rect 1200 2995 1202 3008
rect 1288 2995 1290 3008
rect 1376 2995 1378 3008
rect 1464 2995 1466 3008
rect 1552 2995 1554 3008
rect 1640 2995 1642 3008
rect 1728 2995 1730 3008
rect 1824 2995 1826 3018
rect 1864 2999 1866 3018
rect 2246 3013 2252 3014
rect 2246 3009 2247 3013
rect 2251 3009 2252 3013
rect 2246 3008 2252 3009
rect 2414 3013 2420 3014
rect 2414 3009 2415 3013
rect 2419 3009 2420 3013
rect 2414 3008 2420 3009
rect 2582 3013 2588 3014
rect 2582 3009 2583 3013
rect 2587 3009 2588 3013
rect 2582 3008 2588 3009
rect 2742 3013 2748 3014
rect 2742 3009 2743 3013
rect 2747 3009 2748 3013
rect 2742 3008 2748 3009
rect 2910 3013 2916 3014
rect 2910 3009 2911 3013
rect 2915 3009 2916 3013
rect 2910 3008 2916 3009
rect 3078 3013 3084 3014
rect 3078 3009 3079 3013
rect 3083 3009 3084 3013
rect 3078 3008 3084 3009
rect 2248 2999 2250 3008
rect 2416 2999 2418 3008
rect 2584 2999 2586 3008
rect 2744 2999 2746 3008
rect 2912 2999 2914 3008
rect 3080 2999 3082 3008
rect 3576 2999 3578 3018
rect 1863 2998 1867 2999
rect 111 2994 115 2995
rect 111 2989 115 2990
rect 143 2994 147 2995
rect 143 2989 147 2990
rect 231 2994 235 2995
rect 231 2989 235 2990
rect 319 2994 323 2995
rect 319 2989 323 2990
rect 407 2994 411 2995
rect 407 2989 411 2990
rect 495 2994 499 2995
rect 495 2989 499 2990
rect 583 2994 587 2995
rect 583 2989 587 2990
rect 671 2994 675 2995
rect 671 2989 675 2990
rect 759 2994 763 2995
rect 759 2989 763 2990
rect 847 2994 851 2995
rect 847 2989 851 2990
rect 935 2994 939 2995
rect 935 2989 939 2990
rect 1023 2994 1027 2995
rect 1023 2989 1027 2990
rect 1111 2994 1115 2995
rect 1111 2989 1115 2990
rect 1199 2994 1203 2995
rect 1199 2989 1203 2990
rect 1287 2994 1291 2995
rect 1287 2989 1291 2990
rect 1375 2994 1379 2995
rect 1375 2989 1379 2990
rect 1407 2994 1411 2995
rect 1407 2989 1411 2990
rect 1463 2994 1467 2995
rect 1463 2989 1467 2990
rect 1519 2994 1523 2995
rect 1519 2989 1523 2990
rect 1551 2994 1555 2995
rect 1551 2989 1555 2990
rect 1631 2994 1635 2995
rect 1631 2989 1635 2990
rect 1639 2994 1643 2995
rect 1639 2989 1643 2990
rect 1727 2994 1731 2995
rect 1727 2989 1731 2990
rect 1823 2994 1827 2995
rect 1863 2993 1867 2994
rect 2239 2998 2243 2999
rect 2239 2993 2243 2994
rect 2247 2998 2251 2999
rect 2247 2993 2251 2994
rect 2415 2998 2419 2999
rect 2415 2993 2419 2994
rect 2463 2998 2467 2999
rect 2463 2993 2467 2994
rect 2583 2998 2587 2999
rect 2583 2993 2587 2994
rect 2671 2998 2675 2999
rect 2671 2993 2675 2994
rect 2743 2998 2747 2999
rect 2743 2993 2747 2994
rect 2863 2998 2867 2999
rect 2863 2993 2867 2994
rect 2911 2998 2915 2999
rect 2911 2993 2915 2994
rect 3031 2998 3035 2999
rect 3031 2993 3035 2994
rect 3079 2998 3083 2999
rect 3079 2993 3083 2994
rect 3191 2998 3195 2999
rect 3191 2993 3195 2994
rect 3343 2998 3347 2999
rect 3343 2993 3347 2994
rect 3479 2998 3483 2999
rect 3479 2993 3483 2994
rect 3575 2998 3579 2999
rect 3575 2993 3579 2994
rect 1823 2989 1827 2990
rect 112 2974 114 2989
rect 1408 2984 1410 2989
rect 1520 2984 1522 2989
rect 1632 2984 1634 2989
rect 1728 2984 1730 2989
rect 1406 2983 1412 2984
rect 1406 2979 1407 2983
rect 1411 2979 1412 2983
rect 1406 2978 1412 2979
rect 1518 2983 1524 2984
rect 1518 2979 1519 2983
rect 1523 2979 1524 2983
rect 1518 2978 1524 2979
rect 1630 2983 1636 2984
rect 1630 2979 1631 2983
rect 1635 2979 1636 2983
rect 1630 2978 1636 2979
rect 1726 2983 1732 2984
rect 1726 2979 1727 2983
rect 1731 2979 1732 2983
rect 1726 2978 1732 2979
rect 1824 2974 1826 2989
rect 1864 2978 1866 2993
rect 2240 2988 2242 2993
rect 2464 2988 2466 2993
rect 2672 2988 2674 2993
rect 2864 2988 2866 2993
rect 3032 2988 3034 2993
rect 3192 2988 3194 2993
rect 3344 2988 3346 2993
rect 3480 2988 3482 2993
rect 2238 2987 2244 2988
rect 2238 2983 2239 2987
rect 2243 2983 2244 2987
rect 2238 2982 2244 2983
rect 2462 2987 2468 2988
rect 2462 2983 2463 2987
rect 2467 2983 2468 2987
rect 2462 2982 2468 2983
rect 2670 2987 2676 2988
rect 2670 2983 2671 2987
rect 2675 2983 2676 2987
rect 2670 2982 2676 2983
rect 2862 2987 2868 2988
rect 2862 2983 2863 2987
rect 2867 2983 2868 2987
rect 2862 2982 2868 2983
rect 3030 2987 3036 2988
rect 3030 2983 3031 2987
rect 3035 2983 3036 2987
rect 3030 2982 3036 2983
rect 3190 2987 3196 2988
rect 3190 2983 3191 2987
rect 3195 2983 3196 2987
rect 3190 2982 3196 2983
rect 3342 2987 3348 2988
rect 3342 2983 3343 2987
rect 3347 2983 3348 2987
rect 3342 2982 3348 2983
rect 3478 2987 3484 2988
rect 3478 2983 3479 2987
rect 3483 2983 3484 2987
rect 3478 2982 3484 2983
rect 3576 2978 3578 2993
rect 1862 2977 1868 2978
rect 110 2973 116 2974
rect 110 2969 111 2973
rect 115 2969 116 2973
rect 110 2968 116 2969
rect 1822 2973 1828 2974
rect 1822 2969 1823 2973
rect 1827 2969 1828 2973
rect 1862 2973 1863 2977
rect 1867 2973 1868 2977
rect 1862 2972 1868 2973
rect 3574 2977 3580 2978
rect 3574 2973 3575 2977
rect 3579 2973 3580 2977
rect 3574 2972 3580 2973
rect 1822 2968 1828 2969
rect 1862 2960 1868 2961
rect 110 2956 116 2957
rect 110 2952 111 2956
rect 115 2952 116 2956
rect 110 2951 116 2952
rect 1822 2956 1828 2957
rect 1822 2952 1823 2956
rect 1827 2952 1828 2956
rect 1862 2956 1863 2960
rect 1867 2956 1868 2960
rect 1862 2955 1868 2956
rect 3574 2960 3580 2961
rect 3574 2956 3575 2960
rect 3579 2956 3580 2960
rect 3574 2955 3580 2956
rect 1822 2951 1828 2952
rect 112 2927 114 2951
rect 1414 2943 1420 2944
rect 1414 2939 1415 2943
rect 1419 2939 1420 2943
rect 1414 2938 1420 2939
rect 1526 2943 1532 2944
rect 1526 2939 1527 2943
rect 1531 2939 1532 2943
rect 1526 2938 1532 2939
rect 1638 2943 1644 2944
rect 1638 2939 1639 2943
rect 1643 2939 1644 2943
rect 1638 2938 1644 2939
rect 1734 2943 1740 2944
rect 1734 2939 1735 2943
rect 1739 2939 1740 2943
rect 1734 2938 1740 2939
rect 1416 2927 1418 2938
rect 1528 2927 1530 2938
rect 1640 2927 1642 2938
rect 1736 2927 1738 2938
rect 1824 2927 1826 2951
rect 111 2926 115 2927
rect 111 2921 115 2922
rect 1359 2926 1363 2927
rect 1359 2921 1363 2922
rect 1415 2926 1419 2927
rect 1415 2921 1419 2922
rect 1471 2926 1475 2927
rect 1471 2921 1475 2922
rect 1527 2926 1531 2927
rect 1527 2921 1531 2922
rect 1583 2926 1587 2927
rect 1583 2921 1587 2922
rect 1639 2926 1643 2927
rect 1639 2921 1643 2922
rect 1703 2926 1707 2927
rect 1703 2921 1707 2922
rect 1735 2926 1739 2927
rect 1735 2921 1739 2922
rect 1823 2926 1827 2927
rect 1823 2921 1827 2922
rect 112 2897 114 2921
rect 1360 2910 1362 2921
rect 1472 2910 1474 2921
rect 1584 2910 1586 2921
rect 1704 2910 1706 2921
rect 1358 2909 1364 2910
rect 1358 2905 1359 2909
rect 1363 2905 1364 2909
rect 1358 2904 1364 2905
rect 1470 2909 1476 2910
rect 1470 2905 1471 2909
rect 1475 2905 1476 2909
rect 1470 2904 1476 2905
rect 1582 2909 1588 2910
rect 1582 2905 1583 2909
rect 1587 2905 1588 2909
rect 1582 2904 1588 2905
rect 1702 2909 1708 2910
rect 1702 2905 1703 2909
rect 1707 2905 1708 2909
rect 1702 2904 1708 2905
rect 1824 2897 1826 2921
rect 1864 2915 1866 2955
rect 2246 2947 2252 2948
rect 2246 2943 2247 2947
rect 2251 2943 2252 2947
rect 2246 2942 2252 2943
rect 2470 2947 2476 2948
rect 2470 2943 2471 2947
rect 2475 2943 2476 2947
rect 2470 2942 2476 2943
rect 2678 2947 2684 2948
rect 2678 2943 2679 2947
rect 2683 2943 2684 2947
rect 2678 2942 2684 2943
rect 2870 2947 2876 2948
rect 2870 2943 2871 2947
rect 2875 2943 2876 2947
rect 2870 2942 2876 2943
rect 3038 2947 3044 2948
rect 3038 2943 3039 2947
rect 3043 2943 3044 2947
rect 3038 2942 3044 2943
rect 3198 2947 3204 2948
rect 3198 2943 3199 2947
rect 3203 2943 3204 2947
rect 3198 2942 3204 2943
rect 3350 2947 3356 2948
rect 3350 2943 3351 2947
rect 3355 2943 3356 2947
rect 3350 2942 3356 2943
rect 3486 2947 3492 2948
rect 3486 2943 3487 2947
rect 3491 2943 3492 2947
rect 3486 2942 3492 2943
rect 2248 2915 2250 2942
rect 2472 2915 2474 2942
rect 2680 2915 2682 2942
rect 2872 2915 2874 2942
rect 3040 2915 3042 2942
rect 3200 2915 3202 2942
rect 3352 2915 3354 2942
rect 3488 2915 3490 2942
rect 3576 2915 3578 2955
rect 1863 2914 1867 2915
rect 1863 2909 1867 2910
rect 2239 2914 2243 2915
rect 2239 2909 2243 2910
rect 2247 2914 2251 2915
rect 2247 2909 2251 2910
rect 2463 2914 2467 2915
rect 2463 2909 2467 2910
rect 2471 2914 2475 2915
rect 2471 2909 2475 2910
rect 2671 2914 2675 2915
rect 2671 2909 2675 2910
rect 2679 2914 2683 2915
rect 2679 2909 2683 2910
rect 2855 2914 2859 2915
rect 2855 2909 2859 2910
rect 2871 2914 2875 2915
rect 2871 2909 2875 2910
rect 3023 2914 3027 2915
rect 3023 2909 3027 2910
rect 3039 2914 3043 2915
rect 3039 2909 3043 2910
rect 3183 2914 3187 2915
rect 3183 2909 3187 2910
rect 3199 2914 3203 2915
rect 3199 2909 3203 2910
rect 3335 2914 3339 2915
rect 3335 2909 3339 2910
rect 3351 2914 3355 2915
rect 3351 2909 3355 2910
rect 3487 2914 3491 2915
rect 3487 2909 3491 2910
rect 3575 2914 3579 2915
rect 3575 2909 3579 2910
rect 110 2896 116 2897
rect 110 2892 111 2896
rect 115 2892 116 2896
rect 110 2891 116 2892
rect 1822 2896 1828 2897
rect 1822 2892 1823 2896
rect 1827 2892 1828 2896
rect 1822 2891 1828 2892
rect 1864 2885 1866 2909
rect 2240 2898 2242 2909
rect 2464 2898 2466 2909
rect 2672 2898 2674 2909
rect 2856 2898 2858 2909
rect 3024 2898 3026 2909
rect 3184 2898 3186 2909
rect 3336 2898 3338 2909
rect 3488 2898 3490 2909
rect 2238 2897 2244 2898
rect 2238 2893 2239 2897
rect 2243 2893 2244 2897
rect 2238 2892 2244 2893
rect 2462 2897 2468 2898
rect 2462 2893 2463 2897
rect 2467 2893 2468 2897
rect 2462 2892 2468 2893
rect 2670 2897 2676 2898
rect 2670 2893 2671 2897
rect 2675 2893 2676 2897
rect 2670 2892 2676 2893
rect 2854 2897 2860 2898
rect 2854 2893 2855 2897
rect 2859 2893 2860 2897
rect 2854 2892 2860 2893
rect 3022 2897 3028 2898
rect 3022 2893 3023 2897
rect 3027 2893 3028 2897
rect 3022 2892 3028 2893
rect 3182 2897 3188 2898
rect 3182 2893 3183 2897
rect 3187 2893 3188 2897
rect 3182 2892 3188 2893
rect 3334 2897 3340 2898
rect 3334 2893 3335 2897
rect 3339 2893 3340 2897
rect 3334 2892 3340 2893
rect 3486 2897 3492 2898
rect 3486 2893 3487 2897
rect 3491 2893 3492 2897
rect 3486 2892 3492 2893
rect 3576 2885 3578 2909
rect 1862 2884 1868 2885
rect 1862 2880 1863 2884
rect 1867 2880 1868 2884
rect 110 2879 116 2880
rect 110 2875 111 2879
rect 115 2875 116 2879
rect 110 2874 116 2875
rect 1822 2879 1828 2880
rect 1862 2879 1868 2880
rect 3574 2884 3580 2885
rect 3574 2880 3575 2884
rect 3579 2880 3580 2884
rect 3574 2879 3580 2880
rect 1822 2875 1823 2879
rect 1827 2875 1828 2879
rect 1822 2874 1828 2875
rect 112 2855 114 2874
rect 1350 2869 1356 2870
rect 1350 2865 1351 2869
rect 1355 2865 1356 2869
rect 1350 2864 1356 2865
rect 1462 2869 1468 2870
rect 1462 2865 1463 2869
rect 1467 2865 1468 2869
rect 1462 2864 1468 2865
rect 1574 2869 1580 2870
rect 1574 2865 1575 2869
rect 1579 2865 1580 2869
rect 1574 2864 1580 2865
rect 1694 2869 1700 2870
rect 1694 2865 1695 2869
rect 1699 2865 1700 2869
rect 1694 2864 1700 2865
rect 1352 2855 1354 2864
rect 1464 2855 1466 2864
rect 1576 2855 1578 2864
rect 1696 2855 1698 2864
rect 1824 2855 1826 2874
rect 1862 2867 1868 2868
rect 1862 2863 1863 2867
rect 1867 2863 1868 2867
rect 1862 2862 1868 2863
rect 3574 2867 3580 2868
rect 3574 2863 3575 2867
rect 3579 2863 3580 2867
rect 3574 2862 3580 2863
rect 111 2854 115 2855
rect 111 2849 115 2850
rect 135 2854 139 2855
rect 135 2849 139 2850
rect 223 2854 227 2855
rect 223 2849 227 2850
rect 311 2854 315 2855
rect 311 2849 315 2850
rect 399 2854 403 2855
rect 399 2849 403 2850
rect 487 2854 491 2855
rect 487 2849 491 2850
rect 599 2854 603 2855
rect 599 2849 603 2850
rect 727 2854 731 2855
rect 727 2849 731 2850
rect 863 2854 867 2855
rect 863 2849 867 2850
rect 999 2854 1003 2855
rect 999 2849 1003 2850
rect 1135 2854 1139 2855
rect 1135 2849 1139 2850
rect 1263 2854 1267 2855
rect 1263 2849 1267 2850
rect 1351 2854 1355 2855
rect 1351 2849 1355 2850
rect 1383 2854 1387 2855
rect 1383 2849 1387 2850
rect 1463 2854 1467 2855
rect 1463 2849 1467 2850
rect 1503 2854 1507 2855
rect 1503 2849 1507 2850
rect 1575 2854 1579 2855
rect 1575 2849 1579 2850
rect 1623 2854 1627 2855
rect 1623 2849 1627 2850
rect 1695 2854 1699 2855
rect 1695 2849 1699 2850
rect 1727 2854 1731 2855
rect 1727 2849 1731 2850
rect 1823 2854 1827 2855
rect 1823 2849 1827 2850
rect 112 2834 114 2849
rect 136 2844 138 2849
rect 224 2844 226 2849
rect 312 2844 314 2849
rect 400 2844 402 2849
rect 488 2844 490 2849
rect 600 2844 602 2849
rect 728 2844 730 2849
rect 864 2844 866 2849
rect 1000 2844 1002 2849
rect 1136 2844 1138 2849
rect 1264 2844 1266 2849
rect 1384 2844 1386 2849
rect 1504 2844 1506 2849
rect 1624 2844 1626 2849
rect 1728 2844 1730 2849
rect 134 2843 140 2844
rect 134 2839 135 2843
rect 139 2839 140 2843
rect 134 2838 140 2839
rect 222 2843 228 2844
rect 222 2839 223 2843
rect 227 2839 228 2843
rect 222 2838 228 2839
rect 310 2843 316 2844
rect 310 2839 311 2843
rect 315 2839 316 2843
rect 310 2838 316 2839
rect 398 2843 404 2844
rect 398 2839 399 2843
rect 403 2839 404 2843
rect 398 2838 404 2839
rect 486 2843 492 2844
rect 486 2839 487 2843
rect 491 2839 492 2843
rect 486 2838 492 2839
rect 598 2843 604 2844
rect 598 2839 599 2843
rect 603 2839 604 2843
rect 598 2838 604 2839
rect 726 2843 732 2844
rect 726 2839 727 2843
rect 731 2839 732 2843
rect 726 2838 732 2839
rect 862 2843 868 2844
rect 862 2839 863 2843
rect 867 2839 868 2843
rect 862 2838 868 2839
rect 998 2843 1004 2844
rect 998 2839 999 2843
rect 1003 2839 1004 2843
rect 998 2838 1004 2839
rect 1134 2843 1140 2844
rect 1134 2839 1135 2843
rect 1139 2839 1140 2843
rect 1134 2838 1140 2839
rect 1262 2843 1268 2844
rect 1262 2839 1263 2843
rect 1267 2839 1268 2843
rect 1262 2838 1268 2839
rect 1382 2843 1388 2844
rect 1382 2839 1383 2843
rect 1387 2839 1388 2843
rect 1382 2838 1388 2839
rect 1502 2843 1508 2844
rect 1502 2839 1503 2843
rect 1507 2839 1508 2843
rect 1502 2838 1508 2839
rect 1622 2843 1628 2844
rect 1622 2839 1623 2843
rect 1627 2839 1628 2843
rect 1622 2838 1628 2839
rect 1726 2843 1732 2844
rect 1726 2839 1727 2843
rect 1731 2839 1732 2843
rect 1726 2838 1732 2839
rect 1824 2834 1826 2849
rect 1864 2843 1866 2862
rect 2230 2857 2236 2858
rect 2230 2853 2231 2857
rect 2235 2853 2236 2857
rect 2230 2852 2236 2853
rect 2454 2857 2460 2858
rect 2454 2853 2455 2857
rect 2459 2853 2460 2857
rect 2454 2852 2460 2853
rect 2662 2857 2668 2858
rect 2662 2853 2663 2857
rect 2667 2853 2668 2857
rect 2662 2852 2668 2853
rect 2846 2857 2852 2858
rect 2846 2853 2847 2857
rect 2851 2853 2852 2857
rect 2846 2852 2852 2853
rect 3014 2857 3020 2858
rect 3014 2853 3015 2857
rect 3019 2853 3020 2857
rect 3014 2852 3020 2853
rect 3174 2857 3180 2858
rect 3174 2853 3175 2857
rect 3179 2853 3180 2857
rect 3174 2852 3180 2853
rect 3326 2857 3332 2858
rect 3326 2853 3327 2857
rect 3331 2853 3332 2857
rect 3326 2852 3332 2853
rect 3478 2857 3484 2858
rect 3478 2853 3479 2857
rect 3483 2853 3484 2857
rect 3478 2852 3484 2853
rect 2232 2843 2234 2852
rect 2456 2843 2458 2852
rect 2664 2843 2666 2852
rect 2848 2843 2850 2852
rect 3016 2843 3018 2852
rect 3176 2843 3178 2852
rect 3328 2843 3330 2852
rect 3480 2843 3482 2852
rect 3576 2843 3578 2862
rect 1863 2842 1867 2843
rect 1863 2837 1867 2838
rect 1895 2842 1899 2843
rect 1895 2837 1899 2838
rect 1983 2842 1987 2843
rect 1983 2837 1987 2838
rect 2071 2842 2075 2843
rect 2071 2837 2075 2838
rect 2159 2842 2163 2843
rect 2159 2837 2163 2838
rect 2231 2842 2235 2843
rect 2231 2837 2235 2838
rect 2247 2842 2251 2843
rect 2247 2837 2251 2838
rect 2335 2842 2339 2843
rect 2335 2837 2339 2838
rect 2423 2842 2427 2843
rect 2423 2837 2427 2838
rect 2455 2842 2459 2843
rect 2455 2837 2459 2838
rect 2511 2842 2515 2843
rect 2511 2837 2515 2838
rect 2599 2842 2603 2843
rect 2599 2837 2603 2838
rect 2663 2842 2667 2843
rect 2663 2837 2667 2838
rect 2687 2842 2691 2843
rect 2687 2837 2691 2838
rect 2791 2842 2795 2843
rect 2791 2837 2795 2838
rect 2847 2842 2851 2843
rect 2847 2837 2851 2838
rect 2903 2842 2907 2843
rect 2903 2837 2907 2838
rect 3015 2842 3019 2843
rect 3015 2837 3019 2838
rect 3031 2842 3035 2843
rect 3031 2837 3035 2838
rect 3175 2842 3179 2843
rect 3175 2837 3179 2838
rect 3327 2842 3331 2843
rect 3327 2837 3331 2838
rect 3479 2842 3483 2843
rect 3479 2837 3483 2838
rect 3575 2842 3579 2843
rect 3575 2837 3579 2838
rect 110 2833 116 2834
rect 110 2829 111 2833
rect 115 2829 116 2833
rect 110 2828 116 2829
rect 1822 2833 1828 2834
rect 1822 2829 1823 2833
rect 1827 2829 1828 2833
rect 1822 2828 1828 2829
rect 1864 2822 1866 2837
rect 1896 2832 1898 2837
rect 1984 2832 1986 2837
rect 2072 2832 2074 2837
rect 2160 2832 2162 2837
rect 2248 2832 2250 2837
rect 2336 2832 2338 2837
rect 2424 2832 2426 2837
rect 2512 2832 2514 2837
rect 2600 2832 2602 2837
rect 2688 2832 2690 2837
rect 2792 2832 2794 2837
rect 2904 2832 2906 2837
rect 3032 2832 3034 2837
rect 3176 2832 3178 2837
rect 3328 2832 3330 2837
rect 3480 2832 3482 2837
rect 1894 2831 1900 2832
rect 1894 2827 1895 2831
rect 1899 2827 1900 2831
rect 1894 2826 1900 2827
rect 1982 2831 1988 2832
rect 1982 2827 1983 2831
rect 1987 2827 1988 2831
rect 1982 2826 1988 2827
rect 2070 2831 2076 2832
rect 2070 2827 2071 2831
rect 2075 2827 2076 2831
rect 2070 2826 2076 2827
rect 2158 2831 2164 2832
rect 2158 2827 2159 2831
rect 2163 2827 2164 2831
rect 2158 2826 2164 2827
rect 2246 2831 2252 2832
rect 2246 2827 2247 2831
rect 2251 2827 2252 2831
rect 2246 2826 2252 2827
rect 2334 2831 2340 2832
rect 2334 2827 2335 2831
rect 2339 2827 2340 2831
rect 2334 2826 2340 2827
rect 2422 2831 2428 2832
rect 2422 2827 2423 2831
rect 2427 2827 2428 2831
rect 2422 2826 2428 2827
rect 2510 2831 2516 2832
rect 2510 2827 2511 2831
rect 2515 2827 2516 2831
rect 2510 2826 2516 2827
rect 2598 2831 2604 2832
rect 2598 2827 2599 2831
rect 2603 2827 2604 2831
rect 2598 2826 2604 2827
rect 2686 2831 2692 2832
rect 2686 2827 2687 2831
rect 2691 2827 2692 2831
rect 2686 2826 2692 2827
rect 2790 2831 2796 2832
rect 2790 2827 2791 2831
rect 2795 2827 2796 2831
rect 2790 2826 2796 2827
rect 2902 2831 2908 2832
rect 2902 2827 2903 2831
rect 2907 2827 2908 2831
rect 2902 2826 2908 2827
rect 3030 2831 3036 2832
rect 3030 2827 3031 2831
rect 3035 2827 3036 2831
rect 3030 2826 3036 2827
rect 3174 2831 3180 2832
rect 3174 2827 3175 2831
rect 3179 2827 3180 2831
rect 3174 2826 3180 2827
rect 3326 2831 3332 2832
rect 3326 2827 3327 2831
rect 3331 2827 3332 2831
rect 3326 2826 3332 2827
rect 3478 2831 3484 2832
rect 3478 2827 3479 2831
rect 3483 2827 3484 2831
rect 3478 2826 3484 2827
rect 3576 2822 3578 2837
rect 1862 2821 1868 2822
rect 1862 2817 1863 2821
rect 1867 2817 1868 2821
rect 110 2816 116 2817
rect 110 2812 111 2816
rect 115 2812 116 2816
rect 110 2811 116 2812
rect 1822 2816 1828 2817
rect 1862 2816 1868 2817
rect 3574 2821 3580 2822
rect 3574 2817 3575 2821
rect 3579 2817 3580 2821
rect 3574 2816 3580 2817
rect 1822 2812 1823 2816
rect 1827 2812 1828 2816
rect 1822 2811 1828 2812
rect 112 2787 114 2811
rect 142 2803 148 2804
rect 142 2799 143 2803
rect 147 2799 148 2803
rect 142 2798 148 2799
rect 230 2803 236 2804
rect 230 2799 231 2803
rect 235 2799 236 2803
rect 230 2798 236 2799
rect 318 2803 324 2804
rect 318 2799 319 2803
rect 323 2799 324 2803
rect 318 2798 324 2799
rect 406 2803 412 2804
rect 406 2799 407 2803
rect 411 2799 412 2803
rect 406 2798 412 2799
rect 494 2803 500 2804
rect 494 2799 495 2803
rect 499 2799 500 2803
rect 494 2798 500 2799
rect 606 2803 612 2804
rect 606 2799 607 2803
rect 611 2799 612 2803
rect 606 2798 612 2799
rect 734 2803 740 2804
rect 734 2799 735 2803
rect 739 2799 740 2803
rect 734 2798 740 2799
rect 870 2803 876 2804
rect 870 2799 871 2803
rect 875 2799 876 2803
rect 870 2798 876 2799
rect 1006 2803 1012 2804
rect 1006 2799 1007 2803
rect 1011 2799 1012 2803
rect 1006 2798 1012 2799
rect 1142 2803 1148 2804
rect 1142 2799 1143 2803
rect 1147 2799 1148 2803
rect 1142 2798 1148 2799
rect 1270 2803 1276 2804
rect 1270 2799 1271 2803
rect 1275 2799 1276 2803
rect 1270 2798 1276 2799
rect 1390 2803 1396 2804
rect 1390 2799 1391 2803
rect 1395 2799 1396 2803
rect 1390 2798 1396 2799
rect 1510 2803 1516 2804
rect 1510 2799 1511 2803
rect 1515 2799 1516 2803
rect 1510 2798 1516 2799
rect 1630 2803 1636 2804
rect 1630 2799 1631 2803
rect 1635 2799 1636 2803
rect 1630 2798 1636 2799
rect 1734 2803 1740 2804
rect 1734 2799 1735 2803
rect 1739 2799 1740 2803
rect 1734 2798 1740 2799
rect 144 2787 146 2798
rect 232 2787 234 2798
rect 320 2787 322 2798
rect 408 2787 410 2798
rect 496 2787 498 2798
rect 608 2787 610 2798
rect 736 2787 738 2798
rect 872 2787 874 2798
rect 1008 2787 1010 2798
rect 1144 2787 1146 2798
rect 1272 2787 1274 2798
rect 1392 2787 1394 2798
rect 1512 2787 1514 2798
rect 1632 2787 1634 2798
rect 1736 2787 1738 2798
rect 1824 2787 1826 2811
rect 1862 2804 1868 2805
rect 1862 2800 1863 2804
rect 1867 2800 1868 2804
rect 1862 2799 1868 2800
rect 3574 2804 3580 2805
rect 3574 2800 3575 2804
rect 3579 2800 3580 2804
rect 3574 2799 3580 2800
rect 111 2786 115 2787
rect 111 2781 115 2782
rect 143 2786 147 2787
rect 143 2781 147 2782
rect 191 2786 195 2787
rect 191 2781 195 2782
rect 231 2786 235 2787
rect 231 2781 235 2782
rect 295 2786 299 2787
rect 295 2781 299 2782
rect 319 2786 323 2787
rect 319 2781 323 2782
rect 407 2786 411 2787
rect 407 2781 411 2782
rect 415 2786 419 2787
rect 415 2781 419 2782
rect 495 2786 499 2787
rect 495 2781 499 2782
rect 551 2786 555 2787
rect 551 2781 555 2782
rect 607 2786 611 2787
rect 607 2781 611 2782
rect 687 2786 691 2787
rect 687 2781 691 2782
rect 735 2786 739 2787
rect 735 2781 739 2782
rect 823 2786 827 2787
rect 823 2781 827 2782
rect 871 2786 875 2787
rect 871 2781 875 2782
rect 959 2786 963 2787
rect 959 2781 963 2782
rect 1007 2786 1011 2787
rect 1007 2781 1011 2782
rect 1087 2786 1091 2787
rect 1087 2781 1091 2782
rect 1143 2786 1147 2787
rect 1143 2781 1147 2782
rect 1207 2786 1211 2787
rect 1207 2781 1211 2782
rect 1271 2786 1275 2787
rect 1271 2781 1275 2782
rect 1319 2786 1323 2787
rect 1319 2781 1323 2782
rect 1391 2786 1395 2787
rect 1391 2781 1395 2782
rect 1431 2786 1435 2787
rect 1431 2781 1435 2782
rect 1511 2786 1515 2787
rect 1511 2781 1515 2782
rect 1535 2786 1539 2787
rect 1535 2781 1539 2782
rect 1631 2786 1635 2787
rect 1631 2781 1635 2782
rect 1647 2786 1651 2787
rect 1647 2781 1651 2782
rect 1735 2786 1739 2787
rect 1735 2781 1739 2782
rect 1823 2786 1827 2787
rect 1823 2781 1827 2782
rect 112 2757 114 2781
rect 192 2770 194 2781
rect 296 2770 298 2781
rect 416 2770 418 2781
rect 552 2770 554 2781
rect 688 2770 690 2781
rect 824 2770 826 2781
rect 960 2770 962 2781
rect 1088 2770 1090 2781
rect 1208 2770 1210 2781
rect 1320 2770 1322 2781
rect 1432 2770 1434 2781
rect 1536 2770 1538 2781
rect 1648 2770 1650 2781
rect 1736 2770 1738 2781
rect 190 2769 196 2770
rect 190 2765 191 2769
rect 195 2765 196 2769
rect 190 2764 196 2765
rect 294 2769 300 2770
rect 294 2765 295 2769
rect 299 2765 300 2769
rect 294 2764 300 2765
rect 414 2769 420 2770
rect 414 2765 415 2769
rect 419 2765 420 2769
rect 414 2764 420 2765
rect 550 2769 556 2770
rect 550 2765 551 2769
rect 555 2765 556 2769
rect 550 2764 556 2765
rect 686 2769 692 2770
rect 686 2765 687 2769
rect 691 2765 692 2769
rect 686 2764 692 2765
rect 822 2769 828 2770
rect 822 2765 823 2769
rect 827 2765 828 2769
rect 822 2764 828 2765
rect 958 2769 964 2770
rect 958 2765 959 2769
rect 963 2765 964 2769
rect 958 2764 964 2765
rect 1086 2769 1092 2770
rect 1086 2765 1087 2769
rect 1091 2765 1092 2769
rect 1086 2764 1092 2765
rect 1206 2769 1212 2770
rect 1206 2765 1207 2769
rect 1211 2765 1212 2769
rect 1206 2764 1212 2765
rect 1318 2769 1324 2770
rect 1318 2765 1319 2769
rect 1323 2765 1324 2769
rect 1318 2764 1324 2765
rect 1430 2769 1436 2770
rect 1430 2765 1431 2769
rect 1435 2765 1436 2769
rect 1430 2764 1436 2765
rect 1534 2769 1540 2770
rect 1534 2765 1535 2769
rect 1539 2765 1540 2769
rect 1534 2764 1540 2765
rect 1646 2769 1652 2770
rect 1646 2765 1647 2769
rect 1651 2765 1652 2769
rect 1646 2764 1652 2765
rect 1734 2769 1740 2770
rect 1734 2765 1735 2769
rect 1739 2765 1740 2769
rect 1734 2764 1740 2765
rect 1824 2757 1826 2781
rect 1864 2763 1866 2799
rect 1902 2791 1908 2792
rect 1902 2787 1903 2791
rect 1907 2787 1908 2791
rect 1902 2786 1908 2787
rect 1990 2791 1996 2792
rect 1990 2787 1991 2791
rect 1995 2787 1996 2791
rect 1990 2786 1996 2787
rect 2078 2791 2084 2792
rect 2078 2787 2079 2791
rect 2083 2787 2084 2791
rect 2078 2786 2084 2787
rect 2166 2791 2172 2792
rect 2166 2787 2167 2791
rect 2171 2787 2172 2791
rect 2166 2786 2172 2787
rect 2254 2791 2260 2792
rect 2254 2787 2255 2791
rect 2259 2787 2260 2791
rect 2254 2786 2260 2787
rect 2342 2791 2348 2792
rect 2342 2787 2343 2791
rect 2347 2787 2348 2791
rect 2342 2786 2348 2787
rect 2430 2791 2436 2792
rect 2430 2787 2431 2791
rect 2435 2787 2436 2791
rect 2430 2786 2436 2787
rect 2518 2791 2524 2792
rect 2518 2787 2519 2791
rect 2523 2787 2524 2791
rect 2518 2786 2524 2787
rect 2606 2791 2612 2792
rect 2606 2787 2607 2791
rect 2611 2787 2612 2791
rect 2606 2786 2612 2787
rect 2694 2791 2700 2792
rect 2694 2787 2695 2791
rect 2699 2787 2700 2791
rect 2694 2786 2700 2787
rect 2798 2791 2804 2792
rect 2798 2787 2799 2791
rect 2803 2787 2804 2791
rect 2798 2786 2804 2787
rect 2910 2791 2916 2792
rect 2910 2787 2911 2791
rect 2915 2787 2916 2791
rect 2910 2786 2916 2787
rect 3038 2791 3044 2792
rect 3038 2787 3039 2791
rect 3043 2787 3044 2791
rect 3038 2786 3044 2787
rect 3182 2791 3188 2792
rect 3182 2787 3183 2791
rect 3187 2787 3188 2791
rect 3182 2786 3188 2787
rect 3334 2791 3340 2792
rect 3334 2787 3335 2791
rect 3339 2787 3340 2791
rect 3334 2786 3340 2787
rect 3486 2791 3492 2792
rect 3486 2787 3487 2791
rect 3491 2787 3492 2791
rect 3486 2786 3492 2787
rect 1904 2763 1906 2786
rect 1992 2763 1994 2786
rect 2080 2763 2082 2786
rect 2168 2763 2170 2786
rect 2256 2763 2258 2786
rect 2344 2763 2346 2786
rect 2432 2763 2434 2786
rect 2520 2763 2522 2786
rect 2608 2763 2610 2786
rect 2696 2763 2698 2786
rect 2800 2763 2802 2786
rect 2912 2763 2914 2786
rect 3040 2763 3042 2786
rect 3184 2763 3186 2786
rect 3336 2763 3338 2786
rect 3488 2763 3490 2786
rect 3576 2763 3578 2799
rect 1863 2762 1867 2763
rect 1863 2757 1867 2758
rect 1903 2762 1907 2763
rect 1903 2757 1907 2758
rect 1991 2762 1995 2763
rect 1991 2757 1995 2758
rect 2047 2762 2051 2763
rect 2047 2757 2051 2758
rect 2079 2762 2083 2763
rect 2079 2757 2083 2758
rect 2167 2762 2171 2763
rect 2167 2757 2171 2758
rect 2255 2762 2259 2763
rect 2255 2757 2259 2758
rect 2295 2762 2299 2763
rect 2295 2757 2299 2758
rect 2343 2762 2347 2763
rect 2343 2757 2347 2758
rect 2431 2762 2435 2763
rect 2431 2757 2435 2758
rect 2447 2762 2451 2763
rect 2447 2757 2451 2758
rect 2519 2762 2523 2763
rect 2519 2757 2523 2758
rect 2607 2762 2611 2763
rect 2607 2757 2611 2758
rect 2623 2762 2627 2763
rect 2623 2757 2627 2758
rect 2695 2762 2699 2763
rect 2695 2757 2699 2758
rect 2799 2762 2803 2763
rect 2799 2757 2803 2758
rect 2823 2762 2827 2763
rect 2823 2757 2827 2758
rect 2911 2762 2915 2763
rect 2911 2757 2915 2758
rect 3039 2762 3043 2763
rect 3039 2757 3043 2758
rect 3183 2762 3187 2763
rect 3183 2757 3187 2758
rect 3271 2762 3275 2763
rect 3271 2757 3275 2758
rect 3335 2762 3339 2763
rect 3335 2757 3339 2758
rect 3487 2762 3491 2763
rect 3487 2757 3491 2758
rect 3575 2762 3579 2763
rect 3575 2757 3579 2758
rect 110 2756 116 2757
rect 110 2752 111 2756
rect 115 2752 116 2756
rect 110 2751 116 2752
rect 1822 2756 1828 2757
rect 1822 2752 1823 2756
rect 1827 2752 1828 2756
rect 1822 2751 1828 2752
rect 110 2739 116 2740
rect 110 2735 111 2739
rect 115 2735 116 2739
rect 110 2734 116 2735
rect 1822 2739 1828 2740
rect 1822 2735 1823 2739
rect 1827 2735 1828 2739
rect 1822 2734 1828 2735
rect 112 2711 114 2734
rect 182 2729 188 2730
rect 182 2725 183 2729
rect 187 2725 188 2729
rect 182 2724 188 2725
rect 286 2729 292 2730
rect 286 2725 287 2729
rect 291 2725 292 2729
rect 286 2724 292 2725
rect 406 2729 412 2730
rect 406 2725 407 2729
rect 411 2725 412 2729
rect 406 2724 412 2725
rect 542 2729 548 2730
rect 542 2725 543 2729
rect 547 2725 548 2729
rect 542 2724 548 2725
rect 678 2729 684 2730
rect 678 2725 679 2729
rect 683 2725 684 2729
rect 678 2724 684 2725
rect 814 2729 820 2730
rect 814 2725 815 2729
rect 819 2725 820 2729
rect 814 2724 820 2725
rect 950 2729 956 2730
rect 950 2725 951 2729
rect 955 2725 956 2729
rect 950 2724 956 2725
rect 1078 2729 1084 2730
rect 1078 2725 1079 2729
rect 1083 2725 1084 2729
rect 1078 2724 1084 2725
rect 1198 2729 1204 2730
rect 1198 2725 1199 2729
rect 1203 2725 1204 2729
rect 1198 2724 1204 2725
rect 1310 2729 1316 2730
rect 1310 2725 1311 2729
rect 1315 2725 1316 2729
rect 1310 2724 1316 2725
rect 1422 2729 1428 2730
rect 1422 2725 1423 2729
rect 1427 2725 1428 2729
rect 1422 2724 1428 2725
rect 1526 2729 1532 2730
rect 1526 2725 1527 2729
rect 1531 2725 1532 2729
rect 1526 2724 1532 2725
rect 1638 2729 1644 2730
rect 1638 2725 1639 2729
rect 1643 2725 1644 2729
rect 1638 2724 1644 2725
rect 1726 2729 1732 2730
rect 1726 2725 1727 2729
rect 1731 2725 1732 2729
rect 1726 2724 1732 2725
rect 184 2711 186 2724
rect 288 2711 290 2724
rect 408 2711 410 2724
rect 544 2711 546 2724
rect 680 2711 682 2724
rect 816 2711 818 2724
rect 952 2711 954 2724
rect 1080 2711 1082 2724
rect 1200 2711 1202 2724
rect 1312 2711 1314 2724
rect 1424 2711 1426 2724
rect 1528 2711 1530 2724
rect 1640 2711 1642 2724
rect 1728 2711 1730 2724
rect 1824 2711 1826 2734
rect 1864 2733 1866 2757
rect 2048 2746 2050 2757
rect 2168 2746 2170 2757
rect 2296 2746 2298 2757
rect 2448 2746 2450 2757
rect 2624 2746 2626 2757
rect 2824 2746 2826 2757
rect 3040 2746 3042 2757
rect 3272 2746 3274 2757
rect 3488 2746 3490 2757
rect 2046 2745 2052 2746
rect 2046 2741 2047 2745
rect 2051 2741 2052 2745
rect 2046 2740 2052 2741
rect 2166 2745 2172 2746
rect 2166 2741 2167 2745
rect 2171 2741 2172 2745
rect 2166 2740 2172 2741
rect 2294 2745 2300 2746
rect 2294 2741 2295 2745
rect 2299 2741 2300 2745
rect 2294 2740 2300 2741
rect 2446 2745 2452 2746
rect 2446 2741 2447 2745
rect 2451 2741 2452 2745
rect 2446 2740 2452 2741
rect 2622 2745 2628 2746
rect 2622 2741 2623 2745
rect 2627 2741 2628 2745
rect 2622 2740 2628 2741
rect 2822 2745 2828 2746
rect 2822 2741 2823 2745
rect 2827 2741 2828 2745
rect 2822 2740 2828 2741
rect 3038 2745 3044 2746
rect 3038 2741 3039 2745
rect 3043 2741 3044 2745
rect 3038 2740 3044 2741
rect 3270 2745 3276 2746
rect 3270 2741 3271 2745
rect 3275 2741 3276 2745
rect 3270 2740 3276 2741
rect 3486 2745 3492 2746
rect 3486 2741 3487 2745
rect 3491 2741 3492 2745
rect 3486 2740 3492 2741
rect 3576 2733 3578 2757
rect 1862 2732 1868 2733
rect 1862 2728 1863 2732
rect 1867 2728 1868 2732
rect 1862 2727 1868 2728
rect 3574 2732 3580 2733
rect 3574 2728 3575 2732
rect 3579 2728 3580 2732
rect 3574 2727 3580 2728
rect 1862 2715 1868 2716
rect 1862 2711 1863 2715
rect 1867 2711 1868 2715
rect 111 2710 115 2711
rect 111 2705 115 2706
rect 167 2710 171 2711
rect 167 2705 171 2706
rect 183 2710 187 2711
rect 183 2705 187 2706
rect 279 2710 283 2711
rect 279 2705 283 2706
rect 287 2710 291 2711
rect 287 2705 291 2706
rect 391 2710 395 2711
rect 391 2705 395 2706
rect 407 2710 411 2711
rect 407 2705 411 2706
rect 503 2710 507 2711
rect 503 2705 507 2706
rect 543 2710 547 2711
rect 543 2705 547 2706
rect 615 2710 619 2711
rect 615 2705 619 2706
rect 679 2710 683 2711
rect 679 2705 683 2706
rect 815 2710 819 2711
rect 815 2705 819 2706
rect 951 2710 955 2711
rect 951 2705 955 2706
rect 1079 2710 1083 2711
rect 1079 2705 1083 2706
rect 1199 2710 1203 2711
rect 1199 2705 1203 2706
rect 1311 2710 1315 2711
rect 1311 2705 1315 2706
rect 1423 2710 1427 2711
rect 1423 2705 1427 2706
rect 1527 2710 1531 2711
rect 1527 2705 1531 2706
rect 1639 2710 1643 2711
rect 1639 2705 1643 2706
rect 1727 2710 1731 2711
rect 1727 2705 1731 2706
rect 1823 2710 1827 2711
rect 1862 2710 1868 2711
rect 3574 2715 3580 2716
rect 3574 2711 3575 2715
rect 3579 2711 3580 2715
rect 3574 2710 3580 2711
rect 1823 2705 1827 2706
rect 112 2690 114 2705
rect 168 2700 170 2705
rect 280 2700 282 2705
rect 392 2700 394 2705
rect 504 2700 506 2705
rect 616 2700 618 2705
rect 166 2699 172 2700
rect 166 2695 167 2699
rect 171 2695 172 2699
rect 166 2694 172 2695
rect 278 2699 284 2700
rect 278 2695 279 2699
rect 283 2695 284 2699
rect 278 2694 284 2695
rect 390 2699 396 2700
rect 390 2695 391 2699
rect 395 2695 396 2699
rect 390 2694 396 2695
rect 502 2699 508 2700
rect 502 2695 503 2699
rect 507 2695 508 2699
rect 502 2694 508 2695
rect 614 2699 620 2700
rect 614 2695 615 2699
rect 619 2695 620 2699
rect 614 2694 620 2695
rect 1824 2690 1826 2705
rect 1864 2695 1866 2710
rect 2038 2705 2044 2706
rect 2038 2701 2039 2705
rect 2043 2701 2044 2705
rect 2038 2700 2044 2701
rect 2158 2705 2164 2706
rect 2158 2701 2159 2705
rect 2163 2701 2164 2705
rect 2158 2700 2164 2701
rect 2286 2705 2292 2706
rect 2286 2701 2287 2705
rect 2291 2701 2292 2705
rect 2286 2700 2292 2701
rect 2438 2705 2444 2706
rect 2438 2701 2439 2705
rect 2443 2701 2444 2705
rect 2438 2700 2444 2701
rect 2614 2705 2620 2706
rect 2614 2701 2615 2705
rect 2619 2701 2620 2705
rect 2614 2700 2620 2701
rect 2814 2705 2820 2706
rect 2814 2701 2815 2705
rect 2819 2701 2820 2705
rect 2814 2700 2820 2701
rect 3030 2705 3036 2706
rect 3030 2701 3031 2705
rect 3035 2701 3036 2705
rect 3030 2700 3036 2701
rect 3262 2705 3268 2706
rect 3262 2701 3263 2705
rect 3267 2701 3268 2705
rect 3262 2700 3268 2701
rect 3478 2705 3484 2706
rect 3478 2701 3479 2705
rect 3483 2701 3484 2705
rect 3478 2700 3484 2701
rect 2040 2695 2042 2700
rect 2160 2695 2162 2700
rect 2288 2695 2290 2700
rect 2440 2695 2442 2700
rect 2616 2695 2618 2700
rect 2816 2695 2818 2700
rect 3032 2695 3034 2700
rect 3264 2695 3266 2700
rect 3480 2695 3482 2700
rect 3576 2695 3578 2710
rect 1863 2694 1867 2695
rect 110 2689 116 2690
rect 110 2685 111 2689
rect 115 2685 116 2689
rect 110 2684 116 2685
rect 1822 2689 1828 2690
rect 1863 2689 1867 2690
rect 1943 2694 1947 2695
rect 1943 2689 1947 2690
rect 2039 2694 2043 2695
rect 2039 2689 2043 2690
rect 2055 2694 2059 2695
rect 2055 2689 2059 2690
rect 2159 2694 2163 2695
rect 2159 2689 2163 2690
rect 2167 2694 2171 2695
rect 2167 2689 2171 2690
rect 2287 2694 2291 2695
rect 2287 2689 2291 2690
rect 2407 2694 2411 2695
rect 2407 2689 2411 2690
rect 2439 2694 2443 2695
rect 2439 2689 2443 2690
rect 2519 2694 2523 2695
rect 2519 2689 2523 2690
rect 2615 2694 2619 2695
rect 2615 2689 2619 2690
rect 2631 2694 2635 2695
rect 2631 2689 2635 2690
rect 2735 2694 2739 2695
rect 2735 2689 2739 2690
rect 2815 2694 2819 2695
rect 2815 2689 2819 2690
rect 2847 2694 2851 2695
rect 2847 2689 2851 2690
rect 2959 2694 2963 2695
rect 2959 2689 2963 2690
rect 3031 2694 3035 2695
rect 3031 2689 3035 2690
rect 3071 2694 3075 2695
rect 3071 2689 3075 2690
rect 3263 2694 3267 2695
rect 3263 2689 3267 2690
rect 3479 2694 3483 2695
rect 3479 2689 3483 2690
rect 3575 2694 3579 2695
rect 3575 2689 3579 2690
rect 1822 2685 1823 2689
rect 1827 2685 1828 2689
rect 1822 2684 1828 2685
rect 1864 2674 1866 2689
rect 1944 2684 1946 2689
rect 2056 2684 2058 2689
rect 2168 2684 2170 2689
rect 2288 2684 2290 2689
rect 2408 2684 2410 2689
rect 2520 2684 2522 2689
rect 2632 2684 2634 2689
rect 2736 2684 2738 2689
rect 2848 2684 2850 2689
rect 2960 2684 2962 2689
rect 3072 2684 3074 2689
rect 1942 2683 1948 2684
rect 1942 2679 1943 2683
rect 1947 2679 1948 2683
rect 1942 2678 1948 2679
rect 2054 2683 2060 2684
rect 2054 2679 2055 2683
rect 2059 2679 2060 2683
rect 2054 2678 2060 2679
rect 2166 2683 2172 2684
rect 2166 2679 2167 2683
rect 2171 2679 2172 2683
rect 2166 2678 2172 2679
rect 2286 2683 2292 2684
rect 2286 2679 2287 2683
rect 2291 2679 2292 2683
rect 2286 2678 2292 2679
rect 2406 2683 2412 2684
rect 2406 2679 2407 2683
rect 2411 2679 2412 2683
rect 2406 2678 2412 2679
rect 2518 2683 2524 2684
rect 2518 2679 2519 2683
rect 2523 2679 2524 2683
rect 2518 2678 2524 2679
rect 2630 2683 2636 2684
rect 2630 2679 2631 2683
rect 2635 2679 2636 2683
rect 2630 2678 2636 2679
rect 2734 2683 2740 2684
rect 2734 2679 2735 2683
rect 2739 2679 2740 2683
rect 2734 2678 2740 2679
rect 2846 2683 2852 2684
rect 2846 2679 2847 2683
rect 2851 2679 2852 2683
rect 2846 2678 2852 2679
rect 2958 2683 2964 2684
rect 2958 2679 2959 2683
rect 2963 2679 2964 2683
rect 2958 2678 2964 2679
rect 3070 2683 3076 2684
rect 3070 2679 3071 2683
rect 3075 2679 3076 2683
rect 3070 2678 3076 2679
rect 3576 2674 3578 2689
rect 1862 2673 1868 2674
rect 110 2672 116 2673
rect 110 2668 111 2672
rect 115 2668 116 2672
rect 110 2667 116 2668
rect 1822 2672 1828 2673
rect 1822 2668 1823 2672
rect 1827 2668 1828 2672
rect 1862 2669 1863 2673
rect 1867 2669 1868 2673
rect 1862 2668 1868 2669
rect 3574 2673 3580 2674
rect 3574 2669 3575 2673
rect 3579 2669 3580 2673
rect 3574 2668 3580 2669
rect 1822 2667 1828 2668
rect 112 2627 114 2667
rect 174 2659 180 2660
rect 174 2655 175 2659
rect 179 2655 180 2659
rect 174 2654 180 2655
rect 286 2659 292 2660
rect 286 2655 287 2659
rect 291 2655 292 2659
rect 286 2654 292 2655
rect 398 2659 404 2660
rect 398 2655 399 2659
rect 403 2655 404 2659
rect 398 2654 404 2655
rect 510 2659 516 2660
rect 510 2655 511 2659
rect 515 2655 516 2659
rect 510 2654 516 2655
rect 622 2659 628 2660
rect 622 2655 623 2659
rect 627 2655 628 2659
rect 622 2654 628 2655
rect 176 2627 178 2654
rect 288 2627 290 2654
rect 400 2627 402 2654
rect 512 2627 514 2654
rect 624 2627 626 2654
rect 1824 2627 1826 2667
rect 1862 2656 1868 2657
rect 1862 2652 1863 2656
rect 1867 2652 1868 2656
rect 1862 2651 1868 2652
rect 3574 2656 3580 2657
rect 3574 2652 3575 2656
rect 3579 2652 3580 2656
rect 3574 2651 3580 2652
rect 111 2626 115 2627
rect 111 2621 115 2622
rect 175 2626 179 2627
rect 175 2621 179 2622
rect 223 2626 227 2627
rect 223 2621 227 2622
rect 287 2626 291 2627
rect 287 2621 291 2622
rect 351 2626 355 2627
rect 351 2621 355 2622
rect 399 2626 403 2627
rect 399 2621 403 2622
rect 495 2626 499 2627
rect 495 2621 499 2622
rect 511 2626 515 2627
rect 511 2621 515 2622
rect 623 2626 627 2627
rect 623 2621 627 2622
rect 663 2626 667 2627
rect 663 2621 667 2622
rect 839 2626 843 2627
rect 839 2621 843 2622
rect 1023 2626 1027 2627
rect 1023 2621 1027 2622
rect 1215 2626 1219 2627
rect 1215 2621 1219 2622
rect 1407 2626 1411 2627
rect 1407 2621 1411 2622
rect 1607 2626 1611 2627
rect 1607 2621 1611 2622
rect 1823 2626 1827 2627
rect 1864 2623 1866 2651
rect 1950 2643 1956 2644
rect 1950 2639 1951 2643
rect 1955 2639 1956 2643
rect 1950 2638 1956 2639
rect 2062 2643 2068 2644
rect 2062 2639 2063 2643
rect 2067 2639 2068 2643
rect 2062 2638 2068 2639
rect 2174 2643 2180 2644
rect 2174 2639 2175 2643
rect 2179 2639 2180 2643
rect 2174 2638 2180 2639
rect 2294 2643 2300 2644
rect 2294 2639 2295 2643
rect 2299 2639 2300 2643
rect 2294 2638 2300 2639
rect 2414 2643 2420 2644
rect 2414 2639 2415 2643
rect 2419 2639 2420 2643
rect 2414 2638 2420 2639
rect 2526 2643 2532 2644
rect 2526 2639 2527 2643
rect 2531 2639 2532 2643
rect 2526 2638 2532 2639
rect 2638 2643 2644 2644
rect 2638 2639 2639 2643
rect 2643 2639 2644 2643
rect 2638 2638 2644 2639
rect 2742 2643 2748 2644
rect 2742 2639 2743 2643
rect 2747 2639 2748 2643
rect 2742 2638 2748 2639
rect 2854 2643 2860 2644
rect 2854 2639 2855 2643
rect 2859 2639 2860 2643
rect 2854 2638 2860 2639
rect 2966 2643 2972 2644
rect 2966 2639 2967 2643
rect 2971 2639 2972 2643
rect 2966 2638 2972 2639
rect 3078 2643 3084 2644
rect 3078 2639 3079 2643
rect 3083 2639 3084 2643
rect 3078 2638 3084 2639
rect 1952 2623 1954 2638
rect 2064 2623 2066 2638
rect 2176 2623 2178 2638
rect 2296 2623 2298 2638
rect 2416 2623 2418 2638
rect 2528 2623 2530 2638
rect 2640 2623 2642 2638
rect 2744 2623 2746 2638
rect 2856 2623 2858 2638
rect 2968 2623 2970 2638
rect 3080 2623 3082 2638
rect 3576 2623 3578 2651
rect 1823 2621 1827 2622
rect 1863 2622 1867 2623
rect 112 2597 114 2621
rect 224 2610 226 2621
rect 352 2610 354 2621
rect 496 2610 498 2621
rect 664 2610 666 2621
rect 840 2610 842 2621
rect 1024 2610 1026 2621
rect 1216 2610 1218 2621
rect 1408 2610 1410 2621
rect 1608 2610 1610 2621
rect 222 2609 228 2610
rect 222 2605 223 2609
rect 227 2605 228 2609
rect 222 2604 228 2605
rect 350 2609 356 2610
rect 350 2605 351 2609
rect 355 2605 356 2609
rect 350 2604 356 2605
rect 494 2609 500 2610
rect 494 2605 495 2609
rect 499 2605 500 2609
rect 494 2604 500 2605
rect 662 2609 668 2610
rect 662 2605 663 2609
rect 667 2605 668 2609
rect 662 2604 668 2605
rect 838 2609 844 2610
rect 838 2605 839 2609
rect 843 2605 844 2609
rect 838 2604 844 2605
rect 1022 2609 1028 2610
rect 1022 2605 1023 2609
rect 1027 2605 1028 2609
rect 1022 2604 1028 2605
rect 1214 2609 1220 2610
rect 1214 2605 1215 2609
rect 1219 2605 1220 2609
rect 1214 2604 1220 2605
rect 1406 2609 1412 2610
rect 1406 2605 1407 2609
rect 1411 2605 1412 2609
rect 1406 2604 1412 2605
rect 1606 2609 1612 2610
rect 1606 2605 1607 2609
rect 1611 2605 1612 2609
rect 1606 2604 1612 2605
rect 1824 2597 1826 2621
rect 1863 2617 1867 2618
rect 1895 2622 1899 2623
rect 1895 2617 1899 2618
rect 1951 2622 1955 2623
rect 1951 2617 1955 2618
rect 2063 2622 2067 2623
rect 2063 2617 2067 2618
rect 2071 2622 2075 2623
rect 2071 2617 2075 2618
rect 2175 2622 2179 2623
rect 2175 2617 2179 2618
rect 2263 2622 2267 2623
rect 2263 2617 2267 2618
rect 2295 2622 2299 2623
rect 2295 2617 2299 2618
rect 2415 2622 2419 2623
rect 2415 2617 2419 2618
rect 2463 2622 2467 2623
rect 2463 2617 2467 2618
rect 2527 2622 2531 2623
rect 2527 2617 2531 2618
rect 2639 2622 2643 2623
rect 2639 2617 2643 2618
rect 2663 2622 2667 2623
rect 2663 2617 2667 2618
rect 2743 2622 2747 2623
rect 2743 2617 2747 2618
rect 2855 2622 2859 2623
rect 2855 2617 2859 2618
rect 2871 2622 2875 2623
rect 2871 2617 2875 2618
rect 2967 2622 2971 2623
rect 2967 2617 2971 2618
rect 3079 2622 3083 2623
rect 3079 2617 3083 2618
rect 3295 2622 3299 2623
rect 3295 2617 3299 2618
rect 3487 2622 3491 2623
rect 3487 2617 3491 2618
rect 3575 2622 3579 2623
rect 3575 2617 3579 2618
rect 110 2596 116 2597
rect 110 2592 111 2596
rect 115 2592 116 2596
rect 110 2591 116 2592
rect 1822 2596 1828 2597
rect 1822 2592 1823 2596
rect 1827 2592 1828 2596
rect 1864 2593 1866 2617
rect 1896 2606 1898 2617
rect 2072 2606 2074 2617
rect 2264 2606 2266 2617
rect 2464 2606 2466 2617
rect 2664 2606 2666 2617
rect 2872 2606 2874 2617
rect 3080 2606 3082 2617
rect 3296 2606 3298 2617
rect 3488 2606 3490 2617
rect 1894 2605 1900 2606
rect 1894 2601 1895 2605
rect 1899 2601 1900 2605
rect 1894 2600 1900 2601
rect 2070 2605 2076 2606
rect 2070 2601 2071 2605
rect 2075 2601 2076 2605
rect 2070 2600 2076 2601
rect 2262 2605 2268 2606
rect 2262 2601 2263 2605
rect 2267 2601 2268 2605
rect 2262 2600 2268 2601
rect 2462 2605 2468 2606
rect 2462 2601 2463 2605
rect 2467 2601 2468 2605
rect 2462 2600 2468 2601
rect 2662 2605 2668 2606
rect 2662 2601 2663 2605
rect 2667 2601 2668 2605
rect 2662 2600 2668 2601
rect 2870 2605 2876 2606
rect 2870 2601 2871 2605
rect 2875 2601 2876 2605
rect 2870 2600 2876 2601
rect 3078 2605 3084 2606
rect 3078 2601 3079 2605
rect 3083 2601 3084 2605
rect 3078 2600 3084 2601
rect 3294 2605 3300 2606
rect 3294 2601 3295 2605
rect 3299 2601 3300 2605
rect 3294 2600 3300 2601
rect 3486 2605 3492 2606
rect 3486 2601 3487 2605
rect 3491 2601 3492 2605
rect 3486 2600 3492 2601
rect 3576 2593 3578 2617
rect 1822 2591 1828 2592
rect 1862 2592 1868 2593
rect 1862 2588 1863 2592
rect 1867 2588 1868 2592
rect 1862 2587 1868 2588
rect 3574 2592 3580 2593
rect 3574 2588 3575 2592
rect 3579 2588 3580 2592
rect 3574 2587 3580 2588
rect 110 2579 116 2580
rect 110 2575 111 2579
rect 115 2575 116 2579
rect 110 2574 116 2575
rect 1822 2579 1828 2580
rect 1822 2575 1823 2579
rect 1827 2575 1828 2579
rect 1822 2574 1828 2575
rect 1862 2575 1868 2576
rect 112 2559 114 2574
rect 214 2569 220 2570
rect 214 2565 215 2569
rect 219 2565 220 2569
rect 214 2564 220 2565
rect 342 2569 348 2570
rect 342 2565 343 2569
rect 347 2565 348 2569
rect 342 2564 348 2565
rect 486 2569 492 2570
rect 486 2565 487 2569
rect 491 2565 492 2569
rect 486 2564 492 2565
rect 654 2569 660 2570
rect 654 2565 655 2569
rect 659 2565 660 2569
rect 654 2564 660 2565
rect 830 2569 836 2570
rect 830 2565 831 2569
rect 835 2565 836 2569
rect 830 2564 836 2565
rect 1014 2569 1020 2570
rect 1014 2565 1015 2569
rect 1019 2565 1020 2569
rect 1014 2564 1020 2565
rect 1206 2569 1212 2570
rect 1206 2565 1207 2569
rect 1211 2565 1212 2569
rect 1206 2564 1212 2565
rect 1398 2569 1404 2570
rect 1398 2565 1399 2569
rect 1403 2565 1404 2569
rect 1398 2564 1404 2565
rect 1598 2569 1604 2570
rect 1598 2565 1599 2569
rect 1603 2565 1604 2569
rect 1598 2564 1604 2565
rect 216 2559 218 2564
rect 344 2559 346 2564
rect 488 2559 490 2564
rect 656 2559 658 2564
rect 832 2559 834 2564
rect 1016 2559 1018 2564
rect 1208 2559 1210 2564
rect 1400 2559 1402 2564
rect 1600 2559 1602 2564
rect 1824 2559 1826 2574
rect 1862 2571 1863 2575
rect 1867 2571 1868 2575
rect 1862 2570 1868 2571
rect 3574 2575 3580 2576
rect 3574 2571 3575 2575
rect 3579 2571 3580 2575
rect 3574 2570 3580 2571
rect 111 2558 115 2559
rect 111 2553 115 2554
rect 215 2558 219 2559
rect 215 2553 219 2554
rect 271 2558 275 2559
rect 271 2553 275 2554
rect 343 2558 347 2559
rect 343 2553 347 2554
rect 471 2558 475 2559
rect 471 2553 475 2554
rect 487 2558 491 2559
rect 487 2553 491 2554
rect 655 2558 659 2559
rect 655 2553 659 2554
rect 671 2558 675 2559
rect 671 2553 675 2554
rect 831 2558 835 2559
rect 831 2553 835 2554
rect 855 2558 859 2559
rect 855 2553 859 2554
rect 1015 2558 1019 2559
rect 1015 2553 1019 2554
rect 1023 2558 1027 2559
rect 1023 2553 1027 2554
rect 1175 2558 1179 2559
rect 1175 2553 1179 2554
rect 1207 2558 1211 2559
rect 1207 2553 1211 2554
rect 1319 2558 1323 2559
rect 1319 2553 1323 2554
rect 1399 2558 1403 2559
rect 1399 2553 1403 2554
rect 1455 2558 1459 2559
rect 1455 2553 1459 2554
rect 1591 2558 1595 2559
rect 1591 2553 1595 2554
rect 1599 2558 1603 2559
rect 1599 2553 1603 2554
rect 1727 2558 1731 2559
rect 1727 2553 1731 2554
rect 1823 2558 1827 2559
rect 1864 2555 1866 2570
rect 1886 2565 1892 2566
rect 1886 2561 1887 2565
rect 1891 2561 1892 2565
rect 1886 2560 1892 2561
rect 2062 2565 2068 2566
rect 2062 2561 2063 2565
rect 2067 2561 2068 2565
rect 2062 2560 2068 2561
rect 2254 2565 2260 2566
rect 2254 2561 2255 2565
rect 2259 2561 2260 2565
rect 2254 2560 2260 2561
rect 2454 2565 2460 2566
rect 2454 2561 2455 2565
rect 2459 2561 2460 2565
rect 2454 2560 2460 2561
rect 2654 2565 2660 2566
rect 2654 2561 2655 2565
rect 2659 2561 2660 2565
rect 2654 2560 2660 2561
rect 2862 2565 2868 2566
rect 2862 2561 2863 2565
rect 2867 2561 2868 2565
rect 2862 2560 2868 2561
rect 3070 2565 3076 2566
rect 3070 2561 3071 2565
rect 3075 2561 3076 2565
rect 3070 2560 3076 2561
rect 3286 2565 3292 2566
rect 3286 2561 3287 2565
rect 3291 2561 3292 2565
rect 3286 2560 3292 2561
rect 3478 2565 3484 2566
rect 3478 2561 3479 2565
rect 3483 2561 3484 2565
rect 3478 2560 3484 2561
rect 1888 2555 1890 2560
rect 2064 2555 2066 2560
rect 2256 2555 2258 2560
rect 2456 2555 2458 2560
rect 2656 2555 2658 2560
rect 2864 2555 2866 2560
rect 3072 2555 3074 2560
rect 3288 2555 3290 2560
rect 3480 2555 3482 2560
rect 3576 2555 3578 2570
rect 1823 2553 1827 2554
rect 1863 2554 1867 2555
rect 112 2538 114 2553
rect 272 2548 274 2553
rect 472 2548 474 2553
rect 672 2548 674 2553
rect 856 2548 858 2553
rect 1024 2548 1026 2553
rect 1176 2548 1178 2553
rect 1320 2548 1322 2553
rect 1456 2548 1458 2553
rect 1592 2548 1594 2553
rect 1728 2548 1730 2553
rect 270 2547 276 2548
rect 270 2543 271 2547
rect 275 2543 276 2547
rect 270 2542 276 2543
rect 470 2547 476 2548
rect 470 2543 471 2547
rect 475 2543 476 2547
rect 470 2542 476 2543
rect 670 2547 676 2548
rect 670 2543 671 2547
rect 675 2543 676 2547
rect 670 2542 676 2543
rect 854 2547 860 2548
rect 854 2543 855 2547
rect 859 2543 860 2547
rect 854 2542 860 2543
rect 1022 2547 1028 2548
rect 1022 2543 1023 2547
rect 1027 2543 1028 2547
rect 1022 2542 1028 2543
rect 1174 2547 1180 2548
rect 1174 2543 1175 2547
rect 1179 2543 1180 2547
rect 1174 2542 1180 2543
rect 1318 2547 1324 2548
rect 1318 2543 1319 2547
rect 1323 2543 1324 2547
rect 1318 2542 1324 2543
rect 1454 2547 1460 2548
rect 1454 2543 1455 2547
rect 1459 2543 1460 2547
rect 1454 2542 1460 2543
rect 1590 2547 1596 2548
rect 1590 2543 1591 2547
rect 1595 2543 1596 2547
rect 1590 2542 1596 2543
rect 1726 2547 1732 2548
rect 1726 2543 1727 2547
rect 1731 2543 1732 2547
rect 1726 2542 1732 2543
rect 1824 2538 1826 2553
rect 1863 2549 1867 2550
rect 1887 2554 1891 2555
rect 1887 2549 1891 2550
rect 2039 2554 2043 2555
rect 2039 2549 2043 2550
rect 2063 2554 2067 2555
rect 2063 2549 2067 2550
rect 2215 2554 2219 2555
rect 2215 2549 2219 2550
rect 2255 2554 2259 2555
rect 2255 2549 2259 2550
rect 2399 2554 2403 2555
rect 2399 2549 2403 2550
rect 2455 2554 2459 2555
rect 2455 2549 2459 2550
rect 2575 2554 2579 2555
rect 2575 2549 2579 2550
rect 2655 2554 2659 2555
rect 2655 2549 2659 2550
rect 2743 2554 2747 2555
rect 2743 2549 2747 2550
rect 2863 2554 2867 2555
rect 2863 2549 2867 2550
rect 2903 2554 2907 2555
rect 2903 2549 2907 2550
rect 3055 2554 3059 2555
rect 3055 2549 3059 2550
rect 3071 2554 3075 2555
rect 3071 2549 3075 2550
rect 3199 2554 3203 2555
rect 3199 2549 3203 2550
rect 3287 2554 3291 2555
rect 3287 2549 3291 2550
rect 3343 2554 3347 2555
rect 3343 2549 3347 2550
rect 3479 2554 3483 2555
rect 3479 2549 3483 2550
rect 3575 2554 3579 2555
rect 3575 2549 3579 2550
rect 110 2537 116 2538
rect 110 2533 111 2537
rect 115 2533 116 2537
rect 110 2532 116 2533
rect 1822 2537 1828 2538
rect 1822 2533 1823 2537
rect 1827 2533 1828 2537
rect 1864 2534 1866 2549
rect 1888 2544 1890 2549
rect 2040 2544 2042 2549
rect 2216 2544 2218 2549
rect 2400 2544 2402 2549
rect 2576 2544 2578 2549
rect 2744 2544 2746 2549
rect 2904 2544 2906 2549
rect 3056 2544 3058 2549
rect 3200 2544 3202 2549
rect 3344 2544 3346 2549
rect 3480 2544 3482 2549
rect 1886 2543 1892 2544
rect 1886 2539 1887 2543
rect 1891 2539 1892 2543
rect 1886 2538 1892 2539
rect 2038 2543 2044 2544
rect 2038 2539 2039 2543
rect 2043 2539 2044 2543
rect 2038 2538 2044 2539
rect 2214 2543 2220 2544
rect 2214 2539 2215 2543
rect 2219 2539 2220 2543
rect 2214 2538 2220 2539
rect 2398 2543 2404 2544
rect 2398 2539 2399 2543
rect 2403 2539 2404 2543
rect 2398 2538 2404 2539
rect 2574 2543 2580 2544
rect 2574 2539 2575 2543
rect 2579 2539 2580 2543
rect 2574 2538 2580 2539
rect 2742 2543 2748 2544
rect 2742 2539 2743 2543
rect 2747 2539 2748 2543
rect 2742 2538 2748 2539
rect 2902 2543 2908 2544
rect 2902 2539 2903 2543
rect 2907 2539 2908 2543
rect 2902 2538 2908 2539
rect 3054 2543 3060 2544
rect 3054 2539 3055 2543
rect 3059 2539 3060 2543
rect 3054 2538 3060 2539
rect 3198 2543 3204 2544
rect 3198 2539 3199 2543
rect 3203 2539 3204 2543
rect 3198 2538 3204 2539
rect 3342 2543 3348 2544
rect 3342 2539 3343 2543
rect 3347 2539 3348 2543
rect 3342 2538 3348 2539
rect 3478 2543 3484 2544
rect 3478 2539 3479 2543
rect 3483 2539 3484 2543
rect 3478 2538 3484 2539
rect 3576 2534 3578 2549
rect 1822 2532 1828 2533
rect 1862 2533 1868 2534
rect 1862 2529 1863 2533
rect 1867 2529 1868 2533
rect 1862 2528 1868 2529
rect 3574 2533 3580 2534
rect 3574 2529 3575 2533
rect 3579 2529 3580 2533
rect 3574 2528 3580 2529
rect 110 2520 116 2521
rect 110 2516 111 2520
rect 115 2516 116 2520
rect 110 2515 116 2516
rect 1822 2520 1828 2521
rect 1822 2516 1823 2520
rect 1827 2516 1828 2520
rect 1822 2515 1828 2516
rect 1862 2516 1868 2517
rect 112 2487 114 2515
rect 278 2507 284 2508
rect 278 2503 279 2507
rect 283 2503 284 2507
rect 278 2502 284 2503
rect 478 2507 484 2508
rect 478 2503 479 2507
rect 483 2503 484 2507
rect 478 2502 484 2503
rect 678 2507 684 2508
rect 678 2503 679 2507
rect 683 2503 684 2507
rect 678 2502 684 2503
rect 862 2507 868 2508
rect 862 2503 863 2507
rect 867 2503 868 2507
rect 862 2502 868 2503
rect 1030 2507 1036 2508
rect 1030 2503 1031 2507
rect 1035 2503 1036 2507
rect 1030 2502 1036 2503
rect 1182 2507 1188 2508
rect 1182 2503 1183 2507
rect 1187 2503 1188 2507
rect 1182 2502 1188 2503
rect 1326 2507 1332 2508
rect 1326 2503 1327 2507
rect 1331 2503 1332 2507
rect 1326 2502 1332 2503
rect 1462 2507 1468 2508
rect 1462 2503 1463 2507
rect 1467 2503 1468 2507
rect 1462 2502 1468 2503
rect 1598 2507 1604 2508
rect 1598 2503 1599 2507
rect 1603 2503 1604 2507
rect 1598 2502 1604 2503
rect 1734 2507 1740 2508
rect 1734 2503 1735 2507
rect 1739 2503 1740 2507
rect 1734 2502 1740 2503
rect 280 2487 282 2502
rect 480 2487 482 2502
rect 680 2487 682 2502
rect 864 2487 866 2502
rect 1032 2487 1034 2502
rect 1184 2487 1186 2502
rect 1328 2487 1330 2502
rect 1464 2487 1466 2502
rect 1600 2487 1602 2502
rect 1736 2487 1738 2502
rect 1824 2487 1826 2515
rect 1862 2512 1863 2516
rect 1867 2512 1868 2516
rect 1862 2511 1868 2512
rect 3574 2516 3580 2517
rect 3574 2512 3575 2516
rect 3579 2512 3580 2516
rect 3574 2511 3580 2512
rect 1864 2487 1866 2511
rect 1894 2503 1900 2504
rect 1894 2499 1895 2503
rect 1899 2499 1900 2503
rect 1894 2498 1900 2499
rect 2046 2503 2052 2504
rect 2046 2499 2047 2503
rect 2051 2499 2052 2503
rect 2046 2498 2052 2499
rect 2222 2503 2228 2504
rect 2222 2499 2223 2503
rect 2227 2499 2228 2503
rect 2222 2498 2228 2499
rect 2406 2503 2412 2504
rect 2406 2499 2407 2503
rect 2411 2499 2412 2503
rect 2406 2498 2412 2499
rect 2582 2503 2588 2504
rect 2582 2499 2583 2503
rect 2587 2499 2588 2503
rect 2582 2498 2588 2499
rect 2750 2503 2756 2504
rect 2750 2499 2751 2503
rect 2755 2499 2756 2503
rect 2750 2498 2756 2499
rect 2910 2503 2916 2504
rect 2910 2499 2911 2503
rect 2915 2499 2916 2503
rect 2910 2498 2916 2499
rect 3062 2503 3068 2504
rect 3062 2499 3063 2503
rect 3067 2499 3068 2503
rect 3062 2498 3068 2499
rect 3206 2503 3212 2504
rect 3206 2499 3207 2503
rect 3211 2499 3212 2503
rect 3206 2498 3212 2499
rect 3350 2503 3356 2504
rect 3350 2499 3351 2503
rect 3355 2499 3356 2503
rect 3350 2498 3356 2499
rect 3486 2503 3492 2504
rect 3486 2499 3487 2503
rect 3491 2499 3492 2503
rect 3486 2498 3492 2499
rect 1896 2487 1898 2498
rect 2048 2487 2050 2498
rect 2224 2487 2226 2498
rect 2408 2487 2410 2498
rect 2584 2487 2586 2498
rect 2752 2487 2754 2498
rect 2912 2487 2914 2498
rect 3064 2487 3066 2498
rect 3208 2487 3210 2498
rect 3352 2487 3354 2498
rect 3488 2487 3490 2498
rect 3576 2487 3578 2511
rect 111 2486 115 2487
rect 111 2481 115 2482
rect 183 2486 187 2487
rect 183 2481 187 2482
rect 279 2486 283 2487
rect 279 2481 283 2482
rect 319 2486 323 2487
rect 319 2481 323 2482
rect 463 2486 467 2487
rect 463 2481 467 2482
rect 479 2486 483 2487
rect 479 2481 483 2482
rect 607 2486 611 2487
rect 607 2481 611 2482
rect 679 2486 683 2487
rect 679 2481 683 2482
rect 743 2486 747 2487
rect 743 2481 747 2482
rect 863 2486 867 2487
rect 863 2481 867 2482
rect 879 2486 883 2487
rect 879 2481 883 2482
rect 1007 2486 1011 2487
rect 1007 2481 1011 2482
rect 1031 2486 1035 2487
rect 1031 2481 1035 2482
rect 1127 2486 1131 2487
rect 1127 2481 1131 2482
rect 1183 2486 1187 2487
rect 1183 2481 1187 2482
rect 1239 2486 1243 2487
rect 1239 2481 1243 2482
rect 1327 2486 1331 2487
rect 1327 2481 1331 2482
rect 1343 2486 1347 2487
rect 1343 2481 1347 2482
rect 1447 2486 1451 2487
rect 1447 2481 1451 2482
rect 1463 2486 1467 2487
rect 1463 2481 1467 2482
rect 1551 2486 1555 2487
rect 1551 2481 1555 2482
rect 1599 2486 1603 2487
rect 1599 2481 1603 2482
rect 1647 2486 1651 2487
rect 1647 2481 1651 2482
rect 1735 2486 1739 2487
rect 1735 2481 1739 2482
rect 1823 2486 1827 2487
rect 1823 2481 1827 2482
rect 1863 2486 1867 2487
rect 1863 2481 1867 2482
rect 1895 2486 1899 2487
rect 1895 2481 1899 2482
rect 1991 2486 1995 2487
rect 1991 2481 1995 2482
rect 2047 2486 2051 2487
rect 2047 2481 2051 2482
rect 2127 2486 2131 2487
rect 2127 2481 2131 2482
rect 2223 2486 2227 2487
rect 2223 2481 2227 2482
rect 2279 2486 2283 2487
rect 2279 2481 2283 2482
rect 2407 2486 2411 2487
rect 2407 2481 2411 2482
rect 2439 2486 2443 2487
rect 2439 2481 2443 2482
rect 2583 2486 2587 2487
rect 2583 2481 2587 2482
rect 2599 2486 2603 2487
rect 2599 2481 2603 2482
rect 2751 2486 2755 2487
rect 2751 2481 2755 2482
rect 2767 2486 2771 2487
rect 2767 2481 2771 2482
rect 2911 2486 2915 2487
rect 2911 2481 2915 2482
rect 2943 2486 2947 2487
rect 2943 2481 2947 2482
rect 3063 2486 3067 2487
rect 3063 2481 3067 2482
rect 3119 2486 3123 2487
rect 3119 2481 3123 2482
rect 3207 2486 3211 2487
rect 3207 2481 3211 2482
rect 3295 2486 3299 2487
rect 3295 2481 3299 2482
rect 3351 2486 3355 2487
rect 3351 2481 3355 2482
rect 3471 2486 3475 2487
rect 3471 2481 3475 2482
rect 3487 2486 3491 2487
rect 3487 2481 3491 2482
rect 3575 2486 3579 2487
rect 3575 2481 3579 2482
rect 112 2457 114 2481
rect 184 2470 186 2481
rect 320 2470 322 2481
rect 464 2470 466 2481
rect 608 2470 610 2481
rect 744 2470 746 2481
rect 880 2470 882 2481
rect 1008 2470 1010 2481
rect 1128 2470 1130 2481
rect 1240 2470 1242 2481
rect 1344 2470 1346 2481
rect 1448 2470 1450 2481
rect 1552 2470 1554 2481
rect 1648 2470 1650 2481
rect 1736 2470 1738 2481
rect 182 2469 188 2470
rect 182 2465 183 2469
rect 187 2465 188 2469
rect 182 2464 188 2465
rect 318 2469 324 2470
rect 318 2465 319 2469
rect 323 2465 324 2469
rect 318 2464 324 2465
rect 462 2469 468 2470
rect 462 2465 463 2469
rect 467 2465 468 2469
rect 462 2464 468 2465
rect 606 2469 612 2470
rect 606 2465 607 2469
rect 611 2465 612 2469
rect 606 2464 612 2465
rect 742 2469 748 2470
rect 742 2465 743 2469
rect 747 2465 748 2469
rect 742 2464 748 2465
rect 878 2469 884 2470
rect 878 2465 879 2469
rect 883 2465 884 2469
rect 878 2464 884 2465
rect 1006 2469 1012 2470
rect 1006 2465 1007 2469
rect 1011 2465 1012 2469
rect 1006 2464 1012 2465
rect 1126 2469 1132 2470
rect 1126 2465 1127 2469
rect 1131 2465 1132 2469
rect 1126 2464 1132 2465
rect 1238 2469 1244 2470
rect 1238 2465 1239 2469
rect 1243 2465 1244 2469
rect 1238 2464 1244 2465
rect 1342 2469 1348 2470
rect 1342 2465 1343 2469
rect 1347 2465 1348 2469
rect 1342 2464 1348 2465
rect 1446 2469 1452 2470
rect 1446 2465 1447 2469
rect 1451 2465 1452 2469
rect 1446 2464 1452 2465
rect 1550 2469 1556 2470
rect 1550 2465 1551 2469
rect 1555 2465 1556 2469
rect 1550 2464 1556 2465
rect 1646 2469 1652 2470
rect 1646 2465 1647 2469
rect 1651 2465 1652 2469
rect 1646 2464 1652 2465
rect 1734 2469 1740 2470
rect 1734 2465 1735 2469
rect 1739 2465 1740 2469
rect 1734 2464 1740 2465
rect 1824 2457 1826 2481
rect 1864 2457 1866 2481
rect 1896 2470 1898 2481
rect 1992 2470 1994 2481
rect 2128 2470 2130 2481
rect 2280 2470 2282 2481
rect 2440 2470 2442 2481
rect 2600 2470 2602 2481
rect 2768 2470 2770 2481
rect 2944 2470 2946 2481
rect 3120 2470 3122 2481
rect 3296 2470 3298 2481
rect 3472 2470 3474 2481
rect 1894 2469 1900 2470
rect 1894 2465 1895 2469
rect 1899 2465 1900 2469
rect 1894 2464 1900 2465
rect 1990 2469 1996 2470
rect 1990 2465 1991 2469
rect 1995 2465 1996 2469
rect 1990 2464 1996 2465
rect 2126 2469 2132 2470
rect 2126 2465 2127 2469
rect 2131 2465 2132 2469
rect 2126 2464 2132 2465
rect 2278 2469 2284 2470
rect 2278 2465 2279 2469
rect 2283 2465 2284 2469
rect 2278 2464 2284 2465
rect 2438 2469 2444 2470
rect 2438 2465 2439 2469
rect 2443 2465 2444 2469
rect 2438 2464 2444 2465
rect 2598 2469 2604 2470
rect 2598 2465 2599 2469
rect 2603 2465 2604 2469
rect 2598 2464 2604 2465
rect 2766 2469 2772 2470
rect 2766 2465 2767 2469
rect 2771 2465 2772 2469
rect 2766 2464 2772 2465
rect 2942 2469 2948 2470
rect 2942 2465 2943 2469
rect 2947 2465 2948 2469
rect 2942 2464 2948 2465
rect 3118 2469 3124 2470
rect 3118 2465 3119 2469
rect 3123 2465 3124 2469
rect 3118 2464 3124 2465
rect 3294 2469 3300 2470
rect 3294 2465 3295 2469
rect 3299 2465 3300 2469
rect 3294 2464 3300 2465
rect 3470 2469 3476 2470
rect 3470 2465 3471 2469
rect 3475 2465 3476 2469
rect 3470 2464 3476 2465
rect 3576 2457 3578 2481
rect 110 2456 116 2457
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 110 2451 116 2452
rect 1822 2456 1828 2457
rect 1822 2452 1823 2456
rect 1827 2452 1828 2456
rect 1822 2451 1828 2452
rect 1862 2456 1868 2457
rect 1862 2452 1863 2456
rect 1867 2452 1868 2456
rect 1862 2451 1868 2452
rect 3574 2456 3580 2457
rect 3574 2452 3575 2456
rect 3579 2452 3580 2456
rect 3574 2451 3580 2452
rect 110 2439 116 2440
rect 110 2435 111 2439
rect 115 2435 116 2439
rect 110 2434 116 2435
rect 1822 2439 1828 2440
rect 1822 2435 1823 2439
rect 1827 2435 1828 2439
rect 1822 2434 1828 2435
rect 1862 2439 1868 2440
rect 1862 2435 1863 2439
rect 1867 2435 1868 2439
rect 1862 2434 1868 2435
rect 3574 2439 3580 2440
rect 3574 2435 3575 2439
rect 3579 2435 3580 2439
rect 3574 2434 3580 2435
rect 112 2411 114 2434
rect 174 2429 180 2430
rect 174 2425 175 2429
rect 179 2425 180 2429
rect 174 2424 180 2425
rect 310 2429 316 2430
rect 310 2425 311 2429
rect 315 2425 316 2429
rect 310 2424 316 2425
rect 454 2429 460 2430
rect 454 2425 455 2429
rect 459 2425 460 2429
rect 454 2424 460 2425
rect 598 2429 604 2430
rect 598 2425 599 2429
rect 603 2425 604 2429
rect 598 2424 604 2425
rect 734 2429 740 2430
rect 734 2425 735 2429
rect 739 2425 740 2429
rect 734 2424 740 2425
rect 870 2429 876 2430
rect 870 2425 871 2429
rect 875 2425 876 2429
rect 870 2424 876 2425
rect 998 2429 1004 2430
rect 998 2425 999 2429
rect 1003 2425 1004 2429
rect 998 2424 1004 2425
rect 1118 2429 1124 2430
rect 1118 2425 1119 2429
rect 1123 2425 1124 2429
rect 1118 2424 1124 2425
rect 1230 2429 1236 2430
rect 1230 2425 1231 2429
rect 1235 2425 1236 2429
rect 1230 2424 1236 2425
rect 1334 2429 1340 2430
rect 1334 2425 1335 2429
rect 1339 2425 1340 2429
rect 1334 2424 1340 2425
rect 1438 2429 1444 2430
rect 1438 2425 1439 2429
rect 1443 2425 1444 2429
rect 1438 2424 1444 2425
rect 1542 2429 1548 2430
rect 1542 2425 1543 2429
rect 1547 2425 1548 2429
rect 1542 2424 1548 2425
rect 1638 2429 1644 2430
rect 1638 2425 1639 2429
rect 1643 2425 1644 2429
rect 1638 2424 1644 2425
rect 1726 2429 1732 2430
rect 1726 2425 1727 2429
rect 1731 2425 1732 2429
rect 1726 2424 1732 2425
rect 176 2411 178 2424
rect 312 2411 314 2424
rect 456 2411 458 2424
rect 600 2411 602 2424
rect 736 2411 738 2424
rect 872 2411 874 2424
rect 1000 2411 1002 2424
rect 1120 2411 1122 2424
rect 1232 2411 1234 2424
rect 1336 2411 1338 2424
rect 1440 2411 1442 2424
rect 1544 2411 1546 2424
rect 1640 2411 1642 2424
rect 1728 2411 1730 2424
rect 1824 2411 1826 2434
rect 1864 2411 1866 2434
rect 1886 2429 1892 2430
rect 1886 2425 1887 2429
rect 1891 2425 1892 2429
rect 1886 2424 1892 2425
rect 1982 2429 1988 2430
rect 1982 2425 1983 2429
rect 1987 2425 1988 2429
rect 1982 2424 1988 2425
rect 2118 2429 2124 2430
rect 2118 2425 2119 2429
rect 2123 2425 2124 2429
rect 2118 2424 2124 2425
rect 2270 2429 2276 2430
rect 2270 2425 2271 2429
rect 2275 2425 2276 2429
rect 2270 2424 2276 2425
rect 2430 2429 2436 2430
rect 2430 2425 2431 2429
rect 2435 2425 2436 2429
rect 2430 2424 2436 2425
rect 2590 2429 2596 2430
rect 2590 2425 2591 2429
rect 2595 2425 2596 2429
rect 2590 2424 2596 2425
rect 2758 2429 2764 2430
rect 2758 2425 2759 2429
rect 2763 2425 2764 2429
rect 2758 2424 2764 2425
rect 2934 2429 2940 2430
rect 2934 2425 2935 2429
rect 2939 2425 2940 2429
rect 2934 2424 2940 2425
rect 3110 2429 3116 2430
rect 3110 2425 3111 2429
rect 3115 2425 3116 2429
rect 3110 2424 3116 2425
rect 3286 2429 3292 2430
rect 3286 2425 3287 2429
rect 3291 2425 3292 2429
rect 3286 2424 3292 2425
rect 3462 2429 3468 2430
rect 3462 2425 3463 2429
rect 3467 2425 3468 2429
rect 3462 2424 3468 2425
rect 1888 2411 1890 2424
rect 1984 2411 1986 2424
rect 2120 2411 2122 2424
rect 2272 2411 2274 2424
rect 2432 2411 2434 2424
rect 2592 2411 2594 2424
rect 2760 2411 2762 2424
rect 2936 2411 2938 2424
rect 3112 2411 3114 2424
rect 3288 2411 3290 2424
rect 3464 2411 3466 2424
rect 3576 2411 3578 2434
rect 111 2410 115 2411
rect 111 2405 115 2406
rect 151 2410 155 2411
rect 151 2405 155 2406
rect 175 2410 179 2411
rect 175 2405 179 2406
rect 311 2410 315 2411
rect 311 2405 315 2406
rect 319 2410 323 2411
rect 319 2405 323 2406
rect 455 2410 459 2411
rect 455 2405 459 2406
rect 479 2410 483 2411
rect 479 2405 483 2406
rect 599 2410 603 2411
rect 599 2405 603 2406
rect 639 2410 643 2411
rect 639 2405 643 2406
rect 735 2410 739 2411
rect 735 2405 739 2406
rect 783 2410 787 2411
rect 783 2405 787 2406
rect 871 2410 875 2411
rect 871 2405 875 2406
rect 919 2410 923 2411
rect 919 2405 923 2406
rect 999 2410 1003 2411
rect 999 2405 1003 2406
rect 1047 2410 1051 2411
rect 1047 2405 1051 2406
rect 1119 2410 1123 2411
rect 1119 2405 1123 2406
rect 1175 2410 1179 2411
rect 1175 2405 1179 2406
rect 1231 2410 1235 2411
rect 1231 2405 1235 2406
rect 1303 2410 1307 2411
rect 1303 2405 1307 2406
rect 1335 2410 1339 2411
rect 1335 2405 1339 2406
rect 1431 2410 1435 2411
rect 1431 2405 1435 2406
rect 1439 2410 1443 2411
rect 1439 2405 1443 2406
rect 1543 2410 1547 2411
rect 1543 2405 1547 2406
rect 1639 2410 1643 2411
rect 1639 2405 1643 2406
rect 1727 2410 1731 2411
rect 1727 2405 1731 2406
rect 1823 2410 1827 2411
rect 1823 2405 1827 2406
rect 1863 2410 1867 2411
rect 1863 2405 1867 2406
rect 1887 2410 1891 2411
rect 1887 2405 1891 2406
rect 1983 2410 1987 2411
rect 1983 2405 1987 2406
rect 2119 2410 2123 2411
rect 2119 2405 2123 2406
rect 2271 2410 2275 2411
rect 2271 2405 2275 2406
rect 2351 2410 2355 2411
rect 2351 2405 2355 2406
rect 2431 2410 2435 2411
rect 2431 2405 2435 2406
rect 2503 2410 2507 2411
rect 2503 2405 2507 2406
rect 2591 2410 2595 2411
rect 2591 2405 2595 2406
rect 2655 2410 2659 2411
rect 2655 2405 2659 2406
rect 2759 2410 2763 2411
rect 2759 2405 2763 2406
rect 2807 2410 2811 2411
rect 2807 2405 2811 2406
rect 2935 2410 2939 2411
rect 2935 2405 2939 2406
rect 2967 2410 2971 2411
rect 2967 2405 2971 2406
rect 3111 2410 3115 2411
rect 3111 2405 3115 2406
rect 3135 2410 3139 2411
rect 3135 2405 3139 2406
rect 3287 2410 3291 2411
rect 3287 2405 3291 2406
rect 3303 2410 3307 2411
rect 3303 2405 3307 2406
rect 3463 2410 3467 2411
rect 3463 2405 3467 2406
rect 3471 2410 3475 2411
rect 3471 2405 3475 2406
rect 3575 2410 3579 2411
rect 3575 2405 3579 2406
rect 112 2390 114 2405
rect 152 2400 154 2405
rect 320 2400 322 2405
rect 480 2400 482 2405
rect 640 2400 642 2405
rect 784 2400 786 2405
rect 920 2400 922 2405
rect 1048 2400 1050 2405
rect 1176 2400 1178 2405
rect 1304 2400 1306 2405
rect 1432 2400 1434 2405
rect 150 2399 156 2400
rect 150 2395 151 2399
rect 155 2395 156 2399
rect 150 2394 156 2395
rect 318 2399 324 2400
rect 318 2395 319 2399
rect 323 2395 324 2399
rect 318 2394 324 2395
rect 478 2399 484 2400
rect 478 2395 479 2399
rect 483 2395 484 2399
rect 478 2394 484 2395
rect 638 2399 644 2400
rect 638 2395 639 2399
rect 643 2395 644 2399
rect 638 2394 644 2395
rect 782 2399 788 2400
rect 782 2395 783 2399
rect 787 2395 788 2399
rect 782 2394 788 2395
rect 918 2399 924 2400
rect 918 2395 919 2399
rect 923 2395 924 2399
rect 918 2394 924 2395
rect 1046 2399 1052 2400
rect 1046 2395 1047 2399
rect 1051 2395 1052 2399
rect 1046 2394 1052 2395
rect 1174 2399 1180 2400
rect 1174 2395 1175 2399
rect 1179 2395 1180 2399
rect 1174 2394 1180 2395
rect 1302 2399 1308 2400
rect 1302 2395 1303 2399
rect 1307 2395 1308 2399
rect 1302 2394 1308 2395
rect 1430 2399 1436 2400
rect 1430 2395 1431 2399
rect 1435 2395 1436 2399
rect 1430 2394 1436 2395
rect 1824 2390 1826 2405
rect 1864 2390 1866 2405
rect 2352 2400 2354 2405
rect 2504 2400 2506 2405
rect 2656 2400 2658 2405
rect 2808 2400 2810 2405
rect 2968 2400 2970 2405
rect 3136 2400 3138 2405
rect 3304 2400 3306 2405
rect 3472 2400 3474 2405
rect 2350 2399 2356 2400
rect 2350 2395 2351 2399
rect 2355 2395 2356 2399
rect 2350 2394 2356 2395
rect 2502 2399 2508 2400
rect 2502 2395 2503 2399
rect 2507 2395 2508 2399
rect 2502 2394 2508 2395
rect 2654 2399 2660 2400
rect 2654 2395 2655 2399
rect 2659 2395 2660 2399
rect 2654 2394 2660 2395
rect 2806 2399 2812 2400
rect 2806 2395 2807 2399
rect 2811 2395 2812 2399
rect 2806 2394 2812 2395
rect 2966 2399 2972 2400
rect 2966 2395 2967 2399
rect 2971 2395 2972 2399
rect 2966 2394 2972 2395
rect 3134 2399 3140 2400
rect 3134 2395 3135 2399
rect 3139 2395 3140 2399
rect 3134 2394 3140 2395
rect 3302 2399 3308 2400
rect 3302 2395 3303 2399
rect 3307 2395 3308 2399
rect 3302 2394 3308 2395
rect 3470 2399 3476 2400
rect 3470 2395 3471 2399
rect 3475 2395 3476 2399
rect 3470 2394 3476 2395
rect 3576 2390 3578 2405
rect 110 2389 116 2390
rect 110 2385 111 2389
rect 115 2385 116 2389
rect 110 2384 116 2385
rect 1822 2389 1828 2390
rect 1822 2385 1823 2389
rect 1827 2385 1828 2389
rect 1822 2384 1828 2385
rect 1862 2389 1868 2390
rect 1862 2385 1863 2389
rect 1867 2385 1868 2389
rect 1862 2384 1868 2385
rect 3574 2389 3580 2390
rect 3574 2385 3575 2389
rect 3579 2385 3580 2389
rect 3574 2384 3580 2385
rect 110 2372 116 2373
rect 110 2368 111 2372
rect 115 2368 116 2372
rect 110 2367 116 2368
rect 1822 2372 1828 2373
rect 1822 2368 1823 2372
rect 1827 2368 1828 2372
rect 1822 2367 1828 2368
rect 1862 2372 1868 2373
rect 1862 2368 1863 2372
rect 1867 2368 1868 2372
rect 1862 2367 1868 2368
rect 3574 2372 3580 2373
rect 3574 2368 3575 2372
rect 3579 2368 3580 2372
rect 3574 2367 3580 2368
rect 112 2339 114 2367
rect 158 2359 164 2360
rect 158 2355 159 2359
rect 163 2355 164 2359
rect 158 2354 164 2355
rect 326 2359 332 2360
rect 326 2355 327 2359
rect 331 2355 332 2359
rect 326 2354 332 2355
rect 486 2359 492 2360
rect 486 2355 487 2359
rect 491 2355 492 2359
rect 486 2354 492 2355
rect 646 2359 652 2360
rect 646 2355 647 2359
rect 651 2355 652 2359
rect 646 2354 652 2355
rect 790 2359 796 2360
rect 790 2355 791 2359
rect 795 2355 796 2359
rect 790 2354 796 2355
rect 926 2359 932 2360
rect 926 2355 927 2359
rect 931 2355 932 2359
rect 926 2354 932 2355
rect 1054 2359 1060 2360
rect 1054 2355 1055 2359
rect 1059 2355 1060 2359
rect 1054 2354 1060 2355
rect 1182 2359 1188 2360
rect 1182 2355 1183 2359
rect 1187 2355 1188 2359
rect 1182 2354 1188 2355
rect 1310 2359 1316 2360
rect 1310 2355 1311 2359
rect 1315 2355 1316 2359
rect 1310 2354 1316 2355
rect 1438 2359 1444 2360
rect 1438 2355 1439 2359
rect 1443 2355 1444 2359
rect 1438 2354 1444 2355
rect 160 2339 162 2354
rect 328 2339 330 2354
rect 488 2339 490 2354
rect 648 2339 650 2354
rect 792 2339 794 2354
rect 928 2339 930 2354
rect 1056 2339 1058 2354
rect 1184 2339 1186 2354
rect 1312 2339 1314 2354
rect 1440 2339 1442 2354
rect 1824 2339 1826 2367
rect 1864 2339 1866 2367
rect 2358 2359 2364 2360
rect 2358 2355 2359 2359
rect 2363 2355 2364 2359
rect 2358 2354 2364 2355
rect 2510 2359 2516 2360
rect 2510 2355 2511 2359
rect 2515 2355 2516 2359
rect 2510 2354 2516 2355
rect 2662 2359 2668 2360
rect 2662 2355 2663 2359
rect 2667 2355 2668 2359
rect 2662 2354 2668 2355
rect 2814 2359 2820 2360
rect 2814 2355 2815 2359
rect 2819 2355 2820 2359
rect 2814 2354 2820 2355
rect 2974 2359 2980 2360
rect 2974 2355 2975 2359
rect 2979 2355 2980 2359
rect 2974 2354 2980 2355
rect 3142 2359 3148 2360
rect 3142 2355 3143 2359
rect 3147 2355 3148 2359
rect 3142 2354 3148 2355
rect 3310 2359 3316 2360
rect 3310 2355 3311 2359
rect 3315 2355 3316 2359
rect 3310 2354 3316 2355
rect 3478 2359 3484 2360
rect 3478 2355 3479 2359
rect 3483 2355 3484 2359
rect 3478 2354 3484 2355
rect 2360 2339 2362 2354
rect 2512 2339 2514 2354
rect 2664 2339 2666 2354
rect 2816 2339 2818 2354
rect 2976 2339 2978 2354
rect 3144 2339 3146 2354
rect 3312 2339 3314 2354
rect 3480 2339 3482 2354
rect 3576 2339 3578 2367
rect 111 2338 115 2339
rect 111 2333 115 2334
rect 143 2338 147 2339
rect 143 2333 147 2334
rect 159 2338 163 2339
rect 159 2333 163 2334
rect 263 2338 267 2339
rect 263 2333 267 2334
rect 327 2338 331 2339
rect 327 2333 331 2334
rect 407 2338 411 2339
rect 407 2333 411 2334
rect 487 2338 491 2339
rect 487 2333 491 2334
rect 543 2338 547 2339
rect 543 2333 547 2334
rect 647 2338 651 2339
rect 647 2333 651 2334
rect 679 2338 683 2339
rect 679 2333 683 2334
rect 791 2338 795 2339
rect 791 2333 795 2334
rect 807 2338 811 2339
rect 807 2333 811 2334
rect 927 2338 931 2339
rect 927 2333 931 2334
rect 1039 2338 1043 2339
rect 1039 2333 1043 2334
rect 1055 2338 1059 2339
rect 1055 2333 1059 2334
rect 1159 2338 1163 2339
rect 1159 2333 1163 2334
rect 1183 2338 1187 2339
rect 1183 2333 1187 2334
rect 1279 2338 1283 2339
rect 1279 2333 1283 2334
rect 1311 2338 1315 2339
rect 1311 2333 1315 2334
rect 1439 2338 1443 2339
rect 1439 2333 1443 2334
rect 1823 2338 1827 2339
rect 1823 2333 1827 2334
rect 1863 2338 1867 2339
rect 1863 2333 1867 2334
rect 2351 2338 2355 2339
rect 2351 2333 2355 2334
rect 2359 2338 2363 2339
rect 2359 2333 2363 2334
rect 2447 2338 2451 2339
rect 2447 2333 2451 2334
rect 2511 2338 2515 2339
rect 2511 2333 2515 2334
rect 2559 2338 2563 2339
rect 2559 2333 2563 2334
rect 2663 2338 2667 2339
rect 2663 2333 2667 2334
rect 2703 2338 2707 2339
rect 2703 2333 2707 2334
rect 2815 2338 2819 2339
rect 2815 2333 2819 2334
rect 2879 2338 2883 2339
rect 2879 2333 2883 2334
rect 2975 2338 2979 2339
rect 2975 2333 2979 2334
rect 3079 2338 3083 2339
rect 3079 2333 3083 2334
rect 3143 2338 3147 2339
rect 3143 2333 3147 2334
rect 3287 2338 3291 2339
rect 3287 2333 3291 2334
rect 3311 2338 3315 2339
rect 3311 2333 3315 2334
rect 3479 2338 3483 2339
rect 3479 2333 3483 2334
rect 3487 2338 3491 2339
rect 3487 2333 3491 2334
rect 3575 2338 3579 2339
rect 3575 2333 3579 2334
rect 112 2309 114 2333
rect 144 2322 146 2333
rect 264 2322 266 2333
rect 408 2322 410 2333
rect 544 2322 546 2333
rect 680 2322 682 2333
rect 808 2322 810 2333
rect 928 2322 930 2333
rect 1040 2322 1042 2333
rect 1160 2322 1162 2333
rect 1280 2322 1282 2333
rect 142 2321 148 2322
rect 142 2317 143 2321
rect 147 2317 148 2321
rect 142 2316 148 2317
rect 262 2321 268 2322
rect 262 2317 263 2321
rect 267 2317 268 2321
rect 262 2316 268 2317
rect 406 2321 412 2322
rect 406 2317 407 2321
rect 411 2317 412 2321
rect 406 2316 412 2317
rect 542 2321 548 2322
rect 542 2317 543 2321
rect 547 2317 548 2321
rect 542 2316 548 2317
rect 678 2321 684 2322
rect 678 2317 679 2321
rect 683 2317 684 2321
rect 678 2316 684 2317
rect 806 2321 812 2322
rect 806 2317 807 2321
rect 811 2317 812 2321
rect 806 2316 812 2317
rect 926 2321 932 2322
rect 926 2317 927 2321
rect 931 2317 932 2321
rect 926 2316 932 2317
rect 1038 2321 1044 2322
rect 1038 2317 1039 2321
rect 1043 2317 1044 2321
rect 1038 2316 1044 2317
rect 1158 2321 1164 2322
rect 1158 2317 1159 2321
rect 1163 2317 1164 2321
rect 1158 2316 1164 2317
rect 1278 2321 1284 2322
rect 1278 2317 1279 2321
rect 1283 2317 1284 2321
rect 1278 2316 1284 2317
rect 1824 2309 1826 2333
rect 1864 2309 1866 2333
rect 2352 2322 2354 2333
rect 2448 2322 2450 2333
rect 2560 2322 2562 2333
rect 2704 2322 2706 2333
rect 2880 2322 2882 2333
rect 3080 2322 3082 2333
rect 3288 2322 3290 2333
rect 3488 2322 3490 2333
rect 2350 2321 2356 2322
rect 2350 2317 2351 2321
rect 2355 2317 2356 2321
rect 2350 2316 2356 2317
rect 2446 2321 2452 2322
rect 2446 2317 2447 2321
rect 2451 2317 2452 2321
rect 2446 2316 2452 2317
rect 2558 2321 2564 2322
rect 2558 2317 2559 2321
rect 2563 2317 2564 2321
rect 2558 2316 2564 2317
rect 2702 2321 2708 2322
rect 2702 2317 2703 2321
rect 2707 2317 2708 2321
rect 2702 2316 2708 2317
rect 2878 2321 2884 2322
rect 2878 2317 2879 2321
rect 2883 2317 2884 2321
rect 2878 2316 2884 2317
rect 3078 2321 3084 2322
rect 3078 2317 3079 2321
rect 3083 2317 3084 2321
rect 3078 2316 3084 2317
rect 3286 2321 3292 2322
rect 3286 2317 3287 2321
rect 3291 2317 3292 2321
rect 3286 2316 3292 2317
rect 3486 2321 3492 2322
rect 3486 2317 3487 2321
rect 3491 2317 3492 2321
rect 3486 2316 3492 2317
rect 3576 2309 3578 2333
rect 110 2308 116 2309
rect 110 2304 111 2308
rect 115 2304 116 2308
rect 110 2303 116 2304
rect 1822 2308 1828 2309
rect 1822 2304 1823 2308
rect 1827 2304 1828 2308
rect 1822 2303 1828 2304
rect 1862 2308 1868 2309
rect 1862 2304 1863 2308
rect 1867 2304 1868 2308
rect 1862 2303 1868 2304
rect 3574 2308 3580 2309
rect 3574 2304 3575 2308
rect 3579 2304 3580 2308
rect 3574 2303 3580 2304
rect 110 2291 116 2292
rect 110 2287 111 2291
rect 115 2287 116 2291
rect 110 2286 116 2287
rect 1822 2291 1828 2292
rect 1822 2287 1823 2291
rect 1827 2287 1828 2291
rect 1822 2286 1828 2287
rect 1862 2291 1868 2292
rect 1862 2287 1863 2291
rect 1867 2287 1868 2291
rect 1862 2286 1868 2287
rect 3574 2291 3580 2292
rect 3574 2287 3575 2291
rect 3579 2287 3580 2291
rect 3574 2286 3580 2287
rect 112 2271 114 2286
rect 134 2281 140 2282
rect 134 2277 135 2281
rect 139 2277 140 2281
rect 134 2276 140 2277
rect 254 2281 260 2282
rect 254 2277 255 2281
rect 259 2277 260 2281
rect 254 2276 260 2277
rect 398 2281 404 2282
rect 398 2277 399 2281
rect 403 2277 404 2281
rect 398 2276 404 2277
rect 534 2281 540 2282
rect 534 2277 535 2281
rect 539 2277 540 2281
rect 534 2276 540 2277
rect 670 2281 676 2282
rect 670 2277 671 2281
rect 675 2277 676 2281
rect 670 2276 676 2277
rect 798 2281 804 2282
rect 798 2277 799 2281
rect 803 2277 804 2281
rect 798 2276 804 2277
rect 918 2281 924 2282
rect 918 2277 919 2281
rect 923 2277 924 2281
rect 918 2276 924 2277
rect 1030 2281 1036 2282
rect 1030 2277 1031 2281
rect 1035 2277 1036 2281
rect 1030 2276 1036 2277
rect 1150 2281 1156 2282
rect 1150 2277 1151 2281
rect 1155 2277 1156 2281
rect 1150 2276 1156 2277
rect 1270 2281 1276 2282
rect 1270 2277 1271 2281
rect 1275 2277 1276 2281
rect 1270 2276 1276 2277
rect 136 2271 138 2276
rect 256 2271 258 2276
rect 400 2271 402 2276
rect 536 2271 538 2276
rect 672 2271 674 2276
rect 800 2271 802 2276
rect 920 2271 922 2276
rect 1032 2271 1034 2276
rect 1152 2271 1154 2276
rect 1272 2271 1274 2276
rect 1824 2271 1826 2286
rect 1864 2271 1866 2286
rect 2342 2281 2348 2282
rect 2342 2277 2343 2281
rect 2347 2277 2348 2281
rect 2342 2276 2348 2277
rect 2438 2281 2444 2282
rect 2438 2277 2439 2281
rect 2443 2277 2444 2281
rect 2438 2276 2444 2277
rect 2550 2281 2556 2282
rect 2550 2277 2551 2281
rect 2555 2277 2556 2281
rect 2550 2276 2556 2277
rect 2694 2281 2700 2282
rect 2694 2277 2695 2281
rect 2699 2277 2700 2281
rect 2694 2276 2700 2277
rect 2870 2281 2876 2282
rect 2870 2277 2871 2281
rect 2875 2277 2876 2281
rect 2870 2276 2876 2277
rect 3070 2281 3076 2282
rect 3070 2277 3071 2281
rect 3075 2277 3076 2281
rect 3070 2276 3076 2277
rect 3278 2281 3284 2282
rect 3278 2277 3279 2281
rect 3283 2277 3284 2281
rect 3278 2276 3284 2277
rect 3478 2281 3484 2282
rect 3478 2277 3479 2281
rect 3483 2277 3484 2281
rect 3478 2276 3484 2277
rect 2344 2271 2346 2276
rect 2440 2271 2442 2276
rect 2552 2271 2554 2276
rect 2696 2271 2698 2276
rect 2872 2271 2874 2276
rect 3072 2271 3074 2276
rect 3280 2271 3282 2276
rect 3480 2271 3482 2276
rect 3576 2271 3578 2286
rect 111 2270 115 2271
rect 111 2265 115 2266
rect 135 2270 139 2271
rect 135 2265 139 2266
rect 231 2270 235 2271
rect 231 2265 235 2266
rect 255 2270 259 2271
rect 255 2265 259 2266
rect 351 2270 355 2271
rect 351 2265 355 2266
rect 399 2270 403 2271
rect 399 2265 403 2266
rect 471 2270 475 2271
rect 471 2265 475 2266
rect 535 2270 539 2271
rect 535 2265 539 2266
rect 591 2270 595 2271
rect 591 2265 595 2266
rect 671 2270 675 2271
rect 671 2265 675 2266
rect 711 2270 715 2271
rect 711 2265 715 2266
rect 799 2270 803 2271
rect 799 2265 803 2266
rect 823 2270 827 2271
rect 823 2265 827 2266
rect 919 2270 923 2271
rect 919 2265 923 2266
rect 935 2270 939 2271
rect 935 2265 939 2266
rect 1031 2270 1035 2271
rect 1031 2265 1035 2266
rect 1055 2270 1059 2271
rect 1055 2265 1059 2266
rect 1151 2270 1155 2271
rect 1151 2265 1155 2266
rect 1175 2270 1179 2271
rect 1175 2265 1179 2266
rect 1271 2270 1275 2271
rect 1271 2265 1275 2266
rect 1823 2270 1827 2271
rect 1823 2265 1827 2266
rect 1863 2270 1867 2271
rect 1863 2265 1867 2266
rect 2335 2270 2339 2271
rect 2335 2265 2339 2266
rect 2343 2270 2347 2271
rect 2343 2265 2347 2266
rect 2439 2270 2443 2271
rect 2439 2265 2443 2266
rect 2447 2270 2451 2271
rect 2447 2265 2451 2266
rect 2551 2270 2555 2271
rect 2551 2265 2555 2266
rect 2583 2270 2587 2271
rect 2583 2265 2587 2266
rect 2695 2270 2699 2271
rect 2695 2265 2699 2266
rect 2735 2270 2739 2271
rect 2735 2265 2739 2266
rect 2871 2270 2875 2271
rect 2871 2265 2875 2266
rect 2911 2270 2915 2271
rect 2911 2265 2915 2266
rect 3071 2270 3075 2271
rect 3071 2265 3075 2266
rect 3103 2270 3107 2271
rect 3103 2265 3107 2266
rect 3279 2270 3283 2271
rect 3279 2265 3283 2266
rect 3303 2270 3307 2271
rect 3303 2265 3307 2266
rect 3479 2270 3483 2271
rect 3479 2265 3483 2266
rect 3575 2270 3579 2271
rect 3575 2265 3579 2266
rect 112 2250 114 2265
rect 136 2260 138 2265
rect 232 2260 234 2265
rect 352 2260 354 2265
rect 472 2260 474 2265
rect 592 2260 594 2265
rect 712 2260 714 2265
rect 824 2260 826 2265
rect 936 2260 938 2265
rect 1056 2260 1058 2265
rect 1176 2260 1178 2265
rect 134 2259 140 2260
rect 134 2255 135 2259
rect 139 2255 140 2259
rect 134 2254 140 2255
rect 230 2259 236 2260
rect 230 2255 231 2259
rect 235 2255 236 2259
rect 230 2254 236 2255
rect 350 2259 356 2260
rect 350 2255 351 2259
rect 355 2255 356 2259
rect 350 2254 356 2255
rect 470 2259 476 2260
rect 470 2255 471 2259
rect 475 2255 476 2259
rect 470 2254 476 2255
rect 590 2259 596 2260
rect 590 2255 591 2259
rect 595 2255 596 2259
rect 590 2254 596 2255
rect 710 2259 716 2260
rect 710 2255 711 2259
rect 715 2255 716 2259
rect 710 2254 716 2255
rect 822 2259 828 2260
rect 822 2255 823 2259
rect 827 2255 828 2259
rect 822 2254 828 2255
rect 934 2259 940 2260
rect 934 2255 935 2259
rect 939 2255 940 2259
rect 934 2254 940 2255
rect 1054 2259 1060 2260
rect 1054 2255 1055 2259
rect 1059 2255 1060 2259
rect 1054 2254 1060 2255
rect 1174 2259 1180 2260
rect 1174 2255 1175 2259
rect 1179 2255 1180 2259
rect 1174 2254 1180 2255
rect 1824 2250 1826 2265
rect 1864 2250 1866 2265
rect 2336 2260 2338 2265
rect 2448 2260 2450 2265
rect 2584 2260 2586 2265
rect 2736 2260 2738 2265
rect 2912 2260 2914 2265
rect 3104 2260 3106 2265
rect 3304 2260 3306 2265
rect 3480 2260 3482 2265
rect 2334 2259 2340 2260
rect 2334 2255 2335 2259
rect 2339 2255 2340 2259
rect 2334 2254 2340 2255
rect 2446 2259 2452 2260
rect 2446 2255 2447 2259
rect 2451 2255 2452 2259
rect 2446 2254 2452 2255
rect 2582 2259 2588 2260
rect 2582 2255 2583 2259
rect 2587 2255 2588 2259
rect 2582 2254 2588 2255
rect 2734 2259 2740 2260
rect 2734 2255 2735 2259
rect 2739 2255 2740 2259
rect 2734 2254 2740 2255
rect 2910 2259 2916 2260
rect 2910 2255 2911 2259
rect 2915 2255 2916 2259
rect 2910 2254 2916 2255
rect 3102 2259 3108 2260
rect 3102 2255 3103 2259
rect 3107 2255 3108 2259
rect 3102 2254 3108 2255
rect 3302 2259 3308 2260
rect 3302 2255 3303 2259
rect 3307 2255 3308 2259
rect 3302 2254 3308 2255
rect 3478 2259 3484 2260
rect 3478 2255 3479 2259
rect 3483 2255 3484 2259
rect 3478 2254 3484 2255
rect 3576 2250 3578 2265
rect 110 2249 116 2250
rect 110 2245 111 2249
rect 115 2245 116 2249
rect 110 2244 116 2245
rect 1822 2249 1828 2250
rect 1822 2245 1823 2249
rect 1827 2245 1828 2249
rect 1822 2244 1828 2245
rect 1862 2249 1868 2250
rect 1862 2245 1863 2249
rect 1867 2245 1868 2249
rect 1862 2244 1868 2245
rect 3574 2249 3580 2250
rect 3574 2245 3575 2249
rect 3579 2245 3580 2249
rect 3574 2244 3580 2245
rect 110 2232 116 2233
rect 110 2228 111 2232
rect 115 2228 116 2232
rect 110 2227 116 2228
rect 1822 2232 1828 2233
rect 1822 2228 1823 2232
rect 1827 2228 1828 2232
rect 1822 2227 1828 2228
rect 1862 2232 1868 2233
rect 1862 2228 1863 2232
rect 1867 2228 1868 2232
rect 1862 2227 1868 2228
rect 3574 2232 3580 2233
rect 3574 2228 3575 2232
rect 3579 2228 3580 2232
rect 3574 2227 3580 2228
rect 112 2199 114 2227
rect 142 2219 148 2220
rect 142 2215 143 2219
rect 147 2215 148 2219
rect 142 2214 148 2215
rect 238 2219 244 2220
rect 238 2215 239 2219
rect 243 2215 244 2219
rect 238 2214 244 2215
rect 358 2219 364 2220
rect 358 2215 359 2219
rect 363 2215 364 2219
rect 358 2214 364 2215
rect 478 2219 484 2220
rect 478 2215 479 2219
rect 483 2215 484 2219
rect 478 2214 484 2215
rect 598 2219 604 2220
rect 598 2215 599 2219
rect 603 2215 604 2219
rect 598 2214 604 2215
rect 718 2219 724 2220
rect 718 2215 719 2219
rect 723 2215 724 2219
rect 718 2214 724 2215
rect 830 2219 836 2220
rect 830 2215 831 2219
rect 835 2215 836 2219
rect 830 2214 836 2215
rect 942 2219 948 2220
rect 942 2215 943 2219
rect 947 2215 948 2219
rect 942 2214 948 2215
rect 1062 2219 1068 2220
rect 1062 2215 1063 2219
rect 1067 2215 1068 2219
rect 1062 2214 1068 2215
rect 1182 2219 1188 2220
rect 1182 2215 1183 2219
rect 1187 2215 1188 2219
rect 1182 2214 1188 2215
rect 144 2199 146 2214
rect 240 2199 242 2214
rect 360 2199 362 2214
rect 480 2199 482 2214
rect 600 2199 602 2214
rect 720 2199 722 2214
rect 832 2199 834 2214
rect 944 2199 946 2214
rect 1064 2199 1066 2214
rect 1184 2199 1186 2214
rect 1824 2199 1826 2227
rect 1864 2203 1866 2227
rect 2342 2219 2348 2220
rect 2342 2215 2343 2219
rect 2347 2215 2348 2219
rect 2342 2214 2348 2215
rect 2454 2219 2460 2220
rect 2454 2215 2455 2219
rect 2459 2215 2460 2219
rect 2454 2214 2460 2215
rect 2590 2219 2596 2220
rect 2590 2215 2591 2219
rect 2595 2215 2596 2219
rect 2590 2214 2596 2215
rect 2742 2219 2748 2220
rect 2742 2215 2743 2219
rect 2747 2215 2748 2219
rect 2742 2214 2748 2215
rect 2918 2219 2924 2220
rect 2918 2215 2919 2219
rect 2923 2215 2924 2219
rect 2918 2214 2924 2215
rect 3110 2219 3116 2220
rect 3110 2215 3111 2219
rect 3115 2215 3116 2219
rect 3110 2214 3116 2215
rect 3310 2219 3316 2220
rect 3310 2215 3311 2219
rect 3315 2215 3316 2219
rect 3310 2214 3316 2215
rect 3486 2219 3492 2220
rect 3486 2215 3487 2219
rect 3491 2215 3492 2219
rect 3486 2214 3492 2215
rect 2344 2203 2346 2214
rect 2456 2203 2458 2214
rect 2592 2203 2594 2214
rect 2744 2203 2746 2214
rect 2920 2203 2922 2214
rect 3112 2203 3114 2214
rect 3312 2203 3314 2214
rect 3488 2203 3490 2214
rect 3576 2203 3578 2227
rect 1863 2202 1867 2203
rect 111 2198 115 2199
rect 111 2193 115 2194
rect 143 2198 147 2199
rect 143 2193 147 2194
rect 239 2198 243 2199
rect 239 2193 243 2194
rect 247 2198 251 2199
rect 247 2193 251 2194
rect 359 2198 363 2199
rect 359 2193 363 2194
rect 383 2198 387 2199
rect 383 2193 387 2194
rect 479 2198 483 2199
rect 479 2193 483 2194
rect 519 2198 523 2199
rect 519 2193 523 2194
rect 599 2198 603 2199
rect 599 2193 603 2194
rect 655 2198 659 2199
rect 655 2193 659 2194
rect 719 2198 723 2199
rect 719 2193 723 2194
rect 783 2198 787 2199
rect 783 2193 787 2194
rect 831 2198 835 2199
rect 831 2193 835 2194
rect 911 2198 915 2199
rect 911 2193 915 2194
rect 943 2198 947 2199
rect 943 2193 947 2194
rect 1031 2198 1035 2199
rect 1031 2193 1035 2194
rect 1063 2198 1067 2199
rect 1063 2193 1067 2194
rect 1159 2198 1163 2199
rect 1159 2193 1163 2194
rect 1183 2198 1187 2199
rect 1183 2193 1187 2194
rect 1287 2198 1291 2199
rect 1287 2193 1291 2194
rect 1823 2198 1827 2199
rect 1863 2197 1867 2198
rect 2255 2202 2259 2203
rect 2255 2197 2259 2198
rect 2343 2202 2347 2203
rect 2343 2197 2347 2198
rect 2439 2202 2443 2203
rect 2439 2197 2443 2198
rect 2455 2202 2459 2203
rect 2455 2197 2459 2198
rect 2551 2202 2555 2203
rect 2551 2197 2555 2198
rect 2591 2202 2595 2203
rect 2591 2197 2595 2198
rect 2695 2202 2699 2203
rect 2695 2197 2699 2198
rect 2743 2202 2747 2203
rect 2743 2197 2747 2198
rect 2871 2202 2875 2203
rect 2871 2197 2875 2198
rect 2919 2202 2923 2203
rect 2919 2197 2923 2198
rect 3071 2202 3075 2203
rect 3071 2197 3075 2198
rect 3111 2202 3115 2203
rect 3111 2197 3115 2198
rect 3287 2202 3291 2203
rect 3287 2197 3291 2198
rect 3311 2202 3315 2203
rect 3311 2197 3315 2198
rect 3487 2202 3491 2203
rect 3487 2197 3491 2198
rect 3575 2202 3579 2203
rect 3575 2197 3579 2198
rect 1823 2193 1827 2194
rect 112 2169 114 2193
rect 144 2182 146 2193
rect 248 2182 250 2193
rect 384 2182 386 2193
rect 520 2182 522 2193
rect 656 2182 658 2193
rect 784 2182 786 2193
rect 912 2182 914 2193
rect 1032 2182 1034 2193
rect 1160 2182 1162 2193
rect 1288 2182 1290 2193
rect 142 2181 148 2182
rect 142 2177 143 2181
rect 147 2177 148 2181
rect 142 2176 148 2177
rect 246 2181 252 2182
rect 246 2177 247 2181
rect 251 2177 252 2181
rect 246 2176 252 2177
rect 382 2181 388 2182
rect 382 2177 383 2181
rect 387 2177 388 2181
rect 382 2176 388 2177
rect 518 2181 524 2182
rect 518 2177 519 2181
rect 523 2177 524 2181
rect 518 2176 524 2177
rect 654 2181 660 2182
rect 654 2177 655 2181
rect 659 2177 660 2181
rect 654 2176 660 2177
rect 782 2181 788 2182
rect 782 2177 783 2181
rect 787 2177 788 2181
rect 782 2176 788 2177
rect 910 2181 916 2182
rect 910 2177 911 2181
rect 915 2177 916 2181
rect 910 2176 916 2177
rect 1030 2181 1036 2182
rect 1030 2177 1031 2181
rect 1035 2177 1036 2181
rect 1030 2176 1036 2177
rect 1158 2181 1164 2182
rect 1158 2177 1159 2181
rect 1163 2177 1164 2181
rect 1158 2176 1164 2177
rect 1286 2181 1292 2182
rect 1286 2177 1287 2181
rect 1291 2177 1292 2181
rect 1286 2176 1292 2177
rect 1824 2169 1826 2193
rect 1864 2173 1866 2197
rect 2256 2186 2258 2197
rect 2344 2186 2346 2197
rect 2440 2186 2442 2197
rect 2552 2186 2554 2197
rect 2696 2186 2698 2197
rect 2872 2186 2874 2197
rect 3072 2186 3074 2197
rect 3288 2186 3290 2197
rect 3488 2186 3490 2197
rect 2254 2185 2260 2186
rect 2254 2181 2255 2185
rect 2259 2181 2260 2185
rect 2254 2180 2260 2181
rect 2342 2185 2348 2186
rect 2342 2181 2343 2185
rect 2347 2181 2348 2185
rect 2342 2180 2348 2181
rect 2438 2185 2444 2186
rect 2438 2181 2439 2185
rect 2443 2181 2444 2185
rect 2438 2180 2444 2181
rect 2550 2185 2556 2186
rect 2550 2181 2551 2185
rect 2555 2181 2556 2185
rect 2550 2180 2556 2181
rect 2694 2185 2700 2186
rect 2694 2181 2695 2185
rect 2699 2181 2700 2185
rect 2694 2180 2700 2181
rect 2870 2185 2876 2186
rect 2870 2181 2871 2185
rect 2875 2181 2876 2185
rect 2870 2180 2876 2181
rect 3070 2185 3076 2186
rect 3070 2181 3071 2185
rect 3075 2181 3076 2185
rect 3070 2180 3076 2181
rect 3286 2185 3292 2186
rect 3286 2181 3287 2185
rect 3291 2181 3292 2185
rect 3286 2180 3292 2181
rect 3486 2185 3492 2186
rect 3486 2181 3487 2185
rect 3491 2181 3492 2185
rect 3486 2180 3492 2181
rect 3576 2173 3578 2197
rect 1862 2172 1868 2173
rect 110 2168 116 2169
rect 110 2164 111 2168
rect 115 2164 116 2168
rect 110 2163 116 2164
rect 1822 2168 1828 2169
rect 1822 2164 1823 2168
rect 1827 2164 1828 2168
rect 1862 2168 1863 2172
rect 1867 2168 1868 2172
rect 1862 2167 1868 2168
rect 3574 2172 3580 2173
rect 3574 2168 3575 2172
rect 3579 2168 3580 2172
rect 3574 2167 3580 2168
rect 1822 2163 1828 2164
rect 1862 2155 1868 2156
rect 110 2151 116 2152
rect 110 2147 111 2151
rect 115 2147 116 2151
rect 110 2146 116 2147
rect 1822 2151 1828 2152
rect 1822 2147 1823 2151
rect 1827 2147 1828 2151
rect 1862 2151 1863 2155
rect 1867 2151 1868 2155
rect 1862 2150 1868 2151
rect 3574 2155 3580 2156
rect 3574 2151 3575 2155
rect 3579 2151 3580 2155
rect 3574 2150 3580 2151
rect 1822 2146 1828 2147
rect 112 2123 114 2146
rect 134 2141 140 2142
rect 134 2137 135 2141
rect 139 2137 140 2141
rect 134 2136 140 2137
rect 238 2141 244 2142
rect 238 2137 239 2141
rect 243 2137 244 2141
rect 238 2136 244 2137
rect 374 2141 380 2142
rect 374 2137 375 2141
rect 379 2137 380 2141
rect 374 2136 380 2137
rect 510 2141 516 2142
rect 510 2137 511 2141
rect 515 2137 516 2141
rect 510 2136 516 2137
rect 646 2141 652 2142
rect 646 2137 647 2141
rect 651 2137 652 2141
rect 646 2136 652 2137
rect 774 2141 780 2142
rect 774 2137 775 2141
rect 779 2137 780 2141
rect 774 2136 780 2137
rect 902 2141 908 2142
rect 902 2137 903 2141
rect 907 2137 908 2141
rect 902 2136 908 2137
rect 1022 2141 1028 2142
rect 1022 2137 1023 2141
rect 1027 2137 1028 2141
rect 1022 2136 1028 2137
rect 1150 2141 1156 2142
rect 1150 2137 1151 2141
rect 1155 2137 1156 2141
rect 1150 2136 1156 2137
rect 1278 2141 1284 2142
rect 1278 2137 1279 2141
rect 1283 2137 1284 2141
rect 1278 2136 1284 2137
rect 136 2123 138 2136
rect 240 2123 242 2136
rect 376 2123 378 2136
rect 512 2123 514 2136
rect 648 2123 650 2136
rect 776 2123 778 2136
rect 904 2123 906 2136
rect 1024 2123 1026 2136
rect 1152 2123 1154 2136
rect 1280 2123 1282 2136
rect 1824 2123 1826 2146
rect 1864 2127 1866 2150
rect 2246 2145 2252 2146
rect 2246 2141 2247 2145
rect 2251 2141 2252 2145
rect 2246 2140 2252 2141
rect 2334 2145 2340 2146
rect 2334 2141 2335 2145
rect 2339 2141 2340 2145
rect 2334 2140 2340 2141
rect 2430 2145 2436 2146
rect 2430 2141 2431 2145
rect 2435 2141 2436 2145
rect 2430 2140 2436 2141
rect 2542 2145 2548 2146
rect 2542 2141 2543 2145
rect 2547 2141 2548 2145
rect 2542 2140 2548 2141
rect 2686 2145 2692 2146
rect 2686 2141 2687 2145
rect 2691 2141 2692 2145
rect 2686 2140 2692 2141
rect 2862 2145 2868 2146
rect 2862 2141 2863 2145
rect 2867 2141 2868 2145
rect 2862 2140 2868 2141
rect 3062 2145 3068 2146
rect 3062 2141 3063 2145
rect 3067 2141 3068 2145
rect 3062 2140 3068 2141
rect 3278 2145 3284 2146
rect 3278 2141 3279 2145
rect 3283 2141 3284 2145
rect 3278 2140 3284 2141
rect 3478 2145 3484 2146
rect 3478 2141 3479 2145
rect 3483 2141 3484 2145
rect 3478 2140 3484 2141
rect 2248 2127 2250 2140
rect 2336 2127 2338 2140
rect 2432 2127 2434 2140
rect 2544 2127 2546 2140
rect 2688 2127 2690 2140
rect 2864 2127 2866 2140
rect 3064 2127 3066 2140
rect 3280 2127 3282 2140
rect 3480 2127 3482 2140
rect 3576 2127 3578 2150
rect 1863 2126 1867 2127
rect 111 2122 115 2123
rect 111 2117 115 2118
rect 135 2122 139 2123
rect 135 2117 139 2118
rect 231 2122 235 2123
rect 231 2117 235 2118
rect 239 2122 243 2123
rect 239 2117 243 2118
rect 359 2122 363 2123
rect 359 2117 363 2118
rect 375 2122 379 2123
rect 375 2117 379 2118
rect 479 2122 483 2123
rect 479 2117 483 2118
rect 511 2122 515 2123
rect 511 2117 515 2118
rect 599 2122 603 2123
rect 599 2117 603 2118
rect 647 2122 651 2123
rect 647 2117 651 2118
rect 719 2122 723 2123
rect 719 2117 723 2118
rect 775 2122 779 2123
rect 775 2117 779 2118
rect 831 2122 835 2123
rect 831 2117 835 2118
rect 903 2122 907 2123
rect 903 2117 907 2118
rect 943 2122 947 2123
rect 943 2117 947 2118
rect 1023 2122 1027 2123
rect 1023 2117 1027 2118
rect 1055 2122 1059 2123
rect 1055 2117 1059 2118
rect 1151 2122 1155 2123
rect 1151 2117 1155 2118
rect 1175 2122 1179 2123
rect 1175 2117 1179 2118
rect 1279 2122 1283 2123
rect 1279 2117 1283 2118
rect 1823 2122 1827 2123
rect 1863 2121 1867 2122
rect 2151 2126 2155 2127
rect 2151 2121 2155 2122
rect 2239 2126 2243 2127
rect 2239 2121 2243 2122
rect 2247 2126 2251 2127
rect 2247 2121 2251 2122
rect 2327 2126 2331 2127
rect 2327 2121 2331 2122
rect 2335 2126 2339 2127
rect 2335 2121 2339 2122
rect 2415 2126 2419 2127
rect 2415 2121 2419 2122
rect 2431 2126 2435 2127
rect 2431 2121 2435 2122
rect 2503 2126 2507 2127
rect 2503 2121 2507 2122
rect 2543 2126 2547 2127
rect 2543 2121 2547 2122
rect 2615 2126 2619 2127
rect 2615 2121 2619 2122
rect 2687 2126 2691 2127
rect 2687 2121 2691 2122
rect 2751 2126 2755 2127
rect 2751 2121 2755 2122
rect 2863 2126 2867 2127
rect 2863 2121 2867 2122
rect 2919 2126 2923 2127
rect 2919 2121 2923 2122
rect 3063 2126 3067 2127
rect 3063 2121 3067 2122
rect 3103 2126 3107 2127
rect 3103 2121 3107 2122
rect 3279 2126 3283 2127
rect 3279 2121 3283 2122
rect 3303 2126 3307 2127
rect 3303 2121 3307 2122
rect 3479 2126 3483 2127
rect 3479 2121 3483 2122
rect 3575 2126 3579 2127
rect 3575 2121 3579 2122
rect 1823 2117 1827 2118
rect 112 2102 114 2117
rect 136 2112 138 2117
rect 232 2112 234 2117
rect 360 2112 362 2117
rect 480 2112 482 2117
rect 600 2112 602 2117
rect 720 2112 722 2117
rect 832 2112 834 2117
rect 944 2112 946 2117
rect 1056 2112 1058 2117
rect 1176 2112 1178 2117
rect 134 2111 140 2112
rect 134 2107 135 2111
rect 139 2107 140 2111
rect 134 2106 140 2107
rect 230 2111 236 2112
rect 230 2107 231 2111
rect 235 2107 236 2111
rect 230 2106 236 2107
rect 358 2111 364 2112
rect 358 2107 359 2111
rect 363 2107 364 2111
rect 358 2106 364 2107
rect 478 2111 484 2112
rect 478 2107 479 2111
rect 483 2107 484 2111
rect 478 2106 484 2107
rect 598 2111 604 2112
rect 598 2107 599 2111
rect 603 2107 604 2111
rect 598 2106 604 2107
rect 718 2111 724 2112
rect 718 2107 719 2111
rect 723 2107 724 2111
rect 718 2106 724 2107
rect 830 2111 836 2112
rect 830 2107 831 2111
rect 835 2107 836 2111
rect 830 2106 836 2107
rect 942 2111 948 2112
rect 942 2107 943 2111
rect 947 2107 948 2111
rect 942 2106 948 2107
rect 1054 2111 1060 2112
rect 1054 2107 1055 2111
rect 1059 2107 1060 2111
rect 1054 2106 1060 2107
rect 1174 2111 1180 2112
rect 1174 2107 1175 2111
rect 1179 2107 1180 2111
rect 1174 2106 1180 2107
rect 1824 2102 1826 2117
rect 1864 2106 1866 2121
rect 2152 2116 2154 2121
rect 2240 2116 2242 2121
rect 2328 2116 2330 2121
rect 2416 2116 2418 2121
rect 2504 2116 2506 2121
rect 2616 2116 2618 2121
rect 2752 2116 2754 2121
rect 2920 2116 2922 2121
rect 3104 2116 3106 2121
rect 3304 2116 3306 2121
rect 3480 2116 3482 2121
rect 2150 2115 2156 2116
rect 2150 2111 2151 2115
rect 2155 2111 2156 2115
rect 2150 2110 2156 2111
rect 2238 2115 2244 2116
rect 2238 2111 2239 2115
rect 2243 2111 2244 2115
rect 2238 2110 2244 2111
rect 2326 2115 2332 2116
rect 2326 2111 2327 2115
rect 2331 2111 2332 2115
rect 2326 2110 2332 2111
rect 2414 2115 2420 2116
rect 2414 2111 2415 2115
rect 2419 2111 2420 2115
rect 2414 2110 2420 2111
rect 2502 2115 2508 2116
rect 2502 2111 2503 2115
rect 2507 2111 2508 2115
rect 2502 2110 2508 2111
rect 2614 2115 2620 2116
rect 2614 2111 2615 2115
rect 2619 2111 2620 2115
rect 2614 2110 2620 2111
rect 2750 2115 2756 2116
rect 2750 2111 2751 2115
rect 2755 2111 2756 2115
rect 2750 2110 2756 2111
rect 2918 2115 2924 2116
rect 2918 2111 2919 2115
rect 2923 2111 2924 2115
rect 2918 2110 2924 2111
rect 3102 2115 3108 2116
rect 3102 2111 3103 2115
rect 3107 2111 3108 2115
rect 3102 2110 3108 2111
rect 3302 2115 3308 2116
rect 3302 2111 3303 2115
rect 3307 2111 3308 2115
rect 3302 2110 3308 2111
rect 3478 2115 3484 2116
rect 3478 2111 3479 2115
rect 3483 2111 3484 2115
rect 3478 2110 3484 2111
rect 3576 2106 3578 2121
rect 1862 2105 1868 2106
rect 110 2101 116 2102
rect 110 2097 111 2101
rect 115 2097 116 2101
rect 110 2096 116 2097
rect 1822 2101 1828 2102
rect 1822 2097 1823 2101
rect 1827 2097 1828 2101
rect 1862 2101 1863 2105
rect 1867 2101 1868 2105
rect 1862 2100 1868 2101
rect 3574 2105 3580 2106
rect 3574 2101 3575 2105
rect 3579 2101 3580 2105
rect 3574 2100 3580 2101
rect 1822 2096 1828 2097
rect 1862 2088 1868 2089
rect 110 2084 116 2085
rect 110 2080 111 2084
rect 115 2080 116 2084
rect 110 2079 116 2080
rect 1822 2084 1828 2085
rect 1822 2080 1823 2084
rect 1827 2080 1828 2084
rect 1862 2084 1863 2088
rect 1867 2084 1868 2088
rect 1862 2083 1868 2084
rect 3574 2088 3580 2089
rect 3574 2084 3575 2088
rect 3579 2084 3580 2088
rect 3574 2083 3580 2084
rect 1822 2079 1828 2080
rect 112 2043 114 2079
rect 142 2071 148 2072
rect 142 2067 143 2071
rect 147 2067 148 2071
rect 142 2066 148 2067
rect 238 2071 244 2072
rect 238 2067 239 2071
rect 243 2067 244 2071
rect 238 2066 244 2067
rect 366 2071 372 2072
rect 366 2067 367 2071
rect 371 2067 372 2071
rect 366 2066 372 2067
rect 486 2071 492 2072
rect 486 2067 487 2071
rect 491 2067 492 2071
rect 486 2066 492 2067
rect 606 2071 612 2072
rect 606 2067 607 2071
rect 611 2067 612 2071
rect 606 2066 612 2067
rect 726 2071 732 2072
rect 726 2067 727 2071
rect 731 2067 732 2071
rect 726 2066 732 2067
rect 838 2071 844 2072
rect 838 2067 839 2071
rect 843 2067 844 2071
rect 838 2066 844 2067
rect 950 2071 956 2072
rect 950 2067 951 2071
rect 955 2067 956 2071
rect 950 2066 956 2067
rect 1062 2071 1068 2072
rect 1062 2067 1063 2071
rect 1067 2067 1068 2071
rect 1062 2066 1068 2067
rect 1182 2071 1188 2072
rect 1182 2067 1183 2071
rect 1187 2067 1188 2071
rect 1182 2066 1188 2067
rect 144 2043 146 2066
rect 240 2043 242 2066
rect 368 2043 370 2066
rect 488 2043 490 2066
rect 608 2043 610 2066
rect 728 2043 730 2066
rect 840 2043 842 2066
rect 952 2043 954 2066
rect 1064 2043 1066 2066
rect 1184 2043 1186 2066
rect 1824 2043 1826 2079
rect 1864 2055 1866 2083
rect 2158 2075 2164 2076
rect 2158 2071 2159 2075
rect 2163 2071 2164 2075
rect 2158 2070 2164 2071
rect 2246 2075 2252 2076
rect 2246 2071 2247 2075
rect 2251 2071 2252 2075
rect 2246 2070 2252 2071
rect 2334 2075 2340 2076
rect 2334 2071 2335 2075
rect 2339 2071 2340 2075
rect 2334 2070 2340 2071
rect 2422 2075 2428 2076
rect 2422 2071 2423 2075
rect 2427 2071 2428 2075
rect 2422 2070 2428 2071
rect 2510 2075 2516 2076
rect 2510 2071 2511 2075
rect 2515 2071 2516 2075
rect 2510 2070 2516 2071
rect 2622 2075 2628 2076
rect 2622 2071 2623 2075
rect 2627 2071 2628 2075
rect 2622 2070 2628 2071
rect 2758 2075 2764 2076
rect 2758 2071 2759 2075
rect 2763 2071 2764 2075
rect 2758 2070 2764 2071
rect 2926 2075 2932 2076
rect 2926 2071 2927 2075
rect 2931 2071 2932 2075
rect 2926 2070 2932 2071
rect 3110 2075 3116 2076
rect 3110 2071 3111 2075
rect 3115 2071 3116 2075
rect 3110 2070 3116 2071
rect 3310 2075 3316 2076
rect 3310 2071 3311 2075
rect 3315 2071 3316 2075
rect 3310 2070 3316 2071
rect 3486 2075 3492 2076
rect 3486 2071 3487 2075
rect 3491 2071 3492 2075
rect 3486 2070 3492 2071
rect 2160 2055 2162 2070
rect 2248 2055 2250 2070
rect 2336 2055 2338 2070
rect 2424 2055 2426 2070
rect 2512 2055 2514 2070
rect 2624 2055 2626 2070
rect 2760 2055 2762 2070
rect 2928 2055 2930 2070
rect 3112 2055 3114 2070
rect 3312 2055 3314 2070
rect 3488 2055 3490 2070
rect 3576 2055 3578 2083
rect 1863 2054 1867 2055
rect 1863 2049 1867 2050
rect 1999 2054 2003 2055
rect 1999 2049 2003 2050
rect 2127 2054 2131 2055
rect 2127 2049 2131 2050
rect 2159 2054 2163 2055
rect 2159 2049 2163 2050
rect 2247 2054 2251 2055
rect 2247 2049 2251 2050
rect 2255 2054 2259 2055
rect 2255 2049 2259 2050
rect 2335 2054 2339 2055
rect 2335 2049 2339 2050
rect 2399 2054 2403 2055
rect 2399 2049 2403 2050
rect 2423 2054 2427 2055
rect 2423 2049 2427 2050
rect 2511 2054 2515 2055
rect 2511 2049 2515 2050
rect 2551 2054 2555 2055
rect 2551 2049 2555 2050
rect 2623 2054 2627 2055
rect 2623 2049 2627 2050
rect 2711 2054 2715 2055
rect 2711 2049 2715 2050
rect 2759 2054 2763 2055
rect 2759 2049 2763 2050
rect 2879 2054 2883 2055
rect 2879 2049 2883 2050
rect 2927 2054 2931 2055
rect 2927 2049 2931 2050
rect 3063 2054 3067 2055
rect 3063 2049 3067 2050
rect 3111 2054 3115 2055
rect 3111 2049 3115 2050
rect 3247 2054 3251 2055
rect 3247 2049 3251 2050
rect 3311 2054 3315 2055
rect 3311 2049 3315 2050
rect 3439 2054 3443 2055
rect 3439 2049 3443 2050
rect 3487 2054 3491 2055
rect 3487 2049 3491 2050
rect 3575 2054 3579 2055
rect 3575 2049 3579 2050
rect 111 2042 115 2043
rect 111 2037 115 2038
rect 143 2042 147 2043
rect 143 2037 147 2038
rect 167 2042 171 2043
rect 167 2037 171 2038
rect 239 2042 243 2043
rect 239 2037 243 2038
rect 311 2042 315 2043
rect 311 2037 315 2038
rect 367 2042 371 2043
rect 367 2037 371 2038
rect 447 2042 451 2043
rect 447 2037 451 2038
rect 487 2042 491 2043
rect 487 2037 491 2038
rect 575 2042 579 2043
rect 575 2037 579 2038
rect 607 2042 611 2043
rect 607 2037 611 2038
rect 695 2042 699 2043
rect 695 2037 699 2038
rect 727 2042 731 2043
rect 727 2037 731 2038
rect 807 2042 811 2043
rect 807 2037 811 2038
rect 839 2042 843 2043
rect 839 2037 843 2038
rect 911 2042 915 2043
rect 911 2037 915 2038
rect 951 2042 955 2043
rect 951 2037 955 2038
rect 1015 2042 1019 2043
rect 1015 2037 1019 2038
rect 1063 2042 1067 2043
rect 1063 2037 1067 2038
rect 1119 2042 1123 2043
rect 1119 2037 1123 2038
rect 1183 2042 1187 2043
rect 1183 2037 1187 2038
rect 1223 2042 1227 2043
rect 1223 2037 1227 2038
rect 1327 2042 1331 2043
rect 1327 2037 1331 2038
rect 1823 2042 1827 2043
rect 1823 2037 1827 2038
rect 112 2013 114 2037
rect 168 2026 170 2037
rect 312 2026 314 2037
rect 448 2026 450 2037
rect 576 2026 578 2037
rect 696 2026 698 2037
rect 808 2026 810 2037
rect 912 2026 914 2037
rect 1016 2026 1018 2037
rect 1120 2026 1122 2037
rect 1224 2026 1226 2037
rect 1328 2026 1330 2037
rect 166 2025 172 2026
rect 166 2021 167 2025
rect 171 2021 172 2025
rect 166 2020 172 2021
rect 310 2025 316 2026
rect 310 2021 311 2025
rect 315 2021 316 2025
rect 310 2020 316 2021
rect 446 2025 452 2026
rect 446 2021 447 2025
rect 451 2021 452 2025
rect 446 2020 452 2021
rect 574 2025 580 2026
rect 574 2021 575 2025
rect 579 2021 580 2025
rect 574 2020 580 2021
rect 694 2025 700 2026
rect 694 2021 695 2025
rect 699 2021 700 2025
rect 694 2020 700 2021
rect 806 2025 812 2026
rect 806 2021 807 2025
rect 811 2021 812 2025
rect 806 2020 812 2021
rect 910 2025 916 2026
rect 910 2021 911 2025
rect 915 2021 916 2025
rect 910 2020 916 2021
rect 1014 2025 1020 2026
rect 1014 2021 1015 2025
rect 1019 2021 1020 2025
rect 1014 2020 1020 2021
rect 1118 2025 1124 2026
rect 1118 2021 1119 2025
rect 1123 2021 1124 2025
rect 1118 2020 1124 2021
rect 1222 2025 1228 2026
rect 1222 2021 1223 2025
rect 1227 2021 1228 2025
rect 1222 2020 1228 2021
rect 1326 2025 1332 2026
rect 1326 2021 1327 2025
rect 1331 2021 1332 2025
rect 1326 2020 1332 2021
rect 1824 2013 1826 2037
rect 1864 2025 1866 2049
rect 2000 2038 2002 2049
rect 2128 2038 2130 2049
rect 2256 2038 2258 2049
rect 2400 2038 2402 2049
rect 2552 2038 2554 2049
rect 2712 2038 2714 2049
rect 2880 2038 2882 2049
rect 3064 2038 3066 2049
rect 3248 2038 3250 2049
rect 3440 2038 3442 2049
rect 1998 2037 2004 2038
rect 1998 2033 1999 2037
rect 2003 2033 2004 2037
rect 1998 2032 2004 2033
rect 2126 2037 2132 2038
rect 2126 2033 2127 2037
rect 2131 2033 2132 2037
rect 2126 2032 2132 2033
rect 2254 2037 2260 2038
rect 2254 2033 2255 2037
rect 2259 2033 2260 2037
rect 2254 2032 2260 2033
rect 2398 2037 2404 2038
rect 2398 2033 2399 2037
rect 2403 2033 2404 2037
rect 2398 2032 2404 2033
rect 2550 2037 2556 2038
rect 2550 2033 2551 2037
rect 2555 2033 2556 2037
rect 2550 2032 2556 2033
rect 2710 2037 2716 2038
rect 2710 2033 2711 2037
rect 2715 2033 2716 2037
rect 2710 2032 2716 2033
rect 2878 2037 2884 2038
rect 2878 2033 2879 2037
rect 2883 2033 2884 2037
rect 2878 2032 2884 2033
rect 3062 2037 3068 2038
rect 3062 2033 3063 2037
rect 3067 2033 3068 2037
rect 3062 2032 3068 2033
rect 3246 2037 3252 2038
rect 3246 2033 3247 2037
rect 3251 2033 3252 2037
rect 3246 2032 3252 2033
rect 3438 2037 3444 2038
rect 3438 2033 3439 2037
rect 3443 2033 3444 2037
rect 3438 2032 3444 2033
rect 3576 2025 3578 2049
rect 1862 2024 1868 2025
rect 1862 2020 1863 2024
rect 1867 2020 1868 2024
rect 1862 2019 1868 2020
rect 3574 2024 3580 2025
rect 3574 2020 3575 2024
rect 3579 2020 3580 2024
rect 3574 2019 3580 2020
rect 110 2012 116 2013
rect 110 2008 111 2012
rect 115 2008 116 2012
rect 110 2007 116 2008
rect 1822 2012 1828 2013
rect 1822 2008 1823 2012
rect 1827 2008 1828 2012
rect 1822 2007 1828 2008
rect 1862 2007 1868 2008
rect 1862 2003 1863 2007
rect 1867 2003 1868 2007
rect 1862 2002 1868 2003
rect 3574 2007 3580 2008
rect 3574 2003 3575 2007
rect 3579 2003 3580 2007
rect 3574 2002 3580 2003
rect 110 1995 116 1996
rect 110 1991 111 1995
rect 115 1991 116 1995
rect 110 1990 116 1991
rect 1822 1995 1828 1996
rect 1822 1991 1823 1995
rect 1827 1991 1828 1995
rect 1822 1990 1828 1991
rect 112 1975 114 1990
rect 158 1985 164 1986
rect 158 1981 159 1985
rect 163 1981 164 1985
rect 158 1980 164 1981
rect 302 1985 308 1986
rect 302 1981 303 1985
rect 307 1981 308 1985
rect 302 1980 308 1981
rect 438 1985 444 1986
rect 438 1981 439 1985
rect 443 1981 444 1985
rect 438 1980 444 1981
rect 566 1985 572 1986
rect 566 1981 567 1985
rect 571 1981 572 1985
rect 566 1980 572 1981
rect 686 1985 692 1986
rect 686 1981 687 1985
rect 691 1981 692 1985
rect 686 1980 692 1981
rect 798 1985 804 1986
rect 798 1981 799 1985
rect 803 1981 804 1985
rect 798 1980 804 1981
rect 902 1985 908 1986
rect 902 1981 903 1985
rect 907 1981 908 1985
rect 902 1980 908 1981
rect 1006 1985 1012 1986
rect 1006 1981 1007 1985
rect 1011 1981 1012 1985
rect 1006 1980 1012 1981
rect 1110 1985 1116 1986
rect 1110 1981 1111 1985
rect 1115 1981 1116 1985
rect 1110 1980 1116 1981
rect 1214 1985 1220 1986
rect 1214 1981 1215 1985
rect 1219 1981 1220 1985
rect 1214 1980 1220 1981
rect 1318 1985 1324 1986
rect 1318 1981 1319 1985
rect 1323 1981 1324 1985
rect 1318 1980 1324 1981
rect 160 1975 162 1980
rect 304 1975 306 1980
rect 440 1975 442 1980
rect 568 1975 570 1980
rect 688 1975 690 1980
rect 800 1975 802 1980
rect 904 1975 906 1980
rect 1008 1975 1010 1980
rect 1112 1975 1114 1980
rect 1216 1975 1218 1980
rect 1320 1975 1322 1980
rect 1824 1975 1826 1990
rect 1864 1979 1866 2002
rect 1990 1997 1996 1998
rect 1990 1993 1991 1997
rect 1995 1993 1996 1997
rect 1990 1992 1996 1993
rect 2118 1997 2124 1998
rect 2118 1993 2119 1997
rect 2123 1993 2124 1997
rect 2118 1992 2124 1993
rect 2246 1997 2252 1998
rect 2246 1993 2247 1997
rect 2251 1993 2252 1997
rect 2246 1992 2252 1993
rect 2390 1997 2396 1998
rect 2390 1993 2391 1997
rect 2395 1993 2396 1997
rect 2390 1992 2396 1993
rect 2542 1997 2548 1998
rect 2542 1993 2543 1997
rect 2547 1993 2548 1997
rect 2542 1992 2548 1993
rect 2702 1997 2708 1998
rect 2702 1993 2703 1997
rect 2707 1993 2708 1997
rect 2702 1992 2708 1993
rect 2870 1997 2876 1998
rect 2870 1993 2871 1997
rect 2875 1993 2876 1997
rect 2870 1992 2876 1993
rect 3054 1997 3060 1998
rect 3054 1993 3055 1997
rect 3059 1993 3060 1997
rect 3054 1992 3060 1993
rect 3238 1997 3244 1998
rect 3238 1993 3239 1997
rect 3243 1993 3244 1997
rect 3238 1992 3244 1993
rect 3430 1997 3436 1998
rect 3430 1993 3431 1997
rect 3435 1993 3436 1997
rect 3430 1992 3436 1993
rect 1992 1979 1994 1992
rect 2120 1979 2122 1992
rect 2248 1979 2250 1992
rect 2392 1979 2394 1992
rect 2544 1979 2546 1992
rect 2704 1979 2706 1992
rect 2872 1979 2874 1992
rect 3056 1979 3058 1992
rect 3240 1979 3242 1992
rect 3432 1979 3434 1992
rect 3576 1979 3578 2002
rect 1863 1978 1867 1979
rect 111 1974 115 1975
rect 111 1969 115 1970
rect 159 1974 163 1975
rect 159 1969 163 1970
rect 295 1974 299 1975
rect 295 1969 299 1970
rect 303 1974 307 1975
rect 303 1969 307 1970
rect 439 1974 443 1975
rect 439 1969 443 1970
rect 567 1974 571 1975
rect 567 1969 571 1970
rect 583 1974 587 1975
rect 583 1969 587 1970
rect 687 1974 691 1975
rect 687 1969 691 1970
rect 719 1974 723 1975
rect 719 1969 723 1970
rect 799 1974 803 1975
rect 799 1969 803 1970
rect 855 1974 859 1975
rect 855 1969 859 1970
rect 903 1974 907 1975
rect 903 1969 907 1970
rect 991 1974 995 1975
rect 991 1969 995 1970
rect 1007 1974 1011 1975
rect 1007 1969 1011 1970
rect 1111 1974 1115 1975
rect 1111 1969 1115 1970
rect 1119 1974 1123 1975
rect 1119 1969 1123 1970
rect 1215 1974 1219 1975
rect 1215 1969 1219 1970
rect 1239 1974 1243 1975
rect 1239 1969 1243 1970
rect 1319 1974 1323 1975
rect 1319 1969 1323 1970
rect 1359 1974 1363 1975
rect 1359 1969 1363 1970
rect 1479 1974 1483 1975
rect 1479 1969 1483 1970
rect 1599 1974 1603 1975
rect 1599 1969 1603 1970
rect 1823 1974 1827 1975
rect 1863 1973 1867 1974
rect 1903 1978 1907 1979
rect 1903 1973 1907 1974
rect 1991 1978 1995 1979
rect 1991 1973 1995 1974
rect 2119 1978 2123 1979
rect 2119 1973 2123 1974
rect 2159 1978 2163 1979
rect 2159 1973 2163 1974
rect 2247 1978 2251 1979
rect 2247 1973 2251 1974
rect 2391 1978 2395 1979
rect 2391 1973 2395 1974
rect 2399 1978 2403 1979
rect 2399 1973 2403 1974
rect 2543 1978 2547 1979
rect 2543 1973 2547 1974
rect 2615 1978 2619 1979
rect 2615 1973 2619 1974
rect 2703 1978 2707 1979
rect 2703 1973 2707 1974
rect 2815 1978 2819 1979
rect 2815 1973 2819 1974
rect 2871 1978 2875 1979
rect 2871 1973 2875 1974
rect 2999 1978 3003 1979
rect 2999 1973 3003 1974
rect 3055 1978 3059 1979
rect 3055 1973 3059 1974
rect 3167 1978 3171 1979
rect 3167 1973 3171 1974
rect 3239 1978 3243 1979
rect 3239 1973 3243 1974
rect 3335 1978 3339 1979
rect 3335 1973 3339 1974
rect 3431 1978 3435 1979
rect 3431 1973 3435 1974
rect 3479 1978 3483 1979
rect 3479 1973 3483 1974
rect 3575 1978 3579 1979
rect 3575 1973 3579 1974
rect 1823 1969 1827 1970
rect 112 1954 114 1969
rect 160 1964 162 1969
rect 296 1964 298 1969
rect 440 1964 442 1969
rect 584 1964 586 1969
rect 720 1964 722 1969
rect 856 1964 858 1969
rect 992 1964 994 1969
rect 1120 1964 1122 1969
rect 1240 1964 1242 1969
rect 1360 1964 1362 1969
rect 1480 1964 1482 1969
rect 1600 1964 1602 1969
rect 158 1963 164 1964
rect 158 1959 159 1963
rect 163 1959 164 1963
rect 158 1958 164 1959
rect 294 1963 300 1964
rect 294 1959 295 1963
rect 299 1959 300 1963
rect 294 1958 300 1959
rect 438 1963 444 1964
rect 438 1959 439 1963
rect 443 1959 444 1963
rect 438 1958 444 1959
rect 582 1963 588 1964
rect 582 1959 583 1963
rect 587 1959 588 1963
rect 582 1958 588 1959
rect 718 1963 724 1964
rect 718 1959 719 1963
rect 723 1959 724 1963
rect 718 1958 724 1959
rect 854 1963 860 1964
rect 854 1959 855 1963
rect 859 1959 860 1963
rect 854 1958 860 1959
rect 990 1963 996 1964
rect 990 1959 991 1963
rect 995 1959 996 1963
rect 990 1958 996 1959
rect 1118 1963 1124 1964
rect 1118 1959 1119 1963
rect 1123 1959 1124 1963
rect 1118 1958 1124 1959
rect 1238 1963 1244 1964
rect 1238 1959 1239 1963
rect 1243 1959 1244 1963
rect 1238 1958 1244 1959
rect 1358 1963 1364 1964
rect 1358 1959 1359 1963
rect 1363 1959 1364 1963
rect 1358 1958 1364 1959
rect 1478 1963 1484 1964
rect 1478 1959 1479 1963
rect 1483 1959 1484 1963
rect 1478 1958 1484 1959
rect 1598 1963 1604 1964
rect 1598 1959 1599 1963
rect 1603 1959 1604 1963
rect 1598 1958 1604 1959
rect 1824 1954 1826 1969
rect 1864 1958 1866 1973
rect 1904 1968 1906 1973
rect 2160 1968 2162 1973
rect 2400 1968 2402 1973
rect 2616 1968 2618 1973
rect 2816 1968 2818 1973
rect 3000 1968 3002 1973
rect 3168 1968 3170 1973
rect 3336 1968 3338 1973
rect 3480 1968 3482 1973
rect 1902 1967 1908 1968
rect 1902 1963 1903 1967
rect 1907 1963 1908 1967
rect 1902 1962 1908 1963
rect 2158 1967 2164 1968
rect 2158 1963 2159 1967
rect 2163 1963 2164 1967
rect 2158 1962 2164 1963
rect 2398 1967 2404 1968
rect 2398 1963 2399 1967
rect 2403 1963 2404 1967
rect 2398 1962 2404 1963
rect 2614 1967 2620 1968
rect 2614 1963 2615 1967
rect 2619 1963 2620 1967
rect 2614 1962 2620 1963
rect 2814 1967 2820 1968
rect 2814 1963 2815 1967
rect 2819 1963 2820 1967
rect 2814 1962 2820 1963
rect 2998 1967 3004 1968
rect 2998 1963 2999 1967
rect 3003 1963 3004 1967
rect 2998 1962 3004 1963
rect 3166 1967 3172 1968
rect 3166 1963 3167 1967
rect 3171 1963 3172 1967
rect 3166 1962 3172 1963
rect 3334 1967 3340 1968
rect 3334 1963 3335 1967
rect 3339 1963 3340 1967
rect 3334 1962 3340 1963
rect 3478 1967 3484 1968
rect 3478 1963 3479 1967
rect 3483 1963 3484 1967
rect 3478 1962 3484 1963
rect 3576 1958 3578 1973
rect 1862 1957 1868 1958
rect 110 1953 116 1954
rect 110 1949 111 1953
rect 115 1949 116 1953
rect 110 1948 116 1949
rect 1822 1953 1828 1954
rect 1822 1949 1823 1953
rect 1827 1949 1828 1953
rect 1862 1953 1863 1957
rect 1867 1953 1868 1957
rect 1862 1952 1868 1953
rect 3574 1957 3580 1958
rect 3574 1953 3575 1957
rect 3579 1953 3580 1957
rect 3574 1952 3580 1953
rect 1822 1948 1828 1949
rect 1862 1940 1868 1941
rect 110 1936 116 1937
rect 110 1932 111 1936
rect 115 1932 116 1936
rect 110 1931 116 1932
rect 1822 1936 1828 1937
rect 1822 1932 1823 1936
rect 1827 1932 1828 1936
rect 1862 1936 1863 1940
rect 1867 1936 1868 1940
rect 1862 1935 1868 1936
rect 3574 1940 3580 1941
rect 3574 1936 3575 1940
rect 3579 1936 3580 1940
rect 3574 1935 3580 1936
rect 1822 1931 1828 1932
rect 112 1899 114 1931
rect 166 1923 172 1924
rect 166 1919 167 1923
rect 171 1919 172 1923
rect 166 1918 172 1919
rect 302 1923 308 1924
rect 302 1919 303 1923
rect 307 1919 308 1923
rect 302 1918 308 1919
rect 446 1923 452 1924
rect 446 1919 447 1923
rect 451 1919 452 1923
rect 446 1918 452 1919
rect 590 1923 596 1924
rect 590 1919 591 1923
rect 595 1919 596 1923
rect 590 1918 596 1919
rect 726 1923 732 1924
rect 726 1919 727 1923
rect 731 1919 732 1923
rect 726 1918 732 1919
rect 862 1923 868 1924
rect 862 1919 863 1923
rect 867 1919 868 1923
rect 862 1918 868 1919
rect 998 1923 1004 1924
rect 998 1919 999 1923
rect 1003 1919 1004 1923
rect 998 1918 1004 1919
rect 1126 1923 1132 1924
rect 1126 1919 1127 1923
rect 1131 1919 1132 1923
rect 1126 1918 1132 1919
rect 1246 1923 1252 1924
rect 1246 1919 1247 1923
rect 1251 1919 1252 1923
rect 1246 1918 1252 1919
rect 1366 1923 1372 1924
rect 1366 1919 1367 1923
rect 1371 1919 1372 1923
rect 1366 1918 1372 1919
rect 1486 1923 1492 1924
rect 1486 1919 1487 1923
rect 1491 1919 1492 1923
rect 1486 1918 1492 1919
rect 1606 1923 1612 1924
rect 1606 1919 1607 1923
rect 1611 1919 1612 1923
rect 1606 1918 1612 1919
rect 168 1899 170 1918
rect 304 1899 306 1918
rect 448 1899 450 1918
rect 592 1899 594 1918
rect 728 1899 730 1918
rect 864 1899 866 1918
rect 1000 1899 1002 1918
rect 1128 1899 1130 1918
rect 1248 1899 1250 1918
rect 1368 1899 1370 1918
rect 1488 1899 1490 1918
rect 1608 1899 1610 1918
rect 1824 1899 1826 1931
rect 1864 1911 1866 1935
rect 1910 1927 1916 1928
rect 1910 1923 1911 1927
rect 1915 1923 1916 1927
rect 1910 1922 1916 1923
rect 2166 1927 2172 1928
rect 2166 1923 2167 1927
rect 2171 1923 2172 1927
rect 2166 1922 2172 1923
rect 2406 1927 2412 1928
rect 2406 1923 2407 1927
rect 2411 1923 2412 1927
rect 2406 1922 2412 1923
rect 2622 1927 2628 1928
rect 2622 1923 2623 1927
rect 2627 1923 2628 1927
rect 2622 1922 2628 1923
rect 2822 1927 2828 1928
rect 2822 1923 2823 1927
rect 2827 1923 2828 1927
rect 2822 1922 2828 1923
rect 3006 1927 3012 1928
rect 3006 1923 3007 1927
rect 3011 1923 3012 1927
rect 3006 1922 3012 1923
rect 3174 1927 3180 1928
rect 3174 1923 3175 1927
rect 3179 1923 3180 1927
rect 3174 1922 3180 1923
rect 3342 1927 3348 1928
rect 3342 1923 3343 1927
rect 3347 1923 3348 1927
rect 3342 1922 3348 1923
rect 3486 1927 3492 1928
rect 3486 1923 3487 1927
rect 3491 1923 3492 1927
rect 3486 1922 3492 1923
rect 1912 1911 1914 1922
rect 2168 1911 2170 1922
rect 2408 1911 2410 1922
rect 2624 1911 2626 1922
rect 2824 1911 2826 1922
rect 3008 1911 3010 1922
rect 3176 1911 3178 1922
rect 3344 1911 3346 1922
rect 3488 1911 3490 1922
rect 3576 1911 3578 1935
rect 1863 1910 1867 1911
rect 1863 1905 1867 1906
rect 1895 1910 1899 1911
rect 1895 1905 1899 1906
rect 1911 1910 1915 1911
rect 1911 1905 1915 1906
rect 1983 1910 1987 1911
rect 1983 1905 1987 1906
rect 2071 1910 2075 1911
rect 2071 1905 2075 1906
rect 2167 1910 2171 1911
rect 2167 1905 2171 1906
rect 2295 1910 2299 1911
rect 2295 1905 2299 1906
rect 2407 1910 2411 1911
rect 2407 1905 2411 1906
rect 2447 1910 2451 1911
rect 2447 1905 2451 1906
rect 2607 1910 2611 1911
rect 2607 1905 2611 1906
rect 2623 1910 2627 1911
rect 2623 1905 2627 1906
rect 2767 1910 2771 1911
rect 2767 1905 2771 1906
rect 2823 1910 2827 1911
rect 2823 1905 2827 1906
rect 2919 1910 2923 1911
rect 2919 1905 2923 1906
rect 3007 1910 3011 1911
rect 3007 1905 3011 1906
rect 3071 1910 3075 1911
rect 3071 1905 3075 1906
rect 3175 1910 3179 1911
rect 3175 1905 3179 1906
rect 3215 1910 3219 1911
rect 3215 1905 3219 1906
rect 3343 1910 3347 1911
rect 3343 1905 3347 1906
rect 3359 1910 3363 1911
rect 3359 1905 3363 1906
rect 3487 1910 3491 1911
rect 3487 1905 3491 1906
rect 3575 1910 3579 1911
rect 3575 1905 3579 1906
rect 111 1898 115 1899
rect 111 1893 115 1894
rect 167 1898 171 1899
rect 167 1893 171 1894
rect 223 1898 227 1899
rect 223 1893 227 1894
rect 303 1898 307 1899
rect 303 1893 307 1894
rect 447 1898 451 1899
rect 447 1893 451 1894
rect 479 1898 483 1899
rect 479 1893 483 1894
rect 591 1898 595 1899
rect 591 1893 595 1894
rect 719 1898 723 1899
rect 719 1893 723 1894
rect 727 1898 731 1899
rect 727 1893 731 1894
rect 863 1898 867 1899
rect 863 1893 867 1894
rect 935 1898 939 1899
rect 935 1893 939 1894
rect 999 1898 1003 1899
rect 999 1893 1003 1894
rect 1127 1898 1131 1899
rect 1127 1893 1131 1894
rect 1247 1898 1251 1899
rect 1247 1893 1251 1894
rect 1295 1898 1299 1899
rect 1295 1893 1299 1894
rect 1367 1898 1371 1899
rect 1367 1893 1371 1894
rect 1455 1898 1459 1899
rect 1455 1893 1459 1894
rect 1487 1898 1491 1899
rect 1487 1893 1491 1894
rect 1607 1898 1611 1899
rect 1607 1893 1611 1894
rect 1735 1898 1739 1899
rect 1735 1893 1739 1894
rect 1823 1898 1827 1899
rect 1823 1893 1827 1894
rect 112 1869 114 1893
rect 224 1882 226 1893
rect 480 1882 482 1893
rect 720 1882 722 1893
rect 936 1882 938 1893
rect 1128 1882 1130 1893
rect 1296 1882 1298 1893
rect 1456 1882 1458 1893
rect 1608 1882 1610 1893
rect 1736 1882 1738 1893
rect 222 1881 228 1882
rect 222 1877 223 1881
rect 227 1877 228 1881
rect 222 1876 228 1877
rect 478 1881 484 1882
rect 478 1877 479 1881
rect 483 1877 484 1881
rect 478 1876 484 1877
rect 718 1881 724 1882
rect 718 1877 719 1881
rect 723 1877 724 1881
rect 718 1876 724 1877
rect 934 1881 940 1882
rect 934 1877 935 1881
rect 939 1877 940 1881
rect 934 1876 940 1877
rect 1126 1881 1132 1882
rect 1126 1877 1127 1881
rect 1131 1877 1132 1881
rect 1126 1876 1132 1877
rect 1294 1881 1300 1882
rect 1294 1877 1295 1881
rect 1299 1877 1300 1881
rect 1294 1876 1300 1877
rect 1454 1881 1460 1882
rect 1454 1877 1455 1881
rect 1459 1877 1460 1881
rect 1454 1876 1460 1877
rect 1606 1881 1612 1882
rect 1606 1877 1607 1881
rect 1611 1877 1612 1881
rect 1606 1876 1612 1877
rect 1734 1881 1740 1882
rect 1734 1877 1735 1881
rect 1739 1877 1740 1881
rect 1734 1876 1740 1877
rect 1824 1869 1826 1893
rect 1864 1881 1866 1905
rect 1896 1894 1898 1905
rect 1984 1894 1986 1905
rect 2072 1894 2074 1905
rect 2168 1894 2170 1905
rect 2296 1894 2298 1905
rect 2448 1894 2450 1905
rect 2608 1894 2610 1905
rect 2768 1894 2770 1905
rect 2920 1894 2922 1905
rect 3072 1894 3074 1905
rect 3216 1894 3218 1905
rect 3360 1894 3362 1905
rect 3488 1894 3490 1905
rect 1894 1893 1900 1894
rect 1894 1889 1895 1893
rect 1899 1889 1900 1893
rect 1894 1888 1900 1889
rect 1982 1893 1988 1894
rect 1982 1889 1983 1893
rect 1987 1889 1988 1893
rect 1982 1888 1988 1889
rect 2070 1893 2076 1894
rect 2070 1889 2071 1893
rect 2075 1889 2076 1893
rect 2070 1888 2076 1889
rect 2166 1893 2172 1894
rect 2166 1889 2167 1893
rect 2171 1889 2172 1893
rect 2166 1888 2172 1889
rect 2294 1893 2300 1894
rect 2294 1889 2295 1893
rect 2299 1889 2300 1893
rect 2294 1888 2300 1889
rect 2446 1893 2452 1894
rect 2446 1889 2447 1893
rect 2451 1889 2452 1893
rect 2446 1888 2452 1889
rect 2606 1893 2612 1894
rect 2606 1889 2607 1893
rect 2611 1889 2612 1893
rect 2606 1888 2612 1889
rect 2766 1893 2772 1894
rect 2766 1889 2767 1893
rect 2771 1889 2772 1893
rect 2766 1888 2772 1889
rect 2918 1893 2924 1894
rect 2918 1889 2919 1893
rect 2923 1889 2924 1893
rect 2918 1888 2924 1889
rect 3070 1893 3076 1894
rect 3070 1889 3071 1893
rect 3075 1889 3076 1893
rect 3070 1888 3076 1889
rect 3214 1893 3220 1894
rect 3214 1889 3215 1893
rect 3219 1889 3220 1893
rect 3214 1888 3220 1889
rect 3358 1893 3364 1894
rect 3358 1889 3359 1893
rect 3363 1889 3364 1893
rect 3358 1888 3364 1889
rect 3486 1893 3492 1894
rect 3486 1889 3487 1893
rect 3491 1889 3492 1893
rect 3486 1888 3492 1889
rect 3576 1881 3578 1905
rect 1862 1880 1868 1881
rect 1862 1876 1863 1880
rect 1867 1876 1868 1880
rect 1862 1875 1868 1876
rect 3574 1880 3580 1881
rect 3574 1876 3575 1880
rect 3579 1876 3580 1880
rect 3574 1875 3580 1876
rect 110 1868 116 1869
rect 110 1864 111 1868
rect 115 1864 116 1868
rect 110 1863 116 1864
rect 1822 1868 1828 1869
rect 1822 1864 1823 1868
rect 1827 1864 1828 1868
rect 1822 1863 1828 1864
rect 1862 1863 1868 1864
rect 1862 1859 1863 1863
rect 1867 1859 1868 1863
rect 1862 1858 1868 1859
rect 3574 1863 3580 1864
rect 3574 1859 3575 1863
rect 3579 1859 3580 1863
rect 3574 1858 3580 1859
rect 110 1851 116 1852
rect 110 1847 111 1851
rect 115 1847 116 1851
rect 110 1846 116 1847
rect 1822 1851 1828 1852
rect 1822 1847 1823 1851
rect 1827 1847 1828 1851
rect 1822 1846 1828 1847
rect 112 1831 114 1846
rect 214 1841 220 1842
rect 214 1837 215 1841
rect 219 1837 220 1841
rect 214 1836 220 1837
rect 470 1841 476 1842
rect 470 1837 471 1841
rect 475 1837 476 1841
rect 470 1836 476 1837
rect 710 1841 716 1842
rect 710 1837 711 1841
rect 715 1837 716 1841
rect 710 1836 716 1837
rect 926 1841 932 1842
rect 926 1837 927 1841
rect 931 1837 932 1841
rect 926 1836 932 1837
rect 1118 1841 1124 1842
rect 1118 1837 1119 1841
rect 1123 1837 1124 1841
rect 1118 1836 1124 1837
rect 1286 1841 1292 1842
rect 1286 1837 1287 1841
rect 1291 1837 1292 1841
rect 1286 1836 1292 1837
rect 1446 1841 1452 1842
rect 1446 1837 1447 1841
rect 1451 1837 1452 1841
rect 1446 1836 1452 1837
rect 1598 1841 1604 1842
rect 1598 1837 1599 1841
rect 1603 1837 1604 1841
rect 1598 1836 1604 1837
rect 1726 1841 1732 1842
rect 1726 1837 1727 1841
rect 1731 1837 1732 1841
rect 1726 1836 1732 1837
rect 216 1831 218 1836
rect 472 1831 474 1836
rect 712 1831 714 1836
rect 928 1831 930 1836
rect 1120 1831 1122 1836
rect 1288 1831 1290 1836
rect 1448 1831 1450 1836
rect 1600 1831 1602 1836
rect 1728 1831 1730 1836
rect 1824 1831 1826 1846
rect 1864 1839 1866 1858
rect 1886 1853 1892 1854
rect 1886 1849 1887 1853
rect 1891 1849 1892 1853
rect 1886 1848 1892 1849
rect 1974 1853 1980 1854
rect 1974 1849 1975 1853
rect 1979 1849 1980 1853
rect 1974 1848 1980 1849
rect 2062 1853 2068 1854
rect 2062 1849 2063 1853
rect 2067 1849 2068 1853
rect 2062 1848 2068 1849
rect 2158 1853 2164 1854
rect 2158 1849 2159 1853
rect 2163 1849 2164 1853
rect 2158 1848 2164 1849
rect 2286 1853 2292 1854
rect 2286 1849 2287 1853
rect 2291 1849 2292 1853
rect 2286 1848 2292 1849
rect 2438 1853 2444 1854
rect 2438 1849 2439 1853
rect 2443 1849 2444 1853
rect 2438 1848 2444 1849
rect 2598 1853 2604 1854
rect 2598 1849 2599 1853
rect 2603 1849 2604 1853
rect 2598 1848 2604 1849
rect 2758 1853 2764 1854
rect 2758 1849 2759 1853
rect 2763 1849 2764 1853
rect 2758 1848 2764 1849
rect 2910 1853 2916 1854
rect 2910 1849 2911 1853
rect 2915 1849 2916 1853
rect 2910 1848 2916 1849
rect 3062 1853 3068 1854
rect 3062 1849 3063 1853
rect 3067 1849 3068 1853
rect 3062 1848 3068 1849
rect 3206 1853 3212 1854
rect 3206 1849 3207 1853
rect 3211 1849 3212 1853
rect 3206 1848 3212 1849
rect 3350 1853 3356 1854
rect 3350 1849 3351 1853
rect 3355 1849 3356 1853
rect 3350 1848 3356 1849
rect 3478 1853 3484 1854
rect 3478 1849 3479 1853
rect 3483 1849 3484 1853
rect 3478 1848 3484 1849
rect 1888 1839 1890 1848
rect 1976 1839 1978 1848
rect 2064 1839 2066 1848
rect 2160 1839 2162 1848
rect 2288 1839 2290 1848
rect 2440 1839 2442 1848
rect 2600 1839 2602 1848
rect 2760 1839 2762 1848
rect 2912 1839 2914 1848
rect 3064 1839 3066 1848
rect 3208 1839 3210 1848
rect 3352 1839 3354 1848
rect 3480 1839 3482 1848
rect 3576 1839 3578 1858
rect 1863 1838 1867 1839
rect 1863 1833 1867 1834
rect 1887 1838 1891 1839
rect 1887 1833 1891 1834
rect 1975 1838 1979 1839
rect 1975 1833 1979 1834
rect 1999 1838 2003 1839
rect 1999 1833 2003 1834
rect 2063 1838 2067 1839
rect 2063 1833 2067 1834
rect 2159 1838 2163 1839
rect 2159 1833 2163 1834
rect 2223 1838 2227 1839
rect 2223 1833 2227 1834
rect 2287 1838 2291 1839
rect 2287 1833 2291 1834
rect 2439 1838 2443 1839
rect 2439 1833 2443 1834
rect 2599 1838 2603 1839
rect 2599 1833 2603 1834
rect 2639 1838 2643 1839
rect 2639 1833 2643 1834
rect 2759 1838 2763 1839
rect 2759 1833 2763 1834
rect 2831 1838 2835 1839
rect 2831 1833 2835 1834
rect 2911 1838 2915 1839
rect 2911 1833 2915 1834
rect 3015 1838 3019 1839
rect 3015 1833 3019 1834
rect 3063 1838 3067 1839
rect 3063 1833 3067 1834
rect 3199 1838 3203 1839
rect 3199 1833 3203 1834
rect 3207 1838 3211 1839
rect 3207 1833 3211 1834
rect 3351 1838 3355 1839
rect 3351 1833 3355 1834
rect 3391 1838 3395 1839
rect 3391 1833 3395 1834
rect 3479 1838 3483 1839
rect 3479 1833 3483 1834
rect 3575 1838 3579 1839
rect 3575 1833 3579 1834
rect 111 1830 115 1831
rect 111 1825 115 1826
rect 215 1830 219 1831
rect 215 1825 219 1826
rect 247 1830 251 1831
rect 247 1825 251 1826
rect 415 1830 419 1831
rect 415 1825 419 1826
rect 471 1830 475 1831
rect 471 1825 475 1826
rect 591 1830 595 1831
rect 591 1825 595 1826
rect 711 1830 715 1831
rect 711 1825 715 1826
rect 759 1830 763 1831
rect 759 1825 763 1826
rect 927 1830 931 1831
rect 927 1825 931 1826
rect 1079 1830 1083 1831
rect 1079 1825 1083 1826
rect 1119 1830 1123 1831
rect 1119 1825 1123 1826
rect 1223 1830 1227 1831
rect 1223 1825 1227 1826
rect 1287 1830 1291 1831
rect 1287 1825 1291 1826
rect 1359 1830 1363 1831
rect 1359 1825 1363 1826
rect 1447 1830 1451 1831
rect 1447 1825 1451 1826
rect 1487 1830 1491 1831
rect 1487 1825 1491 1826
rect 1599 1830 1603 1831
rect 1599 1825 1603 1826
rect 1615 1830 1619 1831
rect 1615 1825 1619 1826
rect 1727 1830 1731 1831
rect 1727 1825 1731 1826
rect 1823 1830 1827 1831
rect 1823 1825 1827 1826
rect 112 1810 114 1825
rect 248 1820 250 1825
rect 416 1820 418 1825
rect 592 1820 594 1825
rect 760 1820 762 1825
rect 928 1820 930 1825
rect 1080 1820 1082 1825
rect 1224 1820 1226 1825
rect 1360 1820 1362 1825
rect 1488 1820 1490 1825
rect 1616 1820 1618 1825
rect 1728 1820 1730 1825
rect 246 1819 252 1820
rect 246 1815 247 1819
rect 251 1815 252 1819
rect 246 1814 252 1815
rect 414 1819 420 1820
rect 414 1815 415 1819
rect 419 1815 420 1819
rect 414 1814 420 1815
rect 590 1819 596 1820
rect 590 1815 591 1819
rect 595 1815 596 1819
rect 590 1814 596 1815
rect 758 1819 764 1820
rect 758 1815 759 1819
rect 763 1815 764 1819
rect 758 1814 764 1815
rect 926 1819 932 1820
rect 926 1815 927 1819
rect 931 1815 932 1819
rect 926 1814 932 1815
rect 1078 1819 1084 1820
rect 1078 1815 1079 1819
rect 1083 1815 1084 1819
rect 1078 1814 1084 1815
rect 1222 1819 1228 1820
rect 1222 1815 1223 1819
rect 1227 1815 1228 1819
rect 1222 1814 1228 1815
rect 1358 1819 1364 1820
rect 1358 1815 1359 1819
rect 1363 1815 1364 1819
rect 1358 1814 1364 1815
rect 1486 1819 1492 1820
rect 1486 1815 1487 1819
rect 1491 1815 1492 1819
rect 1486 1814 1492 1815
rect 1614 1819 1620 1820
rect 1614 1815 1615 1819
rect 1619 1815 1620 1819
rect 1614 1814 1620 1815
rect 1726 1819 1732 1820
rect 1726 1815 1727 1819
rect 1731 1815 1732 1819
rect 1726 1814 1732 1815
rect 1824 1810 1826 1825
rect 1864 1818 1866 1833
rect 2000 1828 2002 1833
rect 2224 1828 2226 1833
rect 2440 1828 2442 1833
rect 2640 1828 2642 1833
rect 2832 1828 2834 1833
rect 3016 1828 3018 1833
rect 3200 1828 3202 1833
rect 3392 1828 3394 1833
rect 1998 1827 2004 1828
rect 1998 1823 1999 1827
rect 2003 1823 2004 1827
rect 1998 1822 2004 1823
rect 2222 1827 2228 1828
rect 2222 1823 2223 1827
rect 2227 1823 2228 1827
rect 2222 1822 2228 1823
rect 2438 1827 2444 1828
rect 2438 1823 2439 1827
rect 2443 1823 2444 1827
rect 2438 1822 2444 1823
rect 2638 1827 2644 1828
rect 2638 1823 2639 1827
rect 2643 1823 2644 1827
rect 2638 1822 2644 1823
rect 2830 1827 2836 1828
rect 2830 1823 2831 1827
rect 2835 1823 2836 1827
rect 2830 1822 2836 1823
rect 3014 1827 3020 1828
rect 3014 1823 3015 1827
rect 3019 1823 3020 1827
rect 3014 1822 3020 1823
rect 3198 1827 3204 1828
rect 3198 1823 3199 1827
rect 3203 1823 3204 1827
rect 3198 1822 3204 1823
rect 3390 1827 3396 1828
rect 3390 1823 3391 1827
rect 3395 1823 3396 1827
rect 3390 1822 3396 1823
rect 3576 1818 3578 1833
rect 1862 1817 1868 1818
rect 1862 1813 1863 1817
rect 1867 1813 1868 1817
rect 1862 1812 1868 1813
rect 3574 1817 3580 1818
rect 3574 1813 3575 1817
rect 3579 1813 3580 1817
rect 3574 1812 3580 1813
rect 110 1809 116 1810
rect 110 1805 111 1809
rect 115 1805 116 1809
rect 110 1804 116 1805
rect 1822 1809 1828 1810
rect 1822 1805 1823 1809
rect 1827 1805 1828 1809
rect 1822 1804 1828 1805
rect 1862 1800 1868 1801
rect 1862 1796 1863 1800
rect 1867 1796 1868 1800
rect 1862 1795 1868 1796
rect 3574 1800 3580 1801
rect 3574 1796 3575 1800
rect 3579 1796 3580 1800
rect 3574 1795 3580 1796
rect 110 1792 116 1793
rect 110 1788 111 1792
rect 115 1788 116 1792
rect 110 1787 116 1788
rect 1822 1792 1828 1793
rect 1822 1788 1823 1792
rect 1827 1788 1828 1792
rect 1822 1787 1828 1788
rect 112 1759 114 1787
rect 254 1779 260 1780
rect 254 1775 255 1779
rect 259 1775 260 1779
rect 254 1774 260 1775
rect 422 1779 428 1780
rect 422 1775 423 1779
rect 427 1775 428 1779
rect 422 1774 428 1775
rect 598 1779 604 1780
rect 598 1775 599 1779
rect 603 1775 604 1779
rect 598 1774 604 1775
rect 766 1779 772 1780
rect 766 1775 767 1779
rect 771 1775 772 1779
rect 766 1774 772 1775
rect 934 1779 940 1780
rect 934 1775 935 1779
rect 939 1775 940 1779
rect 934 1774 940 1775
rect 1086 1779 1092 1780
rect 1086 1775 1087 1779
rect 1091 1775 1092 1779
rect 1086 1774 1092 1775
rect 1230 1779 1236 1780
rect 1230 1775 1231 1779
rect 1235 1775 1236 1779
rect 1230 1774 1236 1775
rect 1366 1779 1372 1780
rect 1366 1775 1367 1779
rect 1371 1775 1372 1779
rect 1366 1774 1372 1775
rect 1494 1779 1500 1780
rect 1494 1775 1495 1779
rect 1499 1775 1500 1779
rect 1494 1774 1500 1775
rect 1622 1779 1628 1780
rect 1622 1775 1623 1779
rect 1627 1775 1628 1779
rect 1622 1774 1628 1775
rect 1734 1779 1740 1780
rect 1734 1775 1735 1779
rect 1739 1775 1740 1779
rect 1734 1774 1740 1775
rect 256 1759 258 1774
rect 424 1759 426 1774
rect 600 1759 602 1774
rect 768 1759 770 1774
rect 936 1759 938 1774
rect 1088 1759 1090 1774
rect 1232 1759 1234 1774
rect 1368 1759 1370 1774
rect 1496 1759 1498 1774
rect 1624 1759 1626 1774
rect 1736 1759 1738 1774
rect 1824 1759 1826 1787
rect 1864 1767 1866 1795
rect 2006 1787 2012 1788
rect 2006 1783 2007 1787
rect 2011 1783 2012 1787
rect 2006 1782 2012 1783
rect 2230 1787 2236 1788
rect 2230 1783 2231 1787
rect 2235 1783 2236 1787
rect 2230 1782 2236 1783
rect 2446 1787 2452 1788
rect 2446 1783 2447 1787
rect 2451 1783 2452 1787
rect 2446 1782 2452 1783
rect 2646 1787 2652 1788
rect 2646 1783 2647 1787
rect 2651 1783 2652 1787
rect 2646 1782 2652 1783
rect 2838 1787 2844 1788
rect 2838 1783 2839 1787
rect 2843 1783 2844 1787
rect 2838 1782 2844 1783
rect 3022 1787 3028 1788
rect 3022 1783 3023 1787
rect 3027 1783 3028 1787
rect 3022 1782 3028 1783
rect 3206 1787 3212 1788
rect 3206 1783 3207 1787
rect 3211 1783 3212 1787
rect 3206 1782 3212 1783
rect 3398 1787 3404 1788
rect 3398 1783 3399 1787
rect 3403 1783 3404 1787
rect 3398 1782 3404 1783
rect 2008 1767 2010 1782
rect 2232 1767 2234 1782
rect 2448 1767 2450 1782
rect 2648 1767 2650 1782
rect 2840 1767 2842 1782
rect 3024 1767 3026 1782
rect 3208 1767 3210 1782
rect 3400 1767 3402 1782
rect 3576 1767 3578 1795
rect 1863 1766 1867 1767
rect 1863 1761 1867 1762
rect 1943 1766 1947 1767
rect 1943 1761 1947 1762
rect 2007 1766 2011 1767
rect 2007 1761 2011 1762
rect 2087 1766 2091 1767
rect 2087 1761 2091 1762
rect 2231 1766 2235 1767
rect 2231 1761 2235 1762
rect 2247 1766 2251 1767
rect 2247 1761 2251 1762
rect 2415 1766 2419 1767
rect 2415 1761 2419 1762
rect 2447 1766 2451 1767
rect 2447 1761 2451 1762
rect 2599 1766 2603 1767
rect 2599 1761 2603 1762
rect 2647 1766 2651 1767
rect 2647 1761 2651 1762
rect 2791 1766 2795 1767
rect 2791 1761 2795 1762
rect 2839 1766 2843 1767
rect 2839 1761 2843 1762
rect 2991 1766 2995 1767
rect 2991 1761 2995 1762
rect 3023 1766 3027 1767
rect 3023 1761 3027 1762
rect 3199 1766 3203 1767
rect 3199 1761 3203 1762
rect 3207 1766 3211 1767
rect 3207 1761 3211 1762
rect 3399 1766 3403 1767
rect 3399 1761 3403 1762
rect 3415 1766 3419 1767
rect 3415 1761 3419 1762
rect 3575 1766 3579 1767
rect 3575 1761 3579 1762
rect 111 1758 115 1759
rect 111 1753 115 1754
rect 255 1758 259 1759
rect 255 1753 259 1754
rect 327 1758 331 1759
rect 327 1753 331 1754
rect 423 1758 427 1759
rect 423 1753 427 1754
rect 471 1758 475 1759
rect 471 1753 475 1754
rect 599 1758 603 1759
rect 599 1753 603 1754
rect 615 1758 619 1759
rect 615 1753 619 1754
rect 767 1758 771 1759
rect 767 1753 771 1754
rect 919 1758 923 1759
rect 919 1753 923 1754
rect 935 1758 939 1759
rect 935 1753 939 1754
rect 1071 1758 1075 1759
rect 1071 1753 1075 1754
rect 1087 1758 1091 1759
rect 1087 1753 1091 1754
rect 1223 1758 1227 1759
rect 1223 1753 1227 1754
rect 1231 1758 1235 1759
rect 1231 1753 1235 1754
rect 1367 1758 1371 1759
rect 1367 1753 1371 1754
rect 1375 1758 1379 1759
rect 1375 1753 1379 1754
rect 1495 1758 1499 1759
rect 1495 1753 1499 1754
rect 1527 1758 1531 1759
rect 1527 1753 1531 1754
rect 1623 1758 1627 1759
rect 1623 1753 1627 1754
rect 1687 1758 1691 1759
rect 1687 1753 1691 1754
rect 1735 1758 1739 1759
rect 1735 1753 1739 1754
rect 1823 1758 1827 1759
rect 1823 1753 1827 1754
rect 112 1729 114 1753
rect 328 1742 330 1753
rect 472 1742 474 1753
rect 616 1742 618 1753
rect 768 1742 770 1753
rect 920 1742 922 1753
rect 1072 1742 1074 1753
rect 1224 1742 1226 1753
rect 1376 1742 1378 1753
rect 1528 1742 1530 1753
rect 1688 1742 1690 1753
rect 326 1741 332 1742
rect 326 1737 327 1741
rect 331 1737 332 1741
rect 326 1736 332 1737
rect 470 1741 476 1742
rect 470 1737 471 1741
rect 475 1737 476 1741
rect 470 1736 476 1737
rect 614 1741 620 1742
rect 614 1737 615 1741
rect 619 1737 620 1741
rect 614 1736 620 1737
rect 766 1741 772 1742
rect 766 1737 767 1741
rect 771 1737 772 1741
rect 766 1736 772 1737
rect 918 1741 924 1742
rect 918 1737 919 1741
rect 923 1737 924 1741
rect 918 1736 924 1737
rect 1070 1741 1076 1742
rect 1070 1737 1071 1741
rect 1075 1737 1076 1741
rect 1070 1736 1076 1737
rect 1222 1741 1228 1742
rect 1222 1737 1223 1741
rect 1227 1737 1228 1741
rect 1222 1736 1228 1737
rect 1374 1741 1380 1742
rect 1374 1737 1375 1741
rect 1379 1737 1380 1741
rect 1374 1736 1380 1737
rect 1526 1741 1532 1742
rect 1526 1737 1527 1741
rect 1531 1737 1532 1741
rect 1526 1736 1532 1737
rect 1686 1741 1692 1742
rect 1686 1737 1687 1741
rect 1691 1737 1692 1741
rect 1686 1736 1692 1737
rect 1824 1729 1826 1753
rect 1864 1737 1866 1761
rect 1944 1750 1946 1761
rect 2088 1750 2090 1761
rect 2248 1750 2250 1761
rect 2416 1750 2418 1761
rect 2600 1750 2602 1761
rect 2792 1750 2794 1761
rect 2992 1750 2994 1761
rect 3200 1750 3202 1761
rect 3416 1750 3418 1761
rect 1942 1749 1948 1750
rect 1942 1745 1943 1749
rect 1947 1745 1948 1749
rect 1942 1744 1948 1745
rect 2086 1749 2092 1750
rect 2086 1745 2087 1749
rect 2091 1745 2092 1749
rect 2086 1744 2092 1745
rect 2246 1749 2252 1750
rect 2246 1745 2247 1749
rect 2251 1745 2252 1749
rect 2246 1744 2252 1745
rect 2414 1749 2420 1750
rect 2414 1745 2415 1749
rect 2419 1745 2420 1749
rect 2414 1744 2420 1745
rect 2598 1749 2604 1750
rect 2598 1745 2599 1749
rect 2603 1745 2604 1749
rect 2598 1744 2604 1745
rect 2790 1749 2796 1750
rect 2790 1745 2791 1749
rect 2795 1745 2796 1749
rect 2790 1744 2796 1745
rect 2990 1749 2996 1750
rect 2990 1745 2991 1749
rect 2995 1745 2996 1749
rect 2990 1744 2996 1745
rect 3198 1749 3204 1750
rect 3198 1745 3199 1749
rect 3203 1745 3204 1749
rect 3198 1744 3204 1745
rect 3414 1749 3420 1750
rect 3414 1745 3415 1749
rect 3419 1745 3420 1749
rect 3414 1744 3420 1745
rect 3576 1737 3578 1761
rect 1862 1736 1868 1737
rect 1862 1732 1863 1736
rect 1867 1732 1868 1736
rect 1862 1731 1868 1732
rect 3574 1736 3580 1737
rect 3574 1732 3575 1736
rect 3579 1732 3580 1736
rect 3574 1731 3580 1732
rect 110 1728 116 1729
rect 110 1724 111 1728
rect 115 1724 116 1728
rect 110 1723 116 1724
rect 1822 1728 1828 1729
rect 1822 1724 1823 1728
rect 1827 1724 1828 1728
rect 1822 1723 1828 1724
rect 1862 1719 1868 1720
rect 1862 1715 1863 1719
rect 1867 1715 1868 1719
rect 1862 1714 1868 1715
rect 3574 1719 3580 1720
rect 3574 1715 3575 1719
rect 3579 1715 3580 1719
rect 3574 1714 3580 1715
rect 110 1711 116 1712
rect 110 1707 111 1711
rect 115 1707 116 1711
rect 110 1706 116 1707
rect 1822 1711 1828 1712
rect 1822 1707 1823 1711
rect 1827 1707 1828 1711
rect 1822 1706 1828 1707
rect 112 1687 114 1706
rect 318 1701 324 1702
rect 318 1697 319 1701
rect 323 1697 324 1701
rect 318 1696 324 1697
rect 462 1701 468 1702
rect 462 1697 463 1701
rect 467 1697 468 1701
rect 462 1696 468 1697
rect 606 1701 612 1702
rect 606 1697 607 1701
rect 611 1697 612 1701
rect 606 1696 612 1697
rect 758 1701 764 1702
rect 758 1697 759 1701
rect 763 1697 764 1701
rect 758 1696 764 1697
rect 910 1701 916 1702
rect 910 1697 911 1701
rect 915 1697 916 1701
rect 910 1696 916 1697
rect 1062 1701 1068 1702
rect 1062 1697 1063 1701
rect 1067 1697 1068 1701
rect 1062 1696 1068 1697
rect 1214 1701 1220 1702
rect 1214 1697 1215 1701
rect 1219 1697 1220 1701
rect 1214 1696 1220 1697
rect 1366 1701 1372 1702
rect 1366 1697 1367 1701
rect 1371 1697 1372 1701
rect 1366 1696 1372 1697
rect 1518 1701 1524 1702
rect 1518 1697 1519 1701
rect 1523 1697 1524 1701
rect 1518 1696 1524 1697
rect 1678 1701 1684 1702
rect 1678 1697 1679 1701
rect 1683 1697 1684 1701
rect 1678 1696 1684 1697
rect 320 1687 322 1696
rect 464 1687 466 1696
rect 608 1687 610 1696
rect 760 1687 762 1696
rect 912 1687 914 1696
rect 1064 1687 1066 1696
rect 1216 1687 1218 1696
rect 1368 1687 1370 1696
rect 1520 1687 1522 1696
rect 1680 1687 1682 1696
rect 1824 1687 1826 1706
rect 1864 1695 1866 1714
rect 1934 1709 1940 1710
rect 1934 1705 1935 1709
rect 1939 1705 1940 1709
rect 1934 1704 1940 1705
rect 2078 1709 2084 1710
rect 2078 1705 2079 1709
rect 2083 1705 2084 1709
rect 2078 1704 2084 1705
rect 2238 1709 2244 1710
rect 2238 1705 2239 1709
rect 2243 1705 2244 1709
rect 2238 1704 2244 1705
rect 2406 1709 2412 1710
rect 2406 1705 2407 1709
rect 2411 1705 2412 1709
rect 2406 1704 2412 1705
rect 2590 1709 2596 1710
rect 2590 1705 2591 1709
rect 2595 1705 2596 1709
rect 2590 1704 2596 1705
rect 2782 1709 2788 1710
rect 2782 1705 2783 1709
rect 2787 1705 2788 1709
rect 2782 1704 2788 1705
rect 2982 1709 2988 1710
rect 2982 1705 2983 1709
rect 2987 1705 2988 1709
rect 2982 1704 2988 1705
rect 3190 1709 3196 1710
rect 3190 1705 3191 1709
rect 3195 1705 3196 1709
rect 3190 1704 3196 1705
rect 3406 1709 3412 1710
rect 3406 1705 3407 1709
rect 3411 1705 3412 1709
rect 3406 1704 3412 1705
rect 1936 1695 1938 1704
rect 2080 1695 2082 1704
rect 2240 1695 2242 1704
rect 2408 1695 2410 1704
rect 2592 1695 2594 1704
rect 2784 1695 2786 1704
rect 2984 1695 2986 1704
rect 3192 1695 3194 1704
rect 3408 1695 3410 1704
rect 3576 1695 3578 1714
rect 1863 1694 1867 1695
rect 1863 1689 1867 1690
rect 1911 1694 1915 1695
rect 1911 1689 1915 1690
rect 1935 1694 1939 1695
rect 1935 1689 1939 1690
rect 2031 1694 2035 1695
rect 2031 1689 2035 1690
rect 2079 1694 2083 1695
rect 2079 1689 2083 1690
rect 2151 1694 2155 1695
rect 2151 1689 2155 1690
rect 2239 1694 2243 1695
rect 2239 1689 2243 1690
rect 2271 1694 2275 1695
rect 2271 1689 2275 1690
rect 2399 1694 2403 1695
rect 2399 1689 2403 1690
rect 2407 1694 2411 1695
rect 2407 1689 2411 1690
rect 2543 1694 2547 1695
rect 2543 1689 2547 1690
rect 2591 1694 2595 1695
rect 2591 1689 2595 1690
rect 2695 1694 2699 1695
rect 2695 1689 2699 1690
rect 2783 1694 2787 1695
rect 2783 1689 2787 1690
rect 2863 1694 2867 1695
rect 2863 1689 2867 1690
rect 2983 1694 2987 1695
rect 2983 1689 2987 1690
rect 3047 1694 3051 1695
rect 3047 1689 3051 1690
rect 3191 1694 3195 1695
rect 3191 1689 3195 1690
rect 3239 1694 3243 1695
rect 3239 1689 3243 1690
rect 3407 1694 3411 1695
rect 3407 1689 3411 1690
rect 3431 1694 3435 1695
rect 3431 1689 3435 1690
rect 3575 1694 3579 1695
rect 3575 1689 3579 1690
rect 111 1686 115 1687
rect 111 1681 115 1682
rect 311 1686 315 1687
rect 311 1681 315 1682
rect 319 1686 323 1687
rect 319 1681 323 1682
rect 447 1686 451 1687
rect 447 1681 451 1682
rect 463 1686 467 1687
rect 463 1681 467 1682
rect 591 1686 595 1687
rect 591 1681 595 1682
rect 607 1686 611 1687
rect 607 1681 611 1682
rect 735 1686 739 1687
rect 735 1681 739 1682
rect 759 1686 763 1687
rect 759 1681 763 1682
rect 887 1686 891 1687
rect 887 1681 891 1682
rect 911 1686 915 1687
rect 911 1681 915 1682
rect 1039 1686 1043 1687
rect 1039 1681 1043 1682
rect 1063 1686 1067 1687
rect 1063 1681 1067 1682
rect 1191 1686 1195 1687
rect 1191 1681 1195 1682
rect 1215 1686 1219 1687
rect 1215 1681 1219 1682
rect 1343 1686 1347 1687
rect 1343 1681 1347 1682
rect 1367 1686 1371 1687
rect 1367 1681 1371 1682
rect 1495 1686 1499 1687
rect 1495 1681 1499 1682
rect 1519 1686 1523 1687
rect 1519 1681 1523 1682
rect 1647 1686 1651 1687
rect 1647 1681 1651 1682
rect 1679 1686 1683 1687
rect 1679 1681 1683 1682
rect 1823 1686 1827 1687
rect 1823 1681 1827 1682
rect 112 1666 114 1681
rect 312 1676 314 1681
rect 448 1676 450 1681
rect 592 1676 594 1681
rect 736 1676 738 1681
rect 888 1676 890 1681
rect 1040 1676 1042 1681
rect 1192 1676 1194 1681
rect 1344 1676 1346 1681
rect 1496 1676 1498 1681
rect 1648 1676 1650 1681
rect 310 1675 316 1676
rect 310 1671 311 1675
rect 315 1671 316 1675
rect 310 1670 316 1671
rect 446 1675 452 1676
rect 446 1671 447 1675
rect 451 1671 452 1675
rect 446 1670 452 1671
rect 590 1675 596 1676
rect 590 1671 591 1675
rect 595 1671 596 1675
rect 590 1670 596 1671
rect 734 1675 740 1676
rect 734 1671 735 1675
rect 739 1671 740 1675
rect 734 1670 740 1671
rect 886 1675 892 1676
rect 886 1671 887 1675
rect 891 1671 892 1675
rect 886 1670 892 1671
rect 1038 1675 1044 1676
rect 1038 1671 1039 1675
rect 1043 1671 1044 1675
rect 1038 1670 1044 1671
rect 1190 1675 1196 1676
rect 1190 1671 1191 1675
rect 1195 1671 1196 1675
rect 1190 1670 1196 1671
rect 1342 1675 1348 1676
rect 1342 1671 1343 1675
rect 1347 1671 1348 1675
rect 1342 1670 1348 1671
rect 1494 1675 1500 1676
rect 1494 1671 1495 1675
rect 1499 1671 1500 1675
rect 1494 1670 1500 1671
rect 1646 1675 1652 1676
rect 1646 1671 1647 1675
rect 1651 1671 1652 1675
rect 1646 1670 1652 1671
rect 1824 1666 1826 1681
rect 1864 1674 1866 1689
rect 1912 1684 1914 1689
rect 2032 1684 2034 1689
rect 2152 1684 2154 1689
rect 2272 1684 2274 1689
rect 2400 1684 2402 1689
rect 2544 1684 2546 1689
rect 2696 1684 2698 1689
rect 2864 1684 2866 1689
rect 3048 1684 3050 1689
rect 3240 1684 3242 1689
rect 3432 1684 3434 1689
rect 1910 1683 1916 1684
rect 1910 1679 1911 1683
rect 1915 1679 1916 1683
rect 1910 1678 1916 1679
rect 2030 1683 2036 1684
rect 2030 1679 2031 1683
rect 2035 1679 2036 1683
rect 2030 1678 2036 1679
rect 2150 1683 2156 1684
rect 2150 1679 2151 1683
rect 2155 1679 2156 1683
rect 2150 1678 2156 1679
rect 2270 1683 2276 1684
rect 2270 1679 2271 1683
rect 2275 1679 2276 1683
rect 2270 1678 2276 1679
rect 2398 1683 2404 1684
rect 2398 1679 2399 1683
rect 2403 1679 2404 1683
rect 2398 1678 2404 1679
rect 2542 1683 2548 1684
rect 2542 1679 2543 1683
rect 2547 1679 2548 1683
rect 2542 1678 2548 1679
rect 2694 1683 2700 1684
rect 2694 1679 2695 1683
rect 2699 1679 2700 1683
rect 2694 1678 2700 1679
rect 2862 1683 2868 1684
rect 2862 1679 2863 1683
rect 2867 1679 2868 1683
rect 2862 1678 2868 1679
rect 3046 1683 3052 1684
rect 3046 1679 3047 1683
rect 3051 1679 3052 1683
rect 3046 1678 3052 1679
rect 3238 1683 3244 1684
rect 3238 1679 3239 1683
rect 3243 1679 3244 1683
rect 3238 1678 3244 1679
rect 3430 1683 3436 1684
rect 3430 1679 3431 1683
rect 3435 1679 3436 1683
rect 3430 1678 3436 1679
rect 3576 1674 3578 1689
rect 1862 1673 1868 1674
rect 1862 1669 1863 1673
rect 1867 1669 1868 1673
rect 1862 1668 1868 1669
rect 3574 1673 3580 1674
rect 3574 1669 3575 1673
rect 3579 1669 3580 1673
rect 3574 1668 3580 1669
rect 110 1665 116 1666
rect 110 1661 111 1665
rect 115 1661 116 1665
rect 110 1660 116 1661
rect 1822 1665 1828 1666
rect 1822 1661 1823 1665
rect 1827 1661 1828 1665
rect 1822 1660 1828 1661
rect 1862 1656 1868 1657
rect 1862 1652 1863 1656
rect 1867 1652 1868 1656
rect 1862 1651 1868 1652
rect 3574 1656 3580 1657
rect 3574 1652 3575 1656
rect 3579 1652 3580 1656
rect 3574 1651 3580 1652
rect 110 1648 116 1649
rect 110 1644 111 1648
rect 115 1644 116 1648
rect 110 1643 116 1644
rect 1822 1648 1828 1649
rect 1822 1644 1823 1648
rect 1827 1644 1828 1648
rect 1822 1643 1828 1644
rect 112 1611 114 1643
rect 318 1635 324 1636
rect 318 1631 319 1635
rect 323 1631 324 1635
rect 318 1630 324 1631
rect 454 1635 460 1636
rect 454 1631 455 1635
rect 459 1631 460 1635
rect 454 1630 460 1631
rect 598 1635 604 1636
rect 598 1631 599 1635
rect 603 1631 604 1635
rect 598 1630 604 1631
rect 742 1635 748 1636
rect 742 1631 743 1635
rect 747 1631 748 1635
rect 742 1630 748 1631
rect 894 1635 900 1636
rect 894 1631 895 1635
rect 899 1631 900 1635
rect 894 1630 900 1631
rect 1046 1635 1052 1636
rect 1046 1631 1047 1635
rect 1051 1631 1052 1635
rect 1046 1630 1052 1631
rect 1198 1635 1204 1636
rect 1198 1631 1199 1635
rect 1203 1631 1204 1635
rect 1198 1630 1204 1631
rect 1350 1635 1356 1636
rect 1350 1631 1351 1635
rect 1355 1631 1356 1635
rect 1350 1630 1356 1631
rect 1502 1635 1508 1636
rect 1502 1631 1503 1635
rect 1507 1631 1508 1635
rect 1502 1630 1508 1631
rect 1654 1635 1660 1636
rect 1654 1631 1655 1635
rect 1659 1631 1660 1635
rect 1654 1630 1660 1631
rect 320 1611 322 1630
rect 456 1611 458 1630
rect 600 1611 602 1630
rect 744 1611 746 1630
rect 896 1611 898 1630
rect 1048 1611 1050 1630
rect 1200 1611 1202 1630
rect 1352 1611 1354 1630
rect 1504 1611 1506 1630
rect 1656 1611 1658 1630
rect 1824 1611 1826 1643
rect 1864 1619 1866 1651
rect 1918 1643 1924 1644
rect 1918 1639 1919 1643
rect 1923 1639 1924 1643
rect 1918 1638 1924 1639
rect 2038 1643 2044 1644
rect 2038 1639 2039 1643
rect 2043 1639 2044 1643
rect 2038 1638 2044 1639
rect 2158 1643 2164 1644
rect 2158 1639 2159 1643
rect 2163 1639 2164 1643
rect 2158 1638 2164 1639
rect 2278 1643 2284 1644
rect 2278 1639 2279 1643
rect 2283 1639 2284 1643
rect 2278 1638 2284 1639
rect 2406 1643 2412 1644
rect 2406 1639 2407 1643
rect 2411 1639 2412 1643
rect 2406 1638 2412 1639
rect 2550 1643 2556 1644
rect 2550 1639 2551 1643
rect 2555 1639 2556 1643
rect 2550 1638 2556 1639
rect 2702 1643 2708 1644
rect 2702 1639 2703 1643
rect 2707 1639 2708 1643
rect 2702 1638 2708 1639
rect 2870 1643 2876 1644
rect 2870 1639 2871 1643
rect 2875 1639 2876 1643
rect 2870 1638 2876 1639
rect 3054 1643 3060 1644
rect 3054 1639 3055 1643
rect 3059 1639 3060 1643
rect 3054 1638 3060 1639
rect 3246 1643 3252 1644
rect 3246 1639 3247 1643
rect 3251 1639 3252 1643
rect 3246 1638 3252 1639
rect 3438 1643 3444 1644
rect 3438 1639 3439 1643
rect 3443 1639 3444 1643
rect 3438 1638 3444 1639
rect 1920 1619 1922 1638
rect 2040 1619 2042 1638
rect 2160 1619 2162 1638
rect 2280 1619 2282 1638
rect 2408 1619 2410 1638
rect 2552 1619 2554 1638
rect 2704 1619 2706 1638
rect 2872 1619 2874 1638
rect 3056 1619 3058 1638
rect 3248 1619 3250 1638
rect 3440 1619 3442 1638
rect 3576 1619 3578 1651
rect 1863 1618 1867 1619
rect 1863 1613 1867 1614
rect 1895 1618 1899 1619
rect 1895 1613 1899 1614
rect 1919 1618 1923 1619
rect 1919 1613 1923 1614
rect 2015 1618 2019 1619
rect 2015 1613 2019 1614
rect 2039 1618 2043 1619
rect 2039 1613 2043 1614
rect 2151 1618 2155 1619
rect 2151 1613 2155 1614
rect 2159 1618 2163 1619
rect 2159 1613 2163 1614
rect 2279 1618 2283 1619
rect 2279 1613 2283 1614
rect 2287 1618 2291 1619
rect 2287 1613 2291 1614
rect 2407 1618 2411 1619
rect 2407 1613 2411 1614
rect 2431 1618 2435 1619
rect 2431 1613 2435 1614
rect 2551 1618 2555 1619
rect 2551 1613 2555 1614
rect 2583 1618 2587 1619
rect 2583 1613 2587 1614
rect 2703 1618 2707 1619
rect 2703 1613 2707 1614
rect 2743 1618 2747 1619
rect 2743 1613 2747 1614
rect 2871 1618 2875 1619
rect 2871 1613 2875 1614
rect 2911 1618 2915 1619
rect 2911 1613 2915 1614
rect 3055 1618 3059 1619
rect 3055 1613 3059 1614
rect 3095 1618 3099 1619
rect 3095 1613 3099 1614
rect 3247 1618 3251 1619
rect 3247 1613 3251 1614
rect 3279 1618 3283 1619
rect 3279 1613 3283 1614
rect 3439 1618 3443 1619
rect 3439 1613 3443 1614
rect 3471 1618 3475 1619
rect 3471 1613 3475 1614
rect 3575 1618 3579 1619
rect 3575 1613 3579 1614
rect 111 1610 115 1611
rect 111 1605 115 1606
rect 223 1610 227 1611
rect 223 1605 227 1606
rect 319 1610 323 1611
rect 319 1605 323 1606
rect 351 1610 355 1611
rect 351 1605 355 1606
rect 455 1610 459 1611
rect 455 1605 459 1606
rect 487 1610 491 1611
rect 487 1605 491 1606
rect 599 1610 603 1611
rect 599 1605 603 1606
rect 623 1610 627 1611
rect 623 1605 627 1606
rect 743 1610 747 1611
rect 743 1605 747 1606
rect 759 1610 763 1611
rect 759 1605 763 1606
rect 895 1610 899 1611
rect 895 1605 899 1606
rect 903 1610 907 1611
rect 903 1605 907 1606
rect 1047 1610 1051 1611
rect 1047 1605 1051 1606
rect 1055 1610 1059 1611
rect 1055 1605 1059 1606
rect 1199 1610 1203 1611
rect 1199 1605 1203 1606
rect 1215 1610 1219 1611
rect 1215 1605 1219 1606
rect 1351 1610 1355 1611
rect 1351 1605 1355 1606
rect 1375 1610 1379 1611
rect 1375 1605 1379 1606
rect 1503 1610 1507 1611
rect 1503 1605 1507 1606
rect 1543 1610 1547 1611
rect 1543 1605 1547 1606
rect 1655 1610 1659 1611
rect 1655 1605 1659 1606
rect 1823 1610 1827 1611
rect 1823 1605 1827 1606
rect 112 1581 114 1605
rect 224 1594 226 1605
rect 352 1594 354 1605
rect 488 1594 490 1605
rect 624 1594 626 1605
rect 760 1594 762 1605
rect 904 1594 906 1605
rect 1056 1594 1058 1605
rect 1216 1594 1218 1605
rect 1376 1594 1378 1605
rect 1544 1594 1546 1605
rect 222 1593 228 1594
rect 222 1589 223 1593
rect 227 1589 228 1593
rect 222 1588 228 1589
rect 350 1593 356 1594
rect 350 1589 351 1593
rect 355 1589 356 1593
rect 350 1588 356 1589
rect 486 1593 492 1594
rect 486 1589 487 1593
rect 491 1589 492 1593
rect 486 1588 492 1589
rect 622 1593 628 1594
rect 622 1589 623 1593
rect 627 1589 628 1593
rect 622 1588 628 1589
rect 758 1593 764 1594
rect 758 1589 759 1593
rect 763 1589 764 1593
rect 758 1588 764 1589
rect 902 1593 908 1594
rect 902 1589 903 1593
rect 907 1589 908 1593
rect 902 1588 908 1589
rect 1054 1593 1060 1594
rect 1054 1589 1055 1593
rect 1059 1589 1060 1593
rect 1054 1588 1060 1589
rect 1214 1593 1220 1594
rect 1214 1589 1215 1593
rect 1219 1589 1220 1593
rect 1214 1588 1220 1589
rect 1374 1593 1380 1594
rect 1374 1589 1375 1593
rect 1379 1589 1380 1593
rect 1374 1588 1380 1589
rect 1542 1593 1548 1594
rect 1542 1589 1543 1593
rect 1547 1589 1548 1593
rect 1542 1588 1548 1589
rect 1824 1581 1826 1605
rect 1864 1589 1866 1613
rect 1896 1602 1898 1613
rect 2016 1602 2018 1613
rect 2152 1602 2154 1613
rect 2288 1602 2290 1613
rect 2432 1602 2434 1613
rect 2584 1602 2586 1613
rect 2744 1602 2746 1613
rect 2912 1602 2914 1613
rect 3096 1602 3098 1613
rect 3280 1602 3282 1613
rect 3472 1602 3474 1613
rect 1894 1601 1900 1602
rect 1894 1597 1895 1601
rect 1899 1597 1900 1601
rect 1894 1596 1900 1597
rect 2014 1601 2020 1602
rect 2014 1597 2015 1601
rect 2019 1597 2020 1601
rect 2014 1596 2020 1597
rect 2150 1601 2156 1602
rect 2150 1597 2151 1601
rect 2155 1597 2156 1601
rect 2150 1596 2156 1597
rect 2286 1601 2292 1602
rect 2286 1597 2287 1601
rect 2291 1597 2292 1601
rect 2286 1596 2292 1597
rect 2430 1601 2436 1602
rect 2430 1597 2431 1601
rect 2435 1597 2436 1601
rect 2430 1596 2436 1597
rect 2582 1601 2588 1602
rect 2582 1597 2583 1601
rect 2587 1597 2588 1601
rect 2582 1596 2588 1597
rect 2742 1601 2748 1602
rect 2742 1597 2743 1601
rect 2747 1597 2748 1601
rect 2742 1596 2748 1597
rect 2910 1601 2916 1602
rect 2910 1597 2911 1601
rect 2915 1597 2916 1601
rect 2910 1596 2916 1597
rect 3094 1601 3100 1602
rect 3094 1597 3095 1601
rect 3099 1597 3100 1601
rect 3094 1596 3100 1597
rect 3278 1601 3284 1602
rect 3278 1597 3279 1601
rect 3283 1597 3284 1601
rect 3278 1596 3284 1597
rect 3470 1601 3476 1602
rect 3470 1597 3471 1601
rect 3475 1597 3476 1601
rect 3470 1596 3476 1597
rect 3576 1589 3578 1613
rect 1862 1588 1868 1589
rect 1862 1584 1863 1588
rect 1867 1584 1868 1588
rect 1862 1583 1868 1584
rect 3574 1588 3580 1589
rect 3574 1584 3575 1588
rect 3579 1584 3580 1588
rect 3574 1583 3580 1584
rect 110 1580 116 1581
rect 110 1576 111 1580
rect 115 1576 116 1580
rect 110 1575 116 1576
rect 1822 1580 1828 1581
rect 1822 1576 1823 1580
rect 1827 1576 1828 1580
rect 1822 1575 1828 1576
rect 1862 1571 1868 1572
rect 1862 1567 1863 1571
rect 1867 1567 1868 1571
rect 1862 1566 1868 1567
rect 3574 1571 3580 1572
rect 3574 1567 3575 1571
rect 3579 1567 3580 1571
rect 3574 1566 3580 1567
rect 110 1563 116 1564
rect 110 1559 111 1563
rect 115 1559 116 1563
rect 110 1558 116 1559
rect 1822 1563 1828 1564
rect 1822 1559 1823 1563
rect 1827 1559 1828 1563
rect 1822 1558 1828 1559
rect 112 1539 114 1558
rect 214 1553 220 1554
rect 214 1549 215 1553
rect 219 1549 220 1553
rect 214 1548 220 1549
rect 342 1553 348 1554
rect 342 1549 343 1553
rect 347 1549 348 1553
rect 342 1548 348 1549
rect 478 1553 484 1554
rect 478 1549 479 1553
rect 483 1549 484 1553
rect 478 1548 484 1549
rect 614 1553 620 1554
rect 614 1549 615 1553
rect 619 1549 620 1553
rect 614 1548 620 1549
rect 750 1553 756 1554
rect 750 1549 751 1553
rect 755 1549 756 1553
rect 750 1548 756 1549
rect 894 1553 900 1554
rect 894 1549 895 1553
rect 899 1549 900 1553
rect 894 1548 900 1549
rect 1046 1553 1052 1554
rect 1046 1549 1047 1553
rect 1051 1549 1052 1553
rect 1046 1548 1052 1549
rect 1206 1553 1212 1554
rect 1206 1549 1207 1553
rect 1211 1549 1212 1553
rect 1206 1548 1212 1549
rect 1366 1553 1372 1554
rect 1366 1549 1367 1553
rect 1371 1549 1372 1553
rect 1366 1548 1372 1549
rect 1534 1553 1540 1554
rect 1534 1549 1535 1553
rect 1539 1549 1540 1553
rect 1534 1548 1540 1549
rect 216 1539 218 1548
rect 344 1539 346 1548
rect 480 1539 482 1548
rect 616 1539 618 1548
rect 752 1539 754 1548
rect 896 1539 898 1548
rect 1048 1539 1050 1548
rect 1208 1539 1210 1548
rect 1368 1539 1370 1548
rect 1536 1539 1538 1548
rect 1824 1539 1826 1558
rect 1864 1543 1866 1566
rect 1886 1561 1892 1562
rect 1886 1557 1887 1561
rect 1891 1557 1892 1561
rect 1886 1556 1892 1557
rect 2006 1561 2012 1562
rect 2006 1557 2007 1561
rect 2011 1557 2012 1561
rect 2006 1556 2012 1557
rect 2142 1561 2148 1562
rect 2142 1557 2143 1561
rect 2147 1557 2148 1561
rect 2142 1556 2148 1557
rect 2278 1561 2284 1562
rect 2278 1557 2279 1561
rect 2283 1557 2284 1561
rect 2278 1556 2284 1557
rect 2422 1561 2428 1562
rect 2422 1557 2423 1561
rect 2427 1557 2428 1561
rect 2422 1556 2428 1557
rect 2574 1561 2580 1562
rect 2574 1557 2575 1561
rect 2579 1557 2580 1561
rect 2574 1556 2580 1557
rect 2734 1561 2740 1562
rect 2734 1557 2735 1561
rect 2739 1557 2740 1561
rect 2734 1556 2740 1557
rect 2902 1561 2908 1562
rect 2902 1557 2903 1561
rect 2907 1557 2908 1561
rect 2902 1556 2908 1557
rect 3086 1561 3092 1562
rect 3086 1557 3087 1561
rect 3091 1557 3092 1561
rect 3086 1556 3092 1557
rect 3270 1561 3276 1562
rect 3270 1557 3271 1561
rect 3275 1557 3276 1561
rect 3270 1556 3276 1557
rect 3462 1561 3468 1562
rect 3462 1557 3463 1561
rect 3467 1557 3468 1561
rect 3462 1556 3468 1557
rect 1888 1543 1890 1556
rect 2008 1543 2010 1556
rect 2144 1543 2146 1556
rect 2280 1543 2282 1556
rect 2424 1543 2426 1556
rect 2576 1543 2578 1556
rect 2736 1543 2738 1556
rect 2904 1543 2906 1556
rect 3088 1543 3090 1556
rect 3272 1543 3274 1556
rect 3464 1543 3466 1556
rect 3576 1543 3578 1566
rect 1863 1542 1867 1543
rect 111 1538 115 1539
rect 111 1533 115 1534
rect 135 1538 139 1539
rect 135 1533 139 1534
rect 215 1538 219 1539
rect 215 1533 219 1534
rect 271 1538 275 1539
rect 271 1533 275 1534
rect 343 1538 347 1539
rect 343 1533 347 1534
rect 423 1538 427 1539
rect 423 1533 427 1534
rect 479 1538 483 1539
rect 479 1533 483 1534
rect 583 1538 587 1539
rect 583 1533 587 1534
rect 615 1538 619 1539
rect 615 1533 619 1534
rect 735 1538 739 1539
rect 735 1533 739 1534
rect 751 1538 755 1539
rect 751 1533 755 1534
rect 887 1538 891 1539
rect 887 1533 891 1534
rect 895 1538 899 1539
rect 895 1533 899 1534
rect 1039 1538 1043 1539
rect 1039 1533 1043 1534
rect 1047 1538 1051 1539
rect 1047 1533 1051 1534
rect 1191 1538 1195 1539
rect 1191 1533 1195 1534
rect 1207 1538 1211 1539
rect 1207 1533 1211 1534
rect 1343 1538 1347 1539
rect 1343 1533 1347 1534
rect 1367 1538 1371 1539
rect 1367 1533 1371 1534
rect 1495 1538 1499 1539
rect 1495 1533 1499 1534
rect 1535 1538 1539 1539
rect 1535 1533 1539 1534
rect 1823 1538 1827 1539
rect 1863 1537 1867 1538
rect 1887 1542 1891 1543
rect 1887 1537 1891 1538
rect 2007 1542 2011 1543
rect 2007 1537 2011 1538
rect 2023 1542 2027 1543
rect 2023 1537 2027 1538
rect 2143 1542 2147 1543
rect 2143 1537 2147 1538
rect 2183 1542 2187 1543
rect 2183 1537 2187 1538
rect 2279 1542 2283 1543
rect 2279 1537 2283 1538
rect 2343 1542 2347 1543
rect 2343 1537 2347 1538
rect 2423 1542 2427 1543
rect 2423 1537 2427 1538
rect 2503 1542 2507 1543
rect 2503 1537 2507 1538
rect 2575 1542 2579 1543
rect 2575 1537 2579 1538
rect 2663 1542 2667 1543
rect 2663 1537 2667 1538
rect 2735 1542 2739 1543
rect 2735 1537 2739 1538
rect 2823 1542 2827 1543
rect 2823 1537 2827 1538
rect 2903 1542 2907 1543
rect 2903 1537 2907 1538
rect 2983 1542 2987 1543
rect 2983 1537 2987 1538
rect 3087 1542 3091 1543
rect 3087 1537 3091 1538
rect 3151 1542 3155 1543
rect 3151 1537 3155 1538
rect 3271 1542 3275 1543
rect 3271 1537 3275 1538
rect 3319 1542 3323 1543
rect 3319 1537 3323 1538
rect 3463 1542 3467 1543
rect 3463 1537 3467 1538
rect 3479 1542 3483 1543
rect 3479 1537 3483 1538
rect 3575 1542 3579 1543
rect 3575 1537 3579 1538
rect 1823 1533 1827 1534
rect 112 1518 114 1533
rect 136 1528 138 1533
rect 272 1528 274 1533
rect 424 1528 426 1533
rect 584 1528 586 1533
rect 736 1528 738 1533
rect 888 1528 890 1533
rect 1040 1528 1042 1533
rect 1192 1528 1194 1533
rect 1344 1528 1346 1533
rect 1496 1528 1498 1533
rect 134 1527 140 1528
rect 134 1523 135 1527
rect 139 1523 140 1527
rect 134 1522 140 1523
rect 270 1527 276 1528
rect 270 1523 271 1527
rect 275 1523 276 1527
rect 270 1522 276 1523
rect 422 1527 428 1528
rect 422 1523 423 1527
rect 427 1523 428 1527
rect 422 1522 428 1523
rect 582 1527 588 1528
rect 582 1523 583 1527
rect 587 1523 588 1527
rect 582 1522 588 1523
rect 734 1527 740 1528
rect 734 1523 735 1527
rect 739 1523 740 1527
rect 734 1522 740 1523
rect 886 1527 892 1528
rect 886 1523 887 1527
rect 891 1523 892 1527
rect 886 1522 892 1523
rect 1038 1527 1044 1528
rect 1038 1523 1039 1527
rect 1043 1523 1044 1527
rect 1038 1522 1044 1523
rect 1190 1527 1196 1528
rect 1190 1523 1191 1527
rect 1195 1523 1196 1527
rect 1190 1522 1196 1523
rect 1342 1527 1348 1528
rect 1342 1523 1343 1527
rect 1347 1523 1348 1527
rect 1342 1522 1348 1523
rect 1494 1527 1500 1528
rect 1494 1523 1495 1527
rect 1499 1523 1500 1527
rect 1494 1522 1500 1523
rect 1824 1518 1826 1533
rect 1864 1522 1866 1537
rect 1888 1532 1890 1537
rect 2024 1532 2026 1537
rect 2184 1532 2186 1537
rect 2344 1532 2346 1537
rect 2504 1532 2506 1537
rect 2664 1532 2666 1537
rect 2824 1532 2826 1537
rect 2984 1532 2986 1537
rect 3152 1532 3154 1537
rect 3320 1532 3322 1537
rect 3480 1532 3482 1537
rect 1886 1531 1892 1532
rect 1886 1527 1887 1531
rect 1891 1527 1892 1531
rect 1886 1526 1892 1527
rect 2022 1531 2028 1532
rect 2022 1527 2023 1531
rect 2027 1527 2028 1531
rect 2022 1526 2028 1527
rect 2182 1531 2188 1532
rect 2182 1527 2183 1531
rect 2187 1527 2188 1531
rect 2182 1526 2188 1527
rect 2342 1531 2348 1532
rect 2342 1527 2343 1531
rect 2347 1527 2348 1531
rect 2342 1526 2348 1527
rect 2502 1531 2508 1532
rect 2502 1527 2503 1531
rect 2507 1527 2508 1531
rect 2502 1526 2508 1527
rect 2662 1531 2668 1532
rect 2662 1527 2663 1531
rect 2667 1527 2668 1531
rect 2662 1526 2668 1527
rect 2822 1531 2828 1532
rect 2822 1527 2823 1531
rect 2827 1527 2828 1531
rect 2822 1526 2828 1527
rect 2982 1531 2988 1532
rect 2982 1527 2983 1531
rect 2987 1527 2988 1531
rect 2982 1526 2988 1527
rect 3150 1531 3156 1532
rect 3150 1527 3151 1531
rect 3155 1527 3156 1531
rect 3150 1526 3156 1527
rect 3318 1531 3324 1532
rect 3318 1527 3319 1531
rect 3323 1527 3324 1531
rect 3318 1526 3324 1527
rect 3478 1531 3484 1532
rect 3478 1527 3479 1531
rect 3483 1527 3484 1531
rect 3478 1526 3484 1527
rect 3576 1522 3578 1537
rect 1862 1521 1868 1522
rect 110 1517 116 1518
rect 110 1513 111 1517
rect 115 1513 116 1517
rect 110 1512 116 1513
rect 1822 1517 1828 1518
rect 1822 1513 1823 1517
rect 1827 1513 1828 1517
rect 1862 1517 1863 1521
rect 1867 1517 1868 1521
rect 1862 1516 1868 1517
rect 3574 1521 3580 1522
rect 3574 1517 3575 1521
rect 3579 1517 3580 1521
rect 3574 1516 3580 1517
rect 1822 1512 1828 1513
rect 1862 1504 1868 1505
rect 110 1500 116 1501
rect 110 1496 111 1500
rect 115 1496 116 1500
rect 110 1495 116 1496
rect 1822 1500 1828 1501
rect 1822 1496 1823 1500
rect 1827 1496 1828 1500
rect 1862 1500 1863 1504
rect 1867 1500 1868 1504
rect 1862 1499 1868 1500
rect 3574 1504 3580 1505
rect 3574 1500 3575 1504
rect 3579 1500 3580 1504
rect 3574 1499 3580 1500
rect 1822 1495 1828 1496
rect 112 1463 114 1495
rect 142 1487 148 1488
rect 142 1483 143 1487
rect 147 1483 148 1487
rect 142 1482 148 1483
rect 278 1487 284 1488
rect 278 1483 279 1487
rect 283 1483 284 1487
rect 278 1482 284 1483
rect 430 1487 436 1488
rect 430 1483 431 1487
rect 435 1483 436 1487
rect 430 1482 436 1483
rect 590 1487 596 1488
rect 590 1483 591 1487
rect 595 1483 596 1487
rect 590 1482 596 1483
rect 742 1487 748 1488
rect 742 1483 743 1487
rect 747 1483 748 1487
rect 742 1482 748 1483
rect 894 1487 900 1488
rect 894 1483 895 1487
rect 899 1483 900 1487
rect 894 1482 900 1483
rect 1046 1487 1052 1488
rect 1046 1483 1047 1487
rect 1051 1483 1052 1487
rect 1046 1482 1052 1483
rect 1198 1487 1204 1488
rect 1198 1483 1199 1487
rect 1203 1483 1204 1487
rect 1198 1482 1204 1483
rect 1350 1487 1356 1488
rect 1350 1483 1351 1487
rect 1355 1483 1356 1487
rect 1350 1482 1356 1483
rect 1502 1487 1508 1488
rect 1502 1483 1503 1487
rect 1507 1483 1508 1487
rect 1502 1482 1508 1483
rect 144 1463 146 1482
rect 280 1463 282 1482
rect 432 1463 434 1482
rect 592 1463 594 1482
rect 744 1463 746 1482
rect 896 1463 898 1482
rect 1048 1463 1050 1482
rect 1200 1463 1202 1482
rect 1352 1463 1354 1482
rect 1504 1463 1506 1482
rect 1824 1463 1826 1495
rect 1864 1467 1866 1499
rect 1894 1491 1900 1492
rect 1894 1487 1895 1491
rect 1899 1487 1900 1491
rect 1894 1486 1900 1487
rect 2030 1491 2036 1492
rect 2030 1487 2031 1491
rect 2035 1487 2036 1491
rect 2030 1486 2036 1487
rect 2190 1491 2196 1492
rect 2190 1487 2191 1491
rect 2195 1487 2196 1491
rect 2190 1486 2196 1487
rect 2350 1491 2356 1492
rect 2350 1487 2351 1491
rect 2355 1487 2356 1491
rect 2350 1486 2356 1487
rect 2510 1491 2516 1492
rect 2510 1487 2511 1491
rect 2515 1487 2516 1491
rect 2510 1486 2516 1487
rect 2670 1491 2676 1492
rect 2670 1487 2671 1491
rect 2675 1487 2676 1491
rect 2670 1486 2676 1487
rect 2830 1491 2836 1492
rect 2830 1487 2831 1491
rect 2835 1487 2836 1491
rect 2830 1486 2836 1487
rect 2990 1491 2996 1492
rect 2990 1487 2991 1491
rect 2995 1487 2996 1491
rect 2990 1486 2996 1487
rect 3158 1491 3164 1492
rect 3158 1487 3159 1491
rect 3163 1487 3164 1491
rect 3158 1486 3164 1487
rect 3326 1491 3332 1492
rect 3326 1487 3327 1491
rect 3331 1487 3332 1491
rect 3326 1486 3332 1487
rect 3486 1491 3492 1492
rect 3486 1487 3487 1491
rect 3491 1487 3492 1491
rect 3486 1486 3492 1487
rect 1896 1467 1898 1486
rect 2032 1467 2034 1486
rect 2192 1467 2194 1486
rect 2352 1467 2354 1486
rect 2512 1467 2514 1486
rect 2672 1467 2674 1486
rect 2832 1467 2834 1486
rect 2992 1467 2994 1486
rect 3160 1467 3162 1486
rect 3328 1467 3330 1486
rect 3488 1467 3490 1486
rect 3576 1467 3578 1499
rect 1863 1466 1867 1467
rect 111 1462 115 1463
rect 111 1457 115 1458
rect 143 1462 147 1463
rect 143 1457 147 1458
rect 263 1462 267 1463
rect 263 1457 267 1458
rect 279 1462 283 1463
rect 279 1457 283 1458
rect 399 1462 403 1463
rect 399 1457 403 1458
rect 431 1462 435 1463
rect 431 1457 435 1458
rect 535 1462 539 1463
rect 535 1457 539 1458
rect 591 1462 595 1463
rect 591 1457 595 1458
rect 663 1462 667 1463
rect 663 1457 667 1458
rect 743 1462 747 1463
rect 743 1457 747 1458
rect 791 1462 795 1463
rect 791 1457 795 1458
rect 895 1462 899 1463
rect 895 1457 899 1458
rect 911 1462 915 1463
rect 911 1457 915 1458
rect 1023 1462 1027 1463
rect 1023 1457 1027 1458
rect 1047 1462 1051 1463
rect 1047 1457 1051 1458
rect 1143 1462 1147 1463
rect 1143 1457 1147 1458
rect 1199 1462 1203 1463
rect 1199 1457 1203 1458
rect 1263 1462 1267 1463
rect 1263 1457 1267 1458
rect 1351 1462 1355 1463
rect 1351 1457 1355 1458
rect 1383 1462 1387 1463
rect 1383 1457 1387 1458
rect 1503 1462 1507 1463
rect 1503 1457 1507 1458
rect 1631 1462 1635 1463
rect 1631 1457 1635 1458
rect 1735 1462 1739 1463
rect 1735 1457 1739 1458
rect 1823 1462 1827 1463
rect 1863 1461 1867 1462
rect 1895 1466 1899 1467
rect 1895 1461 1899 1462
rect 2031 1466 2035 1467
rect 2031 1461 2035 1462
rect 2183 1466 2187 1467
rect 2183 1461 2187 1462
rect 2191 1466 2195 1467
rect 2191 1461 2195 1462
rect 2351 1466 2355 1467
rect 2351 1461 2355 1462
rect 2359 1466 2363 1467
rect 2359 1461 2363 1462
rect 2511 1466 2515 1467
rect 2511 1461 2515 1462
rect 2527 1466 2531 1467
rect 2527 1461 2531 1462
rect 2671 1466 2675 1467
rect 2671 1461 2675 1462
rect 2687 1466 2691 1467
rect 2687 1461 2691 1462
rect 2831 1466 2835 1467
rect 2831 1461 2835 1462
rect 2847 1466 2851 1467
rect 2847 1461 2851 1462
rect 2991 1466 2995 1467
rect 2991 1461 2995 1462
rect 3007 1466 3011 1467
rect 3007 1461 3011 1462
rect 3159 1466 3163 1467
rect 3159 1461 3163 1462
rect 3175 1466 3179 1467
rect 3175 1461 3179 1462
rect 3327 1466 3331 1467
rect 3327 1461 3331 1462
rect 3343 1466 3347 1467
rect 3343 1461 3347 1462
rect 3487 1466 3491 1467
rect 3487 1461 3491 1462
rect 3575 1466 3579 1467
rect 3575 1461 3579 1462
rect 1823 1457 1827 1458
rect 112 1433 114 1457
rect 144 1446 146 1457
rect 264 1446 266 1457
rect 400 1446 402 1457
rect 536 1446 538 1457
rect 664 1446 666 1457
rect 792 1446 794 1457
rect 912 1446 914 1457
rect 1024 1446 1026 1457
rect 1144 1446 1146 1457
rect 1264 1446 1266 1457
rect 1384 1446 1386 1457
rect 1504 1446 1506 1457
rect 1632 1446 1634 1457
rect 1736 1446 1738 1457
rect 142 1445 148 1446
rect 142 1441 143 1445
rect 147 1441 148 1445
rect 142 1440 148 1441
rect 262 1445 268 1446
rect 262 1441 263 1445
rect 267 1441 268 1445
rect 262 1440 268 1441
rect 398 1445 404 1446
rect 398 1441 399 1445
rect 403 1441 404 1445
rect 398 1440 404 1441
rect 534 1445 540 1446
rect 534 1441 535 1445
rect 539 1441 540 1445
rect 534 1440 540 1441
rect 662 1445 668 1446
rect 662 1441 663 1445
rect 667 1441 668 1445
rect 662 1440 668 1441
rect 790 1445 796 1446
rect 790 1441 791 1445
rect 795 1441 796 1445
rect 790 1440 796 1441
rect 910 1445 916 1446
rect 910 1441 911 1445
rect 915 1441 916 1445
rect 910 1440 916 1441
rect 1022 1445 1028 1446
rect 1022 1441 1023 1445
rect 1027 1441 1028 1445
rect 1022 1440 1028 1441
rect 1142 1445 1148 1446
rect 1142 1441 1143 1445
rect 1147 1441 1148 1445
rect 1142 1440 1148 1441
rect 1262 1445 1268 1446
rect 1262 1441 1263 1445
rect 1267 1441 1268 1445
rect 1262 1440 1268 1441
rect 1382 1445 1388 1446
rect 1382 1441 1383 1445
rect 1387 1441 1388 1445
rect 1382 1440 1388 1441
rect 1502 1445 1508 1446
rect 1502 1441 1503 1445
rect 1507 1441 1508 1445
rect 1502 1440 1508 1441
rect 1630 1445 1636 1446
rect 1630 1441 1631 1445
rect 1635 1441 1636 1445
rect 1630 1440 1636 1441
rect 1734 1445 1740 1446
rect 1734 1441 1735 1445
rect 1739 1441 1740 1445
rect 1734 1440 1740 1441
rect 1824 1433 1826 1457
rect 1864 1437 1866 1461
rect 2184 1450 2186 1461
rect 2360 1450 2362 1461
rect 2528 1450 2530 1461
rect 2688 1450 2690 1461
rect 2848 1450 2850 1461
rect 3008 1450 3010 1461
rect 3176 1450 3178 1461
rect 3344 1450 3346 1461
rect 3488 1450 3490 1461
rect 2182 1449 2188 1450
rect 2182 1445 2183 1449
rect 2187 1445 2188 1449
rect 2182 1444 2188 1445
rect 2358 1449 2364 1450
rect 2358 1445 2359 1449
rect 2363 1445 2364 1449
rect 2358 1444 2364 1445
rect 2526 1449 2532 1450
rect 2526 1445 2527 1449
rect 2531 1445 2532 1449
rect 2526 1444 2532 1445
rect 2686 1449 2692 1450
rect 2686 1445 2687 1449
rect 2691 1445 2692 1449
rect 2686 1444 2692 1445
rect 2846 1449 2852 1450
rect 2846 1445 2847 1449
rect 2851 1445 2852 1449
rect 2846 1444 2852 1445
rect 3006 1449 3012 1450
rect 3006 1445 3007 1449
rect 3011 1445 3012 1449
rect 3006 1444 3012 1445
rect 3174 1449 3180 1450
rect 3174 1445 3175 1449
rect 3179 1445 3180 1449
rect 3174 1444 3180 1445
rect 3342 1449 3348 1450
rect 3342 1445 3343 1449
rect 3347 1445 3348 1449
rect 3342 1444 3348 1445
rect 3486 1449 3492 1450
rect 3486 1445 3487 1449
rect 3491 1445 3492 1449
rect 3486 1444 3492 1445
rect 3576 1437 3578 1461
rect 1862 1436 1868 1437
rect 110 1432 116 1433
rect 110 1428 111 1432
rect 115 1428 116 1432
rect 110 1427 116 1428
rect 1822 1432 1828 1433
rect 1822 1428 1823 1432
rect 1827 1428 1828 1432
rect 1862 1432 1863 1436
rect 1867 1432 1868 1436
rect 1862 1431 1868 1432
rect 3574 1436 3580 1437
rect 3574 1432 3575 1436
rect 3579 1432 3580 1436
rect 3574 1431 3580 1432
rect 1822 1427 1828 1428
rect 1862 1419 1868 1420
rect 110 1415 116 1416
rect 110 1411 111 1415
rect 115 1411 116 1415
rect 110 1410 116 1411
rect 1822 1415 1828 1416
rect 1822 1411 1823 1415
rect 1827 1411 1828 1415
rect 1862 1415 1863 1419
rect 1867 1415 1868 1419
rect 1862 1414 1868 1415
rect 3574 1419 3580 1420
rect 3574 1415 3575 1419
rect 3579 1415 3580 1419
rect 3574 1414 3580 1415
rect 1822 1410 1828 1411
rect 112 1395 114 1410
rect 134 1405 140 1406
rect 134 1401 135 1405
rect 139 1401 140 1405
rect 134 1400 140 1401
rect 254 1405 260 1406
rect 254 1401 255 1405
rect 259 1401 260 1405
rect 254 1400 260 1401
rect 390 1405 396 1406
rect 390 1401 391 1405
rect 395 1401 396 1405
rect 390 1400 396 1401
rect 526 1405 532 1406
rect 526 1401 527 1405
rect 531 1401 532 1405
rect 526 1400 532 1401
rect 654 1405 660 1406
rect 654 1401 655 1405
rect 659 1401 660 1405
rect 654 1400 660 1401
rect 782 1405 788 1406
rect 782 1401 783 1405
rect 787 1401 788 1405
rect 782 1400 788 1401
rect 902 1405 908 1406
rect 902 1401 903 1405
rect 907 1401 908 1405
rect 902 1400 908 1401
rect 1014 1405 1020 1406
rect 1014 1401 1015 1405
rect 1019 1401 1020 1405
rect 1014 1400 1020 1401
rect 1134 1405 1140 1406
rect 1134 1401 1135 1405
rect 1139 1401 1140 1405
rect 1134 1400 1140 1401
rect 1254 1405 1260 1406
rect 1254 1401 1255 1405
rect 1259 1401 1260 1405
rect 1254 1400 1260 1401
rect 1374 1405 1380 1406
rect 1374 1401 1375 1405
rect 1379 1401 1380 1405
rect 1374 1400 1380 1401
rect 1494 1405 1500 1406
rect 1494 1401 1495 1405
rect 1499 1401 1500 1405
rect 1494 1400 1500 1401
rect 1622 1405 1628 1406
rect 1622 1401 1623 1405
rect 1627 1401 1628 1405
rect 1622 1400 1628 1401
rect 1726 1405 1732 1406
rect 1726 1401 1727 1405
rect 1731 1401 1732 1405
rect 1726 1400 1732 1401
rect 136 1395 138 1400
rect 256 1395 258 1400
rect 392 1395 394 1400
rect 528 1395 530 1400
rect 656 1395 658 1400
rect 784 1395 786 1400
rect 904 1395 906 1400
rect 1016 1395 1018 1400
rect 1136 1395 1138 1400
rect 1256 1395 1258 1400
rect 1376 1395 1378 1400
rect 1496 1395 1498 1400
rect 1624 1395 1626 1400
rect 1728 1395 1730 1400
rect 1824 1395 1826 1410
rect 111 1394 115 1395
rect 111 1389 115 1390
rect 135 1394 139 1395
rect 135 1389 139 1390
rect 255 1394 259 1395
rect 255 1389 259 1390
rect 327 1394 331 1395
rect 327 1389 331 1390
rect 391 1394 395 1395
rect 391 1389 395 1390
rect 527 1394 531 1395
rect 527 1389 531 1390
rect 551 1394 555 1395
rect 551 1389 555 1390
rect 655 1394 659 1395
rect 655 1389 659 1390
rect 783 1394 787 1395
rect 783 1389 787 1390
rect 903 1394 907 1395
rect 903 1389 907 1390
rect 1015 1394 1019 1395
rect 1015 1389 1019 1390
rect 1023 1394 1027 1395
rect 1023 1389 1027 1390
rect 1135 1394 1139 1395
rect 1135 1389 1139 1390
rect 1255 1394 1259 1395
rect 1255 1389 1259 1390
rect 1263 1394 1267 1395
rect 1263 1389 1267 1390
rect 1375 1394 1379 1395
rect 1375 1389 1379 1390
rect 1495 1394 1499 1395
rect 1495 1389 1499 1390
rect 1503 1394 1507 1395
rect 1503 1389 1507 1390
rect 1623 1394 1627 1395
rect 1623 1389 1627 1390
rect 1727 1394 1731 1395
rect 1727 1389 1731 1390
rect 1823 1394 1827 1395
rect 1864 1391 1866 1414
rect 2174 1409 2180 1410
rect 2174 1405 2175 1409
rect 2179 1405 2180 1409
rect 2174 1404 2180 1405
rect 2350 1409 2356 1410
rect 2350 1405 2351 1409
rect 2355 1405 2356 1409
rect 2350 1404 2356 1405
rect 2518 1409 2524 1410
rect 2518 1405 2519 1409
rect 2523 1405 2524 1409
rect 2518 1404 2524 1405
rect 2678 1409 2684 1410
rect 2678 1405 2679 1409
rect 2683 1405 2684 1409
rect 2678 1404 2684 1405
rect 2838 1409 2844 1410
rect 2838 1405 2839 1409
rect 2843 1405 2844 1409
rect 2838 1404 2844 1405
rect 2998 1409 3004 1410
rect 2998 1405 2999 1409
rect 3003 1405 3004 1409
rect 2998 1404 3004 1405
rect 3166 1409 3172 1410
rect 3166 1405 3167 1409
rect 3171 1405 3172 1409
rect 3166 1404 3172 1405
rect 3334 1409 3340 1410
rect 3334 1405 3335 1409
rect 3339 1405 3340 1409
rect 3334 1404 3340 1405
rect 3478 1409 3484 1410
rect 3478 1405 3479 1409
rect 3483 1405 3484 1409
rect 3478 1404 3484 1405
rect 2176 1391 2178 1404
rect 2352 1391 2354 1404
rect 2520 1391 2522 1404
rect 2680 1391 2682 1404
rect 2840 1391 2842 1404
rect 3000 1391 3002 1404
rect 3168 1391 3170 1404
rect 3336 1391 3338 1404
rect 3480 1391 3482 1404
rect 3576 1391 3578 1414
rect 1823 1389 1827 1390
rect 1863 1390 1867 1391
rect 112 1374 114 1389
rect 136 1384 138 1389
rect 328 1384 330 1389
rect 552 1384 554 1389
rect 784 1384 786 1389
rect 1024 1384 1026 1389
rect 1264 1384 1266 1389
rect 1504 1384 1506 1389
rect 1728 1384 1730 1389
rect 134 1383 140 1384
rect 134 1379 135 1383
rect 139 1379 140 1383
rect 134 1378 140 1379
rect 326 1383 332 1384
rect 326 1379 327 1383
rect 331 1379 332 1383
rect 326 1378 332 1379
rect 550 1383 556 1384
rect 550 1379 551 1383
rect 555 1379 556 1383
rect 550 1378 556 1379
rect 782 1383 788 1384
rect 782 1379 783 1383
rect 787 1379 788 1383
rect 782 1378 788 1379
rect 1022 1383 1028 1384
rect 1022 1379 1023 1383
rect 1027 1379 1028 1383
rect 1022 1378 1028 1379
rect 1262 1383 1268 1384
rect 1262 1379 1263 1383
rect 1267 1379 1268 1383
rect 1262 1378 1268 1379
rect 1502 1383 1508 1384
rect 1502 1379 1503 1383
rect 1507 1379 1508 1383
rect 1502 1378 1508 1379
rect 1726 1383 1732 1384
rect 1726 1379 1727 1383
rect 1731 1379 1732 1383
rect 1726 1378 1732 1379
rect 1824 1374 1826 1389
rect 1863 1385 1867 1386
rect 2079 1390 2083 1391
rect 2079 1385 2083 1386
rect 2175 1390 2179 1391
rect 2175 1385 2179 1386
rect 2263 1390 2267 1391
rect 2263 1385 2267 1386
rect 2351 1390 2355 1391
rect 2351 1385 2355 1386
rect 2439 1390 2443 1391
rect 2439 1385 2443 1386
rect 2519 1390 2523 1391
rect 2519 1385 2523 1386
rect 2615 1390 2619 1391
rect 2615 1385 2619 1386
rect 2679 1390 2683 1391
rect 2679 1385 2683 1386
rect 2783 1390 2787 1391
rect 2783 1385 2787 1386
rect 2839 1390 2843 1391
rect 2839 1385 2843 1386
rect 2935 1390 2939 1391
rect 2935 1385 2939 1386
rect 2999 1390 3003 1391
rect 2999 1385 3003 1386
rect 3079 1390 3083 1391
rect 3079 1385 3083 1386
rect 3167 1390 3171 1391
rect 3167 1385 3171 1386
rect 3223 1390 3227 1391
rect 3223 1385 3227 1386
rect 3335 1390 3339 1391
rect 3335 1385 3339 1386
rect 3359 1390 3363 1391
rect 3359 1385 3363 1386
rect 3479 1390 3483 1391
rect 3479 1385 3483 1386
rect 3575 1390 3579 1391
rect 3575 1385 3579 1386
rect 110 1373 116 1374
rect 110 1369 111 1373
rect 115 1369 116 1373
rect 110 1368 116 1369
rect 1822 1373 1828 1374
rect 1822 1369 1823 1373
rect 1827 1369 1828 1373
rect 1864 1370 1866 1385
rect 2080 1380 2082 1385
rect 2264 1380 2266 1385
rect 2440 1380 2442 1385
rect 2616 1380 2618 1385
rect 2784 1380 2786 1385
rect 2936 1380 2938 1385
rect 3080 1380 3082 1385
rect 3224 1380 3226 1385
rect 3360 1380 3362 1385
rect 3480 1380 3482 1385
rect 2078 1379 2084 1380
rect 2078 1375 2079 1379
rect 2083 1375 2084 1379
rect 2078 1374 2084 1375
rect 2262 1379 2268 1380
rect 2262 1375 2263 1379
rect 2267 1375 2268 1379
rect 2262 1374 2268 1375
rect 2438 1379 2444 1380
rect 2438 1375 2439 1379
rect 2443 1375 2444 1379
rect 2438 1374 2444 1375
rect 2614 1379 2620 1380
rect 2614 1375 2615 1379
rect 2619 1375 2620 1379
rect 2614 1374 2620 1375
rect 2782 1379 2788 1380
rect 2782 1375 2783 1379
rect 2787 1375 2788 1379
rect 2782 1374 2788 1375
rect 2934 1379 2940 1380
rect 2934 1375 2935 1379
rect 2939 1375 2940 1379
rect 2934 1374 2940 1375
rect 3078 1379 3084 1380
rect 3078 1375 3079 1379
rect 3083 1375 3084 1379
rect 3078 1374 3084 1375
rect 3222 1379 3228 1380
rect 3222 1375 3223 1379
rect 3227 1375 3228 1379
rect 3222 1374 3228 1375
rect 3358 1379 3364 1380
rect 3358 1375 3359 1379
rect 3363 1375 3364 1379
rect 3358 1374 3364 1375
rect 3478 1379 3484 1380
rect 3478 1375 3479 1379
rect 3483 1375 3484 1379
rect 3478 1374 3484 1375
rect 3576 1370 3578 1385
rect 1822 1368 1828 1369
rect 1862 1369 1868 1370
rect 1862 1365 1863 1369
rect 1867 1365 1868 1369
rect 1862 1364 1868 1365
rect 3574 1369 3580 1370
rect 3574 1365 3575 1369
rect 3579 1365 3580 1369
rect 3574 1364 3580 1365
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 110 1351 116 1352
rect 1822 1356 1828 1357
rect 1822 1352 1823 1356
rect 1827 1352 1828 1356
rect 1822 1351 1828 1352
rect 1862 1352 1868 1353
rect 112 1319 114 1351
rect 142 1343 148 1344
rect 142 1339 143 1343
rect 147 1339 148 1343
rect 142 1338 148 1339
rect 334 1343 340 1344
rect 334 1339 335 1343
rect 339 1339 340 1343
rect 334 1338 340 1339
rect 558 1343 564 1344
rect 558 1339 559 1343
rect 563 1339 564 1343
rect 558 1338 564 1339
rect 790 1343 796 1344
rect 790 1339 791 1343
rect 795 1339 796 1343
rect 790 1338 796 1339
rect 1030 1343 1036 1344
rect 1030 1339 1031 1343
rect 1035 1339 1036 1343
rect 1030 1338 1036 1339
rect 1270 1343 1276 1344
rect 1270 1339 1271 1343
rect 1275 1339 1276 1343
rect 1270 1338 1276 1339
rect 1510 1343 1516 1344
rect 1510 1339 1511 1343
rect 1515 1339 1516 1343
rect 1510 1338 1516 1339
rect 1734 1343 1740 1344
rect 1734 1339 1735 1343
rect 1739 1339 1740 1343
rect 1734 1338 1740 1339
rect 144 1319 146 1338
rect 336 1319 338 1338
rect 560 1319 562 1338
rect 792 1319 794 1338
rect 1032 1319 1034 1338
rect 1272 1319 1274 1338
rect 1512 1319 1514 1338
rect 1736 1319 1738 1338
rect 1824 1319 1826 1351
rect 1862 1348 1863 1352
rect 1867 1348 1868 1352
rect 1862 1347 1868 1348
rect 3574 1352 3580 1353
rect 3574 1348 3575 1352
rect 3579 1348 3580 1352
rect 3574 1347 3580 1348
rect 1864 1323 1866 1347
rect 2086 1339 2092 1340
rect 2086 1335 2087 1339
rect 2091 1335 2092 1339
rect 2086 1334 2092 1335
rect 2270 1339 2276 1340
rect 2270 1335 2271 1339
rect 2275 1335 2276 1339
rect 2270 1334 2276 1335
rect 2446 1339 2452 1340
rect 2446 1335 2447 1339
rect 2451 1335 2452 1339
rect 2446 1334 2452 1335
rect 2622 1339 2628 1340
rect 2622 1335 2623 1339
rect 2627 1335 2628 1339
rect 2622 1334 2628 1335
rect 2790 1339 2796 1340
rect 2790 1335 2791 1339
rect 2795 1335 2796 1339
rect 2790 1334 2796 1335
rect 2942 1339 2948 1340
rect 2942 1335 2943 1339
rect 2947 1335 2948 1339
rect 2942 1334 2948 1335
rect 3086 1339 3092 1340
rect 3086 1335 3087 1339
rect 3091 1335 3092 1339
rect 3086 1334 3092 1335
rect 3230 1339 3236 1340
rect 3230 1335 3231 1339
rect 3235 1335 3236 1339
rect 3230 1334 3236 1335
rect 3366 1339 3372 1340
rect 3366 1335 3367 1339
rect 3371 1335 3372 1339
rect 3366 1334 3372 1335
rect 3486 1339 3492 1340
rect 3486 1335 3487 1339
rect 3491 1335 3492 1339
rect 3486 1334 3492 1335
rect 2088 1323 2090 1334
rect 2272 1323 2274 1334
rect 2448 1323 2450 1334
rect 2624 1323 2626 1334
rect 2792 1323 2794 1334
rect 2944 1323 2946 1334
rect 3088 1323 3090 1334
rect 3232 1323 3234 1334
rect 3368 1323 3370 1334
rect 3488 1323 3490 1334
rect 3576 1323 3578 1347
rect 1863 1322 1867 1323
rect 111 1318 115 1319
rect 111 1313 115 1314
rect 143 1318 147 1319
rect 143 1313 147 1314
rect 327 1318 331 1319
rect 327 1313 331 1314
rect 335 1318 339 1319
rect 335 1313 339 1314
rect 527 1318 531 1319
rect 527 1313 531 1314
rect 559 1318 563 1319
rect 559 1313 563 1314
rect 719 1318 723 1319
rect 719 1313 723 1314
rect 791 1318 795 1319
rect 791 1313 795 1314
rect 903 1318 907 1319
rect 903 1313 907 1314
rect 1031 1318 1035 1319
rect 1031 1313 1035 1314
rect 1071 1318 1075 1319
rect 1071 1313 1075 1314
rect 1231 1318 1235 1319
rect 1231 1313 1235 1314
rect 1271 1318 1275 1319
rect 1271 1313 1275 1314
rect 1383 1318 1387 1319
rect 1383 1313 1387 1314
rect 1511 1318 1515 1319
rect 1511 1313 1515 1314
rect 1535 1318 1539 1319
rect 1535 1313 1539 1314
rect 1687 1318 1691 1319
rect 1687 1313 1691 1314
rect 1735 1318 1739 1319
rect 1735 1313 1739 1314
rect 1823 1318 1827 1319
rect 1863 1317 1867 1318
rect 2087 1322 2091 1323
rect 2087 1317 2091 1318
rect 2271 1322 2275 1323
rect 2271 1317 2275 1318
rect 2311 1322 2315 1323
rect 2311 1317 2315 1318
rect 2447 1322 2451 1323
rect 2447 1317 2451 1318
rect 2519 1322 2523 1323
rect 2519 1317 2523 1318
rect 2623 1322 2627 1323
rect 2623 1317 2627 1318
rect 2711 1322 2715 1323
rect 2711 1317 2715 1318
rect 2791 1322 2795 1323
rect 2791 1317 2795 1318
rect 2887 1322 2891 1323
rect 2887 1317 2891 1318
rect 2943 1322 2947 1323
rect 2943 1317 2947 1318
rect 3047 1322 3051 1323
rect 3047 1317 3051 1318
rect 3087 1322 3091 1323
rect 3087 1317 3091 1318
rect 3199 1322 3203 1323
rect 3199 1317 3203 1318
rect 3231 1322 3235 1323
rect 3231 1317 3235 1318
rect 3351 1322 3355 1323
rect 3351 1317 3355 1318
rect 3367 1322 3371 1323
rect 3367 1317 3371 1318
rect 3487 1322 3491 1323
rect 3487 1317 3491 1318
rect 3575 1322 3579 1323
rect 3575 1317 3579 1318
rect 1823 1313 1827 1314
rect 112 1289 114 1313
rect 144 1302 146 1313
rect 328 1302 330 1313
rect 528 1302 530 1313
rect 720 1302 722 1313
rect 904 1302 906 1313
rect 1072 1302 1074 1313
rect 1232 1302 1234 1313
rect 1384 1302 1386 1313
rect 1536 1302 1538 1313
rect 1688 1302 1690 1313
rect 142 1301 148 1302
rect 142 1297 143 1301
rect 147 1297 148 1301
rect 142 1296 148 1297
rect 326 1301 332 1302
rect 326 1297 327 1301
rect 331 1297 332 1301
rect 326 1296 332 1297
rect 526 1301 532 1302
rect 526 1297 527 1301
rect 531 1297 532 1301
rect 526 1296 532 1297
rect 718 1301 724 1302
rect 718 1297 719 1301
rect 723 1297 724 1301
rect 718 1296 724 1297
rect 902 1301 908 1302
rect 902 1297 903 1301
rect 907 1297 908 1301
rect 902 1296 908 1297
rect 1070 1301 1076 1302
rect 1070 1297 1071 1301
rect 1075 1297 1076 1301
rect 1070 1296 1076 1297
rect 1230 1301 1236 1302
rect 1230 1297 1231 1301
rect 1235 1297 1236 1301
rect 1230 1296 1236 1297
rect 1382 1301 1388 1302
rect 1382 1297 1383 1301
rect 1387 1297 1388 1301
rect 1382 1296 1388 1297
rect 1534 1301 1540 1302
rect 1534 1297 1535 1301
rect 1539 1297 1540 1301
rect 1534 1296 1540 1297
rect 1686 1301 1692 1302
rect 1686 1297 1687 1301
rect 1691 1297 1692 1301
rect 1686 1296 1692 1297
rect 1824 1289 1826 1313
rect 1864 1293 1866 1317
rect 2088 1306 2090 1317
rect 2312 1306 2314 1317
rect 2520 1306 2522 1317
rect 2712 1306 2714 1317
rect 2888 1306 2890 1317
rect 3048 1306 3050 1317
rect 3200 1306 3202 1317
rect 3352 1306 3354 1317
rect 3488 1306 3490 1317
rect 2086 1305 2092 1306
rect 2086 1301 2087 1305
rect 2091 1301 2092 1305
rect 2086 1300 2092 1301
rect 2310 1305 2316 1306
rect 2310 1301 2311 1305
rect 2315 1301 2316 1305
rect 2310 1300 2316 1301
rect 2518 1305 2524 1306
rect 2518 1301 2519 1305
rect 2523 1301 2524 1305
rect 2518 1300 2524 1301
rect 2710 1305 2716 1306
rect 2710 1301 2711 1305
rect 2715 1301 2716 1305
rect 2710 1300 2716 1301
rect 2886 1305 2892 1306
rect 2886 1301 2887 1305
rect 2891 1301 2892 1305
rect 2886 1300 2892 1301
rect 3046 1305 3052 1306
rect 3046 1301 3047 1305
rect 3051 1301 3052 1305
rect 3046 1300 3052 1301
rect 3198 1305 3204 1306
rect 3198 1301 3199 1305
rect 3203 1301 3204 1305
rect 3198 1300 3204 1301
rect 3350 1305 3356 1306
rect 3350 1301 3351 1305
rect 3355 1301 3356 1305
rect 3350 1300 3356 1301
rect 3486 1305 3492 1306
rect 3486 1301 3487 1305
rect 3491 1301 3492 1305
rect 3486 1300 3492 1301
rect 3576 1293 3578 1317
rect 1862 1292 1868 1293
rect 110 1288 116 1289
rect 110 1284 111 1288
rect 115 1284 116 1288
rect 110 1283 116 1284
rect 1822 1288 1828 1289
rect 1822 1284 1823 1288
rect 1827 1284 1828 1288
rect 1862 1288 1863 1292
rect 1867 1288 1868 1292
rect 1862 1287 1868 1288
rect 3574 1292 3580 1293
rect 3574 1288 3575 1292
rect 3579 1288 3580 1292
rect 3574 1287 3580 1288
rect 1822 1283 1828 1284
rect 1862 1275 1868 1276
rect 110 1271 116 1272
rect 110 1267 111 1271
rect 115 1267 116 1271
rect 110 1266 116 1267
rect 1822 1271 1828 1272
rect 1822 1267 1823 1271
rect 1827 1267 1828 1271
rect 1862 1271 1863 1275
rect 1867 1271 1868 1275
rect 1862 1270 1868 1271
rect 3574 1275 3580 1276
rect 3574 1271 3575 1275
rect 3579 1271 3580 1275
rect 3574 1270 3580 1271
rect 1822 1266 1828 1267
rect 112 1247 114 1266
rect 134 1261 140 1262
rect 134 1257 135 1261
rect 139 1257 140 1261
rect 134 1256 140 1257
rect 318 1261 324 1262
rect 318 1257 319 1261
rect 323 1257 324 1261
rect 318 1256 324 1257
rect 518 1261 524 1262
rect 518 1257 519 1261
rect 523 1257 524 1261
rect 518 1256 524 1257
rect 710 1261 716 1262
rect 710 1257 711 1261
rect 715 1257 716 1261
rect 710 1256 716 1257
rect 894 1261 900 1262
rect 894 1257 895 1261
rect 899 1257 900 1261
rect 894 1256 900 1257
rect 1062 1261 1068 1262
rect 1062 1257 1063 1261
rect 1067 1257 1068 1261
rect 1062 1256 1068 1257
rect 1222 1261 1228 1262
rect 1222 1257 1223 1261
rect 1227 1257 1228 1261
rect 1222 1256 1228 1257
rect 1374 1261 1380 1262
rect 1374 1257 1375 1261
rect 1379 1257 1380 1261
rect 1374 1256 1380 1257
rect 1526 1261 1532 1262
rect 1526 1257 1527 1261
rect 1531 1257 1532 1261
rect 1526 1256 1532 1257
rect 1678 1261 1684 1262
rect 1678 1257 1679 1261
rect 1683 1257 1684 1261
rect 1678 1256 1684 1257
rect 136 1247 138 1256
rect 320 1247 322 1256
rect 520 1247 522 1256
rect 712 1247 714 1256
rect 896 1247 898 1256
rect 1064 1247 1066 1256
rect 1224 1247 1226 1256
rect 1376 1247 1378 1256
rect 1528 1247 1530 1256
rect 1680 1247 1682 1256
rect 1824 1247 1826 1266
rect 1864 1251 1866 1270
rect 2078 1265 2084 1266
rect 2078 1261 2079 1265
rect 2083 1261 2084 1265
rect 2078 1260 2084 1261
rect 2302 1265 2308 1266
rect 2302 1261 2303 1265
rect 2307 1261 2308 1265
rect 2302 1260 2308 1261
rect 2510 1265 2516 1266
rect 2510 1261 2511 1265
rect 2515 1261 2516 1265
rect 2510 1260 2516 1261
rect 2702 1265 2708 1266
rect 2702 1261 2703 1265
rect 2707 1261 2708 1265
rect 2702 1260 2708 1261
rect 2878 1265 2884 1266
rect 2878 1261 2879 1265
rect 2883 1261 2884 1265
rect 2878 1260 2884 1261
rect 3038 1265 3044 1266
rect 3038 1261 3039 1265
rect 3043 1261 3044 1265
rect 3038 1260 3044 1261
rect 3190 1265 3196 1266
rect 3190 1261 3191 1265
rect 3195 1261 3196 1265
rect 3190 1260 3196 1261
rect 3342 1265 3348 1266
rect 3342 1261 3343 1265
rect 3347 1261 3348 1265
rect 3342 1260 3348 1261
rect 3478 1265 3484 1266
rect 3478 1261 3479 1265
rect 3483 1261 3484 1265
rect 3478 1260 3484 1261
rect 2080 1251 2082 1260
rect 2304 1251 2306 1260
rect 2512 1251 2514 1260
rect 2704 1251 2706 1260
rect 2880 1251 2882 1260
rect 3040 1251 3042 1260
rect 3192 1251 3194 1260
rect 3344 1251 3346 1260
rect 3480 1251 3482 1260
rect 3576 1251 3578 1270
rect 1863 1250 1867 1251
rect 111 1246 115 1247
rect 111 1241 115 1242
rect 135 1246 139 1247
rect 135 1241 139 1242
rect 295 1246 299 1247
rect 295 1241 299 1242
rect 319 1246 323 1247
rect 319 1241 323 1242
rect 479 1246 483 1247
rect 479 1241 483 1242
rect 519 1246 523 1247
rect 519 1241 523 1242
rect 655 1246 659 1247
rect 655 1241 659 1242
rect 711 1246 715 1247
rect 711 1241 715 1242
rect 815 1246 819 1247
rect 815 1241 819 1242
rect 895 1246 899 1247
rect 895 1241 899 1242
rect 967 1246 971 1247
rect 967 1241 971 1242
rect 1063 1246 1067 1247
rect 1063 1241 1067 1242
rect 1111 1246 1115 1247
rect 1111 1241 1115 1242
rect 1223 1246 1227 1247
rect 1223 1241 1227 1242
rect 1247 1246 1251 1247
rect 1247 1241 1251 1242
rect 1375 1246 1379 1247
rect 1375 1241 1379 1242
rect 1383 1246 1387 1247
rect 1383 1241 1387 1242
rect 1527 1246 1531 1247
rect 1527 1241 1531 1242
rect 1679 1246 1683 1247
rect 1679 1241 1683 1242
rect 1823 1246 1827 1247
rect 1863 1245 1867 1246
rect 1903 1250 1907 1251
rect 1903 1245 1907 1246
rect 1991 1250 1995 1251
rect 1991 1245 1995 1246
rect 2079 1250 2083 1251
rect 2079 1245 2083 1246
rect 2095 1250 2099 1251
rect 2095 1245 2099 1246
rect 2215 1250 2219 1251
rect 2215 1245 2219 1246
rect 2303 1250 2307 1251
rect 2303 1245 2307 1246
rect 2351 1250 2355 1251
rect 2351 1245 2355 1246
rect 2487 1250 2491 1251
rect 2487 1245 2491 1246
rect 2511 1250 2515 1251
rect 2511 1245 2515 1246
rect 2631 1250 2635 1251
rect 2631 1245 2635 1246
rect 2703 1250 2707 1251
rect 2703 1245 2707 1246
rect 2775 1250 2779 1251
rect 2775 1245 2779 1246
rect 2879 1250 2883 1251
rect 2879 1245 2883 1246
rect 2919 1250 2923 1251
rect 2919 1245 2923 1246
rect 3039 1250 3043 1251
rect 3039 1245 3043 1246
rect 3063 1250 3067 1251
rect 3063 1245 3067 1246
rect 3191 1250 3195 1251
rect 3191 1245 3195 1246
rect 3207 1250 3211 1251
rect 3207 1245 3211 1246
rect 3343 1250 3347 1251
rect 3343 1245 3347 1246
rect 3351 1250 3355 1251
rect 3351 1245 3355 1246
rect 3479 1250 3483 1251
rect 3479 1245 3483 1246
rect 3575 1250 3579 1251
rect 3575 1245 3579 1246
rect 1823 1241 1827 1242
rect 112 1226 114 1241
rect 136 1236 138 1241
rect 296 1236 298 1241
rect 480 1236 482 1241
rect 656 1236 658 1241
rect 816 1236 818 1241
rect 968 1236 970 1241
rect 1112 1236 1114 1241
rect 1248 1236 1250 1241
rect 1384 1236 1386 1241
rect 1528 1236 1530 1241
rect 134 1235 140 1236
rect 134 1231 135 1235
rect 139 1231 140 1235
rect 134 1230 140 1231
rect 294 1235 300 1236
rect 294 1231 295 1235
rect 299 1231 300 1235
rect 294 1230 300 1231
rect 478 1235 484 1236
rect 478 1231 479 1235
rect 483 1231 484 1235
rect 478 1230 484 1231
rect 654 1235 660 1236
rect 654 1231 655 1235
rect 659 1231 660 1235
rect 654 1230 660 1231
rect 814 1235 820 1236
rect 814 1231 815 1235
rect 819 1231 820 1235
rect 814 1230 820 1231
rect 966 1235 972 1236
rect 966 1231 967 1235
rect 971 1231 972 1235
rect 966 1230 972 1231
rect 1110 1235 1116 1236
rect 1110 1231 1111 1235
rect 1115 1231 1116 1235
rect 1110 1230 1116 1231
rect 1246 1235 1252 1236
rect 1246 1231 1247 1235
rect 1251 1231 1252 1235
rect 1246 1230 1252 1231
rect 1382 1235 1388 1236
rect 1382 1231 1383 1235
rect 1387 1231 1388 1235
rect 1382 1230 1388 1231
rect 1526 1235 1532 1236
rect 1526 1231 1527 1235
rect 1531 1231 1532 1235
rect 1526 1230 1532 1231
rect 1824 1226 1826 1241
rect 1864 1230 1866 1245
rect 1904 1240 1906 1245
rect 1992 1240 1994 1245
rect 2096 1240 2098 1245
rect 2216 1240 2218 1245
rect 2352 1240 2354 1245
rect 2488 1240 2490 1245
rect 2632 1240 2634 1245
rect 2776 1240 2778 1245
rect 2920 1240 2922 1245
rect 3064 1240 3066 1245
rect 3208 1240 3210 1245
rect 3352 1240 3354 1245
rect 3480 1240 3482 1245
rect 1902 1239 1908 1240
rect 1902 1235 1903 1239
rect 1907 1235 1908 1239
rect 1902 1234 1908 1235
rect 1990 1239 1996 1240
rect 1990 1235 1991 1239
rect 1995 1235 1996 1239
rect 1990 1234 1996 1235
rect 2094 1239 2100 1240
rect 2094 1235 2095 1239
rect 2099 1235 2100 1239
rect 2094 1234 2100 1235
rect 2214 1239 2220 1240
rect 2214 1235 2215 1239
rect 2219 1235 2220 1239
rect 2214 1234 2220 1235
rect 2350 1239 2356 1240
rect 2350 1235 2351 1239
rect 2355 1235 2356 1239
rect 2350 1234 2356 1235
rect 2486 1239 2492 1240
rect 2486 1235 2487 1239
rect 2491 1235 2492 1239
rect 2486 1234 2492 1235
rect 2630 1239 2636 1240
rect 2630 1235 2631 1239
rect 2635 1235 2636 1239
rect 2630 1234 2636 1235
rect 2774 1239 2780 1240
rect 2774 1235 2775 1239
rect 2779 1235 2780 1239
rect 2774 1234 2780 1235
rect 2918 1239 2924 1240
rect 2918 1235 2919 1239
rect 2923 1235 2924 1239
rect 2918 1234 2924 1235
rect 3062 1239 3068 1240
rect 3062 1235 3063 1239
rect 3067 1235 3068 1239
rect 3062 1234 3068 1235
rect 3206 1239 3212 1240
rect 3206 1235 3207 1239
rect 3211 1235 3212 1239
rect 3206 1234 3212 1235
rect 3350 1239 3356 1240
rect 3350 1235 3351 1239
rect 3355 1235 3356 1239
rect 3350 1234 3356 1235
rect 3478 1239 3484 1240
rect 3478 1235 3479 1239
rect 3483 1235 3484 1239
rect 3478 1234 3484 1235
rect 3576 1230 3578 1245
rect 1862 1229 1868 1230
rect 110 1225 116 1226
rect 110 1221 111 1225
rect 115 1221 116 1225
rect 110 1220 116 1221
rect 1822 1225 1828 1226
rect 1822 1221 1823 1225
rect 1827 1221 1828 1225
rect 1862 1225 1863 1229
rect 1867 1225 1868 1229
rect 1862 1224 1868 1225
rect 3574 1229 3580 1230
rect 3574 1225 3575 1229
rect 3579 1225 3580 1229
rect 3574 1224 3580 1225
rect 1822 1220 1828 1221
rect 1862 1212 1868 1213
rect 110 1208 116 1209
rect 110 1204 111 1208
rect 115 1204 116 1208
rect 110 1203 116 1204
rect 1822 1208 1828 1209
rect 1822 1204 1823 1208
rect 1827 1204 1828 1208
rect 1862 1208 1863 1212
rect 1867 1208 1868 1212
rect 1862 1207 1868 1208
rect 3574 1212 3580 1213
rect 3574 1208 3575 1212
rect 3579 1208 3580 1212
rect 3574 1207 3580 1208
rect 1822 1203 1828 1204
rect 112 1175 114 1203
rect 142 1195 148 1196
rect 142 1191 143 1195
rect 147 1191 148 1195
rect 142 1190 148 1191
rect 302 1195 308 1196
rect 302 1191 303 1195
rect 307 1191 308 1195
rect 302 1190 308 1191
rect 486 1195 492 1196
rect 486 1191 487 1195
rect 491 1191 492 1195
rect 486 1190 492 1191
rect 662 1195 668 1196
rect 662 1191 663 1195
rect 667 1191 668 1195
rect 662 1190 668 1191
rect 822 1195 828 1196
rect 822 1191 823 1195
rect 827 1191 828 1195
rect 822 1190 828 1191
rect 974 1195 980 1196
rect 974 1191 975 1195
rect 979 1191 980 1195
rect 974 1190 980 1191
rect 1118 1195 1124 1196
rect 1118 1191 1119 1195
rect 1123 1191 1124 1195
rect 1118 1190 1124 1191
rect 1254 1195 1260 1196
rect 1254 1191 1255 1195
rect 1259 1191 1260 1195
rect 1254 1190 1260 1191
rect 1390 1195 1396 1196
rect 1390 1191 1391 1195
rect 1395 1191 1396 1195
rect 1390 1190 1396 1191
rect 1534 1195 1540 1196
rect 1534 1191 1535 1195
rect 1539 1191 1540 1195
rect 1534 1190 1540 1191
rect 144 1175 146 1190
rect 304 1175 306 1190
rect 488 1175 490 1190
rect 664 1175 666 1190
rect 824 1175 826 1190
rect 976 1175 978 1190
rect 1120 1175 1122 1190
rect 1256 1175 1258 1190
rect 1392 1175 1394 1190
rect 1536 1175 1538 1190
rect 1824 1175 1826 1203
rect 1864 1179 1866 1207
rect 1910 1199 1916 1200
rect 1910 1195 1911 1199
rect 1915 1195 1916 1199
rect 1910 1194 1916 1195
rect 1998 1199 2004 1200
rect 1998 1195 1999 1199
rect 2003 1195 2004 1199
rect 1998 1194 2004 1195
rect 2102 1199 2108 1200
rect 2102 1195 2103 1199
rect 2107 1195 2108 1199
rect 2102 1194 2108 1195
rect 2222 1199 2228 1200
rect 2222 1195 2223 1199
rect 2227 1195 2228 1199
rect 2222 1194 2228 1195
rect 2358 1199 2364 1200
rect 2358 1195 2359 1199
rect 2363 1195 2364 1199
rect 2358 1194 2364 1195
rect 2494 1199 2500 1200
rect 2494 1195 2495 1199
rect 2499 1195 2500 1199
rect 2494 1194 2500 1195
rect 2638 1199 2644 1200
rect 2638 1195 2639 1199
rect 2643 1195 2644 1199
rect 2638 1194 2644 1195
rect 2782 1199 2788 1200
rect 2782 1195 2783 1199
rect 2787 1195 2788 1199
rect 2782 1194 2788 1195
rect 2926 1199 2932 1200
rect 2926 1195 2927 1199
rect 2931 1195 2932 1199
rect 2926 1194 2932 1195
rect 3070 1199 3076 1200
rect 3070 1195 3071 1199
rect 3075 1195 3076 1199
rect 3070 1194 3076 1195
rect 3214 1199 3220 1200
rect 3214 1195 3215 1199
rect 3219 1195 3220 1199
rect 3214 1194 3220 1195
rect 3358 1199 3364 1200
rect 3358 1195 3359 1199
rect 3363 1195 3364 1199
rect 3358 1194 3364 1195
rect 3486 1199 3492 1200
rect 3486 1195 3487 1199
rect 3491 1195 3492 1199
rect 3486 1194 3492 1195
rect 1912 1179 1914 1194
rect 2000 1179 2002 1194
rect 2104 1179 2106 1194
rect 2224 1179 2226 1194
rect 2360 1179 2362 1194
rect 2496 1179 2498 1194
rect 2640 1179 2642 1194
rect 2784 1179 2786 1194
rect 2928 1179 2930 1194
rect 3072 1179 3074 1194
rect 3216 1179 3218 1194
rect 3360 1179 3362 1194
rect 3488 1179 3490 1194
rect 3576 1179 3578 1207
rect 1863 1178 1867 1179
rect 111 1174 115 1175
rect 111 1169 115 1170
rect 143 1174 147 1175
rect 143 1169 147 1170
rect 167 1174 171 1175
rect 167 1169 171 1170
rect 303 1174 307 1175
rect 303 1169 307 1170
rect 319 1174 323 1175
rect 319 1169 323 1170
rect 471 1174 475 1175
rect 471 1169 475 1170
rect 487 1174 491 1175
rect 487 1169 491 1170
rect 615 1174 619 1175
rect 615 1169 619 1170
rect 663 1174 667 1175
rect 663 1169 667 1170
rect 759 1174 763 1175
rect 759 1169 763 1170
rect 823 1174 827 1175
rect 823 1169 827 1170
rect 911 1174 915 1175
rect 911 1169 915 1170
rect 975 1174 979 1175
rect 975 1169 979 1170
rect 1063 1174 1067 1175
rect 1063 1169 1067 1170
rect 1119 1174 1123 1175
rect 1119 1169 1123 1170
rect 1231 1174 1235 1175
rect 1231 1169 1235 1170
rect 1255 1174 1259 1175
rect 1255 1169 1259 1170
rect 1391 1174 1395 1175
rect 1391 1169 1395 1170
rect 1399 1174 1403 1175
rect 1399 1169 1403 1170
rect 1535 1174 1539 1175
rect 1535 1169 1539 1170
rect 1575 1174 1579 1175
rect 1575 1169 1579 1170
rect 1735 1174 1739 1175
rect 1735 1169 1739 1170
rect 1823 1174 1827 1175
rect 1863 1173 1867 1174
rect 1895 1178 1899 1179
rect 1895 1173 1899 1174
rect 1911 1178 1915 1179
rect 1911 1173 1915 1174
rect 1999 1178 2003 1179
rect 1999 1173 2003 1174
rect 2063 1178 2067 1179
rect 2063 1173 2067 1174
rect 2103 1178 2107 1179
rect 2103 1173 2107 1174
rect 2223 1178 2227 1179
rect 2223 1173 2227 1174
rect 2255 1178 2259 1179
rect 2255 1173 2259 1174
rect 2359 1178 2363 1179
rect 2359 1173 2363 1174
rect 2439 1178 2443 1179
rect 2439 1173 2443 1174
rect 2495 1178 2499 1179
rect 2495 1173 2499 1174
rect 2615 1178 2619 1179
rect 2615 1173 2619 1174
rect 2639 1178 2643 1179
rect 2639 1173 2643 1174
rect 2783 1178 2787 1179
rect 2783 1173 2787 1174
rect 2791 1178 2795 1179
rect 2791 1173 2795 1174
rect 2927 1178 2931 1179
rect 2927 1173 2931 1174
rect 2967 1178 2971 1179
rect 2967 1173 2971 1174
rect 3071 1178 3075 1179
rect 3071 1173 3075 1174
rect 3143 1178 3147 1179
rect 3143 1173 3147 1174
rect 3215 1178 3219 1179
rect 3215 1173 3219 1174
rect 3327 1178 3331 1179
rect 3327 1173 3331 1174
rect 3359 1178 3363 1179
rect 3359 1173 3363 1174
rect 3487 1178 3491 1179
rect 3487 1173 3491 1174
rect 3575 1178 3579 1179
rect 3575 1173 3579 1174
rect 1823 1169 1827 1170
rect 112 1145 114 1169
rect 168 1158 170 1169
rect 320 1158 322 1169
rect 472 1158 474 1169
rect 616 1158 618 1169
rect 760 1158 762 1169
rect 912 1158 914 1169
rect 1064 1158 1066 1169
rect 1232 1158 1234 1169
rect 1400 1158 1402 1169
rect 1576 1158 1578 1169
rect 1736 1158 1738 1169
rect 166 1157 172 1158
rect 166 1153 167 1157
rect 171 1153 172 1157
rect 166 1152 172 1153
rect 318 1157 324 1158
rect 318 1153 319 1157
rect 323 1153 324 1157
rect 318 1152 324 1153
rect 470 1157 476 1158
rect 470 1153 471 1157
rect 475 1153 476 1157
rect 470 1152 476 1153
rect 614 1157 620 1158
rect 614 1153 615 1157
rect 619 1153 620 1157
rect 614 1152 620 1153
rect 758 1157 764 1158
rect 758 1153 759 1157
rect 763 1153 764 1157
rect 758 1152 764 1153
rect 910 1157 916 1158
rect 910 1153 911 1157
rect 915 1153 916 1157
rect 910 1152 916 1153
rect 1062 1157 1068 1158
rect 1062 1153 1063 1157
rect 1067 1153 1068 1157
rect 1062 1152 1068 1153
rect 1230 1157 1236 1158
rect 1230 1153 1231 1157
rect 1235 1153 1236 1157
rect 1230 1152 1236 1153
rect 1398 1157 1404 1158
rect 1398 1153 1399 1157
rect 1403 1153 1404 1157
rect 1398 1152 1404 1153
rect 1574 1157 1580 1158
rect 1574 1153 1575 1157
rect 1579 1153 1580 1157
rect 1574 1152 1580 1153
rect 1734 1157 1740 1158
rect 1734 1153 1735 1157
rect 1739 1153 1740 1157
rect 1734 1152 1740 1153
rect 1824 1145 1826 1169
rect 1864 1149 1866 1173
rect 1896 1162 1898 1173
rect 2064 1162 2066 1173
rect 2256 1162 2258 1173
rect 2440 1162 2442 1173
rect 2616 1162 2618 1173
rect 2792 1162 2794 1173
rect 2968 1162 2970 1173
rect 3144 1162 3146 1173
rect 3328 1162 3330 1173
rect 3488 1162 3490 1173
rect 1894 1161 1900 1162
rect 1894 1157 1895 1161
rect 1899 1157 1900 1161
rect 1894 1156 1900 1157
rect 2062 1161 2068 1162
rect 2062 1157 2063 1161
rect 2067 1157 2068 1161
rect 2062 1156 2068 1157
rect 2254 1161 2260 1162
rect 2254 1157 2255 1161
rect 2259 1157 2260 1161
rect 2254 1156 2260 1157
rect 2438 1161 2444 1162
rect 2438 1157 2439 1161
rect 2443 1157 2444 1161
rect 2438 1156 2444 1157
rect 2614 1161 2620 1162
rect 2614 1157 2615 1161
rect 2619 1157 2620 1161
rect 2614 1156 2620 1157
rect 2790 1161 2796 1162
rect 2790 1157 2791 1161
rect 2795 1157 2796 1161
rect 2790 1156 2796 1157
rect 2966 1161 2972 1162
rect 2966 1157 2967 1161
rect 2971 1157 2972 1161
rect 2966 1156 2972 1157
rect 3142 1161 3148 1162
rect 3142 1157 3143 1161
rect 3147 1157 3148 1161
rect 3142 1156 3148 1157
rect 3326 1161 3332 1162
rect 3326 1157 3327 1161
rect 3331 1157 3332 1161
rect 3326 1156 3332 1157
rect 3486 1161 3492 1162
rect 3486 1157 3487 1161
rect 3491 1157 3492 1161
rect 3486 1156 3492 1157
rect 3576 1149 3578 1173
rect 1862 1148 1868 1149
rect 110 1144 116 1145
rect 110 1140 111 1144
rect 115 1140 116 1144
rect 110 1139 116 1140
rect 1822 1144 1828 1145
rect 1822 1140 1823 1144
rect 1827 1140 1828 1144
rect 1862 1144 1863 1148
rect 1867 1144 1868 1148
rect 1862 1143 1868 1144
rect 3574 1148 3580 1149
rect 3574 1144 3575 1148
rect 3579 1144 3580 1148
rect 3574 1143 3580 1144
rect 1822 1139 1828 1140
rect 1862 1131 1868 1132
rect 110 1127 116 1128
rect 110 1123 111 1127
rect 115 1123 116 1127
rect 110 1122 116 1123
rect 1822 1127 1828 1128
rect 1822 1123 1823 1127
rect 1827 1123 1828 1127
rect 1862 1127 1863 1131
rect 1867 1127 1868 1131
rect 1862 1126 1868 1127
rect 3574 1131 3580 1132
rect 3574 1127 3575 1131
rect 3579 1127 3580 1131
rect 3574 1126 3580 1127
rect 1822 1122 1828 1123
rect 112 1103 114 1122
rect 158 1117 164 1118
rect 158 1113 159 1117
rect 163 1113 164 1117
rect 158 1112 164 1113
rect 310 1117 316 1118
rect 310 1113 311 1117
rect 315 1113 316 1117
rect 310 1112 316 1113
rect 462 1117 468 1118
rect 462 1113 463 1117
rect 467 1113 468 1117
rect 462 1112 468 1113
rect 606 1117 612 1118
rect 606 1113 607 1117
rect 611 1113 612 1117
rect 606 1112 612 1113
rect 750 1117 756 1118
rect 750 1113 751 1117
rect 755 1113 756 1117
rect 750 1112 756 1113
rect 902 1117 908 1118
rect 902 1113 903 1117
rect 907 1113 908 1117
rect 902 1112 908 1113
rect 1054 1117 1060 1118
rect 1054 1113 1055 1117
rect 1059 1113 1060 1117
rect 1054 1112 1060 1113
rect 1222 1117 1228 1118
rect 1222 1113 1223 1117
rect 1227 1113 1228 1117
rect 1222 1112 1228 1113
rect 1390 1117 1396 1118
rect 1390 1113 1391 1117
rect 1395 1113 1396 1117
rect 1390 1112 1396 1113
rect 1566 1117 1572 1118
rect 1566 1113 1567 1117
rect 1571 1113 1572 1117
rect 1566 1112 1572 1113
rect 1726 1117 1732 1118
rect 1726 1113 1727 1117
rect 1731 1113 1732 1117
rect 1726 1112 1732 1113
rect 160 1103 162 1112
rect 312 1103 314 1112
rect 464 1103 466 1112
rect 608 1103 610 1112
rect 752 1103 754 1112
rect 904 1103 906 1112
rect 1056 1103 1058 1112
rect 1224 1103 1226 1112
rect 1392 1103 1394 1112
rect 1568 1103 1570 1112
rect 1728 1103 1730 1112
rect 1824 1103 1826 1122
rect 111 1102 115 1103
rect 111 1097 115 1098
rect 159 1102 163 1103
rect 159 1097 163 1098
rect 215 1102 219 1103
rect 215 1097 219 1098
rect 311 1102 315 1103
rect 311 1097 315 1098
rect 327 1102 331 1103
rect 327 1097 331 1098
rect 439 1102 443 1103
rect 439 1097 443 1098
rect 463 1102 467 1103
rect 463 1097 467 1098
rect 559 1102 563 1103
rect 559 1097 563 1098
rect 607 1102 611 1103
rect 607 1097 611 1098
rect 679 1102 683 1103
rect 679 1097 683 1098
rect 751 1102 755 1103
rect 751 1097 755 1098
rect 807 1102 811 1103
rect 807 1097 811 1098
rect 903 1102 907 1103
rect 903 1097 907 1098
rect 943 1102 947 1103
rect 943 1097 947 1098
rect 1055 1102 1059 1103
rect 1055 1097 1059 1098
rect 1087 1102 1091 1103
rect 1087 1097 1091 1098
rect 1223 1102 1227 1103
rect 1223 1097 1227 1098
rect 1247 1102 1251 1103
rect 1247 1097 1251 1098
rect 1391 1102 1395 1103
rect 1391 1097 1395 1098
rect 1407 1102 1411 1103
rect 1407 1097 1411 1098
rect 1567 1102 1571 1103
rect 1567 1097 1571 1098
rect 1575 1102 1579 1103
rect 1575 1097 1579 1098
rect 1727 1102 1731 1103
rect 1727 1097 1731 1098
rect 1823 1102 1827 1103
rect 1864 1099 1866 1126
rect 1886 1121 1892 1122
rect 1886 1117 1887 1121
rect 1891 1117 1892 1121
rect 1886 1116 1892 1117
rect 2054 1121 2060 1122
rect 2054 1117 2055 1121
rect 2059 1117 2060 1121
rect 2054 1116 2060 1117
rect 2246 1121 2252 1122
rect 2246 1117 2247 1121
rect 2251 1117 2252 1121
rect 2246 1116 2252 1117
rect 2430 1121 2436 1122
rect 2430 1117 2431 1121
rect 2435 1117 2436 1121
rect 2430 1116 2436 1117
rect 2606 1121 2612 1122
rect 2606 1117 2607 1121
rect 2611 1117 2612 1121
rect 2606 1116 2612 1117
rect 2782 1121 2788 1122
rect 2782 1117 2783 1121
rect 2787 1117 2788 1121
rect 2782 1116 2788 1117
rect 2958 1121 2964 1122
rect 2958 1117 2959 1121
rect 2963 1117 2964 1121
rect 2958 1116 2964 1117
rect 3134 1121 3140 1122
rect 3134 1117 3135 1121
rect 3139 1117 3140 1121
rect 3134 1116 3140 1117
rect 3318 1121 3324 1122
rect 3318 1117 3319 1121
rect 3323 1117 3324 1121
rect 3318 1116 3324 1117
rect 3478 1121 3484 1122
rect 3478 1117 3479 1121
rect 3483 1117 3484 1121
rect 3478 1116 3484 1117
rect 1888 1099 1890 1116
rect 2056 1099 2058 1116
rect 2248 1099 2250 1116
rect 2432 1099 2434 1116
rect 2608 1099 2610 1116
rect 2784 1099 2786 1116
rect 2960 1099 2962 1116
rect 3136 1099 3138 1116
rect 3320 1099 3322 1116
rect 3480 1099 3482 1116
rect 3576 1099 3578 1126
rect 1823 1097 1827 1098
rect 1863 1098 1867 1099
rect 112 1082 114 1097
rect 216 1092 218 1097
rect 328 1092 330 1097
rect 440 1092 442 1097
rect 560 1092 562 1097
rect 680 1092 682 1097
rect 808 1092 810 1097
rect 944 1092 946 1097
rect 1088 1092 1090 1097
rect 1248 1092 1250 1097
rect 1408 1092 1410 1097
rect 1576 1092 1578 1097
rect 1728 1092 1730 1097
rect 214 1091 220 1092
rect 214 1087 215 1091
rect 219 1087 220 1091
rect 214 1086 220 1087
rect 326 1091 332 1092
rect 326 1087 327 1091
rect 331 1087 332 1091
rect 326 1086 332 1087
rect 438 1091 444 1092
rect 438 1087 439 1091
rect 443 1087 444 1091
rect 438 1086 444 1087
rect 558 1091 564 1092
rect 558 1087 559 1091
rect 563 1087 564 1091
rect 558 1086 564 1087
rect 678 1091 684 1092
rect 678 1087 679 1091
rect 683 1087 684 1091
rect 678 1086 684 1087
rect 806 1091 812 1092
rect 806 1087 807 1091
rect 811 1087 812 1091
rect 806 1086 812 1087
rect 942 1091 948 1092
rect 942 1087 943 1091
rect 947 1087 948 1091
rect 942 1086 948 1087
rect 1086 1091 1092 1092
rect 1086 1087 1087 1091
rect 1091 1087 1092 1091
rect 1086 1086 1092 1087
rect 1246 1091 1252 1092
rect 1246 1087 1247 1091
rect 1251 1087 1252 1091
rect 1246 1086 1252 1087
rect 1406 1091 1412 1092
rect 1406 1087 1407 1091
rect 1411 1087 1412 1091
rect 1406 1086 1412 1087
rect 1574 1091 1580 1092
rect 1574 1087 1575 1091
rect 1579 1087 1580 1091
rect 1574 1086 1580 1087
rect 1726 1091 1732 1092
rect 1726 1087 1727 1091
rect 1731 1087 1732 1091
rect 1726 1086 1732 1087
rect 1824 1082 1826 1097
rect 1863 1093 1867 1094
rect 1887 1098 1891 1099
rect 1887 1093 1891 1094
rect 1935 1098 1939 1099
rect 1935 1093 1939 1094
rect 2055 1098 2059 1099
rect 2055 1093 2059 1094
rect 2095 1098 2099 1099
rect 2095 1093 2099 1094
rect 2247 1098 2251 1099
rect 2247 1093 2251 1094
rect 2407 1098 2411 1099
rect 2407 1093 2411 1094
rect 2431 1098 2435 1099
rect 2431 1093 2435 1094
rect 2567 1098 2571 1099
rect 2567 1093 2571 1094
rect 2607 1098 2611 1099
rect 2607 1093 2611 1094
rect 2735 1098 2739 1099
rect 2735 1093 2739 1094
rect 2783 1098 2787 1099
rect 2783 1093 2787 1094
rect 2911 1098 2915 1099
rect 2911 1093 2915 1094
rect 2959 1098 2963 1099
rect 2959 1093 2963 1094
rect 3095 1098 3099 1099
rect 3095 1093 3099 1094
rect 3135 1098 3139 1099
rect 3135 1093 3139 1094
rect 3287 1098 3291 1099
rect 3287 1093 3291 1094
rect 3319 1098 3323 1099
rect 3319 1093 3323 1094
rect 3479 1098 3483 1099
rect 3479 1093 3483 1094
rect 3575 1098 3579 1099
rect 3575 1093 3579 1094
rect 110 1081 116 1082
rect 110 1077 111 1081
rect 115 1077 116 1081
rect 110 1076 116 1077
rect 1822 1081 1828 1082
rect 1822 1077 1823 1081
rect 1827 1077 1828 1081
rect 1864 1078 1866 1093
rect 1936 1088 1938 1093
rect 2096 1088 2098 1093
rect 2248 1088 2250 1093
rect 2408 1088 2410 1093
rect 2568 1088 2570 1093
rect 2736 1088 2738 1093
rect 2912 1088 2914 1093
rect 3096 1088 3098 1093
rect 3288 1088 3290 1093
rect 3480 1088 3482 1093
rect 1934 1087 1940 1088
rect 1934 1083 1935 1087
rect 1939 1083 1940 1087
rect 1934 1082 1940 1083
rect 2094 1087 2100 1088
rect 2094 1083 2095 1087
rect 2099 1083 2100 1087
rect 2094 1082 2100 1083
rect 2246 1087 2252 1088
rect 2246 1083 2247 1087
rect 2251 1083 2252 1087
rect 2246 1082 2252 1083
rect 2406 1087 2412 1088
rect 2406 1083 2407 1087
rect 2411 1083 2412 1087
rect 2406 1082 2412 1083
rect 2566 1087 2572 1088
rect 2566 1083 2567 1087
rect 2571 1083 2572 1087
rect 2566 1082 2572 1083
rect 2734 1087 2740 1088
rect 2734 1083 2735 1087
rect 2739 1083 2740 1087
rect 2734 1082 2740 1083
rect 2910 1087 2916 1088
rect 2910 1083 2911 1087
rect 2915 1083 2916 1087
rect 2910 1082 2916 1083
rect 3094 1087 3100 1088
rect 3094 1083 3095 1087
rect 3099 1083 3100 1087
rect 3094 1082 3100 1083
rect 3286 1087 3292 1088
rect 3286 1083 3287 1087
rect 3291 1083 3292 1087
rect 3286 1082 3292 1083
rect 3478 1087 3484 1088
rect 3478 1083 3479 1087
rect 3483 1083 3484 1087
rect 3478 1082 3484 1083
rect 3576 1078 3578 1093
rect 1822 1076 1828 1077
rect 1862 1077 1868 1078
rect 1862 1073 1863 1077
rect 1867 1073 1868 1077
rect 1862 1072 1868 1073
rect 3574 1077 3580 1078
rect 3574 1073 3575 1077
rect 3579 1073 3580 1077
rect 3574 1072 3580 1073
rect 110 1064 116 1065
rect 110 1060 111 1064
rect 115 1060 116 1064
rect 110 1059 116 1060
rect 1822 1064 1828 1065
rect 1822 1060 1823 1064
rect 1827 1060 1828 1064
rect 1822 1059 1828 1060
rect 1862 1060 1868 1061
rect 112 1027 114 1059
rect 222 1051 228 1052
rect 222 1047 223 1051
rect 227 1047 228 1051
rect 222 1046 228 1047
rect 334 1051 340 1052
rect 334 1047 335 1051
rect 339 1047 340 1051
rect 334 1046 340 1047
rect 446 1051 452 1052
rect 446 1047 447 1051
rect 451 1047 452 1051
rect 446 1046 452 1047
rect 566 1051 572 1052
rect 566 1047 567 1051
rect 571 1047 572 1051
rect 566 1046 572 1047
rect 686 1051 692 1052
rect 686 1047 687 1051
rect 691 1047 692 1051
rect 686 1046 692 1047
rect 814 1051 820 1052
rect 814 1047 815 1051
rect 819 1047 820 1051
rect 814 1046 820 1047
rect 950 1051 956 1052
rect 950 1047 951 1051
rect 955 1047 956 1051
rect 950 1046 956 1047
rect 1094 1051 1100 1052
rect 1094 1047 1095 1051
rect 1099 1047 1100 1051
rect 1094 1046 1100 1047
rect 1254 1051 1260 1052
rect 1254 1047 1255 1051
rect 1259 1047 1260 1051
rect 1254 1046 1260 1047
rect 1414 1051 1420 1052
rect 1414 1047 1415 1051
rect 1419 1047 1420 1051
rect 1414 1046 1420 1047
rect 1582 1051 1588 1052
rect 1582 1047 1583 1051
rect 1587 1047 1588 1051
rect 1582 1046 1588 1047
rect 1734 1051 1740 1052
rect 1734 1047 1735 1051
rect 1739 1047 1740 1051
rect 1734 1046 1740 1047
rect 224 1027 226 1046
rect 336 1027 338 1046
rect 448 1027 450 1046
rect 568 1027 570 1046
rect 688 1027 690 1046
rect 816 1027 818 1046
rect 952 1027 954 1046
rect 1096 1027 1098 1046
rect 1256 1027 1258 1046
rect 1416 1027 1418 1046
rect 1584 1027 1586 1046
rect 1736 1027 1738 1046
rect 1824 1027 1826 1059
rect 1862 1056 1863 1060
rect 1867 1056 1868 1060
rect 1862 1055 1868 1056
rect 3574 1060 3580 1061
rect 3574 1056 3575 1060
rect 3579 1056 3580 1060
rect 3574 1055 3580 1056
rect 1864 1027 1866 1055
rect 1942 1047 1948 1048
rect 1942 1043 1943 1047
rect 1947 1043 1948 1047
rect 1942 1042 1948 1043
rect 2102 1047 2108 1048
rect 2102 1043 2103 1047
rect 2107 1043 2108 1047
rect 2102 1042 2108 1043
rect 2254 1047 2260 1048
rect 2254 1043 2255 1047
rect 2259 1043 2260 1047
rect 2254 1042 2260 1043
rect 2414 1047 2420 1048
rect 2414 1043 2415 1047
rect 2419 1043 2420 1047
rect 2414 1042 2420 1043
rect 2574 1047 2580 1048
rect 2574 1043 2575 1047
rect 2579 1043 2580 1047
rect 2574 1042 2580 1043
rect 2742 1047 2748 1048
rect 2742 1043 2743 1047
rect 2747 1043 2748 1047
rect 2742 1042 2748 1043
rect 2918 1047 2924 1048
rect 2918 1043 2919 1047
rect 2923 1043 2924 1047
rect 2918 1042 2924 1043
rect 3102 1047 3108 1048
rect 3102 1043 3103 1047
rect 3107 1043 3108 1047
rect 3102 1042 3108 1043
rect 3294 1047 3300 1048
rect 3294 1043 3295 1047
rect 3299 1043 3300 1047
rect 3294 1042 3300 1043
rect 3486 1047 3492 1048
rect 3486 1043 3487 1047
rect 3491 1043 3492 1047
rect 3486 1042 3492 1043
rect 1944 1027 1946 1042
rect 2104 1027 2106 1042
rect 2256 1027 2258 1042
rect 2416 1027 2418 1042
rect 2576 1027 2578 1042
rect 2744 1027 2746 1042
rect 2920 1027 2922 1042
rect 3104 1027 3106 1042
rect 3296 1027 3298 1042
rect 3488 1027 3490 1042
rect 3576 1027 3578 1055
rect 111 1026 115 1027
rect 111 1021 115 1022
rect 223 1026 227 1027
rect 223 1021 227 1022
rect 335 1026 339 1027
rect 335 1021 339 1022
rect 343 1026 347 1027
rect 343 1021 347 1022
rect 431 1026 435 1027
rect 431 1021 435 1022
rect 447 1026 451 1027
rect 447 1021 451 1022
rect 535 1026 539 1027
rect 535 1021 539 1022
rect 567 1026 571 1027
rect 567 1021 571 1022
rect 655 1026 659 1027
rect 655 1021 659 1022
rect 687 1026 691 1027
rect 687 1021 691 1022
rect 791 1026 795 1027
rect 791 1021 795 1022
rect 815 1026 819 1027
rect 815 1021 819 1022
rect 951 1026 955 1027
rect 951 1021 955 1022
rect 1095 1026 1099 1027
rect 1095 1021 1099 1022
rect 1135 1026 1139 1027
rect 1135 1021 1139 1022
rect 1255 1026 1259 1027
rect 1255 1021 1259 1022
rect 1327 1026 1331 1027
rect 1327 1021 1331 1022
rect 1415 1026 1419 1027
rect 1415 1021 1419 1022
rect 1535 1026 1539 1027
rect 1535 1021 1539 1022
rect 1583 1026 1587 1027
rect 1583 1021 1587 1022
rect 1735 1026 1739 1027
rect 1735 1021 1739 1022
rect 1823 1026 1827 1027
rect 1823 1021 1827 1022
rect 1863 1026 1867 1027
rect 1863 1021 1867 1022
rect 1943 1026 1947 1027
rect 1943 1021 1947 1022
rect 2071 1026 2075 1027
rect 2071 1021 2075 1022
rect 2103 1026 2107 1027
rect 2103 1021 2107 1022
rect 2191 1026 2195 1027
rect 2191 1021 2195 1022
rect 2255 1026 2259 1027
rect 2255 1021 2259 1022
rect 2311 1026 2315 1027
rect 2311 1021 2315 1022
rect 2415 1026 2419 1027
rect 2415 1021 2419 1022
rect 2439 1026 2443 1027
rect 2439 1021 2443 1022
rect 2575 1026 2579 1027
rect 2575 1021 2579 1022
rect 2719 1026 2723 1027
rect 2719 1021 2723 1022
rect 2743 1026 2747 1027
rect 2743 1021 2747 1022
rect 2871 1026 2875 1027
rect 2871 1021 2875 1022
rect 2919 1026 2923 1027
rect 2919 1021 2923 1022
rect 3031 1026 3035 1027
rect 3031 1021 3035 1022
rect 3103 1026 3107 1027
rect 3103 1021 3107 1022
rect 3191 1026 3195 1027
rect 3191 1021 3195 1022
rect 3295 1026 3299 1027
rect 3295 1021 3299 1022
rect 3351 1026 3355 1027
rect 3351 1021 3355 1022
rect 3487 1026 3491 1027
rect 3487 1021 3491 1022
rect 3575 1026 3579 1027
rect 3575 1021 3579 1022
rect 112 997 114 1021
rect 344 1010 346 1021
rect 432 1010 434 1021
rect 536 1010 538 1021
rect 656 1010 658 1021
rect 792 1010 794 1021
rect 952 1010 954 1021
rect 1136 1010 1138 1021
rect 1328 1010 1330 1021
rect 1536 1010 1538 1021
rect 1736 1010 1738 1021
rect 342 1009 348 1010
rect 342 1005 343 1009
rect 347 1005 348 1009
rect 342 1004 348 1005
rect 430 1009 436 1010
rect 430 1005 431 1009
rect 435 1005 436 1009
rect 430 1004 436 1005
rect 534 1009 540 1010
rect 534 1005 535 1009
rect 539 1005 540 1009
rect 534 1004 540 1005
rect 654 1009 660 1010
rect 654 1005 655 1009
rect 659 1005 660 1009
rect 654 1004 660 1005
rect 790 1009 796 1010
rect 790 1005 791 1009
rect 795 1005 796 1009
rect 790 1004 796 1005
rect 950 1009 956 1010
rect 950 1005 951 1009
rect 955 1005 956 1009
rect 950 1004 956 1005
rect 1134 1009 1140 1010
rect 1134 1005 1135 1009
rect 1139 1005 1140 1009
rect 1134 1004 1140 1005
rect 1326 1009 1332 1010
rect 1326 1005 1327 1009
rect 1331 1005 1332 1009
rect 1326 1004 1332 1005
rect 1534 1009 1540 1010
rect 1534 1005 1535 1009
rect 1539 1005 1540 1009
rect 1534 1004 1540 1005
rect 1734 1009 1740 1010
rect 1734 1005 1735 1009
rect 1739 1005 1740 1009
rect 1734 1004 1740 1005
rect 1824 997 1826 1021
rect 1864 997 1866 1021
rect 1944 1010 1946 1021
rect 2072 1010 2074 1021
rect 2192 1010 2194 1021
rect 2312 1010 2314 1021
rect 2440 1010 2442 1021
rect 2576 1010 2578 1021
rect 2720 1010 2722 1021
rect 2872 1010 2874 1021
rect 3032 1010 3034 1021
rect 3192 1010 3194 1021
rect 3352 1010 3354 1021
rect 3488 1010 3490 1021
rect 1942 1009 1948 1010
rect 1942 1005 1943 1009
rect 1947 1005 1948 1009
rect 1942 1004 1948 1005
rect 2070 1009 2076 1010
rect 2070 1005 2071 1009
rect 2075 1005 2076 1009
rect 2070 1004 2076 1005
rect 2190 1009 2196 1010
rect 2190 1005 2191 1009
rect 2195 1005 2196 1009
rect 2190 1004 2196 1005
rect 2310 1009 2316 1010
rect 2310 1005 2311 1009
rect 2315 1005 2316 1009
rect 2310 1004 2316 1005
rect 2438 1009 2444 1010
rect 2438 1005 2439 1009
rect 2443 1005 2444 1009
rect 2438 1004 2444 1005
rect 2574 1009 2580 1010
rect 2574 1005 2575 1009
rect 2579 1005 2580 1009
rect 2574 1004 2580 1005
rect 2718 1009 2724 1010
rect 2718 1005 2719 1009
rect 2723 1005 2724 1009
rect 2718 1004 2724 1005
rect 2870 1009 2876 1010
rect 2870 1005 2871 1009
rect 2875 1005 2876 1009
rect 2870 1004 2876 1005
rect 3030 1009 3036 1010
rect 3030 1005 3031 1009
rect 3035 1005 3036 1009
rect 3030 1004 3036 1005
rect 3190 1009 3196 1010
rect 3190 1005 3191 1009
rect 3195 1005 3196 1009
rect 3190 1004 3196 1005
rect 3350 1009 3356 1010
rect 3350 1005 3351 1009
rect 3355 1005 3356 1009
rect 3350 1004 3356 1005
rect 3486 1009 3492 1010
rect 3486 1005 3487 1009
rect 3491 1005 3492 1009
rect 3486 1004 3492 1005
rect 3576 997 3578 1021
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 110 991 116 992
rect 1822 996 1828 997
rect 1822 992 1823 996
rect 1827 992 1828 996
rect 1822 991 1828 992
rect 1862 996 1868 997
rect 1862 992 1863 996
rect 1867 992 1868 996
rect 1862 991 1868 992
rect 3574 996 3580 997
rect 3574 992 3575 996
rect 3579 992 3580 996
rect 3574 991 3580 992
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 110 974 116 975
rect 1822 979 1828 980
rect 1822 975 1823 979
rect 1827 975 1828 979
rect 1822 974 1828 975
rect 1862 979 1868 980
rect 1862 975 1863 979
rect 1867 975 1868 979
rect 1862 974 1868 975
rect 3574 979 3580 980
rect 3574 975 3575 979
rect 3579 975 3580 979
rect 3574 974 3580 975
rect 112 955 114 974
rect 334 969 340 970
rect 334 965 335 969
rect 339 965 340 969
rect 334 964 340 965
rect 422 969 428 970
rect 422 965 423 969
rect 427 965 428 969
rect 422 964 428 965
rect 526 969 532 970
rect 526 965 527 969
rect 531 965 532 969
rect 526 964 532 965
rect 646 969 652 970
rect 646 965 647 969
rect 651 965 652 969
rect 646 964 652 965
rect 782 969 788 970
rect 782 965 783 969
rect 787 965 788 969
rect 782 964 788 965
rect 942 969 948 970
rect 942 965 943 969
rect 947 965 948 969
rect 942 964 948 965
rect 1126 969 1132 970
rect 1126 965 1127 969
rect 1131 965 1132 969
rect 1126 964 1132 965
rect 1318 969 1324 970
rect 1318 965 1319 969
rect 1323 965 1324 969
rect 1318 964 1324 965
rect 1526 969 1532 970
rect 1526 965 1527 969
rect 1531 965 1532 969
rect 1526 964 1532 965
rect 1726 969 1732 970
rect 1726 965 1727 969
rect 1731 965 1732 969
rect 1726 964 1732 965
rect 336 955 338 964
rect 424 955 426 964
rect 528 955 530 964
rect 648 955 650 964
rect 784 955 786 964
rect 944 955 946 964
rect 1128 955 1130 964
rect 1320 955 1322 964
rect 1528 955 1530 964
rect 1728 955 1730 964
rect 1824 955 1826 974
rect 1864 955 1866 974
rect 1934 969 1940 970
rect 1934 965 1935 969
rect 1939 965 1940 969
rect 1934 964 1940 965
rect 2062 969 2068 970
rect 2062 965 2063 969
rect 2067 965 2068 969
rect 2062 964 2068 965
rect 2182 969 2188 970
rect 2182 965 2183 969
rect 2187 965 2188 969
rect 2182 964 2188 965
rect 2302 969 2308 970
rect 2302 965 2303 969
rect 2307 965 2308 969
rect 2302 964 2308 965
rect 2430 969 2436 970
rect 2430 965 2431 969
rect 2435 965 2436 969
rect 2430 964 2436 965
rect 2566 969 2572 970
rect 2566 965 2567 969
rect 2571 965 2572 969
rect 2566 964 2572 965
rect 2710 969 2716 970
rect 2710 965 2711 969
rect 2715 965 2716 969
rect 2710 964 2716 965
rect 2862 969 2868 970
rect 2862 965 2863 969
rect 2867 965 2868 969
rect 2862 964 2868 965
rect 3022 969 3028 970
rect 3022 965 3023 969
rect 3027 965 3028 969
rect 3022 964 3028 965
rect 3182 969 3188 970
rect 3182 965 3183 969
rect 3187 965 3188 969
rect 3182 964 3188 965
rect 3342 969 3348 970
rect 3342 965 3343 969
rect 3347 965 3348 969
rect 3342 964 3348 965
rect 3478 969 3484 970
rect 3478 965 3479 969
rect 3483 965 3484 969
rect 3478 964 3484 965
rect 1936 955 1938 964
rect 2064 955 2066 964
rect 2184 955 2186 964
rect 2304 955 2306 964
rect 2432 955 2434 964
rect 2568 955 2570 964
rect 2712 955 2714 964
rect 2864 955 2866 964
rect 3024 955 3026 964
rect 3184 955 3186 964
rect 3344 955 3346 964
rect 3480 955 3482 964
rect 3576 955 3578 974
rect 111 954 115 955
rect 111 949 115 950
rect 335 954 339 955
rect 335 949 339 950
rect 367 954 371 955
rect 367 949 371 950
rect 423 954 427 955
rect 423 949 427 950
rect 463 954 467 955
rect 463 949 467 950
rect 527 954 531 955
rect 527 949 531 950
rect 575 954 579 955
rect 575 949 579 950
rect 647 954 651 955
rect 647 949 651 950
rect 703 954 707 955
rect 703 949 707 950
rect 783 954 787 955
rect 783 949 787 950
rect 847 954 851 955
rect 847 949 851 950
rect 943 954 947 955
rect 943 949 947 950
rect 1007 954 1011 955
rect 1007 949 1011 950
rect 1127 954 1131 955
rect 1127 949 1131 950
rect 1175 954 1179 955
rect 1175 949 1179 950
rect 1319 954 1323 955
rect 1319 949 1323 950
rect 1351 954 1355 955
rect 1351 949 1355 950
rect 1527 954 1531 955
rect 1527 949 1531 950
rect 1711 954 1715 955
rect 1711 949 1715 950
rect 1727 954 1731 955
rect 1727 949 1731 950
rect 1823 954 1827 955
rect 1823 949 1827 950
rect 1863 954 1867 955
rect 1863 949 1867 950
rect 1887 954 1891 955
rect 1887 949 1891 950
rect 1935 954 1939 955
rect 1935 949 1939 950
rect 2047 954 2051 955
rect 2047 949 2051 950
rect 2063 954 2067 955
rect 2063 949 2067 950
rect 2183 954 2187 955
rect 2183 949 2187 950
rect 2199 954 2203 955
rect 2199 949 2203 950
rect 2303 954 2307 955
rect 2303 949 2307 950
rect 2351 954 2355 955
rect 2351 949 2355 950
rect 2431 954 2435 955
rect 2431 949 2435 950
rect 2495 954 2499 955
rect 2495 949 2499 950
rect 2567 954 2571 955
rect 2567 949 2571 950
rect 2631 954 2635 955
rect 2631 949 2635 950
rect 2711 954 2715 955
rect 2711 949 2715 950
rect 2759 954 2763 955
rect 2759 949 2763 950
rect 2863 954 2867 955
rect 2863 949 2867 950
rect 2887 954 2891 955
rect 2887 949 2891 950
rect 3023 954 3027 955
rect 3023 949 3027 950
rect 3183 954 3187 955
rect 3183 949 3187 950
rect 3343 954 3347 955
rect 3343 949 3347 950
rect 3479 954 3483 955
rect 3479 949 3483 950
rect 3575 954 3579 955
rect 3575 949 3579 950
rect 112 934 114 949
rect 368 944 370 949
rect 464 944 466 949
rect 576 944 578 949
rect 704 944 706 949
rect 848 944 850 949
rect 1008 944 1010 949
rect 1176 944 1178 949
rect 1352 944 1354 949
rect 1528 944 1530 949
rect 1712 944 1714 949
rect 366 943 372 944
rect 366 939 367 943
rect 371 939 372 943
rect 366 938 372 939
rect 462 943 468 944
rect 462 939 463 943
rect 467 939 468 943
rect 462 938 468 939
rect 574 943 580 944
rect 574 939 575 943
rect 579 939 580 943
rect 574 938 580 939
rect 702 943 708 944
rect 702 939 703 943
rect 707 939 708 943
rect 702 938 708 939
rect 846 943 852 944
rect 846 939 847 943
rect 851 939 852 943
rect 846 938 852 939
rect 1006 943 1012 944
rect 1006 939 1007 943
rect 1011 939 1012 943
rect 1006 938 1012 939
rect 1174 943 1180 944
rect 1174 939 1175 943
rect 1179 939 1180 943
rect 1174 938 1180 939
rect 1350 943 1356 944
rect 1350 939 1351 943
rect 1355 939 1356 943
rect 1350 938 1356 939
rect 1526 943 1532 944
rect 1526 939 1527 943
rect 1531 939 1532 943
rect 1526 938 1532 939
rect 1710 943 1716 944
rect 1710 939 1711 943
rect 1715 939 1716 943
rect 1710 938 1716 939
rect 1824 934 1826 949
rect 1864 934 1866 949
rect 1888 944 1890 949
rect 2048 944 2050 949
rect 2200 944 2202 949
rect 2352 944 2354 949
rect 2496 944 2498 949
rect 2632 944 2634 949
rect 2760 944 2762 949
rect 2888 944 2890 949
rect 3024 944 3026 949
rect 1886 943 1892 944
rect 1886 939 1887 943
rect 1891 939 1892 943
rect 1886 938 1892 939
rect 2046 943 2052 944
rect 2046 939 2047 943
rect 2051 939 2052 943
rect 2046 938 2052 939
rect 2198 943 2204 944
rect 2198 939 2199 943
rect 2203 939 2204 943
rect 2198 938 2204 939
rect 2350 943 2356 944
rect 2350 939 2351 943
rect 2355 939 2356 943
rect 2350 938 2356 939
rect 2494 943 2500 944
rect 2494 939 2495 943
rect 2499 939 2500 943
rect 2494 938 2500 939
rect 2630 943 2636 944
rect 2630 939 2631 943
rect 2635 939 2636 943
rect 2630 938 2636 939
rect 2758 943 2764 944
rect 2758 939 2759 943
rect 2763 939 2764 943
rect 2758 938 2764 939
rect 2886 943 2892 944
rect 2886 939 2887 943
rect 2891 939 2892 943
rect 2886 938 2892 939
rect 3022 943 3028 944
rect 3022 939 3023 943
rect 3027 939 3028 943
rect 3022 938 3028 939
rect 3576 934 3578 949
rect 110 933 116 934
rect 110 929 111 933
rect 115 929 116 933
rect 110 928 116 929
rect 1822 933 1828 934
rect 1822 929 1823 933
rect 1827 929 1828 933
rect 1822 928 1828 929
rect 1862 933 1868 934
rect 1862 929 1863 933
rect 1867 929 1868 933
rect 1862 928 1868 929
rect 3574 933 3580 934
rect 3574 929 3575 933
rect 3579 929 3580 933
rect 3574 928 3580 929
rect 110 916 116 917
rect 110 912 111 916
rect 115 912 116 916
rect 110 911 116 912
rect 1822 916 1828 917
rect 1822 912 1823 916
rect 1827 912 1828 916
rect 1822 911 1828 912
rect 1862 916 1868 917
rect 1862 912 1863 916
rect 1867 912 1868 916
rect 1862 911 1868 912
rect 3574 916 3580 917
rect 3574 912 3575 916
rect 3579 912 3580 916
rect 3574 911 3580 912
rect 112 883 114 911
rect 374 903 380 904
rect 374 899 375 903
rect 379 899 380 903
rect 374 898 380 899
rect 470 903 476 904
rect 470 899 471 903
rect 475 899 476 903
rect 470 898 476 899
rect 582 903 588 904
rect 582 899 583 903
rect 587 899 588 903
rect 582 898 588 899
rect 710 903 716 904
rect 710 899 711 903
rect 715 899 716 903
rect 710 898 716 899
rect 854 903 860 904
rect 854 899 855 903
rect 859 899 860 903
rect 854 898 860 899
rect 1014 903 1020 904
rect 1014 899 1015 903
rect 1019 899 1020 903
rect 1014 898 1020 899
rect 1182 903 1188 904
rect 1182 899 1183 903
rect 1187 899 1188 903
rect 1182 898 1188 899
rect 1358 903 1364 904
rect 1358 899 1359 903
rect 1363 899 1364 903
rect 1358 898 1364 899
rect 1534 903 1540 904
rect 1534 899 1535 903
rect 1539 899 1540 903
rect 1534 898 1540 899
rect 1718 903 1724 904
rect 1718 899 1719 903
rect 1723 899 1724 903
rect 1718 898 1724 899
rect 376 883 378 898
rect 472 883 474 898
rect 584 883 586 898
rect 712 883 714 898
rect 856 883 858 898
rect 1016 883 1018 898
rect 1184 883 1186 898
rect 1360 883 1362 898
rect 1536 883 1538 898
rect 1720 883 1722 898
rect 1824 883 1826 911
rect 1864 887 1866 911
rect 1894 903 1900 904
rect 1894 899 1895 903
rect 1899 899 1900 903
rect 1894 898 1900 899
rect 2054 903 2060 904
rect 2054 899 2055 903
rect 2059 899 2060 903
rect 2054 898 2060 899
rect 2206 903 2212 904
rect 2206 899 2207 903
rect 2211 899 2212 903
rect 2206 898 2212 899
rect 2358 903 2364 904
rect 2358 899 2359 903
rect 2363 899 2364 903
rect 2358 898 2364 899
rect 2502 903 2508 904
rect 2502 899 2503 903
rect 2507 899 2508 903
rect 2502 898 2508 899
rect 2638 903 2644 904
rect 2638 899 2639 903
rect 2643 899 2644 903
rect 2638 898 2644 899
rect 2766 903 2772 904
rect 2766 899 2767 903
rect 2771 899 2772 903
rect 2766 898 2772 899
rect 2894 903 2900 904
rect 2894 899 2895 903
rect 2899 899 2900 903
rect 2894 898 2900 899
rect 3030 903 3036 904
rect 3030 899 3031 903
rect 3035 899 3036 903
rect 3030 898 3036 899
rect 1896 887 1898 898
rect 2056 887 2058 898
rect 2208 887 2210 898
rect 2360 887 2362 898
rect 2504 887 2506 898
rect 2640 887 2642 898
rect 2768 887 2770 898
rect 2896 887 2898 898
rect 3032 887 3034 898
rect 3576 887 3578 911
rect 1863 886 1867 887
rect 111 882 115 883
rect 111 877 115 878
rect 343 882 347 883
rect 343 877 347 878
rect 375 882 379 883
rect 375 877 379 878
rect 431 882 435 883
rect 431 877 435 878
rect 471 882 475 883
rect 471 877 475 878
rect 535 882 539 883
rect 535 877 539 878
rect 583 882 587 883
rect 583 877 587 878
rect 647 882 651 883
rect 647 877 651 878
rect 711 882 715 883
rect 711 877 715 878
rect 783 882 787 883
rect 783 877 787 878
rect 855 882 859 883
rect 855 877 859 878
rect 927 882 931 883
rect 927 877 931 878
rect 1015 882 1019 883
rect 1015 877 1019 878
rect 1087 882 1091 883
rect 1087 877 1091 878
rect 1183 882 1187 883
rect 1183 877 1187 878
rect 1263 882 1267 883
rect 1263 877 1267 878
rect 1359 882 1363 883
rect 1359 877 1363 878
rect 1447 882 1451 883
rect 1447 877 1451 878
rect 1535 882 1539 883
rect 1535 877 1539 878
rect 1631 882 1635 883
rect 1631 877 1635 878
rect 1719 882 1723 883
rect 1719 877 1723 878
rect 1823 882 1827 883
rect 1863 881 1867 882
rect 1895 886 1899 887
rect 1895 881 1899 882
rect 2015 886 2019 887
rect 2015 881 2019 882
rect 2055 886 2059 887
rect 2055 881 2059 882
rect 2167 886 2171 887
rect 2167 881 2171 882
rect 2207 886 2211 887
rect 2207 881 2211 882
rect 2319 886 2323 887
rect 2319 881 2323 882
rect 2359 886 2363 887
rect 2359 881 2363 882
rect 2487 886 2491 887
rect 2487 881 2491 882
rect 2503 886 2507 887
rect 2503 881 2507 882
rect 2639 886 2643 887
rect 2639 881 2643 882
rect 2663 886 2667 887
rect 2663 881 2667 882
rect 2767 886 2771 887
rect 2767 881 2771 882
rect 2847 886 2851 887
rect 2847 881 2851 882
rect 2895 886 2899 887
rect 2895 881 2899 882
rect 3031 886 3035 887
rect 3031 881 3035 882
rect 3039 886 3043 887
rect 3039 881 3043 882
rect 3239 886 3243 887
rect 3239 881 3243 882
rect 3439 886 3443 887
rect 3439 881 3443 882
rect 3575 886 3579 887
rect 3575 881 3579 882
rect 1823 877 1827 878
rect 112 853 114 877
rect 344 866 346 877
rect 432 866 434 877
rect 536 866 538 877
rect 648 866 650 877
rect 784 866 786 877
rect 928 866 930 877
rect 1088 866 1090 877
rect 1264 866 1266 877
rect 1448 866 1450 877
rect 1632 866 1634 877
rect 342 865 348 866
rect 342 861 343 865
rect 347 861 348 865
rect 342 860 348 861
rect 430 865 436 866
rect 430 861 431 865
rect 435 861 436 865
rect 430 860 436 861
rect 534 865 540 866
rect 534 861 535 865
rect 539 861 540 865
rect 534 860 540 861
rect 646 865 652 866
rect 646 861 647 865
rect 651 861 652 865
rect 646 860 652 861
rect 782 865 788 866
rect 782 861 783 865
rect 787 861 788 865
rect 782 860 788 861
rect 926 865 932 866
rect 926 861 927 865
rect 931 861 932 865
rect 926 860 932 861
rect 1086 865 1092 866
rect 1086 861 1087 865
rect 1091 861 1092 865
rect 1086 860 1092 861
rect 1262 865 1268 866
rect 1262 861 1263 865
rect 1267 861 1268 865
rect 1262 860 1268 861
rect 1446 865 1452 866
rect 1446 861 1447 865
rect 1451 861 1452 865
rect 1446 860 1452 861
rect 1630 865 1636 866
rect 1630 861 1631 865
rect 1635 861 1636 865
rect 1630 860 1636 861
rect 1824 853 1826 877
rect 1864 857 1866 881
rect 1896 870 1898 881
rect 2016 870 2018 881
rect 2168 870 2170 881
rect 2320 870 2322 881
rect 2488 870 2490 881
rect 2664 870 2666 881
rect 2848 870 2850 881
rect 3040 870 3042 881
rect 3240 870 3242 881
rect 3440 870 3442 881
rect 1894 869 1900 870
rect 1894 865 1895 869
rect 1899 865 1900 869
rect 1894 864 1900 865
rect 2014 869 2020 870
rect 2014 865 2015 869
rect 2019 865 2020 869
rect 2014 864 2020 865
rect 2166 869 2172 870
rect 2166 865 2167 869
rect 2171 865 2172 869
rect 2166 864 2172 865
rect 2318 869 2324 870
rect 2318 865 2319 869
rect 2323 865 2324 869
rect 2318 864 2324 865
rect 2486 869 2492 870
rect 2486 865 2487 869
rect 2491 865 2492 869
rect 2486 864 2492 865
rect 2662 869 2668 870
rect 2662 865 2663 869
rect 2667 865 2668 869
rect 2662 864 2668 865
rect 2846 869 2852 870
rect 2846 865 2847 869
rect 2851 865 2852 869
rect 2846 864 2852 865
rect 3038 869 3044 870
rect 3038 865 3039 869
rect 3043 865 3044 869
rect 3038 864 3044 865
rect 3238 869 3244 870
rect 3238 865 3239 869
rect 3243 865 3244 869
rect 3238 864 3244 865
rect 3438 869 3444 870
rect 3438 865 3439 869
rect 3443 865 3444 869
rect 3438 864 3444 865
rect 3576 857 3578 881
rect 1862 856 1868 857
rect 110 852 116 853
rect 110 848 111 852
rect 115 848 116 852
rect 110 847 116 848
rect 1822 852 1828 853
rect 1822 848 1823 852
rect 1827 848 1828 852
rect 1862 852 1863 856
rect 1867 852 1868 856
rect 1862 851 1868 852
rect 3574 856 3580 857
rect 3574 852 3575 856
rect 3579 852 3580 856
rect 3574 851 3580 852
rect 1822 847 1828 848
rect 1862 839 1868 840
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 110 830 116 831
rect 1822 835 1828 836
rect 1822 831 1823 835
rect 1827 831 1828 835
rect 1862 835 1863 839
rect 1867 835 1868 839
rect 1862 834 1868 835
rect 3574 839 3580 840
rect 3574 835 3575 839
rect 3579 835 3580 839
rect 3574 834 3580 835
rect 1822 830 1828 831
rect 112 815 114 830
rect 334 825 340 826
rect 334 821 335 825
rect 339 821 340 825
rect 334 820 340 821
rect 422 825 428 826
rect 422 821 423 825
rect 427 821 428 825
rect 422 820 428 821
rect 526 825 532 826
rect 526 821 527 825
rect 531 821 532 825
rect 526 820 532 821
rect 638 825 644 826
rect 638 821 639 825
rect 643 821 644 825
rect 638 820 644 821
rect 774 825 780 826
rect 774 821 775 825
rect 779 821 780 825
rect 774 820 780 821
rect 918 825 924 826
rect 918 821 919 825
rect 923 821 924 825
rect 918 820 924 821
rect 1078 825 1084 826
rect 1078 821 1079 825
rect 1083 821 1084 825
rect 1078 820 1084 821
rect 1254 825 1260 826
rect 1254 821 1255 825
rect 1259 821 1260 825
rect 1254 820 1260 821
rect 1438 825 1444 826
rect 1438 821 1439 825
rect 1443 821 1444 825
rect 1438 820 1444 821
rect 1622 825 1628 826
rect 1622 821 1623 825
rect 1627 821 1628 825
rect 1622 820 1628 821
rect 336 815 338 820
rect 424 815 426 820
rect 528 815 530 820
rect 640 815 642 820
rect 776 815 778 820
rect 920 815 922 820
rect 1080 815 1082 820
rect 1256 815 1258 820
rect 1440 815 1442 820
rect 1624 815 1626 820
rect 1824 815 1826 830
rect 1864 819 1866 834
rect 1886 829 1892 830
rect 1886 825 1887 829
rect 1891 825 1892 829
rect 1886 824 1892 825
rect 2006 829 2012 830
rect 2006 825 2007 829
rect 2011 825 2012 829
rect 2006 824 2012 825
rect 2158 829 2164 830
rect 2158 825 2159 829
rect 2163 825 2164 829
rect 2158 824 2164 825
rect 2310 829 2316 830
rect 2310 825 2311 829
rect 2315 825 2316 829
rect 2310 824 2316 825
rect 2478 829 2484 830
rect 2478 825 2479 829
rect 2483 825 2484 829
rect 2478 824 2484 825
rect 2654 829 2660 830
rect 2654 825 2655 829
rect 2659 825 2660 829
rect 2654 824 2660 825
rect 2838 829 2844 830
rect 2838 825 2839 829
rect 2843 825 2844 829
rect 2838 824 2844 825
rect 3030 829 3036 830
rect 3030 825 3031 829
rect 3035 825 3036 829
rect 3030 824 3036 825
rect 3230 829 3236 830
rect 3230 825 3231 829
rect 3235 825 3236 829
rect 3230 824 3236 825
rect 3430 829 3436 830
rect 3430 825 3431 829
rect 3435 825 3436 829
rect 3430 824 3436 825
rect 1888 819 1890 824
rect 2008 819 2010 824
rect 2160 819 2162 824
rect 2312 819 2314 824
rect 2480 819 2482 824
rect 2656 819 2658 824
rect 2840 819 2842 824
rect 3032 819 3034 824
rect 3232 819 3234 824
rect 3432 819 3434 824
rect 3576 819 3578 834
rect 1863 818 1867 819
rect 111 814 115 815
rect 111 809 115 810
rect 287 814 291 815
rect 287 809 291 810
rect 335 814 339 815
rect 335 809 339 810
rect 407 814 411 815
rect 407 809 411 810
rect 423 814 427 815
rect 423 809 427 810
rect 527 814 531 815
rect 527 809 531 810
rect 535 814 539 815
rect 535 809 539 810
rect 639 814 643 815
rect 639 809 643 810
rect 679 814 683 815
rect 679 809 683 810
rect 775 814 779 815
rect 775 809 779 810
rect 823 814 827 815
rect 823 809 827 810
rect 919 814 923 815
rect 919 809 923 810
rect 975 814 979 815
rect 975 809 979 810
rect 1079 814 1083 815
rect 1079 809 1083 810
rect 1127 814 1131 815
rect 1127 809 1131 810
rect 1255 814 1259 815
rect 1255 809 1259 810
rect 1279 814 1283 815
rect 1279 809 1283 810
rect 1439 814 1443 815
rect 1439 809 1443 810
rect 1599 814 1603 815
rect 1599 809 1603 810
rect 1623 814 1627 815
rect 1623 809 1627 810
rect 1823 814 1827 815
rect 1863 813 1867 814
rect 1887 818 1891 819
rect 1887 813 1891 814
rect 1991 818 1995 819
rect 1991 813 1995 814
rect 2007 818 2011 819
rect 2007 813 2011 814
rect 2135 818 2139 819
rect 2135 813 2139 814
rect 2159 818 2163 819
rect 2159 813 2163 814
rect 2287 818 2291 819
rect 2287 813 2291 814
rect 2311 818 2315 819
rect 2311 813 2315 814
rect 2455 818 2459 819
rect 2455 813 2459 814
rect 2479 818 2483 819
rect 2479 813 2483 814
rect 2623 818 2627 819
rect 2623 813 2627 814
rect 2655 818 2659 819
rect 2655 813 2659 814
rect 2799 818 2803 819
rect 2799 813 2803 814
rect 2839 818 2843 819
rect 2839 813 2843 814
rect 2967 818 2971 819
rect 2967 813 2971 814
rect 3031 818 3035 819
rect 3031 813 3035 814
rect 3143 818 3147 819
rect 3143 813 3147 814
rect 3231 818 3235 819
rect 3231 813 3235 814
rect 3319 818 3323 819
rect 3319 813 3323 814
rect 3431 818 3435 819
rect 3431 813 3435 814
rect 3479 818 3483 819
rect 3479 813 3483 814
rect 3575 818 3579 819
rect 3575 813 3579 814
rect 1823 809 1827 810
rect 112 794 114 809
rect 288 804 290 809
rect 408 804 410 809
rect 536 804 538 809
rect 680 804 682 809
rect 824 804 826 809
rect 976 804 978 809
rect 1128 804 1130 809
rect 1280 804 1282 809
rect 1440 804 1442 809
rect 1600 804 1602 809
rect 286 803 292 804
rect 286 799 287 803
rect 291 799 292 803
rect 286 798 292 799
rect 406 803 412 804
rect 406 799 407 803
rect 411 799 412 803
rect 406 798 412 799
rect 534 803 540 804
rect 534 799 535 803
rect 539 799 540 803
rect 534 798 540 799
rect 678 803 684 804
rect 678 799 679 803
rect 683 799 684 803
rect 678 798 684 799
rect 822 803 828 804
rect 822 799 823 803
rect 827 799 828 803
rect 822 798 828 799
rect 974 803 980 804
rect 974 799 975 803
rect 979 799 980 803
rect 974 798 980 799
rect 1126 803 1132 804
rect 1126 799 1127 803
rect 1131 799 1132 803
rect 1126 798 1132 799
rect 1278 803 1284 804
rect 1278 799 1279 803
rect 1283 799 1284 803
rect 1278 798 1284 799
rect 1438 803 1444 804
rect 1438 799 1439 803
rect 1443 799 1444 803
rect 1438 798 1444 799
rect 1598 803 1604 804
rect 1598 799 1599 803
rect 1603 799 1604 803
rect 1598 798 1604 799
rect 1824 794 1826 809
rect 1864 798 1866 813
rect 1888 808 1890 813
rect 1992 808 1994 813
rect 2136 808 2138 813
rect 2288 808 2290 813
rect 2456 808 2458 813
rect 2624 808 2626 813
rect 2800 808 2802 813
rect 2968 808 2970 813
rect 3144 808 3146 813
rect 3320 808 3322 813
rect 3480 808 3482 813
rect 1886 807 1892 808
rect 1886 803 1887 807
rect 1891 803 1892 807
rect 1886 802 1892 803
rect 1990 807 1996 808
rect 1990 803 1991 807
rect 1995 803 1996 807
rect 1990 802 1996 803
rect 2134 807 2140 808
rect 2134 803 2135 807
rect 2139 803 2140 807
rect 2134 802 2140 803
rect 2286 807 2292 808
rect 2286 803 2287 807
rect 2291 803 2292 807
rect 2286 802 2292 803
rect 2454 807 2460 808
rect 2454 803 2455 807
rect 2459 803 2460 807
rect 2454 802 2460 803
rect 2622 807 2628 808
rect 2622 803 2623 807
rect 2627 803 2628 807
rect 2622 802 2628 803
rect 2798 807 2804 808
rect 2798 803 2799 807
rect 2803 803 2804 807
rect 2798 802 2804 803
rect 2966 807 2972 808
rect 2966 803 2967 807
rect 2971 803 2972 807
rect 2966 802 2972 803
rect 3142 807 3148 808
rect 3142 803 3143 807
rect 3147 803 3148 807
rect 3142 802 3148 803
rect 3318 807 3324 808
rect 3318 803 3319 807
rect 3323 803 3324 807
rect 3318 802 3324 803
rect 3478 807 3484 808
rect 3478 803 3479 807
rect 3483 803 3484 807
rect 3478 802 3484 803
rect 3576 798 3578 813
rect 1862 797 1868 798
rect 110 793 116 794
rect 110 789 111 793
rect 115 789 116 793
rect 110 788 116 789
rect 1822 793 1828 794
rect 1822 789 1823 793
rect 1827 789 1828 793
rect 1862 793 1863 797
rect 1867 793 1868 797
rect 1862 792 1868 793
rect 3574 797 3580 798
rect 3574 793 3575 797
rect 3579 793 3580 797
rect 3574 792 3580 793
rect 1822 788 1828 789
rect 1862 780 1868 781
rect 110 776 116 777
rect 110 772 111 776
rect 115 772 116 776
rect 110 771 116 772
rect 1822 776 1828 777
rect 1822 772 1823 776
rect 1827 772 1828 776
rect 1862 776 1863 780
rect 1867 776 1868 780
rect 1862 775 1868 776
rect 3574 780 3580 781
rect 3574 776 3575 780
rect 3579 776 3580 780
rect 3574 775 3580 776
rect 1822 771 1828 772
rect 112 743 114 771
rect 294 763 300 764
rect 294 759 295 763
rect 299 759 300 763
rect 294 758 300 759
rect 414 763 420 764
rect 414 759 415 763
rect 419 759 420 763
rect 414 758 420 759
rect 542 763 548 764
rect 542 759 543 763
rect 547 759 548 763
rect 542 758 548 759
rect 686 763 692 764
rect 686 759 687 763
rect 691 759 692 763
rect 686 758 692 759
rect 830 763 836 764
rect 830 759 831 763
rect 835 759 836 763
rect 830 758 836 759
rect 982 763 988 764
rect 982 759 983 763
rect 987 759 988 763
rect 982 758 988 759
rect 1134 763 1140 764
rect 1134 759 1135 763
rect 1139 759 1140 763
rect 1134 758 1140 759
rect 1286 763 1292 764
rect 1286 759 1287 763
rect 1291 759 1292 763
rect 1286 758 1292 759
rect 1446 763 1452 764
rect 1446 759 1447 763
rect 1451 759 1452 763
rect 1446 758 1452 759
rect 1606 763 1612 764
rect 1606 759 1607 763
rect 1611 759 1612 763
rect 1606 758 1612 759
rect 296 743 298 758
rect 416 743 418 758
rect 544 743 546 758
rect 688 743 690 758
rect 832 743 834 758
rect 984 743 986 758
rect 1136 743 1138 758
rect 1288 743 1290 758
rect 1448 743 1450 758
rect 1608 743 1610 758
rect 1824 743 1826 771
rect 1864 747 1866 775
rect 1894 767 1900 768
rect 1894 763 1895 767
rect 1899 763 1900 767
rect 1894 762 1900 763
rect 1998 767 2004 768
rect 1998 763 1999 767
rect 2003 763 2004 767
rect 1998 762 2004 763
rect 2142 767 2148 768
rect 2142 763 2143 767
rect 2147 763 2148 767
rect 2142 762 2148 763
rect 2294 767 2300 768
rect 2294 763 2295 767
rect 2299 763 2300 767
rect 2294 762 2300 763
rect 2462 767 2468 768
rect 2462 763 2463 767
rect 2467 763 2468 767
rect 2462 762 2468 763
rect 2630 767 2636 768
rect 2630 763 2631 767
rect 2635 763 2636 767
rect 2630 762 2636 763
rect 2806 767 2812 768
rect 2806 763 2807 767
rect 2811 763 2812 767
rect 2806 762 2812 763
rect 2974 767 2980 768
rect 2974 763 2975 767
rect 2979 763 2980 767
rect 2974 762 2980 763
rect 3150 767 3156 768
rect 3150 763 3151 767
rect 3155 763 3156 767
rect 3150 762 3156 763
rect 3326 767 3332 768
rect 3326 763 3327 767
rect 3331 763 3332 767
rect 3326 762 3332 763
rect 3486 767 3492 768
rect 3486 763 3487 767
rect 3491 763 3492 767
rect 3486 762 3492 763
rect 1896 747 1898 762
rect 2000 747 2002 762
rect 2144 747 2146 762
rect 2296 747 2298 762
rect 2464 747 2466 762
rect 2632 747 2634 762
rect 2808 747 2810 762
rect 2976 747 2978 762
rect 3152 747 3154 762
rect 3328 747 3330 762
rect 3488 747 3490 762
rect 3576 747 3578 775
rect 1863 746 1867 747
rect 111 742 115 743
rect 111 737 115 738
rect 215 742 219 743
rect 215 737 219 738
rect 295 742 299 743
rect 295 737 299 738
rect 359 742 363 743
rect 359 737 363 738
rect 415 742 419 743
rect 415 737 419 738
rect 503 742 507 743
rect 503 737 507 738
rect 543 742 547 743
rect 543 737 547 738
rect 647 742 651 743
rect 647 737 651 738
rect 687 742 691 743
rect 687 737 691 738
rect 791 742 795 743
rect 791 737 795 738
rect 831 742 835 743
rect 831 737 835 738
rect 935 742 939 743
rect 935 737 939 738
rect 983 742 987 743
rect 983 737 987 738
rect 1087 742 1091 743
rect 1087 737 1091 738
rect 1135 742 1139 743
rect 1135 737 1139 738
rect 1247 742 1251 743
rect 1247 737 1251 738
rect 1287 742 1291 743
rect 1287 737 1291 738
rect 1415 742 1419 743
rect 1415 737 1419 738
rect 1447 742 1451 743
rect 1447 737 1451 738
rect 1583 742 1587 743
rect 1583 737 1587 738
rect 1607 742 1611 743
rect 1607 737 1611 738
rect 1735 742 1739 743
rect 1735 737 1739 738
rect 1823 742 1827 743
rect 1863 741 1867 742
rect 1895 746 1899 747
rect 1895 741 1899 742
rect 1999 746 2003 747
rect 1999 741 2003 742
rect 2063 746 2067 747
rect 2063 741 2067 742
rect 2143 746 2147 747
rect 2143 741 2147 742
rect 2255 746 2259 747
rect 2255 741 2259 742
rect 2295 746 2299 747
rect 2295 741 2299 742
rect 2447 746 2451 747
rect 2447 741 2451 742
rect 2463 746 2467 747
rect 2463 741 2467 742
rect 2631 746 2635 747
rect 2631 741 2635 742
rect 2639 746 2643 747
rect 2639 741 2643 742
rect 2807 746 2811 747
rect 2807 741 2811 742
rect 2823 746 2827 747
rect 2823 741 2827 742
rect 2975 746 2979 747
rect 2975 741 2979 742
rect 2999 746 3003 747
rect 2999 741 3003 742
rect 3151 746 3155 747
rect 3151 741 3155 742
rect 3167 746 3171 747
rect 3167 741 3171 742
rect 3327 746 3331 747
rect 3327 741 3331 742
rect 3335 746 3339 747
rect 3335 741 3339 742
rect 3487 746 3491 747
rect 3487 741 3491 742
rect 3575 746 3579 747
rect 3575 741 3579 742
rect 1823 737 1827 738
rect 112 713 114 737
rect 216 726 218 737
rect 360 726 362 737
rect 504 726 506 737
rect 648 726 650 737
rect 792 726 794 737
rect 936 726 938 737
rect 1088 726 1090 737
rect 1248 726 1250 737
rect 1416 726 1418 737
rect 1584 726 1586 737
rect 1736 726 1738 737
rect 214 725 220 726
rect 214 721 215 725
rect 219 721 220 725
rect 214 720 220 721
rect 358 725 364 726
rect 358 721 359 725
rect 363 721 364 725
rect 358 720 364 721
rect 502 725 508 726
rect 502 721 503 725
rect 507 721 508 725
rect 502 720 508 721
rect 646 725 652 726
rect 646 721 647 725
rect 651 721 652 725
rect 646 720 652 721
rect 790 725 796 726
rect 790 721 791 725
rect 795 721 796 725
rect 790 720 796 721
rect 934 725 940 726
rect 934 721 935 725
rect 939 721 940 725
rect 934 720 940 721
rect 1086 725 1092 726
rect 1086 721 1087 725
rect 1091 721 1092 725
rect 1086 720 1092 721
rect 1246 725 1252 726
rect 1246 721 1247 725
rect 1251 721 1252 725
rect 1246 720 1252 721
rect 1414 725 1420 726
rect 1414 721 1415 725
rect 1419 721 1420 725
rect 1414 720 1420 721
rect 1582 725 1588 726
rect 1582 721 1583 725
rect 1587 721 1588 725
rect 1582 720 1588 721
rect 1734 725 1740 726
rect 1734 721 1735 725
rect 1739 721 1740 725
rect 1734 720 1740 721
rect 1824 713 1826 737
rect 1864 717 1866 741
rect 1896 730 1898 741
rect 2064 730 2066 741
rect 2256 730 2258 741
rect 2448 730 2450 741
rect 2640 730 2642 741
rect 2824 730 2826 741
rect 3000 730 3002 741
rect 3168 730 3170 741
rect 3336 730 3338 741
rect 3488 730 3490 741
rect 1894 729 1900 730
rect 1894 725 1895 729
rect 1899 725 1900 729
rect 1894 724 1900 725
rect 2062 729 2068 730
rect 2062 725 2063 729
rect 2067 725 2068 729
rect 2062 724 2068 725
rect 2254 729 2260 730
rect 2254 725 2255 729
rect 2259 725 2260 729
rect 2254 724 2260 725
rect 2446 729 2452 730
rect 2446 725 2447 729
rect 2451 725 2452 729
rect 2446 724 2452 725
rect 2638 729 2644 730
rect 2638 725 2639 729
rect 2643 725 2644 729
rect 2638 724 2644 725
rect 2822 729 2828 730
rect 2822 725 2823 729
rect 2827 725 2828 729
rect 2822 724 2828 725
rect 2998 729 3004 730
rect 2998 725 2999 729
rect 3003 725 3004 729
rect 2998 724 3004 725
rect 3166 729 3172 730
rect 3166 725 3167 729
rect 3171 725 3172 729
rect 3166 724 3172 725
rect 3334 729 3340 730
rect 3334 725 3335 729
rect 3339 725 3340 729
rect 3334 724 3340 725
rect 3486 729 3492 730
rect 3486 725 3487 729
rect 3491 725 3492 729
rect 3486 724 3492 725
rect 3576 717 3578 741
rect 1862 716 1868 717
rect 110 712 116 713
rect 110 708 111 712
rect 115 708 116 712
rect 110 707 116 708
rect 1822 712 1828 713
rect 1822 708 1823 712
rect 1827 708 1828 712
rect 1862 712 1863 716
rect 1867 712 1868 716
rect 1862 711 1868 712
rect 3574 716 3580 717
rect 3574 712 3575 716
rect 3579 712 3580 716
rect 3574 711 3580 712
rect 1822 707 1828 708
rect 1862 699 1868 700
rect 110 695 116 696
rect 110 691 111 695
rect 115 691 116 695
rect 110 690 116 691
rect 1822 695 1828 696
rect 1822 691 1823 695
rect 1827 691 1828 695
rect 1862 695 1863 699
rect 1867 695 1868 699
rect 1862 694 1868 695
rect 3574 699 3580 700
rect 3574 695 3575 699
rect 3579 695 3580 699
rect 3574 694 3580 695
rect 1822 690 1828 691
rect 112 675 114 690
rect 206 685 212 686
rect 206 681 207 685
rect 211 681 212 685
rect 206 680 212 681
rect 350 685 356 686
rect 350 681 351 685
rect 355 681 356 685
rect 350 680 356 681
rect 494 685 500 686
rect 494 681 495 685
rect 499 681 500 685
rect 494 680 500 681
rect 638 685 644 686
rect 638 681 639 685
rect 643 681 644 685
rect 638 680 644 681
rect 782 685 788 686
rect 782 681 783 685
rect 787 681 788 685
rect 782 680 788 681
rect 926 685 932 686
rect 926 681 927 685
rect 931 681 932 685
rect 926 680 932 681
rect 1078 685 1084 686
rect 1078 681 1079 685
rect 1083 681 1084 685
rect 1078 680 1084 681
rect 1238 685 1244 686
rect 1238 681 1239 685
rect 1243 681 1244 685
rect 1238 680 1244 681
rect 1406 685 1412 686
rect 1406 681 1407 685
rect 1411 681 1412 685
rect 1406 680 1412 681
rect 1574 685 1580 686
rect 1574 681 1575 685
rect 1579 681 1580 685
rect 1574 680 1580 681
rect 1726 685 1732 686
rect 1726 681 1727 685
rect 1731 681 1732 685
rect 1726 680 1732 681
rect 208 675 210 680
rect 352 675 354 680
rect 496 675 498 680
rect 640 675 642 680
rect 784 675 786 680
rect 928 675 930 680
rect 1080 675 1082 680
rect 1240 675 1242 680
rect 1408 675 1410 680
rect 1576 675 1578 680
rect 1728 675 1730 680
rect 1824 675 1826 690
rect 1864 675 1866 694
rect 1886 689 1892 690
rect 1886 685 1887 689
rect 1891 685 1892 689
rect 1886 684 1892 685
rect 2054 689 2060 690
rect 2054 685 2055 689
rect 2059 685 2060 689
rect 2054 684 2060 685
rect 2246 689 2252 690
rect 2246 685 2247 689
rect 2251 685 2252 689
rect 2246 684 2252 685
rect 2438 689 2444 690
rect 2438 685 2439 689
rect 2443 685 2444 689
rect 2438 684 2444 685
rect 2630 689 2636 690
rect 2630 685 2631 689
rect 2635 685 2636 689
rect 2630 684 2636 685
rect 2814 689 2820 690
rect 2814 685 2815 689
rect 2819 685 2820 689
rect 2814 684 2820 685
rect 2990 689 2996 690
rect 2990 685 2991 689
rect 2995 685 2996 689
rect 2990 684 2996 685
rect 3158 689 3164 690
rect 3158 685 3159 689
rect 3163 685 3164 689
rect 3158 684 3164 685
rect 3326 689 3332 690
rect 3326 685 3327 689
rect 3331 685 3332 689
rect 3326 684 3332 685
rect 3478 689 3484 690
rect 3478 685 3479 689
rect 3483 685 3484 689
rect 3478 684 3484 685
rect 1888 675 1890 684
rect 2056 675 2058 684
rect 2248 675 2250 684
rect 2440 675 2442 684
rect 2632 675 2634 684
rect 2816 675 2818 684
rect 2992 675 2994 684
rect 3160 675 3162 684
rect 3328 675 3330 684
rect 3480 675 3482 684
rect 3576 675 3578 694
rect 111 674 115 675
rect 111 669 115 670
rect 135 674 139 675
rect 135 669 139 670
rect 207 674 211 675
rect 207 669 211 670
rect 295 674 299 675
rect 295 669 299 670
rect 351 674 355 675
rect 351 669 355 670
rect 463 674 467 675
rect 463 669 467 670
rect 495 674 499 675
rect 495 669 499 670
rect 623 674 627 675
rect 623 669 627 670
rect 639 674 643 675
rect 639 669 643 670
rect 775 674 779 675
rect 775 669 779 670
rect 783 674 787 675
rect 783 669 787 670
rect 927 674 931 675
rect 927 669 931 670
rect 1071 674 1075 675
rect 1071 669 1075 670
rect 1079 674 1083 675
rect 1079 669 1083 670
rect 1207 674 1211 675
rect 1207 669 1211 670
rect 1239 674 1243 675
rect 1239 669 1243 670
rect 1343 674 1347 675
rect 1343 669 1347 670
rect 1407 674 1411 675
rect 1407 669 1411 670
rect 1479 674 1483 675
rect 1479 669 1483 670
rect 1575 674 1579 675
rect 1575 669 1579 670
rect 1615 674 1619 675
rect 1615 669 1619 670
rect 1727 674 1731 675
rect 1727 669 1731 670
rect 1823 674 1827 675
rect 1823 669 1827 670
rect 1863 674 1867 675
rect 1863 669 1867 670
rect 1887 674 1891 675
rect 1887 669 1891 670
rect 2055 674 2059 675
rect 2055 669 2059 670
rect 2215 674 2219 675
rect 2215 669 2219 670
rect 2247 674 2251 675
rect 2247 669 2251 670
rect 2359 674 2363 675
rect 2359 669 2363 670
rect 2439 674 2443 675
rect 2439 669 2443 670
rect 2511 674 2515 675
rect 2511 669 2515 670
rect 2631 674 2635 675
rect 2631 669 2635 670
rect 2671 674 2675 675
rect 2671 669 2675 670
rect 2815 674 2819 675
rect 2815 669 2819 670
rect 2831 674 2835 675
rect 2831 669 2835 670
rect 2991 674 2995 675
rect 2991 669 2995 670
rect 3159 674 3163 675
rect 3159 669 3163 670
rect 3327 674 3331 675
rect 3327 669 3331 670
rect 3479 674 3483 675
rect 3479 669 3483 670
rect 3575 674 3579 675
rect 3575 669 3579 670
rect 112 654 114 669
rect 136 664 138 669
rect 296 664 298 669
rect 464 664 466 669
rect 624 664 626 669
rect 776 664 778 669
rect 928 664 930 669
rect 1072 664 1074 669
rect 1208 664 1210 669
rect 1344 664 1346 669
rect 1480 664 1482 669
rect 1616 664 1618 669
rect 1728 664 1730 669
rect 134 663 140 664
rect 134 659 135 663
rect 139 659 140 663
rect 134 658 140 659
rect 294 663 300 664
rect 294 659 295 663
rect 299 659 300 663
rect 294 658 300 659
rect 462 663 468 664
rect 462 659 463 663
rect 467 659 468 663
rect 462 658 468 659
rect 622 663 628 664
rect 622 659 623 663
rect 627 659 628 663
rect 622 658 628 659
rect 774 663 780 664
rect 774 659 775 663
rect 779 659 780 663
rect 774 658 780 659
rect 926 663 932 664
rect 926 659 927 663
rect 931 659 932 663
rect 926 658 932 659
rect 1070 663 1076 664
rect 1070 659 1071 663
rect 1075 659 1076 663
rect 1070 658 1076 659
rect 1206 663 1212 664
rect 1206 659 1207 663
rect 1211 659 1212 663
rect 1206 658 1212 659
rect 1342 663 1348 664
rect 1342 659 1343 663
rect 1347 659 1348 663
rect 1342 658 1348 659
rect 1478 663 1484 664
rect 1478 659 1479 663
rect 1483 659 1484 663
rect 1478 658 1484 659
rect 1614 663 1620 664
rect 1614 659 1615 663
rect 1619 659 1620 663
rect 1614 658 1620 659
rect 1726 663 1732 664
rect 1726 659 1727 663
rect 1731 659 1732 663
rect 1726 658 1732 659
rect 1824 654 1826 669
rect 1864 654 1866 669
rect 2216 664 2218 669
rect 2360 664 2362 669
rect 2512 664 2514 669
rect 2672 664 2674 669
rect 2832 664 2834 669
rect 2992 664 2994 669
rect 3160 664 3162 669
rect 3328 664 3330 669
rect 3480 664 3482 669
rect 2214 663 2220 664
rect 2214 659 2215 663
rect 2219 659 2220 663
rect 2214 658 2220 659
rect 2358 663 2364 664
rect 2358 659 2359 663
rect 2363 659 2364 663
rect 2358 658 2364 659
rect 2510 663 2516 664
rect 2510 659 2511 663
rect 2515 659 2516 663
rect 2510 658 2516 659
rect 2670 663 2676 664
rect 2670 659 2671 663
rect 2675 659 2676 663
rect 2670 658 2676 659
rect 2830 663 2836 664
rect 2830 659 2831 663
rect 2835 659 2836 663
rect 2830 658 2836 659
rect 2990 663 2996 664
rect 2990 659 2991 663
rect 2995 659 2996 663
rect 2990 658 2996 659
rect 3158 663 3164 664
rect 3158 659 3159 663
rect 3163 659 3164 663
rect 3158 658 3164 659
rect 3326 663 3332 664
rect 3326 659 3327 663
rect 3331 659 3332 663
rect 3326 658 3332 659
rect 3478 663 3484 664
rect 3478 659 3479 663
rect 3483 659 3484 663
rect 3478 658 3484 659
rect 3576 654 3578 669
rect 110 653 116 654
rect 110 649 111 653
rect 115 649 116 653
rect 110 648 116 649
rect 1822 653 1828 654
rect 1822 649 1823 653
rect 1827 649 1828 653
rect 1822 648 1828 649
rect 1862 653 1868 654
rect 1862 649 1863 653
rect 1867 649 1868 653
rect 1862 648 1868 649
rect 3574 653 3580 654
rect 3574 649 3575 653
rect 3579 649 3580 653
rect 3574 648 3580 649
rect 110 636 116 637
rect 110 632 111 636
rect 115 632 116 636
rect 110 631 116 632
rect 1822 636 1828 637
rect 1822 632 1823 636
rect 1827 632 1828 636
rect 1822 631 1828 632
rect 1862 636 1868 637
rect 1862 632 1863 636
rect 1867 632 1868 636
rect 1862 631 1868 632
rect 3574 636 3580 637
rect 3574 632 3575 636
rect 3579 632 3580 636
rect 3574 631 3580 632
rect 112 603 114 631
rect 142 623 148 624
rect 142 619 143 623
rect 147 619 148 623
rect 142 618 148 619
rect 302 623 308 624
rect 302 619 303 623
rect 307 619 308 623
rect 302 618 308 619
rect 470 623 476 624
rect 470 619 471 623
rect 475 619 476 623
rect 470 618 476 619
rect 630 623 636 624
rect 630 619 631 623
rect 635 619 636 623
rect 630 618 636 619
rect 782 623 788 624
rect 782 619 783 623
rect 787 619 788 623
rect 782 618 788 619
rect 934 623 940 624
rect 934 619 935 623
rect 939 619 940 623
rect 934 618 940 619
rect 1078 623 1084 624
rect 1078 619 1079 623
rect 1083 619 1084 623
rect 1078 618 1084 619
rect 1214 623 1220 624
rect 1214 619 1215 623
rect 1219 619 1220 623
rect 1214 618 1220 619
rect 1350 623 1356 624
rect 1350 619 1351 623
rect 1355 619 1356 623
rect 1350 618 1356 619
rect 1486 623 1492 624
rect 1486 619 1487 623
rect 1491 619 1492 623
rect 1486 618 1492 619
rect 1622 623 1628 624
rect 1622 619 1623 623
rect 1627 619 1628 623
rect 1622 618 1628 619
rect 1734 623 1740 624
rect 1734 619 1735 623
rect 1739 619 1740 623
rect 1734 618 1740 619
rect 144 603 146 618
rect 304 603 306 618
rect 472 603 474 618
rect 632 603 634 618
rect 784 603 786 618
rect 936 603 938 618
rect 1080 603 1082 618
rect 1216 603 1218 618
rect 1352 603 1354 618
rect 1488 603 1490 618
rect 1624 603 1626 618
rect 1736 603 1738 618
rect 1824 603 1826 631
rect 1864 603 1866 631
rect 2222 623 2228 624
rect 2222 619 2223 623
rect 2227 619 2228 623
rect 2222 618 2228 619
rect 2366 623 2372 624
rect 2366 619 2367 623
rect 2371 619 2372 623
rect 2366 618 2372 619
rect 2518 623 2524 624
rect 2518 619 2519 623
rect 2523 619 2524 623
rect 2518 618 2524 619
rect 2678 623 2684 624
rect 2678 619 2679 623
rect 2683 619 2684 623
rect 2678 618 2684 619
rect 2838 623 2844 624
rect 2838 619 2839 623
rect 2843 619 2844 623
rect 2838 618 2844 619
rect 2998 623 3004 624
rect 2998 619 2999 623
rect 3003 619 3004 623
rect 2998 618 3004 619
rect 3166 623 3172 624
rect 3166 619 3167 623
rect 3171 619 3172 623
rect 3166 618 3172 619
rect 3334 623 3340 624
rect 3334 619 3335 623
rect 3339 619 3340 623
rect 3334 618 3340 619
rect 3486 623 3492 624
rect 3486 619 3487 623
rect 3491 619 3492 623
rect 3486 618 3492 619
rect 2224 603 2226 618
rect 2368 603 2370 618
rect 2520 603 2522 618
rect 2680 603 2682 618
rect 2840 603 2842 618
rect 3000 603 3002 618
rect 3168 603 3170 618
rect 3336 603 3338 618
rect 3488 603 3490 618
rect 3576 603 3578 631
rect 111 602 115 603
rect 111 597 115 598
rect 143 602 147 603
rect 143 597 147 598
rect 303 602 307 603
rect 303 597 307 598
rect 471 602 475 603
rect 471 597 475 598
rect 487 602 491 603
rect 487 597 491 598
rect 631 602 635 603
rect 631 597 635 598
rect 671 602 675 603
rect 671 597 675 598
rect 783 602 787 603
rect 783 597 787 598
rect 847 602 851 603
rect 847 597 851 598
rect 935 602 939 603
rect 935 597 939 598
rect 1023 602 1027 603
rect 1023 597 1027 598
rect 1079 602 1083 603
rect 1079 597 1083 598
rect 1199 602 1203 603
rect 1199 597 1203 598
rect 1215 602 1219 603
rect 1215 597 1219 598
rect 1351 602 1355 603
rect 1351 597 1355 598
rect 1375 602 1379 603
rect 1375 597 1379 598
rect 1487 602 1491 603
rect 1487 597 1491 598
rect 1559 602 1563 603
rect 1559 597 1563 598
rect 1623 602 1627 603
rect 1623 597 1627 598
rect 1735 602 1739 603
rect 1735 597 1739 598
rect 1823 602 1827 603
rect 1823 597 1827 598
rect 1863 602 1867 603
rect 1863 597 1867 598
rect 2199 602 2203 603
rect 2199 597 2203 598
rect 2223 602 2227 603
rect 2223 597 2227 598
rect 2287 602 2291 603
rect 2287 597 2291 598
rect 2367 602 2371 603
rect 2367 597 2371 598
rect 2375 602 2379 603
rect 2375 597 2379 598
rect 2463 602 2467 603
rect 2463 597 2467 598
rect 2519 602 2523 603
rect 2519 597 2523 598
rect 2567 602 2571 603
rect 2567 597 2571 598
rect 2679 602 2683 603
rect 2679 597 2683 598
rect 2815 602 2819 603
rect 2815 597 2819 598
rect 2839 602 2843 603
rect 2839 597 2843 598
rect 2975 602 2979 603
rect 2975 597 2979 598
rect 2999 602 3003 603
rect 2999 597 3003 598
rect 3143 602 3147 603
rect 3143 597 3147 598
rect 3167 602 3171 603
rect 3167 597 3171 598
rect 3327 602 3331 603
rect 3327 597 3331 598
rect 3335 602 3339 603
rect 3335 597 3339 598
rect 3487 602 3491 603
rect 3487 597 3491 598
rect 3575 602 3579 603
rect 3575 597 3579 598
rect 112 573 114 597
rect 144 586 146 597
rect 304 586 306 597
rect 488 586 490 597
rect 672 586 674 597
rect 848 586 850 597
rect 1024 586 1026 597
rect 1200 586 1202 597
rect 1376 586 1378 597
rect 1560 586 1562 597
rect 1736 586 1738 597
rect 142 585 148 586
rect 142 581 143 585
rect 147 581 148 585
rect 142 580 148 581
rect 302 585 308 586
rect 302 581 303 585
rect 307 581 308 585
rect 302 580 308 581
rect 486 585 492 586
rect 486 581 487 585
rect 491 581 492 585
rect 486 580 492 581
rect 670 585 676 586
rect 670 581 671 585
rect 675 581 676 585
rect 670 580 676 581
rect 846 585 852 586
rect 846 581 847 585
rect 851 581 852 585
rect 846 580 852 581
rect 1022 585 1028 586
rect 1022 581 1023 585
rect 1027 581 1028 585
rect 1022 580 1028 581
rect 1198 585 1204 586
rect 1198 581 1199 585
rect 1203 581 1204 585
rect 1198 580 1204 581
rect 1374 585 1380 586
rect 1374 581 1375 585
rect 1379 581 1380 585
rect 1374 580 1380 581
rect 1558 585 1564 586
rect 1558 581 1559 585
rect 1563 581 1564 585
rect 1558 580 1564 581
rect 1734 585 1740 586
rect 1734 581 1735 585
rect 1739 581 1740 585
rect 1734 580 1740 581
rect 1824 573 1826 597
rect 1864 573 1866 597
rect 2200 586 2202 597
rect 2288 586 2290 597
rect 2376 586 2378 597
rect 2464 586 2466 597
rect 2568 586 2570 597
rect 2680 586 2682 597
rect 2816 586 2818 597
rect 2976 586 2978 597
rect 3144 586 3146 597
rect 3328 586 3330 597
rect 3488 586 3490 597
rect 2198 585 2204 586
rect 2198 581 2199 585
rect 2203 581 2204 585
rect 2198 580 2204 581
rect 2286 585 2292 586
rect 2286 581 2287 585
rect 2291 581 2292 585
rect 2286 580 2292 581
rect 2374 585 2380 586
rect 2374 581 2375 585
rect 2379 581 2380 585
rect 2374 580 2380 581
rect 2462 585 2468 586
rect 2462 581 2463 585
rect 2467 581 2468 585
rect 2462 580 2468 581
rect 2566 585 2572 586
rect 2566 581 2567 585
rect 2571 581 2572 585
rect 2566 580 2572 581
rect 2678 585 2684 586
rect 2678 581 2679 585
rect 2683 581 2684 585
rect 2678 580 2684 581
rect 2814 585 2820 586
rect 2814 581 2815 585
rect 2819 581 2820 585
rect 2814 580 2820 581
rect 2974 585 2980 586
rect 2974 581 2975 585
rect 2979 581 2980 585
rect 2974 580 2980 581
rect 3142 585 3148 586
rect 3142 581 3143 585
rect 3147 581 3148 585
rect 3142 580 3148 581
rect 3326 585 3332 586
rect 3326 581 3327 585
rect 3331 581 3332 585
rect 3326 580 3332 581
rect 3486 585 3492 586
rect 3486 581 3487 585
rect 3491 581 3492 585
rect 3486 580 3492 581
rect 3576 573 3578 597
rect 110 572 116 573
rect 110 568 111 572
rect 115 568 116 572
rect 110 567 116 568
rect 1822 572 1828 573
rect 1822 568 1823 572
rect 1827 568 1828 572
rect 1822 567 1828 568
rect 1862 572 1868 573
rect 1862 568 1863 572
rect 1867 568 1868 572
rect 1862 567 1868 568
rect 3574 572 3580 573
rect 3574 568 3575 572
rect 3579 568 3580 572
rect 3574 567 3580 568
rect 110 555 116 556
rect 110 551 111 555
rect 115 551 116 555
rect 110 550 116 551
rect 1822 555 1828 556
rect 1822 551 1823 555
rect 1827 551 1828 555
rect 1822 550 1828 551
rect 1862 555 1868 556
rect 1862 551 1863 555
rect 1867 551 1868 555
rect 1862 550 1868 551
rect 3574 555 3580 556
rect 3574 551 3575 555
rect 3579 551 3580 555
rect 3574 550 3580 551
rect 112 531 114 550
rect 134 545 140 546
rect 134 541 135 545
rect 139 541 140 545
rect 134 540 140 541
rect 294 545 300 546
rect 294 541 295 545
rect 299 541 300 545
rect 294 540 300 541
rect 478 545 484 546
rect 478 541 479 545
rect 483 541 484 545
rect 478 540 484 541
rect 662 545 668 546
rect 662 541 663 545
rect 667 541 668 545
rect 662 540 668 541
rect 838 545 844 546
rect 838 541 839 545
rect 843 541 844 545
rect 838 540 844 541
rect 1014 545 1020 546
rect 1014 541 1015 545
rect 1019 541 1020 545
rect 1014 540 1020 541
rect 1190 545 1196 546
rect 1190 541 1191 545
rect 1195 541 1196 545
rect 1190 540 1196 541
rect 1366 545 1372 546
rect 1366 541 1367 545
rect 1371 541 1372 545
rect 1366 540 1372 541
rect 1550 545 1556 546
rect 1550 541 1551 545
rect 1555 541 1556 545
rect 1550 540 1556 541
rect 1726 545 1732 546
rect 1726 541 1727 545
rect 1731 541 1732 545
rect 1726 540 1732 541
rect 136 531 138 540
rect 296 531 298 540
rect 480 531 482 540
rect 664 531 666 540
rect 840 531 842 540
rect 1016 531 1018 540
rect 1192 531 1194 540
rect 1368 531 1370 540
rect 1552 531 1554 540
rect 1728 531 1730 540
rect 1824 531 1826 550
rect 1864 531 1866 550
rect 2190 545 2196 546
rect 2190 541 2191 545
rect 2195 541 2196 545
rect 2190 540 2196 541
rect 2278 545 2284 546
rect 2278 541 2279 545
rect 2283 541 2284 545
rect 2278 540 2284 541
rect 2366 545 2372 546
rect 2366 541 2367 545
rect 2371 541 2372 545
rect 2366 540 2372 541
rect 2454 545 2460 546
rect 2454 541 2455 545
rect 2459 541 2460 545
rect 2454 540 2460 541
rect 2558 545 2564 546
rect 2558 541 2559 545
rect 2563 541 2564 545
rect 2558 540 2564 541
rect 2670 545 2676 546
rect 2670 541 2671 545
rect 2675 541 2676 545
rect 2670 540 2676 541
rect 2806 545 2812 546
rect 2806 541 2807 545
rect 2811 541 2812 545
rect 2806 540 2812 541
rect 2966 545 2972 546
rect 2966 541 2967 545
rect 2971 541 2972 545
rect 2966 540 2972 541
rect 3134 545 3140 546
rect 3134 541 3135 545
rect 3139 541 3140 545
rect 3134 540 3140 541
rect 3318 545 3324 546
rect 3318 541 3319 545
rect 3323 541 3324 545
rect 3318 540 3324 541
rect 3478 545 3484 546
rect 3478 541 3479 545
rect 3483 541 3484 545
rect 3478 540 3484 541
rect 2192 531 2194 540
rect 2280 531 2282 540
rect 2368 531 2370 540
rect 2456 531 2458 540
rect 2560 531 2562 540
rect 2672 531 2674 540
rect 2808 531 2810 540
rect 2968 531 2970 540
rect 3136 531 3138 540
rect 3320 531 3322 540
rect 3480 531 3482 540
rect 3576 531 3578 550
rect 111 530 115 531
rect 111 525 115 526
rect 135 530 139 531
rect 135 525 139 526
rect 295 530 299 531
rect 295 525 299 526
rect 303 530 307 531
rect 303 525 307 526
rect 479 530 483 531
rect 479 525 483 526
rect 495 530 499 531
rect 495 525 499 526
rect 663 530 667 531
rect 663 525 667 526
rect 679 530 683 531
rect 679 525 683 526
rect 839 530 843 531
rect 839 525 843 526
rect 863 530 867 531
rect 863 525 867 526
rect 1015 530 1019 531
rect 1015 525 1019 526
rect 1031 530 1035 531
rect 1031 525 1035 526
rect 1191 530 1195 531
rect 1191 525 1195 526
rect 1351 530 1355 531
rect 1351 525 1355 526
rect 1367 530 1371 531
rect 1367 525 1371 526
rect 1503 530 1507 531
rect 1503 525 1507 526
rect 1551 530 1555 531
rect 1551 525 1555 526
rect 1663 530 1667 531
rect 1663 525 1667 526
rect 1727 530 1731 531
rect 1727 525 1731 526
rect 1823 530 1827 531
rect 1823 525 1827 526
rect 1863 530 1867 531
rect 1863 525 1867 526
rect 2191 530 2195 531
rect 2191 525 2195 526
rect 2279 530 2283 531
rect 2279 525 2283 526
rect 2303 530 2307 531
rect 2303 525 2307 526
rect 2367 530 2371 531
rect 2367 525 2371 526
rect 2399 530 2403 531
rect 2399 525 2403 526
rect 2455 530 2459 531
rect 2455 525 2459 526
rect 2503 530 2507 531
rect 2503 525 2507 526
rect 2559 530 2563 531
rect 2559 525 2563 526
rect 2607 530 2611 531
rect 2607 525 2611 526
rect 2671 530 2675 531
rect 2671 525 2675 526
rect 2719 530 2723 531
rect 2719 525 2723 526
rect 2807 530 2811 531
rect 2807 525 2811 526
rect 2839 530 2843 531
rect 2839 525 2843 526
rect 2967 530 2971 531
rect 2967 525 2971 526
rect 3095 530 3099 531
rect 3095 525 3099 526
rect 3135 530 3139 531
rect 3135 525 3139 526
rect 3223 530 3227 531
rect 3223 525 3227 526
rect 3319 530 3323 531
rect 3319 525 3323 526
rect 3351 530 3355 531
rect 3351 525 3355 526
rect 3479 530 3483 531
rect 3479 525 3483 526
rect 3575 530 3579 531
rect 3575 525 3579 526
rect 112 510 114 525
rect 136 520 138 525
rect 304 520 306 525
rect 496 520 498 525
rect 680 520 682 525
rect 864 520 866 525
rect 1032 520 1034 525
rect 1192 520 1194 525
rect 1352 520 1354 525
rect 1504 520 1506 525
rect 1664 520 1666 525
rect 134 519 140 520
rect 134 515 135 519
rect 139 515 140 519
rect 134 514 140 515
rect 302 519 308 520
rect 302 515 303 519
rect 307 515 308 519
rect 302 514 308 515
rect 494 519 500 520
rect 494 515 495 519
rect 499 515 500 519
rect 494 514 500 515
rect 678 519 684 520
rect 678 515 679 519
rect 683 515 684 519
rect 678 514 684 515
rect 862 519 868 520
rect 862 515 863 519
rect 867 515 868 519
rect 862 514 868 515
rect 1030 519 1036 520
rect 1030 515 1031 519
rect 1035 515 1036 519
rect 1030 514 1036 515
rect 1190 519 1196 520
rect 1190 515 1191 519
rect 1195 515 1196 519
rect 1190 514 1196 515
rect 1350 519 1356 520
rect 1350 515 1351 519
rect 1355 515 1356 519
rect 1350 514 1356 515
rect 1502 519 1508 520
rect 1502 515 1503 519
rect 1507 515 1508 519
rect 1502 514 1508 515
rect 1662 519 1668 520
rect 1662 515 1663 519
rect 1667 515 1668 519
rect 1662 514 1668 515
rect 1824 510 1826 525
rect 1864 510 1866 525
rect 2304 520 2306 525
rect 2400 520 2402 525
rect 2504 520 2506 525
rect 2608 520 2610 525
rect 2720 520 2722 525
rect 2840 520 2842 525
rect 2968 520 2970 525
rect 3096 520 3098 525
rect 3224 520 3226 525
rect 3352 520 3354 525
rect 3480 520 3482 525
rect 2302 519 2308 520
rect 2302 515 2303 519
rect 2307 515 2308 519
rect 2302 514 2308 515
rect 2398 519 2404 520
rect 2398 515 2399 519
rect 2403 515 2404 519
rect 2398 514 2404 515
rect 2502 519 2508 520
rect 2502 515 2503 519
rect 2507 515 2508 519
rect 2502 514 2508 515
rect 2606 519 2612 520
rect 2606 515 2607 519
rect 2611 515 2612 519
rect 2606 514 2612 515
rect 2718 519 2724 520
rect 2718 515 2719 519
rect 2723 515 2724 519
rect 2718 514 2724 515
rect 2838 519 2844 520
rect 2838 515 2839 519
rect 2843 515 2844 519
rect 2838 514 2844 515
rect 2966 519 2972 520
rect 2966 515 2967 519
rect 2971 515 2972 519
rect 2966 514 2972 515
rect 3094 519 3100 520
rect 3094 515 3095 519
rect 3099 515 3100 519
rect 3094 514 3100 515
rect 3222 519 3228 520
rect 3222 515 3223 519
rect 3227 515 3228 519
rect 3222 514 3228 515
rect 3350 519 3356 520
rect 3350 515 3351 519
rect 3355 515 3356 519
rect 3350 514 3356 515
rect 3478 519 3484 520
rect 3478 515 3479 519
rect 3483 515 3484 519
rect 3478 514 3484 515
rect 3576 510 3578 525
rect 110 509 116 510
rect 110 505 111 509
rect 115 505 116 509
rect 110 504 116 505
rect 1822 509 1828 510
rect 1822 505 1823 509
rect 1827 505 1828 509
rect 1822 504 1828 505
rect 1862 509 1868 510
rect 1862 505 1863 509
rect 1867 505 1868 509
rect 1862 504 1868 505
rect 3574 509 3580 510
rect 3574 505 3575 509
rect 3579 505 3580 509
rect 3574 504 3580 505
rect 110 492 116 493
rect 110 488 111 492
rect 115 488 116 492
rect 110 487 116 488
rect 1822 492 1828 493
rect 1822 488 1823 492
rect 1827 488 1828 492
rect 1822 487 1828 488
rect 1862 492 1868 493
rect 1862 488 1863 492
rect 1867 488 1868 492
rect 1862 487 1868 488
rect 3574 492 3580 493
rect 3574 488 3575 492
rect 3579 488 3580 492
rect 3574 487 3580 488
rect 112 459 114 487
rect 142 479 148 480
rect 142 475 143 479
rect 147 475 148 479
rect 142 474 148 475
rect 310 479 316 480
rect 310 475 311 479
rect 315 475 316 479
rect 310 474 316 475
rect 502 479 508 480
rect 502 475 503 479
rect 507 475 508 479
rect 502 474 508 475
rect 686 479 692 480
rect 686 475 687 479
rect 691 475 692 479
rect 686 474 692 475
rect 870 479 876 480
rect 870 475 871 479
rect 875 475 876 479
rect 870 474 876 475
rect 1038 479 1044 480
rect 1038 475 1039 479
rect 1043 475 1044 479
rect 1038 474 1044 475
rect 1198 479 1204 480
rect 1198 475 1199 479
rect 1203 475 1204 479
rect 1198 474 1204 475
rect 1358 479 1364 480
rect 1358 475 1359 479
rect 1363 475 1364 479
rect 1358 474 1364 475
rect 1510 479 1516 480
rect 1510 475 1511 479
rect 1515 475 1516 479
rect 1510 474 1516 475
rect 1670 479 1676 480
rect 1670 475 1671 479
rect 1675 475 1676 479
rect 1670 474 1676 475
rect 144 459 146 474
rect 312 459 314 474
rect 504 459 506 474
rect 688 459 690 474
rect 872 459 874 474
rect 1040 459 1042 474
rect 1200 459 1202 474
rect 1360 459 1362 474
rect 1512 459 1514 474
rect 1672 459 1674 474
rect 1824 459 1826 487
rect 1864 463 1866 487
rect 2310 479 2316 480
rect 2310 475 2311 479
rect 2315 475 2316 479
rect 2310 474 2316 475
rect 2406 479 2412 480
rect 2406 475 2407 479
rect 2411 475 2412 479
rect 2406 474 2412 475
rect 2510 479 2516 480
rect 2510 475 2511 479
rect 2515 475 2516 479
rect 2510 474 2516 475
rect 2614 479 2620 480
rect 2614 475 2615 479
rect 2619 475 2620 479
rect 2614 474 2620 475
rect 2726 479 2732 480
rect 2726 475 2727 479
rect 2731 475 2732 479
rect 2726 474 2732 475
rect 2846 479 2852 480
rect 2846 475 2847 479
rect 2851 475 2852 479
rect 2846 474 2852 475
rect 2974 479 2980 480
rect 2974 475 2975 479
rect 2979 475 2980 479
rect 2974 474 2980 475
rect 3102 479 3108 480
rect 3102 475 3103 479
rect 3107 475 3108 479
rect 3102 474 3108 475
rect 3230 479 3236 480
rect 3230 475 3231 479
rect 3235 475 3236 479
rect 3230 474 3236 475
rect 3358 479 3364 480
rect 3358 475 3359 479
rect 3363 475 3364 479
rect 3358 474 3364 475
rect 3486 479 3492 480
rect 3486 475 3487 479
rect 3491 475 3492 479
rect 3486 474 3492 475
rect 2312 463 2314 474
rect 2408 463 2410 474
rect 2512 463 2514 474
rect 2616 463 2618 474
rect 2728 463 2730 474
rect 2848 463 2850 474
rect 2976 463 2978 474
rect 3104 463 3106 474
rect 3232 463 3234 474
rect 3360 463 3362 474
rect 3488 463 3490 474
rect 3576 463 3578 487
rect 1863 462 1867 463
rect 111 458 115 459
rect 111 453 115 454
rect 143 458 147 459
rect 143 453 147 454
rect 303 458 307 459
rect 303 453 307 454
rect 311 458 315 459
rect 311 453 315 454
rect 495 458 499 459
rect 495 453 499 454
rect 503 458 507 459
rect 503 453 507 454
rect 687 458 691 459
rect 687 453 691 454
rect 871 458 875 459
rect 871 453 875 454
rect 879 458 883 459
rect 879 453 883 454
rect 1039 458 1043 459
rect 1039 453 1043 454
rect 1055 458 1059 459
rect 1055 453 1059 454
rect 1199 458 1203 459
rect 1199 453 1203 454
rect 1223 458 1227 459
rect 1223 453 1227 454
rect 1359 458 1363 459
rect 1359 453 1363 454
rect 1391 458 1395 459
rect 1391 453 1395 454
rect 1511 458 1515 459
rect 1511 453 1515 454
rect 1559 458 1563 459
rect 1559 453 1563 454
rect 1671 458 1675 459
rect 1671 453 1675 454
rect 1727 458 1731 459
rect 1727 453 1731 454
rect 1823 458 1827 459
rect 1863 457 1867 458
rect 2239 462 2243 463
rect 2239 457 2243 458
rect 2311 462 2315 463
rect 2311 457 2315 458
rect 2327 462 2331 463
rect 2327 457 2331 458
rect 2407 462 2411 463
rect 2407 457 2411 458
rect 2431 462 2435 463
rect 2431 457 2435 458
rect 2511 462 2515 463
rect 2511 457 2515 458
rect 2559 462 2563 463
rect 2559 457 2563 458
rect 2615 462 2619 463
rect 2615 457 2619 458
rect 2695 462 2699 463
rect 2695 457 2699 458
rect 2727 462 2731 463
rect 2727 457 2731 458
rect 2847 462 2851 463
rect 2847 457 2851 458
rect 2975 462 2979 463
rect 2975 457 2979 458
rect 2999 462 3003 463
rect 2999 457 3003 458
rect 3103 462 3107 463
rect 3103 457 3107 458
rect 3159 462 3163 463
rect 3159 457 3163 458
rect 3231 462 3235 463
rect 3231 457 3235 458
rect 3327 462 3331 463
rect 3327 457 3331 458
rect 3359 462 3363 463
rect 3359 457 3363 458
rect 3487 462 3491 463
rect 3487 457 3491 458
rect 3575 462 3579 463
rect 3575 457 3579 458
rect 1823 453 1827 454
rect 112 429 114 453
rect 144 442 146 453
rect 304 442 306 453
rect 496 442 498 453
rect 688 442 690 453
rect 880 442 882 453
rect 1056 442 1058 453
rect 1224 442 1226 453
rect 1392 442 1394 453
rect 1560 442 1562 453
rect 1728 442 1730 453
rect 142 441 148 442
rect 142 437 143 441
rect 147 437 148 441
rect 142 436 148 437
rect 302 441 308 442
rect 302 437 303 441
rect 307 437 308 441
rect 302 436 308 437
rect 494 441 500 442
rect 494 437 495 441
rect 499 437 500 441
rect 494 436 500 437
rect 686 441 692 442
rect 686 437 687 441
rect 691 437 692 441
rect 686 436 692 437
rect 878 441 884 442
rect 878 437 879 441
rect 883 437 884 441
rect 878 436 884 437
rect 1054 441 1060 442
rect 1054 437 1055 441
rect 1059 437 1060 441
rect 1054 436 1060 437
rect 1222 441 1228 442
rect 1222 437 1223 441
rect 1227 437 1228 441
rect 1222 436 1228 437
rect 1390 441 1396 442
rect 1390 437 1391 441
rect 1395 437 1396 441
rect 1390 436 1396 437
rect 1558 441 1564 442
rect 1558 437 1559 441
rect 1563 437 1564 441
rect 1558 436 1564 437
rect 1726 441 1732 442
rect 1726 437 1727 441
rect 1731 437 1732 441
rect 1726 436 1732 437
rect 1824 429 1826 453
rect 1864 433 1866 457
rect 2240 446 2242 457
rect 2328 446 2330 457
rect 2432 446 2434 457
rect 2560 446 2562 457
rect 2696 446 2698 457
rect 2848 446 2850 457
rect 3000 446 3002 457
rect 3160 446 3162 457
rect 3328 446 3330 457
rect 3488 446 3490 457
rect 2238 445 2244 446
rect 2238 441 2239 445
rect 2243 441 2244 445
rect 2238 440 2244 441
rect 2326 445 2332 446
rect 2326 441 2327 445
rect 2331 441 2332 445
rect 2326 440 2332 441
rect 2430 445 2436 446
rect 2430 441 2431 445
rect 2435 441 2436 445
rect 2430 440 2436 441
rect 2558 445 2564 446
rect 2558 441 2559 445
rect 2563 441 2564 445
rect 2558 440 2564 441
rect 2694 445 2700 446
rect 2694 441 2695 445
rect 2699 441 2700 445
rect 2694 440 2700 441
rect 2846 445 2852 446
rect 2846 441 2847 445
rect 2851 441 2852 445
rect 2846 440 2852 441
rect 2998 445 3004 446
rect 2998 441 2999 445
rect 3003 441 3004 445
rect 2998 440 3004 441
rect 3158 445 3164 446
rect 3158 441 3159 445
rect 3163 441 3164 445
rect 3158 440 3164 441
rect 3326 445 3332 446
rect 3326 441 3327 445
rect 3331 441 3332 445
rect 3326 440 3332 441
rect 3486 445 3492 446
rect 3486 441 3487 445
rect 3491 441 3492 445
rect 3486 440 3492 441
rect 3576 433 3578 457
rect 1862 432 1868 433
rect 110 428 116 429
rect 110 424 111 428
rect 115 424 116 428
rect 110 423 116 424
rect 1822 428 1828 429
rect 1822 424 1823 428
rect 1827 424 1828 428
rect 1862 428 1863 432
rect 1867 428 1868 432
rect 1862 427 1868 428
rect 3574 432 3580 433
rect 3574 428 3575 432
rect 3579 428 3580 432
rect 3574 427 3580 428
rect 1822 423 1828 424
rect 1862 415 1868 416
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 110 406 116 407
rect 1822 411 1828 412
rect 1822 407 1823 411
rect 1827 407 1828 411
rect 1862 411 1863 415
rect 1867 411 1868 415
rect 1862 410 1868 411
rect 3574 415 3580 416
rect 3574 411 3575 415
rect 3579 411 3580 415
rect 3574 410 3580 411
rect 1822 406 1828 407
rect 112 391 114 406
rect 134 401 140 402
rect 134 397 135 401
rect 139 397 140 401
rect 134 396 140 397
rect 294 401 300 402
rect 294 397 295 401
rect 299 397 300 401
rect 294 396 300 397
rect 486 401 492 402
rect 486 397 487 401
rect 491 397 492 401
rect 486 396 492 397
rect 678 401 684 402
rect 678 397 679 401
rect 683 397 684 401
rect 678 396 684 397
rect 870 401 876 402
rect 870 397 871 401
rect 875 397 876 401
rect 870 396 876 397
rect 1046 401 1052 402
rect 1046 397 1047 401
rect 1051 397 1052 401
rect 1046 396 1052 397
rect 1214 401 1220 402
rect 1214 397 1215 401
rect 1219 397 1220 401
rect 1214 396 1220 397
rect 1382 401 1388 402
rect 1382 397 1383 401
rect 1387 397 1388 401
rect 1382 396 1388 397
rect 1550 401 1556 402
rect 1550 397 1551 401
rect 1555 397 1556 401
rect 1550 396 1556 397
rect 1718 401 1724 402
rect 1718 397 1719 401
rect 1723 397 1724 401
rect 1718 396 1724 397
rect 136 391 138 396
rect 296 391 298 396
rect 488 391 490 396
rect 680 391 682 396
rect 872 391 874 396
rect 1048 391 1050 396
rect 1216 391 1218 396
rect 1384 391 1386 396
rect 1552 391 1554 396
rect 1720 391 1722 396
rect 1824 391 1826 406
rect 1864 395 1866 410
rect 2230 405 2236 406
rect 2230 401 2231 405
rect 2235 401 2236 405
rect 2230 400 2236 401
rect 2318 405 2324 406
rect 2318 401 2319 405
rect 2323 401 2324 405
rect 2318 400 2324 401
rect 2422 405 2428 406
rect 2422 401 2423 405
rect 2427 401 2428 405
rect 2422 400 2428 401
rect 2550 405 2556 406
rect 2550 401 2551 405
rect 2555 401 2556 405
rect 2550 400 2556 401
rect 2686 405 2692 406
rect 2686 401 2687 405
rect 2691 401 2692 405
rect 2686 400 2692 401
rect 2838 405 2844 406
rect 2838 401 2839 405
rect 2843 401 2844 405
rect 2838 400 2844 401
rect 2990 405 2996 406
rect 2990 401 2991 405
rect 2995 401 2996 405
rect 2990 400 2996 401
rect 3150 405 3156 406
rect 3150 401 3151 405
rect 3155 401 3156 405
rect 3150 400 3156 401
rect 3318 405 3324 406
rect 3318 401 3319 405
rect 3323 401 3324 405
rect 3318 400 3324 401
rect 3478 405 3484 406
rect 3478 401 3479 405
rect 3483 401 3484 405
rect 3478 400 3484 401
rect 2232 395 2234 400
rect 2320 395 2322 400
rect 2424 395 2426 400
rect 2552 395 2554 400
rect 2688 395 2690 400
rect 2840 395 2842 400
rect 2992 395 2994 400
rect 3152 395 3154 400
rect 3320 395 3322 400
rect 3480 395 3482 400
rect 3576 395 3578 410
rect 1863 394 1867 395
rect 111 390 115 391
rect 111 385 115 386
rect 135 390 139 391
rect 135 385 139 386
rect 263 390 267 391
rect 263 385 267 386
rect 295 390 299 391
rect 295 385 299 386
rect 423 390 427 391
rect 423 385 427 386
rect 487 390 491 391
rect 487 385 491 386
rect 591 390 595 391
rect 591 385 595 386
rect 679 390 683 391
rect 679 385 683 386
rect 767 390 771 391
rect 767 385 771 386
rect 871 390 875 391
rect 871 385 875 386
rect 935 390 939 391
rect 935 385 939 386
rect 1047 390 1051 391
rect 1047 385 1051 386
rect 1103 390 1107 391
rect 1103 385 1107 386
rect 1215 390 1219 391
rect 1215 385 1219 386
rect 1263 390 1267 391
rect 1263 385 1267 386
rect 1383 390 1387 391
rect 1383 385 1387 386
rect 1423 390 1427 391
rect 1423 385 1427 386
rect 1551 390 1555 391
rect 1551 385 1555 386
rect 1583 390 1587 391
rect 1583 385 1587 386
rect 1719 390 1723 391
rect 1719 385 1723 386
rect 1727 390 1731 391
rect 1727 385 1731 386
rect 1823 390 1827 391
rect 1863 389 1867 390
rect 2183 394 2187 395
rect 2183 389 2187 390
rect 2231 394 2235 395
rect 2231 389 2235 390
rect 2287 394 2291 395
rect 2287 389 2291 390
rect 2319 394 2323 395
rect 2319 389 2323 390
rect 2399 394 2403 395
rect 2399 389 2403 390
rect 2423 394 2427 395
rect 2423 389 2427 390
rect 2527 394 2531 395
rect 2527 389 2531 390
rect 2551 394 2555 395
rect 2551 389 2555 390
rect 2671 394 2675 395
rect 2671 389 2675 390
rect 2687 394 2691 395
rect 2687 389 2691 390
rect 2815 394 2819 395
rect 2815 389 2819 390
rect 2839 394 2843 395
rect 2839 389 2843 390
rect 2967 394 2971 395
rect 2967 389 2971 390
rect 2991 394 2995 395
rect 2991 389 2995 390
rect 3127 394 3131 395
rect 3127 389 3131 390
rect 3151 394 3155 395
rect 3151 389 3155 390
rect 3295 394 3299 395
rect 3295 389 3299 390
rect 3319 394 3323 395
rect 3319 389 3323 390
rect 3463 394 3467 395
rect 3463 389 3467 390
rect 3479 394 3483 395
rect 3479 389 3483 390
rect 3575 394 3579 395
rect 3575 389 3579 390
rect 1823 385 1827 386
rect 112 370 114 385
rect 136 380 138 385
rect 264 380 266 385
rect 424 380 426 385
rect 592 380 594 385
rect 768 380 770 385
rect 936 380 938 385
rect 1104 380 1106 385
rect 1264 380 1266 385
rect 1424 380 1426 385
rect 1584 380 1586 385
rect 1728 380 1730 385
rect 134 379 140 380
rect 134 375 135 379
rect 139 375 140 379
rect 134 374 140 375
rect 262 379 268 380
rect 262 375 263 379
rect 267 375 268 379
rect 262 374 268 375
rect 422 379 428 380
rect 422 375 423 379
rect 427 375 428 379
rect 422 374 428 375
rect 590 379 596 380
rect 590 375 591 379
rect 595 375 596 379
rect 590 374 596 375
rect 766 379 772 380
rect 766 375 767 379
rect 771 375 772 379
rect 766 374 772 375
rect 934 379 940 380
rect 934 375 935 379
rect 939 375 940 379
rect 934 374 940 375
rect 1102 379 1108 380
rect 1102 375 1103 379
rect 1107 375 1108 379
rect 1102 374 1108 375
rect 1262 379 1268 380
rect 1262 375 1263 379
rect 1267 375 1268 379
rect 1262 374 1268 375
rect 1422 379 1428 380
rect 1422 375 1423 379
rect 1427 375 1428 379
rect 1422 374 1428 375
rect 1582 379 1588 380
rect 1582 375 1583 379
rect 1587 375 1588 379
rect 1582 374 1588 375
rect 1726 379 1732 380
rect 1726 375 1727 379
rect 1731 375 1732 379
rect 1726 374 1732 375
rect 1824 370 1826 385
rect 1864 374 1866 389
rect 2184 384 2186 389
rect 2288 384 2290 389
rect 2400 384 2402 389
rect 2528 384 2530 389
rect 2672 384 2674 389
rect 2816 384 2818 389
rect 2968 384 2970 389
rect 3128 384 3130 389
rect 3296 384 3298 389
rect 3464 384 3466 389
rect 2182 383 2188 384
rect 2182 379 2183 383
rect 2187 379 2188 383
rect 2182 378 2188 379
rect 2286 383 2292 384
rect 2286 379 2287 383
rect 2291 379 2292 383
rect 2286 378 2292 379
rect 2398 383 2404 384
rect 2398 379 2399 383
rect 2403 379 2404 383
rect 2398 378 2404 379
rect 2526 383 2532 384
rect 2526 379 2527 383
rect 2531 379 2532 383
rect 2526 378 2532 379
rect 2670 383 2676 384
rect 2670 379 2671 383
rect 2675 379 2676 383
rect 2670 378 2676 379
rect 2814 383 2820 384
rect 2814 379 2815 383
rect 2819 379 2820 383
rect 2814 378 2820 379
rect 2966 383 2972 384
rect 2966 379 2967 383
rect 2971 379 2972 383
rect 2966 378 2972 379
rect 3126 383 3132 384
rect 3126 379 3127 383
rect 3131 379 3132 383
rect 3126 378 3132 379
rect 3294 383 3300 384
rect 3294 379 3295 383
rect 3299 379 3300 383
rect 3294 378 3300 379
rect 3462 383 3468 384
rect 3462 379 3463 383
rect 3467 379 3468 383
rect 3462 378 3468 379
rect 3576 374 3578 389
rect 1862 373 1868 374
rect 110 369 116 370
rect 110 365 111 369
rect 115 365 116 369
rect 110 364 116 365
rect 1822 369 1828 370
rect 1822 365 1823 369
rect 1827 365 1828 369
rect 1862 369 1863 373
rect 1867 369 1868 373
rect 1862 368 1868 369
rect 3574 373 3580 374
rect 3574 369 3575 373
rect 3579 369 3580 373
rect 3574 368 3580 369
rect 1822 364 1828 365
rect 1862 356 1868 357
rect 110 352 116 353
rect 110 348 111 352
rect 115 348 116 352
rect 110 347 116 348
rect 1822 352 1828 353
rect 1822 348 1823 352
rect 1827 348 1828 352
rect 1862 352 1863 356
rect 1867 352 1868 356
rect 1862 351 1868 352
rect 3574 356 3580 357
rect 3574 352 3575 356
rect 3579 352 3580 356
rect 3574 351 3580 352
rect 1822 347 1828 348
rect 112 323 114 347
rect 142 339 148 340
rect 142 335 143 339
rect 147 335 148 339
rect 142 334 148 335
rect 270 339 276 340
rect 270 335 271 339
rect 275 335 276 339
rect 270 334 276 335
rect 430 339 436 340
rect 430 335 431 339
rect 435 335 436 339
rect 430 334 436 335
rect 598 339 604 340
rect 598 335 599 339
rect 603 335 604 339
rect 598 334 604 335
rect 774 339 780 340
rect 774 335 775 339
rect 779 335 780 339
rect 774 334 780 335
rect 942 339 948 340
rect 942 335 943 339
rect 947 335 948 339
rect 942 334 948 335
rect 1110 339 1116 340
rect 1110 335 1111 339
rect 1115 335 1116 339
rect 1110 334 1116 335
rect 1270 339 1276 340
rect 1270 335 1271 339
rect 1275 335 1276 339
rect 1270 334 1276 335
rect 1430 339 1436 340
rect 1430 335 1431 339
rect 1435 335 1436 339
rect 1430 334 1436 335
rect 1590 339 1596 340
rect 1590 335 1591 339
rect 1595 335 1596 339
rect 1590 334 1596 335
rect 1734 339 1740 340
rect 1734 335 1735 339
rect 1739 335 1740 339
rect 1734 334 1740 335
rect 144 323 146 334
rect 272 323 274 334
rect 432 323 434 334
rect 600 323 602 334
rect 776 323 778 334
rect 944 323 946 334
rect 1112 323 1114 334
rect 1272 323 1274 334
rect 1432 323 1434 334
rect 1592 323 1594 334
rect 1736 323 1738 334
rect 1824 323 1826 347
rect 111 322 115 323
rect 111 317 115 318
rect 143 322 147 323
rect 143 317 147 318
rect 215 322 219 323
rect 215 317 219 318
rect 271 322 275 323
rect 271 317 275 318
rect 351 322 355 323
rect 351 317 355 318
rect 431 322 435 323
rect 431 317 435 318
rect 495 322 499 323
rect 495 317 499 318
rect 599 322 603 323
rect 599 317 603 318
rect 639 322 643 323
rect 639 317 643 318
rect 775 322 779 323
rect 775 317 779 318
rect 791 322 795 323
rect 791 317 795 318
rect 935 322 939 323
rect 935 317 939 318
rect 943 322 947 323
rect 943 317 947 318
rect 1079 322 1083 323
rect 1079 317 1083 318
rect 1111 322 1115 323
rect 1111 317 1115 318
rect 1223 322 1227 323
rect 1223 317 1227 318
rect 1271 322 1275 323
rect 1271 317 1275 318
rect 1359 322 1363 323
rect 1359 317 1363 318
rect 1431 322 1435 323
rect 1431 317 1435 318
rect 1487 322 1491 323
rect 1487 317 1491 318
rect 1591 322 1595 323
rect 1591 317 1595 318
rect 1623 322 1627 323
rect 1623 317 1627 318
rect 1735 322 1739 323
rect 1735 317 1739 318
rect 1823 322 1827 323
rect 1864 319 1866 351
rect 2190 343 2196 344
rect 2190 339 2191 343
rect 2195 339 2196 343
rect 2190 338 2196 339
rect 2294 343 2300 344
rect 2294 339 2295 343
rect 2299 339 2300 343
rect 2294 338 2300 339
rect 2406 343 2412 344
rect 2406 339 2407 343
rect 2411 339 2412 343
rect 2406 338 2412 339
rect 2534 343 2540 344
rect 2534 339 2535 343
rect 2539 339 2540 343
rect 2534 338 2540 339
rect 2678 343 2684 344
rect 2678 339 2679 343
rect 2683 339 2684 343
rect 2678 338 2684 339
rect 2822 343 2828 344
rect 2822 339 2823 343
rect 2827 339 2828 343
rect 2822 338 2828 339
rect 2974 343 2980 344
rect 2974 339 2975 343
rect 2979 339 2980 343
rect 2974 338 2980 339
rect 3134 343 3140 344
rect 3134 339 3135 343
rect 3139 339 3140 343
rect 3134 338 3140 339
rect 3302 343 3308 344
rect 3302 339 3303 343
rect 3307 339 3308 343
rect 3302 338 3308 339
rect 3470 343 3476 344
rect 3470 339 3471 343
rect 3475 339 3476 343
rect 3470 338 3476 339
rect 2192 319 2194 338
rect 2296 319 2298 338
rect 2408 319 2410 338
rect 2536 319 2538 338
rect 2680 319 2682 338
rect 2824 319 2826 338
rect 2976 319 2978 338
rect 3136 319 3138 338
rect 3304 319 3306 338
rect 3472 319 3474 338
rect 3576 319 3578 351
rect 1823 317 1827 318
rect 1863 318 1867 319
rect 112 293 114 317
rect 216 306 218 317
rect 352 306 354 317
rect 496 306 498 317
rect 640 306 642 317
rect 792 306 794 317
rect 936 306 938 317
rect 1080 306 1082 317
rect 1224 306 1226 317
rect 1360 306 1362 317
rect 1488 306 1490 317
rect 1624 306 1626 317
rect 1736 306 1738 317
rect 214 305 220 306
rect 214 301 215 305
rect 219 301 220 305
rect 214 300 220 301
rect 350 305 356 306
rect 350 301 351 305
rect 355 301 356 305
rect 350 300 356 301
rect 494 305 500 306
rect 494 301 495 305
rect 499 301 500 305
rect 494 300 500 301
rect 638 305 644 306
rect 638 301 639 305
rect 643 301 644 305
rect 638 300 644 301
rect 790 305 796 306
rect 790 301 791 305
rect 795 301 796 305
rect 790 300 796 301
rect 934 305 940 306
rect 934 301 935 305
rect 939 301 940 305
rect 934 300 940 301
rect 1078 305 1084 306
rect 1078 301 1079 305
rect 1083 301 1084 305
rect 1078 300 1084 301
rect 1222 305 1228 306
rect 1222 301 1223 305
rect 1227 301 1228 305
rect 1222 300 1228 301
rect 1358 305 1364 306
rect 1358 301 1359 305
rect 1363 301 1364 305
rect 1358 300 1364 301
rect 1486 305 1492 306
rect 1486 301 1487 305
rect 1491 301 1492 305
rect 1486 300 1492 301
rect 1622 305 1628 306
rect 1622 301 1623 305
rect 1627 301 1628 305
rect 1622 300 1628 301
rect 1734 305 1740 306
rect 1734 301 1735 305
rect 1739 301 1740 305
rect 1734 300 1740 301
rect 1824 293 1826 317
rect 1863 313 1867 314
rect 1895 318 1899 319
rect 1895 313 1899 314
rect 2087 318 2091 319
rect 2087 313 2091 314
rect 2191 318 2195 319
rect 2191 313 2195 314
rect 2295 318 2299 319
rect 2295 313 2299 314
rect 2303 318 2307 319
rect 2303 313 2307 314
rect 2407 318 2411 319
rect 2407 313 2411 314
rect 2511 318 2515 319
rect 2511 313 2515 314
rect 2535 318 2539 319
rect 2535 313 2539 314
rect 2679 318 2683 319
rect 2679 313 2683 314
rect 2711 318 2715 319
rect 2711 313 2715 314
rect 2823 318 2827 319
rect 2823 313 2827 314
rect 2903 318 2907 319
rect 2903 313 2907 314
rect 2975 318 2979 319
rect 2975 313 2979 314
rect 3095 318 3099 319
rect 3095 313 3099 314
rect 3135 318 3139 319
rect 3135 313 3139 314
rect 3295 318 3299 319
rect 3295 313 3299 314
rect 3303 318 3307 319
rect 3303 313 3307 314
rect 3471 318 3475 319
rect 3471 313 3475 314
rect 3487 318 3491 319
rect 3487 313 3491 314
rect 3575 318 3579 319
rect 3575 313 3579 314
rect 110 292 116 293
rect 110 288 111 292
rect 115 288 116 292
rect 110 287 116 288
rect 1822 292 1828 293
rect 1822 288 1823 292
rect 1827 288 1828 292
rect 1864 289 1866 313
rect 1896 302 1898 313
rect 2088 302 2090 313
rect 2304 302 2306 313
rect 2512 302 2514 313
rect 2712 302 2714 313
rect 2904 302 2906 313
rect 3096 302 3098 313
rect 3296 302 3298 313
rect 3488 302 3490 313
rect 1894 301 1900 302
rect 1894 297 1895 301
rect 1899 297 1900 301
rect 1894 296 1900 297
rect 2086 301 2092 302
rect 2086 297 2087 301
rect 2091 297 2092 301
rect 2086 296 2092 297
rect 2302 301 2308 302
rect 2302 297 2303 301
rect 2307 297 2308 301
rect 2302 296 2308 297
rect 2510 301 2516 302
rect 2510 297 2511 301
rect 2515 297 2516 301
rect 2510 296 2516 297
rect 2710 301 2716 302
rect 2710 297 2711 301
rect 2715 297 2716 301
rect 2710 296 2716 297
rect 2902 301 2908 302
rect 2902 297 2903 301
rect 2907 297 2908 301
rect 2902 296 2908 297
rect 3094 301 3100 302
rect 3094 297 3095 301
rect 3099 297 3100 301
rect 3094 296 3100 297
rect 3294 301 3300 302
rect 3294 297 3295 301
rect 3299 297 3300 301
rect 3294 296 3300 297
rect 3486 301 3492 302
rect 3486 297 3487 301
rect 3491 297 3492 301
rect 3486 296 3492 297
rect 3576 289 3578 313
rect 1822 287 1828 288
rect 1862 288 1868 289
rect 1862 284 1863 288
rect 1867 284 1868 288
rect 1862 283 1868 284
rect 3574 288 3580 289
rect 3574 284 3575 288
rect 3579 284 3580 288
rect 3574 283 3580 284
rect 110 275 116 276
rect 110 271 111 275
rect 115 271 116 275
rect 110 270 116 271
rect 1822 275 1828 276
rect 1822 271 1823 275
rect 1827 271 1828 275
rect 1822 270 1828 271
rect 1862 271 1868 272
rect 112 247 114 270
rect 206 265 212 266
rect 206 261 207 265
rect 211 261 212 265
rect 206 260 212 261
rect 342 265 348 266
rect 342 261 343 265
rect 347 261 348 265
rect 342 260 348 261
rect 486 265 492 266
rect 486 261 487 265
rect 491 261 492 265
rect 486 260 492 261
rect 630 265 636 266
rect 630 261 631 265
rect 635 261 636 265
rect 630 260 636 261
rect 782 265 788 266
rect 782 261 783 265
rect 787 261 788 265
rect 782 260 788 261
rect 926 265 932 266
rect 926 261 927 265
rect 931 261 932 265
rect 926 260 932 261
rect 1070 265 1076 266
rect 1070 261 1071 265
rect 1075 261 1076 265
rect 1070 260 1076 261
rect 1214 265 1220 266
rect 1214 261 1215 265
rect 1219 261 1220 265
rect 1214 260 1220 261
rect 1350 265 1356 266
rect 1350 261 1351 265
rect 1355 261 1356 265
rect 1350 260 1356 261
rect 1478 265 1484 266
rect 1478 261 1479 265
rect 1483 261 1484 265
rect 1478 260 1484 261
rect 1614 265 1620 266
rect 1614 261 1615 265
rect 1619 261 1620 265
rect 1614 260 1620 261
rect 1726 265 1732 266
rect 1726 261 1727 265
rect 1731 261 1732 265
rect 1726 260 1732 261
rect 208 247 210 260
rect 344 247 346 260
rect 488 247 490 260
rect 632 247 634 260
rect 784 247 786 260
rect 928 247 930 260
rect 1072 247 1074 260
rect 1216 247 1218 260
rect 1352 247 1354 260
rect 1480 247 1482 260
rect 1616 247 1618 260
rect 1728 247 1730 260
rect 1824 247 1826 270
rect 1862 267 1863 271
rect 1867 267 1868 271
rect 1862 266 1868 267
rect 3574 271 3580 272
rect 3574 267 3575 271
rect 3579 267 3580 271
rect 3574 266 3580 267
rect 1864 251 1866 266
rect 1886 261 1892 262
rect 1886 257 1887 261
rect 1891 257 1892 261
rect 1886 256 1892 257
rect 2078 261 2084 262
rect 2078 257 2079 261
rect 2083 257 2084 261
rect 2078 256 2084 257
rect 2294 261 2300 262
rect 2294 257 2295 261
rect 2299 257 2300 261
rect 2294 256 2300 257
rect 2502 261 2508 262
rect 2502 257 2503 261
rect 2507 257 2508 261
rect 2502 256 2508 257
rect 2702 261 2708 262
rect 2702 257 2703 261
rect 2707 257 2708 261
rect 2702 256 2708 257
rect 2894 261 2900 262
rect 2894 257 2895 261
rect 2899 257 2900 261
rect 2894 256 2900 257
rect 3086 261 3092 262
rect 3086 257 3087 261
rect 3091 257 3092 261
rect 3086 256 3092 257
rect 3286 261 3292 262
rect 3286 257 3287 261
rect 3291 257 3292 261
rect 3286 256 3292 257
rect 3478 261 3484 262
rect 3478 257 3479 261
rect 3483 257 3484 261
rect 3478 256 3484 257
rect 1888 251 1890 256
rect 2080 251 2082 256
rect 2296 251 2298 256
rect 2504 251 2506 256
rect 2704 251 2706 256
rect 2896 251 2898 256
rect 3088 251 3090 256
rect 3288 251 3290 256
rect 3480 251 3482 256
rect 3576 251 3578 266
rect 1863 250 1867 251
rect 111 246 115 247
rect 111 241 115 242
rect 207 246 211 247
rect 207 241 211 242
rect 231 246 235 247
rect 231 241 235 242
rect 343 246 347 247
rect 343 241 347 242
rect 359 246 363 247
rect 359 241 363 242
rect 487 246 491 247
rect 487 241 491 242
rect 623 246 627 247
rect 623 241 627 242
rect 631 246 635 247
rect 631 241 635 242
rect 759 246 763 247
rect 759 241 763 242
rect 783 246 787 247
rect 783 241 787 242
rect 895 246 899 247
rect 895 241 899 242
rect 927 246 931 247
rect 927 241 931 242
rect 1031 246 1035 247
rect 1031 241 1035 242
rect 1071 246 1075 247
rect 1071 241 1075 242
rect 1159 246 1163 247
rect 1159 241 1163 242
rect 1215 246 1219 247
rect 1215 241 1219 242
rect 1295 246 1299 247
rect 1295 241 1299 242
rect 1351 246 1355 247
rect 1351 241 1355 242
rect 1431 246 1435 247
rect 1431 241 1435 242
rect 1479 246 1483 247
rect 1479 241 1483 242
rect 1615 246 1619 247
rect 1615 241 1619 242
rect 1727 246 1731 247
rect 1727 241 1731 242
rect 1823 246 1827 247
rect 1863 245 1867 246
rect 1887 250 1891 251
rect 1887 245 1891 246
rect 1999 250 2003 251
rect 1999 245 2003 246
rect 2079 250 2083 251
rect 2079 245 2083 246
rect 2143 250 2147 251
rect 2143 245 2147 246
rect 2295 250 2299 251
rect 2295 245 2299 246
rect 2455 250 2459 251
rect 2455 245 2459 246
rect 2503 250 2507 251
rect 2503 245 2507 246
rect 2615 250 2619 251
rect 2615 245 2619 246
rect 2703 250 2707 251
rect 2703 245 2707 246
rect 2783 250 2787 251
rect 2783 245 2787 246
rect 2895 250 2899 251
rect 2895 245 2899 246
rect 2951 250 2955 251
rect 2951 245 2955 246
rect 3087 250 3091 251
rect 3087 245 3091 246
rect 3127 250 3131 251
rect 3127 245 3131 246
rect 3287 250 3291 251
rect 3287 245 3291 246
rect 3311 250 3315 251
rect 3311 245 3315 246
rect 3479 250 3483 251
rect 3479 245 3483 246
rect 3575 250 3579 251
rect 3575 245 3579 246
rect 1823 241 1827 242
rect 112 226 114 241
rect 232 236 234 241
rect 360 236 362 241
rect 488 236 490 241
rect 624 236 626 241
rect 760 236 762 241
rect 896 236 898 241
rect 1032 236 1034 241
rect 1160 236 1162 241
rect 1296 236 1298 241
rect 1432 236 1434 241
rect 230 235 236 236
rect 230 231 231 235
rect 235 231 236 235
rect 230 230 236 231
rect 358 235 364 236
rect 358 231 359 235
rect 363 231 364 235
rect 358 230 364 231
rect 486 235 492 236
rect 486 231 487 235
rect 491 231 492 235
rect 486 230 492 231
rect 622 235 628 236
rect 622 231 623 235
rect 627 231 628 235
rect 622 230 628 231
rect 758 235 764 236
rect 758 231 759 235
rect 763 231 764 235
rect 758 230 764 231
rect 894 235 900 236
rect 894 231 895 235
rect 899 231 900 235
rect 894 230 900 231
rect 1030 235 1036 236
rect 1030 231 1031 235
rect 1035 231 1036 235
rect 1030 230 1036 231
rect 1158 235 1164 236
rect 1158 231 1159 235
rect 1163 231 1164 235
rect 1158 230 1164 231
rect 1294 235 1300 236
rect 1294 231 1295 235
rect 1299 231 1300 235
rect 1294 230 1300 231
rect 1430 235 1436 236
rect 1430 231 1431 235
rect 1435 231 1436 235
rect 1430 230 1436 231
rect 1824 226 1826 241
rect 1864 230 1866 245
rect 1888 240 1890 245
rect 2000 240 2002 245
rect 2144 240 2146 245
rect 2296 240 2298 245
rect 2456 240 2458 245
rect 2616 240 2618 245
rect 2784 240 2786 245
rect 2952 240 2954 245
rect 3128 240 3130 245
rect 3312 240 3314 245
rect 3480 240 3482 245
rect 1886 239 1892 240
rect 1886 235 1887 239
rect 1891 235 1892 239
rect 1886 234 1892 235
rect 1998 239 2004 240
rect 1998 235 1999 239
rect 2003 235 2004 239
rect 1998 234 2004 235
rect 2142 239 2148 240
rect 2142 235 2143 239
rect 2147 235 2148 239
rect 2142 234 2148 235
rect 2294 239 2300 240
rect 2294 235 2295 239
rect 2299 235 2300 239
rect 2294 234 2300 235
rect 2454 239 2460 240
rect 2454 235 2455 239
rect 2459 235 2460 239
rect 2454 234 2460 235
rect 2614 239 2620 240
rect 2614 235 2615 239
rect 2619 235 2620 239
rect 2614 234 2620 235
rect 2782 239 2788 240
rect 2782 235 2783 239
rect 2787 235 2788 239
rect 2782 234 2788 235
rect 2950 239 2956 240
rect 2950 235 2951 239
rect 2955 235 2956 239
rect 2950 234 2956 235
rect 3126 239 3132 240
rect 3126 235 3127 239
rect 3131 235 3132 239
rect 3126 234 3132 235
rect 3310 239 3316 240
rect 3310 235 3311 239
rect 3315 235 3316 239
rect 3310 234 3316 235
rect 3478 239 3484 240
rect 3478 235 3479 239
rect 3483 235 3484 239
rect 3478 234 3484 235
rect 3576 230 3578 245
rect 1862 229 1868 230
rect 110 225 116 226
rect 110 221 111 225
rect 115 221 116 225
rect 110 220 116 221
rect 1822 225 1828 226
rect 1822 221 1823 225
rect 1827 221 1828 225
rect 1862 225 1863 229
rect 1867 225 1868 229
rect 1862 224 1868 225
rect 3574 229 3580 230
rect 3574 225 3575 229
rect 3579 225 3580 229
rect 3574 224 3580 225
rect 1822 220 1828 221
rect 1862 212 1868 213
rect 110 208 116 209
rect 110 204 111 208
rect 115 204 116 208
rect 110 203 116 204
rect 1822 208 1828 209
rect 1822 204 1823 208
rect 1827 204 1828 208
rect 1862 208 1863 212
rect 1867 208 1868 212
rect 1862 207 1868 208
rect 3574 212 3580 213
rect 3574 208 3575 212
rect 3579 208 3580 212
rect 3574 207 3580 208
rect 1822 203 1828 204
rect 112 155 114 203
rect 238 195 244 196
rect 238 191 239 195
rect 243 191 244 195
rect 238 190 244 191
rect 366 195 372 196
rect 366 191 367 195
rect 371 191 372 195
rect 366 190 372 191
rect 494 195 500 196
rect 494 191 495 195
rect 499 191 500 195
rect 494 190 500 191
rect 630 195 636 196
rect 630 191 631 195
rect 635 191 636 195
rect 630 190 636 191
rect 766 195 772 196
rect 766 191 767 195
rect 771 191 772 195
rect 766 190 772 191
rect 902 195 908 196
rect 902 191 903 195
rect 907 191 908 195
rect 902 190 908 191
rect 1038 195 1044 196
rect 1038 191 1039 195
rect 1043 191 1044 195
rect 1038 190 1044 191
rect 1166 195 1172 196
rect 1166 191 1167 195
rect 1171 191 1172 195
rect 1166 190 1172 191
rect 1302 195 1308 196
rect 1302 191 1303 195
rect 1307 191 1308 195
rect 1302 190 1308 191
rect 1438 195 1444 196
rect 1438 191 1439 195
rect 1443 191 1444 195
rect 1438 190 1444 191
rect 240 155 242 190
rect 368 155 370 190
rect 496 155 498 190
rect 632 155 634 190
rect 768 155 770 190
rect 904 155 906 190
rect 1040 155 1042 190
rect 1168 155 1170 190
rect 1304 155 1306 190
rect 1440 155 1442 190
rect 1824 155 1826 203
rect 1864 155 1866 207
rect 1894 199 1900 200
rect 1894 195 1895 199
rect 1899 195 1900 199
rect 1894 194 1900 195
rect 2006 199 2012 200
rect 2006 195 2007 199
rect 2011 195 2012 199
rect 2006 194 2012 195
rect 2150 199 2156 200
rect 2150 195 2151 199
rect 2155 195 2156 199
rect 2150 194 2156 195
rect 2302 199 2308 200
rect 2302 195 2303 199
rect 2307 195 2308 199
rect 2302 194 2308 195
rect 2462 199 2468 200
rect 2462 195 2463 199
rect 2467 195 2468 199
rect 2462 194 2468 195
rect 2622 199 2628 200
rect 2622 195 2623 199
rect 2627 195 2628 199
rect 2622 194 2628 195
rect 2790 199 2796 200
rect 2790 195 2791 199
rect 2795 195 2796 199
rect 2790 194 2796 195
rect 2958 199 2964 200
rect 2958 195 2959 199
rect 2963 195 2964 199
rect 2958 194 2964 195
rect 3134 199 3140 200
rect 3134 195 3135 199
rect 3139 195 3140 199
rect 3134 194 3140 195
rect 3318 199 3324 200
rect 3318 195 3319 199
rect 3323 195 3324 199
rect 3318 194 3324 195
rect 3486 199 3492 200
rect 3486 195 3487 199
rect 3491 195 3492 199
rect 3486 194 3492 195
rect 1896 155 1898 194
rect 2008 155 2010 194
rect 2152 155 2154 194
rect 2304 155 2306 194
rect 2464 155 2466 194
rect 2624 155 2626 194
rect 2792 155 2794 194
rect 2960 155 2962 194
rect 3136 155 3138 194
rect 3320 155 3322 194
rect 3488 155 3490 194
rect 3576 155 3578 207
rect 111 154 115 155
rect 111 149 115 150
rect 175 154 179 155
rect 175 149 179 150
rect 239 154 243 155
rect 239 149 243 150
rect 263 154 267 155
rect 263 149 267 150
rect 351 154 355 155
rect 351 149 355 150
rect 367 154 371 155
rect 367 149 371 150
rect 439 154 443 155
rect 439 149 443 150
rect 495 154 499 155
rect 495 149 499 150
rect 527 154 531 155
rect 527 149 531 150
rect 615 154 619 155
rect 615 149 619 150
rect 631 154 635 155
rect 631 149 635 150
rect 703 154 707 155
rect 703 149 707 150
rect 767 154 771 155
rect 767 149 771 150
rect 791 154 795 155
rect 791 149 795 150
rect 879 154 883 155
rect 879 149 883 150
rect 903 154 907 155
rect 903 149 907 150
rect 967 154 971 155
rect 967 149 971 150
rect 1039 154 1043 155
rect 1039 149 1043 150
rect 1055 154 1059 155
rect 1055 149 1059 150
rect 1143 154 1147 155
rect 1143 149 1147 150
rect 1167 154 1171 155
rect 1167 149 1171 150
rect 1231 154 1235 155
rect 1231 149 1235 150
rect 1303 154 1307 155
rect 1303 149 1307 150
rect 1319 154 1323 155
rect 1319 149 1323 150
rect 1407 154 1411 155
rect 1407 149 1411 150
rect 1439 154 1443 155
rect 1439 149 1443 150
rect 1503 154 1507 155
rect 1503 149 1507 150
rect 1823 154 1827 155
rect 1823 149 1827 150
rect 1863 154 1867 155
rect 1863 149 1867 150
rect 1895 154 1899 155
rect 1895 149 1899 150
rect 1983 154 1987 155
rect 1983 149 1987 150
rect 2007 154 2011 155
rect 2007 149 2011 150
rect 2071 154 2075 155
rect 2071 149 2075 150
rect 2151 154 2155 155
rect 2151 149 2155 150
rect 2159 154 2163 155
rect 2159 149 2163 150
rect 2247 154 2251 155
rect 2247 149 2251 150
rect 2303 154 2307 155
rect 2303 149 2307 150
rect 2335 154 2339 155
rect 2335 149 2339 150
rect 2439 154 2443 155
rect 2439 149 2443 150
rect 2463 154 2467 155
rect 2463 149 2467 150
rect 2543 154 2547 155
rect 2543 149 2547 150
rect 2623 154 2627 155
rect 2623 149 2627 150
rect 2647 154 2651 155
rect 2647 149 2651 150
rect 2743 154 2747 155
rect 2743 149 2747 150
rect 2791 154 2795 155
rect 2791 149 2795 150
rect 2839 154 2843 155
rect 2839 149 2843 150
rect 2935 154 2939 155
rect 2935 149 2939 150
rect 2959 154 2963 155
rect 2959 149 2963 150
rect 3031 154 3035 155
rect 3031 149 3035 150
rect 3127 154 3131 155
rect 3127 149 3131 150
rect 3135 154 3139 155
rect 3135 149 3139 150
rect 3223 154 3227 155
rect 3223 149 3227 150
rect 3311 154 3315 155
rect 3311 149 3315 150
rect 3319 154 3323 155
rect 3319 149 3323 150
rect 3399 154 3403 155
rect 3399 149 3403 150
rect 3487 154 3491 155
rect 3487 149 3491 150
rect 3575 154 3579 155
rect 3575 149 3579 150
rect 112 125 114 149
rect 176 138 178 149
rect 264 138 266 149
rect 352 138 354 149
rect 440 138 442 149
rect 528 138 530 149
rect 616 138 618 149
rect 704 138 706 149
rect 792 138 794 149
rect 880 138 882 149
rect 968 138 970 149
rect 1056 138 1058 149
rect 1144 138 1146 149
rect 1232 138 1234 149
rect 1320 138 1322 149
rect 1408 138 1410 149
rect 1504 138 1506 149
rect 174 137 180 138
rect 174 133 175 137
rect 179 133 180 137
rect 174 132 180 133
rect 262 137 268 138
rect 262 133 263 137
rect 267 133 268 137
rect 262 132 268 133
rect 350 137 356 138
rect 350 133 351 137
rect 355 133 356 137
rect 350 132 356 133
rect 438 137 444 138
rect 438 133 439 137
rect 443 133 444 137
rect 438 132 444 133
rect 526 137 532 138
rect 526 133 527 137
rect 531 133 532 137
rect 526 132 532 133
rect 614 137 620 138
rect 614 133 615 137
rect 619 133 620 137
rect 614 132 620 133
rect 702 137 708 138
rect 702 133 703 137
rect 707 133 708 137
rect 702 132 708 133
rect 790 137 796 138
rect 790 133 791 137
rect 795 133 796 137
rect 790 132 796 133
rect 878 137 884 138
rect 878 133 879 137
rect 883 133 884 137
rect 878 132 884 133
rect 966 137 972 138
rect 966 133 967 137
rect 971 133 972 137
rect 966 132 972 133
rect 1054 137 1060 138
rect 1054 133 1055 137
rect 1059 133 1060 137
rect 1054 132 1060 133
rect 1142 137 1148 138
rect 1142 133 1143 137
rect 1147 133 1148 137
rect 1142 132 1148 133
rect 1230 137 1236 138
rect 1230 133 1231 137
rect 1235 133 1236 137
rect 1230 132 1236 133
rect 1318 137 1324 138
rect 1318 133 1319 137
rect 1323 133 1324 137
rect 1318 132 1324 133
rect 1406 137 1412 138
rect 1406 133 1407 137
rect 1411 133 1412 137
rect 1406 132 1412 133
rect 1502 137 1508 138
rect 1502 133 1503 137
rect 1507 133 1508 137
rect 1502 132 1508 133
rect 1824 125 1826 149
rect 1864 125 1866 149
rect 1896 138 1898 149
rect 1984 138 1986 149
rect 2072 138 2074 149
rect 2160 138 2162 149
rect 2248 138 2250 149
rect 2336 138 2338 149
rect 2440 138 2442 149
rect 2544 138 2546 149
rect 2648 138 2650 149
rect 2744 138 2746 149
rect 2840 138 2842 149
rect 2936 138 2938 149
rect 3032 138 3034 149
rect 3128 138 3130 149
rect 3224 138 3226 149
rect 3312 138 3314 149
rect 3400 138 3402 149
rect 3488 138 3490 149
rect 1894 137 1900 138
rect 1894 133 1895 137
rect 1899 133 1900 137
rect 1894 132 1900 133
rect 1982 137 1988 138
rect 1982 133 1983 137
rect 1987 133 1988 137
rect 1982 132 1988 133
rect 2070 137 2076 138
rect 2070 133 2071 137
rect 2075 133 2076 137
rect 2070 132 2076 133
rect 2158 137 2164 138
rect 2158 133 2159 137
rect 2163 133 2164 137
rect 2158 132 2164 133
rect 2246 137 2252 138
rect 2246 133 2247 137
rect 2251 133 2252 137
rect 2246 132 2252 133
rect 2334 137 2340 138
rect 2334 133 2335 137
rect 2339 133 2340 137
rect 2334 132 2340 133
rect 2438 137 2444 138
rect 2438 133 2439 137
rect 2443 133 2444 137
rect 2438 132 2444 133
rect 2542 137 2548 138
rect 2542 133 2543 137
rect 2547 133 2548 137
rect 2542 132 2548 133
rect 2646 137 2652 138
rect 2646 133 2647 137
rect 2651 133 2652 137
rect 2646 132 2652 133
rect 2742 137 2748 138
rect 2742 133 2743 137
rect 2747 133 2748 137
rect 2742 132 2748 133
rect 2838 137 2844 138
rect 2838 133 2839 137
rect 2843 133 2844 137
rect 2838 132 2844 133
rect 2934 137 2940 138
rect 2934 133 2935 137
rect 2939 133 2940 137
rect 2934 132 2940 133
rect 3030 137 3036 138
rect 3030 133 3031 137
rect 3035 133 3036 137
rect 3030 132 3036 133
rect 3126 137 3132 138
rect 3126 133 3127 137
rect 3131 133 3132 137
rect 3126 132 3132 133
rect 3222 137 3228 138
rect 3222 133 3223 137
rect 3227 133 3228 137
rect 3222 132 3228 133
rect 3310 137 3316 138
rect 3310 133 3311 137
rect 3315 133 3316 137
rect 3310 132 3316 133
rect 3398 137 3404 138
rect 3398 133 3399 137
rect 3403 133 3404 137
rect 3398 132 3404 133
rect 3486 137 3492 138
rect 3486 133 3487 137
rect 3491 133 3492 137
rect 3486 132 3492 133
rect 3576 125 3578 149
rect 110 124 116 125
rect 110 120 111 124
rect 115 120 116 124
rect 110 119 116 120
rect 1822 124 1828 125
rect 1822 120 1823 124
rect 1827 120 1828 124
rect 1822 119 1828 120
rect 1862 124 1868 125
rect 1862 120 1863 124
rect 1867 120 1868 124
rect 1862 119 1868 120
rect 3574 124 3580 125
rect 3574 120 3575 124
rect 3579 120 3580 124
rect 3574 119 3580 120
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 110 102 116 103
rect 1822 107 1828 108
rect 1822 103 1823 107
rect 1827 103 1828 107
rect 1822 102 1828 103
rect 1862 107 1868 108
rect 1862 103 1863 107
rect 1867 103 1868 107
rect 1862 102 1868 103
rect 3574 107 3580 108
rect 3574 103 3575 107
rect 3579 103 3580 107
rect 3574 102 3580 103
rect 112 87 114 102
rect 166 97 172 98
rect 166 93 167 97
rect 171 93 172 97
rect 166 92 172 93
rect 254 97 260 98
rect 254 93 255 97
rect 259 93 260 97
rect 254 92 260 93
rect 342 97 348 98
rect 342 93 343 97
rect 347 93 348 97
rect 342 92 348 93
rect 430 97 436 98
rect 430 93 431 97
rect 435 93 436 97
rect 430 92 436 93
rect 518 97 524 98
rect 518 93 519 97
rect 523 93 524 97
rect 518 92 524 93
rect 606 97 612 98
rect 606 93 607 97
rect 611 93 612 97
rect 606 92 612 93
rect 694 97 700 98
rect 694 93 695 97
rect 699 93 700 97
rect 694 92 700 93
rect 782 97 788 98
rect 782 93 783 97
rect 787 93 788 97
rect 782 92 788 93
rect 870 97 876 98
rect 870 93 871 97
rect 875 93 876 97
rect 870 92 876 93
rect 958 97 964 98
rect 958 93 959 97
rect 963 93 964 97
rect 958 92 964 93
rect 1046 97 1052 98
rect 1046 93 1047 97
rect 1051 93 1052 97
rect 1046 92 1052 93
rect 1134 97 1140 98
rect 1134 93 1135 97
rect 1139 93 1140 97
rect 1134 92 1140 93
rect 1222 97 1228 98
rect 1222 93 1223 97
rect 1227 93 1228 97
rect 1222 92 1228 93
rect 1310 97 1316 98
rect 1310 93 1311 97
rect 1315 93 1316 97
rect 1310 92 1316 93
rect 1398 97 1404 98
rect 1398 93 1399 97
rect 1403 93 1404 97
rect 1398 92 1404 93
rect 1494 97 1500 98
rect 1494 93 1495 97
rect 1499 93 1500 97
rect 1494 92 1500 93
rect 168 87 170 92
rect 256 87 258 92
rect 344 87 346 92
rect 432 87 434 92
rect 520 87 522 92
rect 608 87 610 92
rect 696 87 698 92
rect 784 87 786 92
rect 872 87 874 92
rect 960 87 962 92
rect 1048 87 1050 92
rect 1136 87 1138 92
rect 1224 87 1226 92
rect 1312 87 1314 92
rect 1400 87 1402 92
rect 1496 87 1498 92
rect 1824 87 1826 102
rect 1864 87 1866 102
rect 1886 97 1892 98
rect 1886 93 1887 97
rect 1891 93 1892 97
rect 1886 92 1892 93
rect 1974 97 1980 98
rect 1974 93 1975 97
rect 1979 93 1980 97
rect 1974 92 1980 93
rect 2062 97 2068 98
rect 2062 93 2063 97
rect 2067 93 2068 97
rect 2062 92 2068 93
rect 2150 97 2156 98
rect 2150 93 2151 97
rect 2155 93 2156 97
rect 2150 92 2156 93
rect 2238 97 2244 98
rect 2238 93 2239 97
rect 2243 93 2244 97
rect 2238 92 2244 93
rect 2326 97 2332 98
rect 2326 93 2327 97
rect 2331 93 2332 97
rect 2326 92 2332 93
rect 2430 97 2436 98
rect 2430 93 2431 97
rect 2435 93 2436 97
rect 2430 92 2436 93
rect 2534 97 2540 98
rect 2534 93 2535 97
rect 2539 93 2540 97
rect 2534 92 2540 93
rect 2638 97 2644 98
rect 2638 93 2639 97
rect 2643 93 2644 97
rect 2638 92 2644 93
rect 2734 97 2740 98
rect 2734 93 2735 97
rect 2739 93 2740 97
rect 2734 92 2740 93
rect 2830 97 2836 98
rect 2830 93 2831 97
rect 2835 93 2836 97
rect 2830 92 2836 93
rect 2926 97 2932 98
rect 2926 93 2927 97
rect 2931 93 2932 97
rect 2926 92 2932 93
rect 3022 97 3028 98
rect 3022 93 3023 97
rect 3027 93 3028 97
rect 3022 92 3028 93
rect 3118 97 3124 98
rect 3118 93 3119 97
rect 3123 93 3124 97
rect 3118 92 3124 93
rect 3214 97 3220 98
rect 3214 93 3215 97
rect 3219 93 3220 97
rect 3214 92 3220 93
rect 3302 97 3308 98
rect 3302 93 3303 97
rect 3307 93 3308 97
rect 3302 92 3308 93
rect 3390 97 3396 98
rect 3390 93 3391 97
rect 3395 93 3396 97
rect 3390 92 3396 93
rect 3478 97 3484 98
rect 3478 93 3479 97
rect 3483 93 3484 97
rect 3478 92 3484 93
rect 1888 87 1890 92
rect 1976 87 1978 92
rect 2064 87 2066 92
rect 2152 87 2154 92
rect 2240 87 2242 92
rect 2328 87 2330 92
rect 2432 87 2434 92
rect 2536 87 2538 92
rect 2640 87 2642 92
rect 2736 87 2738 92
rect 2832 87 2834 92
rect 2928 87 2930 92
rect 3024 87 3026 92
rect 3120 87 3122 92
rect 3216 87 3218 92
rect 3304 87 3306 92
rect 3392 87 3394 92
rect 3480 87 3482 92
rect 3576 87 3578 102
rect 111 86 115 87
rect 111 81 115 82
rect 167 86 171 87
rect 167 81 171 82
rect 255 86 259 87
rect 255 81 259 82
rect 343 86 347 87
rect 343 81 347 82
rect 431 86 435 87
rect 431 81 435 82
rect 519 86 523 87
rect 519 81 523 82
rect 607 86 611 87
rect 607 81 611 82
rect 695 86 699 87
rect 695 81 699 82
rect 783 86 787 87
rect 783 81 787 82
rect 871 86 875 87
rect 871 81 875 82
rect 959 86 963 87
rect 959 81 963 82
rect 1047 86 1051 87
rect 1047 81 1051 82
rect 1135 86 1139 87
rect 1135 81 1139 82
rect 1223 86 1227 87
rect 1223 81 1227 82
rect 1311 86 1315 87
rect 1311 81 1315 82
rect 1399 86 1403 87
rect 1399 81 1403 82
rect 1495 86 1499 87
rect 1495 81 1499 82
rect 1823 86 1827 87
rect 1823 81 1827 82
rect 1863 86 1867 87
rect 1863 81 1867 82
rect 1887 86 1891 87
rect 1887 81 1891 82
rect 1975 86 1979 87
rect 1975 81 1979 82
rect 2063 86 2067 87
rect 2063 81 2067 82
rect 2151 86 2155 87
rect 2151 81 2155 82
rect 2239 86 2243 87
rect 2239 81 2243 82
rect 2327 86 2331 87
rect 2327 81 2331 82
rect 2431 86 2435 87
rect 2431 81 2435 82
rect 2535 86 2539 87
rect 2535 81 2539 82
rect 2639 86 2643 87
rect 2639 81 2643 82
rect 2735 86 2739 87
rect 2735 81 2739 82
rect 2831 86 2835 87
rect 2831 81 2835 82
rect 2927 86 2931 87
rect 2927 81 2931 82
rect 3023 86 3027 87
rect 3023 81 3027 82
rect 3119 86 3123 87
rect 3119 81 3123 82
rect 3215 86 3219 87
rect 3215 81 3219 82
rect 3303 86 3307 87
rect 3303 81 3307 82
rect 3391 86 3395 87
rect 3391 81 3395 82
rect 3479 86 3483 87
rect 3479 81 3483 82
rect 3575 86 3579 87
rect 3575 81 3579 82
<< m4c >>
rect 111 3646 115 3650
rect 239 3646 243 3650
rect 327 3646 331 3650
rect 415 3646 419 3650
rect 503 3646 507 3650
rect 591 3646 595 3650
rect 679 3646 683 3650
rect 1823 3646 1827 3650
rect 1863 3582 1867 3586
rect 1887 3582 1891 3586
rect 1975 3582 1979 3586
rect 2063 3582 2067 3586
rect 2151 3582 2155 3586
rect 2239 3582 2243 3586
rect 2327 3582 2331 3586
rect 2415 3582 2419 3586
rect 2503 3582 2507 3586
rect 2591 3582 2595 3586
rect 2679 3582 2683 3586
rect 2767 3582 2771 3586
rect 2855 3582 2859 3586
rect 2943 3582 2947 3586
rect 3031 3582 3035 3586
rect 3119 3582 3123 3586
rect 3207 3582 3211 3586
rect 3295 3582 3299 3586
rect 3575 3582 3579 3586
rect 111 3570 115 3574
rect 231 3570 235 3574
rect 247 3570 251 3574
rect 319 3570 323 3574
rect 399 3570 403 3574
rect 407 3570 411 3574
rect 495 3570 499 3574
rect 543 3570 547 3574
rect 583 3570 587 3574
rect 671 3570 675 3574
rect 687 3570 691 3574
rect 823 3570 827 3574
rect 951 3570 955 3574
rect 1079 3570 1083 3574
rect 1199 3570 1203 3574
rect 1311 3570 1315 3574
rect 1423 3570 1427 3574
rect 1543 3570 1547 3574
rect 1823 3570 1827 3574
rect 111 3502 115 3506
rect 183 3502 187 3506
rect 255 3502 259 3506
rect 351 3502 355 3506
rect 407 3502 411 3506
rect 519 3502 523 3506
rect 551 3502 555 3506
rect 679 3502 683 3506
rect 695 3502 699 3506
rect 831 3502 835 3506
rect 959 3502 963 3506
rect 967 3502 971 3506
rect 1087 3502 1091 3506
rect 1095 3502 1099 3506
rect 1207 3502 1211 3506
rect 1215 3502 1219 3506
rect 1319 3502 1323 3506
rect 1335 3502 1339 3506
rect 1431 3502 1435 3506
rect 1455 3502 1459 3506
rect 1551 3502 1555 3506
rect 1575 3502 1579 3506
rect 1823 3502 1827 3506
rect 1863 3506 1867 3510
rect 1895 3506 1899 3510
rect 1911 3506 1915 3510
rect 1983 3506 1987 3510
rect 2015 3506 2019 3510
rect 2071 3506 2075 3510
rect 2135 3506 2139 3510
rect 2159 3506 2163 3510
rect 2247 3506 2251 3510
rect 2263 3506 2267 3510
rect 2335 3506 2339 3510
rect 2391 3506 2395 3510
rect 2423 3506 2427 3510
rect 2511 3506 2515 3510
rect 2527 3506 2531 3510
rect 2599 3506 2603 3510
rect 2663 3506 2667 3510
rect 2687 3506 2691 3510
rect 2775 3506 2779 3510
rect 2799 3506 2803 3510
rect 2863 3506 2867 3510
rect 2943 3506 2947 3510
rect 2951 3506 2955 3510
rect 3039 3506 3043 3510
rect 3087 3506 3091 3510
rect 3127 3506 3131 3510
rect 3215 3506 3219 3510
rect 3303 3506 3307 3510
rect 3575 3506 3579 3510
rect 111 3434 115 3438
rect 135 3434 139 3438
rect 175 3434 179 3438
rect 255 3434 259 3438
rect 343 3434 347 3438
rect 415 3434 419 3438
rect 511 3434 515 3438
rect 583 3434 587 3438
rect 671 3434 675 3438
rect 759 3434 763 3438
rect 823 3434 827 3438
rect 935 3434 939 3438
rect 959 3434 963 3438
rect 1087 3434 1091 3438
rect 1111 3434 1115 3438
rect 1207 3434 1211 3438
rect 1295 3434 1299 3438
rect 1327 3434 1331 3438
rect 1447 3434 1451 3438
rect 1479 3434 1483 3438
rect 1567 3434 1571 3438
rect 1823 3434 1827 3438
rect 1863 3430 1867 3434
rect 1903 3430 1907 3434
rect 1911 3430 1915 3434
rect 2007 3430 2011 3434
rect 2071 3430 2075 3434
rect 2127 3430 2131 3434
rect 2223 3430 2227 3434
rect 2255 3430 2259 3434
rect 2367 3430 2371 3434
rect 2383 3430 2387 3434
rect 2503 3430 2507 3434
rect 2519 3430 2523 3434
rect 2631 3430 2635 3434
rect 2655 3430 2659 3434
rect 2759 3430 2763 3434
rect 2791 3430 2795 3434
rect 2887 3430 2891 3434
rect 2935 3430 2939 3434
rect 3023 3430 3027 3434
rect 3079 3430 3083 3434
rect 3575 3430 3579 3434
rect 111 3358 115 3362
rect 143 3358 147 3362
rect 207 3358 211 3362
rect 263 3358 267 3362
rect 367 3358 371 3362
rect 423 3358 427 3362
rect 535 3358 539 3362
rect 591 3358 595 3362
rect 695 3358 699 3362
rect 767 3358 771 3362
rect 855 3358 859 3362
rect 943 3358 947 3362
rect 999 3358 1003 3362
rect 1119 3358 1123 3362
rect 1143 3358 1147 3362
rect 1279 3358 1283 3362
rect 1303 3358 1307 3362
rect 1415 3358 1419 3362
rect 1487 3358 1491 3362
rect 1559 3358 1563 3362
rect 1823 3358 1827 3362
rect 1863 3358 1867 3362
rect 1895 3358 1899 3362
rect 1919 3358 1923 3362
rect 2047 3358 2051 3362
rect 2079 3358 2083 3362
rect 2207 3358 2211 3362
rect 2231 3358 2235 3362
rect 2367 3358 2371 3362
rect 2375 3358 2379 3362
rect 2511 3358 2515 3362
rect 2535 3358 2539 3362
rect 2639 3358 2643 3362
rect 2703 3358 2707 3362
rect 2767 3358 2771 3362
rect 2879 3358 2883 3362
rect 2895 3358 2899 3362
rect 3031 3358 3035 3362
rect 3055 3358 3059 3362
rect 3575 3358 3579 3362
rect 111 3286 115 3290
rect 199 3286 203 3290
rect 255 3286 259 3290
rect 359 3286 363 3290
rect 375 3286 379 3290
rect 511 3286 515 3290
rect 527 3286 531 3290
rect 663 3286 667 3290
rect 687 3286 691 3290
rect 823 3286 827 3290
rect 847 3286 851 3290
rect 991 3286 995 3290
rect 1135 3286 1139 3290
rect 1167 3286 1171 3290
rect 1271 3286 1275 3290
rect 1343 3286 1347 3290
rect 1407 3286 1411 3290
rect 1519 3286 1523 3290
rect 1551 3286 1555 3290
rect 1823 3286 1827 3290
rect 1863 3286 1867 3290
rect 1887 3286 1891 3290
rect 2039 3286 2043 3290
rect 2063 3286 2067 3290
rect 2199 3286 2203 3290
rect 2263 3286 2267 3290
rect 2359 3286 2363 3290
rect 2455 3286 2459 3290
rect 2527 3286 2531 3290
rect 2639 3286 2643 3290
rect 2695 3286 2699 3290
rect 2815 3286 2819 3290
rect 2871 3286 2875 3290
rect 2983 3286 2987 3290
rect 3047 3286 3051 3290
rect 3151 3286 3155 3290
rect 3319 3286 3323 3290
rect 3479 3286 3483 3290
rect 3575 3286 3579 3290
rect 111 3214 115 3218
rect 263 3214 267 3218
rect 383 3214 387 3218
rect 431 3214 435 3218
rect 519 3214 523 3218
rect 551 3214 555 3218
rect 671 3214 675 3218
rect 799 3214 803 3218
rect 831 3214 835 3218
rect 935 3214 939 3218
rect 999 3214 1003 3218
rect 1079 3214 1083 3218
rect 1175 3214 1179 3218
rect 1231 3214 1235 3218
rect 1351 3214 1355 3218
rect 1383 3214 1387 3218
rect 1527 3214 1531 3218
rect 1535 3214 1539 3218
rect 1823 3214 1827 3218
rect 1863 3218 1867 3222
rect 1895 3218 1899 3222
rect 2071 3218 2075 3222
rect 2087 3218 2091 3222
rect 2271 3218 2275 3222
rect 2303 3218 2307 3222
rect 2463 3218 2467 3222
rect 2511 3218 2515 3222
rect 2647 3218 2651 3222
rect 2703 3218 2707 3222
rect 2823 3218 2827 3222
rect 2879 3218 2883 3222
rect 2991 3218 2995 3222
rect 3039 3218 3043 3222
rect 3159 3218 3163 3222
rect 3199 3218 3203 3222
rect 3327 3218 3331 3222
rect 3351 3218 3355 3222
rect 3487 3218 3491 3222
rect 3575 3218 3579 3222
rect 111 3142 115 3146
rect 423 3142 427 3146
rect 463 3142 467 3146
rect 543 3142 547 3146
rect 551 3142 555 3146
rect 639 3142 643 3146
rect 663 3142 667 3146
rect 735 3142 739 3146
rect 791 3142 795 3146
rect 847 3142 851 3146
rect 927 3142 931 3146
rect 967 3142 971 3146
rect 1071 3142 1075 3146
rect 1095 3142 1099 3146
rect 1223 3142 1227 3146
rect 1231 3142 1235 3146
rect 1375 3142 1379 3146
rect 1519 3142 1523 3146
rect 1527 3142 1531 3146
rect 1823 3142 1827 3146
rect 1863 3146 1867 3150
rect 1887 3146 1891 3150
rect 2079 3146 2083 3150
rect 2295 3146 2299 3150
rect 2503 3146 2507 3150
rect 2695 3146 2699 3150
rect 2871 3146 2875 3150
rect 3031 3146 3035 3150
rect 3039 3146 3043 3150
rect 3191 3146 3195 3150
rect 3343 3146 3347 3150
rect 3479 3146 3483 3150
rect 3575 3146 3579 3150
rect 111 3066 115 3070
rect 151 3066 155 3070
rect 239 3066 243 3070
rect 327 3066 331 3070
rect 415 3066 419 3070
rect 471 3066 475 3070
rect 503 3066 507 3070
rect 559 3066 563 3070
rect 591 3066 595 3070
rect 647 3066 651 3070
rect 679 3066 683 3070
rect 743 3066 747 3070
rect 767 3066 771 3070
rect 855 3066 859 3070
rect 943 3066 947 3070
rect 975 3066 979 3070
rect 1031 3066 1035 3070
rect 1103 3066 1107 3070
rect 1119 3066 1123 3070
rect 1207 3066 1211 3070
rect 1239 3066 1243 3070
rect 1295 3066 1299 3070
rect 1383 3066 1387 3070
rect 1471 3066 1475 3070
rect 1527 3066 1531 3070
rect 1559 3066 1563 3070
rect 1647 3066 1651 3070
rect 1735 3066 1739 3070
rect 1823 3066 1827 3070
rect 1863 3066 1867 3070
rect 1895 3066 1899 3070
rect 2087 3066 2091 3070
rect 2255 3066 2259 3070
rect 2303 3066 2307 3070
rect 2423 3066 2427 3070
rect 2511 3066 2515 3070
rect 2591 3066 2595 3070
rect 2703 3066 2707 3070
rect 2751 3066 2755 3070
rect 2879 3066 2883 3070
rect 2919 3066 2923 3070
rect 3047 3066 3051 3070
rect 3087 3066 3091 3070
rect 3199 3066 3203 3070
rect 3351 3066 3355 3070
rect 3487 3066 3491 3070
rect 3575 3066 3579 3070
rect 111 2990 115 2994
rect 143 2990 147 2994
rect 231 2990 235 2994
rect 319 2990 323 2994
rect 407 2990 411 2994
rect 495 2990 499 2994
rect 583 2990 587 2994
rect 671 2990 675 2994
rect 759 2990 763 2994
rect 847 2990 851 2994
rect 935 2990 939 2994
rect 1023 2990 1027 2994
rect 1111 2990 1115 2994
rect 1199 2990 1203 2994
rect 1287 2990 1291 2994
rect 1375 2990 1379 2994
rect 1407 2990 1411 2994
rect 1463 2990 1467 2994
rect 1519 2990 1523 2994
rect 1551 2990 1555 2994
rect 1631 2990 1635 2994
rect 1639 2990 1643 2994
rect 1727 2990 1731 2994
rect 1823 2990 1827 2994
rect 1863 2994 1867 2998
rect 2239 2994 2243 2998
rect 2247 2994 2251 2998
rect 2415 2994 2419 2998
rect 2463 2994 2467 2998
rect 2583 2994 2587 2998
rect 2671 2994 2675 2998
rect 2743 2994 2747 2998
rect 2863 2994 2867 2998
rect 2911 2994 2915 2998
rect 3031 2994 3035 2998
rect 3079 2994 3083 2998
rect 3191 2994 3195 2998
rect 3343 2994 3347 2998
rect 3479 2994 3483 2998
rect 3575 2994 3579 2998
rect 111 2922 115 2926
rect 1359 2922 1363 2926
rect 1415 2922 1419 2926
rect 1471 2922 1475 2926
rect 1527 2922 1531 2926
rect 1583 2922 1587 2926
rect 1639 2922 1643 2926
rect 1703 2922 1707 2926
rect 1735 2922 1739 2926
rect 1823 2922 1827 2926
rect 1863 2910 1867 2914
rect 2239 2910 2243 2914
rect 2247 2910 2251 2914
rect 2463 2910 2467 2914
rect 2471 2910 2475 2914
rect 2671 2910 2675 2914
rect 2679 2910 2683 2914
rect 2855 2910 2859 2914
rect 2871 2910 2875 2914
rect 3023 2910 3027 2914
rect 3039 2910 3043 2914
rect 3183 2910 3187 2914
rect 3199 2910 3203 2914
rect 3335 2910 3339 2914
rect 3351 2910 3355 2914
rect 3487 2910 3491 2914
rect 3575 2910 3579 2914
rect 111 2850 115 2854
rect 135 2850 139 2854
rect 223 2850 227 2854
rect 311 2850 315 2854
rect 399 2850 403 2854
rect 487 2850 491 2854
rect 599 2850 603 2854
rect 727 2850 731 2854
rect 863 2850 867 2854
rect 999 2850 1003 2854
rect 1135 2850 1139 2854
rect 1263 2850 1267 2854
rect 1351 2850 1355 2854
rect 1383 2850 1387 2854
rect 1463 2850 1467 2854
rect 1503 2850 1507 2854
rect 1575 2850 1579 2854
rect 1623 2850 1627 2854
rect 1695 2850 1699 2854
rect 1727 2850 1731 2854
rect 1823 2850 1827 2854
rect 1863 2838 1867 2842
rect 1895 2838 1899 2842
rect 1983 2838 1987 2842
rect 2071 2838 2075 2842
rect 2159 2838 2163 2842
rect 2231 2838 2235 2842
rect 2247 2838 2251 2842
rect 2335 2838 2339 2842
rect 2423 2838 2427 2842
rect 2455 2838 2459 2842
rect 2511 2838 2515 2842
rect 2599 2838 2603 2842
rect 2663 2838 2667 2842
rect 2687 2838 2691 2842
rect 2791 2838 2795 2842
rect 2847 2838 2851 2842
rect 2903 2838 2907 2842
rect 3015 2838 3019 2842
rect 3031 2838 3035 2842
rect 3175 2838 3179 2842
rect 3327 2838 3331 2842
rect 3479 2838 3483 2842
rect 3575 2838 3579 2842
rect 111 2782 115 2786
rect 143 2782 147 2786
rect 191 2782 195 2786
rect 231 2782 235 2786
rect 295 2782 299 2786
rect 319 2782 323 2786
rect 407 2782 411 2786
rect 415 2782 419 2786
rect 495 2782 499 2786
rect 551 2782 555 2786
rect 607 2782 611 2786
rect 687 2782 691 2786
rect 735 2782 739 2786
rect 823 2782 827 2786
rect 871 2782 875 2786
rect 959 2782 963 2786
rect 1007 2782 1011 2786
rect 1087 2782 1091 2786
rect 1143 2782 1147 2786
rect 1207 2782 1211 2786
rect 1271 2782 1275 2786
rect 1319 2782 1323 2786
rect 1391 2782 1395 2786
rect 1431 2782 1435 2786
rect 1511 2782 1515 2786
rect 1535 2782 1539 2786
rect 1631 2782 1635 2786
rect 1647 2782 1651 2786
rect 1735 2782 1739 2786
rect 1823 2782 1827 2786
rect 1863 2758 1867 2762
rect 1903 2758 1907 2762
rect 1991 2758 1995 2762
rect 2047 2758 2051 2762
rect 2079 2758 2083 2762
rect 2167 2758 2171 2762
rect 2255 2758 2259 2762
rect 2295 2758 2299 2762
rect 2343 2758 2347 2762
rect 2431 2758 2435 2762
rect 2447 2758 2451 2762
rect 2519 2758 2523 2762
rect 2607 2758 2611 2762
rect 2623 2758 2627 2762
rect 2695 2758 2699 2762
rect 2799 2758 2803 2762
rect 2823 2758 2827 2762
rect 2911 2758 2915 2762
rect 3039 2758 3043 2762
rect 3183 2758 3187 2762
rect 3271 2758 3275 2762
rect 3335 2758 3339 2762
rect 3487 2758 3491 2762
rect 3575 2758 3579 2762
rect 111 2706 115 2710
rect 167 2706 171 2710
rect 183 2706 187 2710
rect 279 2706 283 2710
rect 287 2706 291 2710
rect 391 2706 395 2710
rect 407 2706 411 2710
rect 503 2706 507 2710
rect 543 2706 547 2710
rect 615 2706 619 2710
rect 679 2706 683 2710
rect 815 2706 819 2710
rect 951 2706 955 2710
rect 1079 2706 1083 2710
rect 1199 2706 1203 2710
rect 1311 2706 1315 2710
rect 1423 2706 1427 2710
rect 1527 2706 1531 2710
rect 1639 2706 1643 2710
rect 1727 2706 1731 2710
rect 1823 2706 1827 2710
rect 1863 2690 1867 2694
rect 1943 2690 1947 2694
rect 2039 2690 2043 2694
rect 2055 2690 2059 2694
rect 2159 2690 2163 2694
rect 2167 2690 2171 2694
rect 2287 2690 2291 2694
rect 2407 2690 2411 2694
rect 2439 2690 2443 2694
rect 2519 2690 2523 2694
rect 2615 2690 2619 2694
rect 2631 2690 2635 2694
rect 2735 2690 2739 2694
rect 2815 2690 2819 2694
rect 2847 2690 2851 2694
rect 2959 2690 2963 2694
rect 3031 2690 3035 2694
rect 3071 2690 3075 2694
rect 3263 2690 3267 2694
rect 3479 2690 3483 2694
rect 3575 2690 3579 2694
rect 111 2622 115 2626
rect 175 2622 179 2626
rect 223 2622 227 2626
rect 287 2622 291 2626
rect 351 2622 355 2626
rect 399 2622 403 2626
rect 495 2622 499 2626
rect 511 2622 515 2626
rect 623 2622 627 2626
rect 663 2622 667 2626
rect 839 2622 843 2626
rect 1023 2622 1027 2626
rect 1215 2622 1219 2626
rect 1407 2622 1411 2626
rect 1607 2622 1611 2626
rect 1823 2622 1827 2626
rect 1863 2618 1867 2622
rect 1895 2618 1899 2622
rect 1951 2618 1955 2622
rect 2063 2618 2067 2622
rect 2071 2618 2075 2622
rect 2175 2618 2179 2622
rect 2263 2618 2267 2622
rect 2295 2618 2299 2622
rect 2415 2618 2419 2622
rect 2463 2618 2467 2622
rect 2527 2618 2531 2622
rect 2639 2618 2643 2622
rect 2663 2618 2667 2622
rect 2743 2618 2747 2622
rect 2855 2618 2859 2622
rect 2871 2618 2875 2622
rect 2967 2618 2971 2622
rect 3079 2618 3083 2622
rect 3295 2618 3299 2622
rect 3487 2618 3491 2622
rect 3575 2618 3579 2622
rect 111 2554 115 2558
rect 215 2554 219 2558
rect 271 2554 275 2558
rect 343 2554 347 2558
rect 471 2554 475 2558
rect 487 2554 491 2558
rect 655 2554 659 2558
rect 671 2554 675 2558
rect 831 2554 835 2558
rect 855 2554 859 2558
rect 1015 2554 1019 2558
rect 1023 2554 1027 2558
rect 1175 2554 1179 2558
rect 1207 2554 1211 2558
rect 1319 2554 1323 2558
rect 1399 2554 1403 2558
rect 1455 2554 1459 2558
rect 1591 2554 1595 2558
rect 1599 2554 1603 2558
rect 1727 2554 1731 2558
rect 1823 2554 1827 2558
rect 1863 2550 1867 2554
rect 1887 2550 1891 2554
rect 2039 2550 2043 2554
rect 2063 2550 2067 2554
rect 2215 2550 2219 2554
rect 2255 2550 2259 2554
rect 2399 2550 2403 2554
rect 2455 2550 2459 2554
rect 2575 2550 2579 2554
rect 2655 2550 2659 2554
rect 2743 2550 2747 2554
rect 2863 2550 2867 2554
rect 2903 2550 2907 2554
rect 3055 2550 3059 2554
rect 3071 2550 3075 2554
rect 3199 2550 3203 2554
rect 3287 2550 3291 2554
rect 3343 2550 3347 2554
rect 3479 2550 3483 2554
rect 3575 2550 3579 2554
rect 111 2482 115 2486
rect 183 2482 187 2486
rect 279 2482 283 2486
rect 319 2482 323 2486
rect 463 2482 467 2486
rect 479 2482 483 2486
rect 607 2482 611 2486
rect 679 2482 683 2486
rect 743 2482 747 2486
rect 863 2482 867 2486
rect 879 2482 883 2486
rect 1007 2482 1011 2486
rect 1031 2482 1035 2486
rect 1127 2482 1131 2486
rect 1183 2482 1187 2486
rect 1239 2482 1243 2486
rect 1327 2482 1331 2486
rect 1343 2482 1347 2486
rect 1447 2482 1451 2486
rect 1463 2482 1467 2486
rect 1551 2482 1555 2486
rect 1599 2482 1603 2486
rect 1647 2482 1651 2486
rect 1735 2482 1739 2486
rect 1823 2482 1827 2486
rect 1863 2482 1867 2486
rect 1895 2482 1899 2486
rect 1991 2482 1995 2486
rect 2047 2482 2051 2486
rect 2127 2482 2131 2486
rect 2223 2482 2227 2486
rect 2279 2482 2283 2486
rect 2407 2482 2411 2486
rect 2439 2482 2443 2486
rect 2583 2482 2587 2486
rect 2599 2482 2603 2486
rect 2751 2482 2755 2486
rect 2767 2482 2771 2486
rect 2911 2482 2915 2486
rect 2943 2482 2947 2486
rect 3063 2482 3067 2486
rect 3119 2482 3123 2486
rect 3207 2482 3211 2486
rect 3295 2482 3299 2486
rect 3351 2482 3355 2486
rect 3471 2482 3475 2486
rect 3487 2482 3491 2486
rect 3575 2482 3579 2486
rect 111 2406 115 2410
rect 151 2406 155 2410
rect 175 2406 179 2410
rect 311 2406 315 2410
rect 319 2406 323 2410
rect 455 2406 459 2410
rect 479 2406 483 2410
rect 599 2406 603 2410
rect 639 2406 643 2410
rect 735 2406 739 2410
rect 783 2406 787 2410
rect 871 2406 875 2410
rect 919 2406 923 2410
rect 999 2406 1003 2410
rect 1047 2406 1051 2410
rect 1119 2406 1123 2410
rect 1175 2406 1179 2410
rect 1231 2406 1235 2410
rect 1303 2406 1307 2410
rect 1335 2406 1339 2410
rect 1431 2406 1435 2410
rect 1439 2406 1443 2410
rect 1543 2406 1547 2410
rect 1639 2406 1643 2410
rect 1727 2406 1731 2410
rect 1823 2406 1827 2410
rect 1863 2406 1867 2410
rect 1887 2406 1891 2410
rect 1983 2406 1987 2410
rect 2119 2406 2123 2410
rect 2271 2406 2275 2410
rect 2351 2406 2355 2410
rect 2431 2406 2435 2410
rect 2503 2406 2507 2410
rect 2591 2406 2595 2410
rect 2655 2406 2659 2410
rect 2759 2406 2763 2410
rect 2807 2406 2811 2410
rect 2935 2406 2939 2410
rect 2967 2406 2971 2410
rect 3111 2406 3115 2410
rect 3135 2406 3139 2410
rect 3287 2406 3291 2410
rect 3303 2406 3307 2410
rect 3463 2406 3467 2410
rect 3471 2406 3475 2410
rect 3575 2406 3579 2410
rect 111 2334 115 2338
rect 143 2334 147 2338
rect 159 2334 163 2338
rect 263 2334 267 2338
rect 327 2334 331 2338
rect 407 2334 411 2338
rect 487 2334 491 2338
rect 543 2334 547 2338
rect 647 2334 651 2338
rect 679 2334 683 2338
rect 791 2334 795 2338
rect 807 2334 811 2338
rect 927 2334 931 2338
rect 1039 2334 1043 2338
rect 1055 2334 1059 2338
rect 1159 2334 1163 2338
rect 1183 2334 1187 2338
rect 1279 2334 1283 2338
rect 1311 2334 1315 2338
rect 1439 2334 1443 2338
rect 1823 2334 1827 2338
rect 1863 2334 1867 2338
rect 2351 2334 2355 2338
rect 2359 2334 2363 2338
rect 2447 2334 2451 2338
rect 2511 2334 2515 2338
rect 2559 2334 2563 2338
rect 2663 2334 2667 2338
rect 2703 2334 2707 2338
rect 2815 2334 2819 2338
rect 2879 2334 2883 2338
rect 2975 2334 2979 2338
rect 3079 2334 3083 2338
rect 3143 2334 3147 2338
rect 3287 2334 3291 2338
rect 3311 2334 3315 2338
rect 3479 2334 3483 2338
rect 3487 2334 3491 2338
rect 3575 2334 3579 2338
rect 111 2266 115 2270
rect 135 2266 139 2270
rect 231 2266 235 2270
rect 255 2266 259 2270
rect 351 2266 355 2270
rect 399 2266 403 2270
rect 471 2266 475 2270
rect 535 2266 539 2270
rect 591 2266 595 2270
rect 671 2266 675 2270
rect 711 2266 715 2270
rect 799 2266 803 2270
rect 823 2266 827 2270
rect 919 2266 923 2270
rect 935 2266 939 2270
rect 1031 2266 1035 2270
rect 1055 2266 1059 2270
rect 1151 2266 1155 2270
rect 1175 2266 1179 2270
rect 1271 2266 1275 2270
rect 1823 2266 1827 2270
rect 1863 2266 1867 2270
rect 2335 2266 2339 2270
rect 2343 2266 2347 2270
rect 2439 2266 2443 2270
rect 2447 2266 2451 2270
rect 2551 2266 2555 2270
rect 2583 2266 2587 2270
rect 2695 2266 2699 2270
rect 2735 2266 2739 2270
rect 2871 2266 2875 2270
rect 2911 2266 2915 2270
rect 3071 2266 3075 2270
rect 3103 2266 3107 2270
rect 3279 2266 3283 2270
rect 3303 2266 3307 2270
rect 3479 2266 3483 2270
rect 3575 2266 3579 2270
rect 111 2194 115 2198
rect 143 2194 147 2198
rect 239 2194 243 2198
rect 247 2194 251 2198
rect 359 2194 363 2198
rect 383 2194 387 2198
rect 479 2194 483 2198
rect 519 2194 523 2198
rect 599 2194 603 2198
rect 655 2194 659 2198
rect 719 2194 723 2198
rect 783 2194 787 2198
rect 831 2194 835 2198
rect 911 2194 915 2198
rect 943 2194 947 2198
rect 1031 2194 1035 2198
rect 1063 2194 1067 2198
rect 1159 2194 1163 2198
rect 1183 2194 1187 2198
rect 1287 2194 1291 2198
rect 1823 2194 1827 2198
rect 1863 2198 1867 2202
rect 2255 2198 2259 2202
rect 2343 2198 2347 2202
rect 2439 2198 2443 2202
rect 2455 2198 2459 2202
rect 2551 2198 2555 2202
rect 2591 2198 2595 2202
rect 2695 2198 2699 2202
rect 2743 2198 2747 2202
rect 2871 2198 2875 2202
rect 2919 2198 2923 2202
rect 3071 2198 3075 2202
rect 3111 2198 3115 2202
rect 3287 2198 3291 2202
rect 3311 2198 3315 2202
rect 3487 2198 3491 2202
rect 3575 2198 3579 2202
rect 111 2118 115 2122
rect 135 2118 139 2122
rect 231 2118 235 2122
rect 239 2118 243 2122
rect 359 2118 363 2122
rect 375 2118 379 2122
rect 479 2118 483 2122
rect 511 2118 515 2122
rect 599 2118 603 2122
rect 647 2118 651 2122
rect 719 2118 723 2122
rect 775 2118 779 2122
rect 831 2118 835 2122
rect 903 2118 907 2122
rect 943 2118 947 2122
rect 1023 2118 1027 2122
rect 1055 2118 1059 2122
rect 1151 2118 1155 2122
rect 1175 2118 1179 2122
rect 1279 2118 1283 2122
rect 1823 2118 1827 2122
rect 1863 2122 1867 2126
rect 2151 2122 2155 2126
rect 2239 2122 2243 2126
rect 2247 2122 2251 2126
rect 2327 2122 2331 2126
rect 2335 2122 2339 2126
rect 2415 2122 2419 2126
rect 2431 2122 2435 2126
rect 2503 2122 2507 2126
rect 2543 2122 2547 2126
rect 2615 2122 2619 2126
rect 2687 2122 2691 2126
rect 2751 2122 2755 2126
rect 2863 2122 2867 2126
rect 2919 2122 2923 2126
rect 3063 2122 3067 2126
rect 3103 2122 3107 2126
rect 3279 2122 3283 2126
rect 3303 2122 3307 2126
rect 3479 2122 3483 2126
rect 3575 2122 3579 2126
rect 1863 2050 1867 2054
rect 1999 2050 2003 2054
rect 2127 2050 2131 2054
rect 2159 2050 2163 2054
rect 2247 2050 2251 2054
rect 2255 2050 2259 2054
rect 2335 2050 2339 2054
rect 2399 2050 2403 2054
rect 2423 2050 2427 2054
rect 2511 2050 2515 2054
rect 2551 2050 2555 2054
rect 2623 2050 2627 2054
rect 2711 2050 2715 2054
rect 2759 2050 2763 2054
rect 2879 2050 2883 2054
rect 2927 2050 2931 2054
rect 3063 2050 3067 2054
rect 3111 2050 3115 2054
rect 3247 2050 3251 2054
rect 3311 2050 3315 2054
rect 3439 2050 3443 2054
rect 3487 2050 3491 2054
rect 3575 2050 3579 2054
rect 111 2038 115 2042
rect 143 2038 147 2042
rect 167 2038 171 2042
rect 239 2038 243 2042
rect 311 2038 315 2042
rect 367 2038 371 2042
rect 447 2038 451 2042
rect 487 2038 491 2042
rect 575 2038 579 2042
rect 607 2038 611 2042
rect 695 2038 699 2042
rect 727 2038 731 2042
rect 807 2038 811 2042
rect 839 2038 843 2042
rect 911 2038 915 2042
rect 951 2038 955 2042
rect 1015 2038 1019 2042
rect 1063 2038 1067 2042
rect 1119 2038 1123 2042
rect 1183 2038 1187 2042
rect 1223 2038 1227 2042
rect 1327 2038 1331 2042
rect 1823 2038 1827 2042
rect 111 1970 115 1974
rect 159 1970 163 1974
rect 295 1970 299 1974
rect 303 1970 307 1974
rect 439 1970 443 1974
rect 567 1970 571 1974
rect 583 1970 587 1974
rect 687 1970 691 1974
rect 719 1970 723 1974
rect 799 1970 803 1974
rect 855 1970 859 1974
rect 903 1970 907 1974
rect 991 1970 995 1974
rect 1007 1970 1011 1974
rect 1111 1970 1115 1974
rect 1119 1970 1123 1974
rect 1215 1970 1219 1974
rect 1239 1970 1243 1974
rect 1319 1970 1323 1974
rect 1359 1970 1363 1974
rect 1479 1970 1483 1974
rect 1599 1970 1603 1974
rect 1823 1970 1827 1974
rect 1863 1974 1867 1978
rect 1903 1974 1907 1978
rect 1991 1974 1995 1978
rect 2119 1974 2123 1978
rect 2159 1974 2163 1978
rect 2247 1974 2251 1978
rect 2391 1974 2395 1978
rect 2399 1974 2403 1978
rect 2543 1974 2547 1978
rect 2615 1974 2619 1978
rect 2703 1974 2707 1978
rect 2815 1974 2819 1978
rect 2871 1974 2875 1978
rect 2999 1974 3003 1978
rect 3055 1974 3059 1978
rect 3167 1974 3171 1978
rect 3239 1974 3243 1978
rect 3335 1974 3339 1978
rect 3431 1974 3435 1978
rect 3479 1974 3483 1978
rect 3575 1974 3579 1978
rect 1863 1906 1867 1910
rect 1895 1906 1899 1910
rect 1911 1906 1915 1910
rect 1983 1906 1987 1910
rect 2071 1906 2075 1910
rect 2167 1906 2171 1910
rect 2295 1906 2299 1910
rect 2407 1906 2411 1910
rect 2447 1906 2451 1910
rect 2607 1906 2611 1910
rect 2623 1906 2627 1910
rect 2767 1906 2771 1910
rect 2823 1906 2827 1910
rect 2919 1906 2923 1910
rect 3007 1906 3011 1910
rect 3071 1906 3075 1910
rect 3175 1906 3179 1910
rect 3215 1906 3219 1910
rect 3343 1906 3347 1910
rect 3359 1906 3363 1910
rect 3487 1906 3491 1910
rect 3575 1906 3579 1910
rect 111 1894 115 1898
rect 167 1894 171 1898
rect 223 1894 227 1898
rect 303 1894 307 1898
rect 447 1894 451 1898
rect 479 1894 483 1898
rect 591 1894 595 1898
rect 719 1894 723 1898
rect 727 1894 731 1898
rect 863 1894 867 1898
rect 935 1894 939 1898
rect 999 1894 1003 1898
rect 1127 1894 1131 1898
rect 1247 1894 1251 1898
rect 1295 1894 1299 1898
rect 1367 1894 1371 1898
rect 1455 1894 1459 1898
rect 1487 1894 1491 1898
rect 1607 1894 1611 1898
rect 1735 1894 1739 1898
rect 1823 1894 1827 1898
rect 1863 1834 1867 1838
rect 1887 1834 1891 1838
rect 1975 1834 1979 1838
rect 1999 1834 2003 1838
rect 2063 1834 2067 1838
rect 2159 1834 2163 1838
rect 2223 1834 2227 1838
rect 2287 1834 2291 1838
rect 2439 1834 2443 1838
rect 2599 1834 2603 1838
rect 2639 1834 2643 1838
rect 2759 1834 2763 1838
rect 2831 1834 2835 1838
rect 2911 1834 2915 1838
rect 3015 1834 3019 1838
rect 3063 1834 3067 1838
rect 3199 1834 3203 1838
rect 3207 1834 3211 1838
rect 3351 1834 3355 1838
rect 3391 1834 3395 1838
rect 3479 1834 3483 1838
rect 3575 1834 3579 1838
rect 111 1826 115 1830
rect 215 1826 219 1830
rect 247 1826 251 1830
rect 415 1826 419 1830
rect 471 1826 475 1830
rect 591 1826 595 1830
rect 711 1826 715 1830
rect 759 1826 763 1830
rect 927 1826 931 1830
rect 1079 1826 1083 1830
rect 1119 1826 1123 1830
rect 1223 1826 1227 1830
rect 1287 1826 1291 1830
rect 1359 1826 1363 1830
rect 1447 1826 1451 1830
rect 1487 1826 1491 1830
rect 1599 1826 1603 1830
rect 1615 1826 1619 1830
rect 1727 1826 1731 1830
rect 1823 1826 1827 1830
rect 1863 1762 1867 1766
rect 1943 1762 1947 1766
rect 2007 1762 2011 1766
rect 2087 1762 2091 1766
rect 2231 1762 2235 1766
rect 2247 1762 2251 1766
rect 2415 1762 2419 1766
rect 2447 1762 2451 1766
rect 2599 1762 2603 1766
rect 2647 1762 2651 1766
rect 2791 1762 2795 1766
rect 2839 1762 2843 1766
rect 2991 1762 2995 1766
rect 3023 1762 3027 1766
rect 3199 1762 3203 1766
rect 3207 1762 3211 1766
rect 3399 1762 3403 1766
rect 3415 1762 3419 1766
rect 3575 1762 3579 1766
rect 111 1754 115 1758
rect 255 1754 259 1758
rect 327 1754 331 1758
rect 423 1754 427 1758
rect 471 1754 475 1758
rect 599 1754 603 1758
rect 615 1754 619 1758
rect 767 1754 771 1758
rect 919 1754 923 1758
rect 935 1754 939 1758
rect 1071 1754 1075 1758
rect 1087 1754 1091 1758
rect 1223 1754 1227 1758
rect 1231 1754 1235 1758
rect 1367 1754 1371 1758
rect 1375 1754 1379 1758
rect 1495 1754 1499 1758
rect 1527 1754 1531 1758
rect 1623 1754 1627 1758
rect 1687 1754 1691 1758
rect 1735 1754 1739 1758
rect 1823 1754 1827 1758
rect 1863 1690 1867 1694
rect 1911 1690 1915 1694
rect 1935 1690 1939 1694
rect 2031 1690 2035 1694
rect 2079 1690 2083 1694
rect 2151 1690 2155 1694
rect 2239 1690 2243 1694
rect 2271 1690 2275 1694
rect 2399 1690 2403 1694
rect 2407 1690 2411 1694
rect 2543 1690 2547 1694
rect 2591 1690 2595 1694
rect 2695 1690 2699 1694
rect 2783 1690 2787 1694
rect 2863 1690 2867 1694
rect 2983 1690 2987 1694
rect 3047 1690 3051 1694
rect 3191 1690 3195 1694
rect 3239 1690 3243 1694
rect 3407 1690 3411 1694
rect 3431 1690 3435 1694
rect 3575 1690 3579 1694
rect 111 1682 115 1686
rect 311 1682 315 1686
rect 319 1682 323 1686
rect 447 1682 451 1686
rect 463 1682 467 1686
rect 591 1682 595 1686
rect 607 1682 611 1686
rect 735 1682 739 1686
rect 759 1682 763 1686
rect 887 1682 891 1686
rect 911 1682 915 1686
rect 1039 1682 1043 1686
rect 1063 1682 1067 1686
rect 1191 1682 1195 1686
rect 1215 1682 1219 1686
rect 1343 1682 1347 1686
rect 1367 1682 1371 1686
rect 1495 1682 1499 1686
rect 1519 1682 1523 1686
rect 1647 1682 1651 1686
rect 1679 1682 1683 1686
rect 1823 1682 1827 1686
rect 1863 1614 1867 1618
rect 1895 1614 1899 1618
rect 1919 1614 1923 1618
rect 2015 1614 2019 1618
rect 2039 1614 2043 1618
rect 2151 1614 2155 1618
rect 2159 1614 2163 1618
rect 2279 1614 2283 1618
rect 2287 1614 2291 1618
rect 2407 1614 2411 1618
rect 2431 1614 2435 1618
rect 2551 1614 2555 1618
rect 2583 1614 2587 1618
rect 2703 1614 2707 1618
rect 2743 1614 2747 1618
rect 2871 1614 2875 1618
rect 2911 1614 2915 1618
rect 3055 1614 3059 1618
rect 3095 1614 3099 1618
rect 3247 1614 3251 1618
rect 3279 1614 3283 1618
rect 3439 1614 3443 1618
rect 3471 1614 3475 1618
rect 3575 1614 3579 1618
rect 111 1606 115 1610
rect 223 1606 227 1610
rect 319 1606 323 1610
rect 351 1606 355 1610
rect 455 1606 459 1610
rect 487 1606 491 1610
rect 599 1606 603 1610
rect 623 1606 627 1610
rect 743 1606 747 1610
rect 759 1606 763 1610
rect 895 1606 899 1610
rect 903 1606 907 1610
rect 1047 1606 1051 1610
rect 1055 1606 1059 1610
rect 1199 1606 1203 1610
rect 1215 1606 1219 1610
rect 1351 1606 1355 1610
rect 1375 1606 1379 1610
rect 1503 1606 1507 1610
rect 1543 1606 1547 1610
rect 1655 1606 1659 1610
rect 1823 1606 1827 1610
rect 111 1534 115 1538
rect 135 1534 139 1538
rect 215 1534 219 1538
rect 271 1534 275 1538
rect 343 1534 347 1538
rect 423 1534 427 1538
rect 479 1534 483 1538
rect 583 1534 587 1538
rect 615 1534 619 1538
rect 735 1534 739 1538
rect 751 1534 755 1538
rect 887 1534 891 1538
rect 895 1534 899 1538
rect 1039 1534 1043 1538
rect 1047 1534 1051 1538
rect 1191 1534 1195 1538
rect 1207 1534 1211 1538
rect 1343 1534 1347 1538
rect 1367 1534 1371 1538
rect 1495 1534 1499 1538
rect 1535 1534 1539 1538
rect 1823 1534 1827 1538
rect 1863 1538 1867 1542
rect 1887 1538 1891 1542
rect 2007 1538 2011 1542
rect 2023 1538 2027 1542
rect 2143 1538 2147 1542
rect 2183 1538 2187 1542
rect 2279 1538 2283 1542
rect 2343 1538 2347 1542
rect 2423 1538 2427 1542
rect 2503 1538 2507 1542
rect 2575 1538 2579 1542
rect 2663 1538 2667 1542
rect 2735 1538 2739 1542
rect 2823 1538 2827 1542
rect 2903 1538 2907 1542
rect 2983 1538 2987 1542
rect 3087 1538 3091 1542
rect 3151 1538 3155 1542
rect 3271 1538 3275 1542
rect 3319 1538 3323 1542
rect 3463 1538 3467 1542
rect 3479 1538 3483 1542
rect 3575 1538 3579 1542
rect 111 1458 115 1462
rect 143 1458 147 1462
rect 263 1458 267 1462
rect 279 1458 283 1462
rect 399 1458 403 1462
rect 431 1458 435 1462
rect 535 1458 539 1462
rect 591 1458 595 1462
rect 663 1458 667 1462
rect 743 1458 747 1462
rect 791 1458 795 1462
rect 895 1458 899 1462
rect 911 1458 915 1462
rect 1023 1458 1027 1462
rect 1047 1458 1051 1462
rect 1143 1458 1147 1462
rect 1199 1458 1203 1462
rect 1263 1458 1267 1462
rect 1351 1458 1355 1462
rect 1383 1458 1387 1462
rect 1503 1458 1507 1462
rect 1631 1458 1635 1462
rect 1735 1458 1739 1462
rect 1823 1458 1827 1462
rect 1863 1462 1867 1466
rect 1895 1462 1899 1466
rect 2031 1462 2035 1466
rect 2183 1462 2187 1466
rect 2191 1462 2195 1466
rect 2351 1462 2355 1466
rect 2359 1462 2363 1466
rect 2511 1462 2515 1466
rect 2527 1462 2531 1466
rect 2671 1462 2675 1466
rect 2687 1462 2691 1466
rect 2831 1462 2835 1466
rect 2847 1462 2851 1466
rect 2991 1462 2995 1466
rect 3007 1462 3011 1466
rect 3159 1462 3163 1466
rect 3175 1462 3179 1466
rect 3327 1462 3331 1466
rect 3343 1462 3347 1466
rect 3487 1462 3491 1466
rect 3575 1462 3579 1466
rect 111 1390 115 1394
rect 135 1390 139 1394
rect 255 1390 259 1394
rect 327 1390 331 1394
rect 391 1390 395 1394
rect 527 1390 531 1394
rect 551 1390 555 1394
rect 655 1390 659 1394
rect 783 1390 787 1394
rect 903 1390 907 1394
rect 1015 1390 1019 1394
rect 1023 1390 1027 1394
rect 1135 1390 1139 1394
rect 1255 1390 1259 1394
rect 1263 1390 1267 1394
rect 1375 1390 1379 1394
rect 1495 1390 1499 1394
rect 1503 1390 1507 1394
rect 1623 1390 1627 1394
rect 1727 1390 1731 1394
rect 1823 1390 1827 1394
rect 1863 1386 1867 1390
rect 2079 1386 2083 1390
rect 2175 1386 2179 1390
rect 2263 1386 2267 1390
rect 2351 1386 2355 1390
rect 2439 1386 2443 1390
rect 2519 1386 2523 1390
rect 2615 1386 2619 1390
rect 2679 1386 2683 1390
rect 2783 1386 2787 1390
rect 2839 1386 2843 1390
rect 2935 1386 2939 1390
rect 2999 1386 3003 1390
rect 3079 1386 3083 1390
rect 3167 1386 3171 1390
rect 3223 1386 3227 1390
rect 3335 1386 3339 1390
rect 3359 1386 3363 1390
rect 3479 1386 3483 1390
rect 3575 1386 3579 1390
rect 111 1314 115 1318
rect 143 1314 147 1318
rect 327 1314 331 1318
rect 335 1314 339 1318
rect 527 1314 531 1318
rect 559 1314 563 1318
rect 719 1314 723 1318
rect 791 1314 795 1318
rect 903 1314 907 1318
rect 1031 1314 1035 1318
rect 1071 1314 1075 1318
rect 1231 1314 1235 1318
rect 1271 1314 1275 1318
rect 1383 1314 1387 1318
rect 1511 1314 1515 1318
rect 1535 1314 1539 1318
rect 1687 1314 1691 1318
rect 1735 1314 1739 1318
rect 1823 1314 1827 1318
rect 1863 1318 1867 1322
rect 2087 1318 2091 1322
rect 2271 1318 2275 1322
rect 2311 1318 2315 1322
rect 2447 1318 2451 1322
rect 2519 1318 2523 1322
rect 2623 1318 2627 1322
rect 2711 1318 2715 1322
rect 2791 1318 2795 1322
rect 2887 1318 2891 1322
rect 2943 1318 2947 1322
rect 3047 1318 3051 1322
rect 3087 1318 3091 1322
rect 3199 1318 3203 1322
rect 3231 1318 3235 1322
rect 3351 1318 3355 1322
rect 3367 1318 3371 1322
rect 3487 1318 3491 1322
rect 3575 1318 3579 1322
rect 111 1242 115 1246
rect 135 1242 139 1246
rect 295 1242 299 1246
rect 319 1242 323 1246
rect 479 1242 483 1246
rect 519 1242 523 1246
rect 655 1242 659 1246
rect 711 1242 715 1246
rect 815 1242 819 1246
rect 895 1242 899 1246
rect 967 1242 971 1246
rect 1063 1242 1067 1246
rect 1111 1242 1115 1246
rect 1223 1242 1227 1246
rect 1247 1242 1251 1246
rect 1375 1242 1379 1246
rect 1383 1242 1387 1246
rect 1527 1242 1531 1246
rect 1679 1242 1683 1246
rect 1823 1242 1827 1246
rect 1863 1246 1867 1250
rect 1903 1246 1907 1250
rect 1991 1246 1995 1250
rect 2079 1246 2083 1250
rect 2095 1246 2099 1250
rect 2215 1246 2219 1250
rect 2303 1246 2307 1250
rect 2351 1246 2355 1250
rect 2487 1246 2491 1250
rect 2511 1246 2515 1250
rect 2631 1246 2635 1250
rect 2703 1246 2707 1250
rect 2775 1246 2779 1250
rect 2879 1246 2883 1250
rect 2919 1246 2923 1250
rect 3039 1246 3043 1250
rect 3063 1246 3067 1250
rect 3191 1246 3195 1250
rect 3207 1246 3211 1250
rect 3343 1246 3347 1250
rect 3351 1246 3355 1250
rect 3479 1246 3483 1250
rect 3575 1246 3579 1250
rect 111 1170 115 1174
rect 143 1170 147 1174
rect 167 1170 171 1174
rect 303 1170 307 1174
rect 319 1170 323 1174
rect 471 1170 475 1174
rect 487 1170 491 1174
rect 615 1170 619 1174
rect 663 1170 667 1174
rect 759 1170 763 1174
rect 823 1170 827 1174
rect 911 1170 915 1174
rect 975 1170 979 1174
rect 1063 1170 1067 1174
rect 1119 1170 1123 1174
rect 1231 1170 1235 1174
rect 1255 1170 1259 1174
rect 1391 1170 1395 1174
rect 1399 1170 1403 1174
rect 1535 1170 1539 1174
rect 1575 1170 1579 1174
rect 1735 1170 1739 1174
rect 1823 1170 1827 1174
rect 1863 1174 1867 1178
rect 1895 1174 1899 1178
rect 1911 1174 1915 1178
rect 1999 1174 2003 1178
rect 2063 1174 2067 1178
rect 2103 1174 2107 1178
rect 2223 1174 2227 1178
rect 2255 1174 2259 1178
rect 2359 1174 2363 1178
rect 2439 1174 2443 1178
rect 2495 1174 2499 1178
rect 2615 1174 2619 1178
rect 2639 1174 2643 1178
rect 2783 1174 2787 1178
rect 2791 1174 2795 1178
rect 2927 1174 2931 1178
rect 2967 1174 2971 1178
rect 3071 1174 3075 1178
rect 3143 1174 3147 1178
rect 3215 1174 3219 1178
rect 3327 1174 3331 1178
rect 3359 1174 3363 1178
rect 3487 1174 3491 1178
rect 3575 1174 3579 1178
rect 111 1098 115 1102
rect 159 1098 163 1102
rect 215 1098 219 1102
rect 311 1098 315 1102
rect 327 1098 331 1102
rect 439 1098 443 1102
rect 463 1098 467 1102
rect 559 1098 563 1102
rect 607 1098 611 1102
rect 679 1098 683 1102
rect 751 1098 755 1102
rect 807 1098 811 1102
rect 903 1098 907 1102
rect 943 1098 947 1102
rect 1055 1098 1059 1102
rect 1087 1098 1091 1102
rect 1223 1098 1227 1102
rect 1247 1098 1251 1102
rect 1391 1098 1395 1102
rect 1407 1098 1411 1102
rect 1567 1098 1571 1102
rect 1575 1098 1579 1102
rect 1727 1098 1731 1102
rect 1823 1098 1827 1102
rect 1863 1094 1867 1098
rect 1887 1094 1891 1098
rect 1935 1094 1939 1098
rect 2055 1094 2059 1098
rect 2095 1094 2099 1098
rect 2247 1094 2251 1098
rect 2407 1094 2411 1098
rect 2431 1094 2435 1098
rect 2567 1094 2571 1098
rect 2607 1094 2611 1098
rect 2735 1094 2739 1098
rect 2783 1094 2787 1098
rect 2911 1094 2915 1098
rect 2959 1094 2963 1098
rect 3095 1094 3099 1098
rect 3135 1094 3139 1098
rect 3287 1094 3291 1098
rect 3319 1094 3323 1098
rect 3479 1094 3483 1098
rect 3575 1094 3579 1098
rect 111 1022 115 1026
rect 223 1022 227 1026
rect 335 1022 339 1026
rect 343 1022 347 1026
rect 431 1022 435 1026
rect 447 1022 451 1026
rect 535 1022 539 1026
rect 567 1022 571 1026
rect 655 1022 659 1026
rect 687 1022 691 1026
rect 791 1022 795 1026
rect 815 1022 819 1026
rect 951 1022 955 1026
rect 1095 1022 1099 1026
rect 1135 1022 1139 1026
rect 1255 1022 1259 1026
rect 1327 1022 1331 1026
rect 1415 1022 1419 1026
rect 1535 1022 1539 1026
rect 1583 1022 1587 1026
rect 1735 1022 1739 1026
rect 1823 1022 1827 1026
rect 1863 1022 1867 1026
rect 1943 1022 1947 1026
rect 2071 1022 2075 1026
rect 2103 1022 2107 1026
rect 2191 1022 2195 1026
rect 2255 1022 2259 1026
rect 2311 1022 2315 1026
rect 2415 1022 2419 1026
rect 2439 1022 2443 1026
rect 2575 1022 2579 1026
rect 2719 1022 2723 1026
rect 2743 1022 2747 1026
rect 2871 1022 2875 1026
rect 2919 1022 2923 1026
rect 3031 1022 3035 1026
rect 3103 1022 3107 1026
rect 3191 1022 3195 1026
rect 3295 1022 3299 1026
rect 3351 1022 3355 1026
rect 3487 1022 3491 1026
rect 3575 1022 3579 1026
rect 111 950 115 954
rect 335 950 339 954
rect 367 950 371 954
rect 423 950 427 954
rect 463 950 467 954
rect 527 950 531 954
rect 575 950 579 954
rect 647 950 651 954
rect 703 950 707 954
rect 783 950 787 954
rect 847 950 851 954
rect 943 950 947 954
rect 1007 950 1011 954
rect 1127 950 1131 954
rect 1175 950 1179 954
rect 1319 950 1323 954
rect 1351 950 1355 954
rect 1527 950 1531 954
rect 1711 950 1715 954
rect 1727 950 1731 954
rect 1823 950 1827 954
rect 1863 950 1867 954
rect 1887 950 1891 954
rect 1935 950 1939 954
rect 2047 950 2051 954
rect 2063 950 2067 954
rect 2183 950 2187 954
rect 2199 950 2203 954
rect 2303 950 2307 954
rect 2351 950 2355 954
rect 2431 950 2435 954
rect 2495 950 2499 954
rect 2567 950 2571 954
rect 2631 950 2635 954
rect 2711 950 2715 954
rect 2759 950 2763 954
rect 2863 950 2867 954
rect 2887 950 2891 954
rect 3023 950 3027 954
rect 3183 950 3187 954
rect 3343 950 3347 954
rect 3479 950 3483 954
rect 3575 950 3579 954
rect 111 878 115 882
rect 343 878 347 882
rect 375 878 379 882
rect 431 878 435 882
rect 471 878 475 882
rect 535 878 539 882
rect 583 878 587 882
rect 647 878 651 882
rect 711 878 715 882
rect 783 878 787 882
rect 855 878 859 882
rect 927 878 931 882
rect 1015 878 1019 882
rect 1087 878 1091 882
rect 1183 878 1187 882
rect 1263 878 1267 882
rect 1359 878 1363 882
rect 1447 878 1451 882
rect 1535 878 1539 882
rect 1631 878 1635 882
rect 1719 878 1723 882
rect 1823 878 1827 882
rect 1863 882 1867 886
rect 1895 882 1899 886
rect 2015 882 2019 886
rect 2055 882 2059 886
rect 2167 882 2171 886
rect 2207 882 2211 886
rect 2319 882 2323 886
rect 2359 882 2363 886
rect 2487 882 2491 886
rect 2503 882 2507 886
rect 2639 882 2643 886
rect 2663 882 2667 886
rect 2767 882 2771 886
rect 2847 882 2851 886
rect 2895 882 2899 886
rect 3031 882 3035 886
rect 3039 882 3043 886
rect 3239 882 3243 886
rect 3439 882 3443 886
rect 3575 882 3579 886
rect 111 810 115 814
rect 287 810 291 814
rect 335 810 339 814
rect 407 810 411 814
rect 423 810 427 814
rect 527 810 531 814
rect 535 810 539 814
rect 639 810 643 814
rect 679 810 683 814
rect 775 810 779 814
rect 823 810 827 814
rect 919 810 923 814
rect 975 810 979 814
rect 1079 810 1083 814
rect 1127 810 1131 814
rect 1255 810 1259 814
rect 1279 810 1283 814
rect 1439 810 1443 814
rect 1599 810 1603 814
rect 1623 810 1627 814
rect 1823 810 1827 814
rect 1863 814 1867 818
rect 1887 814 1891 818
rect 1991 814 1995 818
rect 2007 814 2011 818
rect 2135 814 2139 818
rect 2159 814 2163 818
rect 2287 814 2291 818
rect 2311 814 2315 818
rect 2455 814 2459 818
rect 2479 814 2483 818
rect 2623 814 2627 818
rect 2655 814 2659 818
rect 2799 814 2803 818
rect 2839 814 2843 818
rect 2967 814 2971 818
rect 3031 814 3035 818
rect 3143 814 3147 818
rect 3231 814 3235 818
rect 3319 814 3323 818
rect 3431 814 3435 818
rect 3479 814 3483 818
rect 3575 814 3579 818
rect 111 738 115 742
rect 215 738 219 742
rect 295 738 299 742
rect 359 738 363 742
rect 415 738 419 742
rect 503 738 507 742
rect 543 738 547 742
rect 647 738 651 742
rect 687 738 691 742
rect 791 738 795 742
rect 831 738 835 742
rect 935 738 939 742
rect 983 738 987 742
rect 1087 738 1091 742
rect 1135 738 1139 742
rect 1247 738 1251 742
rect 1287 738 1291 742
rect 1415 738 1419 742
rect 1447 738 1451 742
rect 1583 738 1587 742
rect 1607 738 1611 742
rect 1735 738 1739 742
rect 1823 738 1827 742
rect 1863 742 1867 746
rect 1895 742 1899 746
rect 1999 742 2003 746
rect 2063 742 2067 746
rect 2143 742 2147 746
rect 2255 742 2259 746
rect 2295 742 2299 746
rect 2447 742 2451 746
rect 2463 742 2467 746
rect 2631 742 2635 746
rect 2639 742 2643 746
rect 2807 742 2811 746
rect 2823 742 2827 746
rect 2975 742 2979 746
rect 2999 742 3003 746
rect 3151 742 3155 746
rect 3167 742 3171 746
rect 3327 742 3331 746
rect 3335 742 3339 746
rect 3487 742 3491 746
rect 3575 742 3579 746
rect 111 670 115 674
rect 135 670 139 674
rect 207 670 211 674
rect 295 670 299 674
rect 351 670 355 674
rect 463 670 467 674
rect 495 670 499 674
rect 623 670 627 674
rect 639 670 643 674
rect 775 670 779 674
rect 783 670 787 674
rect 927 670 931 674
rect 1071 670 1075 674
rect 1079 670 1083 674
rect 1207 670 1211 674
rect 1239 670 1243 674
rect 1343 670 1347 674
rect 1407 670 1411 674
rect 1479 670 1483 674
rect 1575 670 1579 674
rect 1615 670 1619 674
rect 1727 670 1731 674
rect 1823 670 1827 674
rect 1863 670 1867 674
rect 1887 670 1891 674
rect 2055 670 2059 674
rect 2215 670 2219 674
rect 2247 670 2251 674
rect 2359 670 2363 674
rect 2439 670 2443 674
rect 2511 670 2515 674
rect 2631 670 2635 674
rect 2671 670 2675 674
rect 2815 670 2819 674
rect 2831 670 2835 674
rect 2991 670 2995 674
rect 3159 670 3163 674
rect 3327 670 3331 674
rect 3479 670 3483 674
rect 3575 670 3579 674
rect 111 598 115 602
rect 143 598 147 602
rect 303 598 307 602
rect 471 598 475 602
rect 487 598 491 602
rect 631 598 635 602
rect 671 598 675 602
rect 783 598 787 602
rect 847 598 851 602
rect 935 598 939 602
rect 1023 598 1027 602
rect 1079 598 1083 602
rect 1199 598 1203 602
rect 1215 598 1219 602
rect 1351 598 1355 602
rect 1375 598 1379 602
rect 1487 598 1491 602
rect 1559 598 1563 602
rect 1623 598 1627 602
rect 1735 598 1739 602
rect 1823 598 1827 602
rect 1863 598 1867 602
rect 2199 598 2203 602
rect 2223 598 2227 602
rect 2287 598 2291 602
rect 2367 598 2371 602
rect 2375 598 2379 602
rect 2463 598 2467 602
rect 2519 598 2523 602
rect 2567 598 2571 602
rect 2679 598 2683 602
rect 2815 598 2819 602
rect 2839 598 2843 602
rect 2975 598 2979 602
rect 2999 598 3003 602
rect 3143 598 3147 602
rect 3167 598 3171 602
rect 3327 598 3331 602
rect 3335 598 3339 602
rect 3487 598 3491 602
rect 3575 598 3579 602
rect 111 526 115 530
rect 135 526 139 530
rect 295 526 299 530
rect 303 526 307 530
rect 479 526 483 530
rect 495 526 499 530
rect 663 526 667 530
rect 679 526 683 530
rect 839 526 843 530
rect 863 526 867 530
rect 1015 526 1019 530
rect 1031 526 1035 530
rect 1191 526 1195 530
rect 1351 526 1355 530
rect 1367 526 1371 530
rect 1503 526 1507 530
rect 1551 526 1555 530
rect 1663 526 1667 530
rect 1727 526 1731 530
rect 1823 526 1827 530
rect 1863 526 1867 530
rect 2191 526 2195 530
rect 2279 526 2283 530
rect 2303 526 2307 530
rect 2367 526 2371 530
rect 2399 526 2403 530
rect 2455 526 2459 530
rect 2503 526 2507 530
rect 2559 526 2563 530
rect 2607 526 2611 530
rect 2671 526 2675 530
rect 2719 526 2723 530
rect 2807 526 2811 530
rect 2839 526 2843 530
rect 2967 526 2971 530
rect 3095 526 3099 530
rect 3135 526 3139 530
rect 3223 526 3227 530
rect 3319 526 3323 530
rect 3351 526 3355 530
rect 3479 526 3483 530
rect 3575 526 3579 530
rect 111 454 115 458
rect 143 454 147 458
rect 303 454 307 458
rect 311 454 315 458
rect 495 454 499 458
rect 503 454 507 458
rect 687 454 691 458
rect 871 454 875 458
rect 879 454 883 458
rect 1039 454 1043 458
rect 1055 454 1059 458
rect 1199 454 1203 458
rect 1223 454 1227 458
rect 1359 454 1363 458
rect 1391 454 1395 458
rect 1511 454 1515 458
rect 1559 454 1563 458
rect 1671 454 1675 458
rect 1727 454 1731 458
rect 1823 454 1827 458
rect 1863 458 1867 462
rect 2239 458 2243 462
rect 2311 458 2315 462
rect 2327 458 2331 462
rect 2407 458 2411 462
rect 2431 458 2435 462
rect 2511 458 2515 462
rect 2559 458 2563 462
rect 2615 458 2619 462
rect 2695 458 2699 462
rect 2727 458 2731 462
rect 2847 458 2851 462
rect 2975 458 2979 462
rect 2999 458 3003 462
rect 3103 458 3107 462
rect 3159 458 3163 462
rect 3231 458 3235 462
rect 3327 458 3331 462
rect 3359 458 3363 462
rect 3487 458 3491 462
rect 3575 458 3579 462
rect 111 386 115 390
rect 135 386 139 390
rect 263 386 267 390
rect 295 386 299 390
rect 423 386 427 390
rect 487 386 491 390
rect 591 386 595 390
rect 679 386 683 390
rect 767 386 771 390
rect 871 386 875 390
rect 935 386 939 390
rect 1047 386 1051 390
rect 1103 386 1107 390
rect 1215 386 1219 390
rect 1263 386 1267 390
rect 1383 386 1387 390
rect 1423 386 1427 390
rect 1551 386 1555 390
rect 1583 386 1587 390
rect 1719 386 1723 390
rect 1727 386 1731 390
rect 1823 386 1827 390
rect 1863 390 1867 394
rect 2183 390 2187 394
rect 2231 390 2235 394
rect 2287 390 2291 394
rect 2319 390 2323 394
rect 2399 390 2403 394
rect 2423 390 2427 394
rect 2527 390 2531 394
rect 2551 390 2555 394
rect 2671 390 2675 394
rect 2687 390 2691 394
rect 2815 390 2819 394
rect 2839 390 2843 394
rect 2967 390 2971 394
rect 2991 390 2995 394
rect 3127 390 3131 394
rect 3151 390 3155 394
rect 3295 390 3299 394
rect 3319 390 3323 394
rect 3463 390 3467 394
rect 3479 390 3483 394
rect 3575 390 3579 394
rect 111 318 115 322
rect 143 318 147 322
rect 215 318 219 322
rect 271 318 275 322
rect 351 318 355 322
rect 431 318 435 322
rect 495 318 499 322
rect 599 318 603 322
rect 639 318 643 322
rect 775 318 779 322
rect 791 318 795 322
rect 935 318 939 322
rect 943 318 947 322
rect 1079 318 1083 322
rect 1111 318 1115 322
rect 1223 318 1227 322
rect 1271 318 1275 322
rect 1359 318 1363 322
rect 1431 318 1435 322
rect 1487 318 1491 322
rect 1591 318 1595 322
rect 1623 318 1627 322
rect 1735 318 1739 322
rect 1823 318 1827 322
rect 1863 314 1867 318
rect 1895 314 1899 318
rect 2087 314 2091 318
rect 2191 314 2195 318
rect 2295 314 2299 318
rect 2303 314 2307 318
rect 2407 314 2411 318
rect 2511 314 2515 318
rect 2535 314 2539 318
rect 2679 314 2683 318
rect 2711 314 2715 318
rect 2823 314 2827 318
rect 2903 314 2907 318
rect 2975 314 2979 318
rect 3095 314 3099 318
rect 3135 314 3139 318
rect 3295 314 3299 318
rect 3303 314 3307 318
rect 3471 314 3475 318
rect 3487 314 3491 318
rect 3575 314 3579 318
rect 111 242 115 246
rect 207 242 211 246
rect 231 242 235 246
rect 343 242 347 246
rect 359 242 363 246
rect 487 242 491 246
rect 623 242 627 246
rect 631 242 635 246
rect 759 242 763 246
rect 783 242 787 246
rect 895 242 899 246
rect 927 242 931 246
rect 1031 242 1035 246
rect 1071 242 1075 246
rect 1159 242 1163 246
rect 1215 242 1219 246
rect 1295 242 1299 246
rect 1351 242 1355 246
rect 1431 242 1435 246
rect 1479 242 1483 246
rect 1615 242 1619 246
rect 1727 242 1731 246
rect 1823 242 1827 246
rect 1863 246 1867 250
rect 1887 246 1891 250
rect 1999 246 2003 250
rect 2079 246 2083 250
rect 2143 246 2147 250
rect 2295 246 2299 250
rect 2455 246 2459 250
rect 2503 246 2507 250
rect 2615 246 2619 250
rect 2703 246 2707 250
rect 2783 246 2787 250
rect 2895 246 2899 250
rect 2951 246 2955 250
rect 3087 246 3091 250
rect 3127 246 3131 250
rect 3287 246 3291 250
rect 3311 246 3315 250
rect 3479 246 3483 250
rect 3575 246 3579 250
rect 111 150 115 154
rect 175 150 179 154
rect 239 150 243 154
rect 263 150 267 154
rect 351 150 355 154
rect 367 150 371 154
rect 439 150 443 154
rect 495 150 499 154
rect 527 150 531 154
rect 615 150 619 154
rect 631 150 635 154
rect 703 150 707 154
rect 767 150 771 154
rect 791 150 795 154
rect 879 150 883 154
rect 903 150 907 154
rect 967 150 971 154
rect 1039 150 1043 154
rect 1055 150 1059 154
rect 1143 150 1147 154
rect 1167 150 1171 154
rect 1231 150 1235 154
rect 1303 150 1307 154
rect 1319 150 1323 154
rect 1407 150 1411 154
rect 1439 150 1443 154
rect 1503 150 1507 154
rect 1823 150 1827 154
rect 1863 150 1867 154
rect 1895 150 1899 154
rect 1983 150 1987 154
rect 2007 150 2011 154
rect 2071 150 2075 154
rect 2151 150 2155 154
rect 2159 150 2163 154
rect 2247 150 2251 154
rect 2303 150 2307 154
rect 2335 150 2339 154
rect 2439 150 2443 154
rect 2463 150 2467 154
rect 2543 150 2547 154
rect 2623 150 2627 154
rect 2647 150 2651 154
rect 2743 150 2747 154
rect 2791 150 2795 154
rect 2839 150 2843 154
rect 2935 150 2939 154
rect 2959 150 2963 154
rect 3031 150 3035 154
rect 3127 150 3131 154
rect 3135 150 3139 154
rect 3223 150 3227 154
rect 3311 150 3315 154
rect 3319 150 3323 154
rect 3399 150 3403 154
rect 3487 150 3491 154
rect 3575 150 3579 154
rect 111 82 115 86
rect 167 82 171 86
rect 255 82 259 86
rect 343 82 347 86
rect 431 82 435 86
rect 519 82 523 86
rect 607 82 611 86
rect 695 82 699 86
rect 783 82 787 86
rect 871 82 875 86
rect 959 82 963 86
rect 1047 82 1051 86
rect 1135 82 1139 86
rect 1223 82 1227 86
rect 1311 82 1315 86
rect 1399 82 1403 86
rect 1495 82 1499 86
rect 1823 82 1827 86
rect 1863 82 1867 86
rect 1887 82 1891 86
rect 1975 82 1979 86
rect 2063 82 2067 86
rect 2151 82 2155 86
rect 2239 82 2243 86
rect 2327 82 2331 86
rect 2431 82 2435 86
rect 2535 82 2539 86
rect 2639 82 2643 86
rect 2735 82 2739 86
rect 2831 82 2835 86
rect 2927 82 2931 86
rect 3023 82 3027 86
rect 3119 82 3123 86
rect 3215 82 3219 86
rect 3303 82 3307 86
rect 3391 82 3395 86
rect 3479 82 3483 86
rect 3575 82 3579 86
<< m4 >>
rect 96 3645 97 3651
rect 103 3650 1847 3651
rect 103 3646 111 3650
rect 115 3646 239 3650
rect 243 3646 327 3650
rect 331 3646 415 3650
rect 419 3646 503 3650
rect 507 3646 591 3650
rect 595 3646 679 3650
rect 683 3646 1823 3650
rect 1827 3646 1847 3650
rect 103 3645 1847 3646
rect 1853 3645 1854 3651
rect 1834 3581 1835 3587
rect 1841 3586 3599 3587
rect 1841 3582 1863 3586
rect 1867 3582 1887 3586
rect 1891 3582 1975 3586
rect 1979 3582 2063 3586
rect 2067 3582 2151 3586
rect 2155 3582 2239 3586
rect 2243 3582 2327 3586
rect 2331 3582 2415 3586
rect 2419 3582 2503 3586
rect 2507 3582 2591 3586
rect 2595 3582 2679 3586
rect 2683 3582 2767 3586
rect 2771 3582 2855 3586
rect 2859 3582 2943 3586
rect 2947 3582 3031 3586
rect 3035 3582 3119 3586
rect 3123 3582 3207 3586
rect 3211 3582 3295 3586
rect 3299 3582 3575 3586
rect 3579 3582 3599 3586
rect 1841 3581 3599 3582
rect 3605 3581 3606 3587
rect 84 3569 85 3575
rect 91 3574 1835 3575
rect 91 3570 111 3574
rect 115 3570 231 3574
rect 235 3570 247 3574
rect 251 3570 319 3574
rect 323 3570 399 3574
rect 403 3570 407 3574
rect 411 3570 495 3574
rect 499 3570 543 3574
rect 547 3570 583 3574
rect 587 3570 671 3574
rect 675 3570 687 3574
rect 691 3570 823 3574
rect 827 3570 951 3574
rect 955 3570 1079 3574
rect 1083 3570 1199 3574
rect 1203 3570 1311 3574
rect 1315 3570 1423 3574
rect 1427 3570 1543 3574
rect 1547 3570 1823 3574
rect 1827 3570 1835 3574
rect 91 3569 1835 3570
rect 1841 3569 1842 3575
rect 1846 3510 3618 3511
rect 1846 3507 1863 3510
rect 96 3501 97 3507
rect 103 3506 1847 3507
rect 103 3502 111 3506
rect 115 3502 183 3506
rect 187 3502 255 3506
rect 259 3502 351 3506
rect 355 3502 407 3506
rect 411 3502 519 3506
rect 523 3502 551 3506
rect 555 3502 679 3506
rect 683 3502 695 3506
rect 699 3502 831 3506
rect 835 3502 959 3506
rect 963 3502 967 3506
rect 971 3502 1087 3506
rect 1091 3502 1095 3506
rect 1099 3502 1207 3506
rect 1211 3502 1215 3506
rect 1219 3502 1319 3506
rect 1323 3502 1335 3506
rect 1339 3502 1431 3506
rect 1435 3502 1455 3506
rect 1459 3502 1551 3506
rect 1555 3502 1575 3506
rect 1579 3502 1823 3506
rect 1827 3502 1847 3506
rect 103 3501 1847 3502
rect 1853 3506 1863 3507
rect 1867 3506 1895 3510
rect 1899 3506 1911 3510
rect 1915 3506 1983 3510
rect 1987 3506 2015 3510
rect 2019 3506 2071 3510
rect 2075 3506 2135 3510
rect 2139 3506 2159 3510
rect 2163 3506 2247 3510
rect 2251 3506 2263 3510
rect 2267 3506 2335 3510
rect 2339 3506 2391 3510
rect 2395 3506 2423 3510
rect 2427 3506 2511 3510
rect 2515 3506 2527 3510
rect 2531 3506 2599 3510
rect 2603 3506 2663 3510
rect 2667 3506 2687 3510
rect 2691 3506 2775 3510
rect 2779 3506 2799 3510
rect 2803 3506 2863 3510
rect 2867 3506 2943 3510
rect 2947 3506 2951 3510
rect 2955 3506 3039 3510
rect 3043 3506 3087 3510
rect 3091 3506 3127 3510
rect 3131 3506 3215 3510
rect 3219 3506 3303 3510
rect 3307 3506 3575 3510
rect 3579 3506 3618 3510
rect 1853 3505 3618 3506
rect 1853 3501 1854 3505
rect 84 3433 85 3439
rect 91 3438 1835 3439
rect 91 3434 111 3438
rect 115 3434 135 3438
rect 139 3434 175 3438
rect 179 3434 255 3438
rect 259 3434 343 3438
rect 347 3434 415 3438
rect 419 3434 511 3438
rect 515 3434 583 3438
rect 587 3434 671 3438
rect 675 3434 759 3438
rect 763 3434 823 3438
rect 827 3434 935 3438
rect 939 3434 959 3438
rect 963 3434 1087 3438
rect 1091 3434 1111 3438
rect 1115 3434 1207 3438
rect 1211 3434 1295 3438
rect 1299 3434 1327 3438
rect 1331 3434 1447 3438
rect 1451 3434 1479 3438
rect 1483 3434 1567 3438
rect 1571 3434 1823 3438
rect 1827 3434 1835 3438
rect 91 3433 1835 3434
rect 1841 3435 1842 3439
rect 1841 3434 3606 3435
rect 1841 3433 1863 3434
rect 1834 3430 1863 3433
rect 1867 3430 1903 3434
rect 1907 3430 1911 3434
rect 1915 3430 2007 3434
rect 2011 3430 2071 3434
rect 2075 3430 2127 3434
rect 2131 3430 2223 3434
rect 2227 3430 2255 3434
rect 2259 3430 2367 3434
rect 2371 3430 2383 3434
rect 2387 3430 2503 3434
rect 2507 3430 2519 3434
rect 2523 3430 2631 3434
rect 2635 3430 2655 3434
rect 2659 3430 2759 3434
rect 2763 3430 2791 3434
rect 2795 3430 2887 3434
rect 2891 3430 2935 3434
rect 2939 3430 3023 3434
rect 3027 3430 3079 3434
rect 3083 3430 3575 3434
rect 3579 3430 3606 3434
rect 1834 3429 3606 3430
rect 96 3357 97 3363
rect 103 3362 1847 3363
rect 103 3358 111 3362
rect 115 3358 143 3362
rect 147 3358 207 3362
rect 211 3358 263 3362
rect 267 3358 367 3362
rect 371 3358 423 3362
rect 427 3358 535 3362
rect 539 3358 591 3362
rect 595 3358 695 3362
rect 699 3358 767 3362
rect 771 3358 855 3362
rect 859 3358 943 3362
rect 947 3358 999 3362
rect 1003 3358 1119 3362
rect 1123 3358 1143 3362
rect 1147 3358 1279 3362
rect 1283 3358 1303 3362
rect 1307 3358 1415 3362
rect 1419 3358 1487 3362
rect 1491 3358 1559 3362
rect 1563 3358 1823 3362
rect 1827 3358 1847 3362
rect 103 3357 1847 3358
rect 1853 3362 3618 3363
rect 1853 3358 1863 3362
rect 1867 3358 1895 3362
rect 1899 3358 1919 3362
rect 1923 3358 2047 3362
rect 2051 3358 2079 3362
rect 2083 3358 2207 3362
rect 2211 3358 2231 3362
rect 2235 3358 2367 3362
rect 2371 3358 2375 3362
rect 2379 3358 2511 3362
rect 2515 3358 2535 3362
rect 2539 3358 2639 3362
rect 2643 3358 2703 3362
rect 2707 3358 2767 3362
rect 2771 3358 2879 3362
rect 2883 3358 2895 3362
rect 2899 3358 3031 3362
rect 3035 3358 3055 3362
rect 3059 3358 3575 3362
rect 3579 3358 3618 3362
rect 1853 3357 3618 3358
rect 84 3285 85 3291
rect 91 3290 1835 3291
rect 91 3286 111 3290
rect 115 3286 199 3290
rect 203 3286 255 3290
rect 259 3286 359 3290
rect 363 3286 375 3290
rect 379 3286 511 3290
rect 515 3286 527 3290
rect 531 3286 663 3290
rect 667 3286 687 3290
rect 691 3286 823 3290
rect 827 3286 847 3290
rect 851 3286 991 3290
rect 995 3286 1135 3290
rect 1139 3286 1167 3290
rect 1171 3286 1271 3290
rect 1275 3286 1343 3290
rect 1347 3286 1407 3290
rect 1411 3286 1519 3290
rect 1523 3286 1551 3290
rect 1555 3286 1823 3290
rect 1827 3286 1835 3290
rect 91 3285 1835 3286
rect 1841 3290 3606 3291
rect 1841 3286 1863 3290
rect 1867 3286 1887 3290
rect 1891 3286 2039 3290
rect 2043 3286 2063 3290
rect 2067 3286 2199 3290
rect 2203 3286 2263 3290
rect 2267 3286 2359 3290
rect 2363 3286 2455 3290
rect 2459 3286 2527 3290
rect 2531 3286 2639 3290
rect 2643 3286 2695 3290
rect 2699 3286 2815 3290
rect 2819 3286 2871 3290
rect 2875 3286 2983 3290
rect 2987 3286 3047 3290
rect 3051 3286 3151 3290
rect 3155 3286 3319 3290
rect 3323 3286 3479 3290
rect 3483 3286 3575 3290
rect 3579 3286 3606 3290
rect 1841 3285 3606 3286
rect 1846 3222 3618 3223
rect 1846 3219 1863 3222
rect 96 3213 97 3219
rect 103 3218 1847 3219
rect 103 3214 111 3218
rect 115 3214 263 3218
rect 267 3214 383 3218
rect 387 3214 431 3218
rect 435 3214 519 3218
rect 523 3214 551 3218
rect 555 3214 671 3218
rect 675 3214 799 3218
rect 803 3214 831 3218
rect 835 3214 935 3218
rect 939 3214 999 3218
rect 1003 3214 1079 3218
rect 1083 3214 1175 3218
rect 1179 3214 1231 3218
rect 1235 3214 1351 3218
rect 1355 3214 1383 3218
rect 1387 3214 1527 3218
rect 1531 3214 1535 3218
rect 1539 3214 1823 3218
rect 1827 3214 1847 3218
rect 103 3213 1847 3214
rect 1853 3218 1863 3219
rect 1867 3218 1895 3222
rect 1899 3218 2071 3222
rect 2075 3218 2087 3222
rect 2091 3218 2271 3222
rect 2275 3218 2303 3222
rect 2307 3218 2463 3222
rect 2467 3218 2511 3222
rect 2515 3218 2647 3222
rect 2651 3218 2703 3222
rect 2707 3218 2823 3222
rect 2827 3218 2879 3222
rect 2883 3218 2991 3222
rect 2995 3218 3039 3222
rect 3043 3218 3159 3222
rect 3163 3218 3199 3222
rect 3203 3218 3327 3222
rect 3331 3218 3351 3222
rect 3355 3218 3487 3222
rect 3491 3218 3575 3222
rect 3579 3218 3618 3222
rect 1853 3217 3618 3218
rect 1853 3213 1854 3217
rect 1834 3150 3606 3151
rect 1834 3147 1863 3150
rect 84 3141 85 3147
rect 91 3146 1835 3147
rect 91 3142 111 3146
rect 115 3142 423 3146
rect 427 3142 463 3146
rect 467 3142 543 3146
rect 547 3142 551 3146
rect 555 3142 639 3146
rect 643 3142 663 3146
rect 667 3142 735 3146
rect 739 3142 791 3146
rect 795 3142 847 3146
rect 851 3142 927 3146
rect 931 3142 967 3146
rect 971 3142 1071 3146
rect 1075 3142 1095 3146
rect 1099 3142 1223 3146
rect 1227 3142 1231 3146
rect 1235 3142 1375 3146
rect 1379 3142 1519 3146
rect 1523 3142 1527 3146
rect 1531 3142 1823 3146
rect 1827 3142 1835 3146
rect 91 3141 1835 3142
rect 1841 3146 1863 3147
rect 1867 3146 1887 3150
rect 1891 3146 2079 3150
rect 2083 3146 2295 3150
rect 2299 3146 2503 3150
rect 2507 3146 2695 3150
rect 2699 3146 2871 3150
rect 2875 3146 3031 3150
rect 3035 3146 3039 3150
rect 3043 3146 3191 3150
rect 3195 3146 3343 3150
rect 3347 3146 3479 3150
rect 3483 3146 3575 3150
rect 3579 3146 3606 3150
rect 1841 3145 3606 3146
rect 1841 3141 1842 3145
rect 96 3065 97 3071
rect 103 3070 1847 3071
rect 103 3066 111 3070
rect 115 3066 151 3070
rect 155 3066 239 3070
rect 243 3066 327 3070
rect 331 3066 415 3070
rect 419 3066 471 3070
rect 475 3066 503 3070
rect 507 3066 559 3070
rect 563 3066 591 3070
rect 595 3066 647 3070
rect 651 3066 679 3070
rect 683 3066 743 3070
rect 747 3066 767 3070
rect 771 3066 855 3070
rect 859 3066 943 3070
rect 947 3066 975 3070
rect 979 3066 1031 3070
rect 1035 3066 1103 3070
rect 1107 3066 1119 3070
rect 1123 3066 1207 3070
rect 1211 3066 1239 3070
rect 1243 3066 1295 3070
rect 1299 3066 1383 3070
rect 1387 3066 1471 3070
rect 1475 3066 1527 3070
rect 1531 3066 1559 3070
rect 1563 3066 1647 3070
rect 1651 3066 1735 3070
rect 1739 3066 1823 3070
rect 1827 3066 1847 3070
rect 103 3065 1847 3066
rect 1853 3070 3618 3071
rect 1853 3066 1863 3070
rect 1867 3066 1895 3070
rect 1899 3066 2087 3070
rect 2091 3066 2255 3070
rect 2259 3066 2303 3070
rect 2307 3066 2423 3070
rect 2427 3066 2511 3070
rect 2515 3066 2591 3070
rect 2595 3066 2703 3070
rect 2707 3066 2751 3070
rect 2755 3066 2879 3070
rect 2883 3066 2919 3070
rect 2923 3066 3047 3070
rect 3051 3066 3087 3070
rect 3091 3066 3199 3070
rect 3203 3066 3351 3070
rect 3355 3066 3487 3070
rect 3491 3066 3575 3070
rect 3579 3066 3618 3070
rect 1853 3065 3618 3066
rect 1834 2998 3606 2999
rect 1834 2995 1863 2998
rect 84 2989 85 2995
rect 91 2994 1835 2995
rect 91 2990 111 2994
rect 115 2990 143 2994
rect 147 2990 231 2994
rect 235 2990 319 2994
rect 323 2990 407 2994
rect 411 2990 495 2994
rect 499 2990 583 2994
rect 587 2990 671 2994
rect 675 2990 759 2994
rect 763 2990 847 2994
rect 851 2990 935 2994
rect 939 2990 1023 2994
rect 1027 2990 1111 2994
rect 1115 2990 1199 2994
rect 1203 2990 1287 2994
rect 1291 2990 1375 2994
rect 1379 2990 1407 2994
rect 1411 2990 1463 2994
rect 1467 2990 1519 2994
rect 1523 2990 1551 2994
rect 1555 2990 1631 2994
rect 1635 2990 1639 2994
rect 1643 2990 1727 2994
rect 1731 2990 1823 2994
rect 1827 2990 1835 2994
rect 91 2989 1835 2990
rect 1841 2994 1863 2995
rect 1867 2994 2239 2998
rect 2243 2994 2247 2998
rect 2251 2994 2415 2998
rect 2419 2994 2463 2998
rect 2467 2994 2583 2998
rect 2587 2994 2671 2998
rect 2675 2994 2743 2998
rect 2747 2994 2863 2998
rect 2867 2994 2911 2998
rect 2915 2994 3031 2998
rect 3035 2994 3079 2998
rect 3083 2994 3191 2998
rect 3195 2994 3343 2998
rect 3347 2994 3479 2998
rect 3483 2994 3575 2998
rect 3579 2994 3606 2998
rect 1841 2993 3606 2994
rect 1841 2989 1842 2993
rect 96 2921 97 2927
rect 103 2926 1847 2927
rect 103 2922 111 2926
rect 115 2922 1359 2926
rect 1363 2922 1415 2926
rect 1419 2922 1471 2926
rect 1475 2922 1527 2926
rect 1531 2922 1583 2926
rect 1587 2922 1639 2926
rect 1643 2922 1703 2926
rect 1707 2922 1735 2926
rect 1739 2922 1823 2926
rect 1827 2922 1847 2926
rect 103 2921 1847 2922
rect 1853 2921 1854 2927
rect 1846 2909 1847 2915
rect 1853 2914 3611 2915
rect 1853 2910 1863 2914
rect 1867 2910 2239 2914
rect 2243 2910 2247 2914
rect 2251 2910 2463 2914
rect 2467 2910 2471 2914
rect 2475 2910 2671 2914
rect 2675 2910 2679 2914
rect 2683 2910 2855 2914
rect 2859 2910 2871 2914
rect 2875 2910 3023 2914
rect 3027 2910 3039 2914
rect 3043 2910 3183 2914
rect 3187 2910 3199 2914
rect 3203 2910 3335 2914
rect 3339 2910 3351 2914
rect 3355 2910 3487 2914
rect 3491 2910 3575 2914
rect 3579 2910 3611 2914
rect 1853 2909 3611 2910
rect 3617 2909 3618 2915
rect 84 2849 85 2855
rect 91 2854 1835 2855
rect 91 2850 111 2854
rect 115 2850 135 2854
rect 139 2850 223 2854
rect 227 2850 311 2854
rect 315 2850 399 2854
rect 403 2850 487 2854
rect 491 2850 599 2854
rect 603 2850 727 2854
rect 731 2850 863 2854
rect 867 2850 999 2854
rect 1003 2850 1135 2854
rect 1139 2850 1263 2854
rect 1267 2850 1351 2854
rect 1355 2850 1383 2854
rect 1387 2850 1463 2854
rect 1467 2850 1503 2854
rect 1507 2850 1575 2854
rect 1579 2850 1623 2854
rect 1627 2850 1695 2854
rect 1699 2850 1727 2854
rect 1731 2850 1823 2854
rect 1827 2850 1835 2854
rect 91 2849 1835 2850
rect 1841 2849 1842 2855
rect 1834 2837 1835 2843
rect 1841 2842 3599 2843
rect 1841 2838 1863 2842
rect 1867 2838 1895 2842
rect 1899 2838 1983 2842
rect 1987 2838 2071 2842
rect 2075 2838 2159 2842
rect 2163 2838 2231 2842
rect 2235 2838 2247 2842
rect 2251 2838 2335 2842
rect 2339 2838 2423 2842
rect 2427 2838 2455 2842
rect 2459 2838 2511 2842
rect 2515 2838 2599 2842
rect 2603 2838 2663 2842
rect 2667 2838 2687 2842
rect 2691 2838 2791 2842
rect 2795 2838 2847 2842
rect 2851 2838 2903 2842
rect 2907 2838 3015 2842
rect 3019 2838 3031 2842
rect 3035 2838 3175 2842
rect 3179 2838 3327 2842
rect 3331 2838 3479 2842
rect 3483 2838 3575 2842
rect 3579 2838 3599 2842
rect 1841 2837 3599 2838
rect 3605 2837 3606 2843
rect 96 2781 97 2787
rect 103 2786 1847 2787
rect 103 2782 111 2786
rect 115 2782 143 2786
rect 147 2782 191 2786
rect 195 2782 231 2786
rect 235 2782 295 2786
rect 299 2782 319 2786
rect 323 2782 407 2786
rect 411 2782 415 2786
rect 419 2782 495 2786
rect 499 2782 551 2786
rect 555 2782 607 2786
rect 611 2782 687 2786
rect 691 2782 735 2786
rect 739 2782 823 2786
rect 827 2782 871 2786
rect 875 2782 959 2786
rect 963 2782 1007 2786
rect 1011 2782 1087 2786
rect 1091 2782 1143 2786
rect 1147 2782 1207 2786
rect 1211 2782 1271 2786
rect 1275 2782 1319 2786
rect 1323 2782 1391 2786
rect 1395 2782 1431 2786
rect 1435 2782 1511 2786
rect 1515 2782 1535 2786
rect 1539 2782 1631 2786
rect 1635 2782 1647 2786
rect 1651 2782 1735 2786
rect 1739 2782 1823 2786
rect 1827 2782 1847 2786
rect 103 2781 1847 2782
rect 1853 2781 1854 2787
rect 1846 2757 1847 2763
rect 1853 2762 3611 2763
rect 1853 2758 1863 2762
rect 1867 2758 1903 2762
rect 1907 2758 1991 2762
rect 1995 2758 2047 2762
rect 2051 2758 2079 2762
rect 2083 2758 2167 2762
rect 2171 2758 2255 2762
rect 2259 2758 2295 2762
rect 2299 2758 2343 2762
rect 2347 2758 2431 2762
rect 2435 2758 2447 2762
rect 2451 2758 2519 2762
rect 2523 2758 2607 2762
rect 2611 2758 2623 2762
rect 2627 2758 2695 2762
rect 2699 2758 2799 2762
rect 2803 2758 2823 2762
rect 2827 2758 2911 2762
rect 2915 2758 3039 2762
rect 3043 2758 3183 2762
rect 3187 2758 3271 2762
rect 3275 2758 3335 2762
rect 3339 2758 3487 2762
rect 3491 2758 3575 2762
rect 3579 2758 3611 2762
rect 1853 2757 3611 2758
rect 3617 2757 3618 2763
rect 84 2705 85 2711
rect 91 2710 1835 2711
rect 91 2706 111 2710
rect 115 2706 167 2710
rect 171 2706 183 2710
rect 187 2706 279 2710
rect 283 2706 287 2710
rect 291 2706 391 2710
rect 395 2706 407 2710
rect 411 2706 503 2710
rect 507 2706 543 2710
rect 547 2706 615 2710
rect 619 2706 679 2710
rect 683 2706 815 2710
rect 819 2706 951 2710
rect 955 2706 1079 2710
rect 1083 2706 1199 2710
rect 1203 2706 1311 2710
rect 1315 2706 1423 2710
rect 1427 2706 1527 2710
rect 1531 2706 1639 2710
rect 1643 2706 1727 2710
rect 1731 2706 1823 2710
rect 1827 2706 1835 2710
rect 91 2705 1835 2706
rect 1841 2705 1842 2711
rect 1834 2689 1835 2695
rect 1841 2694 3599 2695
rect 1841 2690 1863 2694
rect 1867 2690 1943 2694
rect 1947 2690 2039 2694
rect 2043 2690 2055 2694
rect 2059 2690 2159 2694
rect 2163 2690 2167 2694
rect 2171 2690 2287 2694
rect 2291 2690 2407 2694
rect 2411 2690 2439 2694
rect 2443 2690 2519 2694
rect 2523 2690 2615 2694
rect 2619 2690 2631 2694
rect 2635 2690 2735 2694
rect 2739 2690 2815 2694
rect 2819 2690 2847 2694
rect 2851 2690 2959 2694
rect 2963 2690 3031 2694
rect 3035 2690 3071 2694
rect 3075 2690 3263 2694
rect 3267 2690 3479 2694
rect 3483 2690 3575 2694
rect 3579 2690 3599 2694
rect 1841 2689 3599 2690
rect 3605 2689 3606 2695
rect 96 2621 97 2627
rect 103 2626 1847 2627
rect 103 2622 111 2626
rect 115 2622 175 2626
rect 179 2622 223 2626
rect 227 2622 287 2626
rect 291 2622 351 2626
rect 355 2622 399 2626
rect 403 2622 495 2626
rect 499 2622 511 2626
rect 515 2622 623 2626
rect 627 2622 663 2626
rect 667 2622 839 2626
rect 843 2622 1023 2626
rect 1027 2622 1215 2626
rect 1219 2622 1407 2626
rect 1411 2622 1607 2626
rect 1611 2622 1823 2626
rect 1827 2622 1847 2626
rect 103 2621 1847 2622
rect 1853 2623 1854 2627
rect 1853 2622 3618 2623
rect 1853 2621 1863 2622
rect 1846 2618 1863 2621
rect 1867 2618 1895 2622
rect 1899 2618 1951 2622
rect 1955 2618 2063 2622
rect 2067 2618 2071 2622
rect 2075 2618 2175 2622
rect 2179 2618 2263 2622
rect 2267 2618 2295 2622
rect 2299 2618 2415 2622
rect 2419 2618 2463 2622
rect 2467 2618 2527 2622
rect 2531 2618 2639 2622
rect 2643 2618 2663 2622
rect 2667 2618 2743 2622
rect 2747 2618 2855 2622
rect 2859 2618 2871 2622
rect 2875 2618 2967 2622
rect 2971 2618 3079 2622
rect 3083 2618 3295 2622
rect 3299 2618 3487 2622
rect 3491 2618 3575 2622
rect 3579 2618 3618 2622
rect 1846 2617 3618 2618
rect 84 2553 85 2559
rect 91 2558 1835 2559
rect 91 2554 111 2558
rect 115 2554 215 2558
rect 219 2554 271 2558
rect 275 2554 343 2558
rect 347 2554 471 2558
rect 475 2554 487 2558
rect 491 2554 655 2558
rect 659 2554 671 2558
rect 675 2554 831 2558
rect 835 2554 855 2558
rect 859 2554 1015 2558
rect 1019 2554 1023 2558
rect 1027 2554 1175 2558
rect 1179 2554 1207 2558
rect 1211 2554 1319 2558
rect 1323 2554 1399 2558
rect 1403 2554 1455 2558
rect 1459 2554 1591 2558
rect 1595 2554 1599 2558
rect 1603 2554 1727 2558
rect 1731 2554 1823 2558
rect 1827 2554 1835 2558
rect 91 2553 1835 2554
rect 1841 2555 1842 2559
rect 1841 2554 3606 2555
rect 1841 2553 1863 2554
rect 1834 2550 1863 2553
rect 1867 2550 1887 2554
rect 1891 2550 2039 2554
rect 2043 2550 2063 2554
rect 2067 2550 2215 2554
rect 2219 2550 2255 2554
rect 2259 2550 2399 2554
rect 2403 2550 2455 2554
rect 2459 2550 2575 2554
rect 2579 2550 2655 2554
rect 2659 2550 2743 2554
rect 2747 2550 2863 2554
rect 2867 2550 2903 2554
rect 2907 2550 3055 2554
rect 3059 2550 3071 2554
rect 3075 2550 3199 2554
rect 3203 2550 3287 2554
rect 3291 2550 3343 2554
rect 3347 2550 3479 2554
rect 3483 2550 3575 2554
rect 3579 2550 3606 2554
rect 1834 2549 3606 2550
rect 96 2481 97 2487
rect 103 2486 1847 2487
rect 103 2482 111 2486
rect 115 2482 183 2486
rect 187 2482 279 2486
rect 283 2482 319 2486
rect 323 2482 463 2486
rect 467 2482 479 2486
rect 483 2482 607 2486
rect 611 2482 679 2486
rect 683 2482 743 2486
rect 747 2482 863 2486
rect 867 2482 879 2486
rect 883 2482 1007 2486
rect 1011 2482 1031 2486
rect 1035 2482 1127 2486
rect 1131 2482 1183 2486
rect 1187 2482 1239 2486
rect 1243 2482 1327 2486
rect 1331 2482 1343 2486
rect 1347 2482 1447 2486
rect 1451 2482 1463 2486
rect 1467 2482 1551 2486
rect 1555 2482 1599 2486
rect 1603 2482 1647 2486
rect 1651 2482 1735 2486
rect 1739 2482 1823 2486
rect 1827 2482 1847 2486
rect 103 2481 1847 2482
rect 1853 2486 3618 2487
rect 1853 2482 1863 2486
rect 1867 2482 1895 2486
rect 1899 2482 1991 2486
rect 1995 2482 2047 2486
rect 2051 2482 2127 2486
rect 2131 2482 2223 2486
rect 2227 2482 2279 2486
rect 2283 2482 2407 2486
rect 2411 2482 2439 2486
rect 2443 2482 2583 2486
rect 2587 2482 2599 2486
rect 2603 2482 2751 2486
rect 2755 2482 2767 2486
rect 2771 2482 2911 2486
rect 2915 2482 2943 2486
rect 2947 2482 3063 2486
rect 3067 2482 3119 2486
rect 3123 2482 3207 2486
rect 3211 2482 3295 2486
rect 3299 2482 3351 2486
rect 3355 2482 3471 2486
rect 3475 2482 3487 2486
rect 3491 2482 3575 2486
rect 3579 2482 3618 2486
rect 1853 2481 3618 2482
rect 84 2405 85 2411
rect 91 2410 1835 2411
rect 91 2406 111 2410
rect 115 2406 151 2410
rect 155 2406 175 2410
rect 179 2406 311 2410
rect 315 2406 319 2410
rect 323 2406 455 2410
rect 459 2406 479 2410
rect 483 2406 599 2410
rect 603 2406 639 2410
rect 643 2406 735 2410
rect 739 2406 783 2410
rect 787 2406 871 2410
rect 875 2406 919 2410
rect 923 2406 999 2410
rect 1003 2406 1047 2410
rect 1051 2406 1119 2410
rect 1123 2406 1175 2410
rect 1179 2406 1231 2410
rect 1235 2406 1303 2410
rect 1307 2406 1335 2410
rect 1339 2406 1431 2410
rect 1435 2406 1439 2410
rect 1443 2406 1543 2410
rect 1547 2406 1639 2410
rect 1643 2406 1727 2410
rect 1731 2406 1823 2410
rect 1827 2406 1835 2410
rect 91 2405 1835 2406
rect 1841 2410 3606 2411
rect 1841 2406 1863 2410
rect 1867 2406 1887 2410
rect 1891 2406 1983 2410
rect 1987 2406 2119 2410
rect 2123 2406 2271 2410
rect 2275 2406 2351 2410
rect 2355 2406 2431 2410
rect 2435 2406 2503 2410
rect 2507 2406 2591 2410
rect 2595 2406 2655 2410
rect 2659 2406 2759 2410
rect 2763 2406 2807 2410
rect 2811 2406 2935 2410
rect 2939 2406 2967 2410
rect 2971 2406 3111 2410
rect 3115 2406 3135 2410
rect 3139 2406 3287 2410
rect 3291 2406 3303 2410
rect 3307 2406 3463 2410
rect 3467 2406 3471 2410
rect 3475 2406 3575 2410
rect 3579 2406 3606 2410
rect 1841 2405 3606 2406
rect 96 2333 97 2339
rect 103 2338 1847 2339
rect 103 2334 111 2338
rect 115 2334 143 2338
rect 147 2334 159 2338
rect 163 2334 263 2338
rect 267 2334 327 2338
rect 331 2334 407 2338
rect 411 2334 487 2338
rect 491 2334 543 2338
rect 547 2334 647 2338
rect 651 2334 679 2338
rect 683 2334 791 2338
rect 795 2334 807 2338
rect 811 2334 927 2338
rect 931 2334 1039 2338
rect 1043 2334 1055 2338
rect 1059 2334 1159 2338
rect 1163 2334 1183 2338
rect 1187 2334 1279 2338
rect 1283 2334 1311 2338
rect 1315 2334 1439 2338
rect 1443 2334 1823 2338
rect 1827 2334 1847 2338
rect 103 2333 1847 2334
rect 1853 2338 3618 2339
rect 1853 2334 1863 2338
rect 1867 2334 2351 2338
rect 2355 2334 2359 2338
rect 2363 2334 2447 2338
rect 2451 2334 2511 2338
rect 2515 2334 2559 2338
rect 2563 2334 2663 2338
rect 2667 2334 2703 2338
rect 2707 2334 2815 2338
rect 2819 2334 2879 2338
rect 2883 2334 2975 2338
rect 2979 2334 3079 2338
rect 3083 2334 3143 2338
rect 3147 2334 3287 2338
rect 3291 2334 3311 2338
rect 3315 2334 3479 2338
rect 3483 2334 3487 2338
rect 3491 2334 3575 2338
rect 3579 2334 3618 2338
rect 1853 2333 3618 2334
rect 84 2265 85 2271
rect 91 2270 1835 2271
rect 91 2266 111 2270
rect 115 2266 135 2270
rect 139 2266 231 2270
rect 235 2266 255 2270
rect 259 2266 351 2270
rect 355 2266 399 2270
rect 403 2266 471 2270
rect 475 2266 535 2270
rect 539 2266 591 2270
rect 595 2266 671 2270
rect 675 2266 711 2270
rect 715 2266 799 2270
rect 803 2266 823 2270
rect 827 2266 919 2270
rect 923 2266 935 2270
rect 939 2266 1031 2270
rect 1035 2266 1055 2270
rect 1059 2266 1151 2270
rect 1155 2266 1175 2270
rect 1179 2266 1271 2270
rect 1275 2266 1823 2270
rect 1827 2266 1835 2270
rect 91 2265 1835 2266
rect 1841 2270 3606 2271
rect 1841 2266 1863 2270
rect 1867 2266 2335 2270
rect 2339 2266 2343 2270
rect 2347 2266 2439 2270
rect 2443 2266 2447 2270
rect 2451 2266 2551 2270
rect 2555 2266 2583 2270
rect 2587 2266 2695 2270
rect 2699 2266 2735 2270
rect 2739 2266 2871 2270
rect 2875 2266 2911 2270
rect 2915 2266 3071 2270
rect 3075 2266 3103 2270
rect 3107 2266 3279 2270
rect 3283 2266 3303 2270
rect 3307 2266 3479 2270
rect 3483 2266 3575 2270
rect 3579 2266 3606 2270
rect 1841 2265 3606 2266
rect 1846 2202 3618 2203
rect 1846 2199 1863 2202
rect 96 2193 97 2199
rect 103 2198 1847 2199
rect 103 2194 111 2198
rect 115 2194 143 2198
rect 147 2194 239 2198
rect 243 2194 247 2198
rect 251 2194 359 2198
rect 363 2194 383 2198
rect 387 2194 479 2198
rect 483 2194 519 2198
rect 523 2194 599 2198
rect 603 2194 655 2198
rect 659 2194 719 2198
rect 723 2194 783 2198
rect 787 2194 831 2198
rect 835 2194 911 2198
rect 915 2194 943 2198
rect 947 2194 1031 2198
rect 1035 2194 1063 2198
rect 1067 2194 1159 2198
rect 1163 2194 1183 2198
rect 1187 2194 1287 2198
rect 1291 2194 1823 2198
rect 1827 2194 1847 2198
rect 103 2193 1847 2194
rect 1853 2198 1863 2199
rect 1867 2198 2255 2202
rect 2259 2198 2343 2202
rect 2347 2198 2439 2202
rect 2443 2198 2455 2202
rect 2459 2198 2551 2202
rect 2555 2198 2591 2202
rect 2595 2198 2695 2202
rect 2699 2198 2743 2202
rect 2747 2198 2871 2202
rect 2875 2198 2919 2202
rect 2923 2198 3071 2202
rect 3075 2198 3111 2202
rect 3115 2198 3287 2202
rect 3291 2198 3311 2202
rect 3315 2198 3487 2202
rect 3491 2198 3575 2202
rect 3579 2198 3618 2202
rect 1853 2197 3618 2198
rect 1853 2193 1854 2197
rect 1834 2126 3606 2127
rect 1834 2123 1863 2126
rect 84 2117 85 2123
rect 91 2122 1835 2123
rect 91 2118 111 2122
rect 115 2118 135 2122
rect 139 2118 231 2122
rect 235 2118 239 2122
rect 243 2118 359 2122
rect 363 2118 375 2122
rect 379 2118 479 2122
rect 483 2118 511 2122
rect 515 2118 599 2122
rect 603 2118 647 2122
rect 651 2118 719 2122
rect 723 2118 775 2122
rect 779 2118 831 2122
rect 835 2118 903 2122
rect 907 2118 943 2122
rect 947 2118 1023 2122
rect 1027 2118 1055 2122
rect 1059 2118 1151 2122
rect 1155 2118 1175 2122
rect 1179 2118 1279 2122
rect 1283 2118 1823 2122
rect 1827 2118 1835 2122
rect 91 2117 1835 2118
rect 1841 2122 1863 2123
rect 1867 2122 2151 2126
rect 2155 2122 2239 2126
rect 2243 2122 2247 2126
rect 2251 2122 2327 2126
rect 2331 2122 2335 2126
rect 2339 2122 2415 2126
rect 2419 2122 2431 2126
rect 2435 2122 2503 2126
rect 2507 2122 2543 2126
rect 2547 2122 2615 2126
rect 2619 2122 2687 2126
rect 2691 2122 2751 2126
rect 2755 2122 2863 2126
rect 2867 2122 2919 2126
rect 2923 2122 3063 2126
rect 3067 2122 3103 2126
rect 3107 2122 3279 2126
rect 3283 2122 3303 2126
rect 3307 2122 3479 2126
rect 3483 2122 3575 2126
rect 3579 2122 3606 2126
rect 1841 2121 3606 2122
rect 1841 2117 1842 2121
rect 1846 2049 1847 2055
rect 1853 2054 3611 2055
rect 1853 2050 1863 2054
rect 1867 2050 1999 2054
rect 2003 2050 2127 2054
rect 2131 2050 2159 2054
rect 2163 2050 2247 2054
rect 2251 2050 2255 2054
rect 2259 2050 2335 2054
rect 2339 2050 2399 2054
rect 2403 2050 2423 2054
rect 2427 2050 2511 2054
rect 2515 2050 2551 2054
rect 2555 2050 2623 2054
rect 2627 2050 2711 2054
rect 2715 2050 2759 2054
rect 2763 2050 2879 2054
rect 2883 2050 2927 2054
rect 2931 2050 3063 2054
rect 3067 2050 3111 2054
rect 3115 2050 3247 2054
rect 3251 2050 3311 2054
rect 3315 2050 3439 2054
rect 3443 2050 3487 2054
rect 3491 2050 3575 2054
rect 3579 2050 3611 2054
rect 1853 2049 3611 2050
rect 3617 2049 3618 2055
rect 96 2037 97 2043
rect 103 2042 1847 2043
rect 103 2038 111 2042
rect 115 2038 143 2042
rect 147 2038 167 2042
rect 171 2038 239 2042
rect 243 2038 311 2042
rect 315 2038 367 2042
rect 371 2038 447 2042
rect 451 2038 487 2042
rect 491 2038 575 2042
rect 579 2038 607 2042
rect 611 2038 695 2042
rect 699 2038 727 2042
rect 731 2038 807 2042
rect 811 2038 839 2042
rect 843 2038 911 2042
rect 915 2038 951 2042
rect 955 2038 1015 2042
rect 1019 2038 1063 2042
rect 1067 2038 1119 2042
rect 1123 2038 1183 2042
rect 1187 2038 1223 2042
rect 1227 2038 1327 2042
rect 1331 2038 1823 2042
rect 1827 2038 1847 2042
rect 103 2037 1847 2038
rect 1853 2037 1854 2043
rect 1834 1978 3606 1979
rect 1834 1975 1863 1978
rect 84 1969 85 1975
rect 91 1974 1835 1975
rect 91 1970 111 1974
rect 115 1970 159 1974
rect 163 1970 295 1974
rect 299 1970 303 1974
rect 307 1970 439 1974
rect 443 1970 567 1974
rect 571 1970 583 1974
rect 587 1970 687 1974
rect 691 1970 719 1974
rect 723 1970 799 1974
rect 803 1970 855 1974
rect 859 1970 903 1974
rect 907 1970 991 1974
rect 995 1970 1007 1974
rect 1011 1970 1111 1974
rect 1115 1970 1119 1974
rect 1123 1970 1215 1974
rect 1219 1970 1239 1974
rect 1243 1970 1319 1974
rect 1323 1970 1359 1974
rect 1363 1970 1479 1974
rect 1483 1970 1599 1974
rect 1603 1970 1823 1974
rect 1827 1970 1835 1974
rect 91 1969 1835 1970
rect 1841 1974 1863 1975
rect 1867 1974 1903 1978
rect 1907 1974 1991 1978
rect 1995 1974 2119 1978
rect 2123 1974 2159 1978
rect 2163 1974 2247 1978
rect 2251 1974 2391 1978
rect 2395 1974 2399 1978
rect 2403 1974 2543 1978
rect 2547 1974 2615 1978
rect 2619 1974 2703 1978
rect 2707 1974 2815 1978
rect 2819 1974 2871 1978
rect 2875 1974 2999 1978
rect 3003 1974 3055 1978
rect 3059 1974 3167 1978
rect 3171 1974 3239 1978
rect 3243 1974 3335 1978
rect 3339 1974 3431 1978
rect 3435 1974 3479 1978
rect 3483 1974 3575 1978
rect 3579 1974 3606 1978
rect 1841 1973 3606 1974
rect 1841 1969 1842 1973
rect 1846 1905 1847 1911
rect 1853 1910 3611 1911
rect 1853 1906 1863 1910
rect 1867 1906 1895 1910
rect 1899 1906 1911 1910
rect 1915 1906 1983 1910
rect 1987 1906 2071 1910
rect 2075 1906 2167 1910
rect 2171 1906 2295 1910
rect 2299 1906 2407 1910
rect 2411 1906 2447 1910
rect 2451 1906 2607 1910
rect 2611 1906 2623 1910
rect 2627 1906 2767 1910
rect 2771 1906 2823 1910
rect 2827 1906 2919 1910
rect 2923 1906 3007 1910
rect 3011 1906 3071 1910
rect 3075 1906 3175 1910
rect 3179 1906 3215 1910
rect 3219 1906 3343 1910
rect 3347 1906 3359 1910
rect 3363 1906 3487 1910
rect 3491 1906 3575 1910
rect 3579 1906 3611 1910
rect 1853 1905 3611 1906
rect 3617 1905 3618 1911
rect 96 1893 97 1899
rect 103 1898 1847 1899
rect 103 1894 111 1898
rect 115 1894 167 1898
rect 171 1894 223 1898
rect 227 1894 303 1898
rect 307 1894 447 1898
rect 451 1894 479 1898
rect 483 1894 591 1898
rect 595 1894 719 1898
rect 723 1894 727 1898
rect 731 1894 863 1898
rect 867 1894 935 1898
rect 939 1894 999 1898
rect 1003 1894 1127 1898
rect 1131 1894 1247 1898
rect 1251 1894 1295 1898
rect 1299 1894 1367 1898
rect 1371 1894 1455 1898
rect 1459 1894 1487 1898
rect 1491 1894 1607 1898
rect 1611 1894 1735 1898
rect 1739 1894 1823 1898
rect 1827 1894 1847 1898
rect 103 1893 1847 1894
rect 1853 1893 1854 1899
rect 1834 1833 1835 1839
rect 1841 1838 3599 1839
rect 1841 1834 1863 1838
rect 1867 1834 1887 1838
rect 1891 1834 1975 1838
rect 1979 1834 1999 1838
rect 2003 1834 2063 1838
rect 2067 1834 2159 1838
rect 2163 1834 2223 1838
rect 2227 1834 2287 1838
rect 2291 1834 2439 1838
rect 2443 1834 2599 1838
rect 2603 1834 2639 1838
rect 2643 1834 2759 1838
rect 2763 1834 2831 1838
rect 2835 1834 2911 1838
rect 2915 1834 3015 1838
rect 3019 1834 3063 1838
rect 3067 1834 3199 1838
rect 3203 1834 3207 1838
rect 3211 1834 3351 1838
rect 3355 1834 3391 1838
rect 3395 1834 3479 1838
rect 3483 1834 3575 1838
rect 3579 1834 3599 1838
rect 1841 1833 3599 1834
rect 3605 1833 3606 1839
rect 1834 1831 1842 1833
rect 84 1825 85 1831
rect 91 1830 1835 1831
rect 91 1826 111 1830
rect 115 1826 215 1830
rect 219 1826 247 1830
rect 251 1826 415 1830
rect 419 1826 471 1830
rect 475 1826 591 1830
rect 595 1826 711 1830
rect 715 1826 759 1830
rect 763 1826 927 1830
rect 931 1826 1079 1830
rect 1083 1826 1119 1830
rect 1123 1826 1223 1830
rect 1227 1826 1287 1830
rect 1291 1826 1359 1830
rect 1363 1826 1447 1830
rect 1451 1826 1487 1830
rect 1491 1826 1599 1830
rect 1603 1826 1615 1830
rect 1619 1826 1727 1830
rect 1731 1826 1823 1830
rect 1827 1826 1835 1830
rect 91 1825 1835 1826
rect 1841 1825 1842 1831
rect 1846 1761 1847 1767
rect 1853 1766 3611 1767
rect 1853 1762 1863 1766
rect 1867 1762 1943 1766
rect 1947 1762 2007 1766
rect 2011 1762 2087 1766
rect 2091 1762 2231 1766
rect 2235 1762 2247 1766
rect 2251 1762 2415 1766
rect 2419 1762 2447 1766
rect 2451 1762 2599 1766
rect 2603 1762 2647 1766
rect 2651 1762 2791 1766
rect 2795 1762 2839 1766
rect 2843 1762 2991 1766
rect 2995 1762 3023 1766
rect 3027 1762 3199 1766
rect 3203 1762 3207 1766
rect 3211 1762 3399 1766
rect 3403 1762 3415 1766
rect 3419 1762 3575 1766
rect 3579 1762 3611 1766
rect 1853 1761 3611 1762
rect 3617 1761 3618 1767
rect 1846 1759 1854 1761
rect 96 1753 97 1759
rect 103 1758 1847 1759
rect 103 1754 111 1758
rect 115 1754 255 1758
rect 259 1754 327 1758
rect 331 1754 423 1758
rect 427 1754 471 1758
rect 475 1754 599 1758
rect 603 1754 615 1758
rect 619 1754 767 1758
rect 771 1754 919 1758
rect 923 1754 935 1758
rect 939 1754 1071 1758
rect 1075 1754 1087 1758
rect 1091 1754 1223 1758
rect 1227 1754 1231 1758
rect 1235 1754 1367 1758
rect 1371 1754 1375 1758
rect 1379 1754 1495 1758
rect 1499 1754 1527 1758
rect 1531 1754 1623 1758
rect 1627 1754 1687 1758
rect 1691 1754 1735 1758
rect 1739 1754 1823 1758
rect 1827 1754 1847 1758
rect 103 1753 1847 1754
rect 1853 1753 1854 1759
rect 1834 1689 1835 1695
rect 1841 1694 3599 1695
rect 1841 1690 1863 1694
rect 1867 1690 1911 1694
rect 1915 1690 1935 1694
rect 1939 1690 2031 1694
rect 2035 1690 2079 1694
rect 2083 1690 2151 1694
rect 2155 1690 2239 1694
rect 2243 1690 2271 1694
rect 2275 1690 2399 1694
rect 2403 1690 2407 1694
rect 2411 1690 2543 1694
rect 2547 1690 2591 1694
rect 2595 1690 2695 1694
rect 2699 1690 2783 1694
rect 2787 1690 2863 1694
rect 2867 1690 2983 1694
rect 2987 1690 3047 1694
rect 3051 1690 3191 1694
rect 3195 1690 3239 1694
rect 3243 1690 3407 1694
rect 3411 1690 3431 1694
rect 3435 1690 3575 1694
rect 3579 1690 3599 1694
rect 1841 1689 3599 1690
rect 3605 1689 3606 1695
rect 1834 1687 1842 1689
rect 84 1681 85 1687
rect 91 1686 1835 1687
rect 91 1682 111 1686
rect 115 1682 311 1686
rect 315 1682 319 1686
rect 323 1682 447 1686
rect 451 1682 463 1686
rect 467 1682 591 1686
rect 595 1682 607 1686
rect 611 1682 735 1686
rect 739 1682 759 1686
rect 763 1682 887 1686
rect 891 1682 911 1686
rect 915 1682 1039 1686
rect 1043 1682 1063 1686
rect 1067 1682 1191 1686
rect 1195 1682 1215 1686
rect 1219 1682 1343 1686
rect 1347 1682 1367 1686
rect 1371 1682 1495 1686
rect 1499 1682 1519 1686
rect 1523 1682 1647 1686
rect 1651 1682 1679 1686
rect 1683 1682 1823 1686
rect 1827 1682 1835 1686
rect 91 1681 1835 1682
rect 1841 1681 1842 1687
rect 1846 1613 1847 1619
rect 1853 1618 3611 1619
rect 1853 1614 1863 1618
rect 1867 1614 1895 1618
rect 1899 1614 1919 1618
rect 1923 1614 2015 1618
rect 2019 1614 2039 1618
rect 2043 1614 2151 1618
rect 2155 1614 2159 1618
rect 2163 1614 2279 1618
rect 2283 1614 2287 1618
rect 2291 1614 2407 1618
rect 2411 1614 2431 1618
rect 2435 1614 2551 1618
rect 2555 1614 2583 1618
rect 2587 1614 2703 1618
rect 2707 1614 2743 1618
rect 2747 1614 2871 1618
rect 2875 1614 2911 1618
rect 2915 1614 3055 1618
rect 3059 1614 3095 1618
rect 3099 1614 3247 1618
rect 3251 1614 3279 1618
rect 3283 1614 3439 1618
rect 3443 1614 3471 1618
rect 3475 1614 3575 1618
rect 3579 1614 3611 1618
rect 1853 1613 3611 1614
rect 3617 1613 3618 1619
rect 1846 1611 1854 1613
rect 96 1605 97 1611
rect 103 1610 1847 1611
rect 103 1606 111 1610
rect 115 1606 223 1610
rect 227 1606 319 1610
rect 323 1606 351 1610
rect 355 1606 455 1610
rect 459 1606 487 1610
rect 491 1606 599 1610
rect 603 1606 623 1610
rect 627 1606 743 1610
rect 747 1606 759 1610
rect 763 1606 895 1610
rect 899 1606 903 1610
rect 907 1606 1047 1610
rect 1051 1606 1055 1610
rect 1059 1606 1199 1610
rect 1203 1606 1215 1610
rect 1219 1606 1351 1610
rect 1355 1606 1375 1610
rect 1379 1606 1503 1610
rect 1507 1606 1543 1610
rect 1547 1606 1655 1610
rect 1659 1606 1823 1610
rect 1827 1606 1847 1610
rect 103 1605 1847 1606
rect 1853 1605 1854 1611
rect 1834 1542 3606 1543
rect 1834 1539 1863 1542
rect 84 1533 85 1539
rect 91 1538 1835 1539
rect 91 1534 111 1538
rect 115 1534 135 1538
rect 139 1534 215 1538
rect 219 1534 271 1538
rect 275 1534 343 1538
rect 347 1534 423 1538
rect 427 1534 479 1538
rect 483 1534 583 1538
rect 587 1534 615 1538
rect 619 1534 735 1538
rect 739 1534 751 1538
rect 755 1534 887 1538
rect 891 1534 895 1538
rect 899 1534 1039 1538
rect 1043 1534 1047 1538
rect 1051 1534 1191 1538
rect 1195 1534 1207 1538
rect 1211 1534 1343 1538
rect 1347 1534 1367 1538
rect 1371 1534 1495 1538
rect 1499 1534 1535 1538
rect 1539 1534 1823 1538
rect 1827 1534 1835 1538
rect 91 1533 1835 1534
rect 1841 1538 1863 1539
rect 1867 1538 1887 1542
rect 1891 1538 2007 1542
rect 2011 1538 2023 1542
rect 2027 1538 2143 1542
rect 2147 1538 2183 1542
rect 2187 1538 2279 1542
rect 2283 1538 2343 1542
rect 2347 1538 2423 1542
rect 2427 1538 2503 1542
rect 2507 1538 2575 1542
rect 2579 1538 2663 1542
rect 2667 1538 2735 1542
rect 2739 1538 2823 1542
rect 2827 1538 2903 1542
rect 2907 1538 2983 1542
rect 2987 1538 3087 1542
rect 3091 1538 3151 1542
rect 3155 1538 3271 1542
rect 3275 1538 3319 1542
rect 3323 1538 3463 1542
rect 3467 1538 3479 1542
rect 3483 1538 3575 1542
rect 3579 1538 3606 1542
rect 1841 1537 3606 1538
rect 1841 1533 1842 1537
rect 1846 1466 3618 1467
rect 1846 1463 1863 1466
rect 96 1457 97 1463
rect 103 1462 1847 1463
rect 103 1458 111 1462
rect 115 1458 143 1462
rect 147 1458 263 1462
rect 267 1458 279 1462
rect 283 1458 399 1462
rect 403 1458 431 1462
rect 435 1458 535 1462
rect 539 1458 591 1462
rect 595 1458 663 1462
rect 667 1458 743 1462
rect 747 1458 791 1462
rect 795 1458 895 1462
rect 899 1458 911 1462
rect 915 1458 1023 1462
rect 1027 1458 1047 1462
rect 1051 1458 1143 1462
rect 1147 1458 1199 1462
rect 1203 1458 1263 1462
rect 1267 1458 1351 1462
rect 1355 1458 1383 1462
rect 1387 1458 1503 1462
rect 1507 1458 1631 1462
rect 1635 1458 1735 1462
rect 1739 1458 1823 1462
rect 1827 1458 1847 1462
rect 103 1457 1847 1458
rect 1853 1462 1863 1463
rect 1867 1462 1895 1466
rect 1899 1462 2031 1466
rect 2035 1462 2183 1466
rect 2187 1462 2191 1466
rect 2195 1462 2351 1466
rect 2355 1462 2359 1466
rect 2363 1462 2511 1466
rect 2515 1462 2527 1466
rect 2531 1462 2671 1466
rect 2675 1462 2687 1466
rect 2691 1462 2831 1466
rect 2835 1462 2847 1466
rect 2851 1462 2991 1466
rect 2995 1462 3007 1466
rect 3011 1462 3159 1466
rect 3163 1462 3175 1466
rect 3179 1462 3327 1466
rect 3331 1462 3343 1466
rect 3347 1462 3487 1466
rect 3491 1462 3575 1466
rect 3579 1462 3618 1466
rect 1853 1461 3618 1462
rect 1853 1457 1854 1461
rect 84 1389 85 1395
rect 91 1394 1835 1395
rect 91 1390 111 1394
rect 115 1390 135 1394
rect 139 1390 255 1394
rect 259 1390 327 1394
rect 331 1390 391 1394
rect 395 1390 527 1394
rect 531 1390 551 1394
rect 555 1390 655 1394
rect 659 1390 783 1394
rect 787 1390 903 1394
rect 907 1390 1015 1394
rect 1019 1390 1023 1394
rect 1027 1390 1135 1394
rect 1139 1390 1255 1394
rect 1259 1390 1263 1394
rect 1267 1390 1375 1394
rect 1379 1390 1495 1394
rect 1499 1390 1503 1394
rect 1507 1390 1623 1394
rect 1627 1390 1727 1394
rect 1731 1390 1823 1394
rect 1827 1390 1835 1394
rect 91 1389 1835 1390
rect 1841 1391 1842 1395
rect 1841 1390 3606 1391
rect 1841 1389 1863 1390
rect 1834 1386 1863 1389
rect 1867 1386 2079 1390
rect 2083 1386 2175 1390
rect 2179 1386 2263 1390
rect 2267 1386 2351 1390
rect 2355 1386 2439 1390
rect 2443 1386 2519 1390
rect 2523 1386 2615 1390
rect 2619 1386 2679 1390
rect 2683 1386 2783 1390
rect 2787 1386 2839 1390
rect 2843 1386 2935 1390
rect 2939 1386 2999 1390
rect 3003 1386 3079 1390
rect 3083 1386 3167 1390
rect 3171 1386 3223 1390
rect 3227 1386 3335 1390
rect 3339 1386 3359 1390
rect 3363 1386 3479 1390
rect 3483 1386 3575 1390
rect 3579 1386 3606 1390
rect 1834 1385 3606 1386
rect 1846 1322 3618 1323
rect 1846 1319 1863 1322
rect 96 1313 97 1319
rect 103 1318 1847 1319
rect 103 1314 111 1318
rect 115 1314 143 1318
rect 147 1314 327 1318
rect 331 1314 335 1318
rect 339 1314 527 1318
rect 531 1314 559 1318
rect 563 1314 719 1318
rect 723 1314 791 1318
rect 795 1314 903 1318
rect 907 1314 1031 1318
rect 1035 1314 1071 1318
rect 1075 1314 1231 1318
rect 1235 1314 1271 1318
rect 1275 1314 1383 1318
rect 1387 1314 1511 1318
rect 1515 1314 1535 1318
rect 1539 1314 1687 1318
rect 1691 1314 1735 1318
rect 1739 1314 1823 1318
rect 1827 1314 1847 1318
rect 103 1313 1847 1314
rect 1853 1318 1863 1319
rect 1867 1318 2087 1322
rect 2091 1318 2271 1322
rect 2275 1318 2311 1322
rect 2315 1318 2447 1322
rect 2451 1318 2519 1322
rect 2523 1318 2623 1322
rect 2627 1318 2711 1322
rect 2715 1318 2791 1322
rect 2795 1318 2887 1322
rect 2891 1318 2943 1322
rect 2947 1318 3047 1322
rect 3051 1318 3087 1322
rect 3091 1318 3199 1322
rect 3203 1318 3231 1322
rect 3235 1318 3351 1322
rect 3355 1318 3367 1322
rect 3371 1318 3487 1322
rect 3491 1318 3575 1322
rect 3579 1318 3618 1322
rect 1853 1317 3618 1318
rect 1853 1313 1854 1317
rect 1834 1250 3606 1251
rect 1834 1247 1863 1250
rect 84 1241 85 1247
rect 91 1246 1835 1247
rect 91 1242 111 1246
rect 115 1242 135 1246
rect 139 1242 295 1246
rect 299 1242 319 1246
rect 323 1242 479 1246
rect 483 1242 519 1246
rect 523 1242 655 1246
rect 659 1242 711 1246
rect 715 1242 815 1246
rect 819 1242 895 1246
rect 899 1242 967 1246
rect 971 1242 1063 1246
rect 1067 1242 1111 1246
rect 1115 1242 1223 1246
rect 1227 1242 1247 1246
rect 1251 1242 1375 1246
rect 1379 1242 1383 1246
rect 1387 1242 1527 1246
rect 1531 1242 1679 1246
rect 1683 1242 1823 1246
rect 1827 1242 1835 1246
rect 91 1241 1835 1242
rect 1841 1246 1863 1247
rect 1867 1246 1903 1250
rect 1907 1246 1991 1250
rect 1995 1246 2079 1250
rect 2083 1246 2095 1250
rect 2099 1246 2215 1250
rect 2219 1246 2303 1250
rect 2307 1246 2351 1250
rect 2355 1246 2487 1250
rect 2491 1246 2511 1250
rect 2515 1246 2631 1250
rect 2635 1246 2703 1250
rect 2707 1246 2775 1250
rect 2779 1246 2879 1250
rect 2883 1246 2919 1250
rect 2923 1246 3039 1250
rect 3043 1246 3063 1250
rect 3067 1246 3191 1250
rect 3195 1246 3207 1250
rect 3211 1246 3343 1250
rect 3347 1246 3351 1250
rect 3355 1246 3479 1250
rect 3483 1246 3575 1250
rect 3579 1246 3606 1250
rect 1841 1245 3606 1246
rect 1841 1241 1842 1245
rect 1846 1178 3618 1179
rect 1846 1175 1863 1178
rect 96 1169 97 1175
rect 103 1174 1847 1175
rect 103 1170 111 1174
rect 115 1170 143 1174
rect 147 1170 167 1174
rect 171 1170 303 1174
rect 307 1170 319 1174
rect 323 1170 471 1174
rect 475 1170 487 1174
rect 491 1170 615 1174
rect 619 1170 663 1174
rect 667 1170 759 1174
rect 763 1170 823 1174
rect 827 1170 911 1174
rect 915 1170 975 1174
rect 979 1170 1063 1174
rect 1067 1170 1119 1174
rect 1123 1170 1231 1174
rect 1235 1170 1255 1174
rect 1259 1170 1391 1174
rect 1395 1170 1399 1174
rect 1403 1170 1535 1174
rect 1539 1170 1575 1174
rect 1579 1170 1735 1174
rect 1739 1170 1823 1174
rect 1827 1170 1847 1174
rect 103 1169 1847 1170
rect 1853 1174 1863 1175
rect 1867 1174 1895 1178
rect 1899 1174 1911 1178
rect 1915 1174 1999 1178
rect 2003 1174 2063 1178
rect 2067 1174 2103 1178
rect 2107 1174 2223 1178
rect 2227 1174 2255 1178
rect 2259 1174 2359 1178
rect 2363 1174 2439 1178
rect 2443 1174 2495 1178
rect 2499 1174 2615 1178
rect 2619 1174 2639 1178
rect 2643 1174 2783 1178
rect 2787 1174 2791 1178
rect 2795 1174 2927 1178
rect 2931 1174 2967 1178
rect 2971 1174 3071 1178
rect 3075 1174 3143 1178
rect 3147 1174 3215 1178
rect 3219 1174 3327 1178
rect 3331 1174 3359 1178
rect 3363 1174 3487 1178
rect 3491 1174 3575 1178
rect 3579 1174 3618 1178
rect 1853 1173 3618 1174
rect 1853 1169 1854 1173
rect 84 1097 85 1103
rect 91 1102 1835 1103
rect 91 1098 111 1102
rect 115 1098 159 1102
rect 163 1098 215 1102
rect 219 1098 311 1102
rect 315 1098 327 1102
rect 331 1098 439 1102
rect 443 1098 463 1102
rect 467 1098 559 1102
rect 563 1098 607 1102
rect 611 1098 679 1102
rect 683 1098 751 1102
rect 755 1098 807 1102
rect 811 1098 903 1102
rect 907 1098 943 1102
rect 947 1098 1055 1102
rect 1059 1098 1087 1102
rect 1091 1098 1223 1102
rect 1227 1098 1247 1102
rect 1251 1098 1391 1102
rect 1395 1098 1407 1102
rect 1411 1098 1567 1102
rect 1571 1098 1575 1102
rect 1579 1098 1727 1102
rect 1731 1098 1823 1102
rect 1827 1098 1835 1102
rect 91 1097 1835 1098
rect 1841 1099 1842 1103
rect 1841 1098 3606 1099
rect 1841 1097 1863 1098
rect 1834 1094 1863 1097
rect 1867 1094 1887 1098
rect 1891 1094 1935 1098
rect 1939 1094 2055 1098
rect 2059 1094 2095 1098
rect 2099 1094 2247 1098
rect 2251 1094 2407 1098
rect 2411 1094 2431 1098
rect 2435 1094 2567 1098
rect 2571 1094 2607 1098
rect 2611 1094 2735 1098
rect 2739 1094 2783 1098
rect 2787 1094 2911 1098
rect 2915 1094 2959 1098
rect 2963 1094 3095 1098
rect 3099 1094 3135 1098
rect 3139 1094 3287 1098
rect 3291 1094 3319 1098
rect 3323 1094 3479 1098
rect 3483 1094 3575 1098
rect 3579 1094 3606 1098
rect 1834 1093 3606 1094
rect 96 1021 97 1027
rect 103 1026 1847 1027
rect 103 1022 111 1026
rect 115 1022 223 1026
rect 227 1022 335 1026
rect 339 1022 343 1026
rect 347 1022 431 1026
rect 435 1022 447 1026
rect 451 1022 535 1026
rect 539 1022 567 1026
rect 571 1022 655 1026
rect 659 1022 687 1026
rect 691 1022 791 1026
rect 795 1022 815 1026
rect 819 1022 951 1026
rect 955 1022 1095 1026
rect 1099 1022 1135 1026
rect 1139 1022 1255 1026
rect 1259 1022 1327 1026
rect 1331 1022 1415 1026
rect 1419 1022 1535 1026
rect 1539 1022 1583 1026
rect 1587 1022 1735 1026
rect 1739 1022 1823 1026
rect 1827 1022 1847 1026
rect 103 1021 1847 1022
rect 1853 1026 3618 1027
rect 1853 1022 1863 1026
rect 1867 1022 1943 1026
rect 1947 1022 2071 1026
rect 2075 1022 2103 1026
rect 2107 1022 2191 1026
rect 2195 1022 2255 1026
rect 2259 1022 2311 1026
rect 2315 1022 2415 1026
rect 2419 1022 2439 1026
rect 2443 1022 2575 1026
rect 2579 1022 2719 1026
rect 2723 1022 2743 1026
rect 2747 1022 2871 1026
rect 2875 1022 2919 1026
rect 2923 1022 3031 1026
rect 3035 1022 3103 1026
rect 3107 1022 3191 1026
rect 3195 1022 3295 1026
rect 3299 1022 3351 1026
rect 3355 1022 3487 1026
rect 3491 1022 3575 1026
rect 3579 1022 3618 1026
rect 1853 1021 3618 1022
rect 84 949 85 955
rect 91 954 1835 955
rect 91 950 111 954
rect 115 950 335 954
rect 339 950 367 954
rect 371 950 423 954
rect 427 950 463 954
rect 467 950 527 954
rect 531 950 575 954
rect 579 950 647 954
rect 651 950 703 954
rect 707 950 783 954
rect 787 950 847 954
rect 851 950 943 954
rect 947 950 1007 954
rect 1011 950 1127 954
rect 1131 950 1175 954
rect 1179 950 1319 954
rect 1323 950 1351 954
rect 1355 950 1527 954
rect 1531 950 1711 954
rect 1715 950 1727 954
rect 1731 950 1823 954
rect 1827 950 1835 954
rect 91 949 1835 950
rect 1841 954 3606 955
rect 1841 950 1863 954
rect 1867 950 1887 954
rect 1891 950 1935 954
rect 1939 950 2047 954
rect 2051 950 2063 954
rect 2067 950 2183 954
rect 2187 950 2199 954
rect 2203 950 2303 954
rect 2307 950 2351 954
rect 2355 950 2431 954
rect 2435 950 2495 954
rect 2499 950 2567 954
rect 2571 950 2631 954
rect 2635 950 2711 954
rect 2715 950 2759 954
rect 2763 950 2863 954
rect 2867 950 2887 954
rect 2891 950 3023 954
rect 3027 950 3183 954
rect 3187 950 3343 954
rect 3347 950 3479 954
rect 3483 950 3575 954
rect 3579 950 3606 954
rect 1841 949 3606 950
rect 1846 886 3618 887
rect 1846 883 1863 886
rect 96 877 97 883
rect 103 882 1847 883
rect 103 878 111 882
rect 115 878 343 882
rect 347 878 375 882
rect 379 878 431 882
rect 435 878 471 882
rect 475 878 535 882
rect 539 878 583 882
rect 587 878 647 882
rect 651 878 711 882
rect 715 878 783 882
rect 787 878 855 882
rect 859 878 927 882
rect 931 878 1015 882
rect 1019 878 1087 882
rect 1091 878 1183 882
rect 1187 878 1263 882
rect 1267 878 1359 882
rect 1363 878 1447 882
rect 1451 878 1535 882
rect 1539 878 1631 882
rect 1635 878 1719 882
rect 1723 878 1823 882
rect 1827 878 1847 882
rect 103 877 1847 878
rect 1853 882 1863 883
rect 1867 882 1895 886
rect 1899 882 2015 886
rect 2019 882 2055 886
rect 2059 882 2167 886
rect 2171 882 2207 886
rect 2211 882 2319 886
rect 2323 882 2359 886
rect 2363 882 2487 886
rect 2491 882 2503 886
rect 2507 882 2639 886
rect 2643 882 2663 886
rect 2667 882 2767 886
rect 2771 882 2847 886
rect 2851 882 2895 886
rect 2899 882 3031 886
rect 3035 882 3039 886
rect 3043 882 3239 886
rect 3243 882 3439 886
rect 3443 882 3575 886
rect 3579 882 3618 886
rect 1853 881 3618 882
rect 1853 877 1854 881
rect 1834 818 3606 819
rect 1834 815 1863 818
rect 84 809 85 815
rect 91 814 1835 815
rect 91 810 111 814
rect 115 810 287 814
rect 291 810 335 814
rect 339 810 407 814
rect 411 810 423 814
rect 427 810 527 814
rect 531 810 535 814
rect 539 810 639 814
rect 643 810 679 814
rect 683 810 775 814
rect 779 810 823 814
rect 827 810 919 814
rect 923 810 975 814
rect 979 810 1079 814
rect 1083 810 1127 814
rect 1131 810 1255 814
rect 1259 810 1279 814
rect 1283 810 1439 814
rect 1443 810 1599 814
rect 1603 810 1623 814
rect 1627 810 1823 814
rect 1827 810 1835 814
rect 91 809 1835 810
rect 1841 814 1863 815
rect 1867 814 1887 818
rect 1891 814 1991 818
rect 1995 814 2007 818
rect 2011 814 2135 818
rect 2139 814 2159 818
rect 2163 814 2287 818
rect 2291 814 2311 818
rect 2315 814 2455 818
rect 2459 814 2479 818
rect 2483 814 2623 818
rect 2627 814 2655 818
rect 2659 814 2799 818
rect 2803 814 2839 818
rect 2843 814 2967 818
rect 2971 814 3031 818
rect 3035 814 3143 818
rect 3147 814 3231 818
rect 3235 814 3319 818
rect 3323 814 3431 818
rect 3435 814 3479 818
rect 3483 814 3575 818
rect 3579 814 3606 818
rect 1841 813 3606 814
rect 1841 809 1842 813
rect 1846 746 3618 747
rect 1846 743 1863 746
rect 96 737 97 743
rect 103 742 1847 743
rect 103 738 111 742
rect 115 738 215 742
rect 219 738 295 742
rect 299 738 359 742
rect 363 738 415 742
rect 419 738 503 742
rect 507 738 543 742
rect 547 738 647 742
rect 651 738 687 742
rect 691 738 791 742
rect 795 738 831 742
rect 835 738 935 742
rect 939 738 983 742
rect 987 738 1087 742
rect 1091 738 1135 742
rect 1139 738 1247 742
rect 1251 738 1287 742
rect 1291 738 1415 742
rect 1419 738 1447 742
rect 1451 738 1583 742
rect 1587 738 1607 742
rect 1611 738 1735 742
rect 1739 738 1823 742
rect 1827 738 1847 742
rect 103 737 1847 738
rect 1853 742 1863 743
rect 1867 742 1895 746
rect 1899 742 1999 746
rect 2003 742 2063 746
rect 2067 742 2143 746
rect 2147 742 2255 746
rect 2259 742 2295 746
rect 2299 742 2447 746
rect 2451 742 2463 746
rect 2467 742 2631 746
rect 2635 742 2639 746
rect 2643 742 2807 746
rect 2811 742 2823 746
rect 2827 742 2975 746
rect 2979 742 2999 746
rect 3003 742 3151 746
rect 3155 742 3167 746
rect 3171 742 3327 746
rect 3331 742 3335 746
rect 3339 742 3487 746
rect 3491 742 3575 746
rect 3579 742 3618 746
rect 1853 741 3618 742
rect 1853 737 1854 741
rect 84 669 85 675
rect 91 674 1835 675
rect 91 670 111 674
rect 115 670 135 674
rect 139 670 207 674
rect 211 670 295 674
rect 299 670 351 674
rect 355 670 463 674
rect 467 670 495 674
rect 499 670 623 674
rect 627 670 639 674
rect 643 670 775 674
rect 779 670 783 674
rect 787 670 927 674
rect 931 670 1071 674
rect 1075 670 1079 674
rect 1083 670 1207 674
rect 1211 670 1239 674
rect 1243 670 1343 674
rect 1347 670 1407 674
rect 1411 670 1479 674
rect 1483 670 1575 674
rect 1579 670 1615 674
rect 1619 670 1727 674
rect 1731 670 1823 674
rect 1827 670 1835 674
rect 91 669 1835 670
rect 1841 674 3606 675
rect 1841 670 1863 674
rect 1867 670 1887 674
rect 1891 670 2055 674
rect 2059 670 2215 674
rect 2219 670 2247 674
rect 2251 670 2359 674
rect 2363 670 2439 674
rect 2443 670 2511 674
rect 2515 670 2631 674
rect 2635 670 2671 674
rect 2675 670 2815 674
rect 2819 670 2831 674
rect 2835 670 2991 674
rect 2995 670 3159 674
rect 3163 670 3327 674
rect 3331 670 3479 674
rect 3483 670 3575 674
rect 3579 670 3606 674
rect 1841 669 3606 670
rect 96 597 97 603
rect 103 602 1847 603
rect 103 598 111 602
rect 115 598 143 602
rect 147 598 303 602
rect 307 598 471 602
rect 475 598 487 602
rect 491 598 631 602
rect 635 598 671 602
rect 675 598 783 602
rect 787 598 847 602
rect 851 598 935 602
rect 939 598 1023 602
rect 1027 598 1079 602
rect 1083 598 1199 602
rect 1203 598 1215 602
rect 1219 598 1351 602
rect 1355 598 1375 602
rect 1379 598 1487 602
rect 1491 598 1559 602
rect 1563 598 1623 602
rect 1627 598 1735 602
rect 1739 598 1823 602
rect 1827 598 1847 602
rect 103 597 1847 598
rect 1853 602 3618 603
rect 1853 598 1863 602
rect 1867 598 2199 602
rect 2203 598 2223 602
rect 2227 598 2287 602
rect 2291 598 2367 602
rect 2371 598 2375 602
rect 2379 598 2463 602
rect 2467 598 2519 602
rect 2523 598 2567 602
rect 2571 598 2679 602
rect 2683 598 2815 602
rect 2819 598 2839 602
rect 2843 598 2975 602
rect 2979 598 2999 602
rect 3003 598 3143 602
rect 3147 598 3167 602
rect 3171 598 3327 602
rect 3331 598 3335 602
rect 3339 598 3487 602
rect 3491 598 3575 602
rect 3579 598 3618 602
rect 1853 597 3618 598
rect 84 525 85 531
rect 91 530 1835 531
rect 91 526 111 530
rect 115 526 135 530
rect 139 526 295 530
rect 299 526 303 530
rect 307 526 479 530
rect 483 526 495 530
rect 499 526 663 530
rect 667 526 679 530
rect 683 526 839 530
rect 843 526 863 530
rect 867 526 1015 530
rect 1019 526 1031 530
rect 1035 526 1191 530
rect 1195 526 1351 530
rect 1355 526 1367 530
rect 1371 526 1503 530
rect 1507 526 1551 530
rect 1555 526 1663 530
rect 1667 526 1727 530
rect 1731 526 1823 530
rect 1827 526 1835 530
rect 91 525 1835 526
rect 1841 530 3606 531
rect 1841 526 1863 530
rect 1867 526 2191 530
rect 2195 526 2279 530
rect 2283 526 2303 530
rect 2307 526 2367 530
rect 2371 526 2399 530
rect 2403 526 2455 530
rect 2459 526 2503 530
rect 2507 526 2559 530
rect 2563 526 2607 530
rect 2611 526 2671 530
rect 2675 526 2719 530
rect 2723 526 2807 530
rect 2811 526 2839 530
rect 2843 526 2967 530
rect 2971 526 3095 530
rect 3099 526 3135 530
rect 3139 526 3223 530
rect 3227 526 3319 530
rect 3323 526 3351 530
rect 3355 526 3479 530
rect 3483 526 3575 530
rect 3579 526 3606 530
rect 1841 525 3606 526
rect 1846 462 3618 463
rect 1846 459 1863 462
rect 96 453 97 459
rect 103 458 1847 459
rect 103 454 111 458
rect 115 454 143 458
rect 147 454 303 458
rect 307 454 311 458
rect 315 454 495 458
rect 499 454 503 458
rect 507 454 687 458
rect 691 454 871 458
rect 875 454 879 458
rect 883 454 1039 458
rect 1043 454 1055 458
rect 1059 454 1199 458
rect 1203 454 1223 458
rect 1227 454 1359 458
rect 1363 454 1391 458
rect 1395 454 1511 458
rect 1515 454 1559 458
rect 1563 454 1671 458
rect 1675 454 1727 458
rect 1731 454 1823 458
rect 1827 454 1847 458
rect 103 453 1847 454
rect 1853 458 1863 459
rect 1867 458 2239 462
rect 2243 458 2311 462
rect 2315 458 2327 462
rect 2331 458 2407 462
rect 2411 458 2431 462
rect 2435 458 2511 462
rect 2515 458 2559 462
rect 2563 458 2615 462
rect 2619 458 2695 462
rect 2699 458 2727 462
rect 2731 458 2847 462
rect 2851 458 2975 462
rect 2979 458 2999 462
rect 3003 458 3103 462
rect 3107 458 3159 462
rect 3163 458 3231 462
rect 3235 458 3327 462
rect 3331 458 3359 462
rect 3363 458 3487 462
rect 3491 458 3575 462
rect 3579 458 3618 462
rect 1853 457 3618 458
rect 1853 453 1854 457
rect 1834 394 3606 395
rect 1834 391 1863 394
rect 84 385 85 391
rect 91 390 1835 391
rect 91 386 111 390
rect 115 386 135 390
rect 139 386 263 390
rect 267 386 295 390
rect 299 386 423 390
rect 427 386 487 390
rect 491 386 591 390
rect 595 386 679 390
rect 683 386 767 390
rect 771 386 871 390
rect 875 386 935 390
rect 939 386 1047 390
rect 1051 386 1103 390
rect 1107 386 1215 390
rect 1219 386 1263 390
rect 1267 386 1383 390
rect 1387 386 1423 390
rect 1427 386 1551 390
rect 1555 386 1583 390
rect 1587 386 1719 390
rect 1723 386 1727 390
rect 1731 386 1823 390
rect 1827 386 1835 390
rect 91 385 1835 386
rect 1841 390 1863 391
rect 1867 390 2183 394
rect 2187 390 2231 394
rect 2235 390 2287 394
rect 2291 390 2319 394
rect 2323 390 2399 394
rect 2403 390 2423 394
rect 2427 390 2527 394
rect 2531 390 2551 394
rect 2555 390 2671 394
rect 2675 390 2687 394
rect 2691 390 2815 394
rect 2819 390 2839 394
rect 2843 390 2967 394
rect 2971 390 2991 394
rect 2995 390 3127 394
rect 3131 390 3151 394
rect 3155 390 3295 394
rect 3299 390 3319 394
rect 3323 390 3463 394
rect 3467 390 3479 394
rect 3483 390 3575 394
rect 3579 390 3606 394
rect 1841 389 3606 390
rect 1841 385 1842 389
rect 96 317 97 323
rect 103 322 1847 323
rect 103 318 111 322
rect 115 318 143 322
rect 147 318 215 322
rect 219 318 271 322
rect 275 318 351 322
rect 355 318 431 322
rect 435 318 495 322
rect 499 318 599 322
rect 603 318 639 322
rect 643 318 775 322
rect 779 318 791 322
rect 795 318 935 322
rect 939 318 943 322
rect 947 318 1079 322
rect 1083 318 1111 322
rect 1115 318 1223 322
rect 1227 318 1271 322
rect 1275 318 1359 322
rect 1363 318 1431 322
rect 1435 318 1487 322
rect 1491 318 1591 322
rect 1595 318 1623 322
rect 1627 318 1735 322
rect 1739 318 1823 322
rect 1827 318 1847 322
rect 103 317 1847 318
rect 1853 319 1854 323
rect 1853 318 3618 319
rect 1853 317 1863 318
rect 1846 314 1863 317
rect 1867 314 1895 318
rect 1899 314 2087 318
rect 2091 314 2191 318
rect 2195 314 2295 318
rect 2299 314 2303 318
rect 2307 314 2407 318
rect 2411 314 2511 318
rect 2515 314 2535 318
rect 2539 314 2679 318
rect 2683 314 2711 318
rect 2715 314 2823 318
rect 2827 314 2903 318
rect 2907 314 2975 318
rect 2979 314 3095 318
rect 3099 314 3135 318
rect 3139 314 3295 318
rect 3299 314 3303 318
rect 3307 314 3471 318
rect 3475 314 3487 318
rect 3491 314 3575 318
rect 3579 314 3618 318
rect 1846 313 3618 314
rect 1834 250 3606 251
rect 1834 247 1863 250
rect 84 241 85 247
rect 91 246 1835 247
rect 91 242 111 246
rect 115 242 207 246
rect 211 242 231 246
rect 235 242 343 246
rect 347 242 359 246
rect 363 242 487 246
rect 491 242 623 246
rect 627 242 631 246
rect 635 242 759 246
rect 763 242 783 246
rect 787 242 895 246
rect 899 242 927 246
rect 931 242 1031 246
rect 1035 242 1071 246
rect 1075 242 1159 246
rect 1163 242 1215 246
rect 1219 242 1295 246
rect 1299 242 1351 246
rect 1355 242 1431 246
rect 1435 242 1479 246
rect 1483 242 1615 246
rect 1619 242 1727 246
rect 1731 242 1823 246
rect 1827 242 1835 246
rect 91 241 1835 242
rect 1841 246 1863 247
rect 1867 246 1887 250
rect 1891 246 1999 250
rect 2003 246 2079 250
rect 2083 246 2143 250
rect 2147 246 2295 250
rect 2299 246 2455 250
rect 2459 246 2503 250
rect 2507 246 2615 250
rect 2619 246 2703 250
rect 2707 246 2783 250
rect 2787 246 2895 250
rect 2899 246 2951 250
rect 2955 246 3087 250
rect 3091 246 3127 250
rect 3131 246 3287 250
rect 3291 246 3311 250
rect 3315 246 3479 250
rect 3483 246 3575 250
rect 3579 246 3606 250
rect 1841 245 3606 246
rect 1841 241 1842 245
rect 96 149 97 155
rect 103 154 1847 155
rect 103 150 111 154
rect 115 150 175 154
rect 179 150 239 154
rect 243 150 263 154
rect 267 150 351 154
rect 355 150 367 154
rect 371 150 439 154
rect 443 150 495 154
rect 499 150 527 154
rect 531 150 615 154
rect 619 150 631 154
rect 635 150 703 154
rect 707 150 767 154
rect 771 150 791 154
rect 795 150 879 154
rect 883 150 903 154
rect 907 150 967 154
rect 971 150 1039 154
rect 1043 150 1055 154
rect 1059 150 1143 154
rect 1147 150 1167 154
rect 1171 150 1231 154
rect 1235 150 1303 154
rect 1307 150 1319 154
rect 1323 150 1407 154
rect 1411 150 1439 154
rect 1443 150 1503 154
rect 1507 150 1823 154
rect 1827 150 1847 154
rect 103 149 1847 150
rect 1853 154 3618 155
rect 1853 150 1863 154
rect 1867 150 1895 154
rect 1899 150 1983 154
rect 1987 150 2007 154
rect 2011 150 2071 154
rect 2075 150 2151 154
rect 2155 150 2159 154
rect 2163 150 2247 154
rect 2251 150 2303 154
rect 2307 150 2335 154
rect 2339 150 2439 154
rect 2443 150 2463 154
rect 2467 150 2543 154
rect 2547 150 2623 154
rect 2627 150 2647 154
rect 2651 150 2743 154
rect 2747 150 2791 154
rect 2795 150 2839 154
rect 2843 150 2935 154
rect 2939 150 2959 154
rect 2963 150 3031 154
rect 3035 150 3127 154
rect 3131 150 3135 154
rect 3139 150 3223 154
rect 3227 150 3311 154
rect 3315 150 3319 154
rect 3323 150 3399 154
rect 3403 150 3487 154
rect 3491 150 3575 154
rect 3579 150 3618 154
rect 1853 149 3618 150
rect 84 81 85 87
rect 91 86 1835 87
rect 91 82 111 86
rect 115 82 167 86
rect 171 82 255 86
rect 259 82 343 86
rect 347 82 431 86
rect 435 82 519 86
rect 523 82 607 86
rect 611 82 695 86
rect 699 82 783 86
rect 787 82 871 86
rect 875 82 959 86
rect 963 82 1047 86
rect 1051 82 1135 86
rect 1139 82 1223 86
rect 1227 82 1311 86
rect 1315 82 1399 86
rect 1403 82 1495 86
rect 1499 82 1823 86
rect 1827 82 1835 86
rect 91 81 1835 82
rect 1841 86 3606 87
rect 1841 82 1863 86
rect 1867 82 1887 86
rect 1891 82 1975 86
rect 1979 82 2063 86
rect 2067 82 2151 86
rect 2155 82 2239 86
rect 2243 82 2327 86
rect 2331 82 2431 86
rect 2435 82 2535 86
rect 2539 82 2639 86
rect 2643 82 2735 86
rect 2739 82 2831 86
rect 2835 82 2927 86
rect 2931 82 3023 86
rect 3027 82 3119 86
rect 3123 82 3215 86
rect 3219 82 3303 86
rect 3307 82 3391 86
rect 3395 82 3479 86
rect 3483 82 3575 86
rect 3579 82 3606 86
rect 1841 81 3606 82
<< m5c >>
rect 97 3645 103 3651
rect 1847 3645 1853 3651
rect 1835 3581 1841 3587
rect 3599 3581 3605 3587
rect 85 3569 91 3575
rect 1835 3569 1841 3575
rect 97 3501 103 3507
rect 1847 3501 1853 3507
rect 85 3433 91 3439
rect 1835 3433 1841 3439
rect 97 3357 103 3363
rect 1847 3357 1853 3363
rect 85 3285 91 3291
rect 1835 3285 1841 3291
rect 97 3213 103 3219
rect 1847 3213 1853 3219
rect 85 3141 91 3147
rect 1835 3141 1841 3147
rect 97 3065 103 3071
rect 1847 3065 1853 3071
rect 85 2989 91 2995
rect 1835 2989 1841 2995
rect 97 2921 103 2927
rect 1847 2921 1853 2927
rect 1847 2909 1853 2915
rect 3611 2909 3617 2915
rect 85 2849 91 2855
rect 1835 2849 1841 2855
rect 1835 2837 1841 2843
rect 3599 2837 3605 2843
rect 97 2781 103 2787
rect 1847 2781 1853 2787
rect 1847 2757 1853 2763
rect 3611 2757 3617 2763
rect 85 2705 91 2711
rect 1835 2705 1841 2711
rect 1835 2689 1841 2695
rect 3599 2689 3605 2695
rect 97 2621 103 2627
rect 1847 2621 1853 2627
rect 85 2553 91 2559
rect 1835 2553 1841 2559
rect 97 2481 103 2487
rect 1847 2481 1853 2487
rect 85 2405 91 2411
rect 1835 2405 1841 2411
rect 97 2333 103 2339
rect 1847 2333 1853 2339
rect 85 2265 91 2271
rect 1835 2265 1841 2271
rect 97 2193 103 2199
rect 1847 2193 1853 2199
rect 85 2117 91 2123
rect 1835 2117 1841 2123
rect 1847 2049 1853 2055
rect 3611 2049 3617 2055
rect 97 2037 103 2043
rect 1847 2037 1853 2043
rect 85 1969 91 1975
rect 1835 1969 1841 1975
rect 1847 1905 1853 1911
rect 3611 1905 3617 1911
rect 97 1893 103 1899
rect 1847 1893 1853 1899
rect 1835 1833 1841 1839
rect 3599 1833 3605 1839
rect 85 1825 91 1831
rect 1835 1825 1841 1831
rect 1847 1761 1853 1767
rect 3611 1761 3617 1767
rect 97 1753 103 1759
rect 1847 1753 1853 1759
rect 1835 1689 1841 1695
rect 3599 1689 3605 1695
rect 85 1681 91 1687
rect 1835 1681 1841 1687
rect 1847 1613 1853 1619
rect 3611 1613 3617 1619
rect 97 1605 103 1611
rect 1847 1605 1853 1611
rect 85 1533 91 1539
rect 1835 1533 1841 1539
rect 97 1457 103 1463
rect 1847 1457 1853 1463
rect 85 1389 91 1395
rect 1835 1389 1841 1395
rect 97 1313 103 1319
rect 1847 1313 1853 1319
rect 85 1241 91 1247
rect 1835 1241 1841 1247
rect 97 1169 103 1175
rect 1847 1169 1853 1175
rect 85 1097 91 1103
rect 1835 1097 1841 1103
rect 97 1021 103 1027
rect 1847 1021 1853 1027
rect 85 949 91 955
rect 1835 949 1841 955
rect 97 877 103 883
rect 1847 877 1853 883
rect 85 809 91 815
rect 1835 809 1841 815
rect 97 737 103 743
rect 1847 737 1853 743
rect 85 669 91 675
rect 1835 669 1841 675
rect 97 597 103 603
rect 1847 597 1853 603
rect 85 525 91 531
rect 1835 525 1841 531
rect 97 453 103 459
rect 1847 453 1853 459
rect 85 385 91 391
rect 1835 385 1841 391
rect 97 317 103 323
rect 1847 317 1853 323
rect 85 241 91 247
rect 1835 241 1841 247
rect 97 149 103 155
rect 1847 149 1853 155
rect 85 81 91 87
rect 1835 81 1841 87
<< m5 >>
rect 84 3575 92 3672
rect 84 3569 85 3575
rect 91 3569 92 3575
rect 84 3439 92 3569
rect 84 3433 85 3439
rect 91 3433 92 3439
rect 84 3291 92 3433
rect 84 3285 85 3291
rect 91 3285 92 3291
rect 84 3147 92 3285
rect 84 3141 85 3147
rect 91 3141 92 3147
rect 84 2995 92 3141
rect 84 2989 85 2995
rect 91 2989 92 2995
rect 84 2855 92 2989
rect 84 2849 85 2855
rect 91 2849 92 2855
rect 84 2711 92 2849
rect 84 2705 85 2711
rect 91 2705 92 2711
rect 84 2559 92 2705
rect 84 2553 85 2559
rect 91 2553 92 2559
rect 84 2411 92 2553
rect 84 2405 85 2411
rect 91 2405 92 2411
rect 84 2271 92 2405
rect 84 2265 85 2271
rect 91 2265 92 2271
rect 84 2123 92 2265
rect 84 2117 85 2123
rect 91 2117 92 2123
rect 84 1975 92 2117
rect 84 1969 85 1975
rect 91 1969 92 1975
rect 84 1831 92 1969
rect 84 1825 85 1831
rect 91 1825 92 1831
rect 84 1687 92 1825
rect 84 1681 85 1687
rect 91 1681 92 1687
rect 84 1539 92 1681
rect 84 1533 85 1539
rect 91 1533 92 1539
rect 84 1395 92 1533
rect 84 1389 85 1395
rect 91 1389 92 1395
rect 84 1247 92 1389
rect 84 1241 85 1247
rect 91 1241 92 1247
rect 84 1103 92 1241
rect 84 1097 85 1103
rect 91 1097 92 1103
rect 84 955 92 1097
rect 84 949 85 955
rect 91 949 92 955
rect 84 815 92 949
rect 84 809 85 815
rect 91 809 92 815
rect 84 675 92 809
rect 84 669 85 675
rect 91 669 92 675
rect 84 531 92 669
rect 84 525 85 531
rect 91 525 92 531
rect 84 391 92 525
rect 84 385 85 391
rect 91 385 92 391
rect 84 247 92 385
rect 84 241 85 247
rect 91 241 92 247
rect 84 87 92 241
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 3651 104 3672
rect 96 3645 97 3651
rect 103 3645 104 3651
rect 96 3507 104 3645
rect 96 3501 97 3507
rect 103 3501 104 3507
rect 96 3363 104 3501
rect 96 3357 97 3363
rect 103 3357 104 3363
rect 96 3219 104 3357
rect 96 3213 97 3219
rect 103 3213 104 3219
rect 96 3071 104 3213
rect 96 3065 97 3071
rect 103 3065 104 3071
rect 96 2927 104 3065
rect 96 2921 97 2927
rect 103 2921 104 2927
rect 96 2787 104 2921
rect 96 2781 97 2787
rect 103 2781 104 2787
rect 96 2627 104 2781
rect 96 2621 97 2627
rect 103 2621 104 2627
rect 96 2487 104 2621
rect 96 2481 97 2487
rect 103 2481 104 2487
rect 96 2339 104 2481
rect 96 2333 97 2339
rect 103 2333 104 2339
rect 96 2199 104 2333
rect 96 2193 97 2199
rect 103 2193 104 2199
rect 96 2043 104 2193
rect 96 2037 97 2043
rect 103 2037 104 2043
rect 96 1899 104 2037
rect 96 1893 97 1899
rect 103 1893 104 1899
rect 96 1759 104 1893
rect 96 1753 97 1759
rect 103 1753 104 1759
rect 96 1611 104 1753
rect 96 1605 97 1611
rect 103 1605 104 1611
rect 96 1463 104 1605
rect 96 1457 97 1463
rect 103 1457 104 1463
rect 96 1319 104 1457
rect 96 1313 97 1319
rect 103 1313 104 1319
rect 96 1175 104 1313
rect 96 1169 97 1175
rect 103 1169 104 1175
rect 96 1027 104 1169
rect 96 1021 97 1027
rect 103 1021 104 1027
rect 96 883 104 1021
rect 96 877 97 883
rect 103 877 104 883
rect 96 743 104 877
rect 96 737 97 743
rect 103 737 104 743
rect 96 603 104 737
rect 96 597 97 603
rect 103 597 104 603
rect 96 459 104 597
rect 96 453 97 459
rect 103 453 104 459
rect 96 323 104 453
rect 96 317 97 323
rect 103 317 104 323
rect 96 155 104 317
rect 96 149 97 155
rect 103 149 104 155
rect 96 72 104 149
rect 1834 3587 1842 3672
rect 1834 3581 1835 3587
rect 1841 3581 1842 3587
rect 1834 3575 1842 3581
rect 1834 3569 1835 3575
rect 1841 3569 1842 3575
rect 1834 3439 1842 3569
rect 1834 3433 1835 3439
rect 1841 3433 1842 3439
rect 1834 3291 1842 3433
rect 1834 3285 1835 3291
rect 1841 3285 1842 3291
rect 1834 3147 1842 3285
rect 1834 3141 1835 3147
rect 1841 3141 1842 3147
rect 1834 2995 1842 3141
rect 1834 2989 1835 2995
rect 1841 2989 1842 2995
rect 1834 2855 1842 2989
rect 1834 2849 1835 2855
rect 1841 2849 1842 2855
rect 1834 2843 1842 2849
rect 1834 2837 1835 2843
rect 1841 2837 1842 2843
rect 1834 2711 1842 2837
rect 1834 2705 1835 2711
rect 1841 2705 1842 2711
rect 1834 2695 1842 2705
rect 1834 2689 1835 2695
rect 1841 2689 1842 2695
rect 1834 2559 1842 2689
rect 1834 2553 1835 2559
rect 1841 2553 1842 2559
rect 1834 2411 1842 2553
rect 1834 2405 1835 2411
rect 1841 2405 1842 2411
rect 1834 2271 1842 2405
rect 1834 2265 1835 2271
rect 1841 2265 1842 2271
rect 1834 2123 1842 2265
rect 1834 2117 1835 2123
rect 1841 2117 1842 2123
rect 1834 1975 1842 2117
rect 1834 1969 1835 1975
rect 1841 1969 1842 1975
rect 1834 1839 1842 1969
rect 1834 1833 1835 1839
rect 1841 1833 1842 1839
rect 1834 1831 1842 1833
rect 1834 1825 1835 1831
rect 1841 1825 1842 1831
rect 1834 1695 1842 1825
rect 1834 1689 1835 1695
rect 1841 1689 1842 1695
rect 1834 1687 1842 1689
rect 1834 1681 1835 1687
rect 1841 1681 1842 1687
rect 1834 1539 1842 1681
rect 1834 1533 1835 1539
rect 1841 1533 1842 1539
rect 1834 1395 1842 1533
rect 1834 1389 1835 1395
rect 1841 1389 1842 1395
rect 1834 1247 1842 1389
rect 1834 1241 1835 1247
rect 1841 1241 1842 1247
rect 1834 1103 1842 1241
rect 1834 1097 1835 1103
rect 1841 1097 1842 1103
rect 1834 955 1842 1097
rect 1834 949 1835 955
rect 1841 949 1842 955
rect 1834 815 1842 949
rect 1834 809 1835 815
rect 1841 809 1842 815
rect 1834 675 1842 809
rect 1834 669 1835 675
rect 1841 669 1842 675
rect 1834 531 1842 669
rect 1834 525 1835 531
rect 1841 525 1842 531
rect 1834 391 1842 525
rect 1834 385 1835 391
rect 1841 385 1842 391
rect 1834 247 1842 385
rect 1834 241 1835 247
rect 1841 241 1842 247
rect 1834 87 1842 241
rect 1834 81 1835 87
rect 1841 81 1842 87
rect 1834 72 1842 81
rect 1846 3651 1854 3672
rect 1846 3645 1847 3651
rect 1853 3645 1854 3651
rect 1846 3507 1854 3645
rect 1846 3501 1847 3507
rect 1853 3501 1854 3507
rect 1846 3363 1854 3501
rect 1846 3357 1847 3363
rect 1853 3357 1854 3363
rect 1846 3219 1854 3357
rect 1846 3213 1847 3219
rect 1853 3213 1854 3219
rect 1846 3071 1854 3213
rect 1846 3065 1847 3071
rect 1853 3065 1854 3071
rect 1846 2927 1854 3065
rect 1846 2921 1847 2927
rect 1853 2921 1854 2927
rect 1846 2915 1854 2921
rect 1846 2909 1847 2915
rect 1853 2909 1854 2915
rect 1846 2787 1854 2909
rect 1846 2781 1847 2787
rect 1853 2781 1854 2787
rect 1846 2763 1854 2781
rect 1846 2757 1847 2763
rect 1853 2757 1854 2763
rect 1846 2627 1854 2757
rect 1846 2621 1847 2627
rect 1853 2621 1854 2627
rect 1846 2487 1854 2621
rect 1846 2481 1847 2487
rect 1853 2481 1854 2487
rect 1846 2339 1854 2481
rect 1846 2333 1847 2339
rect 1853 2333 1854 2339
rect 1846 2199 1854 2333
rect 1846 2193 1847 2199
rect 1853 2193 1854 2199
rect 1846 2055 1854 2193
rect 1846 2049 1847 2055
rect 1853 2049 1854 2055
rect 1846 2043 1854 2049
rect 1846 2037 1847 2043
rect 1853 2037 1854 2043
rect 1846 1911 1854 2037
rect 1846 1905 1847 1911
rect 1853 1905 1854 1911
rect 1846 1899 1854 1905
rect 1846 1893 1847 1899
rect 1853 1893 1854 1899
rect 1846 1767 1854 1893
rect 1846 1761 1847 1767
rect 1853 1761 1854 1767
rect 1846 1759 1854 1761
rect 1846 1753 1847 1759
rect 1853 1753 1854 1759
rect 1846 1619 1854 1753
rect 1846 1613 1847 1619
rect 1853 1613 1854 1619
rect 1846 1611 1854 1613
rect 1846 1605 1847 1611
rect 1853 1605 1854 1611
rect 1846 1463 1854 1605
rect 1846 1457 1847 1463
rect 1853 1457 1854 1463
rect 1846 1319 1854 1457
rect 1846 1313 1847 1319
rect 1853 1313 1854 1319
rect 1846 1175 1854 1313
rect 1846 1169 1847 1175
rect 1853 1169 1854 1175
rect 1846 1027 1854 1169
rect 1846 1021 1847 1027
rect 1853 1021 1854 1027
rect 1846 883 1854 1021
rect 1846 877 1847 883
rect 1853 877 1854 883
rect 1846 743 1854 877
rect 1846 737 1847 743
rect 1853 737 1854 743
rect 1846 603 1854 737
rect 1846 597 1847 603
rect 1853 597 1854 603
rect 1846 459 1854 597
rect 1846 453 1847 459
rect 1853 453 1854 459
rect 1846 323 1854 453
rect 1846 317 1847 323
rect 1853 317 1854 323
rect 1846 155 1854 317
rect 1846 149 1847 155
rect 1853 149 1854 155
rect 1846 72 1854 149
rect 3598 3587 3606 3672
rect 3598 3581 3599 3587
rect 3605 3581 3606 3587
rect 3598 2843 3606 3581
rect 3598 2837 3599 2843
rect 3605 2837 3606 2843
rect 3598 2695 3606 2837
rect 3598 2689 3599 2695
rect 3605 2689 3606 2695
rect 3598 1839 3606 2689
rect 3598 1833 3599 1839
rect 3605 1833 3606 1839
rect 3598 1695 3606 1833
rect 3598 1689 3599 1695
rect 3605 1689 3606 1695
rect 3598 72 3606 1689
rect 3610 2915 3618 3672
rect 3610 2909 3611 2915
rect 3617 2909 3618 2915
rect 3610 2763 3618 2909
rect 3610 2757 3611 2763
rect 3617 2757 3618 2763
rect 3610 2055 3618 2757
rect 3610 2049 3611 2055
rect 3617 2049 3618 2055
rect 3610 1911 3618 2049
rect 3610 1905 3611 1911
rect 3617 1905 3618 1911
rect 3610 1767 3618 1905
rect 3610 1761 3611 1767
rect 3617 1761 3618 1767
rect 3610 1619 3618 1761
rect 3610 1613 3611 1619
rect 3617 1613 3618 1619
rect 3610 72 3618 1613
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__193
timestamp 1731220588
transform 1 0 3568 0 -1 3568
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220588
transform 1 0 1856 0 -1 3568
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220588
transform 1 0 3568 0 1 3456
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220588
transform 1 0 1856 0 1 3456
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220588
transform 1 0 3568 0 -1 3416
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220588
transform 1 0 1856 0 -1 3416
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220588
transform 1 0 3568 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220588
transform 1 0 1856 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220588
transform 1 0 3568 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220588
transform 1 0 1856 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220588
transform 1 0 3568 0 1 3168
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220588
transform 1 0 1856 0 1 3168
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220588
transform 1 0 3568 0 -1 3132
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220588
transform 1 0 1856 0 -1 3132
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220588
transform 1 0 3568 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220588
transform 1 0 1856 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220588
transform 1 0 3568 0 -1 2980
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220588
transform 1 0 1856 0 -1 2980
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220588
transform 1 0 3568 0 1 2860
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220588
transform 1 0 1856 0 1 2860
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220588
transform 1 0 3568 0 -1 2824
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220588
transform 1 0 1856 0 -1 2824
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220588
transform 1 0 3568 0 1 2708
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220588
transform 1 0 1856 0 1 2708
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220588
transform 1 0 3568 0 -1 2676
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220588
transform 1 0 1856 0 -1 2676
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220588
transform 1 0 3568 0 1 2568
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220588
transform 1 0 1856 0 1 2568
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220588
transform 1 0 3568 0 -1 2536
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220588
transform 1 0 1856 0 -1 2536
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220588
transform 1 0 3568 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220588
transform 1 0 1856 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220588
transform 1 0 3568 0 -1 2392
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220588
transform 1 0 1856 0 -1 2392
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220588
transform 1 0 3568 0 1 2284
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220588
transform 1 0 1856 0 1 2284
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220588
transform 1 0 3568 0 -1 2252
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220588
transform 1 0 1856 0 -1 2252
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220588
transform 1 0 3568 0 1 2148
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220588
transform 1 0 1856 0 1 2148
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220588
transform 1 0 3568 0 -1 2108
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220588
transform 1 0 1856 0 -1 2108
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220588
transform 1 0 3568 0 1 2000
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220588
transform 1 0 1856 0 1 2000
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220588
transform 1 0 3568 0 -1 1960
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220588
transform 1 0 1856 0 -1 1960
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220588
transform 1 0 3568 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220588
transform 1 0 1856 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220588
transform 1 0 3568 0 -1 1820
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220588
transform 1 0 1856 0 -1 1820
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220588
transform 1 0 3568 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220588
transform 1 0 1856 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220588
transform 1 0 3568 0 -1 1676
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220588
transform 1 0 1856 0 -1 1676
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220588
transform 1 0 3568 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220588
transform 1 0 1856 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220588
transform 1 0 3568 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220588
transform 1 0 1856 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220588
transform 1 0 3568 0 1 1412
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220588
transform 1 0 1856 0 1 1412
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220588
transform 1 0 3568 0 -1 1372
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220588
transform 1 0 1856 0 -1 1372
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220588
transform 1 0 3568 0 1 1268
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220588
transform 1 0 1856 0 1 1268
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220588
transform 1 0 3568 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220588
transform 1 0 1856 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220588
transform 1 0 3568 0 1 1124
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220588
transform 1 0 1856 0 1 1124
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220588
transform 1 0 3568 0 -1 1080
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220588
transform 1 0 1856 0 -1 1080
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220588
transform 1 0 3568 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220588
transform 1 0 1856 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220588
transform 1 0 3568 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220588
transform 1 0 1856 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220588
transform 1 0 3568 0 1 832
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220588
transform 1 0 1856 0 1 832
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220588
transform 1 0 3568 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220588
transform 1 0 1856 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220588
transform 1 0 3568 0 1 692
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220588
transform 1 0 1856 0 1 692
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220588
transform 1 0 3568 0 -1 656
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220588
transform 1 0 1856 0 -1 656
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220588
transform 1 0 3568 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220588
transform 1 0 1856 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220588
transform 1 0 3568 0 -1 512
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220588
transform 1 0 1856 0 -1 512
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220588
transform 1 0 3568 0 1 408
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220588
transform 1 0 1856 0 1 408
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220588
transform 1 0 3568 0 -1 376
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220588
transform 1 0 1856 0 -1 376
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220588
transform 1 0 3568 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220588
transform 1 0 1856 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220588
transform 1 0 3568 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220588
transform 1 0 1856 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220588
transform 1 0 3568 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220588
transform 1 0 1856 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220588
transform 1 0 1816 0 1 3596
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220588
transform 1 0 104 0 1 3596
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220588
transform 1 0 1816 0 -1 3556
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220588
transform 1 0 104 0 -1 3556
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220588
transform 1 0 1816 0 1 3452
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220588
transform 1 0 104 0 1 3452
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220588
transform 1 0 1816 0 -1 3420
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220588
transform 1 0 104 0 -1 3420
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220588
transform 1 0 1816 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220588
transform 1 0 104 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220588
transform 1 0 1816 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220588
transform 1 0 104 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220588
transform 1 0 1816 0 1 3164
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220588
transform 1 0 104 0 1 3164
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220588
transform 1 0 1816 0 -1 3128
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220588
transform 1 0 104 0 -1 3128
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220588
transform 1 0 1816 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220588
transform 1 0 104 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220588
transform 1 0 1816 0 -1 2976
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220588
transform 1 0 104 0 -1 2976
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220588
transform 1 0 1816 0 1 2872
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220588
transform 1 0 104 0 1 2872
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220588
transform 1 0 1816 0 -1 2836
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220588
transform 1 0 104 0 -1 2836
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220588
transform 1 0 1816 0 1 2732
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220588
transform 1 0 104 0 1 2732
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220588
transform 1 0 1816 0 -1 2692
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220588
transform 1 0 104 0 -1 2692
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220588
transform 1 0 1816 0 1 2572
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220588
transform 1 0 104 0 1 2572
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220588
transform 1 0 1816 0 -1 2540
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220588
transform 1 0 104 0 -1 2540
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220588
transform 1 0 1816 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220588
transform 1 0 104 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220588
transform 1 0 1816 0 -1 2392
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220588
transform 1 0 104 0 -1 2392
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220588
transform 1 0 1816 0 1 2284
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220588
transform 1 0 104 0 1 2284
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220588
transform 1 0 1816 0 -1 2252
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220588
transform 1 0 104 0 -1 2252
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220588
transform 1 0 1816 0 1 2144
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220588
transform 1 0 104 0 1 2144
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220588
transform 1 0 1816 0 -1 2104
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220588
transform 1 0 104 0 -1 2104
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220588
transform 1 0 1816 0 1 1988
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220588
transform 1 0 104 0 1 1988
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220588
transform 1 0 1816 0 -1 1956
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220588
transform 1 0 104 0 -1 1956
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220588
transform 1 0 1816 0 1 1844
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220588
transform 1 0 104 0 1 1844
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220588
transform 1 0 1816 0 -1 1812
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220588
transform 1 0 104 0 -1 1812
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220588
transform 1 0 1816 0 1 1704
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220588
transform 1 0 104 0 1 1704
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220588
transform 1 0 1816 0 -1 1668
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220588
transform 1 0 104 0 -1 1668
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220588
transform 1 0 1816 0 1 1556
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220588
transform 1 0 104 0 1 1556
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220588
transform 1 0 1816 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220588
transform 1 0 104 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220588
transform 1 0 1816 0 1 1408
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220588
transform 1 0 104 0 1 1408
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220588
transform 1 0 1816 0 -1 1376
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220588
transform 1 0 104 0 -1 1376
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220588
transform 1 0 1816 0 1 1264
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220588
transform 1 0 104 0 1 1264
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220588
transform 1 0 1816 0 -1 1228
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220588
transform 1 0 104 0 -1 1228
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220588
transform 1 0 1816 0 1 1120
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220588
transform 1 0 104 0 1 1120
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220588
transform 1 0 1816 0 -1 1084
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220588
transform 1 0 104 0 -1 1084
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220588
transform 1 0 1816 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220588
transform 1 0 104 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220588
transform 1 0 1816 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220588
transform 1 0 104 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220588
transform 1 0 1816 0 1 828
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220588
transform 1 0 104 0 1 828
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220588
transform 1 0 1816 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220588
transform 1 0 104 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220588
transform 1 0 1816 0 1 688
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220588
transform 1 0 104 0 1 688
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220588
transform 1 0 1816 0 -1 656
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220588
transform 1 0 104 0 -1 656
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220588
transform 1 0 1816 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220588
transform 1 0 104 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220588
transform 1 0 1816 0 -1 512
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220588
transform 1 0 104 0 -1 512
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220588
transform 1 0 1816 0 1 404
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220588
transform 1 0 104 0 1 404
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220588
transform 1 0 1816 0 -1 372
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220588
transform 1 0 104 0 -1 372
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220588
transform 1 0 1816 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220588
transform 1 0 104 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220588
transform 1 0 1816 0 -1 228
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220588
transform 1 0 104 0 -1 228
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220588
transform 1 0 1816 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220588
transform 1 0 104 0 1 100
box 7 3 12 24
use _0_0std_0_0cells_0_0MUX2X1  tst_5999_6
timestamp 1731220588
transform 1 0 3384 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5998_6
timestamp 1731220588
transform 1 0 3472 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5997_6
timestamp 1731220588
transform 1 0 3472 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5996_6
timestamp 1731220588
transform 1 0 3472 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5995_6
timestamp 1731220588
transform 1 0 3472 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5994_6
timestamp 1731220588
transform 1 0 3472 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5993_6
timestamp 1731220588
transform 1 0 3472 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5992_6
timestamp 1731220588
transform 1 0 3472 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5991_6
timestamp 1731220588
transform 1 0 3472 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5990_6
timestamp 1731220588
transform 1 0 3472 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5989_6
timestamp 1731220588
transform 1 0 3424 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5988_6
timestamp 1731220588
transform 1 0 3312 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5987_6
timestamp 1731220588
transform 1 0 3136 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5986_6
timestamp 1731220588
transform 1 0 3320 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5985_6
timestamp 1731220588
transform 1 0 3152 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5984_6
timestamp 1731220588
transform 1 0 2984 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5983_6
timestamp 1731220588
transform 1 0 2984 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5982_6
timestamp 1731220588
transform 1 0 3152 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5981_6
timestamp 1731220588
transform 1 0 3320 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5980_6
timestamp 1731220588
transform 1 0 3312 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5979_6
timestamp 1731220588
transform 1 0 3128 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5978_6
timestamp 1731220588
transform 1 0 3088 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5977_6
timestamp 1731220588
transform 1 0 2960 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5976_6
timestamp 1731220588
transform 1 0 3344 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5975_6
timestamp 1731220588
transform 1 0 3216 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5974_6
timestamp 1731220588
transform 1 0 3144 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5973_6
timestamp 1731220588
transform 1 0 3312 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5972_6
timestamp 1731220588
transform 1 0 3456 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5971_6
timestamp 1731220588
transform 1 0 3288 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5970_6
timestamp 1731220588
transform 1 0 3120 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5969_6
timestamp 1731220588
transform 1 0 3080 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5968_6
timestamp 1731220588
transform 1 0 3280 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5967_6
timestamp 1731220588
transform 1 0 3120 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5966_6
timestamp 1731220588
transform 1 0 3304 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5965_6
timestamp 1731220588
transform 1 0 3296 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5964_6
timestamp 1731220588
transform 1 0 3208 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5963_6
timestamp 1731220588
transform 1 0 3112 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5962_6
timestamp 1731220588
transform 1 0 3016 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5961_6
timestamp 1731220588
transform 1 0 2920 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5960_6
timestamp 1731220588
transform 1 0 2824 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5959_6
timestamp 1731220588
transform 1 0 2728 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5958_6
timestamp 1731220588
transform 1 0 2632 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5957_6
timestamp 1731220588
transform 1 0 2608 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5956_6
timestamp 1731220588
transform 1 0 2776 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5955_6
timestamp 1731220588
transform 1 0 2944 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5954_6
timestamp 1731220588
transform 1 0 2888 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5953_6
timestamp 1731220588
transform 1 0 2696 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5952_6
timestamp 1731220588
transform 1 0 2496 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5951_6
timestamp 1731220588
transform 1 0 2664 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5950_6
timestamp 1731220588
transform 1 0 2808 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5949_6
timestamp 1731220588
transform 1 0 2960 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5948_6
timestamp 1731220588
transform 1 0 2984 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5947_6
timestamp 1731220588
transform 1 0 2832 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5946_6
timestamp 1731220588
transform 1 0 2832 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5945_6
timestamp 1731220588
transform 1 0 2712 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5944_6
timestamp 1731220588
transform 1 0 2664 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5943_6
timestamp 1731220588
transform 1 0 2552 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5942_6
timestamp 1731220588
transform 1 0 2800 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5941_6
timestamp 1731220588
transform 1 0 2960 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5940_6
timestamp 1731220588
transform 1 0 2824 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5939_6
timestamp 1731220588
transform 1 0 2664 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5938_6
timestamp 1731220588
transform 1 0 2624 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5937_6
timestamp 1731220588
transform 1 0 2808 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5936_6
timestamp 1731220588
transform 1 0 2960 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5935_6
timestamp 1731220588
transform 1 0 2792 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5934_6
timestamp 1731220588
transform 1 0 2616 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5933_6
timestamp 1731220588
transform 1 0 2648 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5932_6
timestamp 1731220588
transform 1 0 2832 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5931_6
timestamp 1731220588
transform 1 0 3224 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5930_6
timestamp 1731220588
transform 1 0 3024 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5929_6
timestamp 1731220588
transform 1 0 3016 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5928_6
timestamp 1731220588
transform 1 0 2880 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5927_6
timestamp 1731220588
transform 1 0 2752 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5926_6
timestamp 1731220588
transform 1 0 2624 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5925_6
timestamp 1731220588
transform 1 0 2488 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5924_6
timestamp 1731220588
transform 1 0 3016 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5923_6
timestamp 1731220588
transform 1 0 2856 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5922_6
timestamp 1731220588
transform 1 0 2704 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5921_6
timestamp 1731220588
transform 1 0 2560 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5920_6
timestamp 1731220588
transform 1 0 2560 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5919_6
timestamp 1731220588
transform 1 0 2728 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5918_6
timestamp 1731220588
transform 1 0 2904 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5917_6
timestamp 1731220588
transform 1 0 3088 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5916_6
timestamp 1731220588
transform 1 0 3128 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5915_6
timestamp 1731220588
transform 1 0 2952 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5914_6
timestamp 1731220588
transform 1 0 2776 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5913_6
timestamp 1731220588
transform 1 0 2600 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5912_6
timestamp 1731220588
transform 1 0 2768 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5911_6
timestamp 1731220588
transform 1 0 3200 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5910_6
timestamp 1731220588
transform 1 0 3056 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5909_6
timestamp 1731220588
transform 1 0 2912 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5908_6
timestamp 1731220588
transform 1 0 2872 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5907_6
timestamp 1731220588
transform 1 0 2696 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5906_6
timestamp 1731220588
transform 1 0 3032 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5905_6
timestamp 1731220588
transform 1 0 3184 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5904_6
timestamp 1731220588
transform 1 0 3336 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5903_6
timestamp 1731220588
transform 1 0 3216 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5902_6
timestamp 1731220588
transform 1 0 3072 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5901_6
timestamp 1731220588
transform 1 0 2928 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5900_6
timestamp 1731220588
transform 1 0 2776 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5899_6
timestamp 1731220588
transform 1 0 3328 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5898_6
timestamp 1731220588
transform 1 0 3160 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5897_6
timestamp 1731220588
transform 1 0 2992 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5896_6
timestamp 1731220588
transform 1 0 2832 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5895_6
timestamp 1731220588
transform 1 0 2672 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5894_6
timestamp 1731220588
transform 1 0 3144 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5893_6
timestamp 1731220588
transform 1 0 2976 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5892_6
timestamp 1731220588
transform 1 0 2816 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5891_6
timestamp 1731220588
transform 1 0 2656 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5890_6
timestamp 1731220588
transform 1 0 3080 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5889_6
timestamp 1731220588
transform 1 0 2896 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5888_6
timestamp 1731220588
transform 1 0 2728 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5887_6
timestamp 1731220588
transform 1 0 2568 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5886_6
timestamp 1731220588
transform 1 0 2536 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5885_6
timestamp 1731220588
transform 1 0 2688 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5884_6
timestamp 1731220588
transform 1 0 2856 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5883_6
timestamp 1731220588
transform 1 0 3040 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5882_6
timestamp 1731220588
transform 1 0 2976 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5881_6
timestamp 1731220588
transform 1 0 2776 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5880_6
timestamp 1731220588
transform 1 0 2632 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5879_6
timestamp 1731220588
transform 1 0 2432 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5878_6
timestamp 1731220588
transform 1 0 2824 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5877_6
timestamp 1731220588
transform 1 0 3008 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5876_6
timestamp 1731220588
transform 1 0 3192 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5875_6
timestamp 1731220588
transform 1 0 3184 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5874_6
timestamp 1731220588
transform 1 0 3232 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5873_6
timestamp 1731220588
transform 1 0 3264 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5872_6
timestamp 1731220588
transform 1 0 3312 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5871_6
timestamp 1731220588
transform 1 0 3352 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5870_6
timestamp 1731220588
transform 1 0 3344 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5869_6
timestamp 1731220588
transform 1 0 3312 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5868_6
timestamp 1731220588
transform 1 0 3280 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5867_6
timestamp 1731220588
transform 1 0 3176 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5866_6
timestamp 1731220588
transform 1 0 3336 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5865_6
timestamp 1731220588
transform 1 0 3472 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5864_6
timestamp 1731220588
transform 1 0 3472 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5863_6
timestamp 1731220588
transform 1 0 3472 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5862_6
timestamp 1731220588
transform 1 0 3472 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5861_6
timestamp 1731220588
transform 1 0 3472 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5860_6
timestamp 1731220588
transform 1 0 3472 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5859_6
timestamp 1731220588
transform 1 0 3472 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5858_6
timestamp 1731220588
transform 1 0 3472 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5857_6
timestamp 1731220588
transform 1 0 3456 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5856_6
timestamp 1731220588
transform 1 0 3424 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5855_6
timestamp 1731220588
transform 1 0 3400 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5854_6
timestamp 1731220588
transform 1 0 3384 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5853_6
timestamp 1731220588
transform 1 0 3200 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5852_6
timestamp 1731220588
transform 1 0 3056 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5851_6
timestamp 1731220588
transform 1 0 2904 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5850_6
timestamp 1731220588
transform 1 0 3328 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5849_6
timestamp 1731220588
transform 1 0 3160 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5848_6
timestamp 1731220588
transform 1 0 2992 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5847_6
timestamp 1731220588
transform 1 0 2808 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5846_6
timestamp 1731220588
transform 1 0 2608 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5845_6
timestamp 1731220588
transform 1 0 3232 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5844_6
timestamp 1731220588
transform 1 0 3048 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5843_6
timestamp 1731220588
transform 1 0 2864 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5842_6
timestamp 1731220588
transform 1 0 2696 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5841_6
timestamp 1731220588
transform 1 0 3296 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5840_6
timestamp 1731220588
transform 1 0 3096 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5839_6
timestamp 1731220588
transform 1 0 2912 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5838_6
timestamp 1731220588
transform 1 0 2744 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5837_6
timestamp 1731220588
transform 1 0 2608 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5836_6
timestamp 1731220588
transform 1 0 3272 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5835_6
timestamp 1731220588
transform 1 0 3056 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5834_6
timestamp 1731220588
transform 1 0 2856 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5833_6
timestamp 1731220588
transform 1 0 2680 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5832_6
timestamp 1731220588
transform 1 0 2728 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5831_6
timestamp 1731220588
transform 1 0 3096 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5830_6
timestamp 1731220588
transform 1 0 2904 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5829_6
timestamp 1731220588
transform 1 0 2864 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5828_6
timestamp 1731220588
transform 1 0 2688 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5827_6
timestamp 1731220588
transform 1 0 3064 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5826_6
timestamp 1731220588
transform 1 0 3272 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5825_6
timestamp 1731220588
transform 1 0 3128 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5824_6
timestamp 1731220588
transform 1 0 2960 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5823_6
timestamp 1731220588
transform 1 0 2800 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5822_6
timestamp 1731220588
transform 1 0 2648 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5821_6
timestamp 1731220588
transform 1 0 2752 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5820_6
timestamp 1731220588
transform 1 0 2928 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5819_6
timestamp 1731220588
transform 1 0 3104 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5818_6
timestamp 1731220588
transform 1 0 3048 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5817_6
timestamp 1731220588
transform 1 0 2896 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5816_6
timestamp 1731220588
transform 1 0 2736 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5815_6
timestamp 1731220588
transform 1 0 2856 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5814_6
timestamp 1731220588
transform 1 0 3064 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5813_6
timestamp 1731220588
transform 1 0 3280 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5812_6
timestamp 1731220588
transform 1 0 3192 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5811_6
timestamp 1731220588
transform 1 0 3336 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5810_6
timestamp 1731220588
transform 1 0 3280 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5809_6
timestamp 1731220588
transform 1 0 3296 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5808_6
timestamp 1731220588
transform 1 0 3296 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5807_6
timestamp 1731220588
transform 1 0 3424 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5806_6
timestamp 1731220588
transform 1 0 3344 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5805_6
timestamp 1731220588
transform 1 0 3472 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5804_6
timestamp 1731220588
transform 1 0 3472 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5803_6
timestamp 1731220588
transform 1 0 3472 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5802_6
timestamp 1731220588
transform 1 0 3472 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5801_6
timestamp 1731220588
transform 1 0 3472 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5800_6
timestamp 1731220588
transform 1 0 3472 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5799_6
timestamp 1731220588
transform 1 0 3464 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5798_6
timestamp 1731220588
transform 1 0 3456 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5797_6
timestamp 1731220588
transform 1 0 3472 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5796_6
timestamp 1731220588
transform 1 0 3472 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5795_6
timestamp 1731220588
transform 1 0 3472 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5794_6
timestamp 1731220588
transform 1 0 3472 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5793_6
timestamp 1731220588
transform 1 0 3472 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5792_6
timestamp 1731220588
transform 1 0 3472 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5791_6
timestamp 1731220588
transform 1 0 3472 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5790_6
timestamp 1731220588
transform 1 0 3472 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5789_6
timestamp 1731220588
transform 1 0 3472 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5788_6
timestamp 1731220588
transform 1 0 3312 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5787_6
timestamp 1731220588
transform 1 0 3184 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5786_6
timestamp 1731220588
transform 1 0 3336 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5785_6
timestamp 1731220588
transform 1 0 3336 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5784_6
timestamp 1731220588
transform 1 0 3184 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5783_6
timestamp 1731220588
transform 1 0 3032 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5782_6
timestamp 1731220588
transform 1 0 2864 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5781_6
timestamp 1731220588
transform 1 0 2864 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5780_6
timestamp 1731220588
transform 1 0 3024 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5779_6
timestamp 1731220588
transform 1 0 3144 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5778_6
timestamp 1731220588
transform 1 0 2976 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5777_6
timestamp 1731220588
transform 1 0 2808 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5776_6
timestamp 1731220588
transform 1 0 2864 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5775_6
timestamp 1731220588
transform 1 0 3040 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5774_6
timestamp 1731220588
transform 1 0 3016 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5773_6
timestamp 1731220588
transform 1 0 2880 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5772_6
timestamp 1731220588
transform 1 0 2752 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5771_6
timestamp 1731220588
transform 1 0 2784 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5770_6
timestamp 1731220588
transform 1 0 2928 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5769_6
timestamp 1731220588
transform 1 0 3072 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5768_6
timestamp 1731220588
transform 1 0 3288 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5767_6
timestamp 1731220588
transform 1 0 3200 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5766_6
timestamp 1731220588
transform 1 0 3112 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5765_6
timestamp 1731220588
transform 1 0 3024 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5764_6
timestamp 1731220588
transform 1 0 2936 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5763_6
timestamp 1731220588
transform 1 0 2848 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5762_6
timestamp 1731220588
transform 1 0 2760 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5761_6
timestamp 1731220588
transform 1 0 2672 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5760_6
timestamp 1731220588
transform 1 0 2584 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5759_6
timestamp 1731220588
transform 1 0 2648 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5758_6
timestamp 1731220588
transform 1 0 2624 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5757_6
timestamp 1731220588
transform 1 0 2496 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5756_6
timestamp 1731220588
transform 1 0 2688 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5755_6
timestamp 1731220588
transform 1 0 2632 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5754_6
timestamp 1731220588
transform 1 0 2688 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5753_6
timestamp 1731220588
transform 1 0 2688 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5752_6
timestamp 1731220588
transform 1 0 2576 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5751_6
timestamp 1731220588
transform 1 0 2736 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5750_6
timestamp 1731220588
transform 1 0 3072 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5749_6
timestamp 1731220588
transform 1 0 2904 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5748_6
timestamp 1731220588
transform 1 0 2856 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5747_6
timestamp 1731220588
transform 1 0 2664 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5746_6
timestamp 1731220588
transform 1 0 3024 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5745_6
timestamp 1731220588
transform 1 0 3184 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5744_6
timestamp 1731220588
transform 1 0 3336 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5743_6
timestamp 1731220588
transform 1 0 3320 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5742_6
timestamp 1731220588
transform 1 0 3168 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5741_6
timestamp 1731220588
transform 1 0 3008 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5740_6
timestamp 1731220588
transform 1 0 2840 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5739_6
timestamp 1731220588
transform 1 0 2656 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5738_6
timestamp 1731220588
transform 1 0 3168 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5737_6
timestamp 1731220588
transform 1 0 3320 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5736_6
timestamp 1731220588
transform 1 0 3256 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5735_6
timestamp 1731220588
transform 1 0 3064 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5734_6
timestamp 1731220588
transform 1 0 2952 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5733_6
timestamp 1731220588
transform 1 0 2840 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5732_6
timestamp 1731220588
transform 1 0 2728 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5731_6
timestamp 1731220588
transform 1 0 2624 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5730_6
timestamp 1731220588
transform 1 0 2512 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5729_6
timestamp 1731220588
transform 1 0 2608 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5728_6
timestamp 1731220588
transform 1 0 2808 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5727_6
timestamp 1731220588
transform 1 0 3024 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5726_6
timestamp 1731220588
transform 1 0 3024 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5725_6
timestamp 1731220588
transform 1 0 2896 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5724_6
timestamp 1731220588
transform 1 0 2784 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5723_6
timestamp 1731220588
transform 1 0 2680 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5722_6
timestamp 1731220588
transform 1 0 2592 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5721_6
timestamp 1731220588
transform 1 0 2328 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5720_6
timestamp 1731220588
transform 1 0 2240 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5719_6
timestamp 1731220588
transform 1 0 2152 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5718_6
timestamp 1731220588
transform 1 0 2064 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5717_6
timestamp 1731220588
transform 1 0 1976 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5716_6
timestamp 1731220588
transform 1 0 1888 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5715_6
timestamp 1731220588
transform 1 0 2280 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5714_6
timestamp 1731220588
transform 1 0 2152 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5713_6
timestamp 1731220588
transform 1 0 2032 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5712_6
timestamp 1731220588
transform 1 0 1936 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5711_6
timestamp 1731220588
transform 1 0 2048 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5710_6
timestamp 1731220588
transform 1 0 2160 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5709_6
timestamp 1731220588
transform 1 0 2248 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5708_6
timestamp 1731220588
transform 1 0 2056 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5707_6
timestamp 1731220588
transform 1 0 1880 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5706_6
timestamp 1731220588
transform 1 0 1880 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5705_6
timestamp 1731220588
transform 1 0 2032 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5704_6
timestamp 1731220588
transform 1 0 2208 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5703_6
timestamp 1731220588
transform 1 0 2264 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5702_6
timestamp 1731220588
transform 1 0 2112 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5701_6
timestamp 1731220588
transform 1 0 1976 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5700_6
timestamp 1731220588
transform 1 0 1880 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5699_6
timestamp 1731220588
transform 1 0 1720 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5698_6
timestamp 1731220588
transform 1 0 1632 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5697_6
timestamp 1731220588
transform 1 0 1536 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5696_6
timestamp 1731220588
transform 1 0 1432 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5695_6
timestamp 1731220588
transform 1 0 1328 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5694_6
timestamp 1731220588
transform 1 0 1224 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5693_6
timestamp 1731220588
transform 1 0 1448 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5692_6
timestamp 1731220588
transform 1 0 1584 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5691_6
timestamp 1731220588
transform 1 0 1720 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5690_6
timestamp 1731220588
transform 1 0 1592 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5689_6
timestamp 1731220588
transform 1 0 1392 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5688_6
timestamp 1731220588
transform 1 0 1200 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5687_6
timestamp 1731220588
transform 1 0 1312 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5686_6
timestamp 1731220588
transform 1 0 1168 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5685_6
timestamp 1731220588
transform 1 0 1016 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5684_6
timestamp 1731220588
transform 1 0 992 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5683_6
timestamp 1731220588
transform 1 0 1112 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5682_6
timestamp 1731220588
transform 1 0 1424 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5681_6
timestamp 1731220588
transform 1 0 1296 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5680_6
timestamp 1731220588
transform 1 0 1168 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5679_6
timestamp 1731220588
transform 1 0 1040 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5678_6
timestamp 1731220588
transform 1 0 912 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5677_6
timestamp 1731220588
transform 1 0 1264 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5676_6
timestamp 1731220588
transform 1 0 1144 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5675_6
timestamp 1731220588
transform 1 0 1024 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5674_6
timestamp 1731220588
transform 1 0 912 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5673_6
timestamp 1731220588
transform 1 0 792 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5672_6
timestamp 1731220588
transform 1 0 704 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5671_6
timestamp 1731220588
transform 1 0 816 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5670_6
timestamp 1731220588
transform 1 0 1168 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5669_6
timestamp 1731220588
transform 1 0 1048 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5668_6
timestamp 1731220588
transform 1 0 928 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5667_6
timestamp 1731220588
transform 1 0 896 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5666_6
timestamp 1731220588
transform 1 0 768 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5665_6
timestamp 1731220588
transform 1 0 1016 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5664_6
timestamp 1731220588
transform 1 0 1144 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5663_6
timestamp 1731220588
transform 1 0 1272 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5662_6
timestamp 1731220588
transform 1 0 1168 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5661_6
timestamp 1731220588
transform 1 0 1048 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5660_6
timestamp 1731220588
transform 1 0 936 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5659_6
timestamp 1731220588
transform 1 0 824 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5658_6
timestamp 1731220588
transform 1 0 712 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5657_6
timestamp 1731220588
transform 1 0 792 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5656_6
timestamp 1731220588
transform 1 0 680 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5655_6
timestamp 1731220588
transform 1 0 712 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5654_6
timestamp 1731220588
transform 1 0 704 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5653_6
timestamp 1731220588
transform 1 0 752 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5652_6
timestamp 1731220588
transform 1 0 920 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5651_6
timestamp 1731220588
transform 1 0 904 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5650_6
timestamp 1731220588
transform 1 0 752 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5649_6
timestamp 1731220588
transform 1 0 880 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5648_6
timestamp 1731220588
transform 1 0 728 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5647_6
timestamp 1731220588
transform 1 0 744 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5646_6
timestamp 1731220588
transform 1 0 608 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5645_6
timestamp 1731220588
transform 1 0 576 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5644_6
timestamp 1731220588
transform 1 0 728 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5643_6
timestamp 1731220588
transform 1 0 648 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5642_6
timestamp 1731220588
transform 1 0 520 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5641_6
timestamp 1731220588
transform 1 0 776 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5640_6
timestamp 1731220588
transform 1 0 1016 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5639_6
timestamp 1731220588
transform 1 0 888 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5638_6
timestamp 1731220588
transform 1 0 704 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5637_6
timestamp 1731220588
transform 1 0 512 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5636_6
timestamp 1731220588
transform 1 0 648 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5635_6
timestamp 1731220588
transform 1 0 808 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5634_6
timestamp 1731220588
transform 1 0 744 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5633_6
timestamp 1731220588
transform 1 0 600 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5632_6
timestamp 1731220588
transform 1 0 672 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5631_6
timestamp 1731220588
transform 1 0 640 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5630_6
timestamp 1731220588
transform 1 0 776 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5629_6
timestamp 1731220588
transform 1 0 840 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5628_6
timestamp 1731220588
transform 1 0 696 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5627_6
timestamp 1731220588
transform 1 0 568 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5626_6
timestamp 1731220588
transform 1 0 632 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5625_6
timestamp 1731220588
transform 1 0 768 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5624_6
timestamp 1731220588
transform 1 0 816 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5623_6
timestamp 1731220588
transform 1 0 672 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5622_6
timestamp 1731220588
transform 1 0 632 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5621_6
timestamp 1731220588
transform 1 0 776 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5620_6
timestamp 1731220588
transform 1 0 768 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5619_6
timestamp 1731220588
transform 1 0 616 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5618_6
timestamp 1731220588
transform 1 0 656 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5617_6
timestamp 1731220588
transform 1 0 832 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5616_6
timestamp 1731220588
transform 1 0 672 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5615_6
timestamp 1731220588
transform 1 0 856 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5614_6
timestamp 1731220588
transform 1 0 864 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5613_6
timestamp 1731220588
transform 1 0 672 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5612_6
timestamp 1731220588
transform 1 0 584 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5611_6
timestamp 1731220588
transform 1 0 760 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5610_6
timestamp 1731220588
transform 1 0 776 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5609_6
timestamp 1731220588
transform 1 0 624 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5608_6
timestamp 1731220588
transform 1 0 480 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5607_6
timestamp 1731220588
transform 1 0 616 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5606_6
timestamp 1731220588
transform 1 0 752 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5605_6
timestamp 1731220588
transform 1 0 776 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5604_6
timestamp 1731220588
transform 1 0 688 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5603_6
timestamp 1731220588
transform 1 0 600 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5602_6
timestamp 1731220588
transform 1 0 512 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5601_6
timestamp 1731220588
transform 1 0 424 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5600_6
timestamp 1731220588
transform 1 0 336 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5599_6
timestamp 1731220588
transform 1 0 248 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5598_6
timestamp 1731220588
transform 1 0 160 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5597_6
timestamp 1731220588
transform 1 0 224 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5596_6
timestamp 1731220588
transform 1 0 480 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5595_6
timestamp 1731220588
transform 1 0 352 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5594_6
timestamp 1731220588
transform 1 0 336 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5593_6
timestamp 1731220588
transform 1 0 200 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5592_6
timestamp 1731220588
transform 1 0 128 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5591_6
timestamp 1731220588
transform 1 0 256 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5590_6
timestamp 1731220588
transform 1 0 416 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5589_6
timestamp 1731220588
transform 1 0 480 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5588_6
timestamp 1731220588
transform 1 0 288 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5587_6
timestamp 1731220588
transform 1 0 128 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5586_6
timestamp 1731220588
transform 1 0 128 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5585_6
timestamp 1731220588
transform 1 0 296 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5584_6
timestamp 1731220588
transform 1 0 488 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5583_6
timestamp 1731220588
transform 1 0 472 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5582_6
timestamp 1731220588
transform 1 0 288 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5581_6
timestamp 1731220588
transform 1 0 128 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5580_6
timestamp 1731220588
transform 1 0 128 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5579_6
timestamp 1731220588
transform 1 0 288 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5578_6
timestamp 1731220588
transform 1 0 456 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5577_6
timestamp 1731220588
transform 1 0 488 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5576_6
timestamp 1731220588
transform 1 0 344 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5575_6
timestamp 1731220588
transform 1 0 200 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5574_6
timestamp 1731220588
transform 1 0 280 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5573_6
timestamp 1731220588
transform 1 0 528 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5572_6
timestamp 1731220588
transform 1 0 400 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5571_6
timestamp 1731220588
transform 1 0 328 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5570_6
timestamp 1731220588
transform 1 0 416 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5569_6
timestamp 1731220588
transform 1 0 520 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5568_6
timestamp 1731220588
transform 1 0 456 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5567_6
timestamp 1731220588
transform 1 0 360 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5566_6
timestamp 1731220588
transform 1 0 328 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5565_6
timestamp 1731220588
transform 1 0 416 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5564_6
timestamp 1731220588
transform 1 0 520 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5563_6
timestamp 1731220588
transform 1 0 552 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5562_6
timestamp 1731220588
transform 1 0 432 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5561_6
timestamp 1731220588
transform 1 0 320 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5560_6
timestamp 1731220588
transform 1 0 208 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5559_6
timestamp 1731220588
transform 1 0 152 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5558_6
timestamp 1731220588
transform 1 0 304 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5557_6
timestamp 1731220588
transform 1 0 456 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5556_6
timestamp 1731220588
transform 1 0 472 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5555_6
timestamp 1731220588
transform 1 0 288 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5554_6
timestamp 1731220588
transform 1 0 128 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5553_6
timestamp 1731220588
transform 1 0 312 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5552_6
timestamp 1731220588
transform 1 0 128 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5551_6
timestamp 1731220588
transform 1 0 128 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5550_6
timestamp 1731220588
transform 1 0 320 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5549_6
timestamp 1731220588
transform 1 0 544 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5548_6
timestamp 1731220588
transform 1 0 384 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5547_6
timestamp 1731220588
transform 1 0 248 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5546_6
timestamp 1731220588
transform 1 0 128 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5545_6
timestamp 1731220588
transform 1 0 128 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5544_6
timestamp 1731220588
transform 1 0 264 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5543_6
timestamp 1731220588
transform 1 0 416 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5542_6
timestamp 1731220588
transform 1 0 472 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5541_6
timestamp 1731220588
transform 1 0 336 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5540_6
timestamp 1731220588
transform 1 0 208 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5539_6
timestamp 1731220588
transform 1 0 304 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5538_6
timestamp 1731220588
transform 1 0 440 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5537_6
timestamp 1731220588
transform 1 0 584 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5536_6
timestamp 1731220588
transform 1 0 456 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5535_6
timestamp 1731220588
transform 1 0 312 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5534_6
timestamp 1731220588
transform 1 0 600 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5533_6
timestamp 1731220588
transform 1 0 584 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5532_6
timestamp 1731220588
transform 1 0 408 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5531_6
timestamp 1731220588
transform 1 0 240 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5530_6
timestamp 1731220588
transform 1 0 208 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5529_6
timestamp 1731220588
transform 1 0 464 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5528_6
timestamp 1731220588
transform 1 0 288 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5527_6
timestamp 1731220588
transform 1 0 152 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5526_6
timestamp 1731220588
transform 1 0 152 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5525_6
timestamp 1731220588
transform 1 0 128 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5524_6
timestamp 1731220588
transform 1 0 224 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5523_6
timestamp 1731220588
transform 1 0 232 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5522_6
timestamp 1731220588
transform 1 0 128 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5521_6
timestamp 1731220588
transform 1 0 128 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5520_6
timestamp 1731220588
transform 1 0 224 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5519_6
timestamp 1731220588
transform 1 0 344 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5518_6
timestamp 1731220588
transform 1 0 248 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5517_6
timestamp 1731220588
transform 1 0 128 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5516_6
timestamp 1731220588
transform 1 0 144 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5515_6
timestamp 1731220588
transform 1 0 312 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5514_6
timestamp 1731220588
transform 1 0 448 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5513_6
timestamp 1731220588
transform 1 0 304 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5512_6
timestamp 1731220588
transform 1 0 168 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5511_6
timestamp 1731220588
transform 1 0 264 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5510_6
timestamp 1731220588
transform 1 0 464 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5509_6
timestamp 1731220588
transform 1 0 480 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5508_6
timestamp 1731220588
transform 1 0 336 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5507_6
timestamp 1731220588
transform 1 0 208 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5506_6
timestamp 1731220588
transform 1 0 160 0 -1 2708
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5505_6
timestamp 1731220588
transform 1 0 272 0 -1 2708
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5504_6
timestamp 1731220588
transform 1 0 384 0 -1 2708
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5503_6
timestamp 1731220588
transform 1 0 400 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5502_6
timestamp 1731220588
transform 1 0 280 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5501_6
timestamp 1731220588
transform 1 0 176 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5500_6
timestamp 1731220588
transform 1 0 128 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5499_6
timestamp 1731220588
transform 1 0 216 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5498_6
timestamp 1731220588
transform 1 0 304 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5497_6
timestamp 1731220588
transform 1 0 392 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5496_6
timestamp 1731220588
transform 1 0 480 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5495_6
timestamp 1731220588
transform 1 0 592 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5494_6
timestamp 1731220588
transform 1 0 720 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5493_6
timestamp 1731220588
transform 1 0 992 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5492_6
timestamp 1731220588
transform 1 0 856 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5491_6
timestamp 1731220588
transform 1 0 808 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5490_6
timestamp 1731220588
transform 1 0 672 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5489_6
timestamp 1731220588
transform 1 0 536 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5488_6
timestamp 1731220588
transform 1 0 496 0 -1 2708
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5487_6
timestamp 1731220588
transform 1 0 608 0 -1 2708
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5486_6
timestamp 1731220588
transform 1 0 648 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5485_6
timestamp 1731220588
transform 1 0 824 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5484_6
timestamp 1731220588
transform 1 0 1008 0 1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5483_6
timestamp 1731220588
transform 1 0 848 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5482_6
timestamp 1731220588
transform 1 0 664 0 -1 2556
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5481_6
timestamp 1731220588
transform 1 0 864 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5480_6
timestamp 1731220588
transform 1 0 728 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5479_6
timestamp 1731220588
transform 1 0 592 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5478_6
timestamp 1731220588
transform 1 0 472 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5477_6
timestamp 1731220588
transform 1 0 632 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5476_6
timestamp 1731220588
transform 1 0 776 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5475_6
timestamp 1731220588
transform 1 0 664 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5474_6
timestamp 1731220588
transform 1 0 528 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5473_6
timestamp 1731220588
transform 1 0 392 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5472_6
timestamp 1731220588
transform 1 0 464 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5471_6
timestamp 1731220588
transform 1 0 584 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5470_6
timestamp 1731220588
transform 1 0 640 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5469_6
timestamp 1731220588
transform 1 0 504 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5468_6
timestamp 1731220588
transform 1 0 368 0 1 2128
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5467_6
timestamp 1731220588
transform 1 0 352 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5466_6
timestamp 1731220588
transform 1 0 472 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5465_6
timestamp 1731220588
transform 1 0 592 0 -1 2120
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5464_6
timestamp 1731220588
transform 1 0 560 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5463_6
timestamp 1731220588
transform 1 0 432 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5462_6
timestamp 1731220588
transform 1 0 296 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5461_6
timestamp 1731220588
transform 1 0 432 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5460_6
timestamp 1731220588
transform 1 0 576 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5459_6
timestamp 1731220588
transform 1 0 848 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5458_6
timestamp 1731220588
transform 1 0 984 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5457_6
timestamp 1731220588
transform 1 0 896 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5456_6
timestamp 1731220588
transform 1 0 1000 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5455_6
timestamp 1731220588
transform 1 0 1104 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5454_6
timestamp 1731220588
transform 1 0 1208 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5453_6
timestamp 1731220588
transform 1 0 1312 0 1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5452_6
timestamp 1731220588
transform 1 0 1232 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5451_6
timestamp 1731220588
transform 1 0 1112 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5450_6
timestamp 1731220588
transform 1 0 1352 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5449_6
timestamp 1731220588
transform 1 0 1472 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5448_6
timestamp 1731220588
transform 1 0 1592 0 -1 1972
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5447_6
timestamp 1731220588
transform 1 0 1592 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5446_6
timestamp 1731220588
transform 1 0 1440 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5445_6
timestamp 1731220588
transform 1 0 1280 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5444_6
timestamp 1731220588
transform 1 0 1112 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5443_6
timestamp 1731220588
transform 1 0 920 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5442_6
timestamp 1731220588
transform 1 0 1072 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5441_6
timestamp 1731220588
transform 1 0 1216 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5440_6
timestamp 1731220588
transform 1 0 1352 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5439_6
timestamp 1731220588
transform 1 0 1360 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5438_6
timestamp 1731220588
transform 1 0 1208 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5437_6
timestamp 1731220588
transform 1 0 1056 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5436_6
timestamp 1731220588
transform 1 0 1032 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5435_6
timestamp 1731220588
transform 1 0 1184 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5434_6
timestamp 1731220588
transform 1 0 1200 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5433_6
timestamp 1731220588
transform 1 0 1040 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5432_6
timestamp 1731220588
transform 1 0 888 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5431_6
timestamp 1731220588
transform 1 0 880 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5430_6
timestamp 1731220588
transform 1 0 1032 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5429_6
timestamp 1731220588
transform 1 0 1008 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5428_6
timestamp 1731220588
transform 1 0 896 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5427_6
timestamp 1731220588
transform 1 0 776 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5426_6
timestamp 1731220588
transform 1 0 1128 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5425_6
timestamp 1731220588
transform 1 0 1248 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5424_6
timestamp 1731220588
transform 1 0 1488 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5423_6
timestamp 1731220588
transform 1 0 1368 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5422_6
timestamp 1731220588
transform 1 0 1336 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5421_6
timestamp 1731220588
transform 1 0 1184 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5420_6
timestamp 1731220588
transform 1 0 1488 0 -1 1536
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5419_6
timestamp 1731220588
transform 1 0 1528 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5418_6
timestamp 1731220588
transform 1 0 1360 0 1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5417_6
timestamp 1731220588
transform 1 0 1336 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5416_6
timestamp 1731220588
transform 1 0 1488 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5415_6
timestamp 1731220588
transform 1 0 1640 0 -1 1684
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5414_6
timestamp 1731220588
transform 1 0 1672 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5413_6
timestamp 1731220588
transform 1 0 1512 0 1 1688
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5412_6
timestamp 1731220588
transform 1 0 1480 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5411_6
timestamp 1731220588
transform 1 0 1608 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5410_6
timestamp 1731220588
transform 1 0 1720 0 -1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5409_6
timestamp 1731220588
transform 1 0 1720 0 1 1828
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5408_6
timestamp 1731220588
transform 1 0 1880 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5407_6
timestamp 1731220588
transform 1 0 2056 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5406_6
timestamp 1731220588
transform 1 0 1968 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5405_6
timestamp 1731220588
transform 1 0 1896 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5404_6
timestamp 1731220588
transform 1 0 2432 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5403_6
timestamp 1731220588
transform 1 0 2280 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5402_6
timestamp 1731220588
transform 1 0 2152 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5401_6
timestamp 1731220588
transform 1 0 1992 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5400_6
timestamp 1731220588
transform 1 0 1928 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5399_6
timestamp 1731220588
transform 1 0 2072 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5398_6
timestamp 1731220588
transform 1 0 2232 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5397_6
timestamp 1731220588
transform 1 0 2144 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5396_6
timestamp 1731220588
transform 1 0 2024 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5395_6
timestamp 1731220588
transform 1 0 1904 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5394_6
timestamp 1731220588
transform 1 0 1880 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5393_6
timestamp 1731220588
transform 1 0 2000 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5392_6
timestamp 1731220588
transform 1 0 2136 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5391_6
timestamp 1731220588
transform 1 0 2016 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5390_6
timestamp 1731220588
transform 1 0 1880 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5389_6
timestamp 1731220588
transform 1 0 1720 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5388_6
timestamp 1731220588
transform 1 0 1616 0 1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5387_6
timestamp 1731220588
transform 1 0 1496 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5386_6
timestamp 1731220588
transform 1 0 1256 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5385_6
timestamp 1731220588
transform 1 0 1720 0 -1 1392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5384_6
timestamp 1731220588
transform 1 0 1672 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5383_6
timestamp 1731220588
transform 1 0 1520 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5382_6
timestamp 1731220588
transform 1 0 1368 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5381_6
timestamp 1731220588
transform 1 0 1216 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5380_6
timestamp 1731220588
transform 1 0 1056 0 1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5379_6
timestamp 1731220588
transform 1 0 1520 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5378_6
timestamp 1731220588
transform 1 0 1376 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5377_6
timestamp 1731220588
transform 1 0 1240 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5376_6
timestamp 1731220588
transform 1 0 1104 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5375_6
timestamp 1731220588
transform 1 0 960 0 -1 1244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5374_6
timestamp 1731220588
transform 1 0 1560 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5373_6
timestamp 1731220588
transform 1 0 1384 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5372_6
timestamp 1731220588
transform 1 0 1216 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5371_6
timestamp 1731220588
transform 1 0 1048 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5370_6
timestamp 1731220588
transform 1 0 896 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5369_6
timestamp 1731220588
transform 1 0 1400 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5368_6
timestamp 1731220588
transform 1 0 1240 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5367_6
timestamp 1731220588
transform 1 0 1080 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5366_6
timestamp 1731220588
transform 1 0 936 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5365_6
timestamp 1731220588
transform 1 0 800 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5364_6
timestamp 1731220588
transform 1 0 936 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5363_6
timestamp 1731220588
transform 1 0 1120 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5362_6
timestamp 1731220588
transform 1 0 1312 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5361_6
timestamp 1731220588
transform 1 0 1168 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5360_6
timestamp 1731220588
transform 1 0 1000 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5359_6
timestamp 1731220588
transform 1 0 912 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5358_6
timestamp 1731220588
transform 1 0 1072 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5357_6
timestamp 1731220588
transform 1 0 1248 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5356_6
timestamp 1731220588
transform 1 0 1120 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5355_6
timestamp 1731220588
transform 1 0 968 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5354_6
timestamp 1731220588
transform 1 0 920 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5353_6
timestamp 1731220588
transform 1 0 1232 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5352_6
timestamp 1731220588
transform 1 0 1072 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5351_6
timestamp 1731220588
transform 1 0 1064 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5350_6
timestamp 1731220588
transform 1 0 920 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5349_6
timestamp 1731220588
transform 1 0 1008 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5348_6
timestamp 1731220588
transform 1 0 1024 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5347_6
timestamp 1731220588
transform 1 0 1040 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5346_6
timestamp 1731220588
transform 1 0 1096 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5345_6
timestamp 1731220588
transform 1 0 928 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5344_6
timestamp 1731220588
transform 1 0 920 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5343_6
timestamp 1731220588
transform 1 0 1064 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5342_6
timestamp 1731220588
transform 1 0 1024 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5341_6
timestamp 1731220588
transform 1 0 888 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5340_6
timestamp 1731220588
transform 1 0 864 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5339_6
timestamp 1731220588
transform 1 0 952 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5338_6
timestamp 1731220588
transform 1 0 1040 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5337_6
timestamp 1731220588
transform 1 0 1128 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5336_6
timestamp 1731220588
transform 1 0 1216 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5335_6
timestamp 1731220588
transform 1 0 1488 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5334_6
timestamp 1731220588
transform 1 0 1392 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5333_6
timestamp 1731220588
transform 1 0 1304 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5332_6
timestamp 1731220588
transform 1 0 1288 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5331_6
timestamp 1731220588
transform 1 0 1152 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5330_6
timestamp 1731220588
transform 1 0 1424 0 -1 244
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5329_6
timestamp 1731220588
transform 1 0 1472 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5328_6
timestamp 1731220588
transform 1 0 1344 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5327_6
timestamp 1731220588
transform 1 0 1208 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5326_6
timestamp 1731220588
transform 1 0 1256 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5325_6
timestamp 1731220588
transform 1 0 1208 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5324_6
timestamp 1731220588
transform 1 0 1376 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5323_6
timestamp 1731220588
transform 1 0 1344 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5322_6
timestamp 1731220588
transform 1 0 1184 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5321_6
timestamp 1731220588
transform 1 0 1184 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5320_6
timestamp 1731220588
transform 1 0 1360 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5319_6
timestamp 1731220588
transform 1 0 1336 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5318_6
timestamp 1731220588
transform 1 0 1200 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5317_6
timestamp 1731220588
transform 1 0 1472 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5316_6
timestamp 1731220588
transform 1 0 1568 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5315_6
timestamp 1731220588
transform 1 0 1400 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5314_6
timestamp 1731220588
transform 1 0 1272 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5313_6
timestamp 1731220588
transform 1 0 1592 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5312_6
timestamp 1731220588
transform 1 0 1432 0 -1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5311_6
timestamp 1731220588
transform 1 0 1432 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5310_6
timestamp 1731220588
transform 1 0 1616 0 1 812
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5309_6
timestamp 1731220588
transform 1 0 1520 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5308_6
timestamp 1731220588
transform 1 0 1344 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5307_6
timestamp 1731220588
transform 1 0 1704 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5306_6
timestamp 1731220588
transform 1 0 1720 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5305_6
timestamp 1731220588
transform 1 0 1520 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5304_6
timestamp 1731220588
transform 1 0 1568 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5303_6
timestamp 1731220588
transform 1 0 1720 0 -1 1100
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5302_6
timestamp 1731220588
transform 1 0 1720 0 1 1104
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5301_6
timestamp 1731220588
transform 1 0 1880 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5300_6
timestamp 1731220588
transform 1 0 1896 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5299_6
timestamp 1731220588
transform 1 0 1984 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5298_6
timestamp 1731220588
transform 1 0 2208 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5297_6
timestamp 1731220588
transform 1 0 2344 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5296_6
timestamp 1731220588
transform 1 0 2624 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5295_6
timestamp 1731220588
transform 1 0 2480 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5294_6
timestamp 1731220588
transform 1 0 2424 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5293_6
timestamp 1731220588
transform 1 0 2400 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5292_6
timestamp 1731220588
transform 1 0 2240 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5291_6
timestamp 1731220588
transform 1 0 2424 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5290_6
timestamp 1731220588
transform 1 0 2296 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5289_6
timestamp 1731220588
transform 1 0 2176 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5288_6
timestamp 1731220588
transform 1 0 2056 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5287_6
timestamp 1731220588
transform 1 0 2192 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5286_6
timestamp 1731220588
transform 1 0 2344 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5285_6
timestamp 1731220588
transform 1 0 2472 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5284_6
timestamp 1731220588
transform 1 0 2304 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5283_6
timestamp 1731220588
transform 1 0 2152 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5282_6
timestamp 1731220588
transform 1 0 2128 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5281_6
timestamp 1731220588
transform 1 0 1984 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5280_6
timestamp 1731220588
transform 1 0 2280 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5279_6
timestamp 1731220588
transform 1 0 2448 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5278_6
timestamp 1731220588
transform 1 0 2432 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5277_6
timestamp 1731220588
transform 1 0 2240 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5276_6
timestamp 1731220588
transform 1 0 2048 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5275_6
timestamp 1731220588
transform 1 0 2208 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5274_6
timestamp 1731220588
transform 1 0 2352 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5273_6
timestamp 1731220588
transform 1 0 2504 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5272_6
timestamp 1731220588
transform 1 0 2448 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5271_6
timestamp 1731220588
transform 1 0 2360 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5270_6
timestamp 1731220588
transform 1 0 2272 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5269_6
timestamp 1731220588
transform 1 0 2184 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5268_6
timestamp 1731220588
transform 1 0 2296 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5267_6
timestamp 1731220588
transform 1 0 2392 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5266_6
timestamp 1731220588
transform 1 0 2496 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5265_6
timestamp 1731220588
transform 1 0 2600 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5264_6
timestamp 1731220588
transform 1 0 2680 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5263_6
timestamp 1731220588
transform 1 0 2544 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5262_6
timestamp 1731220588
transform 1 0 2416 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5261_6
timestamp 1731220588
transform 1 0 2312 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5260_6
timestamp 1731220588
transform 1 0 2224 0 1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5259_6
timestamp 1731220588
transform 1 0 2520 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5258_6
timestamp 1731220588
transform 1 0 2392 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5257_6
timestamp 1731220588
transform 1 0 2280 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5256_6
timestamp 1731220588
transform 1 0 2176 0 -1 392
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5255_6
timestamp 1731220588
transform 1 0 2072 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5254_6
timestamp 1731220588
transform 1 0 2288 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5253_6
timestamp 1731220588
transform 1 0 2288 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5252_6
timestamp 1731220588
transform 1 0 2448 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5251_6
timestamp 1731220588
transform 1 0 2528 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5250_6
timestamp 1731220588
transform 1 0 2424 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5249_6
timestamp 1731220588
transform 1 0 2320 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5248_6
timestamp 1731220588
transform 1 0 2232 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5247_6
timestamp 1731220588
transform 1 0 2144 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5246_6
timestamp 1731220588
transform 1 0 2056 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5245_6
timestamp 1731220588
transform 1 0 1968 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5244_6
timestamp 1731220588
transform 1 0 1880 0 1 84
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5243_6
timestamp 1731220588
transform 1 0 2136 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5242_6
timestamp 1731220588
transform 1 0 1992 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5241_6
timestamp 1731220588
transform 1 0 1880 0 -1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5240_6
timestamp 1731220588
transform 1 0 1880 0 1 248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5239_6
timestamp 1731220588
transform 1 0 1720 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5238_6
timestamp 1731220588
transform 1 0 1608 0 1 252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5237_6
timestamp 1731220588
transform 1 0 1576 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5236_6
timestamp 1731220588
transform 1 0 1416 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5235_6
timestamp 1731220588
transform 1 0 1720 0 -1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5234_6
timestamp 1731220588
transform 1 0 1712 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5233_6
timestamp 1731220588
transform 1 0 1544 0 1 388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5232_6
timestamp 1731220588
transform 1 0 1496 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5231_6
timestamp 1731220588
transform 1 0 1656 0 -1 528
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5230_6
timestamp 1731220588
transform 1 0 1720 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5229_6
timestamp 1731220588
transform 1 0 1544 0 1 532
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5228_6
timestamp 1731220588
transform 1 0 1608 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5227_6
timestamp 1731220588
transform 1 0 1720 0 -1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5226_6
timestamp 1731220588
transform 1 0 1720 0 1 672
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5225_6
timestamp 1731220588
transform 1 0 1880 0 1 676
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5224_6
timestamp 1731220588
transform 1 0 1880 0 -1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5223_6
timestamp 1731220588
transform 1 0 1880 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5222_6
timestamp 1731220588
transform 1 0 2000 0 1 816
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5221_6
timestamp 1731220588
transform 1 0 2040 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5220_6
timestamp 1731220588
transform 1 0 1880 0 -1 952
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5219_6
timestamp 1731220588
transform 1 0 1928 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5218_6
timestamp 1731220588
transform 1 0 1928 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5217_6
timestamp 1731220588
transform 1 0 2088 0 -1 1096
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5216_6
timestamp 1731220588
transform 1 0 2240 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5215_6
timestamp 1731220588
transform 1 0 2048 0 1 1108
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5214_6
timestamp 1731220588
transform 1 0 2088 0 -1 1248
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5213_6
timestamp 1731220588
transform 1 0 2072 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5212_6
timestamp 1731220588
transform 1 0 2504 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5211_6
timestamp 1731220588
transform 1 0 2296 0 1 1252
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5210_6
timestamp 1731220588
transform 1 0 2256 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5209_6
timestamp 1731220588
transform 1 0 2072 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5208_6
timestamp 1731220588
transform 1 0 2608 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5207_6
timestamp 1731220588
transform 1 0 2432 0 -1 1388
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5206_6
timestamp 1731220588
transform 1 0 2344 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5205_6
timestamp 1731220588
transform 1 0 2168 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5204_6
timestamp 1731220588
transform 1 0 2512 0 1 1396
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5203_6
timestamp 1731220588
transform 1 0 2496 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5202_6
timestamp 1731220588
transform 1 0 2336 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5201_6
timestamp 1731220588
transform 1 0 2176 0 -1 1540
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5200_6
timestamp 1731220588
transform 1 0 2272 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5199_6
timestamp 1731220588
transform 1 0 2416 0 1 1548
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5198_6
timestamp 1731220588
transform 1 0 2392 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5197_6
timestamp 1731220588
transform 1 0 2264 0 -1 1692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5196_6
timestamp 1731220588
transform 1 0 2584 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5195_6
timestamp 1731220588
transform 1 0 2400 0 1 1696
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5194_6
timestamp 1731220588
transform 1 0 2216 0 -1 1836
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5193_6
timestamp 1731220588
transform 1 0 2752 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5192_6
timestamp 1731220588
transform 1 0 2592 0 1 1840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5191_6
timestamp 1731220588
transform 1 0 2392 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5190_6
timestamp 1731220588
transform 1 0 2152 0 -1 1976
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5189_6
timestamp 1731220588
transform 1 0 2112 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5188_6
timestamp 1731220588
transform 1 0 1984 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5187_6
timestamp 1731220588
transform 1 0 2536 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5186_6
timestamp 1731220588
transform 1 0 2384 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5185_6
timestamp 1731220588
transform 1 0 2240 0 1 1984
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5184_6
timestamp 1731220588
transform 1 0 2232 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5183_6
timestamp 1731220588
transform 1 0 2144 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5182_6
timestamp 1731220588
transform 1 0 2496 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5181_6
timestamp 1731220588
transform 1 0 2408 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5180_6
timestamp 1731220588
transform 1 0 2320 0 -1 2124
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5179_6
timestamp 1731220588
transform 1 0 2240 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5178_6
timestamp 1731220588
transform 1 0 2328 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5177_6
timestamp 1731220588
transform 1 0 2424 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5176_6
timestamp 1731220588
transform 1 0 2536 0 1 2132
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5175_6
timestamp 1731220588
transform 1 0 2576 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5174_6
timestamp 1731220588
transform 1 0 2440 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5173_6
timestamp 1731220588
transform 1 0 2328 0 -1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5172_6
timestamp 1731220588
transform 1 0 2336 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5171_6
timestamp 1731220588
transform 1 0 2432 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5170_6
timestamp 1731220588
transform 1 0 2544 0 1 2268
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5169_6
timestamp 1731220588
transform 1 0 2496 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5168_6
timestamp 1731220588
transform 1 0 2344 0 -1 2408
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5167_6
timestamp 1731220588
transform 1 0 2424 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5166_6
timestamp 1731220588
transform 1 0 2584 0 1 2416
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5165_6
timestamp 1731220588
transform 1 0 2568 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5164_6
timestamp 1731220588
transform 1 0 2392 0 -1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5163_6
timestamp 1731220588
transform 1 0 2648 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5162_6
timestamp 1731220588
transform 1 0 2448 0 1 2552
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5161_6
timestamp 1731220588
transform 1 0 2400 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5160_6
timestamp 1731220588
transform 1 0 2280 0 -1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5159_6
timestamp 1731220588
transform 1 0 2432 0 1 2692
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5158_6
timestamp 1731220588
transform 1 0 2416 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5157_6
timestamp 1731220588
transform 1 0 2504 0 -1 2840
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5156_6
timestamp 1731220588
transform 1 0 2448 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5155_6
timestamp 1731220588
transform 1 0 2224 0 1 2844
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5154_6
timestamp 1731220588
transform 1 0 2232 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5153_6
timestamp 1731220588
transform 1 0 2456 0 -1 2996
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5152_6
timestamp 1731220588
transform 1 0 2408 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5151_6
timestamp 1731220588
transform 1 0 2240 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5150_6
timestamp 1731220588
transform 1 0 2288 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5149_6
timestamp 1731220588
transform 1 0 2496 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5148_6
timestamp 1731220588
transform 1 0 2496 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5147_6
timestamp 1731220588
transform 1 0 2288 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5146_6
timestamp 1731220588
transform 1 0 2256 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5145_6
timestamp 1731220588
transform 1 0 2448 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5144_6
timestamp 1731220588
transform 1 0 2520 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5143_6
timestamp 1731220588
transform 1 0 2352 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5142_6
timestamp 1731220588
transform 1 0 2192 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5141_6
timestamp 1731220588
transform 1 0 2216 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5140_6
timestamp 1731220588
transform 1 0 2360 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5139_6
timestamp 1731220588
transform 1 0 2248 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5138_6
timestamp 1731220588
transform 1 0 2376 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5137_6
timestamp 1731220588
transform 1 0 2512 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5136_6
timestamp 1731220588
transform 1 0 2496 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5135_6
timestamp 1731220588
transform 1 0 2408 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5134_6
timestamp 1731220588
transform 1 0 2320 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5133_6
timestamp 1731220588
transform 1 0 2232 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5132_6
timestamp 1731220588
transform 1 0 2144 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5131_6
timestamp 1731220588
transform 1 0 2056 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5130_6
timestamp 1731220588
transform 1 0 1968 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5129_6
timestamp 1731220588
transform 1 0 1880 0 -1 3584
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5128_6
timestamp 1731220588
transform 1 0 1896 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5127_6
timestamp 1731220588
transform 1 0 2000 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5126_6
timestamp 1731220588
transform 1 0 2120 0 1 3440
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5125_6
timestamp 1731220588
transform 1 0 2064 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5124_6
timestamp 1731220588
transform 1 0 1904 0 -1 3432
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5123_6
timestamp 1731220588
transform 1 0 1880 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5122_6
timestamp 1731220588
transform 1 0 2032 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5121_6
timestamp 1731220588
transform 1 0 2056 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5120_6
timestamp 1731220588
transform 1 0 1880 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5119_6
timestamp 1731220588
transform 1 0 1880 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5118_6
timestamp 1731220588
transform 1 0 2072 0 1 3152
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5117_6
timestamp 1731220588
transform 1 0 2072 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5116_6
timestamp 1731220588
transform 1 0 1880 0 -1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5115_6
timestamp 1731220588
transform 1 0 1720 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5114_6
timestamp 1731220588
transform 1 0 1632 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5113_6
timestamp 1731220588
transform 1 0 1624 0 -1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5112_6
timestamp 1731220588
transform 1 0 1720 0 -1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5111_6
timestamp 1731220588
transform 1 0 1688 0 1 2856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5110_6
timestamp 1731220588
transform 1 0 1616 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5109_6
timestamp 1731220588
transform 1 0 1496 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5108_6
timestamp 1731220588
transform 1 0 1720 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5107_6
timestamp 1731220588
transform 1 0 1720 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5106_6
timestamp 1731220588
transform 1 0 1632 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5105_6
timestamp 1731220588
transform 1 0 1520 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5104_6
timestamp 1731220588
transform 1 0 1416 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5103_6
timestamp 1731220588
transform 1 0 1304 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5102_6
timestamp 1731220588
transform 1 0 1192 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5101_6
timestamp 1731220588
transform 1 0 1072 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_5100_6
timestamp 1731220588
transform 1 0 944 0 1 2716
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_599_6
timestamp 1731220588
transform 1 0 1128 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_598_6
timestamp 1731220588
transform 1 0 1256 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_597_6
timestamp 1731220588
transform 1 0 1376 0 -1 2852
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_596_6
timestamp 1731220588
transform 1 0 1344 0 1 2856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_595_6
timestamp 1731220588
transform 1 0 1568 0 1 2856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_594_6
timestamp 1731220588
transform 1 0 1456 0 1 2856
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_593_6
timestamp 1731220588
transform 1 0 1400 0 -1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_592_6
timestamp 1731220588
transform 1 0 1512 0 -1 2992
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_591_6
timestamp 1731220588
transform 1 0 1456 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_590_6
timestamp 1731220588
transform 1 0 1544 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_589_6
timestamp 1731220588
transform 1 0 1512 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_588_6
timestamp 1731220588
transform 1 0 1368 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_587_6
timestamp 1731220588
transform 1 0 1368 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_586_6
timestamp 1731220588
transform 1 0 1520 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_585_6
timestamp 1731220588
transform 1 0 1512 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_584_6
timestamp 1731220588
transform 1 0 1336 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_583_6
timestamp 1731220588
transform 1 0 1264 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_582_6
timestamp 1731220588
transform 1 0 1400 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_581_6
timestamp 1731220588
transform 1 0 1544 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_580_6
timestamp 1731220588
transform 1 0 1472 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_579_6
timestamp 1731220588
transform 1 0 1288 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_578_6
timestamp 1731220588
transform 1 0 1560 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_577_6
timestamp 1731220588
transform 1 0 1440 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_576_6
timestamp 1731220588
transform 1 0 1320 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_575_6
timestamp 1731220588
transform 1 0 1200 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_574_6
timestamp 1731220588
transform 1 0 1536 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_573_6
timestamp 1731220588
transform 1 0 1416 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_572_6
timestamp 1731220588
transform 1 0 1304 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_571_6
timestamp 1731220588
transform 1 0 1192 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_570_6
timestamp 1731220588
transform 1 0 1072 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_569_6
timestamp 1731220588
transform 1 0 944 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_568_6
timestamp 1731220588
transform 1 0 816 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_567_6
timestamp 1731220588
transform 1 0 816 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_566_6
timestamp 1731220588
transform 1 0 1080 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_565_6
timestamp 1731220588
transform 1 0 952 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_564_6
timestamp 1731220588
transform 1 0 928 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_563_6
timestamp 1731220588
transform 1 0 1104 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_562_6
timestamp 1731220588
transform 1 0 1128 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_561_6
timestamp 1731220588
transform 1 0 984 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_560_6
timestamp 1731220588
transform 1 0 840 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_559_6
timestamp 1731220588
transform 1 0 984 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_558_6
timestamp 1731220588
transform 1 0 1160 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_557_6
timestamp 1731220588
transform 1 0 1216 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_556_6
timestamp 1731220588
transform 1 0 1064 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_555_6
timestamp 1731220588
transform 1 0 920 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_554_6
timestamp 1731220588
transform 1 0 1088 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_553_6
timestamp 1731220588
transform 1 0 1224 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_552_6
timestamp 1731220588
transform 1 0 1368 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_551_6
timestamp 1731220588
transform 1 0 1280 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_550_6
timestamp 1731220588
transform 1 0 1192 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_549_6
timestamp 1731220588
transform 1 0 1104 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_548_6
timestamp 1731220588
transform 1 0 1016 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_547_6
timestamp 1731220588
transform 1 0 928 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_546_6
timestamp 1731220588
transform 1 0 840 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_545_6
timestamp 1731220588
transform 1 0 752 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_544_6
timestamp 1731220588
transform 1 0 664 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_543_6
timestamp 1731220588
transform 1 0 576 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_542_6
timestamp 1731220588
transform 1 0 488 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_541_6
timestamp 1731220588
transform 1 0 400 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_540_6
timestamp 1731220588
transform 1 0 312 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_539_6
timestamp 1731220588
transform 1 0 224 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_538_6
timestamp 1731220588
transform 1 0 136 0 1 3000
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_537_6
timestamp 1731220588
transform 1 0 960 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_536_6
timestamp 1731220588
transform 1 0 840 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_535_6
timestamp 1731220588
transform 1 0 728 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_534_6
timestamp 1731220588
transform 1 0 632 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_533_6
timestamp 1731220588
transform 1 0 544 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_532_6
timestamp 1731220588
transform 1 0 456 0 -1 3144
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_531_6
timestamp 1731220588
transform 1 0 784 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_530_6
timestamp 1731220588
transform 1 0 656 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_529_6
timestamp 1731220588
transform 1 0 536 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_528_6
timestamp 1731220588
transform 1 0 416 0 1 3148
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_527_6
timestamp 1731220588
transform 1 0 816 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_526_6
timestamp 1731220588
transform 1 0 656 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_525_6
timestamp 1731220588
transform 1 0 504 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_524_6
timestamp 1731220588
transform 1 0 368 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_523_6
timestamp 1731220588
transform 1 0 248 0 -1 3288
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_522_6
timestamp 1731220588
transform 1 0 680 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_521_6
timestamp 1731220588
transform 1 0 520 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_520_6
timestamp 1731220588
transform 1 0 352 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_519_6
timestamp 1731220588
transform 1 0 192 0 1 3292
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_518_6
timestamp 1731220588
transform 1 0 752 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_517_6
timestamp 1731220588
transform 1 0 576 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_516_6
timestamp 1731220588
transform 1 0 408 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_515_6
timestamp 1731220588
transform 1 0 248 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_514_6
timestamp 1731220588
transform 1 0 128 0 -1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_513_6
timestamp 1731220588
transform 1 0 168 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_512_6
timestamp 1731220588
transform 1 0 336 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_511_6
timestamp 1731220588
transform 1 0 504 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_510_6
timestamp 1731220588
transform 1 0 664 0 1 3436
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_59_6
timestamp 1731220588
transform 1 0 680 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_58_6
timestamp 1731220588
transform 1 0 536 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_57_6
timestamp 1731220588
transform 1 0 392 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_56_6
timestamp 1731220588
transform 1 0 240 0 -1 3572
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_55_6
timestamp 1731220588
transform 1 0 224 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_54_6
timestamp 1731220588
transform 1 0 312 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_53_6
timestamp 1731220588
transform 1 0 400 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_52_6
timestamp 1731220588
transform 1 0 488 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_51_6
timestamp 1731220588
transform 1 0 576 0 1 3580
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  tst_50_6
timestamp 1731220588
transform 1 0 664 0 1 3580
box 8 4 80 64
<< end >>
