magic
tech sky130l
timestamp 1730421333
<< ndiffusion >>
rect 8 23 13 24
rect 8 20 9 23
rect 12 20 13 23
rect 8 18 13 20
rect 15 22 20 24
rect 15 19 16 22
rect 19 19 20 22
rect 15 18 20 19
rect 22 23 27 24
rect 22 20 23 23
rect 26 20 27 23
rect 22 18 27 20
rect 29 23 44 24
rect 29 20 40 23
rect 43 20 44 23
rect 29 18 44 20
<< ndc >>
rect 9 20 12 23
rect 16 19 19 22
rect 23 20 26 23
rect 40 20 43 23
<< ntransistor >>
rect 13 18 15 24
rect 20 18 22 24
rect 27 18 29 24
<< pdiffusion >>
rect 8 39 13 46
rect 8 36 9 39
rect 12 36 13 39
rect 8 31 13 36
rect 15 31 20 46
rect 22 39 26 46
rect 22 37 27 39
rect 22 34 23 37
rect 26 34 27 37
rect 22 31 27 34
rect 29 37 34 39
rect 29 35 44 37
rect 29 32 40 35
rect 43 32 44 35
rect 29 31 44 32
<< pdc >>
rect 9 36 12 39
rect 23 34 26 37
rect 40 32 43 35
<< ptransistor >>
rect 13 31 15 46
rect 20 31 22 46
rect 27 31 29 39
<< polysilicon >>
rect 10 53 15 54
rect 10 50 11 53
rect 14 50 15 53
rect 10 49 15 50
rect 18 53 23 54
rect 18 50 19 53
rect 22 50 23 53
rect 18 49 23 50
rect 13 46 15 49
rect 20 46 22 49
rect 27 39 29 41
rect 13 24 15 31
rect 20 24 22 31
rect 27 24 29 31
rect 13 16 15 18
rect 20 16 22 18
rect 27 8 29 18
rect 25 7 30 8
rect 25 4 26 7
rect 29 4 30 7
rect 25 3 30 4
<< pc >>
rect 11 50 14 53
rect 19 50 22 53
rect 26 4 29 7
<< m1 >>
rect 10 53 15 54
rect 10 50 11 53
rect 14 50 15 53
rect 10 49 15 50
rect 18 53 22 54
rect 18 50 19 53
rect 18 49 22 50
rect 25 49 26 52
rect 25 48 29 49
rect 32 48 36 52
rect 25 44 28 48
rect 23 41 28 44
rect 9 39 12 40
rect 9 31 12 36
rect 23 37 26 41
rect 23 33 26 34
rect 8 23 13 24
rect 8 20 9 23
rect 12 20 13 23
rect 8 19 13 20
rect 16 22 19 28
rect 22 23 27 24
rect 22 20 23 23
rect 26 20 27 23
rect 22 19 27 20
rect 33 23 36 48
rect 33 19 36 20
rect 40 35 43 36
rect 40 23 43 32
rect 8 15 12 16
rect 11 12 12 15
rect 16 7 19 19
rect 40 15 43 20
rect 25 7 30 8
rect 25 4 26 7
rect 29 4 30 7
rect 25 3 30 4
<< m2c >>
rect 26 49 29 52
rect 9 28 12 31
rect 16 28 19 31
rect 9 20 12 23
rect 23 20 26 23
rect 33 20 36 23
rect 8 12 11 15
rect 40 12 43 15
rect 16 4 19 7
rect 26 4 29 7
<< m2 >>
rect 25 52 30 53
rect 25 49 26 52
rect 29 49 30 52
rect 25 48 30 49
rect 8 31 20 32
rect 8 28 9 31
rect 12 28 16 31
rect 19 28 20 31
rect 8 27 20 28
rect 8 23 13 24
rect 8 20 9 23
rect 12 22 13 23
rect 22 23 27 24
rect 22 22 23 23
rect 12 20 23 22
rect 26 22 27 23
rect 32 23 37 24
rect 32 22 33 23
rect 26 20 33 22
rect 36 20 37 23
rect 8 19 37 20
rect 7 15 12 16
rect 39 15 44 16
rect 7 12 8 15
rect 11 12 40 15
rect 43 12 44 15
rect 7 11 12 12
rect 39 11 44 12
rect 15 7 30 8
rect 15 4 16 7
rect 19 4 26 7
rect 29 4 30 7
rect 15 3 30 4
<< labels >>
rlabel space 0 0 48 56 6 prboundary
rlabel ndiffusion 44 21 44 21 3 Y
rlabel pdiffusion 44 33 44 33 3 Y
rlabel ndiffusion 30 19 30 19 3 Y
rlabel ndiffusion 30 21 30 21 3 Y
rlabel ndiffusion 30 24 30 24 3 Y
rlabel pdiffusion 30 32 30 32 3 Y
rlabel pdiffusion 30 33 30 33 3 Y
rlabel pdiffusion 30 36 30 36 3 Y
rlabel pdiffusion 30 38 30 38 3 Y
rlabel pdiffusion 27 35 27 35 3 Vdd
rlabel polysilicon 28 40 28 40 3 _Y
rlabel polysilicon 23 51 23 51 3 A
rlabel ntransistor 28 19 28 19 3 _Y
rlabel polysilicon 28 25 28 25 3 _Y
rlabel ptransistor 28 32 28 32 3 _Y
rlabel polysilicon 21 47 21 47 3 A
rlabel ndiffusion 23 19 23 19 3 GND
rlabel ndiffusion 20 20 20 20 3 _Y
rlabel pdiffusion 23 32 23 32 3 Vdd
rlabel pdiffusion 23 35 23 35 3 Vdd
rlabel pdiffusion 23 38 23 38 3 Vdd
rlabel pdiffusion 23 40 23 40 3 Vdd
rlabel polysilicon 28 9 28 9 3 _Y
rlabel polysilicon 21 17 21 17 3 A
rlabel ntransistor 21 19 21 19 3 A
rlabel polysilicon 21 25 21 25 3 A
rlabel ptransistor 21 32 21 32 3 A
rlabel ndiffusion 16 19 16 19 3 _Y
rlabel ndiffusion 16 20 16 20 3 _Y
rlabel ndiffusion 16 23 16 23 3 _Y
rlabel pdiffusion 13 37 13 37 3 _Y
rlabel polysilicon 14 47 14 47 3 B
rlabel polysilicon 14 17 14 17 3 B
rlabel ntransistor 14 19 14 19 3 B
rlabel polysilicon 14 25 14 25 3 B
rlabel ptransistor 14 32 14 32 3 B
rlabel ndiffusion 9 19 9 19 3 GND
rlabel pdiffusion 9 37 9 37 3 _Y
rlabel pdiffusion 9 40 9 40 3 _Y
rlabel ndc 41 21 41 21 3 Y
port 1 e
rlabel m1 41 24 41 24 3 Y
port 1 e
rlabel pdc 41 33 41 33 3 Y
port 1 e
rlabel m1 41 36 41 36 3 Y
port 1 e
rlabel m1 33 49 33 49 3 GND
rlabel m1 41 16 41 16 3 Y
port 1 e
rlabel m1 34 20 34 20 3 GND
rlabel m1 34 24 34 24 3 GND
rlabel m1 26 45 26 45 3 Vdd
rlabel m1 26 49 26 49 3 Vdd
rlabel m1 26 5 26 5 3 _Y
rlabel m1 26 8 26 8 3 _Y
rlabel m1 24 34 24 34 3 Vdd
rlabel pdc 24 35 24 35 3 Vdd
rlabel m1 24 38 24 38 3 Vdd
rlabel m1 24 42 24 42 3 Vdd
rlabel m1 26 4 26 4 3 _Y
rlabel m1 23 20 23 20 3 GND
rlabel m1 23 21 23 21 3 GND
rlabel m1 17 23 17 23 3 _Y
rlabel pc 20 51 20 51 3 A
port 2 e
rlabel m1 15 51 15 51 3 B
port 3 e
rlabel m1 17 8 17 8 3 _Y
rlabel m1 19 50 19 50 3 A
port 2 e
rlabel m1 19 51 19 51 3 A
port 2 e
rlabel m1 19 54 19 54 3 A
port 2 e
rlabel pc 12 51 12 51 3 B
port 3 e
rlabel ndc 17 20 17 20 3 _Y
rlabel m1 11 50 11 50 3 B
port 3 e
rlabel m1 11 51 11 51 3 B
port 3 e
rlabel m1 11 54 11 54 3 B
port 3 e
rlabel m1 10 32 10 32 3 _Y
rlabel pdc 10 37 10 37 3 _Y
rlabel m1 10 40 10 40 3 _Y
rlabel m1 9 16 9 16 3 Y
port 1 e
rlabel m2 30 5 30 5 3 _Y
rlabel m2 37 21 37 21 3 GND
rlabel m2 33 23 33 23 3 GND
rlabel m2c 27 5 27 5 3 _Y
rlabel m2c 34 21 34 21 3 GND
rlabel m2 20 5 20 5 3 _Y
rlabel m2 40 12 40 12 3 Y
port 1 e
rlabel m2 27 21 27 21 3 GND
rlabel m2 27 23 27 23 3 GND
rlabel m2 23 23 23 23 3 GND
rlabel m2 33 24 33 24 3 GND
rlabel m2 20 29 20 29 3 _Y
rlabel m2c 17 5 17 5 3 _Y
rlabel m2 44 13 44 13 3 Y
port 1 e
rlabel m2c 24 21 24 21 3 GND
rlabel m2c 17 29 17 29 3 _Y
rlabel m2 16 4 16 4 3 _Y
rlabel m2 16 5 16 5 3 _Y
rlabel m2 16 8 16 8 3 _Y
rlabel m2c 41 13 41 13 3 Y
port 1 e
rlabel m2 13 21 13 21 3 GND
rlabel m2 13 23 13 23 3 GND
rlabel m2 23 24 23 24 3 GND
rlabel m2 13 29 13 29 3 _Y
rlabel m2 12 13 12 13 3 Y
port 1 e
rlabel m2 40 16 40 16 3 Y
port 1 e
rlabel m2c 10 21 10 21 3 GND
rlabel m2c 10 29 10 29 3 _Y
rlabel m2c 9 13 9 13 3 Y
port 1 e
rlabel m2 9 20 9 20 3 GND
rlabel m2 9 21 9 21 3 GND
rlabel m2 9 24 9 24 3 GND
rlabel m2 9 28 9 28 3 _Y
rlabel m2 9 29 9 29 3 _Y
rlabel m2 9 32 9 32 3 _Y
rlabel m2 8 12 8 12 3 Y
port 1 e
rlabel m2 8 13 8 13 3 Y
port 1 e
rlabel m2 8 16 8 16 3 Y
port 1 e
<< end >>
