magic
tech sky130l
timestamp 1730814361
<< m1 >>
rect 2352 1203 2356 1303
rect 2352 1183 2356 1199
rect 2352 1123 2356 1179
rect 2352 1103 2356 1119
<< m2c >>
rect 1671 3293 1675 3297
rect 3191 3293 3195 3297
rect 1671 3275 1675 3279
rect 3191 3275 3195 3279
rect 3064 3271 3068 3275
rect 1671 3257 1675 3261
rect 3008 3259 3012 3263
rect 2160 3255 2164 3259
rect 2296 3255 2300 3259
rect 2432 3255 2436 3259
rect 2576 3255 2580 3259
rect 2720 3255 2724 3259
rect 2864 3255 2868 3259
rect 3191 3257 3195 3261
rect 1671 3239 1675 3243
rect 3191 3239 3195 3243
rect 1671 3213 1675 3217
rect 3191 3213 3195 3217
rect 1671 3195 1675 3199
rect 2552 3195 2556 3199
rect 2736 3195 2740 3199
rect 3191 3195 3195 3199
rect 2008 3191 2012 3195
rect 2184 3191 2188 3195
rect 2368 3191 2372 3195
rect 2928 3191 2932 3195
rect 3120 3191 3124 3195
rect 1671 3177 1675 3181
rect 2048 3179 2052 3183
rect 2704 3179 2708 3183
rect 3168 3179 3172 3183
rect 1856 3175 1860 3179
rect 2256 3175 2260 3179
rect 2472 3175 2476 3179
rect 2944 3175 2948 3179
rect 3191 3177 3195 3181
rect 1671 3159 1675 3163
rect 3191 3159 3195 3163
rect 1671 3133 1675 3137
rect 3191 3133 3195 3137
rect 111 3117 115 3121
rect 1608 3119 1612 3123
rect 816 3115 820 3119
rect 1088 3115 1092 3119
rect 1360 3115 1364 3119
rect 1631 3117 1635 3121
rect 1671 3115 1675 3119
rect 1704 3115 1708 3119
rect 1872 3115 1876 3119
rect 2032 3115 2036 3119
rect 2520 3115 2524 3119
rect 3191 3115 3195 3119
rect 2192 3111 2196 3115
rect 2352 3111 2356 3115
rect 111 3099 115 3103
rect 1631 3099 1635 3103
rect 1671 3097 1675 3101
rect 2192 3099 2196 3103
rect 2424 3099 2428 3103
rect 2664 3099 2668 3103
rect 1968 3095 1972 3099
rect 2912 3095 2916 3099
rect 3168 3095 3172 3099
rect 3191 3097 3195 3101
rect 1671 3079 1675 3083
rect 3191 3079 3195 3083
rect 111 3069 115 3073
rect 1631 3069 1635 3073
rect 111 3051 115 3055
rect 840 3051 844 3055
rect 1088 3051 1092 3055
rect 1432 3051 1436 3055
rect 1552 3051 1556 3055
rect 1631 3051 1635 3055
rect 1671 3053 1675 3057
rect 3191 3053 3195 3057
rect 712 3047 716 3051
rect 968 3047 972 3051
rect 1208 3047 1212 3051
rect 1320 3047 1324 3051
rect 1671 3035 1675 3039
rect 1880 3035 1884 3039
rect 2640 3035 2644 3039
rect 3168 3035 3172 3039
rect 3191 3035 3195 3039
rect 2120 3031 2124 3035
rect 2376 3031 2380 3035
rect 2912 3031 2916 3035
rect 111 3025 115 3029
rect 632 3027 636 3031
rect 792 3027 796 3031
rect 936 3027 940 3031
rect 1072 3027 1076 3031
rect 1200 3025 1204 3029
rect 1448 3027 1452 3031
rect 1320 3023 1324 3027
rect 1631 3025 1635 3029
rect 1671 3017 1675 3021
rect 2296 3019 2300 3023
rect 2632 3019 2636 3023
rect 1800 3015 1804 3019
rect 1968 3015 1972 3019
rect 2136 3015 2140 3019
rect 2464 3015 2468 3019
rect 3191 3017 3195 3021
rect 111 3007 115 3011
rect 1631 3007 1635 3011
rect 1671 2999 1675 3003
rect 3191 2999 3195 3003
rect 111 2977 115 2981
rect 1631 2977 1635 2981
rect 1671 2973 1675 2977
rect 3191 2973 3195 2977
rect 111 2959 115 2963
rect 792 2959 796 2963
rect 928 2959 932 2963
rect 1064 2959 1068 2963
rect 1200 2959 1204 2963
rect 1631 2959 1635 2963
rect 528 2955 532 2959
rect 656 2955 660 2959
rect 1344 2955 1348 2959
rect 1671 2955 1675 2959
rect 1712 2955 1716 2959
rect 1912 2955 1916 2959
rect 2376 2955 2380 2959
rect 2632 2955 2636 2959
rect 3168 2955 3172 2959
rect 3191 2955 3195 2959
rect 2136 2951 2140 2955
rect 2896 2951 2900 2955
rect 111 2933 115 2937
rect 608 2935 612 2939
rect 1448 2935 1452 2939
rect 1671 2937 1675 2941
rect 1704 2939 1708 2943
rect 2528 2939 2532 2943
rect 3144 2939 3148 2943
rect 448 2931 452 2935
rect 768 2931 772 2935
rect 936 2931 940 2935
rect 1104 2931 1108 2935
rect 1272 2931 1276 2935
rect 1608 2931 1612 2935
rect 1631 2933 1635 2937
rect 1944 2935 1948 2939
rect 2232 2935 2236 2939
rect 2832 2935 2836 2939
rect 3191 2937 3195 2941
rect 1671 2919 1675 2923
rect 3191 2919 3195 2923
rect 111 2915 115 2919
rect 1631 2915 1635 2919
rect 1671 2893 1675 2897
rect 3191 2893 3195 2897
rect 111 2889 115 2893
rect 1631 2889 1635 2893
rect 1671 2875 1675 2879
rect 2304 2875 2308 2879
rect 2560 2875 2564 2879
rect 3191 2875 3195 2879
rect 111 2871 115 2875
rect 1600 2871 1604 2875
rect 1631 2871 1635 2875
rect 2824 2871 2828 2875
rect 3088 2871 3092 2875
rect 344 2867 348 2871
rect 480 2867 484 2871
rect 632 2867 636 2871
rect 800 2867 804 2871
rect 984 2867 988 2871
rect 1184 2867 1188 2871
rect 1392 2867 1396 2871
rect 1671 2857 1675 2861
rect 2216 2859 2220 2863
rect 2544 2859 2548 2863
rect 3120 2859 3124 2863
rect 2384 2855 2388 2859
rect 2688 2855 2692 2859
rect 2832 2855 2836 2859
rect 2976 2855 2980 2859
rect 3191 2857 3195 2861
rect 111 2845 115 2849
rect 264 2843 268 2847
rect 424 2843 428 2847
rect 568 2843 572 2847
rect 704 2843 708 2847
rect 832 2843 836 2847
rect 960 2843 964 2847
rect 1096 2843 1100 2847
rect 1631 2845 1635 2849
rect 1671 2839 1675 2843
rect 3191 2839 3195 2843
rect 111 2827 115 2831
rect 1631 2827 1635 2831
rect 1671 2805 1675 2809
rect 3191 2805 3195 2809
rect 111 2793 115 2797
rect 1631 2793 1635 2797
rect 1671 2787 1675 2791
rect 2312 2787 2316 2791
rect 2488 2787 2492 2791
rect 3191 2787 3195 2791
rect 2136 2783 2140 2787
rect 2664 2783 2668 2787
rect 2840 2783 2844 2787
rect 3016 2783 3020 2787
rect 3168 2783 3172 2787
rect 111 2775 115 2779
rect 408 2775 412 2779
rect 528 2775 532 2779
rect 648 2775 652 2779
rect 760 2775 764 2779
rect 872 2775 876 2779
rect 992 2775 996 2779
rect 1631 2775 1635 2779
rect 160 2771 164 2775
rect 288 2771 292 2775
rect 1671 2769 1675 2773
rect 2384 2771 2388 2775
rect 2544 2771 2548 2775
rect 2048 2767 2052 2771
rect 2216 2767 2220 2771
rect 2712 2767 2716 2771
rect 2880 2767 2884 2771
rect 3191 2769 3195 2773
rect 1671 2751 1675 2755
rect 3191 2751 3195 2755
rect 111 2745 115 2749
rect 144 2747 148 2751
rect 632 2747 636 2751
rect 848 2747 852 2751
rect 1576 2747 1580 2751
rect 272 2743 276 2747
rect 440 2743 444 2747
rect 1080 2743 1084 2747
rect 1328 2743 1332 2747
rect 1631 2745 1635 2749
rect 111 2727 115 2731
rect 1631 2727 1635 2731
rect 1671 2721 1675 2725
rect 3191 2721 3195 2725
rect 1671 2703 1675 2707
rect 2584 2703 2588 2707
rect 2784 2703 2788 2707
rect 3191 2703 3195 2707
rect 2024 2699 2028 2703
rect 2208 2699 2212 2703
rect 2392 2699 2396 2703
rect 2984 2699 2988 2703
rect 3168 2699 3172 2703
rect 111 2689 115 2693
rect 1631 2689 1635 2693
rect 1671 2677 1675 2681
rect 2368 2679 2372 2683
rect 2560 2679 2564 2683
rect 2768 2679 2772 2683
rect 2008 2675 2012 2679
rect 2184 2675 2188 2679
rect 2976 2677 2980 2681
rect 3168 2675 3172 2679
rect 3191 2677 3195 2681
rect 111 2671 115 2675
rect 712 2671 716 2675
rect 968 2671 972 2675
rect 1320 2671 1324 2675
rect 1432 2671 1436 2675
rect 1552 2671 1556 2675
rect 1631 2671 1635 2675
rect 840 2667 844 2671
rect 1088 2667 1092 2671
rect 1208 2667 1212 2671
rect 1671 2659 1675 2663
rect 3191 2659 3195 2663
rect 111 2645 115 2649
rect 616 2647 620 2651
rect 744 2647 748 2651
rect 1328 2647 1332 2651
rect 1448 2647 1452 2651
rect 864 2643 868 2647
rect 984 2643 988 2647
rect 1104 2643 1108 2647
rect 1216 2643 1220 2647
rect 1631 2645 1635 2649
rect 1671 2633 1675 2637
rect 3191 2633 3195 2637
rect 111 2627 115 2631
rect 1631 2627 1635 2631
rect 1671 2615 1675 2619
rect 2304 2615 2308 2619
rect 2696 2615 2700 2619
rect 3191 2615 3195 2619
rect 1920 2611 1924 2615
rect 2112 2611 2116 2615
rect 2496 2611 2500 2615
rect 1671 2597 1675 2601
rect 2448 2599 2452 2603
rect 2680 2599 2684 2603
rect 1832 2595 1836 2599
rect 2024 2595 2028 2599
rect 2224 2595 2228 2599
rect 2928 2595 2932 2599
rect 3168 2595 3172 2599
rect 3191 2597 3195 2601
rect 111 2589 115 2593
rect 1631 2589 1635 2593
rect 1671 2579 1675 2583
rect 3191 2579 3195 2583
rect 111 2571 115 2575
rect 880 2571 884 2575
rect 1000 2571 1004 2575
rect 1224 2571 1228 2575
rect 1344 2571 1348 2575
rect 1631 2571 1635 2575
rect 512 2567 516 2571
rect 640 2567 644 2571
rect 760 2567 764 2571
rect 1112 2567 1116 2571
rect 1671 2549 1675 2553
rect 3191 2549 3195 2553
rect 111 2541 115 2545
rect 784 2543 788 2547
rect 904 2543 908 2547
rect 1016 2543 1020 2547
rect 1248 2543 1252 2547
rect 408 2539 412 2543
rect 536 2539 540 2543
rect 664 2539 668 2543
rect 1128 2539 1132 2543
rect 1631 2541 1635 2545
rect 1671 2531 1675 2535
rect 2064 2531 2068 2535
rect 2224 2531 2228 2535
rect 3191 2531 3195 2535
rect 1744 2527 1748 2531
rect 1904 2527 1908 2531
rect 2384 2527 2388 2531
rect 2544 2527 2548 2531
rect 111 2523 115 2527
rect 1631 2523 1635 2527
rect 1671 2509 1675 2513
rect 1704 2511 1708 2515
rect 2328 2511 2332 2515
rect 2592 2511 2596 2515
rect 1872 2507 1876 2511
rect 2088 2507 2092 2511
rect 2864 2507 2868 2511
rect 3144 2507 3148 2511
rect 3191 2509 3195 2513
rect 1671 2491 1675 2495
rect 3191 2491 3195 2495
rect 111 2485 115 2489
rect 1631 2485 1635 2489
rect 111 2467 115 2471
rect 872 2467 876 2471
rect 1048 2467 1052 2471
rect 1432 2467 1436 2471
rect 1608 2467 1612 2471
rect 1631 2467 1635 2471
rect 312 2463 316 2467
rect 440 2463 444 2467
rect 568 2463 572 2467
rect 712 2463 716 2467
rect 1232 2463 1236 2467
rect 1671 2457 1675 2461
rect 3191 2457 3195 2461
rect 111 2445 115 2449
rect 960 2447 964 2451
rect 1168 2447 1172 2451
rect 1384 2447 1388 2451
rect 1600 2449 1604 2453
rect 208 2443 212 2447
rect 336 2443 340 2447
rect 464 2443 468 2447
rect 608 2443 612 2447
rect 776 2443 780 2447
rect 1631 2445 1635 2449
rect 1671 2439 1675 2443
rect 2328 2439 2332 2443
rect 2576 2439 2580 2443
rect 2832 2439 2836 2443
rect 3191 2439 3195 2443
rect 3088 2435 3092 2439
rect 111 2427 115 2431
rect 1631 2427 1635 2431
rect 1671 2421 1675 2425
rect 2240 2423 2244 2427
rect 2552 2423 2556 2427
rect 2832 2423 2836 2427
rect 2400 2419 2404 2423
rect 2696 2419 2700 2423
rect 2976 2419 2980 2423
rect 3120 2419 3124 2423
rect 3191 2421 3195 2425
rect 1671 2403 1675 2407
rect 3191 2403 3195 2407
rect 111 2385 115 2389
rect 1631 2385 1635 2389
rect 111 2367 115 2371
rect 144 2363 148 2367
rect 248 2363 252 2367
rect 368 2363 372 2367
rect 488 2363 492 2367
rect 600 2365 604 2369
rect 1631 2367 1635 2371
rect 1671 2369 1675 2373
rect 3191 2369 3195 2373
rect 712 2363 716 2367
rect 824 2363 828 2367
rect 944 2363 948 2367
rect 1671 2351 1675 2355
rect 2320 2351 2324 2355
rect 2664 2351 2668 2355
rect 3016 2351 3020 2355
rect 3191 2351 3195 2355
rect 2152 2347 2156 2351
rect 2488 2347 2492 2351
rect 2840 2347 2844 2351
rect 3168 2347 3172 2351
rect 111 2341 115 2345
rect 984 2343 988 2347
rect 1376 2343 1380 2347
rect 1576 2343 1580 2347
rect 144 2339 148 2343
rect 352 2339 356 2343
rect 576 2339 580 2343
rect 784 2339 788 2343
rect 1184 2339 1188 2343
rect 1631 2341 1635 2345
rect 1671 2333 1675 2337
rect 2344 2335 2348 2339
rect 2632 2335 2636 2339
rect 2776 2335 2780 2339
rect 2928 2335 2932 2339
rect 2192 2331 2196 2335
rect 2488 2331 2492 2335
rect 3191 2333 3195 2337
rect 111 2323 115 2327
rect 1631 2323 1635 2327
rect 1671 2315 1675 2319
rect 3191 2315 3195 2319
rect 111 2285 115 2289
rect 1631 2285 1635 2289
rect 1671 2285 1675 2289
rect 3191 2285 3195 2289
rect 111 2267 115 2271
rect 912 2267 916 2271
rect 1032 2267 1036 2271
rect 1152 2267 1156 2271
rect 1264 2267 1268 2271
rect 1496 2267 1500 2271
rect 1631 2267 1635 2271
rect 1671 2267 1675 2271
rect 2104 2269 2108 2273
rect 2800 2267 2804 2271
rect 2992 2267 2996 2271
rect 3191 2267 3195 2271
rect 664 2263 668 2267
rect 792 2263 796 2267
rect 1376 2263 1380 2267
rect 2272 2263 2276 2267
rect 2440 2263 2444 2267
rect 2616 2263 2620 2267
rect 3168 2263 3172 2267
rect 1671 2249 1675 2253
rect 2472 2251 2476 2255
rect 2616 2251 2620 2255
rect 2768 2251 2772 2255
rect 2024 2247 2028 2251
rect 2176 2247 2180 2251
rect 2328 2247 2332 2251
rect 3191 2249 3195 2253
rect 111 2237 115 2241
rect 816 2239 820 2243
rect 1056 2241 1060 2245
rect 1168 2241 1172 2245
rect 1280 2239 1284 2243
rect 1400 2239 1404 2243
rect 560 2235 564 2239
rect 688 2235 692 2239
rect 936 2235 940 2239
rect 1631 2237 1635 2241
rect 1671 2231 1675 2235
rect 3191 2231 3195 2235
rect 111 2219 115 2223
rect 1631 2219 1635 2223
rect 1671 2201 1675 2205
rect 3191 2201 3195 2205
rect 111 2185 115 2189
rect 1631 2185 1635 2189
rect 1671 2183 1675 2187
rect 2112 2185 2116 2189
rect 2728 2183 2732 2187
rect 2960 2183 2964 2187
rect 3191 2183 3195 2187
rect 1936 2179 1940 2183
rect 2304 2179 2308 2183
rect 2512 2179 2516 2183
rect 3168 2179 3172 2183
rect 111 2167 115 2171
rect 1064 2167 1068 2171
rect 1176 2167 1180 2171
rect 1296 2167 1300 2171
rect 1631 2167 1635 2171
rect 464 2163 468 2167
rect 592 2163 596 2167
rect 712 2163 716 2167
rect 832 2163 836 2167
rect 952 2163 956 2167
rect 1671 2165 1675 2169
rect 1856 2167 1860 2171
rect 2008 2167 2012 2171
rect 2160 2167 2164 2171
rect 2456 2167 2460 2171
rect 2608 2167 2612 2171
rect 2304 2163 2308 2167
rect 3191 2165 3195 2169
rect 1671 2147 1675 2151
rect 3191 2147 3195 2151
rect 111 2137 115 2141
rect 360 2135 364 2139
rect 488 2135 492 2139
rect 608 2135 612 2139
rect 728 2135 732 2139
rect 848 2135 852 2139
rect 960 2135 964 2139
rect 1072 2135 1076 2139
rect 1192 2135 1196 2139
rect 1631 2137 1635 2141
rect 111 2119 115 2123
rect 1631 2119 1635 2123
rect 1671 2117 1675 2121
rect 3191 2117 3195 2121
rect 1671 2099 1675 2103
rect 2080 2099 2084 2103
rect 2472 2099 2476 2103
rect 2696 2099 2700 2103
rect 2936 2099 2940 2103
rect 3191 2099 3195 2103
rect 1768 2095 1772 2099
rect 1920 2095 1924 2099
rect 2264 2095 2268 2099
rect 3168 2095 3172 2099
rect 111 2081 115 2085
rect 1631 2081 1635 2085
rect 1671 2081 1675 2085
rect 1832 2083 1836 2087
rect 1976 2083 1980 2087
rect 2120 2083 2124 2087
rect 2416 2083 2420 2087
rect 1704 2079 1708 2083
rect 2264 2079 2268 2083
rect 3191 2081 3195 2085
rect 111 2063 115 2067
rect 632 2063 636 2067
rect 1096 2063 1100 2067
rect 1631 2063 1635 2067
rect 1671 2063 1675 2067
rect 3191 2063 3195 2067
rect 256 2059 260 2063
rect 384 2059 388 2063
rect 512 2059 516 2063
rect 752 2059 756 2063
rect 864 2059 868 2063
rect 976 2059 980 2063
rect 111 2037 115 2041
rect 1192 2039 1196 2043
rect 184 2035 188 2039
rect 376 2035 380 2039
rect 568 2035 572 2039
rect 768 2035 772 2039
rect 976 2035 980 2039
rect 1408 2035 1412 2039
rect 1608 2035 1612 2039
rect 1631 2037 1635 2041
rect 1671 2037 1675 2041
rect 3191 2037 3195 2041
rect 111 2019 115 2023
rect 1631 2019 1635 2023
rect 1671 2019 1675 2023
rect 1704 2019 1708 2023
rect 2048 2019 2052 2023
rect 2416 2019 2420 2023
rect 2776 2019 2780 2023
rect 3191 2019 3195 2023
rect 3144 2015 3148 2019
rect 111 1993 115 1997
rect 1631 1993 1635 1997
rect 1671 1993 1675 1997
rect 2424 1995 2428 1999
rect 2712 1995 2716 1999
rect 2848 1995 2852 1999
rect 2272 1991 2276 1995
rect 2568 1991 2572 1995
rect 2984 1991 2988 1995
rect 3120 1991 3124 1995
rect 3191 1993 3195 1997
rect 111 1975 115 1979
rect 240 1975 244 1979
rect 360 1975 364 1979
rect 472 1975 476 1979
rect 584 1975 588 1979
rect 1631 1975 1635 1979
rect 1671 1975 1675 1979
rect 3191 1975 3195 1979
rect 144 1971 148 1975
rect 696 1971 700 1975
rect 808 1971 812 1975
rect 920 1971 924 1975
rect 111 1949 115 1953
rect 864 1951 868 1955
rect 1576 1951 1580 1955
rect 736 1947 740 1951
rect 992 1947 996 1951
rect 1112 1947 1116 1951
rect 1232 1947 1236 1951
rect 1344 1947 1348 1951
rect 1456 1947 1460 1951
rect 1631 1949 1635 1953
rect 1671 1949 1675 1953
rect 3191 1949 3195 1953
rect 111 1931 115 1935
rect 1631 1931 1635 1935
rect 1671 1931 1675 1935
rect 2400 1931 2404 1935
rect 2552 1931 2556 1935
rect 2704 1931 2708 1935
rect 2856 1931 2860 1935
rect 3008 1931 3012 1935
rect 3191 1931 3195 1935
rect 2248 1927 2252 1931
rect 1671 1909 1675 1913
rect 2648 1911 2652 1915
rect 2824 1911 2828 1915
rect 3008 1911 3012 1915
rect 3168 1911 3172 1915
rect 2160 1907 2164 1911
rect 2320 1907 2324 1911
rect 2480 1907 2484 1911
rect 3191 1909 3195 1913
rect 111 1893 115 1897
rect 1631 1893 1635 1897
rect 1671 1891 1675 1895
rect 3191 1891 3195 1895
rect 111 1875 115 1879
rect 888 1875 892 1879
rect 1008 1875 1012 1879
rect 1128 1875 1132 1879
rect 1240 1875 1244 1879
rect 1352 1875 1356 1879
rect 1472 1875 1476 1879
rect 1631 1875 1635 1879
rect 640 1871 644 1875
rect 768 1871 772 1875
rect 1671 1861 1675 1865
rect 3191 1861 3195 1865
rect 111 1845 115 1849
rect 536 1847 540 1851
rect 1136 1847 1140 1851
rect 1256 1847 1260 1851
rect 664 1843 668 1847
rect 784 1843 788 1847
rect 904 1843 908 1847
rect 1024 1843 1028 1847
rect 1376 1843 1380 1847
rect 1631 1845 1635 1849
rect 1671 1843 1675 1847
rect 2248 1843 2252 1847
rect 2424 1843 2428 1847
rect 2608 1843 2612 1847
rect 2800 1843 2804 1847
rect 2992 1843 2996 1847
rect 3168 1843 3172 1847
rect 3191 1843 3195 1847
rect 2080 1839 2084 1843
rect 111 1827 115 1831
rect 1631 1827 1635 1831
rect 1671 1825 1675 1829
rect 2592 1827 2596 1831
rect 2744 1827 2748 1831
rect 1992 1823 1996 1827
rect 2144 1823 2148 1827
rect 2296 1823 2300 1827
rect 2440 1823 2444 1827
rect 3191 1825 3195 1829
rect 1671 1807 1675 1811
rect 3191 1807 3195 1811
rect 111 1793 115 1797
rect 1631 1793 1635 1797
rect 1671 1781 1675 1785
rect 3191 1781 3195 1785
rect 111 1775 115 1779
rect 688 1775 692 1779
rect 808 1775 812 1779
rect 928 1775 932 1779
rect 1040 1775 1044 1779
rect 1152 1775 1156 1779
rect 1272 1775 1276 1779
rect 1631 1775 1635 1779
rect 432 1771 436 1775
rect 560 1771 564 1775
rect 1671 1763 1675 1767
rect 1912 1763 1916 1767
rect 2088 1763 2092 1767
rect 2280 1763 2284 1767
rect 2496 1763 2500 1767
rect 2720 1763 2724 1767
rect 2952 1763 2956 1767
rect 3168 1763 3172 1767
rect 3191 1763 3195 1767
rect 111 1745 115 1749
rect 336 1743 340 1747
rect 464 1743 468 1747
rect 584 1743 588 1747
rect 704 1743 708 1747
rect 824 1745 828 1749
rect 936 1743 940 1747
rect 1048 1743 1052 1747
rect 1168 1743 1172 1747
rect 1631 1745 1635 1749
rect 1671 1737 1675 1741
rect 3168 1739 3172 1743
rect 1824 1735 1828 1739
rect 1976 1735 1980 1739
rect 2136 1735 2140 1739
rect 2312 1735 2316 1739
rect 2512 1735 2516 1739
rect 2720 1735 2724 1739
rect 2944 1735 2948 1739
rect 3191 1737 3195 1741
rect 111 1727 115 1731
rect 1631 1727 1635 1731
rect 1671 1719 1675 1723
rect 3191 1719 3195 1723
rect 1671 1693 1675 1697
rect 3191 1693 3195 1697
rect 111 1689 115 1693
rect 1631 1689 1635 1693
rect 1671 1675 1675 1679
rect 1888 1675 1892 1679
rect 2032 1675 2036 1679
rect 2320 1675 2324 1679
rect 2472 1675 2476 1679
rect 3191 1675 3195 1679
rect 111 1671 115 1675
rect 720 1671 724 1675
rect 832 1671 836 1675
rect 952 1671 956 1675
rect 1631 1671 1635 1675
rect 1744 1671 1748 1675
rect 2176 1671 2180 1675
rect 232 1667 236 1671
rect 360 1667 364 1671
rect 480 1667 484 1671
rect 600 1667 604 1671
rect 1072 1667 1076 1671
rect 1671 1657 1675 1661
rect 1704 1659 1708 1663
rect 1904 1659 1908 1663
rect 3144 1659 3148 1663
rect 2136 1655 2140 1659
rect 2376 1655 2380 1659
rect 2624 1655 2628 1659
rect 2880 1655 2884 1659
rect 3191 1657 3195 1661
rect 111 1641 115 1645
rect 392 1643 396 1647
rect 720 1643 724 1647
rect 928 1643 932 1647
rect 1152 1643 1156 1647
rect 1608 1643 1612 1647
rect 144 1639 148 1643
rect 256 1639 260 1643
rect 544 1639 548 1643
rect 1392 1639 1396 1643
rect 1631 1641 1635 1645
rect 1671 1639 1675 1643
rect 3191 1639 3195 1643
rect 111 1623 115 1627
rect 1631 1623 1635 1627
rect 1671 1609 1675 1613
rect 3191 1609 3195 1613
rect 111 1589 115 1593
rect 1631 1589 1635 1593
rect 1671 1591 1675 1595
rect 3120 1591 3124 1595
rect 3191 1591 3195 1595
rect 2328 1587 2332 1591
rect 2528 1587 2532 1591
rect 2720 1587 2724 1591
rect 2920 1587 2924 1591
rect 111 1571 115 1575
rect 144 1571 148 1575
rect 312 1571 316 1575
rect 512 1571 516 1575
rect 704 1571 708 1575
rect 1072 1571 1076 1575
rect 1248 1571 1252 1575
rect 1631 1571 1635 1575
rect 1671 1573 1675 1577
rect 2280 1575 2284 1579
rect 2424 1571 2428 1575
rect 2568 1571 2572 1575
rect 2704 1571 2708 1575
rect 2848 1571 2852 1575
rect 2992 1571 2996 1575
rect 3191 1573 3195 1577
rect 896 1567 900 1571
rect 1424 1567 1428 1571
rect 1600 1567 1604 1571
rect 1671 1555 1675 1559
rect 3191 1555 3195 1559
rect 111 1541 115 1545
rect 688 1543 692 1547
rect 1056 1543 1060 1547
rect 1176 1543 1180 1547
rect 1288 1543 1292 1547
rect 816 1539 820 1543
rect 936 1539 940 1543
rect 1408 1539 1412 1543
rect 1528 1539 1532 1543
rect 1631 1541 1635 1545
rect 111 1523 115 1527
rect 1631 1523 1635 1527
rect 1671 1521 1675 1525
rect 3191 1521 3195 1525
rect 1671 1503 1675 1507
rect 2288 1503 2292 1507
rect 2400 1503 2404 1507
rect 2624 1503 2628 1507
rect 2744 1503 2748 1507
rect 2864 1503 2868 1507
rect 3120 1503 3124 1507
rect 3191 1503 3195 1507
rect 2176 1499 2180 1503
rect 2512 1499 2516 1503
rect 2992 1499 2996 1503
rect 111 1489 115 1493
rect 1631 1489 1635 1493
rect 1671 1481 1675 1485
rect 2240 1483 2244 1487
rect 2384 1483 2388 1487
rect 2520 1483 2524 1487
rect 2664 1483 2668 1487
rect 2808 1483 2812 1487
rect 2096 1479 2100 1483
rect 3191 1481 3195 1485
rect 111 1471 115 1475
rect 1304 1471 1308 1475
rect 1424 1471 1428 1475
rect 1631 1471 1635 1475
rect 584 1467 588 1471
rect 712 1467 716 1471
rect 840 1467 844 1471
rect 960 1467 964 1471
rect 1080 1467 1084 1471
rect 1192 1467 1196 1471
rect 1671 1463 1675 1467
rect 3191 1463 3195 1467
rect 111 1441 115 1445
rect 976 1443 980 1447
rect 1200 1443 1204 1447
rect 1320 1443 1324 1447
rect 488 1439 492 1443
rect 616 1439 620 1443
rect 736 1439 740 1443
rect 856 1439 860 1443
rect 1088 1439 1092 1443
rect 1631 1441 1635 1445
rect 1671 1433 1675 1437
rect 3191 1433 3195 1437
rect 111 1423 115 1427
rect 1631 1423 1635 1427
rect 1671 1415 1675 1419
rect 2104 1417 2108 1421
rect 2216 1415 2220 1419
rect 2344 1415 2348 1419
rect 2488 1415 2492 1419
rect 2648 1415 2652 1419
rect 3008 1415 3012 1419
rect 3168 1415 3172 1419
rect 3191 1415 3195 1419
rect 1992 1411 1996 1415
rect 2824 1411 2828 1415
rect 111 1385 115 1389
rect 1631 1385 1635 1389
rect 1671 1381 1675 1385
rect 2248 1383 2252 1387
rect 2400 1383 2404 1387
rect 2576 1383 2580 1387
rect 2776 1383 2780 1387
rect 2984 1383 2988 1387
rect 3168 1383 3172 1387
rect 1888 1379 1892 1383
rect 2000 1379 2004 1383
rect 2112 1379 2116 1383
rect 3191 1381 3195 1385
rect 111 1367 115 1371
rect 1224 1367 1228 1371
rect 1631 1367 1635 1371
rect 384 1363 388 1367
rect 512 1363 516 1367
rect 632 1363 636 1367
rect 752 1363 756 1367
rect 872 1363 876 1367
rect 984 1363 988 1367
rect 1104 1363 1108 1367
rect 1671 1363 1675 1367
rect 3191 1363 3195 1367
rect 111 1341 115 1345
rect 280 1339 284 1343
rect 408 1339 412 1343
rect 536 1339 540 1343
rect 656 1339 660 1343
rect 776 1339 780 1343
rect 888 1339 892 1343
rect 1000 1339 1004 1343
rect 1120 1339 1124 1343
rect 1631 1341 1635 1345
rect 111 1323 115 1327
rect 1631 1323 1635 1327
rect 1671 1325 1675 1329
rect 3191 1325 3195 1329
rect 1671 1307 1675 1311
rect 1896 1307 1900 1311
rect 2000 1307 2004 1311
rect 2104 1309 2108 1313
rect 2416 1307 2420 1311
rect 2520 1307 2524 1311
rect 3191 1307 3195 1311
rect 1784 1303 1788 1307
rect 2208 1303 2212 1307
rect 2312 1303 2316 1307
rect 2352 1303 2356 1307
rect 111 1285 115 1289
rect 1631 1285 1635 1289
rect 1671 1281 1675 1285
rect 1944 1283 1948 1287
rect 2112 1283 2116 1287
rect 2304 1285 2308 1289
rect 1704 1279 1708 1283
rect 1800 1279 1804 1283
rect 111 1267 115 1271
rect 312 1267 316 1271
rect 552 1267 556 1271
rect 1631 1267 1635 1271
rect 184 1263 188 1267
rect 432 1263 436 1267
rect 672 1263 676 1267
rect 784 1263 788 1267
rect 896 1263 900 1267
rect 1016 1263 1020 1267
rect 1671 1263 1675 1267
rect 111 1237 115 1241
rect 512 1239 516 1243
rect 144 1235 148 1239
rect 240 1235 244 1239
rect 368 1235 372 1239
rect 672 1235 676 1239
rect 840 1235 844 1239
rect 1024 1235 1028 1239
rect 1216 1235 1220 1239
rect 1416 1235 1420 1239
rect 1608 1235 1612 1239
rect 1631 1237 1635 1241
rect 111 1219 115 1223
rect 1631 1219 1635 1223
rect 1671 1221 1675 1225
rect 1671 1203 1675 1207
rect 1704 1203 1708 1207
rect 1992 1203 1996 1207
rect 2504 1283 2508 1287
rect 2944 1283 2948 1287
rect 3168 1283 3172 1287
rect 2720 1279 2724 1283
rect 3191 1281 3195 1285
rect 3191 1263 3195 1267
rect 3191 1221 3195 1225
rect 3144 1203 3148 1207
rect 3191 1203 3195 1207
rect 2264 1199 2268 1203
rect 2352 1199 2356 1203
rect 2504 1199 2508 1203
rect 2720 1199 2724 1203
rect 2928 1199 2932 1203
rect 111 1185 115 1189
rect 1631 1185 1635 1189
rect 1671 1181 1675 1185
rect 2256 1183 2260 1187
rect 2704 1183 2708 1187
rect 2856 1183 2860 1187
rect 2352 1179 2356 1183
rect 2408 1179 2412 1183
rect 2560 1179 2564 1183
rect 3008 1179 3012 1183
rect 3191 1181 3195 1185
rect 111 1167 115 1171
rect 1232 1167 1236 1171
rect 1576 1167 1580 1171
rect 1631 1167 1635 1171
rect 736 1163 740 1167
rect 864 1163 868 1167
rect 992 1163 996 1167
rect 1112 1163 1116 1167
rect 1344 1163 1348 1167
rect 1456 1163 1460 1167
rect 1671 1163 1675 1167
rect 111 1137 115 1141
rect 640 1135 644 1139
rect 768 1135 772 1139
rect 888 1135 892 1139
rect 1008 1135 1012 1139
rect 1128 1135 1132 1139
rect 1240 1135 1244 1139
rect 1352 1135 1356 1139
rect 1472 1135 1476 1139
rect 1631 1137 1635 1141
rect 1671 1137 1675 1141
rect 3191 1163 3195 1167
rect 3191 1137 3195 1141
rect 111 1119 115 1123
rect 1631 1119 1635 1123
rect 1671 1119 1675 1123
rect 2344 1119 2348 1123
rect 2352 1119 2356 1123
rect 2504 1119 2508 1123
rect 2664 1119 2668 1123
rect 2824 1119 2828 1123
rect 2984 1119 2988 1123
rect 3144 1119 3148 1123
rect 3191 1119 3195 1123
rect 2184 1115 2188 1119
rect 1671 1097 1675 1101
rect 2336 1099 2340 1103
rect 2352 1099 2356 1103
rect 2488 1099 2492 1103
rect 2648 1099 2652 1103
rect 2824 1099 2828 1103
rect 2080 1095 2084 1099
rect 2200 1095 2204 1099
rect 3008 1095 3012 1099
rect 3168 1095 3172 1099
rect 3191 1097 3195 1101
rect 111 1081 115 1085
rect 1631 1081 1635 1085
rect 1671 1079 1675 1083
rect 3191 1079 3195 1083
rect 111 1063 115 1067
rect 784 1063 788 1067
rect 1376 1063 1380 1067
rect 1631 1063 1635 1067
rect 536 1059 540 1063
rect 664 1059 668 1063
rect 904 1059 908 1063
rect 1024 1059 1028 1063
rect 1136 1059 1140 1063
rect 1256 1059 1260 1063
rect 111 1037 115 1041
rect 688 1039 692 1043
rect 1671 1041 1675 1045
rect 3191 1041 3195 1045
rect 432 1035 436 1039
rect 560 1035 564 1039
rect 808 1035 812 1039
rect 928 1035 932 1039
rect 1040 1035 1044 1039
rect 1152 1035 1156 1039
rect 1272 1035 1276 1039
rect 1631 1037 1635 1041
rect 1671 1023 1675 1027
rect 2352 1023 2356 1027
rect 2832 1023 2836 1027
rect 3008 1023 3012 1027
rect 3168 1023 3172 1027
rect 3191 1023 3195 1027
rect 111 1019 115 1023
rect 1631 1019 1635 1023
rect 1984 1019 1988 1023
rect 2104 1019 2108 1023
rect 2224 1019 2228 1023
rect 2496 1019 2500 1023
rect 2656 1019 2660 1023
rect 1671 1001 1675 1005
rect 2056 1003 2060 1007
rect 2208 1003 2212 1007
rect 2352 1003 2356 1007
rect 1904 999 1908 1003
rect 2504 999 2508 1003
rect 2656 999 2660 1003
rect 3191 1001 3195 1005
rect 111 981 115 985
rect 1631 981 1635 985
rect 1671 983 1675 987
rect 3191 983 3195 987
rect 111 963 115 967
rect 584 963 588 967
rect 704 963 708 967
rect 1631 963 1635 967
rect 336 959 340 963
rect 464 959 468 963
rect 824 959 828 963
rect 936 959 940 963
rect 1048 959 1052 963
rect 1168 959 1172 963
rect 1671 957 1675 961
rect 3191 957 3195 961
rect 1671 939 1675 943
rect 2264 939 2268 943
rect 2704 939 2708 943
rect 2944 939 2948 943
rect 3168 939 3172 943
rect 3191 939 3195 943
rect 111 933 115 937
rect 232 935 236 939
rect 360 931 364 935
rect 480 931 484 935
rect 600 931 604 935
rect 720 931 724 935
rect 832 931 836 935
rect 952 931 956 935
rect 1072 931 1076 935
rect 1631 933 1635 937
rect 1800 935 1804 939
rect 1928 935 1932 939
rect 2080 935 2084 939
rect 2472 935 2476 939
rect 111 915 115 919
rect 1631 915 1635 919
rect 1671 913 1675 917
rect 2232 915 2236 919
rect 2448 915 2452 919
rect 2680 915 2684 919
rect 2920 915 2924 919
rect 3168 915 3172 919
rect 1728 911 1732 915
rect 1880 911 1884 915
rect 2048 911 2052 915
rect 3191 913 3195 917
rect 1671 895 1675 899
rect 3191 895 3195 899
rect 111 877 115 881
rect 1631 877 1635 881
rect 1671 869 1675 873
rect 3191 869 3195 873
rect 111 859 115 863
rect 256 859 260 863
rect 1631 859 1635 863
rect 144 855 148 859
rect 392 855 396 859
rect 544 855 548 859
rect 720 855 724 859
rect 928 855 932 859
rect 1152 855 1156 859
rect 1392 855 1396 859
rect 1608 855 1612 859
rect 1671 851 1675 855
rect 1704 851 1708 855
rect 2024 851 2028 855
rect 2376 851 2380 855
rect 3096 851 3100 855
rect 3191 851 3195 855
rect 2736 847 2740 851
rect 111 837 115 841
rect 144 839 148 843
rect 312 839 316 843
rect 512 839 516 843
rect 1608 839 1612 843
rect 704 835 708 839
rect 888 835 892 839
rect 1056 835 1060 839
rect 1208 835 1212 839
rect 1344 835 1348 839
rect 1480 835 1484 839
rect 1631 837 1635 841
rect 111 819 115 823
rect 1631 819 1635 823
rect 1671 821 1675 825
rect 2448 823 2452 827
rect 2288 819 2292 823
rect 2592 819 2596 823
rect 2728 821 2732 825
rect 3120 823 3124 827
rect 2856 819 2860 823
rect 2984 819 2988 823
rect 3191 821 3195 825
rect 1671 803 1675 807
rect 3191 803 3195 807
rect 111 777 115 781
rect 1631 777 1635 781
rect 1671 773 1675 777
rect 3191 773 3195 777
rect 111 759 115 763
rect 1408 759 1412 763
rect 1528 759 1532 763
rect 1631 759 1635 763
rect 688 755 692 759
rect 816 755 820 759
rect 936 755 940 759
rect 1056 755 1060 759
rect 1176 755 1180 759
rect 1288 755 1292 759
rect 1671 755 1675 759
rect 2368 755 2372 759
rect 2520 755 2524 759
rect 2928 755 2932 759
rect 3056 755 3060 759
rect 3191 755 3195 759
rect 2208 751 2212 755
rect 2664 751 2668 755
rect 2800 751 2804 755
rect 3168 751 3172 755
rect 111 733 115 737
rect 1424 735 1428 739
rect 584 731 588 735
rect 712 731 716 735
rect 840 731 844 735
rect 960 731 964 735
rect 1080 731 1084 735
rect 1192 731 1196 735
rect 1304 731 1308 735
rect 1631 733 1635 737
rect 1671 733 1675 737
rect 2928 735 2932 739
rect 2136 731 2140 735
rect 2296 731 2300 735
rect 2456 731 2460 735
rect 2608 731 2612 735
rect 2768 731 2772 735
rect 3191 733 3195 737
rect 111 715 115 719
rect 1631 715 1635 719
rect 1671 715 1675 719
rect 3191 715 3195 719
rect 1671 689 1675 693
rect 3191 689 3195 693
rect 111 677 115 681
rect 1631 677 1635 681
rect 1671 671 1675 675
rect 3000 671 3004 675
rect 3168 671 3172 675
rect 3191 671 3195 675
rect 2032 667 2036 671
rect 2160 667 2164 671
rect 2304 667 2308 671
rect 2456 667 2460 671
rect 2624 667 2628 671
rect 2808 667 2812 671
rect 111 659 115 663
rect 1200 659 1204 663
rect 1320 659 1324 663
rect 1631 659 1635 663
rect 488 655 492 659
rect 616 655 620 659
rect 736 655 740 659
rect 856 655 860 659
rect 976 655 980 659
rect 1088 655 1092 659
rect 1671 645 1675 649
rect 2768 647 2772 651
rect 1928 643 1932 647
rect 2056 643 2060 647
rect 2192 643 2196 647
rect 2336 643 2340 647
rect 2480 643 2484 647
rect 2624 643 2628 647
rect 3191 645 3195 649
rect 111 629 115 633
rect 752 631 756 635
rect 1224 631 1228 635
rect 384 627 388 631
rect 512 627 516 631
rect 632 627 636 631
rect 872 627 876 631
rect 984 627 988 631
rect 1104 627 1108 631
rect 1631 629 1635 633
rect 1671 627 1675 631
rect 3191 627 3195 631
rect 111 611 115 615
rect 1631 611 1635 615
rect 1671 597 1675 601
rect 3191 597 3195 601
rect 111 577 115 581
rect 1631 577 1635 581
rect 1671 579 1675 583
rect 2192 579 2196 583
rect 2760 579 2764 583
rect 2968 581 2972 585
rect 3168 579 3172 583
rect 3191 579 3195 583
rect 1856 575 1860 579
rect 2024 575 2028 579
rect 2368 575 2372 579
rect 2560 575 2564 579
rect 111 559 115 563
rect 776 559 780 563
rect 1631 559 1635 563
rect 1671 561 1675 565
rect 1776 563 1780 567
rect 2256 563 2260 567
rect 2416 563 2420 567
rect 1936 559 1940 563
rect 2096 559 2100 563
rect 2576 559 2580 563
rect 3191 561 3195 565
rect 280 555 284 559
rect 408 555 412 559
rect 536 555 540 559
rect 656 555 660 559
rect 888 555 892 559
rect 1000 555 1004 559
rect 1120 555 1124 559
rect 1671 543 1675 547
rect 3191 543 3195 547
rect 111 529 115 533
rect 432 531 436 535
rect 784 531 788 535
rect 184 527 188 531
rect 312 527 316 531
rect 552 527 556 531
rect 672 527 676 531
rect 896 527 900 531
rect 1016 527 1020 531
rect 1631 529 1635 533
rect 1671 517 1675 521
rect 3191 517 3195 521
rect 111 511 115 515
rect 1631 511 1635 515
rect 1671 499 1675 503
rect 1896 499 1900 503
rect 2112 499 2116 503
rect 2352 499 2356 503
rect 3144 499 3148 503
rect 3191 499 3195 503
rect 1704 495 1708 499
rect 2608 495 2612 499
rect 2872 495 2876 499
rect 111 473 115 477
rect 1631 473 1635 477
rect 1671 473 1675 477
rect 1704 475 1708 479
rect 2032 475 2036 479
rect 2392 475 2396 479
rect 3120 475 3124 479
rect 2752 471 2756 475
rect 3191 473 3195 477
rect 111 455 115 459
rect 144 455 148 459
rect 240 455 244 459
rect 368 455 372 459
rect 512 455 516 459
rect 664 453 668 457
rect 1144 455 1148 459
rect 1631 455 1635 459
rect 1671 455 1675 459
rect 3191 455 3195 459
rect 824 451 828 455
rect 984 451 988 455
rect 1304 451 1308 455
rect 1464 451 1468 455
rect 1608 451 1612 455
rect 111 425 115 429
rect 1112 427 1116 431
rect 1232 427 1236 431
rect 1456 429 1460 433
rect 1576 427 1580 431
rect 736 423 740 427
rect 864 423 868 427
rect 992 423 996 427
rect 1344 423 1348 427
rect 1631 425 1635 429
rect 1671 425 1675 429
rect 3191 425 3195 429
rect 111 407 115 411
rect 1631 407 1635 411
rect 1671 407 1675 411
rect 2864 407 2868 411
rect 3096 407 3100 411
rect 3191 407 3195 411
rect 2256 403 2260 407
rect 2384 403 2388 407
rect 2512 403 2516 407
rect 2632 403 2636 407
rect 2752 403 2756 407
rect 2976 403 2980 407
rect 1671 377 1675 381
rect 2672 379 2676 383
rect 2800 379 2804 383
rect 2928 379 2932 383
rect 111 373 115 377
rect 1631 373 1635 377
rect 2160 375 2164 379
rect 2288 375 2292 379
rect 2416 375 2420 379
rect 2544 375 2548 379
rect 3056 375 3060 379
rect 3168 375 3172 379
rect 3191 377 3195 381
rect 1671 359 1675 363
rect 3191 359 3195 363
rect 111 355 115 359
rect 656 355 660 359
rect 1472 355 1476 359
rect 1631 355 1635 359
rect 816 351 820 355
rect 960 351 964 355
rect 1096 351 1100 355
rect 1224 351 1228 355
rect 1344 351 1348 355
rect 111 333 115 337
rect 952 335 956 339
rect 1088 335 1092 339
rect 1232 335 1236 339
rect 1376 335 1380 339
rect 552 331 556 335
rect 680 331 684 335
rect 816 331 820 335
rect 1631 333 1635 337
rect 1671 321 1675 325
rect 3191 321 3195 325
rect 111 315 115 319
rect 1631 315 1635 319
rect 1671 303 1675 307
rect 2440 303 2444 307
rect 2872 303 2876 307
rect 3032 303 3036 307
rect 3168 303 3172 307
rect 3191 303 3195 307
rect 2056 299 2060 303
rect 2184 299 2188 303
rect 2312 299 2316 303
rect 2576 299 2580 303
rect 2720 299 2724 303
rect 111 285 115 289
rect 1631 285 1635 289
rect 1671 277 1675 281
rect 2560 279 2564 283
rect 2672 279 2676 283
rect 2792 279 2796 283
rect 1952 275 1956 279
rect 2080 275 2084 279
rect 2208 275 2212 279
rect 2328 275 2332 279
rect 2448 275 2452 279
rect 3191 277 3195 281
rect 111 267 115 271
rect 472 267 476 271
rect 776 267 780 271
rect 1296 267 1300 271
rect 1631 267 1635 271
rect 632 263 636 267
rect 912 263 916 267
rect 1040 263 1044 267
rect 1168 263 1172 267
rect 1671 259 1675 263
rect 3191 259 3195 263
rect 111 245 115 249
rect 368 247 372 251
rect 496 243 500 247
rect 632 243 636 247
rect 768 245 772 249
rect 904 247 908 251
rect 1192 247 1196 251
rect 1048 243 1052 247
rect 1631 245 1635 249
rect 111 227 115 231
rect 1631 227 1635 231
rect 1671 221 1675 225
rect 3191 221 3195 225
rect 1671 203 1675 207
rect 2776 203 2780 207
rect 2976 203 2980 207
rect 3168 203 3172 207
rect 3191 203 3195 207
rect 111 197 115 201
rect 1631 197 1635 201
rect 1856 199 1860 203
rect 1984 199 1988 203
rect 2112 199 2116 203
rect 2256 199 2260 203
rect 2416 199 2420 203
rect 2592 199 2596 203
rect 111 179 115 183
rect 288 179 292 183
rect 456 179 460 183
rect 952 179 956 183
rect 1631 179 1635 183
rect 624 175 628 179
rect 784 175 788 179
rect 1120 175 1124 179
rect 1671 173 1675 177
rect 2152 175 2156 179
rect 2320 175 2324 179
rect 2504 175 2508 179
rect 1752 171 1756 175
rect 1880 171 1884 175
rect 2008 171 2012 175
rect 2712 173 2716 177
rect 2928 175 2932 179
rect 3144 175 3148 179
rect 3191 173 3195 177
rect 111 161 115 165
rect 208 163 212 167
rect 376 163 380 167
rect 1040 163 1044 167
rect 544 159 548 163
rect 704 159 708 163
rect 872 159 876 163
rect 1631 161 1635 165
rect 1671 155 1675 159
rect 3191 155 3195 159
rect 111 143 115 147
rect 1631 143 1635 147
rect 1671 113 1675 117
rect 3191 113 3195 117
rect 111 105 115 109
rect 1631 105 1635 109
rect 1671 95 1675 99
rect 2360 95 2364 99
rect 2528 95 2532 99
rect 2720 95 2724 99
rect 2920 95 2924 99
rect 3120 95 3124 99
rect 3191 95 3195 99
rect 1704 91 1708 95
rect 1824 91 1828 95
rect 1952 91 1956 95
rect 2080 91 2084 95
rect 2208 91 2212 95
rect 111 87 115 91
rect 144 87 148 91
rect 200 87 204 91
rect 296 87 300 91
rect 392 87 396 91
rect 488 87 492 91
rect 592 87 596 91
rect 704 87 708 91
rect 824 87 828 91
rect 952 87 956 91
rect 1088 87 1092 91
rect 1224 87 1228 91
rect 1360 87 1364 91
rect 1496 87 1500 91
rect 1608 87 1612 91
rect 1631 87 1635 91
<< m2 >>
rect 3054 3304 3060 3305
rect 3054 3300 3055 3304
rect 3059 3300 3060 3304
rect 3054 3299 3060 3300
rect 1670 3297 1676 3298
rect 1670 3293 1671 3297
rect 1675 3293 1676 3297
rect 1670 3292 1676 3293
rect 3190 3297 3196 3298
rect 3190 3293 3191 3297
rect 3195 3293 3196 3297
rect 3190 3292 3196 3293
rect 1670 3279 1676 3280
rect 1670 3275 1671 3279
rect 1675 3275 1676 3279
rect 3190 3279 3196 3280
rect 1670 3274 1676 3275
rect 3054 3275 3060 3276
rect 3054 3271 3055 3275
rect 3059 3271 3060 3275
rect 3054 3270 3060 3271
rect 3063 3275 3069 3276
rect 3063 3271 3064 3275
rect 3068 3274 3069 3275
rect 3118 3275 3124 3276
rect 3118 3274 3119 3275
rect 3068 3272 3119 3274
rect 3068 3271 3069 3272
rect 3063 3270 3069 3271
rect 3118 3271 3119 3272
rect 3123 3271 3124 3275
rect 3190 3275 3191 3279
rect 3195 3275 3196 3279
rect 3190 3274 3196 3275
rect 3118 3270 3124 3271
rect 2150 3265 2156 3266
rect 1670 3261 1676 3262
rect 1670 3257 1671 3261
rect 1675 3257 1676 3261
rect 2150 3261 2151 3265
rect 2155 3261 2156 3265
rect 2150 3260 2156 3261
rect 2286 3265 2292 3266
rect 2286 3261 2287 3265
rect 2291 3261 2292 3265
rect 2286 3260 2292 3261
rect 2422 3265 2428 3266
rect 2422 3261 2423 3265
rect 2427 3261 2428 3265
rect 2422 3260 2428 3261
rect 2566 3265 2572 3266
rect 2566 3261 2567 3265
rect 2571 3261 2572 3265
rect 2566 3260 2572 3261
rect 2710 3265 2716 3266
rect 2710 3261 2711 3265
rect 2715 3261 2716 3265
rect 2710 3260 2716 3261
rect 2854 3265 2860 3266
rect 2854 3261 2855 3265
rect 2859 3261 2860 3265
rect 2854 3260 2860 3261
rect 2998 3265 3004 3266
rect 2998 3261 2999 3265
rect 3003 3261 3004 3265
rect 2998 3260 3004 3261
rect 3007 3263 3013 3264
rect 1670 3256 1676 3257
rect 2159 3259 2165 3260
rect 2159 3255 2160 3259
rect 2164 3258 2165 3259
rect 2182 3259 2188 3260
rect 2182 3258 2183 3259
rect 2164 3256 2183 3258
rect 2164 3255 2165 3256
rect 2159 3254 2165 3255
rect 2182 3255 2183 3256
rect 2187 3255 2188 3259
rect 2182 3254 2188 3255
rect 2295 3259 2301 3260
rect 2295 3255 2296 3259
rect 2300 3258 2301 3259
rect 2431 3259 2437 3260
rect 2431 3258 2432 3259
rect 2300 3256 2432 3258
rect 2300 3255 2301 3256
rect 2295 3254 2301 3255
rect 2431 3255 2432 3256
rect 2436 3258 2437 3259
rect 2554 3259 2560 3260
rect 2554 3258 2555 3259
rect 2436 3256 2555 3258
rect 2436 3255 2437 3256
rect 2431 3254 2437 3255
rect 2554 3255 2555 3256
rect 2559 3258 2560 3259
rect 2575 3259 2581 3260
rect 2575 3258 2576 3259
rect 2559 3256 2576 3258
rect 2559 3255 2560 3256
rect 2554 3254 2560 3255
rect 2575 3255 2576 3256
rect 2580 3258 2581 3259
rect 2719 3259 2725 3260
rect 2719 3258 2720 3259
rect 2580 3256 2720 3258
rect 2580 3255 2581 3256
rect 2575 3254 2581 3255
rect 2719 3255 2720 3256
rect 2724 3258 2725 3259
rect 2734 3259 2740 3260
rect 2734 3258 2735 3259
rect 2724 3256 2735 3258
rect 2724 3255 2725 3256
rect 2719 3254 2725 3255
rect 2734 3255 2735 3256
rect 2739 3258 2740 3259
rect 2863 3259 2869 3260
rect 2863 3258 2864 3259
rect 2739 3256 2864 3258
rect 2739 3255 2740 3256
rect 2734 3254 2740 3255
rect 2863 3255 2864 3256
rect 2868 3258 2869 3259
rect 3007 3259 3008 3263
rect 3012 3262 3013 3263
rect 3064 3262 3066 3270
rect 3012 3260 3066 3262
rect 3190 3261 3196 3262
rect 3012 3259 3013 3260
rect 3007 3258 3013 3259
rect 2868 3256 3010 3258
rect 3190 3257 3191 3261
rect 3195 3257 3196 3261
rect 3190 3256 3196 3257
rect 2868 3255 2869 3256
rect 2863 3254 2869 3255
rect 1670 3243 1676 3244
rect 1670 3239 1671 3243
rect 1675 3239 1676 3243
rect 1670 3238 1676 3239
rect 3190 3243 3196 3244
rect 3190 3239 3191 3243
rect 3195 3239 3196 3243
rect 3190 3238 3196 3239
rect 2150 3236 2156 3237
rect 2150 3232 2151 3236
rect 2155 3232 2156 3236
rect 2150 3231 2156 3232
rect 2286 3236 2292 3237
rect 2286 3232 2287 3236
rect 2291 3232 2292 3236
rect 2286 3231 2292 3232
rect 2422 3236 2428 3237
rect 2422 3232 2423 3236
rect 2427 3232 2428 3236
rect 2422 3231 2428 3232
rect 2566 3236 2572 3237
rect 2566 3232 2567 3236
rect 2571 3232 2572 3236
rect 2566 3231 2572 3232
rect 2710 3236 2716 3237
rect 2710 3232 2711 3236
rect 2715 3232 2716 3236
rect 2710 3231 2716 3232
rect 2854 3236 2860 3237
rect 2854 3232 2855 3236
rect 2859 3232 2860 3236
rect 2854 3231 2860 3232
rect 2998 3236 3004 3237
rect 2998 3232 2999 3236
rect 3003 3232 3004 3236
rect 2998 3231 3004 3232
rect 1998 3224 2004 3225
rect 1998 3220 1999 3224
rect 2003 3220 2004 3224
rect 1998 3219 2004 3220
rect 2174 3224 2180 3225
rect 2174 3220 2175 3224
rect 2179 3220 2180 3224
rect 2174 3219 2180 3220
rect 2358 3224 2364 3225
rect 2358 3220 2359 3224
rect 2363 3220 2364 3224
rect 2358 3219 2364 3220
rect 2542 3224 2548 3225
rect 2542 3220 2543 3224
rect 2547 3220 2548 3224
rect 2542 3219 2548 3220
rect 2726 3224 2732 3225
rect 2726 3220 2727 3224
rect 2731 3220 2732 3224
rect 2726 3219 2732 3220
rect 2918 3224 2924 3225
rect 2918 3220 2919 3224
rect 2923 3220 2924 3224
rect 2918 3219 2924 3220
rect 3110 3224 3116 3225
rect 3110 3220 3111 3224
rect 3115 3220 3116 3224
rect 3110 3219 3116 3220
rect 1670 3217 1676 3218
rect 1670 3213 1671 3217
rect 1675 3213 1676 3217
rect 1670 3212 1676 3213
rect 3190 3217 3196 3218
rect 3190 3213 3191 3217
rect 3195 3213 3196 3217
rect 3190 3212 3196 3213
rect 1670 3199 1676 3200
rect 1670 3195 1671 3199
rect 1675 3195 1676 3199
rect 2551 3199 2560 3200
rect 1670 3194 1676 3195
rect 1998 3195 2004 3196
rect 1998 3191 1999 3195
rect 2003 3191 2004 3195
rect 1998 3190 2004 3191
rect 2007 3195 2013 3196
rect 2007 3191 2008 3195
rect 2012 3194 2013 3195
rect 2046 3195 2052 3196
rect 2046 3194 2047 3195
rect 2012 3192 2047 3194
rect 2012 3191 2013 3192
rect 2007 3190 2013 3191
rect 2046 3191 2047 3192
rect 2051 3191 2052 3195
rect 2046 3190 2052 3191
rect 2174 3195 2180 3196
rect 2174 3191 2175 3195
rect 2179 3191 2180 3195
rect 2174 3190 2180 3191
rect 2182 3195 2189 3196
rect 2182 3191 2183 3195
rect 2188 3194 2189 3195
rect 2234 3195 2240 3196
rect 2234 3194 2235 3195
rect 2188 3192 2235 3194
rect 2188 3191 2189 3192
rect 2182 3190 2189 3191
rect 2234 3191 2235 3192
rect 2239 3191 2240 3195
rect 2234 3190 2240 3191
rect 2358 3195 2364 3196
rect 2358 3191 2359 3195
rect 2363 3191 2364 3195
rect 2358 3190 2364 3191
rect 2367 3195 2373 3196
rect 2367 3191 2368 3195
rect 2372 3194 2373 3195
rect 2542 3195 2548 3196
rect 2372 3192 2378 3194
rect 2372 3191 2373 3192
rect 2367 3190 2373 3191
rect 1846 3185 1852 3186
rect 1670 3181 1676 3182
rect 1670 3177 1671 3181
rect 1675 3177 1676 3181
rect 1846 3181 1847 3185
rect 1851 3181 1852 3185
rect 1846 3180 1852 3181
rect 2038 3185 2044 3186
rect 2038 3181 2039 3185
rect 2043 3181 2044 3185
rect 2246 3185 2252 3186
rect 2038 3180 2044 3181
rect 2046 3183 2053 3184
rect 1670 3176 1676 3177
rect 1854 3179 1861 3180
rect 1854 3175 1855 3179
rect 1860 3175 1861 3179
rect 2046 3179 2047 3183
rect 2052 3182 2053 3183
rect 2182 3183 2188 3184
rect 2182 3182 2183 3183
rect 2052 3180 2183 3182
rect 2052 3179 2053 3180
rect 2046 3178 2053 3179
rect 2182 3179 2183 3180
rect 2187 3179 2188 3183
rect 2246 3181 2247 3185
rect 2251 3181 2252 3185
rect 2246 3180 2252 3181
rect 2182 3178 2188 3179
rect 2234 3179 2240 3180
rect 1854 3174 1861 3175
rect 2234 3175 2235 3179
rect 2239 3178 2240 3179
rect 2255 3179 2261 3180
rect 2255 3178 2256 3179
rect 2239 3176 2256 3178
rect 2239 3175 2240 3176
rect 2234 3174 2240 3175
rect 2255 3175 2256 3176
rect 2260 3178 2261 3179
rect 2376 3178 2378 3192
rect 2542 3191 2543 3195
rect 2547 3191 2548 3195
rect 2551 3195 2552 3199
rect 2559 3195 2560 3199
rect 2734 3199 2741 3200
rect 2551 3194 2560 3195
rect 2726 3195 2732 3196
rect 2542 3190 2548 3191
rect 2726 3191 2727 3195
rect 2731 3191 2732 3195
rect 2734 3195 2735 3199
rect 2740 3195 2741 3199
rect 3190 3199 3196 3200
rect 2734 3194 2741 3195
rect 2918 3195 2924 3196
rect 2726 3190 2732 3191
rect 2918 3191 2919 3195
rect 2923 3191 2924 3195
rect 2918 3190 2924 3191
rect 2926 3195 2933 3196
rect 2926 3191 2927 3195
rect 2932 3191 2933 3195
rect 2926 3190 2933 3191
rect 3110 3195 3116 3196
rect 3110 3191 3111 3195
rect 3115 3191 3116 3195
rect 3110 3190 3116 3191
rect 3118 3195 3125 3196
rect 3118 3191 3119 3195
rect 3124 3194 3125 3195
rect 3190 3195 3191 3199
rect 3195 3195 3196 3199
rect 3190 3194 3196 3195
rect 3124 3192 3170 3194
rect 3124 3191 3125 3192
rect 3118 3190 3125 3191
rect 2462 3185 2468 3186
rect 2462 3181 2463 3185
rect 2467 3181 2468 3185
rect 2462 3180 2468 3181
rect 2694 3185 2700 3186
rect 2694 3181 2695 3185
rect 2699 3181 2700 3185
rect 2934 3185 2940 3186
rect 2694 3180 2700 3181
rect 2702 3183 2709 3184
rect 2471 3179 2477 3180
rect 2471 3178 2472 3179
rect 2260 3176 2472 3178
rect 2260 3175 2261 3176
rect 2255 3174 2261 3175
rect 2471 3175 2472 3176
rect 2476 3178 2477 3179
rect 2554 3179 2560 3180
rect 2554 3178 2555 3179
rect 2476 3176 2555 3178
rect 2476 3175 2477 3176
rect 2471 3174 2477 3175
rect 2554 3175 2555 3176
rect 2559 3175 2560 3179
rect 2702 3179 2703 3183
rect 2708 3182 2709 3183
rect 2734 3183 2740 3184
rect 2734 3182 2735 3183
rect 2708 3180 2735 3182
rect 2708 3179 2709 3180
rect 2702 3178 2709 3179
rect 2734 3179 2735 3180
rect 2739 3179 2740 3183
rect 2934 3181 2935 3185
rect 2939 3181 2940 3185
rect 2934 3180 2940 3181
rect 3158 3185 3164 3186
rect 3158 3181 3159 3185
rect 3163 3181 3164 3185
rect 3168 3184 3170 3192
rect 3158 3180 3164 3181
rect 3167 3183 3173 3184
rect 2734 3178 2740 3179
rect 2926 3179 2932 3180
rect 2554 3174 2560 3175
rect 2926 3175 2927 3179
rect 2931 3178 2932 3179
rect 2943 3179 2949 3180
rect 2943 3178 2944 3179
rect 2931 3176 2944 3178
rect 2931 3175 2932 3176
rect 2926 3174 2932 3175
rect 2943 3175 2944 3176
rect 2948 3175 2949 3179
rect 3167 3179 3168 3183
rect 3172 3179 3173 3183
rect 3167 3178 3173 3179
rect 3190 3181 3196 3182
rect 3190 3177 3191 3181
rect 3195 3177 3196 3181
rect 3190 3176 3196 3177
rect 2943 3174 2949 3175
rect 1670 3163 1676 3164
rect 1670 3159 1671 3163
rect 1675 3159 1676 3163
rect 1670 3158 1676 3159
rect 3190 3163 3196 3164
rect 3190 3159 3191 3163
rect 3195 3159 3196 3163
rect 3190 3158 3196 3159
rect 1846 3156 1852 3157
rect 1846 3152 1847 3156
rect 1851 3152 1852 3156
rect 1846 3151 1852 3152
rect 2038 3156 2044 3157
rect 2038 3152 2039 3156
rect 2043 3152 2044 3156
rect 2038 3151 2044 3152
rect 2246 3156 2252 3157
rect 2246 3152 2247 3156
rect 2251 3152 2252 3156
rect 2246 3151 2252 3152
rect 2462 3156 2468 3157
rect 2462 3152 2463 3156
rect 2467 3152 2468 3156
rect 2462 3151 2468 3152
rect 2694 3156 2700 3157
rect 2694 3152 2695 3156
rect 2699 3152 2700 3156
rect 2694 3151 2700 3152
rect 2934 3156 2940 3157
rect 2934 3152 2935 3156
rect 2939 3152 2940 3156
rect 2934 3151 2940 3152
rect 3158 3156 3164 3157
rect 3158 3152 3159 3156
rect 3163 3152 3164 3156
rect 3158 3151 3164 3152
rect 1694 3144 1700 3145
rect 1694 3140 1695 3144
rect 1699 3140 1700 3144
rect 1694 3139 1700 3140
rect 1862 3144 1868 3145
rect 1862 3140 1863 3144
rect 1867 3140 1868 3144
rect 1862 3139 1868 3140
rect 2022 3144 2028 3145
rect 2022 3140 2023 3144
rect 2027 3140 2028 3144
rect 2022 3139 2028 3140
rect 2182 3144 2188 3145
rect 2182 3140 2183 3144
rect 2187 3140 2188 3144
rect 2182 3139 2188 3140
rect 2342 3144 2348 3145
rect 2342 3140 2343 3144
rect 2347 3140 2348 3144
rect 2342 3139 2348 3140
rect 2510 3144 2516 3145
rect 2510 3140 2511 3144
rect 2515 3140 2516 3144
rect 2510 3139 2516 3140
rect 1670 3137 1676 3138
rect 1670 3133 1671 3137
rect 1675 3133 1676 3137
rect 1670 3132 1676 3133
rect 3190 3137 3196 3138
rect 3190 3133 3191 3137
rect 3195 3133 3196 3137
rect 3190 3132 3196 3133
rect 1854 3127 1860 3128
rect 1854 3126 1855 3127
rect 806 3125 812 3126
rect 110 3121 116 3122
rect 110 3117 111 3121
rect 115 3117 116 3121
rect 806 3121 807 3125
rect 811 3121 812 3125
rect 806 3120 812 3121
rect 1078 3125 1084 3126
rect 1078 3121 1079 3125
rect 1083 3121 1084 3125
rect 1078 3120 1084 3121
rect 1350 3125 1356 3126
rect 1350 3121 1351 3125
rect 1355 3121 1356 3125
rect 1350 3120 1356 3121
rect 1598 3125 1604 3126
rect 1598 3121 1599 3125
rect 1603 3121 1604 3125
rect 1609 3124 1855 3126
rect 1598 3120 1604 3121
rect 1607 3123 1613 3124
rect 110 3116 116 3117
rect 815 3119 821 3120
rect 815 3115 816 3119
rect 820 3118 821 3119
rect 838 3119 844 3120
rect 838 3118 839 3119
rect 820 3116 839 3118
rect 820 3115 821 3116
rect 815 3114 821 3115
rect 838 3115 839 3116
rect 843 3115 844 3119
rect 838 3114 844 3115
rect 1086 3119 1093 3120
rect 1086 3115 1087 3119
rect 1092 3115 1093 3119
rect 1086 3114 1093 3115
rect 1342 3119 1348 3120
rect 1342 3115 1343 3119
rect 1347 3118 1348 3119
rect 1359 3119 1365 3120
rect 1359 3118 1360 3119
rect 1347 3116 1360 3118
rect 1347 3115 1348 3116
rect 1342 3114 1348 3115
rect 1359 3115 1360 3116
rect 1364 3115 1365 3119
rect 1607 3119 1608 3123
rect 1612 3119 1613 3123
rect 1607 3118 1613 3119
rect 1630 3121 1636 3122
rect 1630 3117 1631 3121
rect 1635 3117 1636 3121
rect 1704 3120 1706 3124
rect 1854 3123 1855 3124
rect 1859 3126 1860 3127
rect 1859 3124 1875 3126
rect 1859 3123 1860 3124
rect 1854 3122 1860 3123
rect 1873 3120 1875 3124
rect 1630 3116 1636 3117
rect 1670 3119 1676 3120
rect 1359 3114 1365 3115
rect 1670 3115 1671 3119
rect 1675 3115 1676 3119
rect 1703 3119 1709 3120
rect 1670 3114 1676 3115
rect 1694 3115 1700 3116
rect 1694 3111 1695 3115
rect 1699 3111 1700 3115
rect 1703 3115 1704 3119
rect 1708 3115 1709 3119
rect 1871 3119 1877 3120
rect 1703 3114 1709 3115
rect 1862 3115 1868 3116
rect 1694 3110 1700 3111
rect 1862 3111 1863 3115
rect 1867 3111 1868 3115
rect 1871 3115 1872 3119
rect 1876 3115 1877 3119
rect 2031 3119 2037 3120
rect 1871 3114 1877 3115
rect 2022 3115 2028 3116
rect 1862 3110 1868 3111
rect 1873 3106 1875 3114
rect 2022 3111 2023 3115
rect 2027 3111 2028 3115
rect 2031 3115 2032 3119
rect 2036 3118 2037 3119
rect 2046 3119 2052 3120
rect 2046 3118 2047 3119
rect 2036 3116 2047 3118
rect 2036 3115 2037 3116
rect 2031 3114 2037 3115
rect 2046 3115 2047 3116
rect 2051 3115 2052 3119
rect 2519 3119 2525 3120
rect 2046 3114 2052 3115
rect 2182 3115 2188 3116
rect 2022 3110 2028 3111
rect 2182 3111 2183 3115
rect 2187 3111 2188 3115
rect 2182 3110 2188 3111
rect 2191 3115 2197 3116
rect 2191 3111 2192 3115
rect 2196 3114 2197 3115
rect 2234 3115 2240 3116
rect 2234 3114 2235 3115
rect 2196 3112 2235 3114
rect 2196 3111 2197 3112
rect 2191 3110 2197 3111
rect 2234 3111 2235 3112
rect 2239 3111 2240 3115
rect 2234 3110 2240 3111
rect 2342 3115 2348 3116
rect 2342 3111 2343 3115
rect 2347 3111 2348 3115
rect 2342 3110 2348 3111
rect 2351 3115 2357 3116
rect 2351 3111 2352 3115
rect 2356 3114 2357 3115
rect 2510 3115 2516 3116
rect 2356 3112 2426 3114
rect 2356 3111 2357 3112
rect 2351 3110 2357 3111
rect 1878 3107 1884 3108
rect 1878 3106 1879 3107
rect 1873 3104 1879 3106
rect 110 3103 116 3104
rect 110 3099 111 3103
rect 115 3099 116 3103
rect 110 3098 116 3099
rect 1630 3103 1636 3104
rect 1630 3099 1631 3103
rect 1635 3099 1636 3103
rect 1878 3103 1879 3104
rect 1883 3103 1884 3107
rect 1878 3102 1884 3103
rect 1958 3105 1964 3106
rect 1630 3098 1636 3099
rect 1670 3101 1676 3102
rect 1670 3097 1671 3101
rect 1675 3097 1676 3101
rect 1958 3101 1959 3105
rect 1963 3101 1964 3105
rect 1958 3100 1964 3101
rect 2182 3105 2188 3106
rect 2182 3101 2183 3105
rect 2187 3101 2188 3105
rect 2192 3104 2194 3110
rect 2414 3105 2420 3106
rect 2182 3100 2188 3101
rect 2191 3103 2197 3104
rect 806 3096 812 3097
rect 806 3092 807 3096
rect 811 3092 812 3096
rect 806 3091 812 3092
rect 1078 3096 1084 3097
rect 1078 3092 1079 3096
rect 1083 3092 1084 3096
rect 1078 3091 1084 3092
rect 1350 3096 1356 3097
rect 1350 3092 1351 3096
rect 1355 3092 1356 3096
rect 1350 3091 1356 3092
rect 1598 3096 1604 3097
rect 1670 3096 1676 3097
rect 1878 3099 1884 3100
rect 1598 3092 1599 3096
rect 1603 3092 1604 3096
rect 1878 3095 1879 3099
rect 1883 3098 1884 3099
rect 1967 3099 1973 3100
rect 1967 3098 1968 3099
rect 1883 3096 1968 3098
rect 1883 3095 1884 3096
rect 1878 3094 1884 3095
rect 1967 3095 1968 3096
rect 1972 3098 1973 3099
rect 2046 3099 2052 3100
rect 2046 3098 2047 3099
rect 1972 3096 2047 3098
rect 1972 3095 1973 3096
rect 1967 3094 1973 3095
rect 2046 3095 2047 3096
rect 2051 3095 2052 3099
rect 2191 3099 2192 3103
rect 2196 3099 2197 3103
rect 2414 3101 2415 3105
rect 2419 3101 2420 3105
rect 2424 3104 2426 3112
rect 2510 3111 2511 3115
rect 2515 3111 2516 3115
rect 2519 3115 2520 3119
rect 2524 3118 2525 3119
rect 2554 3119 2560 3120
rect 2554 3118 2555 3119
rect 2524 3116 2555 3118
rect 2524 3115 2525 3116
rect 2519 3114 2525 3115
rect 2554 3115 2555 3116
rect 2559 3115 2560 3119
rect 2554 3114 2560 3115
rect 3190 3119 3196 3120
rect 3190 3115 3191 3119
rect 3195 3115 3196 3119
rect 3190 3114 3196 3115
rect 2510 3110 2516 3111
rect 2414 3100 2420 3101
rect 2423 3103 2429 3104
rect 2191 3098 2197 3099
rect 2423 3099 2424 3103
rect 2428 3102 2429 3103
rect 2520 3102 2522 3114
rect 2428 3100 2522 3102
rect 2654 3105 2660 3106
rect 2654 3101 2655 3105
rect 2659 3101 2660 3105
rect 2902 3105 2908 3106
rect 2654 3100 2660 3101
rect 2662 3103 2669 3104
rect 2428 3099 2429 3100
rect 2423 3098 2429 3099
rect 2662 3099 2663 3103
rect 2668 3102 2669 3103
rect 2702 3103 2708 3104
rect 2702 3102 2703 3103
rect 2668 3100 2703 3102
rect 2668 3099 2669 3100
rect 2662 3098 2669 3099
rect 2702 3099 2703 3100
rect 2707 3099 2708 3103
rect 2902 3101 2903 3105
rect 2907 3101 2908 3105
rect 2902 3100 2908 3101
rect 3158 3105 3164 3106
rect 3158 3101 3159 3105
rect 3163 3101 3164 3105
rect 3158 3100 3164 3101
rect 3190 3101 3196 3102
rect 2702 3098 2708 3099
rect 2910 3099 2917 3100
rect 2046 3094 2052 3095
rect 2910 3095 2911 3099
rect 2916 3098 2917 3099
rect 2926 3099 2932 3100
rect 2926 3098 2927 3099
rect 2916 3096 2927 3098
rect 2916 3095 2917 3096
rect 2910 3094 2917 3095
rect 2926 3095 2927 3096
rect 2931 3095 2932 3099
rect 2926 3094 2932 3095
rect 3166 3099 3173 3100
rect 3166 3095 3167 3099
rect 3172 3095 3173 3099
rect 3190 3097 3191 3101
rect 3195 3097 3196 3101
rect 3190 3096 3196 3097
rect 3166 3094 3173 3095
rect 1598 3091 1604 3092
rect 1670 3083 1676 3084
rect 702 3080 708 3081
rect 702 3076 703 3080
rect 707 3076 708 3080
rect 702 3075 708 3076
rect 830 3080 836 3081
rect 830 3076 831 3080
rect 835 3076 836 3080
rect 830 3075 836 3076
rect 958 3080 964 3081
rect 958 3076 959 3080
rect 963 3076 964 3080
rect 958 3075 964 3076
rect 1078 3080 1084 3081
rect 1078 3076 1079 3080
rect 1083 3076 1084 3080
rect 1078 3075 1084 3076
rect 1198 3080 1204 3081
rect 1198 3076 1199 3080
rect 1203 3076 1204 3080
rect 1198 3075 1204 3076
rect 1310 3080 1316 3081
rect 1310 3076 1311 3080
rect 1315 3076 1316 3080
rect 1310 3075 1316 3076
rect 1422 3080 1428 3081
rect 1422 3076 1423 3080
rect 1427 3076 1428 3080
rect 1422 3075 1428 3076
rect 1542 3080 1548 3081
rect 1542 3076 1543 3080
rect 1547 3076 1548 3080
rect 1670 3079 1671 3083
rect 1675 3079 1676 3083
rect 1670 3078 1676 3079
rect 3190 3083 3196 3084
rect 3190 3079 3191 3083
rect 3195 3079 3196 3083
rect 3190 3078 3196 3079
rect 1542 3075 1548 3076
rect 1958 3076 1964 3077
rect 110 3073 116 3074
rect 110 3069 111 3073
rect 115 3069 116 3073
rect 110 3068 116 3069
rect 1630 3073 1636 3074
rect 1630 3069 1631 3073
rect 1635 3069 1636 3073
rect 1958 3072 1959 3076
rect 1963 3072 1964 3076
rect 1958 3071 1964 3072
rect 2182 3076 2188 3077
rect 2182 3072 2183 3076
rect 2187 3072 2188 3076
rect 2182 3071 2188 3072
rect 2414 3076 2420 3077
rect 2414 3072 2415 3076
rect 2419 3072 2420 3076
rect 2414 3071 2420 3072
rect 2654 3076 2660 3077
rect 2654 3072 2655 3076
rect 2659 3072 2660 3076
rect 2654 3071 2660 3072
rect 2902 3076 2908 3077
rect 2902 3072 2903 3076
rect 2907 3072 2908 3076
rect 2902 3071 2908 3072
rect 3158 3076 3164 3077
rect 3158 3072 3159 3076
rect 3163 3072 3164 3076
rect 3158 3071 3164 3072
rect 1630 3068 1636 3069
rect 1870 3064 1876 3065
rect 1870 3060 1871 3064
rect 1875 3060 1876 3064
rect 1870 3059 1876 3060
rect 2110 3064 2116 3065
rect 2110 3060 2111 3064
rect 2115 3060 2116 3064
rect 2110 3059 2116 3060
rect 2366 3064 2372 3065
rect 2366 3060 2367 3064
rect 2371 3060 2372 3064
rect 2366 3059 2372 3060
rect 2630 3064 2636 3065
rect 2630 3060 2631 3064
rect 2635 3060 2636 3064
rect 2630 3059 2636 3060
rect 2902 3064 2908 3065
rect 2902 3060 2903 3064
rect 2907 3060 2908 3064
rect 2902 3059 2908 3060
rect 3158 3064 3164 3065
rect 3158 3060 3159 3064
rect 3163 3060 3164 3064
rect 3158 3059 3164 3060
rect 1456 3056 1554 3058
rect 1670 3057 1676 3058
rect 110 3055 116 3056
rect 110 3051 111 3055
rect 115 3051 116 3055
rect 838 3055 845 3056
rect 110 3050 116 3051
rect 702 3051 708 3052
rect 702 3047 703 3051
rect 707 3047 708 3051
rect 702 3046 708 3047
rect 710 3051 717 3052
rect 710 3047 711 3051
rect 716 3047 717 3051
rect 710 3046 717 3047
rect 830 3051 836 3052
rect 830 3047 831 3051
rect 835 3047 836 3051
rect 838 3051 839 3055
rect 844 3051 845 3055
rect 1086 3055 1093 3056
rect 838 3050 845 3051
rect 958 3051 964 3052
rect 830 3046 836 3047
rect 958 3047 959 3051
rect 963 3047 964 3051
rect 958 3046 964 3047
rect 966 3051 973 3052
rect 966 3047 967 3051
rect 972 3047 973 3051
rect 966 3046 973 3047
rect 1078 3051 1084 3052
rect 1078 3047 1079 3051
rect 1083 3047 1084 3051
rect 1086 3051 1087 3055
rect 1092 3051 1093 3055
rect 1431 3055 1437 3056
rect 1086 3050 1093 3051
rect 1198 3051 1204 3052
rect 1078 3046 1084 3047
rect 1198 3047 1199 3051
rect 1203 3047 1204 3051
rect 1198 3046 1204 3047
rect 1206 3051 1213 3052
rect 1206 3047 1207 3051
rect 1212 3047 1213 3051
rect 1206 3046 1213 3047
rect 1310 3051 1316 3052
rect 1310 3047 1311 3051
rect 1315 3047 1316 3051
rect 1310 3046 1316 3047
rect 1318 3051 1325 3052
rect 1318 3047 1319 3051
rect 1324 3047 1325 3051
rect 1318 3046 1325 3047
rect 1422 3051 1428 3052
rect 1422 3047 1423 3051
rect 1427 3047 1428 3051
rect 1431 3051 1432 3055
rect 1436 3054 1437 3055
rect 1446 3055 1452 3056
rect 1446 3054 1447 3055
rect 1436 3052 1447 3054
rect 1436 3051 1437 3052
rect 1431 3050 1437 3051
rect 1446 3051 1447 3052
rect 1451 3054 1452 3055
rect 1456 3054 1458 3056
rect 1451 3052 1458 3054
rect 1551 3055 1557 3056
rect 1451 3051 1452 3052
rect 1446 3050 1452 3051
rect 1542 3051 1548 3052
rect 1422 3046 1428 3047
rect 1542 3047 1543 3051
rect 1547 3047 1548 3051
rect 1551 3051 1552 3055
rect 1556 3051 1557 3055
rect 1551 3050 1557 3051
rect 1630 3055 1636 3056
rect 1630 3051 1631 3055
rect 1635 3051 1636 3055
rect 1670 3053 1671 3057
rect 1675 3053 1676 3057
rect 1670 3052 1676 3053
rect 3190 3057 3196 3058
rect 3190 3053 3191 3057
rect 3195 3053 3196 3057
rect 3190 3052 3196 3053
rect 1630 3050 1636 3051
rect 1542 3046 1548 3047
rect 1670 3039 1676 3040
rect 1670 3035 1671 3039
rect 1675 3035 1676 3039
rect 1878 3039 1885 3040
rect 1670 3034 1676 3035
rect 1870 3035 1876 3036
rect 622 3033 628 3034
rect 110 3029 116 3030
rect 110 3025 111 3029
rect 115 3025 116 3029
rect 622 3029 623 3033
rect 627 3029 628 3033
rect 782 3033 788 3034
rect 622 3028 628 3029
rect 630 3031 637 3032
rect 630 3027 631 3031
rect 636 3030 637 3031
rect 710 3031 716 3032
rect 710 3030 711 3031
rect 636 3028 711 3030
rect 636 3027 637 3028
rect 630 3026 637 3027
rect 710 3027 711 3028
rect 715 3027 716 3031
rect 782 3029 783 3033
rect 787 3029 788 3033
rect 926 3033 932 3034
rect 782 3028 788 3029
rect 790 3031 797 3032
rect 710 3026 716 3027
rect 790 3027 791 3031
rect 796 3030 797 3031
rect 838 3031 844 3032
rect 838 3030 839 3031
rect 796 3028 839 3030
rect 796 3027 797 3028
rect 790 3026 797 3027
rect 838 3027 839 3028
rect 843 3027 844 3031
rect 926 3029 927 3033
rect 931 3029 932 3033
rect 1062 3033 1068 3034
rect 926 3028 932 3029
rect 934 3031 941 3032
rect 838 3026 844 3027
rect 934 3027 935 3031
rect 940 3030 941 3031
rect 966 3031 972 3032
rect 966 3030 967 3031
rect 940 3028 967 3030
rect 940 3027 941 3028
rect 934 3026 941 3027
rect 966 3027 967 3028
rect 971 3027 972 3031
rect 1062 3029 1063 3033
rect 1067 3029 1068 3033
rect 1190 3033 1196 3034
rect 1062 3028 1068 3029
rect 1071 3031 1077 3032
rect 966 3026 972 3027
rect 1071 3027 1072 3031
rect 1076 3030 1077 3031
rect 1086 3031 1092 3032
rect 1086 3030 1087 3031
rect 1076 3028 1087 3030
rect 1076 3027 1077 3028
rect 1071 3026 1077 3027
rect 1086 3027 1087 3028
rect 1091 3027 1092 3031
rect 1190 3029 1191 3033
rect 1195 3029 1196 3033
rect 1310 3033 1316 3034
rect 1190 3028 1196 3029
rect 1199 3029 1205 3030
rect 1199 3028 1200 3029
rect 1086 3026 1092 3027
rect 1198 3027 1200 3028
rect 110 3024 116 3025
rect 1198 3023 1199 3027
rect 1204 3025 1205 3029
rect 1310 3029 1311 3033
rect 1315 3029 1316 3033
rect 1310 3028 1316 3029
rect 1438 3033 1444 3034
rect 1438 3029 1439 3033
rect 1443 3029 1444 3033
rect 1438 3028 1444 3029
rect 1446 3031 1453 3032
rect 1203 3024 1205 3025
rect 1318 3027 1325 3028
rect 1203 3023 1204 3024
rect 1198 3022 1204 3023
rect 1318 3023 1319 3027
rect 1324 3026 1325 3027
rect 1342 3027 1348 3028
rect 1342 3026 1343 3027
rect 1324 3024 1343 3026
rect 1324 3023 1325 3024
rect 1318 3022 1325 3023
rect 1342 3023 1343 3024
rect 1347 3023 1348 3027
rect 1446 3027 1447 3031
rect 1452 3027 1453 3031
rect 1870 3031 1871 3035
rect 1875 3031 1876 3035
rect 1878 3035 1879 3039
rect 1884 3035 1885 3039
rect 2639 3039 2645 3040
rect 1878 3034 1885 3035
rect 2110 3035 2116 3036
rect 1870 3030 1876 3031
rect 2110 3031 2111 3035
rect 2115 3031 2116 3035
rect 2110 3030 2116 3031
rect 2119 3035 2125 3036
rect 2119 3031 2120 3035
rect 2124 3034 2125 3035
rect 2134 3035 2140 3036
rect 2134 3034 2135 3035
rect 2124 3032 2135 3034
rect 2124 3031 2125 3032
rect 2119 3030 2125 3031
rect 2134 3031 2135 3032
rect 2139 3031 2140 3035
rect 2134 3030 2140 3031
rect 2366 3035 2372 3036
rect 2366 3031 2367 3035
rect 2371 3031 2372 3035
rect 2366 3030 2372 3031
rect 2375 3035 2381 3036
rect 2375 3031 2376 3035
rect 2380 3034 2381 3035
rect 2630 3035 2636 3036
rect 2380 3031 2382 3034
rect 2375 3030 2382 3031
rect 2630 3031 2631 3035
rect 2635 3031 2636 3035
rect 2639 3035 2640 3039
rect 2644 3038 2645 3039
rect 2662 3039 2668 3040
rect 2662 3038 2663 3039
rect 2644 3036 2663 3038
rect 2644 3035 2645 3036
rect 2639 3034 2645 3035
rect 2662 3035 2663 3036
rect 2667 3035 2668 3039
rect 3166 3039 3173 3040
rect 2662 3034 2668 3035
rect 2902 3035 2908 3036
rect 2630 3030 2636 3031
rect 1446 3026 1453 3027
rect 1630 3029 1636 3030
rect 1630 3025 1631 3029
rect 1635 3025 1636 3029
rect 1630 3024 1636 3025
rect 1790 3025 1796 3026
rect 1342 3022 1348 3023
rect 1670 3021 1676 3022
rect 1670 3017 1671 3021
rect 1675 3017 1676 3021
rect 1790 3021 1791 3025
rect 1795 3021 1796 3025
rect 1790 3020 1796 3021
rect 1958 3025 1964 3026
rect 1958 3021 1959 3025
rect 1963 3021 1964 3025
rect 1958 3020 1964 3021
rect 2126 3025 2132 3026
rect 2126 3021 2127 3025
rect 2131 3021 2132 3025
rect 2126 3020 2132 3021
rect 2286 3025 2292 3026
rect 2286 3021 2287 3025
rect 2291 3021 2292 3025
rect 2286 3020 2292 3021
rect 2294 3023 2301 3024
rect 1670 3016 1676 3017
rect 1714 3019 1720 3020
rect 1714 3015 1715 3019
rect 1719 3018 1720 3019
rect 1799 3019 1805 3020
rect 1799 3018 1800 3019
rect 1719 3016 1800 3018
rect 1719 3015 1720 3016
rect 1714 3014 1720 3015
rect 1799 3015 1800 3016
rect 1804 3015 1805 3019
rect 1799 3014 1805 3015
rect 1878 3019 1884 3020
rect 1878 3015 1879 3019
rect 1883 3018 1884 3019
rect 1910 3019 1916 3020
rect 1910 3018 1911 3019
rect 1883 3016 1911 3018
rect 1883 3015 1884 3016
rect 1878 3014 1884 3015
rect 1910 3015 1911 3016
rect 1915 3018 1916 3019
rect 1967 3019 1973 3020
rect 1967 3018 1968 3019
rect 1915 3016 1968 3018
rect 1915 3015 1916 3016
rect 1910 3014 1916 3015
rect 1967 3015 1968 3016
rect 1972 3015 1973 3019
rect 1967 3014 1973 3015
rect 2134 3019 2141 3020
rect 2134 3015 2135 3019
rect 2140 3015 2141 3019
rect 2294 3019 2295 3023
rect 2300 3022 2301 3023
rect 2380 3022 2382 3030
rect 2300 3020 2382 3022
rect 2454 3025 2460 3026
rect 2454 3021 2455 3025
rect 2459 3021 2460 3025
rect 2454 3020 2460 3021
rect 2622 3025 2628 3026
rect 2622 3021 2623 3025
rect 2627 3021 2628 3025
rect 2622 3020 2628 3021
rect 2631 3023 2637 3024
rect 2631 3020 2632 3023
rect 2300 3019 2301 3020
rect 2294 3018 2301 3019
rect 2378 3019 2384 3020
rect 2134 3014 2141 3015
rect 2378 3015 2379 3019
rect 2383 3018 2384 3019
rect 2463 3019 2469 3020
rect 2463 3018 2464 3019
rect 2383 3016 2464 3018
rect 2383 3015 2384 3016
rect 2378 3014 2384 3015
rect 2463 3015 2464 3016
rect 2468 3018 2469 3019
rect 2526 3019 2532 3020
rect 2526 3018 2527 3019
rect 2468 3016 2527 3018
rect 2468 3015 2469 3016
rect 2463 3014 2469 3015
rect 2526 3015 2527 3016
rect 2531 3018 2532 3019
rect 2630 3019 2632 3020
rect 2636 3022 2637 3023
rect 2640 3022 2642 3034
rect 2902 3031 2903 3035
rect 2907 3031 2908 3035
rect 2902 3030 2908 3031
rect 2910 3035 2917 3036
rect 2910 3031 2911 3035
rect 2916 3031 2917 3035
rect 2910 3030 2917 3031
rect 3158 3035 3164 3036
rect 3158 3031 3159 3035
rect 3163 3031 3164 3035
rect 3166 3035 3167 3039
rect 3172 3035 3173 3039
rect 3166 3034 3173 3035
rect 3190 3039 3196 3040
rect 3190 3035 3191 3039
rect 3195 3035 3196 3039
rect 3190 3034 3196 3035
rect 3158 3030 3164 3031
rect 2636 3020 2642 3022
rect 3190 3021 3196 3022
rect 2636 3019 2637 3020
rect 2630 3018 2631 3019
rect 2531 3016 2631 3018
rect 2531 3015 2532 3016
rect 2526 3014 2532 3015
rect 2630 3015 2631 3016
rect 2635 3018 2637 3019
rect 2635 3015 2636 3018
rect 3190 3017 3191 3021
rect 3195 3017 3196 3021
rect 3190 3016 3196 3017
rect 2630 3014 2636 3015
rect 110 3011 116 3012
rect 110 3007 111 3011
rect 115 3007 116 3011
rect 110 3006 116 3007
rect 1630 3011 1636 3012
rect 1630 3007 1631 3011
rect 1635 3007 1636 3011
rect 1630 3006 1636 3007
rect 622 3004 628 3005
rect 622 3000 623 3004
rect 627 3000 628 3004
rect 622 2999 628 3000
rect 782 3004 788 3005
rect 782 3000 783 3004
rect 787 3000 788 3004
rect 782 2999 788 3000
rect 926 3004 932 3005
rect 926 3000 927 3004
rect 931 3000 932 3004
rect 926 2999 932 3000
rect 1062 3004 1068 3005
rect 1062 3000 1063 3004
rect 1067 3000 1068 3004
rect 1062 2999 1068 3000
rect 1190 3004 1196 3005
rect 1190 3000 1191 3004
rect 1195 3000 1196 3004
rect 1190 2999 1196 3000
rect 1310 3004 1316 3005
rect 1310 3000 1311 3004
rect 1315 3000 1316 3004
rect 1310 2999 1316 3000
rect 1438 3004 1444 3005
rect 1438 3000 1439 3004
rect 1443 3000 1444 3004
rect 1438 2999 1444 3000
rect 1670 3003 1676 3004
rect 1670 2999 1671 3003
rect 1675 2999 1676 3003
rect 1670 2998 1676 2999
rect 3190 3003 3196 3004
rect 3190 2999 3191 3003
rect 3195 2999 3196 3003
rect 3190 2998 3196 2999
rect 1790 2996 1796 2997
rect 1790 2992 1791 2996
rect 1795 2992 1796 2996
rect 1790 2991 1796 2992
rect 1958 2996 1964 2997
rect 1958 2992 1959 2996
rect 1963 2992 1964 2996
rect 1958 2991 1964 2992
rect 2126 2996 2132 2997
rect 2126 2992 2127 2996
rect 2131 2992 2132 2996
rect 2126 2991 2132 2992
rect 2286 2996 2292 2997
rect 2286 2992 2287 2996
rect 2291 2992 2292 2996
rect 2286 2991 2292 2992
rect 2454 2996 2460 2997
rect 2454 2992 2455 2996
rect 2459 2992 2460 2996
rect 2454 2991 2460 2992
rect 2622 2996 2628 2997
rect 2622 2992 2623 2996
rect 2627 2992 2628 2996
rect 2622 2991 2628 2992
rect 518 2988 524 2989
rect 518 2984 519 2988
rect 523 2984 524 2988
rect 518 2983 524 2984
rect 646 2988 652 2989
rect 646 2984 647 2988
rect 651 2984 652 2988
rect 646 2983 652 2984
rect 782 2988 788 2989
rect 782 2984 783 2988
rect 787 2984 788 2988
rect 782 2983 788 2984
rect 918 2988 924 2989
rect 918 2984 919 2988
rect 923 2984 924 2988
rect 918 2983 924 2984
rect 1054 2988 1060 2989
rect 1054 2984 1055 2988
rect 1059 2984 1060 2988
rect 1054 2983 1060 2984
rect 1190 2988 1196 2989
rect 1190 2984 1191 2988
rect 1195 2984 1196 2988
rect 1190 2983 1196 2984
rect 1334 2988 1340 2989
rect 1334 2984 1335 2988
rect 1339 2984 1340 2988
rect 1334 2983 1340 2984
rect 1702 2984 1708 2985
rect 110 2981 116 2982
rect 110 2977 111 2981
rect 115 2977 116 2981
rect 110 2976 116 2977
rect 1630 2981 1636 2982
rect 1630 2977 1631 2981
rect 1635 2977 1636 2981
rect 1702 2980 1703 2984
rect 1707 2980 1708 2984
rect 1702 2979 1708 2980
rect 1902 2984 1908 2985
rect 1902 2980 1903 2984
rect 1907 2980 1908 2984
rect 1902 2979 1908 2980
rect 2126 2984 2132 2985
rect 2126 2980 2127 2984
rect 2131 2980 2132 2984
rect 2126 2979 2132 2980
rect 2366 2984 2372 2985
rect 2366 2980 2367 2984
rect 2371 2980 2372 2984
rect 2366 2979 2372 2980
rect 2622 2984 2628 2985
rect 2622 2980 2623 2984
rect 2627 2980 2628 2984
rect 2622 2979 2628 2980
rect 2886 2984 2892 2985
rect 2886 2980 2887 2984
rect 2891 2980 2892 2984
rect 2886 2979 2892 2980
rect 3158 2984 3164 2985
rect 3158 2980 3159 2984
rect 3163 2980 3164 2984
rect 3158 2979 3164 2980
rect 1630 2976 1636 2977
rect 1670 2977 1676 2978
rect 1670 2973 1671 2977
rect 1675 2973 1676 2977
rect 1670 2972 1676 2973
rect 3190 2977 3196 2978
rect 3190 2973 3191 2977
rect 3195 2973 3196 2977
rect 3190 2972 3196 2973
rect 1198 2967 1204 2968
rect 1198 2966 1199 2967
rect 1104 2964 1199 2966
rect 110 2963 116 2964
rect 110 2959 111 2963
rect 115 2959 116 2963
rect 790 2963 797 2964
rect 110 2958 116 2959
rect 518 2959 524 2960
rect 518 2955 519 2959
rect 523 2955 524 2959
rect 518 2954 524 2955
rect 527 2959 533 2960
rect 527 2955 528 2959
rect 532 2955 533 2959
rect 527 2954 533 2955
rect 646 2959 652 2960
rect 646 2955 647 2959
rect 651 2955 652 2959
rect 646 2954 652 2955
rect 655 2959 661 2960
rect 655 2955 656 2959
rect 660 2955 661 2959
rect 655 2954 661 2955
rect 782 2959 788 2960
rect 782 2955 783 2959
rect 787 2955 788 2959
rect 790 2959 791 2963
rect 796 2962 797 2963
rect 802 2963 808 2964
rect 802 2962 803 2963
rect 796 2960 803 2962
rect 796 2959 797 2960
rect 790 2958 797 2959
rect 802 2959 803 2960
rect 807 2959 808 2963
rect 927 2963 933 2964
rect 802 2958 808 2959
rect 918 2959 924 2960
rect 782 2954 788 2955
rect 918 2955 919 2959
rect 923 2955 924 2959
rect 927 2959 928 2963
rect 932 2959 933 2963
rect 1063 2963 1069 2964
rect 927 2958 933 2959
rect 1054 2959 1060 2960
rect 918 2954 924 2955
rect 1054 2955 1055 2959
rect 1059 2955 1060 2959
rect 1063 2959 1064 2963
rect 1068 2962 1069 2963
rect 1086 2963 1092 2964
rect 1086 2962 1087 2963
rect 1068 2960 1087 2962
rect 1068 2959 1069 2960
rect 1063 2958 1069 2959
rect 1086 2959 1087 2960
rect 1091 2962 1092 2963
rect 1102 2963 1108 2964
rect 1102 2962 1103 2963
rect 1091 2960 1103 2962
rect 1091 2959 1092 2960
rect 1086 2958 1092 2959
rect 1102 2959 1103 2960
rect 1107 2959 1108 2963
rect 1198 2963 1199 2964
rect 1203 2964 1204 2967
rect 1203 2963 1205 2964
rect 1198 2962 1200 2963
rect 1102 2958 1108 2959
rect 1190 2959 1196 2960
rect 1054 2954 1060 2955
rect 1190 2955 1191 2959
rect 1195 2955 1196 2959
rect 1199 2959 1200 2962
rect 1204 2959 1205 2963
rect 1630 2963 1636 2964
rect 1199 2958 1205 2959
rect 1334 2959 1340 2960
rect 1190 2954 1196 2955
rect 1334 2955 1335 2959
rect 1339 2955 1340 2959
rect 1334 2954 1340 2955
rect 1342 2959 1349 2960
rect 1342 2955 1343 2959
rect 1348 2955 1349 2959
rect 1630 2959 1631 2963
rect 1635 2959 1636 2963
rect 1630 2958 1636 2959
rect 1670 2959 1676 2960
rect 1342 2954 1349 2955
rect 1670 2955 1671 2959
rect 1675 2955 1676 2959
rect 1711 2959 1720 2960
rect 1670 2954 1676 2955
rect 1702 2955 1708 2956
rect 478 2951 484 2952
rect 478 2947 479 2951
rect 483 2950 484 2951
rect 529 2950 531 2954
rect 630 2951 636 2952
rect 630 2950 631 2951
rect 483 2948 631 2950
rect 483 2947 484 2948
rect 478 2946 484 2947
rect 438 2941 444 2942
rect 110 2937 116 2938
rect 110 2933 111 2937
rect 115 2933 116 2937
rect 438 2937 439 2941
rect 443 2937 444 2941
rect 438 2936 444 2937
rect 598 2941 604 2942
rect 598 2937 599 2941
rect 603 2937 604 2941
rect 609 2940 611 2948
rect 630 2947 631 2948
rect 635 2950 636 2951
rect 657 2950 659 2954
rect 1702 2951 1703 2955
rect 1707 2951 1708 2955
rect 1711 2955 1712 2959
rect 1719 2955 1720 2959
rect 1910 2959 1917 2960
rect 1711 2954 1720 2955
rect 1902 2955 1908 2956
rect 1702 2950 1708 2951
rect 1902 2951 1903 2955
rect 1907 2951 1908 2955
rect 1910 2955 1911 2959
rect 1916 2955 1917 2959
rect 2375 2959 2384 2960
rect 1910 2954 1917 2955
rect 2126 2955 2132 2956
rect 1902 2950 1908 2951
rect 2126 2951 2127 2955
rect 2131 2951 2132 2955
rect 2126 2950 2132 2951
rect 2134 2955 2141 2956
rect 2134 2951 2135 2955
rect 2140 2954 2141 2955
rect 2230 2955 2236 2956
rect 2230 2954 2231 2955
rect 2140 2952 2231 2954
rect 2140 2951 2141 2952
rect 2134 2950 2141 2951
rect 2230 2951 2231 2952
rect 2235 2951 2236 2955
rect 2230 2950 2236 2951
rect 2366 2955 2372 2956
rect 2366 2951 2367 2955
rect 2371 2951 2372 2955
rect 2375 2955 2376 2959
rect 2383 2955 2384 2959
rect 2630 2959 2637 2960
rect 2375 2954 2384 2955
rect 2622 2955 2628 2956
rect 2366 2950 2372 2951
rect 2622 2951 2623 2955
rect 2627 2951 2628 2955
rect 2630 2955 2631 2959
rect 2636 2955 2637 2959
rect 3166 2959 3173 2960
rect 2630 2954 2637 2955
rect 2886 2955 2892 2956
rect 2622 2950 2628 2951
rect 2886 2951 2887 2955
rect 2891 2951 2892 2955
rect 2886 2950 2892 2951
rect 2895 2955 2901 2956
rect 2895 2951 2896 2955
rect 2900 2954 2901 2955
rect 2910 2955 2916 2956
rect 2910 2954 2911 2955
rect 2900 2952 2911 2954
rect 2900 2951 2901 2952
rect 2895 2950 2901 2951
rect 2910 2951 2911 2952
rect 2915 2951 2916 2955
rect 2910 2950 2916 2951
rect 3158 2955 3164 2956
rect 3158 2951 3159 2955
rect 3163 2951 3164 2955
rect 3166 2955 3167 2959
rect 3172 2955 3173 2959
rect 3166 2954 3173 2955
rect 3190 2959 3196 2960
rect 3190 2955 3191 2959
rect 3195 2955 3196 2959
rect 3190 2954 3196 2955
rect 3158 2950 3164 2951
rect 635 2948 681 2950
rect 635 2947 636 2948
rect 630 2946 636 2947
rect 598 2936 604 2937
rect 607 2939 613 2940
rect 110 2932 116 2933
rect 447 2935 453 2936
rect 447 2931 448 2935
rect 452 2934 453 2935
rect 478 2935 484 2936
rect 478 2934 479 2935
rect 452 2932 479 2934
rect 452 2931 453 2932
rect 447 2930 453 2931
rect 478 2931 479 2932
rect 483 2931 484 2935
rect 607 2935 608 2939
rect 612 2935 613 2939
rect 607 2934 613 2935
rect 679 2934 681 2948
rect 2896 2946 2898 2950
rect 1694 2945 1700 2946
rect 758 2941 764 2942
rect 758 2937 759 2941
rect 763 2937 764 2941
rect 758 2936 764 2937
rect 926 2941 932 2942
rect 926 2937 927 2941
rect 931 2937 932 2941
rect 926 2936 932 2937
rect 1094 2941 1100 2942
rect 1094 2937 1095 2941
rect 1099 2937 1100 2941
rect 1094 2936 1100 2937
rect 1262 2941 1268 2942
rect 1262 2937 1263 2941
rect 1267 2937 1268 2941
rect 1262 2936 1268 2937
rect 1438 2941 1444 2942
rect 1438 2937 1439 2941
rect 1443 2937 1444 2941
rect 1598 2941 1604 2942
rect 1438 2936 1444 2937
rect 1446 2939 1453 2940
rect 767 2935 773 2936
rect 767 2934 768 2935
rect 679 2932 768 2934
rect 478 2930 484 2931
rect 767 2931 768 2932
rect 772 2934 773 2935
rect 802 2935 808 2936
rect 802 2934 803 2935
rect 772 2932 803 2934
rect 772 2931 773 2932
rect 767 2930 773 2931
rect 802 2931 803 2932
rect 807 2931 808 2935
rect 802 2930 808 2931
rect 934 2935 941 2936
rect 934 2931 935 2935
rect 940 2931 941 2935
rect 934 2930 941 2931
rect 1102 2935 1109 2936
rect 1102 2931 1103 2935
rect 1108 2931 1109 2935
rect 1102 2930 1109 2931
rect 1271 2935 1277 2936
rect 1271 2931 1272 2935
rect 1276 2934 1277 2935
rect 1342 2935 1348 2936
rect 1342 2934 1343 2935
rect 1276 2932 1343 2934
rect 1276 2931 1277 2932
rect 1271 2930 1277 2931
rect 1342 2931 1343 2932
rect 1347 2934 1348 2935
rect 1446 2935 1447 2939
rect 1452 2935 1453 2939
rect 1598 2937 1599 2941
rect 1603 2937 1604 2941
rect 1670 2941 1676 2942
rect 1598 2936 1604 2937
rect 1630 2937 1636 2938
rect 1446 2934 1453 2935
rect 1607 2935 1613 2936
rect 1347 2932 1450 2934
rect 1347 2931 1348 2932
rect 1342 2930 1348 2931
rect 1607 2931 1608 2935
rect 1612 2934 1613 2935
rect 1612 2932 1614 2934
rect 1630 2933 1631 2937
rect 1635 2933 1636 2937
rect 1670 2937 1671 2941
rect 1675 2937 1676 2941
rect 1694 2941 1695 2945
rect 1699 2941 1700 2945
rect 1934 2945 1940 2946
rect 1694 2940 1700 2941
rect 1703 2943 1709 2944
rect 1703 2939 1704 2943
rect 1708 2942 1709 2943
rect 1714 2943 1720 2944
rect 1714 2942 1715 2943
rect 1708 2940 1715 2942
rect 1708 2939 1709 2940
rect 1703 2938 1709 2939
rect 1714 2939 1715 2940
rect 1719 2939 1720 2943
rect 1934 2941 1935 2945
rect 1939 2941 1940 2945
rect 1934 2940 1940 2941
rect 2222 2945 2228 2946
rect 2222 2941 2223 2945
rect 2227 2941 2228 2945
rect 2518 2945 2524 2946
rect 2294 2943 2300 2944
rect 2294 2942 2295 2943
rect 2222 2940 2228 2941
rect 2239 2940 2295 2942
rect 1714 2938 1720 2939
rect 1910 2939 1916 2940
rect 1670 2936 1676 2937
rect 1630 2932 1636 2933
rect 1612 2931 1616 2932
rect 1607 2930 1611 2931
rect 1610 2927 1611 2930
rect 1615 2930 1616 2931
rect 1704 2930 1706 2938
rect 1910 2935 1911 2939
rect 1915 2938 1916 2939
rect 1943 2939 1949 2940
rect 1943 2938 1944 2939
rect 1915 2936 1944 2938
rect 1915 2935 1916 2936
rect 1910 2934 1916 2935
rect 1943 2935 1944 2936
rect 1948 2935 1949 2939
rect 1943 2934 1949 2935
rect 2230 2939 2237 2940
rect 2230 2935 2231 2939
rect 2236 2938 2237 2939
rect 2239 2938 2241 2940
rect 2294 2939 2295 2940
rect 2299 2939 2300 2943
rect 2518 2941 2519 2945
rect 2523 2941 2524 2945
rect 2822 2945 2828 2946
rect 2518 2940 2524 2941
rect 2526 2943 2533 2944
rect 2294 2938 2300 2939
rect 2526 2939 2527 2943
rect 2532 2939 2533 2943
rect 2822 2941 2823 2945
rect 2827 2941 2828 2945
rect 2822 2940 2828 2941
rect 2839 2944 2898 2946
rect 3134 2945 3140 2946
rect 2839 2940 2841 2944
rect 3134 2941 3135 2945
rect 3139 2941 3140 2945
rect 3134 2940 3140 2941
rect 3142 2943 3149 2944
rect 2526 2938 2533 2939
rect 2831 2939 2841 2940
rect 2236 2936 2241 2938
rect 2236 2935 2237 2936
rect 2230 2934 2237 2935
rect 2831 2935 2832 2939
rect 2839 2936 2841 2939
rect 3142 2939 3143 2943
rect 3148 2942 3149 2943
rect 3166 2943 3172 2944
rect 3166 2942 3167 2943
rect 3148 2940 3167 2942
rect 3148 2939 3149 2940
rect 3142 2938 3149 2939
rect 3166 2939 3167 2940
rect 3171 2939 3172 2943
rect 3166 2938 3172 2939
rect 3190 2941 3196 2942
rect 3190 2937 3191 2941
rect 3195 2937 3196 2941
rect 3190 2936 3196 2937
rect 2839 2935 2840 2936
rect 2831 2934 2840 2935
rect 1615 2928 1706 2930
rect 1615 2927 1616 2928
rect 1610 2926 1616 2927
rect 1670 2923 1676 2924
rect 110 2919 116 2920
rect 110 2915 111 2919
rect 115 2915 116 2919
rect 110 2914 116 2915
rect 1630 2919 1636 2920
rect 1630 2915 1631 2919
rect 1635 2915 1636 2919
rect 1670 2919 1671 2923
rect 1675 2919 1676 2923
rect 1670 2918 1676 2919
rect 3190 2923 3196 2924
rect 3190 2919 3191 2923
rect 3195 2919 3196 2923
rect 3190 2918 3196 2919
rect 1630 2914 1636 2915
rect 1694 2916 1700 2917
rect 438 2912 444 2913
rect 438 2908 439 2912
rect 443 2908 444 2912
rect 438 2907 444 2908
rect 598 2912 604 2913
rect 598 2908 599 2912
rect 603 2908 604 2912
rect 598 2907 604 2908
rect 758 2912 764 2913
rect 758 2908 759 2912
rect 763 2908 764 2912
rect 758 2907 764 2908
rect 926 2912 932 2913
rect 926 2908 927 2912
rect 931 2908 932 2912
rect 926 2907 932 2908
rect 1094 2912 1100 2913
rect 1094 2908 1095 2912
rect 1099 2908 1100 2912
rect 1094 2907 1100 2908
rect 1262 2912 1268 2913
rect 1262 2908 1263 2912
rect 1267 2908 1268 2912
rect 1262 2907 1268 2908
rect 1438 2912 1444 2913
rect 1438 2908 1439 2912
rect 1443 2908 1444 2912
rect 1438 2907 1444 2908
rect 1598 2912 1604 2913
rect 1598 2908 1599 2912
rect 1603 2908 1604 2912
rect 1694 2912 1695 2916
rect 1699 2912 1700 2916
rect 1694 2911 1700 2912
rect 1934 2916 1940 2917
rect 1934 2912 1935 2916
rect 1939 2912 1940 2916
rect 1934 2911 1940 2912
rect 2222 2916 2228 2917
rect 2222 2912 2223 2916
rect 2227 2912 2228 2916
rect 2222 2911 2228 2912
rect 2518 2916 2524 2917
rect 2518 2912 2519 2916
rect 2523 2912 2524 2916
rect 2518 2911 2524 2912
rect 2822 2916 2828 2917
rect 2822 2912 2823 2916
rect 2827 2912 2828 2916
rect 2822 2911 2828 2912
rect 3134 2916 3140 2917
rect 3134 2912 3135 2916
rect 3139 2912 3140 2916
rect 3134 2911 3140 2912
rect 1598 2907 1604 2908
rect 2294 2904 2300 2905
rect 334 2900 340 2901
rect 334 2896 335 2900
rect 339 2896 340 2900
rect 334 2895 340 2896
rect 470 2900 476 2901
rect 470 2896 471 2900
rect 475 2896 476 2900
rect 470 2895 476 2896
rect 622 2900 628 2901
rect 622 2896 623 2900
rect 627 2896 628 2900
rect 622 2895 628 2896
rect 790 2900 796 2901
rect 790 2896 791 2900
rect 795 2896 796 2900
rect 790 2895 796 2896
rect 974 2900 980 2901
rect 974 2896 975 2900
rect 979 2896 980 2900
rect 974 2895 980 2896
rect 1174 2900 1180 2901
rect 1174 2896 1175 2900
rect 1179 2896 1180 2900
rect 1174 2895 1180 2896
rect 1382 2900 1388 2901
rect 1382 2896 1383 2900
rect 1387 2896 1388 2900
rect 1382 2895 1388 2896
rect 1590 2900 1596 2901
rect 1590 2896 1591 2900
rect 1595 2896 1596 2900
rect 2294 2900 2295 2904
rect 2299 2900 2300 2904
rect 2294 2899 2300 2900
rect 2550 2904 2556 2905
rect 2550 2900 2551 2904
rect 2555 2900 2556 2904
rect 2550 2899 2556 2900
rect 2814 2904 2820 2905
rect 2814 2900 2815 2904
rect 2819 2900 2820 2904
rect 2814 2899 2820 2900
rect 3078 2904 3084 2905
rect 3078 2900 3079 2904
rect 3083 2900 3084 2904
rect 3078 2899 3084 2900
rect 1590 2895 1596 2896
rect 1670 2897 1676 2898
rect 110 2893 116 2894
rect 110 2889 111 2893
rect 115 2889 116 2893
rect 110 2888 116 2889
rect 1630 2893 1636 2894
rect 1630 2889 1631 2893
rect 1635 2889 1636 2893
rect 1670 2893 1671 2897
rect 1675 2893 1676 2897
rect 1670 2892 1676 2893
rect 3190 2897 3196 2898
rect 3190 2893 3191 2897
rect 3195 2893 3196 2897
rect 3190 2892 3196 2893
rect 1630 2888 1636 2889
rect 2526 2883 2532 2884
rect 1670 2879 1676 2880
rect 110 2875 116 2876
rect 110 2871 111 2875
rect 115 2871 116 2875
rect 1599 2875 1605 2876
rect 110 2870 116 2871
rect 334 2871 340 2872
rect 334 2867 335 2871
rect 339 2867 340 2871
rect 334 2866 340 2867
rect 343 2871 349 2872
rect 343 2867 344 2871
rect 348 2867 349 2871
rect 343 2866 349 2867
rect 470 2871 476 2872
rect 470 2867 471 2871
rect 475 2867 476 2871
rect 470 2866 476 2867
rect 478 2871 485 2872
rect 478 2867 479 2871
rect 484 2867 485 2871
rect 478 2866 485 2867
rect 622 2871 628 2872
rect 622 2867 623 2871
rect 627 2867 628 2871
rect 622 2866 628 2867
rect 631 2871 637 2872
rect 631 2867 632 2871
rect 636 2870 637 2871
rect 702 2871 708 2872
rect 702 2870 703 2871
rect 636 2868 703 2870
rect 636 2867 637 2868
rect 631 2866 637 2867
rect 702 2867 703 2868
rect 707 2867 708 2871
rect 702 2866 708 2867
rect 790 2871 796 2872
rect 790 2867 791 2871
rect 795 2867 796 2871
rect 790 2866 796 2867
rect 799 2871 808 2872
rect 799 2867 800 2871
rect 807 2867 808 2871
rect 799 2866 808 2867
rect 974 2871 980 2872
rect 974 2867 975 2871
rect 979 2867 980 2871
rect 974 2866 980 2867
rect 982 2871 989 2872
rect 982 2867 983 2871
rect 988 2867 989 2871
rect 982 2866 989 2867
rect 1174 2871 1180 2872
rect 1174 2867 1175 2871
rect 1179 2867 1180 2871
rect 1174 2866 1180 2867
rect 1183 2871 1189 2872
rect 1183 2867 1184 2871
rect 1188 2867 1189 2871
rect 1183 2866 1189 2867
rect 1382 2871 1388 2872
rect 1382 2867 1383 2871
rect 1387 2867 1388 2871
rect 1382 2866 1388 2867
rect 1391 2871 1397 2872
rect 1391 2867 1392 2871
rect 1396 2867 1397 2871
rect 1391 2866 1397 2867
rect 1590 2871 1596 2872
rect 1590 2867 1591 2871
rect 1595 2867 1596 2871
rect 1599 2871 1600 2875
rect 1604 2874 1605 2875
rect 1610 2875 1616 2876
rect 1610 2874 1611 2875
rect 1604 2872 1611 2874
rect 1604 2871 1605 2872
rect 1599 2870 1605 2871
rect 1610 2871 1611 2872
rect 1615 2871 1616 2875
rect 1610 2870 1616 2871
rect 1630 2875 1636 2876
rect 1630 2871 1631 2875
rect 1635 2871 1636 2875
rect 1670 2875 1671 2879
rect 1675 2875 1676 2879
rect 2302 2879 2309 2880
rect 1670 2874 1676 2875
rect 2294 2875 2300 2876
rect 1630 2870 1636 2871
rect 2294 2871 2295 2875
rect 2299 2871 2300 2875
rect 2302 2875 2303 2879
rect 2308 2875 2309 2879
rect 2526 2879 2527 2883
rect 2531 2882 2532 2883
rect 2542 2883 2548 2884
rect 2542 2882 2543 2883
rect 2531 2880 2543 2882
rect 2531 2879 2532 2880
rect 2526 2878 2532 2879
rect 2542 2879 2543 2880
rect 2547 2882 2548 2883
rect 2547 2880 2562 2882
rect 2547 2879 2548 2880
rect 2542 2878 2548 2879
rect 2559 2879 2565 2880
rect 2302 2874 2309 2875
rect 2550 2875 2556 2876
rect 2294 2870 2300 2871
rect 2550 2871 2551 2875
rect 2555 2871 2556 2875
rect 2559 2875 2560 2879
rect 2564 2875 2565 2879
rect 3190 2879 3196 2880
rect 2559 2874 2565 2875
rect 2814 2875 2820 2876
rect 2550 2870 2556 2871
rect 2814 2871 2815 2875
rect 2819 2871 2820 2875
rect 2814 2870 2820 2871
rect 2823 2875 2829 2876
rect 2823 2871 2824 2875
rect 2828 2874 2829 2875
rect 2834 2875 2840 2876
rect 2834 2874 2835 2875
rect 2828 2872 2835 2874
rect 2828 2871 2829 2872
rect 2823 2870 2829 2871
rect 2834 2871 2835 2872
rect 2839 2871 2840 2875
rect 2834 2870 2840 2871
rect 3078 2875 3084 2876
rect 3078 2871 3079 2875
rect 3083 2871 3084 2875
rect 3078 2870 3084 2871
rect 3087 2875 3093 2876
rect 3087 2871 3088 2875
rect 3092 2874 3093 2875
rect 3190 2875 3191 2879
rect 3195 2875 3196 2879
rect 3190 2874 3196 2875
rect 3092 2872 3122 2874
rect 3092 2871 3093 2872
rect 3087 2870 3093 2871
rect 1590 2866 1596 2867
rect 286 2863 292 2864
rect 286 2859 287 2863
rect 291 2862 292 2863
rect 345 2862 347 2866
rect 291 2860 347 2862
rect 1094 2863 1100 2864
rect 291 2859 292 2860
rect 286 2858 292 2859
rect 1094 2859 1095 2863
rect 1099 2862 1100 2863
rect 1102 2863 1108 2864
rect 1102 2862 1103 2863
rect 1099 2860 1103 2862
rect 1099 2859 1100 2860
rect 1094 2858 1100 2859
rect 1102 2859 1103 2860
rect 1107 2862 1108 2863
rect 1184 2862 1186 2866
rect 1107 2860 1186 2862
rect 1342 2863 1348 2864
rect 1107 2859 1108 2860
rect 1102 2858 1108 2859
rect 1342 2859 1343 2863
rect 1347 2862 1348 2863
rect 1392 2862 1394 2866
rect 2206 2865 2212 2866
rect 1347 2860 1394 2862
rect 1670 2861 1676 2862
rect 1347 2859 1348 2860
rect 1342 2858 1348 2859
rect 1670 2857 1671 2861
rect 1675 2857 1676 2861
rect 2206 2861 2207 2865
rect 2211 2861 2212 2865
rect 2374 2865 2380 2866
rect 2206 2860 2212 2861
rect 2215 2863 2221 2864
rect 2215 2859 2216 2863
rect 2220 2862 2221 2863
rect 2302 2863 2308 2864
rect 2302 2862 2303 2863
rect 2220 2860 2303 2862
rect 2220 2859 2221 2860
rect 2215 2858 2221 2859
rect 2302 2859 2303 2860
rect 2307 2859 2308 2863
rect 2374 2861 2375 2865
rect 2379 2861 2380 2865
rect 2374 2860 2380 2861
rect 2534 2865 2540 2866
rect 2534 2861 2535 2865
rect 2539 2861 2540 2865
rect 2678 2865 2684 2866
rect 2534 2860 2540 2861
rect 2542 2863 2549 2864
rect 2302 2858 2308 2859
rect 2382 2859 2389 2860
rect 1670 2856 1676 2857
rect 2382 2855 2383 2859
rect 2388 2855 2389 2859
rect 2542 2859 2543 2863
rect 2548 2859 2549 2863
rect 2678 2861 2679 2865
rect 2683 2861 2684 2865
rect 2678 2860 2684 2861
rect 2822 2865 2828 2866
rect 2822 2861 2823 2865
rect 2827 2861 2828 2865
rect 2822 2860 2828 2861
rect 2966 2865 2972 2866
rect 2966 2861 2967 2865
rect 2971 2861 2972 2865
rect 2966 2860 2972 2861
rect 3110 2865 3116 2866
rect 3110 2861 3111 2865
rect 3115 2861 3116 2865
rect 3120 2864 3122 2872
rect 3110 2860 3116 2861
rect 3119 2863 3125 2864
rect 2542 2858 2549 2859
rect 2686 2859 2693 2860
rect 2382 2854 2389 2855
rect 2686 2855 2687 2859
rect 2692 2855 2693 2859
rect 2686 2854 2693 2855
rect 2831 2859 2840 2860
rect 2831 2855 2832 2859
rect 2839 2855 2840 2859
rect 2831 2854 2840 2855
rect 2974 2859 2981 2860
rect 2974 2855 2975 2859
rect 2980 2855 2981 2859
rect 3119 2859 3120 2863
rect 3124 2862 3125 2863
rect 3142 2863 3148 2864
rect 3142 2862 3143 2863
rect 3124 2860 3143 2862
rect 3124 2859 3125 2860
rect 3119 2858 3125 2859
rect 3142 2859 3143 2860
rect 3147 2862 3148 2863
rect 3166 2863 3172 2864
rect 3166 2862 3167 2863
rect 3147 2860 3167 2862
rect 3147 2859 3148 2860
rect 3142 2858 3148 2859
rect 3166 2859 3167 2860
rect 3171 2859 3172 2863
rect 3166 2858 3172 2859
rect 3190 2861 3196 2862
rect 3190 2857 3191 2861
rect 3195 2857 3196 2861
rect 3190 2856 3196 2857
rect 2974 2854 2981 2855
rect 254 2853 260 2854
rect 110 2849 116 2850
rect 110 2845 111 2849
rect 115 2845 116 2849
rect 254 2849 255 2853
rect 259 2849 260 2853
rect 254 2848 260 2849
rect 414 2853 420 2854
rect 414 2849 415 2853
rect 419 2849 420 2853
rect 414 2848 420 2849
rect 558 2853 564 2854
rect 558 2849 559 2853
rect 563 2849 564 2853
rect 558 2848 564 2849
rect 694 2853 700 2854
rect 694 2849 695 2853
rect 699 2849 700 2853
rect 694 2848 700 2849
rect 822 2853 828 2854
rect 822 2849 823 2853
rect 827 2849 828 2853
rect 822 2848 828 2849
rect 950 2853 956 2854
rect 950 2849 951 2853
rect 955 2849 956 2853
rect 950 2848 956 2849
rect 1086 2853 1092 2854
rect 1086 2849 1087 2853
rect 1091 2849 1092 2853
rect 1086 2848 1092 2849
rect 1630 2849 1636 2850
rect 110 2844 116 2845
rect 263 2847 269 2848
rect 263 2843 264 2847
rect 268 2846 269 2847
rect 286 2847 292 2848
rect 286 2846 287 2847
rect 268 2844 287 2846
rect 268 2843 269 2844
rect 263 2842 269 2843
rect 286 2843 287 2844
rect 291 2843 292 2847
rect 286 2842 292 2843
rect 422 2847 429 2848
rect 422 2843 423 2847
rect 428 2846 429 2847
rect 478 2847 484 2848
rect 478 2846 479 2847
rect 428 2844 479 2846
rect 428 2843 429 2844
rect 422 2842 429 2843
rect 478 2843 479 2844
rect 483 2846 484 2847
rect 567 2847 573 2848
rect 567 2846 568 2847
rect 483 2844 568 2846
rect 483 2843 484 2844
rect 478 2842 484 2843
rect 567 2843 568 2844
rect 572 2843 573 2847
rect 567 2842 573 2843
rect 702 2847 709 2848
rect 702 2843 703 2847
rect 708 2843 709 2847
rect 702 2842 709 2843
rect 802 2847 808 2848
rect 802 2843 803 2847
rect 807 2846 808 2847
rect 831 2847 837 2848
rect 831 2846 832 2847
rect 807 2844 832 2846
rect 807 2843 808 2844
rect 802 2842 808 2843
rect 831 2843 832 2844
rect 836 2846 837 2847
rect 870 2847 876 2848
rect 870 2846 871 2847
rect 836 2844 871 2846
rect 836 2843 837 2844
rect 831 2842 837 2843
rect 870 2843 871 2844
rect 875 2846 876 2847
rect 934 2847 940 2848
rect 934 2846 935 2847
rect 875 2844 935 2846
rect 875 2843 876 2844
rect 870 2842 876 2843
rect 934 2843 935 2844
rect 939 2846 940 2847
rect 959 2847 965 2848
rect 959 2846 960 2847
rect 939 2844 960 2846
rect 939 2843 940 2844
rect 934 2842 940 2843
rect 959 2843 960 2844
rect 964 2846 965 2847
rect 982 2847 988 2848
rect 982 2846 983 2847
rect 964 2844 983 2846
rect 964 2843 965 2844
rect 959 2842 965 2843
rect 982 2843 983 2844
rect 987 2843 988 2847
rect 982 2842 988 2843
rect 1094 2847 1101 2848
rect 1094 2843 1095 2847
rect 1100 2843 1101 2847
rect 1630 2845 1631 2849
rect 1635 2845 1636 2849
rect 1630 2844 1636 2845
rect 1094 2842 1101 2843
rect 1670 2843 1676 2844
rect 1670 2839 1671 2843
rect 1675 2839 1676 2843
rect 1670 2838 1676 2839
rect 3190 2843 3196 2844
rect 3190 2839 3191 2843
rect 3195 2839 3196 2843
rect 3190 2838 3196 2839
rect 2206 2836 2212 2837
rect 2206 2832 2207 2836
rect 2211 2832 2212 2836
rect 110 2831 116 2832
rect 110 2827 111 2831
rect 115 2827 116 2831
rect 110 2826 116 2827
rect 1630 2831 1636 2832
rect 2206 2831 2212 2832
rect 2374 2836 2380 2837
rect 2374 2832 2375 2836
rect 2379 2832 2380 2836
rect 2374 2831 2380 2832
rect 2534 2836 2540 2837
rect 2534 2832 2535 2836
rect 2539 2832 2540 2836
rect 2534 2831 2540 2832
rect 2678 2836 2684 2837
rect 2678 2832 2679 2836
rect 2683 2832 2684 2836
rect 2678 2831 2684 2832
rect 2822 2836 2828 2837
rect 2822 2832 2823 2836
rect 2827 2832 2828 2836
rect 2822 2831 2828 2832
rect 2966 2836 2972 2837
rect 2966 2832 2967 2836
rect 2971 2832 2972 2836
rect 2966 2831 2972 2832
rect 3110 2836 3116 2837
rect 3110 2832 3111 2836
rect 3115 2832 3116 2836
rect 3110 2831 3116 2832
rect 1630 2827 1631 2831
rect 1635 2827 1636 2831
rect 1630 2826 1636 2827
rect 254 2824 260 2825
rect 254 2820 255 2824
rect 259 2820 260 2824
rect 254 2819 260 2820
rect 414 2824 420 2825
rect 414 2820 415 2824
rect 419 2820 420 2824
rect 414 2819 420 2820
rect 558 2824 564 2825
rect 558 2820 559 2824
rect 563 2820 564 2824
rect 558 2819 564 2820
rect 694 2824 700 2825
rect 694 2820 695 2824
rect 699 2820 700 2824
rect 694 2819 700 2820
rect 822 2824 828 2825
rect 822 2820 823 2824
rect 827 2820 828 2824
rect 822 2819 828 2820
rect 950 2824 956 2825
rect 950 2820 951 2824
rect 955 2820 956 2824
rect 950 2819 956 2820
rect 1086 2824 1092 2825
rect 1086 2820 1087 2824
rect 1091 2820 1092 2824
rect 1086 2819 1092 2820
rect 2126 2816 2132 2817
rect 2126 2812 2127 2816
rect 2131 2812 2132 2816
rect 2126 2811 2132 2812
rect 2302 2816 2308 2817
rect 2302 2812 2303 2816
rect 2307 2812 2308 2816
rect 2302 2811 2308 2812
rect 2478 2816 2484 2817
rect 2478 2812 2479 2816
rect 2483 2812 2484 2816
rect 2478 2811 2484 2812
rect 2654 2816 2660 2817
rect 2654 2812 2655 2816
rect 2659 2812 2660 2816
rect 2654 2811 2660 2812
rect 2830 2816 2836 2817
rect 2830 2812 2831 2816
rect 2835 2812 2836 2816
rect 2830 2811 2836 2812
rect 3006 2816 3012 2817
rect 3006 2812 3007 2816
rect 3011 2812 3012 2816
rect 3006 2811 3012 2812
rect 3158 2816 3164 2817
rect 3158 2812 3159 2816
rect 3163 2812 3164 2816
rect 3158 2811 3164 2812
rect 1670 2809 1676 2810
rect 1670 2805 1671 2809
rect 1675 2805 1676 2809
rect 150 2804 156 2805
rect 150 2800 151 2804
rect 155 2800 156 2804
rect 150 2799 156 2800
rect 278 2804 284 2805
rect 278 2800 279 2804
rect 283 2800 284 2804
rect 278 2799 284 2800
rect 398 2804 404 2805
rect 398 2800 399 2804
rect 403 2800 404 2804
rect 398 2799 404 2800
rect 518 2804 524 2805
rect 518 2800 519 2804
rect 523 2800 524 2804
rect 518 2799 524 2800
rect 638 2804 644 2805
rect 638 2800 639 2804
rect 643 2800 644 2804
rect 638 2799 644 2800
rect 750 2804 756 2805
rect 750 2800 751 2804
rect 755 2800 756 2804
rect 750 2799 756 2800
rect 862 2804 868 2805
rect 862 2800 863 2804
rect 867 2800 868 2804
rect 862 2799 868 2800
rect 982 2804 988 2805
rect 1670 2804 1676 2805
rect 3190 2809 3196 2810
rect 3190 2805 3191 2809
rect 3195 2805 3196 2809
rect 3190 2804 3196 2805
rect 982 2800 983 2804
rect 987 2800 988 2804
rect 982 2799 988 2800
rect 110 2797 116 2798
rect 110 2793 111 2797
rect 115 2793 116 2797
rect 110 2792 116 2793
rect 1630 2797 1636 2798
rect 1630 2793 1631 2797
rect 1635 2793 1636 2797
rect 2974 2795 2980 2796
rect 1630 2792 1636 2793
rect 2384 2792 2491 2794
rect 1670 2791 1676 2792
rect 1670 2787 1671 2791
rect 1675 2787 1676 2791
rect 2310 2791 2317 2792
rect 1670 2786 1676 2787
rect 2126 2787 2132 2788
rect 286 2783 292 2784
rect 110 2779 116 2780
rect 110 2775 111 2779
rect 115 2775 116 2779
rect 286 2779 287 2783
rect 291 2782 292 2783
rect 422 2783 428 2784
rect 422 2782 423 2783
rect 291 2780 423 2782
rect 291 2779 292 2780
rect 286 2778 292 2779
rect 407 2779 413 2780
rect 110 2774 116 2775
rect 150 2775 156 2776
rect 150 2771 151 2775
rect 155 2771 156 2775
rect 150 2770 156 2771
rect 158 2775 165 2776
rect 158 2771 159 2775
rect 164 2771 165 2775
rect 158 2770 165 2771
rect 278 2775 284 2776
rect 278 2771 279 2775
rect 283 2771 284 2775
rect 278 2770 284 2771
rect 286 2775 293 2776
rect 286 2771 287 2775
rect 292 2771 293 2775
rect 286 2770 293 2771
rect 398 2775 404 2776
rect 398 2771 399 2775
rect 403 2771 404 2775
rect 407 2775 408 2779
rect 412 2775 413 2779
rect 422 2779 423 2780
rect 427 2782 428 2783
rect 630 2783 636 2784
rect 630 2782 631 2783
rect 427 2780 631 2782
rect 427 2779 428 2780
rect 422 2778 428 2779
rect 527 2779 533 2780
rect 407 2774 413 2775
rect 518 2775 524 2776
rect 398 2770 404 2771
rect 518 2771 519 2775
rect 523 2771 524 2775
rect 527 2775 528 2779
rect 532 2775 533 2779
rect 630 2779 631 2780
rect 635 2782 636 2783
rect 702 2783 708 2784
rect 702 2782 703 2783
rect 635 2780 703 2782
rect 635 2779 636 2780
rect 630 2778 636 2779
rect 647 2779 653 2780
rect 527 2774 533 2775
rect 638 2775 644 2776
rect 518 2770 524 2771
rect 638 2771 639 2775
rect 643 2771 644 2775
rect 647 2775 648 2779
rect 652 2775 653 2779
rect 702 2779 703 2780
rect 707 2782 708 2783
rect 2126 2783 2127 2787
rect 2131 2783 2132 2787
rect 2126 2782 2132 2783
rect 2135 2787 2141 2788
rect 2135 2783 2136 2787
rect 2140 2783 2141 2787
rect 2135 2782 2141 2783
rect 2302 2787 2308 2788
rect 2302 2783 2303 2787
rect 2307 2783 2308 2787
rect 2310 2787 2311 2791
rect 2316 2790 2317 2791
rect 2350 2791 2356 2792
rect 2350 2790 2351 2791
rect 2316 2788 2351 2790
rect 2316 2787 2317 2788
rect 2310 2786 2317 2787
rect 2350 2787 2351 2788
rect 2355 2790 2356 2791
rect 2382 2791 2388 2792
rect 2382 2790 2383 2791
rect 2355 2788 2383 2790
rect 2355 2787 2356 2788
rect 2350 2786 2356 2787
rect 2382 2787 2383 2788
rect 2387 2787 2388 2791
rect 2487 2791 2493 2792
rect 2382 2786 2388 2787
rect 2478 2787 2484 2788
rect 2302 2782 2308 2783
rect 2478 2783 2479 2787
rect 2483 2783 2484 2787
rect 2487 2787 2488 2791
rect 2492 2787 2493 2791
rect 2974 2791 2975 2795
rect 2979 2794 2980 2795
rect 2979 2792 3018 2794
rect 2979 2791 2980 2792
rect 2974 2790 2980 2791
rect 3016 2788 3018 2792
rect 3190 2791 3196 2792
rect 2487 2786 2493 2787
rect 2654 2787 2660 2788
rect 2478 2782 2484 2783
rect 2489 2782 2491 2786
rect 2654 2783 2655 2787
rect 2659 2783 2660 2787
rect 2654 2782 2660 2783
rect 2663 2787 2669 2788
rect 2663 2783 2664 2787
rect 2668 2786 2669 2787
rect 2686 2787 2692 2788
rect 2686 2786 2687 2787
rect 2668 2784 2687 2786
rect 2668 2783 2669 2784
rect 2663 2782 2669 2783
rect 2686 2783 2687 2784
rect 2691 2786 2692 2787
rect 2830 2787 2836 2788
rect 2691 2784 2714 2786
rect 2691 2783 2692 2784
rect 2686 2782 2692 2783
rect 707 2780 762 2782
rect 976 2780 994 2782
rect 707 2779 708 2780
rect 702 2778 708 2779
rect 759 2779 765 2780
rect 647 2774 653 2775
rect 750 2775 756 2776
rect 638 2770 644 2771
rect 750 2771 751 2775
rect 755 2771 756 2775
rect 759 2775 760 2779
rect 764 2775 765 2779
rect 870 2779 877 2780
rect 759 2774 765 2775
rect 862 2775 868 2776
rect 750 2770 756 2771
rect 862 2771 863 2775
rect 867 2771 868 2775
rect 870 2775 871 2779
rect 876 2778 877 2779
rect 966 2779 972 2780
rect 966 2778 967 2779
rect 876 2776 967 2778
rect 876 2775 877 2776
rect 870 2774 877 2775
rect 966 2775 967 2776
rect 971 2778 972 2779
rect 976 2778 978 2780
rect 971 2776 978 2778
rect 991 2779 997 2780
rect 971 2775 972 2776
rect 966 2774 972 2775
rect 982 2775 988 2776
rect 862 2770 868 2771
rect 982 2771 983 2775
rect 987 2771 988 2775
rect 991 2775 992 2779
rect 996 2775 997 2779
rect 991 2774 997 2775
rect 1630 2779 1636 2780
rect 1630 2775 1631 2779
rect 1635 2775 1636 2779
rect 1630 2774 1636 2775
rect 2038 2777 2044 2778
rect 982 2770 988 2771
rect 1670 2773 1676 2774
rect 1670 2769 1671 2773
rect 1675 2769 1676 2773
rect 2038 2773 2039 2777
rect 2043 2773 2044 2777
rect 2038 2772 2044 2773
rect 1670 2768 1676 2769
rect 2022 2771 2028 2772
rect 2022 2767 2023 2771
rect 2027 2770 2028 2771
rect 2047 2771 2053 2772
rect 2047 2770 2048 2771
rect 2027 2768 2048 2770
rect 2027 2767 2028 2768
rect 2022 2766 2028 2767
rect 2047 2767 2048 2768
rect 2052 2770 2053 2771
rect 2136 2770 2138 2782
rect 2489 2780 2546 2782
rect 2206 2777 2212 2778
rect 2206 2773 2207 2777
rect 2211 2773 2212 2777
rect 2206 2772 2212 2773
rect 2374 2777 2380 2778
rect 2374 2773 2375 2777
rect 2379 2773 2380 2777
rect 2534 2777 2540 2778
rect 2374 2772 2380 2773
rect 2382 2775 2389 2776
rect 2215 2771 2221 2772
rect 2215 2770 2216 2771
rect 2052 2768 2216 2770
rect 2052 2767 2053 2768
rect 2047 2766 2053 2767
rect 2215 2767 2216 2768
rect 2220 2770 2221 2771
rect 2230 2771 2236 2772
rect 2230 2770 2231 2771
rect 2220 2768 2231 2770
rect 2220 2767 2221 2768
rect 2215 2766 2221 2767
rect 2230 2767 2231 2768
rect 2235 2767 2236 2771
rect 2382 2771 2383 2775
rect 2388 2771 2389 2775
rect 2534 2773 2535 2777
rect 2539 2773 2540 2777
rect 2544 2776 2546 2780
rect 2702 2777 2708 2778
rect 2534 2772 2540 2773
rect 2543 2775 2549 2776
rect 2382 2770 2389 2771
rect 2543 2771 2544 2775
rect 2548 2774 2549 2775
rect 2558 2775 2564 2776
rect 2558 2774 2559 2775
rect 2548 2772 2559 2774
rect 2548 2771 2549 2772
rect 2543 2770 2549 2771
rect 2558 2771 2559 2772
rect 2563 2771 2564 2775
rect 2702 2773 2703 2777
rect 2707 2773 2708 2777
rect 2702 2772 2708 2773
rect 2712 2772 2714 2784
rect 2830 2783 2831 2787
rect 2835 2783 2836 2787
rect 2830 2782 2836 2783
rect 2838 2787 2845 2788
rect 2838 2783 2839 2787
rect 2844 2783 2845 2787
rect 2838 2782 2845 2783
rect 3006 2787 3012 2788
rect 3006 2783 3007 2787
rect 3011 2783 3012 2787
rect 3006 2782 3012 2783
rect 3014 2787 3021 2788
rect 3014 2783 3015 2787
rect 3020 2783 3021 2787
rect 3014 2782 3021 2783
rect 3158 2787 3164 2788
rect 3158 2783 3159 2787
rect 3163 2783 3164 2787
rect 3158 2782 3164 2783
rect 3166 2787 3173 2788
rect 3166 2783 3167 2787
rect 3172 2783 3173 2787
rect 3190 2787 3191 2791
rect 3195 2787 3196 2791
rect 3190 2786 3196 2787
rect 3166 2782 3173 2783
rect 2870 2777 2876 2778
rect 2870 2773 2871 2777
rect 2875 2773 2876 2777
rect 2870 2772 2876 2773
rect 3190 2773 3196 2774
rect 2558 2770 2564 2771
rect 2711 2771 2717 2772
rect 2230 2766 2236 2767
rect 2711 2767 2712 2771
rect 2716 2770 2717 2771
rect 2838 2771 2844 2772
rect 2838 2770 2839 2771
rect 2716 2768 2839 2770
rect 2716 2767 2717 2768
rect 2711 2766 2717 2767
rect 2838 2767 2839 2768
rect 2843 2770 2844 2771
rect 2879 2771 2885 2772
rect 2879 2770 2880 2771
rect 2843 2768 2880 2770
rect 2843 2767 2844 2768
rect 2838 2766 2844 2767
rect 2879 2767 2880 2768
rect 2884 2767 2885 2771
rect 3190 2769 3191 2773
rect 3195 2769 3196 2773
rect 3190 2768 3196 2769
rect 2879 2766 2885 2767
rect 1670 2755 1676 2756
rect 134 2753 140 2754
rect 110 2749 116 2750
rect 110 2745 111 2749
rect 115 2745 116 2749
rect 134 2749 135 2753
rect 139 2749 140 2753
rect 262 2753 268 2754
rect 134 2748 140 2749
rect 143 2751 149 2752
rect 143 2747 144 2751
rect 148 2750 149 2751
rect 158 2751 164 2752
rect 158 2750 159 2751
rect 148 2748 159 2750
rect 148 2747 149 2748
rect 143 2746 149 2747
rect 158 2747 159 2748
rect 163 2747 164 2751
rect 262 2749 263 2753
rect 267 2749 268 2753
rect 262 2748 268 2749
rect 430 2753 436 2754
rect 430 2749 431 2753
rect 435 2749 436 2753
rect 430 2748 436 2749
rect 622 2753 628 2754
rect 622 2749 623 2753
rect 627 2749 628 2753
rect 838 2753 844 2754
rect 622 2748 628 2749
rect 630 2751 637 2752
rect 158 2746 164 2747
rect 271 2747 277 2748
rect 271 2746 272 2747
rect 110 2744 116 2745
rect 160 2744 272 2746
rect 271 2743 272 2744
rect 276 2746 277 2747
rect 286 2747 292 2748
rect 286 2746 287 2747
rect 276 2744 287 2746
rect 276 2743 277 2744
rect 271 2742 277 2743
rect 286 2743 287 2744
rect 291 2743 292 2747
rect 286 2742 292 2743
rect 422 2747 428 2748
rect 422 2743 423 2747
rect 427 2746 428 2747
rect 439 2747 445 2748
rect 439 2746 440 2747
rect 427 2744 440 2746
rect 427 2743 428 2744
rect 422 2742 428 2743
rect 439 2743 440 2744
rect 444 2743 445 2747
rect 630 2747 631 2751
rect 636 2747 637 2751
rect 838 2749 839 2753
rect 843 2749 844 2753
rect 1070 2753 1076 2754
rect 838 2748 844 2749
rect 847 2751 853 2752
rect 630 2746 637 2747
rect 847 2747 848 2751
rect 852 2750 853 2751
rect 870 2751 876 2752
rect 870 2750 871 2751
rect 852 2748 871 2750
rect 852 2747 853 2748
rect 847 2746 853 2747
rect 870 2747 871 2748
rect 875 2747 876 2751
rect 1070 2749 1071 2753
rect 1075 2749 1076 2753
rect 1070 2748 1076 2749
rect 1318 2753 1324 2754
rect 1318 2749 1319 2753
rect 1323 2749 1324 2753
rect 1318 2748 1324 2749
rect 1566 2753 1572 2754
rect 1566 2749 1567 2753
rect 1571 2749 1572 2753
rect 1566 2748 1572 2749
rect 1574 2751 1581 2752
rect 870 2746 876 2747
rect 1079 2747 1085 2748
rect 439 2742 445 2743
rect 1079 2743 1080 2747
rect 1084 2746 1085 2747
rect 1102 2747 1108 2748
rect 1102 2746 1103 2747
rect 1084 2744 1103 2746
rect 1084 2743 1085 2744
rect 1079 2742 1085 2743
rect 1102 2743 1103 2744
rect 1107 2743 1108 2747
rect 1102 2742 1108 2743
rect 1327 2747 1333 2748
rect 1327 2743 1328 2747
rect 1332 2746 1333 2747
rect 1342 2747 1348 2748
rect 1342 2746 1343 2747
rect 1332 2744 1343 2746
rect 1332 2743 1333 2744
rect 1327 2742 1333 2743
rect 1342 2743 1343 2744
rect 1347 2743 1348 2747
rect 1574 2747 1575 2751
rect 1580 2750 1581 2751
rect 1610 2751 1616 2752
rect 1610 2750 1611 2751
rect 1580 2748 1611 2750
rect 1580 2747 1581 2748
rect 1574 2746 1581 2747
rect 1610 2747 1611 2748
rect 1615 2747 1616 2751
rect 1670 2751 1671 2755
rect 1675 2751 1676 2755
rect 1670 2750 1676 2751
rect 3190 2755 3196 2756
rect 3190 2751 3191 2755
rect 3195 2751 3196 2755
rect 3190 2750 3196 2751
rect 1610 2746 1616 2747
rect 1630 2749 1636 2750
rect 1630 2745 1631 2749
rect 1635 2745 1636 2749
rect 1630 2744 1636 2745
rect 2038 2748 2044 2749
rect 2038 2744 2039 2748
rect 2043 2744 2044 2748
rect 2038 2743 2044 2744
rect 2206 2748 2212 2749
rect 2206 2744 2207 2748
rect 2211 2744 2212 2748
rect 2206 2743 2212 2744
rect 2374 2748 2380 2749
rect 2374 2744 2375 2748
rect 2379 2744 2380 2748
rect 2374 2743 2380 2744
rect 2534 2748 2540 2749
rect 2534 2744 2535 2748
rect 2539 2744 2540 2748
rect 2534 2743 2540 2744
rect 2702 2748 2708 2749
rect 2702 2744 2703 2748
rect 2707 2744 2708 2748
rect 2702 2743 2708 2744
rect 2870 2748 2876 2749
rect 2870 2744 2871 2748
rect 2875 2744 2876 2748
rect 2870 2743 2876 2744
rect 1342 2742 1348 2743
rect 2014 2732 2020 2733
rect 110 2731 116 2732
rect 110 2727 111 2731
rect 115 2727 116 2731
rect 110 2726 116 2727
rect 1630 2731 1636 2732
rect 1630 2727 1631 2731
rect 1635 2727 1636 2731
rect 2014 2728 2015 2732
rect 2019 2728 2020 2732
rect 2014 2727 2020 2728
rect 2198 2732 2204 2733
rect 2198 2728 2199 2732
rect 2203 2728 2204 2732
rect 2198 2727 2204 2728
rect 2382 2732 2388 2733
rect 2382 2728 2383 2732
rect 2387 2728 2388 2732
rect 2382 2727 2388 2728
rect 2574 2732 2580 2733
rect 2574 2728 2575 2732
rect 2579 2728 2580 2732
rect 2574 2727 2580 2728
rect 2774 2732 2780 2733
rect 2774 2728 2775 2732
rect 2779 2728 2780 2732
rect 2774 2727 2780 2728
rect 2974 2732 2980 2733
rect 2974 2728 2975 2732
rect 2979 2728 2980 2732
rect 2974 2727 2980 2728
rect 3158 2732 3164 2733
rect 3158 2728 3159 2732
rect 3163 2728 3164 2732
rect 3158 2727 3164 2728
rect 1630 2726 1636 2727
rect 1670 2725 1676 2726
rect 134 2724 140 2725
rect 134 2720 135 2724
rect 139 2720 140 2724
rect 134 2719 140 2720
rect 262 2724 268 2725
rect 262 2720 263 2724
rect 267 2720 268 2724
rect 262 2719 268 2720
rect 430 2724 436 2725
rect 430 2720 431 2724
rect 435 2720 436 2724
rect 430 2719 436 2720
rect 622 2724 628 2725
rect 622 2720 623 2724
rect 627 2720 628 2724
rect 622 2719 628 2720
rect 838 2724 844 2725
rect 838 2720 839 2724
rect 843 2720 844 2724
rect 838 2719 844 2720
rect 1070 2724 1076 2725
rect 1070 2720 1071 2724
rect 1075 2720 1076 2724
rect 1070 2719 1076 2720
rect 1318 2724 1324 2725
rect 1318 2720 1319 2724
rect 1323 2720 1324 2724
rect 1318 2719 1324 2720
rect 1566 2724 1572 2725
rect 1566 2720 1567 2724
rect 1571 2720 1572 2724
rect 1670 2721 1671 2725
rect 1675 2721 1676 2725
rect 1670 2720 1676 2721
rect 3190 2725 3196 2726
rect 3190 2721 3191 2725
rect 3195 2721 3196 2725
rect 3190 2720 3196 2721
rect 1566 2719 1572 2720
rect 2558 2711 2564 2712
rect 1670 2707 1676 2708
rect 1670 2703 1671 2707
rect 1675 2703 1676 2707
rect 2558 2707 2559 2711
rect 2563 2710 2564 2711
rect 2563 2708 2586 2710
rect 2563 2707 2564 2708
rect 2558 2706 2564 2707
rect 2583 2707 2589 2708
rect 1670 2702 1676 2703
rect 2014 2703 2020 2704
rect 702 2700 708 2701
rect 702 2696 703 2700
rect 707 2696 708 2700
rect 702 2695 708 2696
rect 830 2700 836 2701
rect 830 2696 831 2700
rect 835 2696 836 2700
rect 830 2695 836 2696
rect 958 2700 964 2701
rect 958 2696 959 2700
rect 963 2696 964 2700
rect 958 2695 964 2696
rect 1078 2700 1084 2701
rect 1078 2696 1079 2700
rect 1083 2696 1084 2700
rect 1078 2695 1084 2696
rect 1198 2700 1204 2701
rect 1198 2696 1199 2700
rect 1203 2696 1204 2700
rect 1198 2695 1204 2696
rect 1310 2700 1316 2701
rect 1310 2696 1311 2700
rect 1315 2696 1316 2700
rect 1310 2695 1316 2696
rect 1422 2700 1428 2701
rect 1422 2696 1423 2700
rect 1427 2696 1428 2700
rect 1422 2695 1428 2696
rect 1542 2700 1548 2701
rect 1542 2696 1543 2700
rect 1547 2696 1548 2700
rect 2014 2699 2015 2703
rect 2019 2699 2020 2703
rect 2014 2698 2020 2699
rect 2022 2703 2029 2704
rect 2022 2699 2023 2703
rect 2028 2699 2029 2703
rect 2022 2698 2029 2699
rect 2198 2703 2204 2704
rect 2198 2699 2199 2703
rect 2203 2699 2204 2703
rect 2198 2698 2204 2699
rect 2206 2703 2213 2704
rect 2206 2699 2207 2703
rect 2212 2699 2213 2703
rect 2206 2698 2213 2699
rect 2382 2703 2388 2704
rect 2382 2699 2383 2703
rect 2387 2699 2388 2703
rect 2382 2698 2388 2699
rect 2390 2703 2397 2704
rect 2390 2699 2391 2703
rect 2396 2702 2397 2703
rect 2446 2703 2452 2704
rect 2446 2702 2447 2703
rect 2396 2700 2447 2702
rect 2396 2699 2397 2700
rect 2390 2698 2397 2699
rect 2446 2699 2447 2700
rect 2451 2699 2452 2703
rect 2446 2698 2452 2699
rect 2574 2703 2580 2704
rect 2574 2699 2575 2703
rect 2579 2699 2580 2703
rect 2583 2703 2584 2707
rect 2588 2703 2589 2707
rect 2782 2707 2789 2708
rect 2583 2702 2589 2703
rect 2774 2703 2780 2704
rect 2574 2698 2580 2699
rect 2774 2699 2775 2703
rect 2779 2699 2780 2703
rect 2782 2703 2783 2707
rect 2788 2706 2789 2707
rect 2838 2707 2844 2708
rect 2838 2706 2839 2707
rect 2788 2704 2839 2706
rect 2788 2703 2789 2704
rect 2782 2702 2789 2703
rect 2838 2703 2839 2704
rect 2843 2706 2844 2707
rect 2926 2707 2932 2708
rect 2926 2706 2927 2707
rect 2843 2704 2927 2706
rect 2843 2703 2844 2704
rect 2838 2702 2844 2703
rect 2926 2703 2927 2704
rect 2931 2703 2932 2707
rect 3190 2707 3196 2708
rect 2926 2702 2932 2703
rect 2974 2703 2980 2704
rect 2774 2698 2780 2699
rect 2974 2699 2975 2703
rect 2979 2699 2980 2703
rect 2974 2698 2980 2699
rect 2983 2703 2989 2704
rect 2983 2699 2984 2703
rect 2988 2702 2989 2703
rect 3014 2703 3020 2704
rect 3014 2702 3015 2703
rect 2988 2700 3015 2702
rect 2988 2699 2989 2700
rect 2983 2698 2989 2699
rect 3014 2699 3015 2700
rect 3019 2699 3020 2703
rect 3014 2698 3020 2699
rect 3158 2703 3164 2704
rect 3158 2699 3159 2703
rect 3163 2699 3164 2703
rect 3158 2698 3164 2699
rect 3166 2703 3173 2704
rect 3166 2699 3167 2703
rect 3172 2699 3173 2703
rect 3190 2703 3191 2707
rect 3195 2703 3196 2707
rect 3190 2702 3196 2703
rect 3166 2698 3173 2699
rect 1542 2695 1548 2696
rect 2985 2694 2987 2698
rect 110 2693 116 2694
rect 110 2689 111 2693
rect 115 2689 116 2693
rect 110 2688 116 2689
rect 1630 2693 1636 2694
rect 1630 2689 1631 2693
rect 1635 2689 1636 2693
rect 1630 2688 1636 2689
rect 2976 2692 2987 2694
rect 1998 2685 2004 2686
rect 1670 2681 1676 2682
rect 630 2679 636 2680
rect 110 2675 116 2676
rect 110 2671 111 2675
rect 115 2671 116 2675
rect 630 2675 631 2679
rect 635 2678 636 2679
rect 1342 2679 1348 2680
rect 635 2676 714 2678
rect 635 2675 636 2676
rect 630 2674 636 2675
rect 711 2675 717 2676
rect 110 2670 116 2671
rect 702 2671 708 2672
rect 702 2667 703 2671
rect 707 2667 708 2671
rect 711 2671 712 2675
rect 716 2674 717 2675
rect 742 2675 748 2676
rect 742 2674 743 2675
rect 716 2672 743 2674
rect 716 2671 717 2672
rect 711 2670 717 2671
rect 742 2671 743 2672
rect 747 2671 748 2675
rect 966 2675 973 2676
rect 742 2670 748 2671
rect 830 2671 836 2672
rect 702 2666 708 2667
rect 830 2667 831 2671
rect 835 2667 836 2671
rect 830 2666 836 2667
rect 839 2671 845 2672
rect 839 2667 840 2671
rect 844 2670 845 2671
rect 862 2671 868 2672
rect 862 2670 863 2671
rect 844 2668 863 2670
rect 844 2667 845 2668
rect 839 2666 845 2667
rect 862 2667 863 2668
rect 867 2667 868 2671
rect 862 2666 868 2667
rect 958 2671 964 2672
rect 958 2667 959 2671
rect 963 2667 964 2671
rect 966 2671 967 2675
rect 972 2671 973 2675
rect 1319 2675 1325 2676
rect 966 2670 973 2671
rect 1078 2671 1084 2672
rect 958 2666 964 2667
rect 1078 2667 1079 2671
rect 1083 2667 1084 2671
rect 1078 2666 1084 2667
rect 1087 2671 1093 2672
rect 1087 2667 1088 2671
rect 1092 2670 1093 2671
rect 1102 2671 1108 2672
rect 1102 2670 1103 2671
rect 1092 2668 1103 2670
rect 1092 2667 1093 2668
rect 1087 2666 1093 2667
rect 1102 2667 1103 2668
rect 1107 2667 1108 2671
rect 1102 2666 1108 2667
rect 1198 2671 1204 2672
rect 1198 2667 1199 2671
rect 1203 2667 1204 2671
rect 1198 2666 1204 2667
rect 1206 2671 1213 2672
rect 1206 2667 1207 2671
rect 1212 2667 1213 2671
rect 1206 2666 1213 2667
rect 1310 2671 1316 2672
rect 1310 2667 1311 2671
rect 1315 2667 1316 2671
rect 1319 2671 1320 2675
rect 1324 2674 1325 2675
rect 1342 2675 1343 2679
rect 1347 2678 1348 2679
rect 1446 2679 1452 2680
rect 1446 2678 1447 2679
rect 1347 2676 1447 2678
rect 1347 2675 1348 2676
rect 1342 2674 1348 2675
rect 1431 2675 1438 2676
rect 1324 2672 1346 2674
rect 1324 2671 1325 2672
rect 1319 2670 1325 2671
rect 1422 2671 1428 2672
rect 1310 2666 1316 2667
rect 1422 2667 1423 2671
rect 1427 2667 1428 2671
rect 1431 2671 1432 2675
rect 1436 2672 1438 2675
rect 1446 2675 1447 2676
rect 1451 2678 1452 2679
rect 1451 2676 1554 2678
rect 1670 2677 1671 2681
rect 1675 2677 1676 2681
rect 1998 2681 1999 2685
rect 2003 2681 2004 2685
rect 1998 2680 2004 2681
rect 2174 2685 2180 2686
rect 2174 2681 2175 2685
rect 2179 2681 2180 2685
rect 2174 2680 2180 2681
rect 2358 2685 2364 2686
rect 2358 2681 2359 2685
rect 2363 2681 2364 2685
rect 2550 2685 2556 2686
rect 2358 2680 2364 2681
rect 2367 2683 2373 2684
rect 1670 2676 1676 2677
rect 2006 2679 2013 2680
rect 1451 2675 1452 2676
rect 1446 2674 1452 2675
rect 1551 2675 1557 2676
rect 1436 2671 1437 2672
rect 1431 2670 1437 2671
rect 1542 2671 1548 2672
rect 1422 2666 1428 2667
rect 1542 2667 1543 2671
rect 1547 2667 1548 2671
rect 1551 2671 1552 2675
rect 1556 2674 1557 2675
rect 1574 2675 1580 2676
rect 1574 2674 1575 2675
rect 1556 2672 1575 2674
rect 1556 2671 1557 2672
rect 1551 2670 1557 2671
rect 1574 2671 1575 2672
rect 1579 2671 1580 2675
rect 1574 2670 1580 2671
rect 1630 2675 1636 2676
rect 1630 2671 1631 2675
rect 1635 2671 1636 2675
rect 2006 2675 2007 2679
rect 2012 2678 2013 2679
rect 2022 2679 2028 2680
rect 2022 2678 2023 2679
rect 2012 2676 2023 2678
rect 2012 2675 2013 2676
rect 2006 2674 2013 2675
rect 2022 2675 2023 2676
rect 2027 2678 2028 2679
rect 2183 2679 2189 2680
rect 2183 2678 2184 2679
rect 2027 2676 2184 2678
rect 2027 2675 2028 2676
rect 2022 2674 2028 2675
rect 2183 2675 2184 2676
rect 2188 2678 2189 2679
rect 2206 2679 2212 2680
rect 2206 2678 2207 2679
rect 2188 2676 2207 2678
rect 2188 2675 2189 2676
rect 2183 2674 2189 2675
rect 2206 2675 2207 2676
rect 2211 2675 2212 2679
rect 2206 2674 2212 2675
rect 2350 2679 2356 2680
rect 2350 2675 2351 2679
rect 2355 2678 2356 2679
rect 2367 2679 2368 2683
rect 2372 2682 2373 2683
rect 2390 2683 2396 2684
rect 2390 2682 2391 2683
rect 2372 2680 2391 2682
rect 2372 2679 2373 2680
rect 2367 2678 2373 2679
rect 2390 2679 2391 2680
rect 2395 2679 2396 2683
rect 2550 2681 2551 2685
rect 2555 2681 2556 2685
rect 2758 2685 2764 2686
rect 2550 2680 2556 2681
rect 2558 2683 2565 2684
rect 2390 2678 2396 2679
rect 2558 2679 2559 2683
rect 2564 2679 2565 2683
rect 2758 2681 2759 2685
rect 2763 2681 2764 2685
rect 2966 2685 2972 2686
rect 2758 2680 2764 2681
rect 2767 2683 2773 2684
rect 2558 2678 2565 2679
rect 2767 2679 2768 2683
rect 2772 2682 2773 2683
rect 2782 2683 2788 2684
rect 2782 2682 2783 2683
rect 2772 2680 2783 2682
rect 2772 2679 2773 2680
rect 2767 2678 2773 2679
rect 2782 2679 2783 2680
rect 2787 2679 2788 2683
rect 2966 2681 2967 2685
rect 2971 2681 2972 2685
rect 2976 2682 2978 2692
rect 3158 2685 3164 2686
rect 2966 2680 2972 2681
rect 2975 2681 2981 2682
rect 2782 2678 2788 2679
rect 2926 2679 2932 2680
rect 2355 2676 2371 2678
rect 2355 2675 2356 2676
rect 2350 2674 2356 2675
rect 2926 2675 2927 2679
rect 2931 2678 2932 2679
rect 2975 2678 2976 2681
rect 2931 2677 2976 2678
rect 2980 2677 2981 2681
rect 3158 2681 3159 2685
rect 3163 2681 3164 2685
rect 3158 2680 3164 2681
rect 3190 2681 3196 2682
rect 2931 2676 2981 2677
rect 3166 2679 3173 2680
rect 2931 2675 2932 2676
rect 2926 2674 2932 2675
rect 3166 2675 3167 2679
rect 3172 2675 3173 2679
rect 3190 2677 3191 2681
rect 3195 2677 3196 2681
rect 3190 2676 3196 2677
rect 3166 2674 3173 2675
rect 1630 2670 1636 2671
rect 1542 2666 1548 2667
rect 1670 2663 1676 2664
rect 1670 2659 1671 2663
rect 1675 2659 1676 2663
rect 1670 2658 1676 2659
rect 3190 2663 3196 2664
rect 3190 2659 3191 2663
rect 3195 2659 3196 2663
rect 3190 2658 3196 2659
rect 1998 2656 2004 2657
rect 606 2653 612 2654
rect 110 2649 116 2650
rect 110 2645 111 2649
rect 115 2645 116 2649
rect 606 2649 607 2653
rect 611 2649 612 2653
rect 734 2653 740 2654
rect 606 2648 612 2649
rect 615 2651 621 2652
rect 615 2647 616 2651
rect 620 2650 621 2651
rect 630 2651 636 2652
rect 630 2650 631 2651
rect 620 2648 631 2650
rect 620 2647 621 2648
rect 615 2646 621 2647
rect 630 2647 631 2648
rect 635 2647 636 2651
rect 734 2649 735 2653
rect 739 2649 740 2653
rect 854 2653 860 2654
rect 734 2648 740 2649
rect 742 2651 749 2652
rect 630 2646 636 2647
rect 742 2647 743 2651
rect 748 2647 749 2651
rect 854 2649 855 2653
rect 859 2649 860 2653
rect 854 2648 860 2649
rect 974 2653 980 2654
rect 974 2649 975 2653
rect 979 2649 980 2653
rect 974 2648 980 2649
rect 1094 2653 1100 2654
rect 1094 2649 1095 2653
rect 1099 2649 1100 2653
rect 1094 2648 1100 2649
rect 1206 2653 1212 2654
rect 1206 2649 1207 2653
rect 1211 2649 1212 2653
rect 1206 2648 1212 2649
rect 1318 2653 1324 2654
rect 1318 2649 1319 2653
rect 1323 2649 1324 2653
rect 1438 2653 1444 2654
rect 1318 2648 1324 2649
rect 1327 2651 1333 2652
rect 742 2646 749 2647
rect 862 2647 869 2648
rect 110 2644 116 2645
rect 862 2643 863 2647
rect 868 2643 869 2647
rect 862 2642 869 2643
rect 966 2647 972 2648
rect 966 2643 967 2647
rect 971 2646 972 2647
rect 983 2647 989 2648
rect 983 2646 984 2647
rect 971 2644 984 2646
rect 971 2643 972 2644
rect 966 2642 972 2643
rect 983 2643 984 2644
rect 988 2646 989 2647
rect 1102 2647 1109 2648
rect 1102 2646 1103 2647
rect 988 2644 1103 2646
rect 988 2643 989 2644
rect 983 2642 989 2643
rect 1102 2643 1103 2644
rect 1108 2646 1109 2647
rect 1214 2647 1221 2648
rect 1214 2646 1215 2647
rect 1108 2644 1215 2646
rect 1108 2643 1109 2644
rect 1102 2642 1109 2643
rect 1214 2643 1215 2644
rect 1220 2643 1221 2647
rect 1327 2647 1328 2651
rect 1332 2650 1333 2651
rect 1342 2651 1348 2652
rect 1342 2650 1343 2651
rect 1332 2648 1343 2650
rect 1332 2647 1333 2648
rect 1327 2646 1333 2647
rect 1342 2647 1343 2648
rect 1347 2647 1348 2651
rect 1438 2649 1439 2653
rect 1443 2649 1444 2653
rect 1998 2652 1999 2656
rect 2003 2652 2004 2656
rect 1438 2648 1444 2649
rect 1446 2651 1453 2652
rect 1998 2651 2004 2652
rect 2174 2656 2180 2657
rect 2174 2652 2175 2656
rect 2179 2652 2180 2656
rect 2174 2651 2180 2652
rect 2358 2656 2364 2657
rect 2358 2652 2359 2656
rect 2363 2652 2364 2656
rect 2358 2651 2364 2652
rect 2550 2656 2556 2657
rect 2550 2652 2551 2656
rect 2555 2652 2556 2656
rect 2550 2651 2556 2652
rect 2758 2656 2764 2657
rect 2758 2652 2759 2656
rect 2763 2652 2764 2656
rect 2758 2651 2764 2652
rect 2966 2656 2972 2657
rect 2966 2652 2967 2656
rect 2971 2652 2972 2656
rect 2966 2651 2972 2652
rect 3158 2656 3164 2657
rect 3158 2652 3159 2656
rect 3163 2652 3164 2656
rect 3158 2651 3164 2652
rect 1342 2646 1348 2647
rect 1446 2647 1447 2651
rect 1452 2647 1453 2651
rect 1446 2646 1453 2647
rect 1630 2649 1636 2650
rect 1630 2645 1631 2649
rect 1635 2645 1636 2649
rect 1630 2644 1636 2645
rect 1910 2644 1916 2645
rect 1214 2642 1221 2643
rect 1910 2640 1911 2644
rect 1915 2640 1916 2644
rect 1910 2639 1916 2640
rect 2102 2644 2108 2645
rect 2102 2640 2103 2644
rect 2107 2640 2108 2644
rect 2102 2639 2108 2640
rect 2294 2644 2300 2645
rect 2294 2640 2295 2644
rect 2299 2640 2300 2644
rect 2294 2639 2300 2640
rect 2486 2644 2492 2645
rect 2486 2640 2487 2644
rect 2491 2640 2492 2644
rect 2486 2639 2492 2640
rect 2686 2644 2692 2645
rect 2686 2640 2687 2644
rect 2691 2640 2692 2644
rect 2686 2639 2692 2640
rect 1670 2637 1676 2638
rect 1670 2633 1671 2637
rect 1675 2633 1676 2637
rect 1670 2632 1676 2633
rect 3190 2637 3196 2638
rect 3190 2633 3191 2637
rect 3195 2633 3196 2637
rect 3190 2632 3196 2633
rect 110 2631 116 2632
rect 110 2627 111 2631
rect 115 2627 116 2631
rect 110 2626 116 2627
rect 1630 2631 1636 2632
rect 1630 2627 1631 2631
rect 1635 2627 1636 2631
rect 1630 2626 1636 2627
rect 606 2624 612 2625
rect 606 2620 607 2624
rect 611 2620 612 2624
rect 606 2619 612 2620
rect 734 2624 740 2625
rect 734 2620 735 2624
rect 739 2620 740 2624
rect 734 2619 740 2620
rect 854 2624 860 2625
rect 854 2620 855 2624
rect 859 2620 860 2624
rect 854 2619 860 2620
rect 974 2624 980 2625
rect 974 2620 975 2624
rect 979 2620 980 2624
rect 974 2619 980 2620
rect 1094 2624 1100 2625
rect 1094 2620 1095 2624
rect 1099 2620 1100 2624
rect 1094 2619 1100 2620
rect 1206 2624 1212 2625
rect 1206 2620 1207 2624
rect 1211 2620 1212 2624
rect 1206 2619 1212 2620
rect 1318 2624 1324 2625
rect 1318 2620 1319 2624
rect 1323 2620 1324 2624
rect 1318 2619 1324 2620
rect 1438 2624 1444 2625
rect 1438 2620 1439 2624
rect 1443 2620 1444 2624
rect 1438 2619 1444 2620
rect 1670 2619 1676 2620
rect 1670 2615 1671 2619
rect 1675 2615 1676 2619
rect 2303 2619 2309 2620
rect 1670 2614 1676 2615
rect 1910 2615 1916 2616
rect 1910 2611 1911 2615
rect 1915 2611 1916 2615
rect 1910 2610 1916 2611
rect 1918 2615 1925 2616
rect 1918 2611 1919 2615
rect 1924 2611 1925 2615
rect 1918 2610 1925 2611
rect 2102 2615 2108 2616
rect 2102 2611 2103 2615
rect 2107 2611 2108 2615
rect 2102 2610 2108 2611
rect 2111 2615 2117 2616
rect 2111 2611 2112 2615
rect 2116 2611 2117 2615
rect 2111 2610 2117 2611
rect 2294 2615 2300 2616
rect 2294 2611 2295 2615
rect 2299 2611 2300 2615
rect 2303 2615 2304 2619
rect 2308 2618 2309 2619
rect 2326 2619 2332 2620
rect 2326 2618 2327 2619
rect 2308 2616 2327 2618
rect 2308 2615 2309 2616
rect 2303 2614 2309 2615
rect 2326 2615 2327 2616
rect 2331 2618 2332 2619
rect 2350 2619 2356 2620
rect 2350 2618 2351 2619
rect 2331 2616 2351 2618
rect 2331 2615 2332 2616
rect 2326 2614 2332 2615
rect 2350 2615 2351 2616
rect 2355 2615 2356 2619
rect 2695 2619 2701 2620
rect 2350 2614 2356 2615
rect 2486 2615 2492 2616
rect 2294 2610 2300 2611
rect 2486 2611 2487 2615
rect 2491 2611 2492 2615
rect 2486 2610 2492 2611
rect 2495 2615 2501 2616
rect 2495 2611 2496 2615
rect 2500 2614 2501 2615
rect 2686 2615 2692 2616
rect 2500 2612 2682 2614
rect 2500 2611 2501 2612
rect 2495 2610 2501 2611
rect 2112 2606 2114 2610
rect 1822 2605 1828 2606
rect 1670 2601 1676 2602
rect 502 2600 508 2601
rect 502 2596 503 2600
rect 507 2596 508 2600
rect 502 2595 508 2596
rect 630 2600 636 2601
rect 630 2596 631 2600
rect 635 2596 636 2600
rect 630 2595 636 2596
rect 750 2600 756 2601
rect 750 2596 751 2600
rect 755 2596 756 2600
rect 750 2595 756 2596
rect 870 2600 876 2601
rect 870 2596 871 2600
rect 875 2596 876 2600
rect 870 2595 876 2596
rect 990 2600 996 2601
rect 990 2596 991 2600
rect 995 2596 996 2600
rect 990 2595 996 2596
rect 1102 2600 1108 2601
rect 1102 2596 1103 2600
rect 1107 2596 1108 2600
rect 1102 2595 1108 2596
rect 1214 2600 1220 2601
rect 1214 2596 1215 2600
rect 1219 2596 1220 2600
rect 1214 2595 1220 2596
rect 1334 2600 1340 2601
rect 1334 2596 1335 2600
rect 1339 2596 1340 2600
rect 1670 2597 1671 2601
rect 1675 2597 1676 2601
rect 1822 2601 1823 2605
rect 1827 2601 1828 2605
rect 1822 2600 1828 2601
rect 2014 2605 2020 2606
rect 2014 2601 2015 2605
rect 2019 2601 2020 2605
rect 2014 2600 2020 2601
rect 2064 2604 2114 2606
rect 2214 2605 2220 2606
rect 2064 2600 2066 2604
rect 2214 2601 2215 2605
rect 2219 2601 2220 2605
rect 2214 2600 2220 2601
rect 2438 2605 2444 2606
rect 2438 2601 2439 2605
rect 2443 2601 2444 2605
rect 2438 2600 2444 2601
rect 2446 2603 2453 2604
rect 1670 2596 1676 2597
rect 1830 2599 1837 2600
rect 1334 2595 1340 2596
rect 1830 2595 1831 2599
rect 1836 2595 1837 2599
rect 1830 2594 1837 2595
rect 1918 2599 1924 2600
rect 1918 2595 1919 2599
rect 1923 2598 1924 2599
rect 2006 2599 2012 2600
rect 2006 2598 2007 2599
rect 1923 2596 2007 2598
rect 1923 2595 1924 2596
rect 1918 2594 1924 2595
rect 2006 2595 2007 2596
rect 2011 2598 2012 2599
rect 2023 2599 2029 2600
rect 2023 2598 2024 2599
rect 2011 2596 2024 2598
rect 2011 2595 2012 2596
rect 2006 2594 2012 2595
rect 2023 2595 2024 2596
rect 2028 2598 2029 2599
rect 2062 2599 2068 2600
rect 2062 2598 2063 2599
rect 2028 2596 2063 2598
rect 2028 2595 2029 2596
rect 2023 2594 2029 2595
rect 2062 2595 2063 2596
rect 2067 2595 2068 2599
rect 2062 2594 2068 2595
rect 2206 2599 2212 2600
rect 2206 2595 2207 2599
rect 2211 2598 2212 2599
rect 2222 2599 2229 2600
rect 2222 2598 2223 2599
rect 2211 2596 2223 2598
rect 2211 2595 2212 2596
rect 2206 2594 2212 2595
rect 2222 2595 2223 2596
rect 2228 2595 2229 2599
rect 2446 2599 2447 2603
rect 2452 2602 2453 2603
rect 2496 2602 2498 2610
rect 2452 2600 2498 2602
rect 2670 2605 2676 2606
rect 2670 2601 2671 2605
rect 2675 2601 2676 2605
rect 2680 2604 2682 2612
rect 2686 2611 2687 2615
rect 2691 2611 2692 2615
rect 2695 2615 2696 2619
rect 2700 2618 2701 2619
rect 2782 2619 2788 2620
rect 2782 2618 2783 2619
rect 2700 2616 2783 2618
rect 2700 2615 2701 2616
rect 2695 2614 2701 2615
rect 2782 2615 2783 2616
rect 2787 2615 2788 2619
rect 2782 2614 2788 2615
rect 3190 2619 3196 2620
rect 3190 2615 3191 2619
rect 3195 2615 3196 2619
rect 3190 2614 3196 2615
rect 2686 2610 2692 2611
rect 2670 2600 2676 2601
rect 2679 2603 2685 2604
rect 2452 2599 2453 2600
rect 2446 2598 2453 2599
rect 2679 2599 2680 2603
rect 2684 2602 2685 2603
rect 2696 2602 2698 2614
rect 2684 2600 2698 2602
rect 2918 2605 2924 2606
rect 2918 2601 2919 2605
rect 2923 2601 2924 2605
rect 2918 2600 2924 2601
rect 3158 2605 3164 2606
rect 3158 2601 3159 2605
rect 3163 2601 3164 2605
rect 3158 2600 3164 2601
rect 3190 2601 3196 2602
rect 2684 2599 2685 2600
rect 2679 2598 2685 2599
rect 2926 2599 2933 2600
rect 2222 2594 2229 2595
rect 2926 2595 2927 2599
rect 2932 2595 2933 2599
rect 2926 2594 2933 2595
rect 3142 2599 3148 2600
rect 3142 2595 3143 2599
rect 3147 2598 3148 2599
rect 3166 2599 3173 2600
rect 3166 2598 3167 2599
rect 3147 2596 3167 2598
rect 3147 2595 3148 2596
rect 3142 2594 3148 2595
rect 3166 2595 3167 2596
rect 3172 2595 3173 2599
rect 3190 2597 3191 2601
rect 3195 2597 3196 2601
rect 3190 2596 3196 2597
rect 3166 2594 3173 2595
rect 110 2593 116 2594
rect 110 2589 111 2593
rect 115 2589 116 2593
rect 110 2588 116 2589
rect 1630 2593 1636 2594
rect 1630 2589 1631 2593
rect 1635 2589 1636 2593
rect 1630 2588 1636 2589
rect 1670 2583 1676 2584
rect 862 2579 868 2580
rect 110 2575 116 2576
rect 110 2571 111 2575
rect 115 2571 116 2575
rect 862 2575 863 2579
rect 867 2578 868 2579
rect 902 2579 908 2580
rect 902 2578 903 2579
rect 867 2576 903 2578
rect 867 2575 868 2576
rect 862 2574 868 2575
rect 879 2575 885 2576
rect 110 2570 116 2571
rect 502 2571 508 2572
rect 502 2567 503 2571
rect 507 2567 508 2571
rect 502 2566 508 2567
rect 510 2571 517 2572
rect 510 2567 511 2571
rect 516 2567 517 2571
rect 510 2566 517 2567
rect 630 2571 636 2572
rect 630 2567 631 2571
rect 635 2567 636 2571
rect 630 2566 636 2567
rect 638 2571 645 2572
rect 638 2567 639 2571
rect 644 2567 645 2571
rect 638 2566 645 2567
rect 750 2571 756 2572
rect 750 2567 751 2571
rect 755 2567 756 2571
rect 750 2566 756 2567
rect 759 2571 765 2572
rect 759 2567 760 2571
rect 764 2570 765 2571
rect 782 2571 788 2572
rect 782 2570 783 2571
rect 764 2568 783 2570
rect 764 2567 765 2568
rect 759 2566 765 2567
rect 782 2567 783 2568
rect 787 2567 788 2571
rect 782 2566 788 2567
rect 870 2571 876 2572
rect 870 2567 871 2571
rect 875 2567 876 2571
rect 879 2571 880 2575
rect 884 2571 885 2575
rect 902 2575 903 2576
rect 907 2578 908 2579
rect 1670 2579 1671 2583
rect 1675 2579 1676 2583
rect 1670 2578 1676 2579
rect 3190 2583 3196 2584
rect 3190 2579 3191 2583
rect 3195 2579 3196 2583
rect 3190 2578 3196 2579
rect 907 2576 1002 2578
rect 1280 2576 1346 2578
rect 1822 2576 1828 2577
rect 907 2575 908 2576
rect 902 2574 908 2575
rect 999 2575 1005 2576
rect 879 2570 885 2571
rect 990 2571 996 2572
rect 870 2566 876 2567
rect 990 2567 991 2571
rect 995 2567 996 2571
rect 999 2571 1000 2575
rect 1004 2574 1005 2575
rect 1014 2575 1020 2576
rect 1014 2574 1015 2575
rect 1004 2572 1015 2574
rect 1004 2571 1005 2572
rect 999 2570 1005 2571
rect 1014 2571 1015 2572
rect 1019 2571 1020 2575
rect 1222 2575 1229 2576
rect 1014 2570 1020 2571
rect 1102 2571 1108 2572
rect 990 2566 996 2567
rect 1102 2567 1103 2571
rect 1107 2567 1108 2571
rect 1102 2566 1108 2567
rect 1111 2571 1117 2572
rect 1111 2567 1112 2571
rect 1116 2570 1117 2571
rect 1126 2571 1132 2572
rect 1126 2570 1127 2571
rect 1116 2568 1127 2570
rect 1116 2567 1117 2568
rect 1111 2566 1117 2567
rect 1126 2567 1127 2568
rect 1131 2567 1132 2571
rect 1126 2566 1132 2567
rect 1214 2571 1220 2572
rect 1214 2567 1215 2571
rect 1219 2567 1220 2571
rect 1222 2571 1223 2575
rect 1228 2574 1229 2575
rect 1246 2575 1252 2576
rect 1246 2574 1247 2575
rect 1228 2572 1247 2574
rect 1228 2571 1229 2572
rect 1222 2570 1229 2571
rect 1246 2571 1247 2572
rect 1251 2574 1252 2575
rect 1280 2574 1282 2576
rect 1251 2572 1282 2574
rect 1342 2575 1349 2576
rect 1251 2571 1252 2572
rect 1246 2570 1252 2571
rect 1334 2571 1340 2572
rect 1214 2566 1220 2567
rect 1334 2567 1335 2571
rect 1339 2567 1340 2571
rect 1342 2571 1343 2575
rect 1348 2571 1349 2575
rect 1342 2570 1349 2571
rect 1630 2575 1636 2576
rect 1630 2571 1631 2575
rect 1635 2571 1636 2575
rect 1822 2572 1823 2576
rect 1827 2572 1828 2576
rect 1822 2571 1828 2572
rect 2014 2576 2020 2577
rect 2014 2572 2015 2576
rect 2019 2572 2020 2576
rect 2014 2571 2020 2572
rect 2214 2576 2220 2577
rect 2214 2572 2215 2576
rect 2219 2572 2220 2576
rect 2214 2571 2220 2572
rect 2438 2576 2444 2577
rect 2438 2572 2439 2576
rect 2443 2572 2444 2576
rect 2438 2571 2444 2572
rect 2670 2576 2676 2577
rect 2670 2572 2671 2576
rect 2675 2572 2676 2576
rect 2670 2571 2676 2572
rect 2918 2576 2924 2577
rect 2918 2572 2919 2576
rect 2923 2572 2924 2576
rect 2918 2571 2924 2572
rect 3158 2576 3164 2577
rect 3158 2572 3159 2576
rect 3163 2572 3164 2576
rect 3158 2571 3164 2572
rect 1630 2570 1636 2571
rect 1334 2566 1340 2567
rect 1734 2560 1740 2561
rect 1734 2556 1735 2560
rect 1739 2556 1740 2560
rect 1734 2555 1740 2556
rect 1894 2560 1900 2561
rect 1894 2556 1895 2560
rect 1899 2556 1900 2560
rect 1894 2555 1900 2556
rect 2054 2560 2060 2561
rect 2054 2556 2055 2560
rect 2059 2556 2060 2560
rect 2054 2555 2060 2556
rect 2214 2560 2220 2561
rect 2214 2556 2215 2560
rect 2219 2556 2220 2560
rect 2214 2555 2220 2556
rect 2374 2560 2380 2561
rect 2374 2556 2375 2560
rect 2379 2556 2380 2560
rect 2374 2555 2380 2556
rect 2534 2560 2540 2561
rect 2534 2556 2535 2560
rect 2539 2556 2540 2560
rect 2534 2555 2540 2556
rect 1670 2553 1676 2554
rect 398 2549 404 2550
rect 110 2545 116 2546
rect 110 2541 111 2545
rect 115 2541 116 2545
rect 398 2545 399 2549
rect 403 2545 404 2549
rect 398 2544 404 2545
rect 526 2549 532 2550
rect 526 2545 527 2549
rect 531 2545 532 2549
rect 526 2544 532 2545
rect 654 2549 660 2550
rect 654 2545 655 2549
rect 659 2545 660 2549
rect 654 2544 660 2545
rect 774 2549 780 2550
rect 774 2545 775 2549
rect 779 2545 780 2549
rect 894 2549 900 2550
rect 774 2544 780 2545
rect 782 2547 789 2548
rect 110 2540 116 2541
rect 407 2543 413 2544
rect 407 2539 408 2543
rect 412 2542 413 2543
rect 442 2543 448 2544
rect 442 2542 443 2543
rect 412 2540 443 2542
rect 412 2539 413 2540
rect 407 2538 413 2539
rect 442 2539 443 2540
rect 447 2542 448 2543
rect 510 2543 516 2544
rect 510 2542 511 2543
rect 447 2540 511 2542
rect 447 2539 448 2540
rect 442 2538 448 2539
rect 510 2539 511 2540
rect 515 2542 516 2543
rect 535 2543 541 2544
rect 535 2542 536 2543
rect 515 2540 536 2542
rect 515 2539 516 2540
rect 510 2538 516 2539
rect 535 2539 536 2540
rect 540 2542 541 2543
rect 638 2543 644 2544
rect 638 2542 639 2543
rect 540 2540 639 2542
rect 540 2539 541 2540
rect 535 2538 541 2539
rect 638 2539 639 2540
rect 643 2542 644 2543
rect 663 2543 669 2544
rect 663 2542 664 2543
rect 643 2540 664 2542
rect 643 2539 644 2540
rect 638 2538 644 2539
rect 663 2539 664 2540
rect 668 2539 669 2543
rect 782 2543 783 2547
rect 788 2546 789 2547
rect 862 2547 868 2548
rect 862 2546 863 2547
rect 788 2544 863 2546
rect 788 2543 789 2544
rect 782 2542 789 2543
rect 862 2543 863 2544
rect 867 2543 868 2547
rect 894 2545 895 2549
rect 899 2545 900 2549
rect 1006 2549 1012 2550
rect 894 2544 900 2545
rect 902 2547 909 2548
rect 862 2542 868 2543
rect 902 2543 903 2547
rect 908 2543 909 2547
rect 1006 2545 1007 2549
rect 1011 2545 1012 2549
rect 1118 2549 1124 2550
rect 1006 2544 1012 2545
rect 1014 2547 1021 2548
rect 902 2542 909 2543
rect 1014 2543 1015 2547
rect 1020 2546 1021 2547
rect 1020 2544 1041 2546
rect 1118 2545 1119 2549
rect 1123 2545 1124 2549
rect 1118 2544 1124 2545
rect 1238 2549 1244 2550
rect 1238 2545 1239 2549
rect 1243 2545 1244 2549
rect 1670 2549 1671 2553
rect 1675 2549 1676 2553
rect 1670 2548 1676 2549
rect 3190 2553 3196 2554
rect 3190 2549 3191 2553
rect 3195 2549 3196 2553
rect 3190 2548 3196 2549
rect 1238 2544 1244 2545
rect 1246 2547 1253 2548
rect 1020 2543 1021 2544
rect 1014 2542 1021 2543
rect 1039 2542 1041 2544
rect 1126 2543 1133 2544
rect 1126 2542 1127 2543
rect 1039 2540 1127 2542
rect 663 2538 669 2539
rect 1126 2539 1127 2540
rect 1132 2542 1133 2543
rect 1246 2543 1247 2547
rect 1252 2543 1253 2547
rect 1246 2542 1253 2543
rect 1630 2545 1636 2546
rect 1132 2540 1250 2542
rect 1630 2541 1631 2545
rect 1635 2541 1636 2545
rect 1630 2540 1636 2541
rect 1132 2539 1133 2540
rect 1126 2538 1133 2539
rect 1670 2535 1676 2536
rect 1670 2531 1671 2535
rect 1675 2531 1676 2535
rect 2062 2535 2069 2536
rect 1670 2530 1676 2531
rect 1734 2531 1740 2532
rect 110 2527 116 2528
rect 110 2523 111 2527
rect 115 2523 116 2527
rect 110 2522 116 2523
rect 1630 2527 1636 2528
rect 1630 2523 1631 2527
rect 1635 2523 1636 2527
rect 1734 2527 1735 2531
rect 1739 2527 1740 2531
rect 1734 2526 1740 2527
rect 1743 2531 1749 2532
rect 1743 2527 1744 2531
rect 1748 2527 1749 2531
rect 1743 2526 1749 2527
rect 1894 2531 1900 2532
rect 1894 2527 1895 2531
rect 1899 2527 1900 2531
rect 1894 2526 1900 2527
rect 1902 2531 1909 2532
rect 1902 2527 1903 2531
rect 1908 2530 1909 2531
rect 1918 2531 1924 2532
rect 1918 2530 1919 2531
rect 1908 2528 1919 2530
rect 1908 2527 1909 2528
rect 1902 2526 1909 2527
rect 1918 2527 1919 2528
rect 1923 2527 1924 2531
rect 1918 2526 1924 2527
rect 2054 2531 2060 2532
rect 2054 2527 2055 2531
rect 2059 2527 2060 2531
rect 2062 2531 2063 2535
rect 2068 2531 2069 2535
rect 2222 2535 2229 2536
rect 2062 2530 2069 2531
rect 2214 2531 2220 2532
rect 2054 2526 2060 2527
rect 2214 2527 2215 2531
rect 2219 2527 2220 2531
rect 2222 2531 2223 2535
rect 2228 2531 2229 2535
rect 3190 2535 3196 2536
rect 2222 2530 2229 2531
rect 2374 2531 2380 2532
rect 2214 2526 2220 2527
rect 2374 2527 2375 2531
rect 2379 2527 2380 2531
rect 2374 2526 2380 2527
rect 2383 2531 2389 2532
rect 2383 2527 2384 2531
rect 2388 2527 2389 2531
rect 2383 2526 2389 2527
rect 2534 2531 2540 2532
rect 2534 2527 2535 2531
rect 2539 2527 2540 2531
rect 2534 2526 2540 2527
rect 2543 2531 2549 2532
rect 2543 2527 2544 2531
rect 2548 2527 2549 2531
rect 3190 2531 3191 2535
rect 3195 2531 3196 2535
rect 3190 2530 3196 2531
rect 2543 2526 2549 2527
rect 1630 2522 1636 2523
rect 398 2520 404 2521
rect 398 2516 399 2520
rect 403 2516 404 2520
rect 398 2515 404 2516
rect 526 2520 532 2521
rect 526 2516 527 2520
rect 531 2516 532 2520
rect 526 2515 532 2516
rect 654 2520 660 2521
rect 654 2516 655 2520
rect 659 2516 660 2520
rect 654 2515 660 2516
rect 774 2520 780 2521
rect 774 2516 775 2520
rect 779 2516 780 2520
rect 774 2515 780 2516
rect 894 2520 900 2521
rect 894 2516 895 2520
rect 899 2516 900 2520
rect 894 2515 900 2516
rect 1006 2520 1012 2521
rect 1006 2516 1007 2520
rect 1011 2516 1012 2520
rect 1006 2515 1012 2516
rect 1118 2520 1124 2521
rect 1118 2516 1119 2520
rect 1123 2516 1124 2520
rect 1118 2515 1124 2516
rect 1238 2520 1244 2521
rect 1238 2516 1239 2520
rect 1243 2516 1244 2520
rect 1238 2515 1244 2516
rect 1694 2517 1700 2518
rect 1670 2513 1676 2514
rect 1670 2509 1671 2513
rect 1675 2509 1676 2513
rect 1694 2513 1695 2517
rect 1699 2513 1700 2517
rect 1694 2512 1700 2513
rect 1703 2515 1709 2516
rect 1703 2511 1704 2515
rect 1708 2514 1709 2515
rect 1744 2514 1746 2526
rect 2384 2522 2386 2526
rect 2544 2522 2546 2526
rect 2574 2523 2580 2524
rect 2574 2522 2575 2523
rect 2359 2520 2575 2522
rect 1708 2512 1746 2514
rect 1862 2517 1868 2518
rect 1862 2513 1863 2517
rect 1867 2513 1868 2517
rect 1862 2512 1868 2513
rect 2078 2517 2084 2518
rect 2078 2513 2079 2517
rect 2083 2513 2084 2517
rect 2078 2512 2084 2513
rect 2318 2517 2324 2518
rect 2318 2513 2319 2517
rect 2323 2513 2324 2517
rect 2318 2512 2324 2513
rect 2326 2515 2333 2516
rect 1708 2511 1709 2512
rect 1703 2510 1709 2511
rect 1744 2510 1746 2512
rect 1830 2511 1836 2512
rect 1830 2510 1831 2511
rect 1670 2508 1676 2509
rect 1744 2508 1831 2510
rect 1830 2507 1831 2508
rect 1835 2510 1836 2511
rect 1871 2511 1877 2512
rect 1871 2510 1872 2511
rect 1835 2508 1872 2510
rect 1835 2507 1836 2508
rect 1830 2506 1836 2507
rect 1871 2507 1872 2508
rect 1876 2510 1877 2511
rect 1902 2511 1908 2512
rect 1902 2510 1903 2511
rect 1876 2508 1903 2510
rect 1876 2507 1877 2508
rect 1871 2506 1877 2507
rect 1902 2507 1903 2508
rect 1907 2507 1908 2511
rect 1902 2506 1908 2507
rect 2062 2511 2068 2512
rect 2062 2507 2063 2511
rect 2067 2510 2068 2511
rect 2087 2511 2093 2512
rect 2087 2510 2088 2511
rect 2067 2508 2088 2510
rect 2067 2507 2068 2508
rect 2062 2506 2068 2507
rect 2087 2507 2088 2508
rect 2092 2507 2093 2511
rect 2326 2511 2327 2515
rect 2332 2514 2333 2515
rect 2359 2514 2361 2520
rect 2574 2519 2575 2520
rect 2579 2522 2580 2523
rect 2579 2520 2594 2522
rect 2579 2519 2580 2520
rect 2574 2518 2580 2519
rect 2332 2512 2361 2514
rect 2582 2517 2588 2518
rect 2582 2513 2583 2517
rect 2587 2513 2588 2517
rect 2592 2516 2594 2520
rect 2854 2517 2860 2518
rect 2582 2512 2588 2513
rect 2591 2515 2597 2516
rect 2332 2511 2333 2512
rect 2326 2510 2333 2511
rect 2591 2511 2592 2515
rect 2596 2511 2597 2515
rect 2854 2513 2855 2517
rect 2859 2513 2860 2517
rect 2854 2512 2860 2513
rect 3134 2517 3140 2518
rect 3134 2513 3135 2517
rect 3139 2513 3140 2517
rect 3134 2512 3140 2513
rect 3190 2513 3196 2514
rect 2591 2510 2597 2511
rect 2862 2511 2869 2512
rect 2087 2506 2093 2507
rect 2862 2507 2863 2511
rect 2868 2510 2869 2511
rect 2926 2511 2932 2512
rect 2926 2510 2927 2511
rect 2868 2508 2927 2510
rect 2868 2507 2869 2508
rect 2862 2506 2869 2507
rect 2926 2507 2927 2508
rect 2931 2510 2932 2511
rect 2974 2511 2980 2512
rect 2974 2510 2975 2511
rect 2931 2508 2975 2510
rect 2931 2507 2932 2508
rect 2926 2506 2932 2507
rect 2974 2507 2975 2508
rect 2979 2507 2980 2511
rect 2974 2506 2980 2507
rect 3142 2511 3149 2512
rect 3142 2507 3143 2511
rect 3148 2507 3149 2511
rect 3190 2509 3191 2513
rect 3195 2509 3196 2513
rect 3190 2508 3196 2509
rect 3142 2506 3149 2507
rect 302 2496 308 2497
rect 302 2492 303 2496
rect 307 2492 308 2496
rect 302 2491 308 2492
rect 430 2496 436 2497
rect 430 2492 431 2496
rect 435 2492 436 2496
rect 430 2491 436 2492
rect 558 2496 564 2497
rect 558 2492 559 2496
rect 563 2492 564 2496
rect 558 2491 564 2492
rect 702 2496 708 2497
rect 702 2492 703 2496
rect 707 2492 708 2496
rect 702 2491 708 2492
rect 862 2496 868 2497
rect 862 2492 863 2496
rect 867 2492 868 2496
rect 862 2491 868 2492
rect 1038 2496 1044 2497
rect 1038 2492 1039 2496
rect 1043 2492 1044 2496
rect 1038 2491 1044 2492
rect 1222 2496 1228 2497
rect 1222 2492 1223 2496
rect 1227 2492 1228 2496
rect 1222 2491 1228 2492
rect 1422 2496 1428 2497
rect 1422 2492 1423 2496
rect 1427 2492 1428 2496
rect 1422 2491 1428 2492
rect 1598 2496 1604 2497
rect 1598 2492 1599 2496
rect 1603 2492 1604 2496
rect 1598 2491 1604 2492
rect 1670 2495 1676 2496
rect 1670 2491 1671 2495
rect 1675 2491 1676 2495
rect 1670 2490 1676 2491
rect 3190 2495 3196 2496
rect 3190 2491 3191 2495
rect 3195 2491 3196 2495
rect 3190 2490 3196 2491
rect 110 2489 116 2490
rect 110 2485 111 2489
rect 115 2485 116 2489
rect 110 2484 116 2485
rect 1630 2489 1636 2490
rect 1630 2485 1631 2489
rect 1635 2485 1636 2489
rect 1630 2484 1636 2485
rect 1694 2488 1700 2489
rect 1694 2484 1695 2488
rect 1699 2484 1700 2488
rect 1694 2483 1700 2484
rect 1862 2488 1868 2489
rect 1862 2484 1863 2488
rect 1867 2484 1868 2488
rect 1862 2483 1868 2484
rect 2078 2488 2084 2489
rect 2078 2484 2079 2488
rect 2083 2484 2084 2488
rect 2078 2483 2084 2484
rect 2318 2488 2324 2489
rect 2318 2484 2319 2488
rect 2323 2484 2324 2488
rect 2318 2483 2324 2484
rect 2582 2488 2588 2489
rect 2582 2484 2583 2488
rect 2587 2484 2588 2488
rect 2582 2483 2588 2484
rect 2854 2488 2860 2489
rect 2854 2484 2855 2488
rect 2859 2484 2860 2488
rect 2854 2483 2860 2484
rect 3134 2488 3140 2489
rect 3134 2484 3135 2488
rect 3139 2484 3140 2488
rect 3134 2483 3140 2484
rect 1382 2475 1388 2476
rect 1382 2474 1383 2475
rect 1248 2472 1383 2474
rect 110 2471 116 2472
rect 110 2467 111 2471
rect 115 2467 116 2471
rect 871 2471 877 2472
rect 110 2466 116 2467
rect 302 2467 308 2468
rect 302 2463 303 2467
rect 307 2463 308 2467
rect 302 2462 308 2463
rect 310 2467 317 2468
rect 310 2463 311 2467
rect 316 2463 317 2467
rect 310 2462 317 2463
rect 430 2467 436 2468
rect 430 2463 431 2467
rect 435 2463 436 2467
rect 430 2462 436 2463
rect 438 2467 445 2468
rect 438 2463 439 2467
rect 444 2463 445 2467
rect 438 2462 445 2463
rect 558 2467 564 2468
rect 558 2463 559 2467
rect 563 2463 564 2467
rect 558 2462 564 2463
rect 567 2467 573 2468
rect 567 2463 568 2467
rect 572 2466 573 2467
rect 610 2467 616 2468
rect 610 2466 611 2467
rect 572 2464 611 2466
rect 572 2463 573 2464
rect 567 2462 573 2463
rect 610 2463 611 2464
rect 615 2463 616 2467
rect 610 2462 616 2463
rect 702 2467 708 2468
rect 702 2463 703 2467
rect 707 2463 708 2467
rect 702 2462 708 2463
rect 711 2467 717 2468
rect 711 2463 712 2467
rect 716 2466 717 2467
rect 774 2467 780 2468
rect 774 2466 775 2467
rect 716 2464 775 2466
rect 716 2463 717 2464
rect 711 2462 717 2463
rect 774 2463 775 2464
rect 779 2463 780 2467
rect 774 2462 780 2463
rect 862 2467 868 2468
rect 862 2463 863 2467
rect 867 2463 868 2467
rect 871 2467 872 2471
rect 876 2470 877 2471
rect 902 2471 908 2472
rect 902 2470 903 2471
rect 876 2468 903 2470
rect 876 2467 877 2468
rect 871 2466 877 2467
rect 902 2467 903 2468
rect 907 2467 908 2471
rect 1046 2471 1053 2472
rect 902 2466 908 2467
rect 1038 2467 1044 2468
rect 862 2462 868 2463
rect 1038 2463 1039 2467
rect 1043 2463 1044 2467
rect 1046 2467 1047 2471
rect 1052 2470 1053 2471
rect 1126 2471 1132 2472
rect 1126 2470 1127 2471
rect 1052 2468 1127 2470
rect 1052 2467 1053 2468
rect 1046 2466 1053 2467
rect 1126 2467 1127 2468
rect 1131 2467 1132 2471
rect 1248 2468 1250 2472
rect 1382 2471 1383 2472
rect 1387 2474 1388 2475
rect 1574 2475 1580 2476
rect 1574 2474 1575 2475
rect 1387 2472 1575 2474
rect 1387 2471 1388 2472
rect 1382 2470 1388 2471
rect 1431 2471 1437 2472
rect 1126 2466 1132 2467
rect 1222 2467 1228 2468
rect 1038 2462 1044 2463
rect 1222 2463 1223 2467
rect 1227 2463 1228 2467
rect 1222 2462 1228 2463
rect 1231 2467 1237 2468
rect 1231 2463 1232 2467
rect 1236 2466 1237 2467
rect 1246 2467 1252 2468
rect 1246 2466 1247 2467
rect 1236 2464 1247 2466
rect 1236 2463 1237 2464
rect 1231 2462 1237 2463
rect 1246 2463 1247 2464
rect 1251 2463 1252 2467
rect 1246 2462 1252 2463
rect 1422 2467 1428 2468
rect 1422 2463 1423 2467
rect 1427 2463 1428 2467
rect 1431 2467 1432 2471
rect 1436 2467 1437 2471
rect 1574 2471 1575 2472
rect 1579 2474 1580 2475
rect 1579 2472 1610 2474
rect 1579 2471 1580 2472
rect 1574 2470 1580 2471
rect 1607 2471 1613 2472
rect 1431 2466 1437 2467
rect 1598 2467 1604 2468
rect 1422 2462 1428 2463
rect 1598 2463 1599 2467
rect 1603 2463 1604 2467
rect 1607 2467 1608 2471
rect 1612 2467 1613 2471
rect 1607 2466 1613 2467
rect 1630 2471 1636 2472
rect 1630 2467 1631 2471
rect 1635 2467 1636 2471
rect 1630 2466 1636 2467
rect 2318 2468 2324 2469
rect 1598 2462 1604 2463
rect 1608 2454 1610 2466
rect 2318 2464 2319 2468
rect 2323 2464 2324 2468
rect 2318 2463 2324 2464
rect 2566 2468 2572 2469
rect 2566 2464 2567 2468
rect 2571 2464 2572 2468
rect 2566 2463 2572 2464
rect 2822 2468 2828 2469
rect 2822 2464 2823 2468
rect 2827 2464 2828 2468
rect 2822 2463 2828 2464
rect 3078 2468 3084 2469
rect 3078 2464 3079 2468
rect 3083 2464 3084 2468
rect 3078 2463 3084 2464
rect 1670 2461 1676 2462
rect 1670 2457 1671 2461
rect 1675 2457 1676 2461
rect 1670 2456 1676 2457
rect 3190 2461 3196 2462
rect 3190 2457 3191 2461
rect 3195 2457 3196 2461
rect 3190 2456 3196 2457
rect 198 2453 204 2454
rect 110 2449 116 2450
rect 110 2445 111 2449
rect 115 2445 116 2449
rect 198 2449 199 2453
rect 203 2449 204 2453
rect 198 2448 204 2449
rect 326 2453 332 2454
rect 326 2449 327 2453
rect 331 2449 332 2453
rect 326 2448 332 2449
rect 454 2453 460 2454
rect 454 2449 455 2453
rect 459 2449 460 2453
rect 454 2448 460 2449
rect 598 2453 604 2454
rect 598 2449 599 2453
rect 603 2449 604 2453
rect 598 2448 604 2449
rect 766 2453 772 2454
rect 766 2449 767 2453
rect 771 2449 772 2453
rect 766 2448 772 2449
rect 950 2453 956 2454
rect 950 2449 951 2453
rect 955 2449 956 2453
rect 1158 2453 1164 2454
rect 950 2448 956 2449
rect 959 2451 965 2452
rect 110 2444 116 2445
rect 207 2447 213 2448
rect 207 2443 208 2447
rect 212 2446 213 2447
rect 246 2447 252 2448
rect 246 2446 247 2447
rect 212 2444 247 2446
rect 212 2443 213 2444
rect 207 2442 213 2443
rect 246 2443 247 2444
rect 251 2446 252 2447
rect 310 2447 316 2448
rect 310 2446 311 2447
rect 251 2444 311 2446
rect 251 2443 252 2444
rect 246 2442 252 2443
rect 310 2443 311 2444
rect 315 2446 316 2447
rect 335 2447 341 2448
rect 335 2446 336 2447
rect 315 2444 336 2446
rect 315 2443 316 2444
rect 310 2442 316 2443
rect 335 2443 336 2444
rect 340 2446 341 2447
rect 438 2447 444 2448
rect 438 2446 439 2447
rect 340 2444 439 2446
rect 340 2443 341 2444
rect 335 2442 341 2443
rect 438 2443 439 2444
rect 443 2446 444 2447
rect 463 2447 469 2448
rect 463 2446 464 2447
rect 443 2444 464 2446
rect 443 2443 444 2444
rect 438 2442 444 2443
rect 463 2443 464 2444
rect 468 2443 469 2447
rect 463 2442 469 2443
rect 607 2447 616 2448
rect 607 2443 608 2447
rect 615 2443 616 2447
rect 607 2442 616 2443
rect 774 2447 781 2448
rect 774 2443 775 2447
rect 780 2443 781 2447
rect 959 2447 960 2451
rect 964 2450 965 2451
rect 1046 2451 1052 2452
rect 1046 2450 1047 2451
rect 964 2448 1047 2450
rect 964 2447 965 2448
rect 959 2446 965 2447
rect 1046 2447 1047 2448
rect 1051 2447 1052 2451
rect 1158 2449 1159 2453
rect 1163 2449 1164 2453
rect 1374 2453 1380 2454
rect 1158 2448 1164 2449
rect 1167 2451 1173 2452
rect 1046 2446 1052 2447
rect 1167 2447 1168 2451
rect 1172 2450 1173 2451
rect 1182 2451 1188 2452
rect 1182 2450 1183 2451
rect 1172 2448 1183 2450
rect 1172 2447 1173 2448
rect 1167 2446 1173 2447
rect 1182 2447 1183 2448
rect 1187 2450 1188 2451
rect 1246 2451 1252 2452
rect 1246 2450 1247 2451
rect 1187 2448 1247 2450
rect 1187 2447 1188 2448
rect 1182 2446 1188 2447
rect 1246 2447 1247 2448
rect 1251 2447 1252 2451
rect 1374 2449 1375 2453
rect 1379 2449 1380 2453
rect 1590 2453 1596 2454
rect 1374 2448 1380 2449
rect 1382 2451 1389 2452
rect 1246 2446 1252 2447
rect 1382 2447 1383 2451
rect 1388 2447 1389 2451
rect 1590 2449 1591 2453
rect 1595 2449 1596 2453
rect 1590 2448 1596 2449
rect 1599 2453 1610 2454
rect 1599 2449 1600 2453
rect 1604 2452 1610 2453
rect 1604 2449 1605 2452
rect 1599 2448 1605 2449
rect 1630 2449 1636 2450
rect 1382 2446 1389 2447
rect 1630 2445 1631 2449
rect 1635 2445 1636 2449
rect 1630 2444 1636 2445
rect 774 2442 781 2443
rect 1670 2443 1676 2444
rect 1670 2439 1671 2443
rect 1675 2439 1676 2443
rect 2326 2443 2333 2444
rect 1670 2438 1676 2439
rect 2318 2439 2324 2440
rect 2318 2435 2319 2439
rect 2323 2435 2324 2439
rect 2326 2439 2327 2443
rect 2332 2439 2333 2443
rect 2574 2443 2581 2444
rect 2326 2438 2333 2439
rect 2566 2439 2572 2440
rect 2318 2434 2324 2435
rect 2566 2435 2567 2439
rect 2571 2435 2572 2439
rect 2574 2439 2575 2443
rect 2580 2439 2581 2443
rect 2831 2443 2837 2444
rect 2574 2438 2581 2439
rect 2822 2439 2828 2440
rect 2566 2434 2572 2435
rect 2822 2435 2823 2439
rect 2827 2435 2828 2439
rect 2831 2439 2832 2443
rect 2836 2442 2837 2443
rect 2862 2443 2868 2444
rect 2862 2442 2863 2443
rect 2836 2440 2863 2442
rect 2836 2439 2837 2440
rect 2831 2438 2837 2439
rect 2862 2439 2863 2440
rect 2867 2439 2868 2443
rect 3190 2443 3196 2444
rect 2862 2438 2868 2439
rect 3078 2439 3084 2440
rect 2822 2434 2828 2435
rect 110 2431 116 2432
rect 110 2427 111 2431
rect 115 2427 116 2431
rect 110 2426 116 2427
rect 1630 2431 1636 2432
rect 1630 2427 1631 2431
rect 1635 2427 1636 2431
rect 1630 2426 1636 2427
rect 2230 2429 2236 2430
rect 1670 2425 1676 2426
rect 198 2424 204 2425
rect 198 2420 199 2424
rect 203 2420 204 2424
rect 198 2419 204 2420
rect 326 2424 332 2425
rect 326 2420 327 2424
rect 331 2420 332 2424
rect 326 2419 332 2420
rect 454 2424 460 2425
rect 454 2420 455 2424
rect 459 2420 460 2424
rect 454 2419 460 2420
rect 598 2424 604 2425
rect 598 2420 599 2424
rect 603 2420 604 2424
rect 598 2419 604 2420
rect 766 2424 772 2425
rect 766 2420 767 2424
rect 771 2420 772 2424
rect 766 2419 772 2420
rect 950 2424 956 2425
rect 950 2420 951 2424
rect 955 2420 956 2424
rect 950 2419 956 2420
rect 1158 2424 1164 2425
rect 1158 2420 1159 2424
rect 1163 2420 1164 2424
rect 1158 2419 1164 2420
rect 1374 2424 1380 2425
rect 1374 2420 1375 2424
rect 1379 2420 1380 2424
rect 1374 2419 1380 2420
rect 1590 2424 1596 2425
rect 1590 2420 1591 2424
rect 1595 2420 1596 2424
rect 1670 2421 1671 2425
rect 1675 2421 1676 2425
rect 2230 2425 2231 2429
rect 2235 2425 2236 2429
rect 2390 2429 2396 2430
rect 2230 2424 2236 2425
rect 2238 2427 2245 2428
rect 2238 2423 2239 2427
rect 2244 2426 2245 2427
rect 2326 2427 2332 2428
rect 2326 2426 2327 2427
rect 2244 2424 2327 2426
rect 2244 2423 2245 2424
rect 2238 2422 2245 2423
rect 2326 2423 2327 2424
rect 2331 2426 2332 2427
rect 2342 2427 2348 2428
rect 2342 2426 2343 2427
rect 2331 2424 2343 2426
rect 2331 2423 2332 2424
rect 2326 2422 2332 2423
rect 2342 2423 2343 2424
rect 2347 2426 2348 2427
rect 2347 2424 2361 2426
rect 2390 2425 2391 2429
rect 2395 2425 2396 2429
rect 2390 2424 2396 2425
rect 2542 2429 2548 2430
rect 2542 2425 2543 2429
rect 2547 2425 2548 2429
rect 2686 2429 2692 2430
rect 2542 2424 2548 2425
rect 2551 2427 2557 2428
rect 2347 2423 2348 2424
rect 2342 2422 2348 2423
rect 2359 2422 2361 2424
rect 2399 2423 2405 2424
rect 2399 2422 2400 2423
rect 1670 2420 1676 2421
rect 2359 2420 2400 2422
rect 1590 2419 1596 2420
rect 2399 2419 2400 2420
rect 2404 2419 2405 2423
rect 2551 2423 2552 2427
rect 2556 2426 2557 2427
rect 2574 2427 2580 2428
rect 2574 2426 2575 2427
rect 2556 2424 2575 2426
rect 2556 2423 2557 2424
rect 2551 2422 2557 2423
rect 2574 2423 2575 2424
rect 2579 2423 2580 2427
rect 2686 2425 2687 2429
rect 2691 2425 2692 2429
rect 2686 2424 2692 2425
rect 2822 2429 2828 2430
rect 2822 2425 2823 2429
rect 2827 2425 2828 2429
rect 2833 2428 2835 2438
rect 3078 2435 3079 2439
rect 3083 2435 3084 2439
rect 3078 2434 3084 2435
rect 3087 2439 3093 2440
rect 3087 2435 3088 2439
rect 3092 2438 3093 2439
rect 3190 2439 3191 2443
rect 3195 2439 3196 2443
rect 3190 2438 3196 2439
rect 3092 2436 3123 2438
rect 3092 2435 3093 2436
rect 3087 2434 3093 2435
rect 2966 2429 2972 2430
rect 2822 2424 2828 2425
rect 2831 2427 2837 2428
rect 2574 2422 2580 2423
rect 2666 2423 2672 2424
rect 2399 2418 2405 2419
rect 2666 2419 2667 2423
rect 2671 2422 2672 2423
rect 2695 2423 2701 2424
rect 2695 2422 2696 2423
rect 2671 2420 2696 2422
rect 2671 2419 2672 2420
rect 2666 2418 2672 2419
rect 2695 2419 2696 2420
rect 2700 2422 2701 2423
rect 2831 2423 2832 2427
rect 2836 2423 2837 2427
rect 2966 2425 2967 2429
rect 2971 2425 2972 2429
rect 2966 2424 2972 2425
rect 3110 2429 3116 2430
rect 3110 2425 3111 2429
rect 3115 2425 3116 2429
rect 3110 2424 3116 2425
rect 3121 2424 3123 2436
rect 3190 2425 3196 2426
rect 2831 2422 2837 2423
rect 2974 2423 2981 2424
rect 2700 2420 2835 2422
rect 2700 2419 2701 2420
rect 2695 2418 2701 2419
rect 2974 2419 2975 2423
rect 2980 2422 2981 2423
rect 3014 2423 3020 2424
rect 3014 2422 3015 2423
rect 2980 2420 3015 2422
rect 2980 2419 2981 2420
rect 2974 2418 2981 2419
rect 3014 2419 3015 2420
rect 3019 2419 3020 2423
rect 3014 2418 3020 2419
rect 3119 2423 3125 2424
rect 3119 2419 3120 2423
rect 3124 2422 3125 2423
rect 3142 2423 3148 2424
rect 3142 2422 3143 2423
rect 3124 2420 3143 2422
rect 3124 2419 3125 2420
rect 3119 2418 3125 2419
rect 3142 2419 3143 2420
rect 3147 2422 3148 2423
rect 3166 2423 3172 2424
rect 3166 2422 3167 2423
rect 3147 2420 3167 2422
rect 3147 2419 3148 2420
rect 3142 2418 3148 2419
rect 3166 2419 3167 2420
rect 3171 2419 3172 2423
rect 3190 2421 3191 2425
rect 3195 2421 3196 2425
rect 3190 2420 3196 2421
rect 3166 2418 3172 2419
rect 1670 2407 1676 2408
rect 1670 2403 1671 2407
rect 1675 2403 1676 2407
rect 1670 2402 1676 2403
rect 3190 2407 3196 2408
rect 3190 2403 3191 2407
rect 3195 2403 3196 2407
rect 3190 2402 3196 2403
rect 2230 2400 2236 2401
rect 134 2396 140 2397
rect 134 2392 135 2396
rect 139 2392 140 2396
rect 134 2391 140 2392
rect 238 2396 244 2397
rect 238 2392 239 2396
rect 243 2392 244 2396
rect 238 2391 244 2392
rect 358 2396 364 2397
rect 358 2392 359 2396
rect 363 2392 364 2396
rect 358 2391 364 2392
rect 478 2396 484 2397
rect 478 2392 479 2396
rect 483 2392 484 2396
rect 478 2391 484 2392
rect 590 2396 596 2397
rect 590 2392 591 2396
rect 595 2392 596 2396
rect 590 2391 596 2392
rect 702 2396 708 2397
rect 702 2392 703 2396
rect 707 2392 708 2396
rect 702 2391 708 2392
rect 814 2396 820 2397
rect 814 2392 815 2396
rect 819 2392 820 2396
rect 814 2391 820 2392
rect 934 2396 940 2397
rect 934 2392 935 2396
rect 939 2392 940 2396
rect 2230 2396 2231 2400
rect 2235 2396 2236 2400
rect 2230 2395 2236 2396
rect 2390 2400 2396 2401
rect 2390 2396 2391 2400
rect 2395 2396 2396 2400
rect 2390 2395 2396 2396
rect 2542 2400 2548 2401
rect 2542 2396 2543 2400
rect 2547 2396 2548 2400
rect 2542 2395 2548 2396
rect 2686 2400 2692 2401
rect 2686 2396 2687 2400
rect 2691 2396 2692 2400
rect 2686 2395 2692 2396
rect 2822 2400 2828 2401
rect 2822 2396 2823 2400
rect 2827 2396 2828 2400
rect 2822 2395 2828 2396
rect 2966 2400 2972 2401
rect 2966 2396 2967 2400
rect 2971 2396 2972 2400
rect 2966 2395 2972 2396
rect 3110 2400 3116 2401
rect 3110 2396 3111 2400
rect 3115 2396 3116 2400
rect 3110 2395 3116 2396
rect 934 2391 940 2392
rect 110 2389 116 2390
rect 110 2385 111 2389
rect 115 2385 116 2389
rect 110 2384 116 2385
rect 1630 2389 1636 2390
rect 1630 2385 1631 2389
rect 1635 2385 1636 2389
rect 1630 2384 1636 2385
rect 2142 2380 2148 2381
rect 610 2379 616 2380
rect 610 2378 611 2379
rect 600 2376 611 2378
rect 600 2374 602 2376
rect 610 2375 611 2376
rect 615 2375 616 2379
rect 2142 2376 2143 2380
rect 2147 2376 2148 2380
rect 2142 2375 2148 2376
rect 2310 2380 2316 2381
rect 2310 2376 2311 2380
rect 2315 2376 2316 2380
rect 2310 2375 2316 2376
rect 2478 2380 2484 2381
rect 2478 2376 2479 2380
rect 2483 2376 2484 2380
rect 2478 2375 2484 2376
rect 2654 2380 2660 2381
rect 2654 2376 2655 2380
rect 2659 2376 2660 2380
rect 2654 2375 2660 2376
rect 2830 2380 2836 2381
rect 2830 2376 2831 2380
rect 2835 2376 2836 2380
rect 2830 2375 2836 2376
rect 3006 2380 3012 2381
rect 3006 2376 3007 2380
rect 3011 2376 3012 2380
rect 3006 2375 3012 2376
rect 3158 2380 3164 2381
rect 3158 2376 3159 2380
rect 3163 2376 3164 2380
rect 3158 2375 3164 2376
rect 610 2374 616 2375
rect 576 2372 602 2374
rect 1670 2373 1676 2374
rect 110 2371 116 2372
rect 110 2367 111 2371
rect 115 2367 116 2371
rect 576 2368 578 2372
rect 600 2370 602 2372
rect 1630 2371 1636 2372
rect 599 2369 605 2370
rect 110 2366 116 2367
rect 134 2367 140 2368
rect 134 2363 135 2367
rect 139 2363 140 2367
rect 134 2362 140 2363
rect 142 2367 149 2368
rect 142 2363 143 2367
rect 148 2363 149 2367
rect 142 2362 149 2363
rect 238 2367 244 2368
rect 238 2363 239 2367
rect 243 2363 244 2367
rect 238 2362 244 2363
rect 246 2367 253 2368
rect 246 2363 247 2367
rect 252 2363 253 2367
rect 246 2362 253 2363
rect 358 2367 364 2368
rect 358 2363 359 2367
rect 363 2363 364 2367
rect 358 2362 364 2363
rect 366 2367 373 2368
rect 366 2363 367 2367
rect 372 2363 373 2367
rect 366 2362 373 2363
rect 478 2367 484 2368
rect 478 2363 479 2367
rect 483 2363 484 2367
rect 478 2362 484 2363
rect 487 2367 493 2368
rect 487 2363 488 2367
rect 492 2366 493 2367
rect 574 2367 580 2368
rect 574 2366 575 2367
rect 492 2364 575 2366
rect 492 2363 493 2364
rect 487 2362 493 2363
rect 574 2363 575 2364
rect 579 2363 580 2367
rect 574 2362 580 2363
rect 590 2367 596 2368
rect 590 2363 591 2367
rect 595 2363 596 2367
rect 599 2365 600 2369
rect 604 2365 605 2369
rect 599 2364 605 2365
rect 702 2367 708 2368
rect 590 2362 596 2363
rect 702 2363 703 2367
rect 707 2363 708 2367
rect 702 2362 708 2363
rect 711 2367 717 2368
rect 711 2363 712 2367
rect 716 2366 717 2367
rect 774 2367 780 2368
rect 774 2366 775 2367
rect 716 2364 775 2366
rect 716 2363 717 2364
rect 711 2362 717 2363
rect 774 2363 775 2364
rect 779 2366 780 2367
rect 814 2367 820 2368
rect 779 2364 794 2366
rect 779 2363 780 2364
rect 774 2362 780 2363
rect 792 2360 794 2364
rect 814 2363 815 2367
rect 819 2363 820 2367
rect 814 2362 820 2363
rect 823 2367 829 2368
rect 823 2363 824 2367
rect 828 2363 829 2367
rect 823 2362 829 2363
rect 934 2367 940 2368
rect 934 2363 935 2367
rect 939 2363 940 2367
rect 934 2362 940 2363
rect 942 2367 949 2368
rect 942 2363 943 2367
rect 948 2366 949 2367
rect 982 2367 988 2368
rect 982 2366 983 2367
rect 948 2364 983 2366
rect 948 2363 949 2364
rect 942 2362 949 2363
rect 982 2363 983 2364
rect 987 2363 988 2367
rect 1630 2367 1631 2371
rect 1635 2367 1636 2371
rect 1670 2369 1671 2373
rect 1675 2369 1676 2373
rect 1670 2368 1676 2369
rect 3190 2373 3196 2374
rect 3190 2369 3191 2373
rect 3195 2369 3196 2373
rect 3190 2368 3196 2369
rect 1630 2366 1636 2367
rect 982 2362 988 2363
rect 790 2359 796 2360
rect 790 2355 791 2359
rect 795 2358 796 2359
rect 824 2358 826 2362
rect 3166 2359 3172 2360
rect 3166 2358 3167 2359
rect 795 2356 826 2358
rect 3017 2356 3167 2358
rect 795 2355 796 2356
rect 790 2354 796 2355
rect 1670 2355 1676 2356
rect 1670 2351 1671 2355
rect 1675 2351 1676 2355
rect 2238 2355 2244 2356
rect 2238 2354 2239 2355
rect 2196 2352 2239 2354
rect 1670 2350 1676 2351
rect 2142 2351 2148 2352
rect 134 2349 140 2350
rect 110 2345 116 2346
rect 110 2341 111 2345
rect 115 2341 116 2345
rect 134 2345 135 2349
rect 139 2345 140 2349
rect 134 2344 140 2345
rect 342 2349 348 2350
rect 342 2345 343 2349
rect 347 2345 348 2349
rect 342 2344 348 2345
rect 566 2349 572 2350
rect 566 2345 567 2349
rect 571 2345 572 2349
rect 566 2344 572 2345
rect 774 2349 780 2350
rect 774 2345 775 2349
rect 779 2345 780 2349
rect 774 2344 780 2345
rect 974 2349 980 2350
rect 974 2345 975 2349
rect 979 2345 980 2349
rect 1174 2349 1180 2350
rect 974 2344 980 2345
rect 982 2347 989 2348
rect 110 2340 116 2341
rect 142 2343 149 2344
rect 142 2339 143 2343
rect 148 2342 149 2343
rect 182 2343 188 2344
rect 182 2342 183 2343
rect 148 2340 183 2342
rect 148 2339 149 2340
rect 142 2338 149 2339
rect 182 2339 183 2340
rect 187 2342 188 2343
rect 246 2343 252 2344
rect 246 2342 247 2343
rect 187 2340 247 2342
rect 187 2339 188 2340
rect 182 2338 188 2339
rect 246 2339 247 2340
rect 251 2342 252 2343
rect 351 2343 357 2344
rect 351 2342 352 2343
rect 251 2340 352 2342
rect 251 2339 252 2340
rect 246 2338 252 2339
rect 351 2339 352 2340
rect 356 2342 357 2343
rect 366 2343 372 2344
rect 366 2342 367 2343
rect 356 2340 367 2342
rect 356 2339 357 2340
rect 351 2338 357 2339
rect 366 2339 367 2340
rect 371 2339 372 2343
rect 366 2338 372 2339
rect 574 2343 581 2344
rect 574 2339 575 2343
rect 580 2339 581 2343
rect 574 2338 581 2339
rect 782 2343 789 2344
rect 782 2339 783 2343
rect 788 2339 789 2343
rect 982 2343 983 2347
rect 988 2343 989 2347
rect 1174 2345 1175 2349
rect 1179 2345 1180 2349
rect 1174 2344 1180 2345
rect 1366 2349 1372 2350
rect 1366 2345 1367 2349
rect 1371 2345 1372 2349
rect 1566 2349 1572 2350
rect 1366 2344 1372 2345
rect 1374 2347 1381 2348
rect 982 2342 989 2343
rect 1166 2343 1172 2344
rect 782 2338 789 2339
rect 1166 2339 1167 2343
rect 1171 2342 1172 2343
rect 1182 2343 1189 2344
rect 1182 2342 1183 2343
rect 1171 2340 1183 2342
rect 1171 2339 1172 2340
rect 1166 2338 1172 2339
rect 1182 2339 1183 2340
rect 1188 2339 1189 2343
rect 1374 2343 1375 2347
rect 1380 2343 1381 2347
rect 1566 2345 1567 2349
rect 1571 2345 1572 2349
rect 1566 2344 1572 2345
rect 1574 2347 1581 2348
rect 1374 2342 1381 2343
rect 1574 2343 1575 2347
rect 1580 2343 1581 2347
rect 2142 2347 2143 2351
rect 2147 2347 2148 2351
rect 2142 2346 2148 2347
rect 2151 2351 2157 2352
rect 2151 2347 2152 2351
rect 2156 2350 2157 2351
rect 2174 2351 2180 2352
rect 2174 2350 2175 2351
rect 2156 2348 2175 2350
rect 2156 2347 2157 2348
rect 2151 2346 2157 2347
rect 2174 2347 2175 2348
rect 2179 2350 2180 2351
rect 2196 2350 2198 2352
rect 2238 2351 2239 2352
rect 2243 2351 2244 2355
rect 2319 2355 2325 2356
rect 2238 2350 2244 2351
rect 2310 2351 2316 2352
rect 2179 2348 2198 2350
rect 2179 2347 2180 2348
rect 2174 2346 2180 2347
rect 2310 2347 2311 2351
rect 2315 2347 2316 2351
rect 2319 2351 2320 2355
rect 2324 2354 2325 2355
rect 2342 2355 2348 2356
rect 2342 2354 2343 2355
rect 2324 2352 2343 2354
rect 2324 2351 2325 2352
rect 2319 2350 2325 2351
rect 2342 2351 2343 2352
rect 2347 2351 2348 2355
rect 2663 2355 2672 2356
rect 2342 2350 2348 2351
rect 2478 2351 2484 2352
rect 2310 2346 2316 2347
rect 2478 2347 2479 2351
rect 2483 2347 2484 2351
rect 2478 2346 2484 2347
rect 2487 2351 2493 2352
rect 2487 2347 2488 2351
rect 2492 2347 2493 2351
rect 2487 2346 2493 2347
rect 2654 2351 2660 2352
rect 2654 2347 2655 2351
rect 2659 2347 2660 2351
rect 2663 2351 2664 2355
rect 2671 2351 2672 2355
rect 3014 2355 3021 2356
rect 2663 2350 2672 2351
rect 2830 2351 2836 2352
rect 2654 2346 2660 2347
rect 2830 2347 2831 2351
rect 2835 2347 2836 2351
rect 2830 2346 2836 2347
rect 2839 2351 2845 2352
rect 2839 2347 2840 2351
rect 2844 2350 2845 2351
rect 3006 2351 3012 2352
rect 2844 2348 2931 2350
rect 2844 2347 2845 2348
rect 2839 2346 2845 2347
rect 1574 2342 1581 2343
rect 1630 2345 1636 2346
rect 1630 2341 1631 2345
rect 1635 2341 1636 2345
rect 1630 2340 1636 2341
rect 2182 2341 2188 2342
rect 1182 2338 1189 2339
rect 1670 2337 1676 2338
rect 1670 2333 1671 2337
rect 1675 2333 1676 2337
rect 2182 2337 2183 2341
rect 2187 2337 2188 2341
rect 2182 2336 2188 2337
rect 2334 2341 2340 2342
rect 2334 2337 2335 2341
rect 2339 2337 2340 2341
rect 2478 2341 2484 2342
rect 2334 2336 2340 2337
rect 2342 2339 2349 2340
rect 1670 2332 1676 2333
rect 2174 2335 2180 2336
rect 2174 2331 2175 2335
rect 2179 2334 2180 2335
rect 2191 2335 2197 2336
rect 2191 2334 2192 2335
rect 2179 2332 2192 2334
rect 2179 2331 2180 2332
rect 2174 2330 2180 2331
rect 2191 2331 2192 2332
rect 2196 2331 2197 2335
rect 2342 2335 2343 2339
rect 2348 2335 2349 2339
rect 2478 2337 2479 2341
rect 2483 2337 2484 2341
rect 2478 2336 2484 2337
rect 2488 2336 2490 2346
rect 2622 2341 2628 2342
rect 2622 2337 2623 2341
rect 2627 2337 2628 2341
rect 2766 2341 2772 2342
rect 2622 2336 2628 2337
rect 2630 2339 2637 2340
rect 2342 2334 2349 2335
rect 2486 2335 2493 2336
rect 2191 2330 2197 2331
rect 2486 2331 2487 2335
rect 2492 2334 2493 2335
rect 2630 2335 2631 2339
rect 2636 2338 2637 2339
rect 2666 2339 2672 2340
rect 2666 2338 2667 2339
rect 2636 2336 2667 2338
rect 2636 2335 2637 2336
rect 2630 2334 2637 2335
rect 2666 2335 2667 2336
rect 2671 2335 2672 2339
rect 2766 2337 2767 2341
rect 2771 2337 2772 2341
rect 2766 2336 2772 2337
rect 2775 2339 2781 2340
rect 2666 2334 2672 2335
rect 2775 2335 2776 2339
rect 2780 2338 2781 2339
rect 2798 2339 2804 2340
rect 2798 2338 2799 2339
rect 2780 2336 2799 2338
rect 2780 2335 2781 2336
rect 2775 2334 2781 2335
rect 2798 2335 2799 2336
rect 2803 2338 2804 2339
rect 2839 2338 2841 2346
rect 2803 2336 2841 2338
rect 2918 2341 2924 2342
rect 2918 2337 2919 2341
rect 2923 2337 2924 2341
rect 2929 2340 2931 2348
rect 3006 2347 3007 2351
rect 3011 2347 3012 2351
rect 3014 2351 3015 2355
rect 3020 2351 3021 2355
rect 3166 2355 3167 2356
rect 3171 2355 3172 2359
rect 3166 2354 3172 2355
rect 3190 2355 3196 2356
rect 3014 2350 3021 2351
rect 3158 2351 3164 2352
rect 3006 2346 3012 2347
rect 3158 2347 3159 2351
rect 3163 2347 3164 2351
rect 3158 2346 3164 2347
rect 3166 2351 3173 2352
rect 3166 2347 3167 2351
rect 3172 2347 3173 2351
rect 3190 2351 3191 2355
rect 3195 2351 3196 2355
rect 3190 2350 3196 2351
rect 3166 2346 3173 2347
rect 2918 2336 2924 2337
rect 2927 2339 2933 2340
rect 2803 2335 2804 2336
rect 2798 2334 2804 2335
rect 2927 2335 2928 2339
rect 2932 2338 2933 2339
rect 3014 2339 3020 2340
rect 3014 2338 3015 2339
rect 2932 2336 3015 2338
rect 2932 2335 2933 2336
rect 2927 2334 2933 2335
rect 3014 2335 3015 2336
rect 3019 2335 3020 2339
rect 3014 2334 3020 2335
rect 3190 2337 3196 2338
rect 2492 2332 2634 2334
rect 3190 2333 3191 2337
rect 3195 2333 3196 2337
rect 3190 2332 3196 2333
rect 2492 2331 2493 2332
rect 2486 2330 2493 2331
rect 110 2327 116 2328
rect 110 2323 111 2327
rect 115 2323 116 2327
rect 110 2322 116 2323
rect 1630 2327 1636 2328
rect 1630 2323 1631 2327
rect 1635 2323 1636 2327
rect 1630 2322 1636 2323
rect 134 2320 140 2321
rect 134 2316 135 2320
rect 139 2316 140 2320
rect 134 2315 140 2316
rect 342 2320 348 2321
rect 342 2316 343 2320
rect 347 2316 348 2320
rect 342 2315 348 2316
rect 566 2320 572 2321
rect 566 2316 567 2320
rect 571 2316 572 2320
rect 566 2315 572 2316
rect 774 2320 780 2321
rect 774 2316 775 2320
rect 779 2316 780 2320
rect 774 2315 780 2316
rect 974 2320 980 2321
rect 974 2316 975 2320
rect 979 2316 980 2320
rect 974 2315 980 2316
rect 1174 2320 1180 2321
rect 1174 2316 1175 2320
rect 1179 2316 1180 2320
rect 1174 2315 1180 2316
rect 1366 2320 1372 2321
rect 1366 2316 1367 2320
rect 1371 2316 1372 2320
rect 1366 2315 1372 2316
rect 1566 2320 1572 2321
rect 1566 2316 1567 2320
rect 1571 2316 1572 2320
rect 1566 2315 1572 2316
rect 1670 2319 1676 2320
rect 1670 2315 1671 2319
rect 1675 2315 1676 2319
rect 1670 2314 1676 2315
rect 3190 2319 3196 2320
rect 3190 2315 3191 2319
rect 3195 2315 3196 2319
rect 3190 2314 3196 2315
rect 2182 2312 2188 2313
rect 2182 2308 2183 2312
rect 2187 2308 2188 2312
rect 2182 2307 2188 2308
rect 2334 2312 2340 2313
rect 2334 2308 2335 2312
rect 2339 2308 2340 2312
rect 2334 2307 2340 2308
rect 2478 2312 2484 2313
rect 2478 2308 2479 2312
rect 2483 2308 2484 2312
rect 2478 2307 2484 2308
rect 2622 2312 2628 2313
rect 2622 2308 2623 2312
rect 2627 2308 2628 2312
rect 2622 2307 2628 2308
rect 2766 2312 2772 2313
rect 2766 2308 2767 2312
rect 2771 2308 2772 2312
rect 2766 2307 2772 2308
rect 2918 2312 2924 2313
rect 2918 2308 2919 2312
rect 2923 2308 2924 2312
rect 2918 2307 2924 2308
rect 654 2296 660 2297
rect 654 2292 655 2296
rect 659 2292 660 2296
rect 654 2291 660 2292
rect 782 2296 788 2297
rect 782 2292 783 2296
rect 787 2292 788 2296
rect 782 2291 788 2292
rect 902 2296 908 2297
rect 902 2292 903 2296
rect 907 2292 908 2296
rect 902 2291 908 2292
rect 1022 2296 1028 2297
rect 1022 2292 1023 2296
rect 1027 2292 1028 2296
rect 1022 2291 1028 2292
rect 1142 2296 1148 2297
rect 1142 2292 1143 2296
rect 1147 2292 1148 2296
rect 1142 2291 1148 2292
rect 1254 2296 1260 2297
rect 1254 2292 1255 2296
rect 1259 2292 1260 2296
rect 1254 2291 1260 2292
rect 1366 2296 1372 2297
rect 1366 2292 1367 2296
rect 1371 2292 1372 2296
rect 1366 2291 1372 2292
rect 1486 2296 1492 2297
rect 1486 2292 1487 2296
rect 1491 2292 1492 2296
rect 1486 2291 1492 2292
rect 2094 2296 2100 2297
rect 2094 2292 2095 2296
rect 2099 2292 2100 2296
rect 2094 2291 2100 2292
rect 2262 2296 2268 2297
rect 2262 2292 2263 2296
rect 2267 2292 2268 2296
rect 2262 2291 2268 2292
rect 2430 2296 2436 2297
rect 2430 2292 2431 2296
rect 2435 2292 2436 2296
rect 2430 2291 2436 2292
rect 2606 2296 2612 2297
rect 2606 2292 2607 2296
rect 2611 2292 2612 2296
rect 2606 2291 2612 2292
rect 2790 2296 2796 2297
rect 2790 2292 2791 2296
rect 2795 2292 2796 2296
rect 2790 2291 2796 2292
rect 2982 2296 2988 2297
rect 2982 2292 2983 2296
rect 2987 2292 2988 2296
rect 2982 2291 2988 2292
rect 3158 2296 3164 2297
rect 3158 2292 3159 2296
rect 3163 2292 3164 2296
rect 3158 2291 3164 2292
rect 110 2289 116 2290
rect 110 2285 111 2289
rect 115 2285 116 2289
rect 110 2284 116 2285
rect 1630 2289 1636 2290
rect 1630 2285 1631 2289
rect 1635 2285 1636 2289
rect 1630 2284 1636 2285
rect 1670 2289 1676 2290
rect 1670 2285 1671 2289
rect 1675 2285 1676 2289
rect 1670 2284 1676 2285
rect 3190 2289 3196 2290
rect 3190 2285 3191 2289
rect 3195 2285 3196 2289
rect 3190 2284 3196 2285
rect 1398 2275 1404 2276
rect 952 2272 1034 2274
rect 1056 2272 1154 2274
rect 1168 2272 1266 2274
rect 110 2271 116 2272
rect 110 2267 111 2271
rect 115 2267 116 2271
rect 911 2271 917 2272
rect 110 2266 116 2267
rect 654 2267 660 2268
rect 654 2263 655 2267
rect 659 2263 660 2267
rect 654 2262 660 2263
rect 662 2267 669 2268
rect 662 2263 663 2267
rect 668 2263 669 2267
rect 662 2262 669 2263
rect 782 2267 788 2268
rect 782 2263 783 2267
rect 787 2263 788 2267
rect 782 2262 788 2263
rect 790 2267 797 2268
rect 790 2263 791 2267
rect 796 2266 797 2267
rect 814 2267 820 2268
rect 814 2266 815 2267
rect 796 2264 815 2266
rect 796 2263 797 2264
rect 790 2262 797 2263
rect 814 2263 815 2264
rect 819 2263 820 2267
rect 814 2262 820 2263
rect 902 2267 908 2268
rect 902 2263 903 2267
rect 907 2263 908 2267
rect 911 2267 912 2271
rect 916 2270 917 2271
rect 942 2271 948 2272
rect 942 2270 943 2271
rect 916 2268 943 2270
rect 916 2267 917 2268
rect 911 2266 917 2267
rect 942 2267 943 2268
rect 947 2270 948 2271
rect 950 2271 956 2272
rect 950 2270 951 2271
rect 947 2268 951 2270
rect 947 2267 948 2268
rect 942 2266 948 2267
rect 950 2267 951 2268
rect 955 2267 956 2271
rect 1031 2271 1037 2272
rect 950 2266 956 2267
rect 1022 2267 1028 2268
rect 902 2262 908 2263
rect 1022 2263 1023 2267
rect 1027 2263 1028 2267
rect 1031 2267 1032 2271
rect 1036 2270 1037 2271
rect 1054 2271 1060 2272
rect 1054 2270 1055 2271
rect 1036 2268 1055 2270
rect 1036 2267 1037 2268
rect 1031 2266 1037 2267
rect 1054 2267 1055 2268
rect 1059 2267 1060 2271
rect 1151 2271 1157 2272
rect 1054 2266 1060 2267
rect 1142 2267 1148 2268
rect 1022 2262 1028 2263
rect 1142 2263 1143 2267
rect 1147 2263 1148 2267
rect 1151 2267 1152 2271
rect 1156 2270 1157 2271
rect 1166 2271 1172 2272
rect 1166 2270 1167 2271
rect 1156 2268 1167 2270
rect 1156 2267 1157 2268
rect 1151 2266 1157 2267
rect 1166 2267 1167 2268
rect 1171 2267 1172 2271
rect 1263 2271 1269 2272
rect 1166 2266 1172 2267
rect 1254 2267 1260 2268
rect 1142 2262 1148 2263
rect 1254 2263 1255 2267
rect 1259 2263 1260 2267
rect 1263 2267 1264 2271
rect 1268 2270 1269 2271
rect 1278 2271 1284 2272
rect 1278 2270 1279 2271
rect 1268 2268 1279 2270
rect 1268 2267 1269 2268
rect 1263 2266 1269 2267
rect 1278 2267 1279 2268
rect 1283 2267 1284 2271
rect 1398 2271 1399 2275
rect 1403 2274 1404 2275
rect 2022 2275 2028 2276
rect 1403 2272 1498 2274
rect 1403 2271 1404 2272
rect 1398 2270 1404 2271
rect 1495 2271 1501 2272
rect 1278 2266 1284 2267
rect 1366 2267 1372 2268
rect 1254 2262 1260 2263
rect 1366 2263 1367 2267
rect 1371 2263 1372 2267
rect 1366 2262 1372 2263
rect 1374 2267 1381 2268
rect 1374 2263 1375 2267
rect 1380 2266 1381 2267
rect 1399 2266 1401 2270
rect 1380 2264 1401 2266
rect 1486 2267 1492 2268
rect 1380 2263 1381 2264
rect 1374 2262 1381 2263
rect 1486 2263 1487 2267
rect 1491 2263 1492 2267
rect 1495 2267 1496 2271
rect 1500 2267 1501 2271
rect 1495 2266 1501 2267
rect 1630 2271 1636 2272
rect 1630 2267 1631 2271
rect 1635 2267 1636 2271
rect 1630 2266 1636 2267
rect 1670 2271 1676 2272
rect 1670 2267 1671 2271
rect 1675 2267 1676 2271
rect 2022 2271 2023 2275
rect 2027 2274 2028 2275
rect 2027 2273 2109 2274
rect 2027 2272 2104 2273
rect 2027 2271 2028 2272
rect 2022 2270 2028 2271
rect 2103 2269 2104 2272
rect 2108 2269 2109 2273
rect 2103 2268 2109 2269
rect 2798 2271 2805 2272
rect 1670 2266 1676 2267
rect 2094 2267 2100 2268
rect 1486 2262 1492 2263
rect 2094 2263 2095 2267
rect 2099 2263 2100 2267
rect 2094 2262 2100 2263
rect 2262 2267 2268 2268
rect 2262 2263 2263 2267
rect 2267 2263 2268 2267
rect 2262 2262 2268 2263
rect 2271 2267 2277 2268
rect 2271 2263 2272 2267
rect 2276 2266 2277 2267
rect 2302 2267 2308 2268
rect 2302 2266 2303 2267
rect 2276 2264 2303 2266
rect 2276 2263 2277 2264
rect 2271 2262 2277 2263
rect 2302 2263 2303 2264
rect 2307 2263 2308 2267
rect 2302 2262 2308 2263
rect 2430 2267 2436 2268
rect 2430 2263 2431 2267
rect 2435 2263 2436 2267
rect 2430 2262 2436 2263
rect 2439 2267 2445 2268
rect 2439 2263 2440 2267
rect 2444 2266 2445 2267
rect 2486 2267 2492 2268
rect 2486 2266 2487 2267
rect 2444 2264 2487 2266
rect 2444 2263 2445 2264
rect 2439 2262 2445 2263
rect 2486 2263 2487 2264
rect 2491 2263 2492 2267
rect 2486 2262 2492 2263
rect 2606 2267 2612 2268
rect 2606 2263 2607 2267
rect 2611 2263 2612 2267
rect 2606 2262 2612 2263
rect 2615 2267 2621 2268
rect 2615 2263 2616 2267
rect 2620 2266 2621 2267
rect 2630 2267 2636 2268
rect 2630 2266 2631 2267
rect 2620 2264 2631 2266
rect 2620 2263 2621 2264
rect 2615 2262 2621 2263
rect 2630 2263 2631 2264
rect 2635 2263 2636 2267
rect 2630 2262 2636 2263
rect 2790 2267 2796 2268
rect 2790 2263 2791 2267
rect 2795 2263 2796 2267
rect 2798 2267 2799 2271
rect 2804 2267 2805 2271
rect 2990 2271 2997 2272
rect 2798 2266 2805 2267
rect 2982 2267 2988 2268
rect 2790 2262 2796 2263
rect 2982 2263 2983 2267
rect 2987 2263 2988 2267
rect 2990 2267 2991 2271
rect 2996 2270 2997 2271
rect 3014 2271 3020 2272
rect 3014 2270 3015 2271
rect 2996 2268 3015 2270
rect 2996 2267 2997 2268
rect 2990 2266 2997 2267
rect 3014 2267 3015 2268
rect 3019 2267 3020 2271
rect 3190 2271 3196 2272
rect 3014 2266 3020 2267
rect 3158 2267 3164 2268
rect 2982 2262 2988 2263
rect 3158 2263 3159 2267
rect 3163 2263 3164 2267
rect 3158 2262 3164 2263
rect 3166 2267 3173 2268
rect 3166 2263 3167 2267
rect 3172 2263 3173 2267
rect 3190 2267 3191 2271
rect 3195 2267 3196 2271
rect 3190 2266 3196 2267
rect 3166 2262 3173 2263
rect 2014 2257 2020 2258
rect 1670 2253 1676 2254
rect 1670 2249 1671 2253
rect 1675 2249 1676 2253
rect 2014 2253 2015 2257
rect 2019 2253 2020 2257
rect 2014 2252 2020 2253
rect 2166 2257 2172 2258
rect 2166 2253 2167 2257
rect 2171 2253 2172 2257
rect 2166 2252 2172 2253
rect 2318 2257 2324 2258
rect 2318 2253 2319 2257
rect 2323 2253 2324 2257
rect 2318 2252 2324 2253
rect 2462 2257 2468 2258
rect 2462 2253 2463 2257
rect 2467 2253 2468 2257
rect 2606 2257 2612 2258
rect 2462 2252 2468 2253
rect 2471 2255 2477 2256
rect 1670 2248 1676 2249
rect 2022 2251 2029 2252
rect 1054 2247 1060 2248
rect 550 2245 556 2246
rect 110 2241 116 2242
rect 110 2237 111 2241
rect 115 2237 116 2241
rect 550 2241 551 2245
rect 555 2241 556 2245
rect 550 2240 556 2241
rect 678 2245 684 2246
rect 678 2241 679 2245
rect 683 2241 684 2245
rect 678 2240 684 2241
rect 806 2245 812 2246
rect 806 2241 807 2245
rect 811 2241 812 2245
rect 926 2245 932 2246
rect 806 2240 812 2241
rect 814 2243 821 2244
rect 110 2236 116 2237
rect 559 2239 565 2240
rect 559 2235 560 2239
rect 564 2238 565 2239
rect 574 2239 580 2240
rect 574 2238 575 2239
rect 564 2236 575 2238
rect 564 2235 565 2236
rect 559 2234 565 2235
rect 574 2235 575 2236
rect 579 2238 580 2239
rect 606 2239 612 2240
rect 606 2238 607 2239
rect 579 2236 607 2238
rect 579 2235 580 2236
rect 574 2234 580 2235
rect 606 2235 607 2236
rect 611 2238 612 2239
rect 662 2239 668 2240
rect 662 2238 663 2239
rect 611 2236 663 2238
rect 611 2235 612 2236
rect 606 2234 612 2235
rect 662 2235 663 2236
rect 667 2238 668 2239
rect 687 2239 693 2240
rect 687 2238 688 2239
rect 667 2236 688 2238
rect 667 2235 668 2236
rect 662 2234 668 2235
rect 687 2235 688 2236
rect 692 2235 693 2239
rect 814 2239 815 2243
rect 820 2239 821 2243
rect 926 2241 927 2245
rect 931 2241 932 2245
rect 926 2240 932 2241
rect 1046 2245 1052 2246
rect 1046 2241 1047 2245
rect 1051 2241 1052 2245
rect 1054 2243 1055 2247
rect 1059 2246 1060 2247
rect 1166 2247 1172 2248
rect 1059 2245 1061 2246
rect 1054 2242 1056 2243
rect 1046 2240 1052 2241
rect 1055 2241 1056 2242
rect 1060 2241 1061 2245
rect 1055 2240 1061 2241
rect 1158 2245 1164 2246
rect 1158 2241 1159 2245
rect 1163 2241 1164 2245
rect 1166 2243 1167 2247
rect 1171 2246 1172 2247
rect 2022 2247 2023 2251
rect 2028 2247 2029 2251
rect 2022 2246 2029 2247
rect 2174 2251 2181 2252
rect 2174 2247 2175 2251
rect 2180 2247 2181 2251
rect 2174 2246 2181 2247
rect 2302 2251 2308 2252
rect 2302 2247 2303 2251
rect 2307 2250 2308 2251
rect 2327 2251 2333 2252
rect 2327 2250 2328 2251
rect 2307 2248 2328 2250
rect 2307 2247 2308 2248
rect 2302 2246 2308 2247
rect 2327 2247 2328 2248
rect 2332 2250 2333 2251
rect 2471 2251 2472 2255
rect 2476 2254 2477 2255
rect 2486 2255 2492 2256
rect 2486 2254 2487 2255
rect 2476 2252 2487 2254
rect 2476 2251 2477 2252
rect 2471 2250 2477 2251
rect 2486 2251 2487 2252
rect 2491 2251 2492 2255
rect 2606 2253 2607 2257
rect 2611 2253 2612 2257
rect 2617 2256 2619 2262
rect 2758 2257 2764 2258
rect 2606 2252 2612 2253
rect 2614 2255 2621 2256
rect 2486 2250 2492 2251
rect 2614 2251 2615 2255
rect 2620 2251 2621 2255
rect 2758 2253 2759 2257
rect 2763 2253 2764 2257
rect 2758 2252 2764 2253
rect 2766 2255 2773 2256
rect 2614 2250 2621 2251
rect 2766 2251 2767 2255
rect 2772 2254 2773 2255
rect 2798 2255 2804 2256
rect 2798 2254 2799 2255
rect 2772 2252 2799 2254
rect 2772 2251 2773 2252
rect 2766 2250 2773 2251
rect 2798 2251 2799 2252
rect 2803 2251 2804 2255
rect 2798 2250 2804 2251
rect 3190 2253 3196 2254
rect 2332 2248 2474 2250
rect 3190 2249 3191 2253
rect 3195 2249 3196 2253
rect 3190 2248 3196 2249
rect 2332 2247 2333 2248
rect 2327 2246 2333 2247
rect 1171 2245 1173 2246
rect 1166 2242 1168 2243
rect 1158 2240 1164 2241
rect 1167 2241 1168 2242
rect 1172 2241 1173 2245
rect 1167 2240 1173 2241
rect 1270 2245 1276 2246
rect 1270 2241 1271 2245
rect 1275 2241 1276 2245
rect 1390 2245 1396 2246
rect 1270 2240 1276 2241
rect 1278 2243 1285 2244
rect 814 2238 821 2239
rect 935 2239 941 2240
rect 687 2234 693 2235
rect 935 2235 936 2239
rect 940 2238 941 2239
rect 950 2239 956 2240
rect 950 2238 951 2239
rect 940 2236 951 2238
rect 940 2235 941 2236
rect 935 2234 941 2235
rect 950 2235 951 2236
rect 955 2235 956 2239
rect 1278 2239 1279 2243
rect 1284 2239 1285 2243
rect 1390 2241 1391 2245
rect 1395 2241 1396 2245
rect 1390 2240 1396 2241
rect 1398 2243 1405 2244
rect 1278 2238 1285 2239
rect 1398 2239 1399 2243
rect 1404 2239 1405 2243
rect 1398 2238 1405 2239
rect 1630 2241 1636 2242
rect 1630 2237 1631 2241
rect 1635 2237 1636 2241
rect 1630 2236 1636 2237
rect 950 2234 956 2235
rect 1670 2235 1676 2236
rect 1670 2231 1671 2235
rect 1675 2231 1676 2235
rect 1670 2230 1676 2231
rect 3190 2235 3196 2236
rect 3190 2231 3191 2235
rect 3195 2231 3196 2235
rect 3190 2230 3196 2231
rect 2014 2228 2020 2229
rect 2014 2224 2015 2228
rect 2019 2224 2020 2228
rect 110 2223 116 2224
rect 110 2219 111 2223
rect 115 2219 116 2223
rect 110 2218 116 2219
rect 1630 2223 1636 2224
rect 2014 2223 2020 2224
rect 2166 2228 2172 2229
rect 2166 2224 2167 2228
rect 2171 2224 2172 2228
rect 2166 2223 2172 2224
rect 2318 2228 2324 2229
rect 2318 2224 2319 2228
rect 2323 2224 2324 2228
rect 2318 2223 2324 2224
rect 2462 2228 2468 2229
rect 2462 2224 2463 2228
rect 2467 2224 2468 2228
rect 2462 2223 2468 2224
rect 2606 2228 2612 2229
rect 2606 2224 2607 2228
rect 2611 2224 2612 2228
rect 2606 2223 2612 2224
rect 2758 2228 2764 2229
rect 2758 2224 2759 2228
rect 2763 2224 2764 2228
rect 2758 2223 2764 2224
rect 1630 2219 1631 2223
rect 1635 2219 1636 2223
rect 1630 2218 1636 2219
rect 550 2216 556 2217
rect 550 2212 551 2216
rect 555 2212 556 2216
rect 550 2211 556 2212
rect 678 2216 684 2217
rect 678 2212 679 2216
rect 683 2212 684 2216
rect 678 2211 684 2212
rect 806 2216 812 2217
rect 806 2212 807 2216
rect 811 2212 812 2216
rect 806 2211 812 2212
rect 926 2216 932 2217
rect 926 2212 927 2216
rect 931 2212 932 2216
rect 926 2211 932 2212
rect 1046 2216 1052 2217
rect 1046 2212 1047 2216
rect 1051 2212 1052 2216
rect 1046 2211 1052 2212
rect 1158 2216 1164 2217
rect 1158 2212 1159 2216
rect 1163 2212 1164 2216
rect 1158 2211 1164 2212
rect 1270 2216 1276 2217
rect 1270 2212 1271 2216
rect 1275 2212 1276 2216
rect 1270 2211 1276 2212
rect 1390 2216 1396 2217
rect 1390 2212 1391 2216
rect 1395 2212 1396 2216
rect 1390 2211 1396 2212
rect 1926 2212 1932 2213
rect 1926 2208 1927 2212
rect 1931 2208 1932 2212
rect 1926 2207 1932 2208
rect 2102 2212 2108 2213
rect 2102 2208 2103 2212
rect 2107 2208 2108 2212
rect 2102 2207 2108 2208
rect 2294 2212 2300 2213
rect 2294 2208 2295 2212
rect 2299 2208 2300 2212
rect 2294 2207 2300 2208
rect 2502 2212 2508 2213
rect 2502 2208 2503 2212
rect 2507 2208 2508 2212
rect 2502 2207 2508 2208
rect 2718 2212 2724 2213
rect 2718 2208 2719 2212
rect 2723 2208 2724 2212
rect 2718 2207 2724 2208
rect 2950 2212 2956 2213
rect 2950 2208 2951 2212
rect 2955 2208 2956 2212
rect 2950 2207 2956 2208
rect 3158 2212 3164 2213
rect 3158 2208 3159 2212
rect 3163 2208 3164 2212
rect 3158 2207 3164 2208
rect 1670 2205 1676 2206
rect 1670 2201 1671 2205
rect 1675 2201 1676 2205
rect 1670 2200 1676 2201
rect 3190 2205 3196 2206
rect 3190 2201 3191 2205
rect 3195 2201 3196 2205
rect 3190 2200 3196 2201
rect 454 2196 460 2197
rect 454 2192 455 2196
rect 459 2192 460 2196
rect 454 2191 460 2192
rect 582 2196 588 2197
rect 582 2192 583 2196
rect 587 2192 588 2196
rect 582 2191 588 2192
rect 702 2196 708 2197
rect 702 2192 703 2196
rect 707 2192 708 2196
rect 702 2191 708 2192
rect 822 2196 828 2197
rect 822 2192 823 2196
rect 827 2192 828 2196
rect 822 2191 828 2192
rect 942 2196 948 2197
rect 942 2192 943 2196
rect 947 2192 948 2196
rect 942 2191 948 2192
rect 1054 2196 1060 2197
rect 1054 2192 1055 2196
rect 1059 2192 1060 2196
rect 1054 2191 1060 2192
rect 1166 2196 1172 2197
rect 1166 2192 1167 2196
rect 1171 2192 1172 2196
rect 1166 2191 1172 2192
rect 1286 2196 1292 2197
rect 1286 2192 1287 2196
rect 1291 2192 1292 2196
rect 1286 2191 1292 2192
rect 2022 2195 2028 2196
rect 2022 2191 2023 2195
rect 2027 2194 2028 2195
rect 2027 2192 2118 2194
rect 2027 2191 2028 2192
rect 2022 2190 2028 2191
rect 2116 2191 2124 2192
rect 2116 2190 2119 2191
rect 110 2189 116 2190
rect 110 2185 111 2189
rect 115 2185 116 2189
rect 110 2184 116 2185
rect 1630 2189 1636 2190
rect 1630 2185 1631 2189
rect 1635 2185 1636 2189
rect 2111 2189 2119 2190
rect 1630 2184 1636 2185
rect 1670 2187 1676 2188
rect 1670 2183 1671 2187
rect 1675 2183 1676 2187
rect 2111 2185 2112 2189
rect 2116 2187 2119 2189
rect 2123 2190 2124 2191
rect 2174 2191 2180 2192
rect 2174 2190 2175 2191
rect 2123 2188 2175 2190
rect 2123 2187 2124 2188
rect 2116 2186 2124 2187
rect 2174 2187 2175 2188
rect 2179 2187 2180 2191
rect 2174 2186 2180 2187
rect 2726 2187 2733 2188
rect 2116 2185 2117 2186
rect 2111 2184 2117 2185
rect 1670 2182 1676 2183
rect 1926 2183 1932 2184
rect 1926 2179 1927 2183
rect 1931 2179 1932 2183
rect 1926 2178 1932 2179
rect 1935 2183 1941 2184
rect 1935 2179 1936 2183
rect 1940 2182 1941 2183
rect 2022 2183 2028 2184
rect 2022 2182 2023 2183
rect 1940 2180 2023 2182
rect 1940 2179 1941 2180
rect 1935 2178 1941 2179
rect 2022 2179 2023 2180
rect 2027 2179 2028 2183
rect 2022 2178 2028 2179
rect 2102 2183 2108 2184
rect 2102 2179 2103 2183
rect 2107 2179 2108 2183
rect 2102 2178 2108 2179
rect 2294 2183 2300 2184
rect 2294 2179 2295 2183
rect 2299 2179 2300 2183
rect 2294 2178 2300 2179
rect 2302 2183 2309 2184
rect 2302 2179 2303 2183
rect 2308 2179 2309 2183
rect 2302 2178 2309 2179
rect 2502 2183 2508 2184
rect 2502 2179 2503 2183
rect 2507 2179 2508 2183
rect 2502 2178 2508 2179
rect 2511 2183 2517 2184
rect 2511 2179 2512 2183
rect 2516 2182 2517 2183
rect 2614 2183 2620 2184
rect 2614 2182 2615 2183
rect 2516 2180 2615 2182
rect 2516 2179 2517 2180
rect 2511 2178 2517 2179
rect 1278 2175 1284 2176
rect 110 2171 116 2172
rect 110 2167 111 2171
rect 115 2167 116 2171
rect 1062 2171 1069 2172
rect 110 2166 116 2167
rect 454 2167 460 2168
rect 454 2163 455 2167
rect 459 2163 460 2167
rect 454 2162 460 2163
rect 462 2167 469 2168
rect 462 2163 463 2167
rect 468 2163 469 2167
rect 462 2162 469 2163
rect 582 2167 588 2168
rect 582 2163 583 2167
rect 587 2163 588 2167
rect 582 2162 588 2163
rect 591 2167 597 2168
rect 591 2163 592 2167
rect 596 2166 597 2167
rect 606 2167 612 2168
rect 606 2166 607 2167
rect 596 2164 607 2166
rect 596 2163 597 2164
rect 591 2162 597 2163
rect 606 2163 607 2164
rect 611 2163 612 2167
rect 606 2162 612 2163
rect 702 2167 708 2168
rect 702 2163 703 2167
rect 707 2163 708 2167
rect 702 2162 708 2163
rect 710 2167 717 2168
rect 710 2163 711 2167
rect 716 2163 717 2167
rect 710 2162 717 2163
rect 822 2167 828 2168
rect 822 2163 823 2167
rect 827 2163 828 2167
rect 822 2162 828 2163
rect 831 2167 837 2168
rect 831 2163 832 2167
rect 836 2166 837 2167
rect 862 2167 868 2168
rect 862 2166 863 2167
rect 836 2164 863 2166
rect 836 2163 837 2164
rect 831 2162 837 2163
rect 862 2163 863 2164
rect 867 2163 868 2167
rect 862 2162 868 2163
rect 942 2167 948 2168
rect 942 2163 943 2167
rect 947 2163 948 2167
rect 942 2162 948 2163
rect 950 2167 957 2168
rect 950 2163 951 2167
rect 956 2166 957 2167
rect 974 2167 980 2168
rect 974 2166 975 2167
rect 956 2164 975 2166
rect 956 2163 957 2164
rect 950 2162 957 2163
rect 974 2163 975 2164
rect 979 2163 980 2167
rect 974 2162 980 2163
rect 1054 2167 1060 2168
rect 1054 2163 1055 2167
rect 1059 2163 1060 2167
rect 1062 2167 1063 2171
rect 1068 2167 1069 2171
rect 1174 2171 1181 2172
rect 1062 2166 1069 2167
rect 1166 2167 1172 2168
rect 1054 2162 1060 2163
rect 1166 2163 1167 2167
rect 1171 2163 1172 2167
rect 1174 2167 1175 2171
rect 1180 2167 1181 2171
rect 1278 2171 1279 2175
rect 1283 2174 1284 2175
rect 1283 2172 1298 2174
rect 1846 2173 1852 2174
rect 1283 2171 1284 2172
rect 1278 2170 1284 2171
rect 1295 2171 1301 2172
rect 1174 2166 1181 2167
rect 1286 2167 1292 2168
rect 1166 2162 1172 2163
rect 1286 2163 1287 2167
rect 1291 2163 1292 2167
rect 1295 2167 1296 2171
rect 1300 2167 1301 2171
rect 1295 2166 1301 2167
rect 1630 2171 1636 2172
rect 1630 2167 1631 2171
rect 1635 2167 1636 2171
rect 1630 2166 1636 2167
rect 1670 2169 1676 2170
rect 1670 2165 1671 2169
rect 1675 2165 1676 2169
rect 1846 2169 1847 2173
rect 1851 2169 1852 2173
rect 1846 2168 1852 2169
rect 1855 2171 1861 2172
rect 1855 2167 1856 2171
rect 1860 2170 1861 2171
rect 1936 2170 1938 2178
rect 1860 2168 1938 2170
rect 1998 2173 2004 2174
rect 1998 2169 1999 2173
rect 2003 2169 2004 2173
rect 2150 2173 2156 2174
rect 1998 2168 2004 2169
rect 2007 2171 2013 2172
rect 1860 2167 1861 2168
rect 1855 2166 1861 2167
rect 2007 2167 2008 2171
rect 2012 2170 2013 2171
rect 2022 2171 2028 2172
rect 2022 2170 2023 2171
rect 2012 2168 2023 2170
rect 2012 2167 2013 2168
rect 2007 2166 2013 2167
rect 2022 2167 2023 2168
rect 2027 2167 2028 2171
rect 2150 2169 2151 2173
rect 2155 2169 2156 2173
rect 2294 2173 2300 2174
rect 2150 2168 2156 2169
rect 2159 2171 2165 2172
rect 2022 2166 2028 2167
rect 2159 2167 2160 2171
rect 2164 2170 2165 2171
rect 2174 2171 2180 2172
rect 2174 2170 2175 2171
rect 2164 2168 2175 2170
rect 2164 2167 2165 2168
rect 2159 2166 2165 2167
rect 2174 2167 2175 2168
rect 2179 2167 2180 2171
rect 2294 2169 2295 2173
rect 2299 2169 2300 2173
rect 2294 2168 2300 2169
rect 2446 2173 2452 2174
rect 2446 2169 2447 2173
rect 2451 2169 2452 2173
rect 2446 2168 2452 2169
rect 2455 2171 2461 2172
rect 2174 2166 2180 2167
rect 2302 2167 2309 2168
rect 1670 2164 1676 2165
rect 1286 2162 1292 2163
rect 2302 2163 2303 2167
rect 2308 2163 2309 2167
rect 2455 2167 2456 2171
rect 2460 2170 2461 2171
rect 2470 2171 2476 2172
rect 2470 2170 2471 2171
rect 2460 2168 2471 2170
rect 2460 2167 2461 2168
rect 2455 2166 2461 2167
rect 2470 2167 2471 2168
rect 2475 2170 2476 2171
rect 2513 2170 2515 2178
rect 2475 2168 2515 2170
rect 2598 2173 2604 2174
rect 2598 2169 2599 2173
rect 2603 2169 2604 2173
rect 2609 2172 2611 2180
rect 2614 2179 2615 2180
rect 2619 2179 2620 2183
rect 2614 2178 2620 2179
rect 2718 2183 2724 2184
rect 2718 2179 2719 2183
rect 2723 2179 2724 2183
rect 2726 2183 2727 2187
rect 2732 2186 2733 2187
rect 2766 2187 2772 2188
rect 2766 2186 2767 2187
rect 2732 2184 2767 2186
rect 2732 2183 2733 2184
rect 2726 2182 2733 2183
rect 2766 2183 2767 2184
rect 2771 2183 2772 2187
rect 2958 2187 2965 2188
rect 2766 2182 2772 2183
rect 2950 2183 2956 2184
rect 2718 2178 2724 2179
rect 2950 2179 2951 2183
rect 2955 2179 2956 2183
rect 2958 2183 2959 2187
rect 2964 2186 2965 2187
rect 2990 2187 2996 2188
rect 2990 2186 2991 2187
rect 2964 2184 2991 2186
rect 2964 2183 2965 2184
rect 2958 2182 2965 2183
rect 2990 2183 2991 2184
rect 2995 2183 2996 2187
rect 3190 2187 3196 2188
rect 2990 2182 2996 2183
rect 3158 2183 3164 2184
rect 2950 2178 2956 2179
rect 3158 2179 3159 2183
rect 3163 2179 3164 2183
rect 3158 2178 3164 2179
rect 3166 2183 3173 2184
rect 3166 2179 3167 2183
rect 3172 2179 3173 2183
rect 3190 2183 3191 2187
rect 3195 2183 3196 2187
rect 3190 2182 3196 2183
rect 3166 2178 3173 2179
rect 2598 2168 2604 2169
rect 2607 2171 2613 2172
rect 2475 2167 2476 2168
rect 2470 2166 2476 2167
rect 2607 2167 2608 2171
rect 2612 2167 2613 2171
rect 2607 2166 2613 2167
rect 3190 2169 3196 2170
rect 3190 2165 3191 2169
rect 3195 2165 3196 2169
rect 3190 2164 3196 2165
rect 2302 2162 2309 2163
rect 1670 2151 1676 2152
rect 1670 2147 1671 2151
rect 1675 2147 1676 2151
rect 1670 2146 1676 2147
rect 3190 2151 3196 2152
rect 3190 2147 3191 2151
rect 3195 2147 3196 2151
rect 3190 2146 3196 2147
rect 350 2145 356 2146
rect 110 2141 116 2142
rect 110 2137 111 2141
rect 115 2137 116 2141
rect 350 2141 351 2145
rect 355 2141 356 2145
rect 350 2140 356 2141
rect 478 2145 484 2146
rect 478 2141 479 2145
rect 483 2141 484 2145
rect 478 2140 484 2141
rect 598 2145 604 2146
rect 598 2141 599 2145
rect 603 2141 604 2145
rect 598 2140 604 2141
rect 718 2145 724 2146
rect 718 2141 719 2145
rect 723 2141 724 2145
rect 718 2140 724 2141
rect 838 2145 844 2146
rect 838 2141 839 2145
rect 843 2141 844 2145
rect 838 2140 844 2141
rect 950 2145 956 2146
rect 950 2141 951 2145
rect 955 2141 956 2145
rect 950 2140 956 2141
rect 1062 2145 1068 2146
rect 1062 2141 1063 2145
rect 1067 2141 1068 2145
rect 1062 2140 1068 2141
rect 1182 2145 1188 2146
rect 1182 2141 1183 2145
rect 1187 2141 1188 2145
rect 1846 2144 1852 2145
rect 1182 2140 1188 2141
rect 1630 2141 1636 2142
rect 110 2136 116 2137
rect 359 2139 365 2140
rect 359 2135 360 2139
rect 364 2138 365 2139
rect 382 2139 388 2140
rect 382 2138 383 2139
rect 364 2136 383 2138
rect 364 2135 365 2136
rect 359 2134 365 2135
rect 382 2135 383 2136
rect 387 2138 388 2139
rect 462 2139 468 2140
rect 462 2138 463 2139
rect 387 2136 463 2138
rect 387 2135 388 2136
rect 382 2134 388 2135
rect 462 2135 463 2136
rect 467 2138 468 2139
rect 487 2139 493 2140
rect 487 2138 488 2139
rect 467 2136 488 2138
rect 467 2135 468 2136
rect 462 2134 468 2135
rect 487 2135 488 2136
rect 492 2135 493 2139
rect 487 2134 493 2135
rect 606 2139 613 2140
rect 606 2135 607 2139
rect 612 2138 613 2139
rect 710 2139 716 2140
rect 710 2138 711 2139
rect 612 2136 711 2138
rect 612 2135 613 2136
rect 606 2134 613 2135
rect 710 2135 711 2136
rect 715 2138 716 2139
rect 727 2139 733 2140
rect 727 2138 728 2139
rect 715 2136 728 2138
rect 715 2135 716 2136
rect 710 2134 716 2135
rect 727 2135 728 2136
rect 732 2135 733 2139
rect 727 2134 733 2135
rect 847 2139 853 2140
rect 847 2135 848 2139
rect 852 2138 853 2139
rect 862 2139 868 2140
rect 862 2138 863 2139
rect 852 2136 863 2138
rect 852 2135 853 2136
rect 847 2134 853 2135
rect 862 2135 863 2136
rect 867 2135 868 2139
rect 862 2134 868 2135
rect 959 2139 965 2140
rect 959 2135 960 2139
rect 964 2138 965 2139
rect 974 2139 980 2140
rect 974 2138 975 2139
rect 964 2136 975 2138
rect 964 2135 965 2136
rect 959 2134 965 2135
rect 974 2135 975 2136
rect 979 2138 980 2139
rect 1070 2139 1077 2140
rect 1070 2138 1071 2139
rect 979 2136 1071 2138
rect 979 2135 980 2136
rect 974 2134 980 2135
rect 1070 2135 1071 2136
rect 1076 2135 1077 2139
rect 1070 2134 1077 2135
rect 1174 2139 1180 2140
rect 1174 2135 1175 2139
rect 1179 2138 1180 2139
rect 1191 2139 1197 2140
rect 1191 2138 1192 2139
rect 1179 2136 1192 2138
rect 1179 2135 1180 2136
rect 1174 2134 1180 2135
rect 1191 2135 1192 2136
rect 1196 2135 1197 2139
rect 1630 2137 1631 2141
rect 1635 2137 1636 2141
rect 1846 2140 1847 2144
rect 1851 2140 1852 2144
rect 1846 2139 1852 2140
rect 1998 2144 2004 2145
rect 1998 2140 1999 2144
rect 2003 2140 2004 2144
rect 1998 2139 2004 2140
rect 2150 2144 2156 2145
rect 2150 2140 2151 2144
rect 2155 2140 2156 2144
rect 2150 2139 2156 2140
rect 2294 2144 2300 2145
rect 2294 2140 2295 2144
rect 2299 2140 2300 2144
rect 2294 2139 2300 2140
rect 2446 2144 2452 2145
rect 2446 2140 2447 2144
rect 2451 2140 2452 2144
rect 2446 2139 2452 2140
rect 2598 2144 2604 2145
rect 2598 2140 2599 2144
rect 2603 2140 2604 2144
rect 2598 2139 2604 2140
rect 1630 2136 1636 2137
rect 1191 2134 1197 2135
rect 1758 2128 1764 2129
rect 1758 2124 1759 2128
rect 1763 2124 1764 2128
rect 110 2123 116 2124
rect 110 2119 111 2123
rect 115 2119 116 2123
rect 110 2118 116 2119
rect 1630 2123 1636 2124
rect 1758 2123 1764 2124
rect 1910 2128 1916 2129
rect 1910 2124 1911 2128
rect 1915 2124 1916 2128
rect 1910 2123 1916 2124
rect 2070 2128 2076 2129
rect 2070 2124 2071 2128
rect 2075 2124 2076 2128
rect 2070 2123 2076 2124
rect 2254 2128 2260 2129
rect 2254 2124 2255 2128
rect 2259 2124 2260 2128
rect 2254 2123 2260 2124
rect 2462 2128 2468 2129
rect 2462 2124 2463 2128
rect 2467 2124 2468 2128
rect 2462 2123 2468 2124
rect 2686 2128 2692 2129
rect 2686 2124 2687 2128
rect 2691 2124 2692 2128
rect 2686 2123 2692 2124
rect 2926 2128 2932 2129
rect 2926 2124 2927 2128
rect 2931 2124 2932 2128
rect 2926 2123 2932 2124
rect 3158 2128 3164 2129
rect 3158 2124 3159 2128
rect 3163 2124 3164 2128
rect 3158 2123 3164 2124
rect 1630 2119 1631 2123
rect 1635 2119 1636 2123
rect 1630 2118 1636 2119
rect 1670 2121 1676 2122
rect 1670 2117 1671 2121
rect 1675 2117 1676 2121
rect 350 2116 356 2117
rect 350 2112 351 2116
rect 355 2112 356 2116
rect 350 2111 356 2112
rect 478 2116 484 2117
rect 478 2112 479 2116
rect 483 2112 484 2116
rect 478 2111 484 2112
rect 598 2116 604 2117
rect 598 2112 599 2116
rect 603 2112 604 2116
rect 598 2111 604 2112
rect 718 2116 724 2117
rect 718 2112 719 2116
rect 723 2112 724 2116
rect 718 2111 724 2112
rect 838 2116 844 2117
rect 838 2112 839 2116
rect 843 2112 844 2116
rect 838 2111 844 2112
rect 950 2116 956 2117
rect 950 2112 951 2116
rect 955 2112 956 2116
rect 950 2111 956 2112
rect 1062 2116 1068 2117
rect 1062 2112 1063 2116
rect 1067 2112 1068 2116
rect 1062 2111 1068 2112
rect 1182 2116 1188 2117
rect 1670 2116 1676 2117
rect 3190 2121 3196 2122
rect 3190 2117 3191 2121
rect 3195 2117 3196 2121
rect 3190 2116 3196 2117
rect 1182 2112 1183 2116
rect 1187 2112 1188 2116
rect 1182 2111 1188 2112
rect 1670 2103 1676 2104
rect 1670 2099 1671 2103
rect 1675 2099 1676 2103
rect 2079 2103 2085 2104
rect 1670 2098 1676 2099
rect 1758 2099 1764 2100
rect 1758 2095 1759 2099
rect 1763 2095 1764 2099
rect 1758 2094 1764 2095
rect 1767 2099 1773 2100
rect 1767 2095 1768 2099
rect 1772 2098 1773 2099
rect 1910 2099 1916 2100
rect 1772 2096 1834 2098
rect 1772 2095 1773 2096
rect 1767 2094 1773 2095
rect 246 2092 252 2093
rect 246 2088 247 2092
rect 251 2088 252 2092
rect 246 2087 252 2088
rect 374 2092 380 2093
rect 374 2088 375 2092
rect 379 2088 380 2092
rect 374 2087 380 2088
rect 502 2092 508 2093
rect 502 2088 503 2092
rect 507 2088 508 2092
rect 502 2087 508 2088
rect 622 2092 628 2093
rect 622 2088 623 2092
rect 627 2088 628 2092
rect 622 2087 628 2088
rect 742 2092 748 2093
rect 742 2088 743 2092
rect 747 2088 748 2092
rect 742 2087 748 2088
rect 854 2092 860 2093
rect 854 2088 855 2092
rect 859 2088 860 2092
rect 854 2087 860 2088
rect 966 2092 972 2093
rect 966 2088 967 2092
rect 971 2088 972 2092
rect 966 2087 972 2088
rect 1086 2092 1092 2093
rect 1086 2088 1087 2092
rect 1091 2088 1092 2092
rect 1086 2087 1092 2088
rect 1694 2089 1700 2090
rect 110 2085 116 2086
rect 110 2081 111 2085
rect 115 2081 116 2085
rect 110 2080 116 2081
rect 1630 2085 1636 2086
rect 1630 2081 1631 2085
rect 1635 2081 1636 2085
rect 1630 2080 1636 2081
rect 1670 2085 1676 2086
rect 1670 2081 1671 2085
rect 1675 2081 1676 2085
rect 1694 2085 1695 2089
rect 1699 2085 1700 2089
rect 1694 2084 1700 2085
rect 1822 2089 1828 2090
rect 1822 2085 1823 2089
rect 1827 2085 1828 2089
rect 1832 2088 1834 2096
rect 1910 2095 1911 2099
rect 1915 2095 1916 2099
rect 1910 2094 1916 2095
rect 1919 2099 1925 2100
rect 1919 2095 1920 2099
rect 1924 2098 1925 2099
rect 2070 2099 2076 2100
rect 1924 2096 1978 2098
rect 1924 2095 1925 2096
rect 1919 2094 1925 2095
rect 1822 2084 1828 2085
rect 1831 2087 1837 2088
rect 1670 2080 1676 2081
rect 1702 2083 1709 2084
rect 1702 2079 1703 2083
rect 1708 2079 1709 2083
rect 1831 2083 1832 2087
rect 1836 2086 1837 2087
rect 1920 2086 1922 2094
rect 1836 2084 1922 2086
rect 1966 2089 1972 2090
rect 1966 2085 1967 2089
rect 1971 2085 1972 2089
rect 1976 2088 1978 2096
rect 2070 2095 2071 2099
rect 2075 2095 2076 2099
rect 2079 2099 2080 2103
rect 2084 2102 2085 2103
rect 2118 2103 2124 2104
rect 2118 2102 2119 2103
rect 2084 2100 2119 2102
rect 2084 2099 2085 2100
rect 2079 2098 2085 2099
rect 2118 2099 2119 2100
rect 2123 2099 2124 2103
rect 2470 2103 2477 2104
rect 2118 2098 2124 2099
rect 2254 2099 2260 2100
rect 2070 2094 2076 2095
rect 2254 2095 2255 2099
rect 2259 2095 2260 2099
rect 2254 2094 2260 2095
rect 2263 2099 2269 2100
rect 2263 2095 2264 2099
rect 2268 2098 2269 2099
rect 2302 2099 2308 2100
rect 2302 2098 2303 2099
rect 2268 2096 2303 2098
rect 2268 2095 2269 2096
rect 2263 2094 2269 2095
rect 2302 2095 2303 2096
rect 2307 2095 2308 2099
rect 2302 2094 2308 2095
rect 2462 2099 2468 2100
rect 2462 2095 2463 2099
rect 2467 2095 2468 2099
rect 2470 2099 2471 2103
rect 2476 2099 2477 2103
rect 2695 2103 2701 2104
rect 2470 2098 2477 2099
rect 2686 2099 2692 2100
rect 2462 2094 2468 2095
rect 2686 2095 2687 2099
rect 2691 2095 2692 2099
rect 2695 2099 2696 2103
rect 2700 2102 2701 2103
rect 2726 2103 2732 2104
rect 2726 2102 2727 2103
rect 2700 2100 2727 2102
rect 2700 2099 2701 2100
rect 2695 2098 2701 2099
rect 2726 2099 2727 2100
rect 2731 2099 2732 2103
rect 2935 2103 2941 2104
rect 2726 2098 2732 2099
rect 2926 2099 2932 2100
rect 2686 2094 2692 2095
rect 2926 2095 2927 2099
rect 2931 2095 2932 2099
rect 2935 2099 2936 2103
rect 2940 2102 2941 2103
rect 2958 2103 2964 2104
rect 2958 2102 2959 2103
rect 2940 2100 2959 2102
rect 2940 2099 2941 2100
rect 2935 2098 2941 2099
rect 2958 2099 2959 2100
rect 2963 2099 2964 2103
rect 3190 2103 3196 2104
rect 2958 2098 2964 2099
rect 3158 2099 3164 2100
rect 2926 2094 2932 2095
rect 3158 2095 3159 2099
rect 3163 2095 3164 2099
rect 3158 2094 3164 2095
rect 3166 2099 3173 2100
rect 3166 2095 3167 2099
rect 3172 2095 3173 2099
rect 3190 2099 3191 2103
rect 3195 2099 3196 2103
rect 3190 2098 3196 2099
rect 3166 2094 3173 2095
rect 2110 2089 2116 2090
rect 1966 2084 1972 2085
rect 1975 2087 1981 2088
rect 1836 2083 1837 2084
rect 1831 2082 1837 2083
rect 1975 2083 1976 2087
rect 1980 2086 1981 2087
rect 2022 2087 2028 2088
rect 2022 2086 2023 2087
rect 1980 2084 2023 2086
rect 1980 2083 1981 2084
rect 1975 2082 1981 2083
rect 2022 2083 2023 2084
rect 2027 2083 2028 2087
rect 2110 2085 2111 2089
rect 2115 2085 2116 2089
rect 2254 2089 2260 2090
rect 2110 2084 2116 2085
rect 2118 2087 2125 2088
rect 2022 2082 2028 2083
rect 2118 2083 2119 2087
rect 2124 2083 2125 2087
rect 2254 2085 2255 2089
rect 2259 2085 2260 2089
rect 2254 2084 2260 2085
rect 2265 2084 2267 2094
rect 2406 2089 2412 2090
rect 2406 2085 2407 2089
rect 2411 2085 2412 2089
rect 2406 2084 2412 2085
rect 2414 2087 2421 2088
rect 2118 2082 2125 2083
rect 2246 2083 2252 2084
rect 1702 2078 1709 2079
rect 2246 2079 2247 2083
rect 2251 2082 2252 2083
rect 2263 2083 2269 2084
rect 2263 2082 2264 2083
rect 2251 2080 2264 2082
rect 2251 2079 2252 2080
rect 2246 2078 2252 2079
rect 2263 2079 2264 2080
rect 2268 2079 2269 2083
rect 2414 2083 2415 2087
rect 2420 2086 2421 2087
rect 2470 2087 2476 2088
rect 2470 2086 2471 2087
rect 2420 2084 2471 2086
rect 2420 2083 2421 2084
rect 2414 2082 2421 2083
rect 2470 2083 2471 2084
rect 2475 2083 2476 2087
rect 2470 2082 2476 2083
rect 3190 2085 3196 2086
rect 3190 2081 3191 2085
rect 3195 2081 3196 2085
rect 3190 2080 3196 2081
rect 2263 2078 2269 2079
rect 606 2071 612 2072
rect 606 2070 607 2071
rect 568 2068 607 2070
rect 110 2067 116 2068
rect 110 2063 111 2067
rect 115 2063 116 2067
rect 568 2064 570 2068
rect 606 2067 607 2068
rect 611 2070 612 2071
rect 1070 2071 1076 2072
rect 611 2068 635 2070
rect 611 2067 612 2068
rect 606 2066 612 2067
rect 631 2067 637 2068
rect 110 2062 116 2063
rect 246 2063 252 2064
rect 246 2059 247 2063
rect 251 2059 252 2063
rect 246 2058 252 2059
rect 254 2063 261 2064
rect 254 2059 255 2063
rect 260 2059 261 2063
rect 254 2058 261 2059
rect 374 2063 380 2064
rect 374 2059 375 2063
rect 379 2059 380 2063
rect 374 2058 380 2059
rect 382 2063 389 2064
rect 382 2059 383 2063
rect 388 2059 389 2063
rect 382 2058 389 2059
rect 502 2063 508 2064
rect 502 2059 503 2063
rect 507 2059 508 2063
rect 502 2058 508 2059
rect 511 2063 517 2064
rect 511 2059 512 2063
rect 516 2062 517 2063
rect 566 2063 572 2064
rect 566 2062 567 2063
rect 516 2060 567 2062
rect 516 2059 517 2060
rect 511 2058 517 2059
rect 566 2059 567 2060
rect 571 2059 572 2063
rect 566 2058 572 2059
rect 622 2063 628 2064
rect 622 2059 623 2063
rect 627 2059 628 2063
rect 631 2063 632 2067
rect 636 2063 637 2067
rect 1070 2067 1071 2071
rect 1075 2070 1076 2071
rect 1075 2068 1098 2070
rect 1075 2067 1076 2068
rect 1070 2066 1076 2067
rect 1095 2067 1101 2068
rect 631 2062 637 2063
rect 742 2063 748 2064
rect 622 2058 628 2059
rect 742 2059 743 2063
rect 747 2059 748 2063
rect 742 2058 748 2059
rect 751 2063 757 2064
rect 751 2059 752 2063
rect 756 2062 757 2063
rect 766 2063 772 2064
rect 766 2062 767 2063
rect 756 2060 767 2062
rect 756 2059 757 2060
rect 751 2058 757 2059
rect 766 2059 767 2060
rect 771 2059 772 2063
rect 766 2058 772 2059
rect 854 2063 860 2064
rect 854 2059 855 2063
rect 859 2059 860 2063
rect 854 2058 860 2059
rect 862 2063 869 2064
rect 862 2059 863 2063
rect 868 2059 869 2063
rect 862 2058 869 2059
rect 966 2063 972 2064
rect 966 2059 967 2063
rect 971 2059 972 2063
rect 966 2058 972 2059
rect 974 2063 981 2064
rect 974 2059 975 2063
rect 980 2059 981 2063
rect 974 2058 981 2059
rect 1086 2063 1092 2064
rect 1086 2059 1087 2063
rect 1091 2059 1092 2063
rect 1095 2063 1096 2067
rect 1100 2066 1101 2067
rect 1190 2067 1196 2068
rect 1190 2066 1191 2067
rect 1100 2064 1191 2066
rect 1100 2063 1101 2064
rect 1095 2062 1101 2063
rect 1190 2063 1191 2064
rect 1195 2063 1196 2067
rect 1190 2062 1196 2063
rect 1630 2067 1636 2068
rect 1630 2063 1631 2067
rect 1635 2063 1636 2067
rect 1630 2062 1636 2063
rect 1670 2067 1676 2068
rect 1670 2063 1671 2067
rect 1675 2063 1676 2067
rect 1670 2062 1676 2063
rect 3190 2067 3196 2068
rect 3190 2063 3191 2067
rect 3195 2063 3196 2067
rect 3190 2062 3196 2063
rect 1086 2058 1092 2059
rect 1694 2060 1700 2061
rect 1694 2056 1695 2060
rect 1699 2056 1700 2060
rect 1694 2055 1700 2056
rect 1822 2060 1828 2061
rect 1822 2056 1823 2060
rect 1827 2056 1828 2060
rect 1822 2055 1828 2056
rect 1966 2060 1972 2061
rect 1966 2056 1967 2060
rect 1971 2056 1972 2060
rect 1966 2055 1972 2056
rect 2110 2060 2116 2061
rect 2110 2056 2111 2060
rect 2115 2056 2116 2060
rect 2110 2055 2116 2056
rect 2254 2060 2260 2061
rect 2254 2056 2255 2060
rect 2259 2056 2260 2060
rect 2254 2055 2260 2056
rect 2406 2060 2412 2061
rect 2406 2056 2407 2060
rect 2411 2056 2412 2060
rect 2406 2055 2412 2056
rect 1694 2048 1700 2049
rect 174 2045 180 2046
rect 110 2041 116 2042
rect 110 2037 111 2041
rect 115 2037 116 2041
rect 174 2041 175 2045
rect 179 2041 180 2045
rect 174 2040 180 2041
rect 366 2045 372 2046
rect 366 2041 367 2045
rect 371 2041 372 2045
rect 366 2040 372 2041
rect 558 2045 564 2046
rect 558 2041 559 2045
rect 563 2041 564 2045
rect 558 2040 564 2041
rect 758 2045 764 2046
rect 758 2041 759 2045
rect 763 2041 764 2045
rect 758 2040 764 2041
rect 966 2045 972 2046
rect 966 2041 967 2045
rect 971 2041 972 2045
rect 966 2040 972 2041
rect 1182 2045 1188 2046
rect 1182 2041 1183 2045
rect 1187 2041 1188 2045
rect 1398 2045 1404 2046
rect 1182 2040 1188 2041
rect 1190 2043 1197 2044
rect 110 2036 116 2037
rect 182 2039 189 2040
rect 182 2035 183 2039
rect 188 2035 189 2039
rect 182 2034 189 2035
rect 375 2039 381 2040
rect 375 2035 376 2039
rect 380 2035 381 2039
rect 375 2034 381 2035
rect 566 2039 573 2040
rect 566 2035 567 2039
rect 572 2035 573 2039
rect 566 2034 573 2035
rect 766 2039 773 2040
rect 766 2035 767 2039
rect 772 2035 773 2039
rect 766 2034 773 2035
rect 918 2039 924 2040
rect 918 2035 919 2039
rect 923 2038 924 2039
rect 974 2039 981 2040
rect 974 2038 975 2039
rect 923 2036 975 2038
rect 923 2035 924 2036
rect 918 2034 924 2035
rect 974 2035 975 2036
rect 980 2035 981 2039
rect 1190 2039 1191 2043
rect 1196 2039 1197 2043
rect 1398 2041 1399 2045
rect 1403 2041 1404 2045
rect 1398 2040 1404 2041
rect 1598 2045 1604 2046
rect 1598 2041 1599 2045
rect 1603 2041 1604 2045
rect 1694 2044 1695 2048
rect 1699 2044 1700 2048
rect 1694 2043 1700 2044
rect 2038 2048 2044 2049
rect 2038 2044 2039 2048
rect 2043 2044 2044 2048
rect 2038 2043 2044 2044
rect 2406 2048 2412 2049
rect 2406 2044 2407 2048
rect 2411 2044 2412 2048
rect 2406 2043 2412 2044
rect 2766 2048 2772 2049
rect 2766 2044 2767 2048
rect 2771 2044 2772 2048
rect 2766 2043 2772 2044
rect 3134 2048 3140 2049
rect 3134 2044 3135 2048
rect 3139 2044 3140 2048
rect 3134 2043 3140 2044
rect 1598 2040 1604 2041
rect 1630 2041 1636 2042
rect 1190 2038 1197 2039
rect 1407 2039 1416 2040
rect 974 2034 981 2035
rect 1407 2035 1408 2039
rect 1415 2035 1416 2039
rect 1407 2034 1416 2035
rect 1607 2039 1613 2040
rect 1607 2035 1608 2039
rect 1612 2038 1613 2039
rect 1612 2036 1614 2038
rect 1630 2037 1631 2041
rect 1635 2037 1636 2041
rect 1630 2036 1636 2037
rect 1670 2041 1676 2042
rect 1670 2037 1671 2041
rect 1675 2037 1676 2041
rect 1670 2036 1676 2037
rect 3190 2041 3196 2042
rect 3190 2037 3191 2041
rect 3195 2037 3196 2041
rect 3190 2036 3196 2037
rect 1612 2035 1616 2036
rect 1607 2034 1611 2035
rect 1610 2031 1611 2034
rect 1615 2034 1616 2035
rect 1702 2035 1708 2036
rect 1702 2034 1703 2035
rect 1615 2032 1703 2034
rect 1615 2031 1616 2032
rect 1610 2030 1616 2031
rect 1702 2031 1703 2032
rect 1707 2031 1708 2035
rect 1702 2030 1708 2031
rect 2022 2027 2028 2028
rect 110 2023 116 2024
rect 110 2019 111 2023
rect 115 2019 116 2023
rect 110 2018 116 2019
rect 1630 2023 1636 2024
rect 1630 2019 1631 2023
rect 1635 2019 1636 2023
rect 1630 2018 1636 2019
rect 1670 2023 1676 2024
rect 1670 2019 1671 2023
rect 1675 2019 1676 2023
rect 1702 2023 1709 2024
rect 1670 2018 1676 2019
rect 1694 2019 1700 2020
rect 174 2016 180 2017
rect 174 2012 175 2016
rect 179 2012 180 2016
rect 174 2011 180 2012
rect 366 2016 372 2017
rect 366 2012 367 2016
rect 371 2012 372 2016
rect 366 2011 372 2012
rect 558 2016 564 2017
rect 558 2012 559 2016
rect 563 2012 564 2016
rect 558 2011 564 2012
rect 758 2016 764 2017
rect 758 2012 759 2016
rect 763 2012 764 2016
rect 758 2011 764 2012
rect 966 2016 972 2017
rect 966 2012 967 2016
rect 971 2012 972 2016
rect 966 2011 972 2012
rect 1182 2016 1188 2017
rect 1182 2012 1183 2016
rect 1187 2012 1188 2016
rect 1182 2011 1188 2012
rect 1398 2016 1404 2017
rect 1398 2012 1399 2016
rect 1403 2012 1404 2016
rect 1398 2011 1404 2012
rect 1598 2016 1604 2017
rect 1598 2012 1599 2016
rect 1603 2012 1604 2016
rect 1694 2015 1695 2019
rect 1699 2015 1700 2019
rect 1702 2019 1703 2023
rect 1708 2019 1709 2023
rect 2022 2023 2023 2027
rect 2027 2026 2028 2027
rect 2726 2027 2732 2028
rect 2027 2024 2050 2026
rect 2027 2023 2028 2024
rect 2022 2022 2028 2023
rect 2047 2023 2053 2024
rect 1702 2018 1709 2019
rect 2038 2019 2044 2020
rect 1694 2014 1700 2015
rect 2038 2015 2039 2019
rect 2043 2015 2044 2019
rect 2047 2019 2048 2023
rect 2052 2019 2053 2023
rect 2414 2023 2421 2024
rect 2047 2018 2053 2019
rect 2406 2019 2412 2020
rect 2038 2014 2044 2015
rect 2406 2015 2407 2019
rect 2411 2015 2412 2019
rect 2414 2019 2415 2023
rect 2420 2019 2421 2023
rect 2726 2023 2727 2027
rect 2731 2026 2732 2027
rect 2731 2024 2779 2026
rect 2731 2023 2732 2024
rect 2726 2022 2732 2023
rect 2775 2023 2781 2024
rect 2414 2018 2421 2019
rect 2766 2019 2772 2020
rect 2406 2014 2412 2015
rect 2766 2015 2767 2019
rect 2771 2015 2772 2019
rect 2775 2019 2776 2023
rect 2780 2022 2781 2023
rect 2854 2023 2860 2024
rect 2854 2022 2855 2023
rect 2780 2020 2855 2022
rect 2780 2019 2781 2020
rect 2775 2018 2781 2019
rect 2854 2019 2855 2020
rect 2859 2019 2860 2023
rect 3190 2023 3196 2024
rect 2854 2018 2860 2019
rect 3134 2019 3140 2020
rect 2766 2014 2772 2015
rect 3134 2015 3135 2019
rect 3139 2015 3140 2019
rect 3134 2014 3140 2015
rect 3142 2019 3149 2020
rect 3142 2015 3143 2019
rect 3148 2015 3149 2019
rect 3190 2019 3191 2023
rect 3195 2019 3196 2023
rect 3190 2018 3196 2019
rect 3142 2014 3149 2015
rect 1598 2011 1604 2012
rect 134 2004 140 2005
rect 134 2000 135 2004
rect 139 2000 140 2004
rect 134 1999 140 2000
rect 230 2004 236 2005
rect 230 2000 231 2004
rect 235 2000 236 2004
rect 230 1999 236 2000
rect 350 2004 356 2005
rect 350 2000 351 2004
rect 355 2000 356 2004
rect 350 1999 356 2000
rect 462 2004 468 2005
rect 462 2000 463 2004
rect 467 2000 468 2004
rect 462 1999 468 2000
rect 574 2004 580 2005
rect 574 2000 575 2004
rect 579 2000 580 2004
rect 574 1999 580 2000
rect 686 2004 692 2005
rect 686 2000 687 2004
rect 691 2000 692 2004
rect 686 1999 692 2000
rect 798 2004 804 2005
rect 798 2000 799 2004
rect 803 2000 804 2004
rect 798 1999 804 2000
rect 910 2004 916 2005
rect 910 2000 911 2004
rect 915 2000 916 2004
rect 910 1999 916 2000
rect 2262 2001 2268 2002
rect 110 1997 116 1998
rect 110 1993 111 1997
rect 115 1993 116 1997
rect 110 1992 116 1993
rect 1630 1997 1636 1998
rect 1630 1993 1631 1997
rect 1635 1993 1636 1997
rect 1630 1992 1636 1993
rect 1670 1997 1676 1998
rect 1670 1993 1671 1997
rect 1675 1993 1676 1997
rect 2262 1997 2263 2001
rect 2267 1997 2268 2001
rect 2262 1996 2268 1997
rect 2414 2001 2420 2002
rect 2414 1997 2415 2001
rect 2419 1997 2420 2001
rect 2558 2001 2564 2002
rect 2414 1996 2420 1997
rect 2422 1999 2429 2000
rect 1670 1992 1676 1993
rect 2246 1995 2252 1996
rect 2246 1991 2247 1995
rect 2251 1994 2252 1995
rect 2271 1995 2277 1996
rect 2271 1994 2272 1995
rect 2251 1992 2272 1994
rect 2251 1991 2252 1992
rect 2246 1990 2252 1991
rect 2271 1991 2272 1992
rect 2276 1991 2277 1995
rect 2422 1995 2423 1999
rect 2428 1998 2429 1999
rect 2428 1996 2510 1998
rect 2558 1997 2559 2001
rect 2563 1997 2564 2001
rect 2558 1996 2564 1997
rect 2702 2001 2708 2002
rect 2702 1997 2703 2001
rect 2707 1997 2708 2001
rect 2838 2001 2844 2002
rect 2702 1996 2708 1997
rect 2711 1999 2717 2000
rect 2428 1995 2429 1996
rect 2422 1994 2429 1995
rect 2508 1994 2510 1996
rect 2550 1995 2556 1996
rect 2550 1994 2551 1995
rect 2508 1992 2551 1994
rect 2271 1990 2277 1991
rect 2550 1991 2551 1992
rect 2555 1994 2556 1995
rect 2567 1995 2573 1996
rect 2567 1994 2568 1995
rect 2555 1992 2568 1994
rect 2555 1991 2556 1992
rect 2550 1990 2556 1991
rect 2567 1991 2568 1992
rect 2572 1991 2573 1995
rect 2711 1995 2712 1999
rect 2716 1998 2717 1999
rect 2726 1999 2732 2000
rect 2726 1998 2727 1999
rect 2716 1996 2727 1998
rect 2716 1995 2717 1996
rect 2711 1994 2717 1995
rect 2726 1995 2727 1996
rect 2731 1995 2732 1999
rect 2838 1997 2839 2001
rect 2843 1997 2844 2001
rect 2974 2001 2980 2002
rect 2838 1996 2844 1997
rect 2847 1999 2853 2000
rect 2726 1994 2732 1995
rect 2847 1995 2848 1999
rect 2852 1998 2853 1999
rect 2852 1996 2862 1998
rect 2974 1997 2975 2001
rect 2979 1997 2980 2001
rect 2974 1996 2980 1997
rect 3110 2001 3116 2002
rect 3110 1997 3111 2001
rect 3115 1997 3116 2001
rect 3110 1996 3116 1997
rect 3190 1997 3196 1998
rect 2852 1995 2853 1996
rect 2847 1994 2853 1995
rect 2858 1995 2864 1996
rect 2567 1990 2573 1991
rect 2858 1991 2859 1995
rect 2863 1994 2864 1995
rect 2983 1995 2989 1996
rect 2983 1994 2984 1995
rect 2863 1992 2984 1994
rect 2863 1991 2864 1992
rect 2858 1990 2864 1991
rect 2983 1991 2984 1992
rect 2988 1994 2989 1995
rect 3006 1995 3012 1996
rect 3006 1994 3007 1995
rect 2988 1992 3007 1994
rect 2988 1991 2989 1992
rect 2983 1990 2989 1991
rect 3006 1991 3007 1992
rect 3011 1991 3012 1995
rect 3006 1990 3012 1991
rect 3119 1995 3125 1996
rect 3119 1991 3120 1995
rect 3124 1994 3125 1995
rect 3142 1995 3148 1996
rect 3142 1994 3143 1995
rect 3124 1992 3143 1994
rect 3124 1991 3125 1992
rect 3119 1990 3125 1991
rect 3142 1991 3143 1992
rect 3147 1994 3148 1995
rect 3166 1995 3172 1996
rect 3166 1994 3167 1995
rect 3147 1992 3167 1994
rect 3147 1991 3148 1992
rect 3142 1990 3148 1991
rect 3166 1991 3167 1992
rect 3171 1991 3172 1995
rect 3190 1993 3191 1997
rect 3195 1993 3196 1997
rect 3190 1992 3196 1993
rect 3166 1990 3172 1991
rect 182 1983 188 1984
rect 182 1982 183 1983
rect 145 1980 183 1982
rect 110 1979 116 1980
rect 110 1975 111 1979
rect 115 1975 116 1979
rect 145 1976 147 1980
rect 182 1979 183 1980
rect 187 1982 188 1983
rect 254 1983 260 1984
rect 254 1982 255 1983
rect 187 1980 255 1982
rect 187 1979 188 1980
rect 182 1978 188 1979
rect 239 1979 245 1980
rect 110 1974 116 1975
rect 134 1975 140 1976
rect 134 1971 135 1975
rect 139 1971 140 1975
rect 134 1970 140 1971
rect 142 1975 149 1976
rect 142 1971 143 1975
rect 148 1971 149 1975
rect 142 1970 149 1971
rect 230 1975 236 1976
rect 230 1971 231 1975
rect 235 1971 236 1975
rect 239 1975 240 1979
rect 244 1975 245 1979
rect 254 1979 255 1980
rect 259 1982 260 1983
rect 374 1983 380 1984
rect 374 1982 375 1983
rect 259 1980 375 1982
rect 259 1979 260 1980
rect 254 1978 260 1979
rect 359 1979 365 1980
rect 239 1974 245 1975
rect 350 1975 356 1976
rect 230 1970 236 1971
rect 350 1971 351 1975
rect 355 1971 356 1975
rect 359 1975 360 1979
rect 364 1975 365 1979
rect 374 1979 375 1980
rect 379 1982 380 1983
rect 566 1983 572 1984
rect 566 1982 567 1983
rect 379 1980 567 1982
rect 379 1979 380 1980
rect 374 1978 380 1979
rect 471 1979 477 1980
rect 359 1974 365 1975
rect 462 1975 468 1976
rect 350 1970 356 1971
rect 462 1971 463 1975
rect 467 1971 468 1975
rect 471 1975 472 1979
rect 476 1975 477 1979
rect 566 1979 567 1980
rect 571 1982 572 1983
rect 571 1980 587 1982
rect 571 1979 572 1980
rect 566 1978 572 1979
rect 583 1979 589 1980
rect 471 1974 477 1975
rect 574 1975 580 1976
rect 462 1970 468 1971
rect 574 1971 575 1975
rect 579 1971 580 1975
rect 583 1975 584 1979
rect 588 1975 589 1979
rect 1630 1979 1636 1980
rect 583 1974 589 1975
rect 686 1975 692 1976
rect 574 1970 580 1971
rect 686 1971 687 1975
rect 691 1971 692 1975
rect 686 1970 692 1971
rect 695 1975 701 1976
rect 695 1971 696 1975
rect 700 1971 701 1975
rect 695 1970 701 1971
rect 798 1975 804 1976
rect 798 1971 799 1975
rect 803 1971 804 1975
rect 798 1970 804 1971
rect 807 1975 813 1976
rect 807 1971 808 1975
rect 812 1971 813 1975
rect 807 1970 813 1971
rect 910 1975 916 1976
rect 910 1971 911 1975
rect 915 1971 916 1975
rect 910 1970 916 1971
rect 918 1975 925 1976
rect 918 1971 919 1975
rect 924 1971 925 1975
rect 1630 1975 1631 1979
rect 1635 1975 1636 1979
rect 1630 1974 1636 1975
rect 1670 1979 1676 1980
rect 1670 1975 1671 1979
rect 1675 1975 1676 1979
rect 1670 1974 1676 1975
rect 3190 1979 3196 1980
rect 3190 1975 3191 1979
rect 3195 1975 3196 1979
rect 3190 1974 3196 1975
rect 918 1970 925 1971
rect 2262 1972 2268 1973
rect 697 1966 699 1970
rect 766 1967 772 1968
rect 766 1966 767 1967
rect 697 1964 767 1966
rect 766 1963 767 1964
rect 771 1966 772 1967
rect 809 1966 811 1970
rect 2262 1968 2263 1972
rect 2267 1968 2268 1972
rect 2262 1967 2268 1968
rect 2414 1972 2420 1973
rect 2414 1968 2415 1972
rect 2419 1968 2420 1972
rect 2414 1967 2420 1968
rect 2558 1972 2564 1973
rect 2558 1968 2559 1972
rect 2563 1968 2564 1972
rect 2558 1967 2564 1968
rect 2702 1972 2708 1973
rect 2702 1968 2703 1972
rect 2707 1968 2708 1972
rect 2702 1967 2708 1968
rect 2838 1972 2844 1973
rect 2838 1968 2839 1972
rect 2843 1968 2844 1972
rect 2838 1967 2844 1968
rect 2974 1972 2980 1973
rect 2974 1968 2975 1972
rect 2979 1968 2980 1972
rect 2974 1967 2980 1968
rect 3110 1972 3116 1973
rect 3110 1968 3111 1972
rect 3115 1968 3116 1972
rect 3110 1967 3116 1968
rect 771 1964 811 1966
rect 771 1963 772 1964
rect 766 1962 772 1963
rect 809 1962 811 1964
rect 862 1963 868 1964
rect 862 1962 863 1963
rect 809 1960 863 1962
rect 862 1959 863 1960
rect 867 1959 868 1963
rect 862 1958 868 1959
rect 2238 1960 2244 1961
rect 726 1957 732 1958
rect 110 1953 116 1954
rect 110 1949 111 1953
rect 115 1949 116 1953
rect 726 1953 727 1957
rect 731 1953 732 1957
rect 726 1952 732 1953
rect 854 1957 860 1958
rect 854 1953 855 1957
rect 859 1953 860 1957
rect 865 1956 867 1958
rect 982 1957 988 1958
rect 854 1952 860 1953
rect 863 1955 869 1956
rect 110 1948 116 1949
rect 735 1951 741 1952
rect 735 1947 736 1951
rect 740 1950 741 1951
rect 766 1951 772 1952
rect 766 1950 767 1951
rect 740 1948 767 1950
rect 740 1947 741 1948
rect 735 1946 741 1947
rect 766 1947 767 1948
rect 771 1947 772 1951
rect 863 1951 864 1955
rect 868 1954 869 1955
rect 886 1955 892 1956
rect 886 1954 887 1955
rect 868 1952 887 1954
rect 868 1951 869 1952
rect 863 1950 869 1951
rect 886 1951 887 1952
rect 891 1951 892 1955
rect 982 1953 983 1957
rect 987 1953 988 1957
rect 982 1952 988 1953
rect 1102 1957 1108 1958
rect 1102 1953 1103 1957
rect 1107 1953 1108 1957
rect 1102 1952 1108 1953
rect 1222 1957 1228 1958
rect 1222 1953 1223 1957
rect 1227 1953 1228 1957
rect 1222 1952 1228 1953
rect 1334 1957 1340 1958
rect 1334 1953 1335 1957
rect 1339 1953 1340 1957
rect 1446 1957 1452 1958
rect 1334 1952 1340 1953
rect 1399 1952 1414 1954
rect 1446 1953 1447 1957
rect 1451 1953 1452 1957
rect 1446 1952 1452 1953
rect 1566 1957 1572 1958
rect 1566 1953 1567 1957
rect 1571 1953 1572 1957
rect 2238 1956 2239 1960
rect 2243 1956 2244 1960
rect 1566 1952 1572 1953
rect 1575 1955 1581 1956
rect 886 1950 892 1951
rect 918 1951 924 1952
rect 918 1950 919 1951
rect 888 1948 919 1950
rect 766 1946 772 1947
rect 918 1947 919 1948
rect 923 1950 924 1951
rect 991 1951 997 1952
rect 991 1950 992 1951
rect 923 1948 992 1950
rect 923 1947 924 1948
rect 918 1946 924 1947
rect 991 1947 992 1948
rect 996 1950 997 1951
rect 1006 1951 1012 1952
rect 1006 1950 1007 1951
rect 996 1948 1007 1950
rect 996 1947 997 1948
rect 991 1946 997 1947
rect 1006 1947 1007 1948
rect 1011 1950 1012 1951
rect 1111 1951 1117 1952
rect 1111 1950 1112 1951
rect 1011 1948 1112 1950
rect 1011 1947 1012 1948
rect 1006 1946 1012 1947
rect 1111 1947 1112 1948
rect 1116 1950 1117 1951
rect 1126 1951 1132 1952
rect 1126 1950 1127 1951
rect 1116 1948 1127 1950
rect 1116 1947 1117 1948
rect 1111 1946 1117 1947
rect 1126 1947 1127 1948
rect 1131 1950 1132 1951
rect 1231 1951 1237 1952
rect 1231 1950 1232 1951
rect 1131 1948 1232 1950
rect 1131 1947 1132 1948
rect 1126 1946 1132 1947
rect 1231 1947 1232 1948
rect 1236 1947 1237 1951
rect 1343 1951 1349 1952
rect 1231 1946 1237 1947
rect 1242 1947 1248 1948
rect 1242 1946 1243 1947
rect 1232 1944 1243 1946
rect 1242 1943 1243 1944
rect 1247 1946 1248 1947
rect 1343 1947 1344 1951
rect 1348 1947 1349 1951
rect 1343 1946 1349 1947
rect 1354 1947 1360 1948
rect 1354 1946 1355 1947
rect 1247 1944 1355 1946
rect 1247 1943 1248 1944
rect 1242 1942 1248 1943
rect 1354 1943 1355 1944
rect 1359 1946 1360 1947
rect 1399 1946 1401 1952
rect 1410 1951 1416 1952
rect 1410 1947 1411 1951
rect 1415 1950 1416 1951
rect 1455 1951 1461 1952
rect 1455 1950 1456 1951
rect 1415 1948 1456 1950
rect 1415 1947 1416 1948
rect 1410 1946 1416 1947
rect 1455 1947 1456 1948
rect 1460 1950 1461 1951
rect 1470 1951 1476 1952
rect 1470 1950 1471 1951
rect 1460 1948 1471 1950
rect 1460 1947 1461 1948
rect 1455 1946 1461 1947
rect 1470 1947 1471 1948
rect 1475 1950 1476 1951
rect 1575 1951 1576 1955
rect 1580 1954 1581 1955
rect 1610 1955 1616 1956
rect 2238 1955 2244 1956
rect 2390 1960 2396 1961
rect 2390 1956 2391 1960
rect 2395 1956 2396 1960
rect 2390 1955 2396 1956
rect 2542 1960 2548 1961
rect 2542 1956 2543 1960
rect 2547 1956 2548 1960
rect 2542 1955 2548 1956
rect 2694 1960 2700 1961
rect 2694 1956 2695 1960
rect 2699 1956 2700 1960
rect 2694 1955 2700 1956
rect 2846 1960 2852 1961
rect 2846 1956 2847 1960
rect 2851 1956 2852 1960
rect 2846 1955 2852 1956
rect 2998 1960 3004 1961
rect 2998 1956 2999 1960
rect 3003 1956 3004 1960
rect 2998 1955 3004 1956
rect 1610 1954 1611 1955
rect 1580 1952 1611 1954
rect 1580 1951 1581 1952
rect 1575 1950 1581 1951
rect 1610 1951 1611 1952
rect 1615 1951 1616 1955
rect 1610 1950 1616 1951
rect 1630 1953 1636 1954
rect 1475 1948 1578 1950
rect 1630 1949 1631 1953
rect 1635 1949 1636 1953
rect 1630 1948 1636 1949
rect 1670 1953 1676 1954
rect 1670 1949 1671 1953
rect 1675 1949 1676 1953
rect 1670 1948 1676 1949
rect 3190 1953 3196 1954
rect 3190 1949 3191 1953
rect 3195 1949 3196 1953
rect 3190 1948 3196 1949
rect 1475 1947 1476 1948
rect 1470 1946 1476 1947
rect 1359 1944 1401 1946
rect 1359 1943 1360 1944
rect 1354 1942 1360 1943
rect 110 1935 116 1936
rect 110 1931 111 1935
rect 115 1931 116 1935
rect 110 1930 116 1931
rect 1630 1935 1636 1936
rect 1630 1931 1631 1935
rect 1635 1931 1636 1935
rect 1630 1930 1636 1931
rect 1670 1935 1676 1936
rect 1670 1931 1671 1935
rect 1675 1931 1676 1935
rect 2399 1935 2405 1936
rect 1670 1930 1676 1931
rect 2238 1931 2244 1932
rect 726 1928 732 1929
rect 726 1924 727 1928
rect 731 1924 732 1928
rect 726 1923 732 1924
rect 854 1928 860 1929
rect 854 1924 855 1928
rect 859 1924 860 1928
rect 854 1923 860 1924
rect 982 1928 988 1929
rect 982 1924 983 1928
rect 987 1924 988 1928
rect 982 1923 988 1924
rect 1102 1928 1108 1929
rect 1102 1924 1103 1928
rect 1107 1924 1108 1928
rect 1102 1923 1108 1924
rect 1222 1928 1228 1929
rect 1222 1924 1223 1928
rect 1227 1924 1228 1928
rect 1222 1923 1228 1924
rect 1334 1928 1340 1929
rect 1334 1924 1335 1928
rect 1339 1924 1340 1928
rect 1334 1923 1340 1924
rect 1446 1928 1452 1929
rect 1446 1924 1447 1928
rect 1451 1924 1452 1928
rect 1446 1923 1452 1924
rect 1566 1928 1572 1929
rect 1566 1924 1567 1928
rect 1571 1924 1572 1928
rect 2238 1927 2239 1931
rect 2243 1927 2244 1931
rect 2238 1926 2244 1927
rect 2246 1931 2253 1932
rect 2246 1927 2247 1931
rect 2252 1927 2253 1931
rect 2246 1926 2253 1927
rect 2390 1931 2396 1932
rect 2390 1927 2391 1931
rect 2395 1927 2396 1931
rect 2399 1931 2400 1935
rect 2404 1934 2405 1935
rect 2422 1935 2428 1936
rect 2422 1934 2423 1935
rect 2404 1932 2423 1934
rect 2404 1931 2405 1932
rect 2399 1930 2405 1931
rect 2422 1931 2423 1932
rect 2427 1931 2428 1935
rect 2550 1935 2557 1936
rect 2422 1930 2428 1931
rect 2542 1931 2548 1932
rect 2390 1926 2396 1927
rect 2542 1927 2543 1931
rect 2547 1927 2548 1931
rect 2550 1931 2551 1935
rect 2556 1931 2557 1935
rect 2702 1935 2709 1936
rect 2550 1930 2557 1931
rect 2694 1931 2700 1932
rect 2542 1926 2548 1927
rect 2694 1927 2695 1931
rect 2699 1927 2700 1931
rect 2702 1931 2703 1935
rect 2708 1934 2709 1935
rect 2726 1935 2732 1936
rect 2726 1934 2727 1935
rect 2708 1932 2727 1934
rect 2708 1931 2709 1932
rect 2702 1930 2709 1931
rect 2726 1931 2727 1932
rect 2731 1931 2732 1935
rect 2854 1935 2861 1936
rect 2726 1930 2732 1931
rect 2846 1931 2852 1932
rect 2694 1926 2700 1927
rect 2846 1927 2847 1931
rect 2851 1927 2852 1931
rect 2854 1931 2855 1935
rect 2860 1931 2861 1935
rect 3006 1935 3013 1936
rect 2854 1930 2861 1931
rect 2998 1931 3004 1932
rect 2846 1926 2852 1927
rect 2998 1927 2999 1931
rect 3003 1927 3004 1931
rect 3006 1931 3007 1935
rect 3012 1931 3013 1935
rect 3006 1930 3013 1931
rect 3190 1935 3196 1936
rect 3190 1931 3191 1935
rect 3195 1931 3196 1935
rect 3190 1930 3196 1931
rect 2998 1926 3004 1927
rect 1566 1923 1572 1924
rect 2150 1917 2156 1918
rect 1670 1913 1676 1914
rect 1670 1909 1671 1913
rect 1675 1909 1676 1913
rect 2150 1913 2151 1917
rect 2155 1913 2156 1917
rect 2150 1912 2156 1913
rect 2310 1917 2316 1918
rect 2310 1913 2311 1917
rect 2315 1913 2316 1917
rect 2310 1912 2316 1913
rect 2470 1917 2476 1918
rect 2470 1913 2471 1917
rect 2475 1913 2476 1917
rect 2470 1912 2476 1913
rect 2638 1917 2644 1918
rect 2638 1913 2639 1917
rect 2643 1913 2644 1917
rect 2814 1917 2820 1918
rect 2638 1912 2644 1913
rect 2647 1915 2653 1916
rect 1670 1908 1676 1909
rect 2158 1911 2165 1912
rect 2158 1907 2159 1911
rect 2164 1907 2165 1911
rect 2158 1906 2165 1907
rect 2246 1911 2252 1912
rect 2246 1907 2247 1911
rect 2251 1910 2252 1911
rect 2319 1911 2325 1912
rect 2319 1910 2320 1911
rect 2251 1908 2320 1910
rect 2251 1907 2252 1908
rect 2246 1906 2252 1907
rect 2319 1907 2320 1908
rect 2324 1907 2325 1911
rect 2319 1906 2325 1907
rect 2422 1911 2428 1912
rect 2422 1907 2423 1911
rect 2427 1910 2428 1911
rect 2479 1911 2485 1912
rect 2479 1910 2480 1911
rect 2427 1908 2480 1910
rect 2427 1907 2428 1908
rect 2422 1906 2428 1907
rect 2479 1907 2480 1908
rect 2484 1907 2485 1911
rect 2647 1911 2648 1915
rect 2652 1914 2653 1915
rect 2702 1915 2708 1916
rect 2702 1914 2703 1915
rect 2652 1912 2703 1914
rect 2652 1911 2653 1912
rect 2647 1910 2653 1911
rect 2702 1911 2703 1912
rect 2707 1911 2708 1915
rect 2814 1913 2815 1917
rect 2819 1913 2820 1917
rect 2998 1917 3004 1918
rect 2814 1912 2820 1913
rect 2822 1915 2829 1916
rect 2702 1910 2708 1911
rect 2822 1911 2823 1915
rect 2828 1914 2829 1915
rect 2854 1915 2860 1916
rect 2854 1914 2855 1915
rect 2828 1912 2855 1914
rect 2828 1911 2829 1912
rect 2822 1910 2829 1911
rect 2854 1911 2855 1912
rect 2859 1911 2860 1915
rect 2998 1913 2999 1917
rect 3003 1913 3004 1917
rect 3158 1917 3164 1918
rect 2998 1912 3004 1913
rect 3006 1915 3013 1916
rect 2854 1910 2860 1911
rect 3006 1911 3007 1915
rect 3012 1911 3013 1915
rect 3158 1913 3159 1917
rect 3163 1913 3164 1917
rect 3158 1912 3164 1913
rect 3166 1915 3173 1916
rect 3006 1910 3013 1911
rect 3166 1911 3167 1915
rect 3172 1911 3173 1915
rect 3166 1910 3173 1911
rect 3190 1913 3196 1914
rect 3190 1909 3191 1913
rect 3195 1909 3196 1913
rect 3190 1908 3196 1909
rect 2479 1906 2485 1907
rect 630 1904 636 1905
rect 630 1900 631 1904
rect 635 1900 636 1904
rect 630 1899 636 1900
rect 758 1904 764 1905
rect 758 1900 759 1904
rect 763 1900 764 1904
rect 758 1899 764 1900
rect 878 1904 884 1905
rect 878 1900 879 1904
rect 883 1900 884 1904
rect 878 1899 884 1900
rect 998 1904 1004 1905
rect 998 1900 999 1904
rect 1003 1900 1004 1904
rect 998 1899 1004 1900
rect 1118 1904 1124 1905
rect 1118 1900 1119 1904
rect 1123 1900 1124 1904
rect 1118 1899 1124 1900
rect 1230 1904 1236 1905
rect 1230 1900 1231 1904
rect 1235 1900 1236 1904
rect 1230 1899 1236 1900
rect 1342 1904 1348 1905
rect 1342 1900 1343 1904
rect 1347 1900 1348 1904
rect 1342 1899 1348 1900
rect 1462 1904 1468 1905
rect 1462 1900 1463 1904
rect 1467 1900 1468 1904
rect 1462 1899 1468 1900
rect 110 1897 116 1898
rect 110 1893 111 1897
rect 115 1893 116 1897
rect 110 1892 116 1893
rect 1630 1897 1636 1898
rect 1630 1893 1631 1897
rect 1635 1893 1636 1897
rect 1630 1892 1636 1893
rect 1670 1895 1676 1896
rect 1670 1891 1671 1895
rect 1675 1891 1676 1895
rect 1670 1890 1676 1891
rect 3190 1895 3196 1896
rect 3190 1891 3191 1895
rect 3195 1891 3196 1895
rect 3190 1890 3196 1891
rect 2150 1888 2156 1889
rect 2150 1884 2151 1888
rect 2155 1884 2156 1888
rect 2150 1883 2156 1884
rect 2310 1888 2316 1889
rect 2310 1884 2311 1888
rect 2315 1884 2316 1888
rect 2310 1883 2316 1884
rect 2470 1888 2476 1889
rect 2470 1884 2471 1888
rect 2475 1884 2476 1888
rect 2470 1883 2476 1884
rect 2638 1888 2644 1889
rect 2638 1884 2639 1888
rect 2643 1884 2644 1888
rect 2638 1883 2644 1884
rect 2814 1888 2820 1889
rect 2814 1884 2815 1888
rect 2819 1884 2820 1888
rect 2814 1883 2820 1884
rect 2998 1888 3004 1889
rect 2998 1884 2999 1888
rect 3003 1884 3004 1888
rect 2998 1883 3004 1884
rect 3158 1888 3164 1889
rect 3158 1884 3159 1888
rect 3163 1884 3164 1888
rect 3158 1883 3164 1884
rect 110 1879 116 1880
rect 110 1875 111 1879
rect 115 1875 116 1879
rect 886 1879 893 1880
rect 110 1874 116 1875
rect 630 1875 636 1876
rect 630 1871 631 1875
rect 635 1871 636 1875
rect 630 1870 636 1871
rect 638 1875 645 1876
rect 638 1871 639 1875
rect 644 1871 645 1875
rect 638 1870 645 1871
rect 758 1875 764 1876
rect 758 1871 759 1875
rect 763 1871 764 1875
rect 758 1870 764 1871
rect 766 1875 773 1876
rect 766 1871 767 1875
rect 772 1871 773 1875
rect 766 1870 773 1871
rect 878 1875 884 1876
rect 878 1871 879 1875
rect 883 1871 884 1875
rect 886 1875 887 1879
rect 892 1875 893 1879
rect 1006 1879 1013 1880
rect 886 1874 893 1875
rect 998 1875 1004 1876
rect 878 1870 884 1871
rect 998 1871 999 1875
rect 1003 1871 1004 1875
rect 1006 1875 1007 1879
rect 1012 1875 1013 1879
rect 1126 1879 1133 1880
rect 1006 1874 1013 1875
rect 1118 1875 1124 1876
rect 998 1870 1004 1871
rect 1118 1871 1119 1875
rect 1123 1871 1124 1875
rect 1126 1875 1127 1879
rect 1132 1875 1133 1879
rect 1239 1879 1248 1880
rect 1126 1874 1133 1875
rect 1230 1875 1236 1876
rect 1118 1870 1124 1871
rect 1230 1871 1231 1875
rect 1235 1871 1236 1875
rect 1239 1875 1240 1879
rect 1247 1878 1248 1879
rect 1254 1879 1260 1880
rect 1254 1878 1255 1879
rect 1247 1876 1255 1878
rect 1247 1875 1248 1876
rect 1239 1874 1248 1875
rect 1254 1875 1255 1876
rect 1259 1875 1260 1879
rect 1351 1879 1360 1880
rect 1254 1874 1260 1875
rect 1342 1875 1348 1876
rect 1230 1870 1236 1871
rect 1342 1871 1343 1875
rect 1347 1871 1348 1875
rect 1351 1875 1352 1879
rect 1359 1875 1360 1879
rect 1470 1879 1477 1880
rect 1351 1874 1360 1875
rect 1462 1875 1468 1876
rect 1342 1870 1348 1871
rect 1462 1871 1463 1875
rect 1467 1871 1468 1875
rect 1470 1875 1471 1879
rect 1476 1875 1477 1879
rect 1470 1874 1477 1875
rect 1630 1879 1636 1880
rect 1630 1875 1631 1879
rect 1635 1875 1636 1879
rect 1630 1874 1636 1875
rect 1462 1870 1468 1871
rect 2070 1872 2076 1873
rect 2070 1868 2071 1872
rect 2075 1868 2076 1872
rect 2070 1867 2076 1868
rect 2238 1872 2244 1873
rect 2238 1868 2239 1872
rect 2243 1868 2244 1872
rect 2238 1867 2244 1868
rect 2414 1872 2420 1873
rect 2414 1868 2415 1872
rect 2419 1868 2420 1872
rect 2414 1867 2420 1868
rect 2598 1872 2604 1873
rect 2598 1868 2599 1872
rect 2603 1868 2604 1872
rect 2598 1867 2604 1868
rect 2790 1872 2796 1873
rect 2790 1868 2791 1872
rect 2795 1868 2796 1872
rect 2790 1867 2796 1868
rect 2982 1872 2988 1873
rect 2982 1868 2983 1872
rect 2987 1868 2988 1872
rect 2982 1867 2988 1868
rect 3158 1872 3164 1873
rect 3158 1868 3159 1872
rect 3163 1868 3164 1872
rect 3158 1867 3164 1868
rect 1670 1865 1676 1866
rect 1670 1861 1671 1865
rect 1675 1861 1676 1865
rect 1670 1860 1676 1861
rect 3190 1865 3196 1866
rect 3190 1861 3191 1865
rect 3195 1861 3196 1865
rect 3190 1860 3196 1861
rect 526 1853 532 1854
rect 110 1849 116 1850
rect 110 1845 111 1849
rect 115 1845 116 1849
rect 526 1849 527 1853
rect 531 1849 532 1853
rect 654 1853 660 1854
rect 526 1848 532 1849
rect 535 1851 541 1852
rect 535 1847 536 1851
rect 540 1850 541 1851
rect 638 1851 644 1852
rect 638 1850 639 1851
rect 540 1848 639 1850
rect 540 1847 541 1848
rect 535 1846 541 1847
rect 638 1847 639 1848
rect 643 1847 644 1851
rect 654 1849 655 1853
rect 659 1849 660 1853
rect 654 1848 660 1849
rect 774 1853 780 1854
rect 774 1849 775 1853
rect 779 1849 780 1853
rect 774 1848 780 1849
rect 894 1853 900 1854
rect 894 1849 895 1853
rect 899 1849 900 1853
rect 894 1848 900 1849
rect 1014 1853 1020 1854
rect 1014 1849 1015 1853
rect 1019 1849 1020 1853
rect 1014 1848 1020 1849
rect 1126 1853 1132 1854
rect 1126 1849 1127 1853
rect 1131 1849 1132 1853
rect 1246 1853 1252 1854
rect 1126 1848 1132 1849
rect 1134 1851 1141 1852
rect 638 1846 644 1847
rect 663 1847 669 1848
rect 663 1846 664 1847
rect 110 1844 116 1845
rect 640 1844 664 1846
rect 663 1843 664 1844
rect 668 1846 669 1847
rect 686 1847 692 1848
rect 686 1846 687 1847
rect 668 1844 687 1846
rect 668 1843 669 1844
rect 663 1842 669 1843
rect 686 1843 687 1844
rect 691 1846 692 1847
rect 766 1847 772 1848
rect 766 1846 767 1847
rect 691 1844 767 1846
rect 691 1843 692 1844
rect 686 1842 692 1843
rect 766 1843 767 1844
rect 771 1846 772 1847
rect 783 1847 789 1848
rect 783 1846 784 1847
rect 771 1844 784 1846
rect 771 1843 772 1844
rect 766 1842 772 1843
rect 783 1843 784 1844
rect 788 1846 789 1847
rect 806 1847 812 1848
rect 806 1846 807 1847
rect 788 1844 807 1846
rect 788 1843 789 1844
rect 783 1842 789 1843
rect 806 1843 807 1844
rect 811 1843 812 1847
rect 806 1842 812 1843
rect 886 1847 892 1848
rect 886 1843 887 1847
rect 891 1846 892 1847
rect 903 1847 909 1848
rect 903 1846 904 1847
rect 891 1844 904 1846
rect 891 1843 892 1844
rect 886 1842 892 1843
rect 903 1843 904 1844
rect 908 1846 909 1847
rect 926 1847 932 1848
rect 926 1846 927 1847
rect 908 1844 927 1846
rect 908 1843 909 1844
rect 903 1842 909 1843
rect 926 1843 927 1844
rect 931 1843 932 1847
rect 926 1842 932 1843
rect 1006 1847 1012 1848
rect 1006 1843 1007 1847
rect 1011 1846 1012 1847
rect 1023 1847 1029 1848
rect 1023 1846 1024 1847
rect 1011 1844 1024 1846
rect 1011 1843 1012 1844
rect 1006 1842 1012 1843
rect 1023 1843 1024 1844
rect 1028 1846 1029 1847
rect 1038 1847 1044 1848
rect 1038 1846 1039 1847
rect 1028 1844 1039 1846
rect 1028 1843 1029 1844
rect 1023 1842 1029 1843
rect 1038 1843 1039 1844
rect 1043 1843 1044 1847
rect 1134 1847 1135 1851
rect 1140 1847 1141 1851
rect 1246 1849 1247 1853
rect 1251 1849 1252 1853
rect 1366 1853 1372 1854
rect 1246 1848 1252 1849
rect 1254 1851 1261 1852
rect 1134 1846 1141 1847
rect 1254 1847 1255 1851
rect 1260 1847 1261 1851
rect 1366 1849 1367 1853
rect 1371 1849 1372 1853
rect 2158 1851 2164 1852
rect 1366 1848 1372 1849
rect 1630 1849 1636 1850
rect 1254 1846 1261 1847
rect 1354 1847 1360 1848
rect 1038 1842 1044 1843
rect 1354 1843 1355 1847
rect 1359 1846 1360 1847
rect 1375 1847 1381 1848
rect 1375 1846 1376 1847
rect 1359 1844 1376 1846
rect 1359 1843 1360 1844
rect 1354 1842 1360 1843
rect 1375 1843 1376 1844
rect 1380 1843 1381 1847
rect 1630 1845 1631 1849
rect 1635 1845 1636 1849
rect 1630 1844 1636 1845
rect 1670 1847 1676 1848
rect 1375 1842 1381 1843
rect 1670 1843 1671 1847
rect 1675 1843 1676 1847
rect 2158 1847 2159 1851
rect 2163 1850 2164 1851
rect 2246 1851 2252 1852
rect 2246 1850 2247 1851
rect 2163 1848 2247 1850
rect 2163 1847 2164 1848
rect 2158 1846 2164 1847
rect 2246 1847 2247 1848
rect 2251 1848 2252 1851
rect 2550 1851 2556 1852
rect 2251 1847 2253 1848
rect 2246 1846 2248 1847
rect 1670 1842 1676 1843
rect 2070 1843 2076 1844
rect 2070 1839 2071 1843
rect 2075 1839 2076 1843
rect 2070 1838 2076 1839
rect 2078 1843 2085 1844
rect 2078 1839 2079 1843
rect 2084 1839 2085 1843
rect 2078 1838 2085 1839
rect 2238 1843 2244 1844
rect 2238 1839 2239 1843
rect 2243 1839 2244 1843
rect 2247 1843 2248 1846
rect 2252 1843 2253 1847
rect 2422 1847 2429 1848
rect 2247 1842 2253 1843
rect 2414 1843 2420 1844
rect 2238 1838 2244 1839
rect 2414 1839 2415 1843
rect 2419 1839 2420 1843
rect 2422 1843 2423 1847
rect 2428 1843 2429 1847
rect 2550 1847 2551 1851
rect 2555 1850 2556 1851
rect 2590 1851 2596 1852
rect 2590 1850 2591 1851
rect 2555 1848 2591 1850
rect 2555 1847 2556 1848
rect 2550 1846 2556 1847
rect 2590 1847 2591 1848
rect 2595 1850 2596 1851
rect 2595 1848 2611 1850
rect 2595 1847 2596 1848
rect 2590 1846 2596 1847
rect 2607 1847 2613 1848
rect 2422 1842 2429 1843
rect 2598 1843 2604 1844
rect 2414 1838 2420 1839
rect 2598 1839 2599 1843
rect 2603 1839 2604 1843
rect 2607 1843 2608 1847
rect 2612 1843 2613 1847
rect 2799 1847 2805 1848
rect 2607 1842 2613 1843
rect 2790 1843 2796 1844
rect 2598 1838 2604 1839
rect 2790 1839 2791 1843
rect 2795 1839 2796 1843
rect 2799 1843 2800 1847
rect 2804 1846 2805 1847
rect 2822 1847 2828 1848
rect 2822 1846 2823 1847
rect 2804 1844 2823 1846
rect 2804 1843 2805 1844
rect 2799 1842 2805 1843
rect 2822 1843 2823 1844
rect 2827 1843 2828 1847
rect 2991 1847 2997 1848
rect 2822 1842 2828 1843
rect 2982 1843 2988 1844
rect 2790 1838 2796 1839
rect 1982 1833 1988 1834
rect 110 1831 116 1832
rect 110 1827 111 1831
rect 115 1827 116 1831
rect 110 1826 116 1827
rect 1630 1831 1636 1832
rect 1630 1827 1631 1831
rect 1635 1827 1636 1831
rect 1630 1826 1636 1827
rect 1670 1829 1676 1830
rect 1670 1825 1671 1829
rect 1675 1825 1676 1829
rect 1982 1829 1983 1833
rect 1987 1829 1988 1833
rect 1982 1828 1988 1829
rect 2134 1833 2140 1834
rect 2134 1829 2135 1833
rect 2139 1829 2140 1833
rect 2134 1828 2140 1829
rect 2286 1833 2292 1834
rect 2286 1829 2287 1833
rect 2291 1829 2292 1833
rect 2286 1828 2292 1829
rect 2430 1833 2436 1834
rect 2430 1829 2431 1833
rect 2435 1829 2436 1833
rect 2430 1828 2436 1829
rect 2582 1833 2588 1834
rect 2582 1829 2583 1833
rect 2587 1829 2588 1833
rect 2734 1833 2740 1834
rect 2582 1828 2588 1829
rect 2590 1831 2597 1832
rect 526 1824 532 1825
rect 526 1820 527 1824
rect 531 1820 532 1824
rect 526 1819 532 1820
rect 654 1824 660 1825
rect 654 1820 655 1824
rect 659 1820 660 1824
rect 654 1819 660 1820
rect 774 1824 780 1825
rect 774 1820 775 1824
rect 779 1820 780 1824
rect 774 1819 780 1820
rect 894 1824 900 1825
rect 894 1820 895 1824
rect 899 1820 900 1824
rect 894 1819 900 1820
rect 1014 1824 1020 1825
rect 1014 1820 1015 1824
rect 1019 1820 1020 1824
rect 1014 1819 1020 1820
rect 1126 1824 1132 1825
rect 1126 1820 1127 1824
rect 1131 1820 1132 1824
rect 1126 1819 1132 1820
rect 1246 1824 1252 1825
rect 1246 1820 1247 1824
rect 1251 1820 1252 1824
rect 1246 1819 1252 1820
rect 1366 1824 1372 1825
rect 1670 1824 1676 1825
rect 1990 1827 1997 1828
rect 1366 1820 1367 1824
rect 1371 1820 1372 1824
rect 1990 1823 1991 1827
rect 1996 1823 1997 1827
rect 1990 1822 1997 1823
rect 2086 1827 2092 1828
rect 2086 1823 2087 1827
rect 2091 1826 2092 1827
rect 2143 1827 2149 1828
rect 2143 1826 2144 1827
rect 2091 1824 2144 1826
rect 2091 1823 2092 1824
rect 2086 1822 2092 1823
rect 2143 1823 2144 1824
rect 2148 1826 2149 1827
rect 2158 1827 2164 1828
rect 2158 1826 2159 1827
rect 2148 1824 2159 1826
rect 2148 1823 2149 1824
rect 2143 1822 2149 1823
rect 2158 1823 2159 1824
rect 2163 1823 2164 1827
rect 2158 1822 2164 1823
rect 2246 1827 2252 1828
rect 2246 1823 2247 1827
rect 2251 1826 2252 1827
rect 2295 1827 2301 1828
rect 2295 1826 2296 1827
rect 2251 1824 2296 1826
rect 2251 1823 2252 1824
rect 2246 1822 2252 1823
rect 2295 1823 2296 1824
rect 2300 1823 2301 1827
rect 2295 1822 2301 1823
rect 2422 1827 2428 1828
rect 2422 1823 2423 1827
rect 2427 1826 2428 1827
rect 2439 1827 2445 1828
rect 2439 1826 2440 1827
rect 2427 1824 2440 1826
rect 2427 1823 2428 1824
rect 2422 1822 2428 1823
rect 2439 1823 2440 1824
rect 2444 1826 2445 1827
rect 2494 1827 2500 1828
rect 2494 1826 2495 1827
rect 2444 1824 2495 1826
rect 2444 1823 2445 1824
rect 2439 1822 2445 1823
rect 2494 1823 2495 1824
rect 2499 1823 2500 1827
rect 2590 1827 2591 1831
rect 2596 1827 2597 1831
rect 2734 1829 2735 1833
rect 2739 1829 2740 1833
rect 2734 1828 2740 1829
rect 2742 1831 2749 1832
rect 2590 1826 2597 1827
rect 2742 1827 2743 1831
rect 2748 1830 2749 1831
rect 2801 1830 2803 1842
rect 2982 1839 2983 1843
rect 2987 1839 2988 1843
rect 2991 1843 2992 1847
rect 2996 1846 2997 1847
rect 3006 1847 3012 1848
rect 3006 1846 3007 1847
rect 2996 1844 3007 1846
rect 2996 1843 2997 1844
rect 2991 1842 2997 1843
rect 3006 1843 3007 1844
rect 3011 1843 3012 1847
rect 3166 1847 3173 1848
rect 3006 1842 3012 1843
rect 3158 1843 3164 1844
rect 2982 1838 2988 1839
rect 3158 1839 3159 1843
rect 3163 1839 3164 1843
rect 3166 1843 3167 1847
rect 3172 1843 3173 1847
rect 3166 1842 3173 1843
rect 3190 1847 3196 1848
rect 3190 1843 3191 1847
rect 3195 1843 3196 1847
rect 3190 1842 3196 1843
rect 3158 1838 3164 1839
rect 2748 1828 2803 1830
rect 3190 1829 3196 1830
rect 2748 1827 2749 1828
rect 2742 1826 2749 1827
rect 3190 1825 3191 1829
rect 3195 1825 3196 1829
rect 3190 1824 3196 1825
rect 2494 1822 2500 1823
rect 1366 1819 1372 1820
rect 1670 1811 1676 1812
rect 1670 1807 1671 1811
rect 1675 1807 1676 1811
rect 1670 1806 1676 1807
rect 3190 1811 3196 1812
rect 3190 1807 3191 1811
rect 3195 1807 3196 1811
rect 3190 1806 3196 1807
rect 422 1804 428 1805
rect 422 1800 423 1804
rect 427 1800 428 1804
rect 422 1799 428 1800
rect 550 1804 556 1805
rect 550 1800 551 1804
rect 555 1800 556 1804
rect 550 1799 556 1800
rect 678 1804 684 1805
rect 678 1800 679 1804
rect 683 1800 684 1804
rect 678 1799 684 1800
rect 798 1804 804 1805
rect 798 1800 799 1804
rect 803 1800 804 1804
rect 798 1799 804 1800
rect 918 1804 924 1805
rect 918 1800 919 1804
rect 923 1800 924 1804
rect 918 1799 924 1800
rect 1030 1804 1036 1805
rect 1030 1800 1031 1804
rect 1035 1800 1036 1804
rect 1030 1799 1036 1800
rect 1142 1804 1148 1805
rect 1142 1800 1143 1804
rect 1147 1800 1148 1804
rect 1142 1799 1148 1800
rect 1262 1804 1268 1805
rect 1262 1800 1263 1804
rect 1267 1800 1268 1804
rect 1262 1799 1268 1800
rect 1982 1804 1988 1805
rect 1982 1800 1983 1804
rect 1987 1800 1988 1804
rect 1982 1799 1988 1800
rect 2134 1804 2140 1805
rect 2134 1800 2135 1804
rect 2139 1800 2140 1804
rect 2134 1799 2140 1800
rect 2286 1804 2292 1805
rect 2286 1800 2287 1804
rect 2291 1800 2292 1804
rect 2286 1799 2292 1800
rect 2430 1804 2436 1805
rect 2430 1800 2431 1804
rect 2435 1800 2436 1804
rect 2430 1799 2436 1800
rect 2582 1804 2588 1805
rect 2582 1800 2583 1804
rect 2587 1800 2588 1804
rect 2582 1799 2588 1800
rect 2734 1804 2740 1805
rect 2734 1800 2735 1804
rect 2739 1800 2740 1804
rect 2734 1799 2740 1800
rect 110 1797 116 1798
rect 110 1793 111 1797
rect 115 1793 116 1797
rect 110 1792 116 1793
rect 1630 1797 1636 1798
rect 1630 1793 1631 1797
rect 1635 1793 1636 1797
rect 1630 1792 1636 1793
rect 1902 1792 1908 1793
rect 1902 1788 1903 1792
rect 1907 1788 1908 1792
rect 1902 1787 1908 1788
rect 2078 1792 2084 1793
rect 2078 1788 2079 1792
rect 2083 1788 2084 1792
rect 2078 1787 2084 1788
rect 2270 1792 2276 1793
rect 2270 1788 2271 1792
rect 2275 1788 2276 1792
rect 2270 1787 2276 1788
rect 2486 1792 2492 1793
rect 2486 1788 2487 1792
rect 2491 1788 2492 1792
rect 2486 1787 2492 1788
rect 2710 1792 2716 1793
rect 2710 1788 2711 1792
rect 2715 1788 2716 1792
rect 2710 1787 2716 1788
rect 2942 1792 2948 1793
rect 2942 1788 2943 1792
rect 2947 1788 2948 1792
rect 2942 1787 2948 1788
rect 3158 1792 3164 1793
rect 3158 1788 3159 1792
rect 3163 1788 3164 1792
rect 3158 1787 3164 1788
rect 1670 1785 1676 1786
rect 1134 1783 1140 1784
rect 110 1779 116 1780
rect 110 1775 111 1779
rect 115 1775 116 1779
rect 686 1779 693 1780
rect 110 1774 116 1775
rect 422 1775 428 1776
rect 422 1771 423 1775
rect 427 1771 428 1775
rect 422 1770 428 1771
rect 430 1775 437 1776
rect 430 1771 431 1775
rect 436 1771 437 1775
rect 430 1770 437 1771
rect 550 1775 556 1776
rect 550 1771 551 1775
rect 555 1771 556 1775
rect 550 1770 556 1771
rect 558 1775 565 1776
rect 558 1771 559 1775
rect 564 1771 565 1775
rect 558 1770 565 1771
rect 678 1775 684 1776
rect 678 1771 679 1775
rect 683 1771 684 1775
rect 686 1775 687 1779
rect 692 1775 693 1779
rect 806 1779 813 1780
rect 686 1774 693 1775
rect 798 1775 804 1776
rect 678 1770 684 1771
rect 798 1771 799 1775
rect 803 1771 804 1775
rect 806 1775 807 1779
rect 812 1775 813 1779
rect 926 1779 933 1780
rect 806 1774 813 1775
rect 918 1775 924 1776
rect 798 1770 804 1771
rect 918 1771 919 1775
rect 923 1771 924 1775
rect 926 1775 927 1779
rect 932 1775 933 1779
rect 1038 1779 1045 1780
rect 926 1774 933 1775
rect 1030 1775 1036 1776
rect 918 1770 924 1771
rect 1030 1771 1031 1775
rect 1035 1771 1036 1775
rect 1038 1775 1039 1779
rect 1044 1775 1045 1779
rect 1134 1779 1135 1783
rect 1139 1782 1140 1783
rect 1254 1783 1260 1784
rect 1139 1780 1154 1782
rect 1139 1779 1140 1780
rect 1134 1778 1140 1779
rect 1151 1779 1157 1780
rect 1038 1774 1045 1775
rect 1142 1775 1148 1776
rect 1030 1770 1036 1771
rect 1142 1771 1143 1775
rect 1147 1771 1148 1775
rect 1151 1775 1152 1779
rect 1156 1775 1157 1779
rect 1254 1779 1255 1783
rect 1259 1782 1260 1783
rect 1259 1780 1274 1782
rect 1670 1781 1671 1785
rect 1675 1781 1676 1785
rect 1670 1780 1676 1781
rect 3190 1785 3196 1786
rect 3190 1781 3191 1785
rect 3195 1781 3196 1785
rect 3190 1780 3196 1781
rect 1259 1779 1260 1780
rect 1254 1778 1260 1779
rect 1271 1779 1277 1780
rect 1151 1774 1157 1775
rect 1262 1775 1268 1776
rect 1142 1770 1148 1771
rect 1262 1771 1263 1775
rect 1267 1771 1268 1775
rect 1271 1775 1272 1779
rect 1276 1775 1277 1779
rect 1271 1774 1277 1775
rect 1630 1779 1636 1780
rect 1630 1775 1631 1779
rect 1635 1775 1636 1779
rect 1630 1774 1636 1775
rect 1262 1770 1268 1771
rect 2086 1771 2092 1772
rect 2086 1770 2087 1771
rect 1992 1768 2087 1770
rect 1670 1767 1676 1768
rect 1670 1763 1671 1767
rect 1675 1763 1676 1767
rect 1911 1767 1917 1768
rect 1670 1762 1676 1763
rect 1902 1763 1908 1764
rect 1902 1759 1903 1763
rect 1907 1759 1908 1763
rect 1911 1763 1912 1767
rect 1916 1766 1917 1767
rect 1990 1767 1996 1768
rect 1990 1766 1991 1767
rect 1916 1764 1991 1766
rect 1916 1763 1917 1764
rect 1911 1762 1917 1763
rect 1990 1763 1991 1764
rect 1995 1763 1996 1767
rect 2086 1767 2087 1768
rect 2091 1768 2092 1771
rect 2246 1771 2252 1772
rect 2091 1767 2093 1768
rect 2086 1766 2088 1767
rect 1990 1762 1996 1763
rect 2078 1763 2084 1764
rect 1902 1758 1908 1759
rect 2078 1759 2079 1763
rect 2083 1759 2084 1763
rect 2087 1763 2088 1766
rect 2092 1763 2093 1767
rect 2246 1767 2247 1771
rect 2251 1770 2252 1771
rect 2251 1768 2283 1770
rect 2251 1767 2252 1768
rect 2246 1766 2252 1767
rect 2279 1767 2285 1768
rect 2087 1762 2093 1763
rect 2270 1763 2276 1764
rect 2078 1758 2084 1759
rect 2270 1759 2271 1763
rect 2275 1759 2276 1763
rect 2279 1763 2280 1767
rect 2284 1763 2285 1767
rect 2494 1767 2501 1768
rect 2279 1762 2285 1763
rect 2486 1763 2492 1764
rect 2270 1758 2276 1759
rect 2486 1759 2487 1763
rect 2491 1759 2492 1763
rect 2494 1763 2495 1767
rect 2500 1763 2501 1767
rect 2719 1767 2725 1768
rect 2494 1762 2501 1763
rect 2710 1763 2716 1764
rect 2486 1758 2492 1759
rect 2710 1759 2711 1763
rect 2715 1759 2716 1763
rect 2719 1763 2720 1767
rect 2724 1766 2725 1767
rect 2742 1767 2748 1768
rect 2742 1766 2743 1767
rect 2724 1764 2743 1766
rect 2724 1763 2725 1764
rect 2719 1762 2725 1763
rect 2742 1763 2743 1764
rect 2747 1763 2748 1767
rect 2950 1767 2957 1768
rect 2742 1762 2748 1763
rect 2942 1763 2948 1764
rect 2710 1758 2716 1759
rect 2942 1759 2943 1763
rect 2947 1759 2948 1763
rect 2950 1763 2951 1767
rect 2956 1766 2957 1767
rect 3006 1767 3012 1768
rect 3006 1766 3007 1767
rect 2956 1764 3007 1766
rect 2956 1763 2957 1764
rect 2950 1762 2957 1763
rect 3006 1763 3007 1764
rect 3011 1763 3012 1767
rect 3166 1767 3173 1768
rect 3006 1762 3012 1763
rect 3158 1763 3164 1764
rect 2942 1758 2948 1759
rect 3158 1759 3159 1763
rect 3163 1759 3164 1763
rect 3166 1763 3167 1767
rect 3172 1763 3173 1767
rect 3166 1762 3173 1763
rect 3190 1767 3196 1768
rect 3190 1763 3191 1767
rect 3195 1763 3196 1767
rect 3190 1762 3196 1763
rect 3158 1758 3164 1759
rect 326 1753 332 1754
rect 110 1749 116 1750
rect 110 1745 111 1749
rect 115 1745 116 1749
rect 326 1749 327 1753
rect 331 1749 332 1753
rect 326 1748 332 1749
rect 454 1753 460 1754
rect 454 1749 455 1753
rect 459 1749 460 1753
rect 454 1748 460 1749
rect 574 1753 580 1754
rect 574 1749 575 1753
rect 579 1749 580 1753
rect 574 1748 580 1749
rect 694 1753 700 1754
rect 694 1749 695 1753
rect 699 1749 700 1753
rect 694 1748 700 1749
rect 814 1753 820 1754
rect 814 1749 815 1753
rect 819 1749 820 1753
rect 926 1753 932 1754
rect 814 1748 820 1749
rect 823 1749 829 1750
rect 823 1748 824 1749
rect 110 1744 116 1745
rect 334 1747 341 1748
rect 334 1743 335 1747
rect 340 1746 341 1747
rect 430 1747 436 1748
rect 430 1746 431 1747
rect 340 1744 431 1746
rect 340 1743 341 1744
rect 334 1742 341 1743
rect 430 1743 431 1744
rect 435 1746 436 1747
rect 463 1747 469 1748
rect 463 1746 464 1747
rect 435 1744 464 1746
rect 435 1743 436 1744
rect 430 1742 436 1743
rect 463 1743 464 1744
rect 468 1746 469 1747
rect 558 1747 564 1748
rect 558 1746 559 1747
rect 468 1744 559 1746
rect 468 1743 469 1744
rect 463 1742 469 1743
rect 558 1743 559 1744
rect 563 1746 564 1747
rect 583 1747 589 1748
rect 583 1746 584 1747
rect 563 1744 584 1746
rect 563 1743 564 1744
rect 558 1742 564 1743
rect 583 1743 584 1744
rect 588 1746 589 1747
rect 703 1747 709 1748
rect 703 1746 704 1747
rect 588 1744 704 1746
rect 588 1743 589 1744
rect 583 1742 589 1743
rect 703 1743 704 1744
rect 708 1746 709 1747
rect 718 1747 724 1748
rect 718 1746 719 1747
rect 708 1744 719 1746
rect 708 1743 709 1744
rect 703 1742 709 1743
rect 718 1743 719 1744
rect 723 1746 724 1747
rect 822 1747 824 1748
rect 822 1746 823 1747
rect 723 1744 823 1746
rect 828 1745 829 1749
rect 926 1749 927 1753
rect 931 1749 932 1753
rect 926 1748 932 1749
rect 1038 1753 1044 1754
rect 1038 1749 1039 1753
rect 1043 1749 1044 1753
rect 1038 1748 1044 1749
rect 1158 1753 1164 1754
rect 1158 1749 1159 1753
rect 1163 1749 1164 1753
rect 1158 1748 1164 1749
rect 1630 1749 1636 1750
rect 723 1743 724 1744
rect 718 1742 724 1743
rect 822 1743 823 1744
rect 827 1744 829 1745
rect 935 1747 941 1748
rect 827 1743 828 1744
rect 822 1742 828 1743
rect 935 1743 936 1747
rect 940 1746 941 1747
rect 950 1747 956 1748
rect 950 1746 951 1747
rect 940 1744 951 1746
rect 940 1743 941 1744
rect 935 1742 941 1743
rect 950 1743 951 1744
rect 955 1746 956 1747
rect 1047 1747 1053 1748
rect 1047 1746 1048 1747
rect 955 1744 1048 1746
rect 955 1743 956 1744
rect 950 1742 956 1743
rect 1047 1743 1048 1744
rect 1052 1743 1053 1747
rect 1047 1742 1053 1743
rect 1166 1747 1173 1748
rect 1166 1743 1167 1747
rect 1172 1743 1173 1747
rect 1630 1745 1631 1749
rect 1635 1745 1636 1749
rect 1630 1744 1636 1745
rect 1814 1745 1820 1746
rect 1166 1742 1173 1743
rect 1670 1741 1676 1742
rect 1670 1737 1671 1741
rect 1675 1737 1676 1741
rect 1814 1741 1815 1745
rect 1819 1741 1820 1745
rect 1814 1740 1820 1741
rect 1966 1745 1972 1746
rect 1966 1741 1967 1745
rect 1971 1741 1972 1745
rect 1966 1740 1972 1741
rect 2126 1745 2132 1746
rect 2126 1741 2127 1745
rect 2131 1741 2132 1745
rect 2126 1740 2132 1741
rect 2302 1745 2308 1746
rect 2302 1741 2303 1745
rect 2307 1741 2308 1745
rect 2302 1740 2308 1741
rect 2502 1745 2508 1746
rect 2502 1741 2503 1745
rect 2507 1741 2508 1745
rect 2502 1740 2508 1741
rect 2710 1745 2716 1746
rect 2710 1741 2711 1745
rect 2715 1741 2716 1745
rect 2710 1740 2716 1741
rect 2934 1745 2940 1746
rect 2934 1741 2935 1745
rect 2939 1741 2940 1745
rect 2934 1740 2940 1741
rect 3158 1745 3164 1746
rect 3158 1741 3159 1745
rect 3163 1741 3164 1745
rect 3158 1740 3164 1741
rect 3166 1743 3173 1744
rect 1670 1736 1676 1737
rect 1822 1739 1829 1740
rect 1822 1735 1823 1739
rect 1828 1738 1829 1739
rect 1975 1739 1981 1740
rect 1975 1738 1976 1739
rect 1828 1736 1976 1738
rect 1828 1735 1829 1736
rect 1822 1734 1829 1735
rect 1975 1735 1976 1736
rect 1980 1738 1981 1739
rect 2030 1739 2036 1740
rect 2030 1738 2031 1739
rect 1980 1736 2031 1738
rect 1980 1735 1981 1736
rect 1975 1734 1981 1735
rect 2030 1735 2031 1736
rect 2035 1738 2036 1739
rect 2135 1739 2141 1740
rect 2135 1738 2136 1739
rect 2035 1736 2136 1738
rect 2035 1735 2036 1736
rect 2030 1734 2036 1735
rect 2135 1735 2136 1736
rect 2140 1735 2141 1739
rect 2135 1734 2141 1735
rect 2311 1739 2317 1740
rect 2311 1735 2312 1739
rect 2316 1738 2317 1739
rect 2322 1739 2328 1740
rect 2322 1738 2323 1739
rect 2316 1736 2323 1738
rect 2316 1735 2317 1736
rect 2311 1734 2317 1735
rect 2322 1735 2323 1736
rect 2327 1735 2328 1739
rect 2322 1734 2328 1735
rect 2474 1739 2480 1740
rect 2474 1735 2475 1739
rect 2479 1738 2480 1739
rect 2511 1739 2517 1740
rect 2511 1738 2512 1739
rect 2479 1736 2512 1738
rect 2479 1735 2480 1736
rect 2474 1734 2480 1735
rect 2511 1735 2512 1736
rect 2516 1738 2517 1739
rect 2718 1739 2725 1740
rect 2718 1738 2719 1739
rect 2516 1736 2719 1738
rect 2516 1735 2517 1736
rect 2511 1734 2517 1735
rect 2718 1735 2719 1736
rect 2724 1735 2725 1739
rect 2718 1734 2725 1735
rect 2943 1739 2949 1740
rect 2943 1735 2944 1739
rect 2948 1735 2949 1739
rect 3166 1739 3167 1743
rect 3172 1739 3173 1743
rect 3166 1738 3173 1739
rect 3190 1741 3196 1742
rect 3190 1737 3191 1741
rect 3195 1737 3196 1741
rect 3190 1736 3196 1737
rect 2943 1734 2949 1735
rect 110 1731 116 1732
rect 110 1727 111 1731
rect 115 1727 116 1731
rect 110 1726 116 1727
rect 1630 1731 1636 1732
rect 1630 1727 1631 1731
rect 1635 1727 1636 1731
rect 1630 1726 1636 1727
rect 326 1724 332 1725
rect 326 1720 327 1724
rect 331 1720 332 1724
rect 326 1719 332 1720
rect 454 1724 460 1725
rect 454 1720 455 1724
rect 459 1720 460 1724
rect 454 1719 460 1720
rect 574 1724 580 1725
rect 574 1720 575 1724
rect 579 1720 580 1724
rect 574 1719 580 1720
rect 694 1724 700 1725
rect 694 1720 695 1724
rect 699 1720 700 1724
rect 694 1719 700 1720
rect 814 1724 820 1725
rect 814 1720 815 1724
rect 819 1720 820 1724
rect 814 1719 820 1720
rect 926 1724 932 1725
rect 926 1720 927 1724
rect 931 1720 932 1724
rect 926 1719 932 1720
rect 1038 1724 1044 1725
rect 1038 1720 1039 1724
rect 1043 1720 1044 1724
rect 1038 1719 1044 1720
rect 1158 1724 1164 1725
rect 1158 1720 1159 1724
rect 1163 1720 1164 1724
rect 1158 1719 1164 1720
rect 1670 1723 1676 1724
rect 1670 1719 1671 1723
rect 1675 1719 1676 1723
rect 1670 1718 1676 1719
rect 3190 1723 3196 1724
rect 3190 1719 3191 1723
rect 3195 1719 3196 1723
rect 3190 1718 3196 1719
rect 1814 1716 1820 1717
rect 1814 1712 1815 1716
rect 1819 1712 1820 1716
rect 1814 1711 1820 1712
rect 1966 1716 1972 1717
rect 1966 1712 1967 1716
rect 1971 1712 1972 1716
rect 1966 1711 1972 1712
rect 2126 1716 2132 1717
rect 2126 1712 2127 1716
rect 2131 1712 2132 1716
rect 2126 1711 2132 1712
rect 2302 1716 2308 1717
rect 2302 1712 2303 1716
rect 2307 1712 2308 1716
rect 2302 1711 2308 1712
rect 2502 1716 2508 1717
rect 2502 1712 2503 1716
rect 2507 1712 2508 1716
rect 2502 1711 2508 1712
rect 2710 1716 2716 1717
rect 2710 1712 2711 1716
rect 2715 1712 2716 1716
rect 2710 1711 2716 1712
rect 2934 1716 2940 1717
rect 2934 1712 2935 1716
rect 2939 1712 2940 1716
rect 2934 1711 2940 1712
rect 3158 1716 3164 1717
rect 3158 1712 3159 1716
rect 3163 1712 3164 1716
rect 3158 1711 3164 1712
rect 1734 1704 1740 1705
rect 222 1700 228 1701
rect 222 1696 223 1700
rect 227 1696 228 1700
rect 222 1695 228 1696
rect 350 1700 356 1701
rect 350 1696 351 1700
rect 355 1696 356 1700
rect 350 1695 356 1696
rect 470 1700 476 1701
rect 470 1696 471 1700
rect 475 1696 476 1700
rect 470 1695 476 1696
rect 590 1700 596 1701
rect 590 1696 591 1700
rect 595 1696 596 1700
rect 590 1695 596 1696
rect 710 1700 716 1701
rect 710 1696 711 1700
rect 715 1696 716 1700
rect 710 1695 716 1696
rect 822 1700 828 1701
rect 822 1696 823 1700
rect 827 1696 828 1700
rect 822 1695 828 1696
rect 942 1700 948 1701
rect 942 1696 943 1700
rect 947 1696 948 1700
rect 942 1695 948 1696
rect 1062 1700 1068 1701
rect 1062 1696 1063 1700
rect 1067 1696 1068 1700
rect 1734 1700 1735 1704
rect 1739 1700 1740 1704
rect 1734 1699 1740 1700
rect 1878 1704 1884 1705
rect 1878 1700 1879 1704
rect 1883 1700 1884 1704
rect 1878 1699 1884 1700
rect 2022 1704 2028 1705
rect 2022 1700 2023 1704
rect 2027 1700 2028 1704
rect 2022 1699 2028 1700
rect 2166 1704 2172 1705
rect 2166 1700 2167 1704
rect 2171 1700 2172 1704
rect 2166 1699 2172 1700
rect 2310 1704 2316 1705
rect 2310 1700 2311 1704
rect 2315 1700 2316 1704
rect 2310 1699 2316 1700
rect 2462 1704 2468 1705
rect 2462 1700 2463 1704
rect 2467 1700 2468 1704
rect 2462 1699 2468 1700
rect 1062 1695 1068 1696
rect 1670 1697 1676 1698
rect 110 1693 116 1694
rect 110 1689 111 1693
rect 115 1689 116 1693
rect 110 1688 116 1689
rect 1630 1693 1636 1694
rect 1630 1689 1631 1693
rect 1635 1689 1636 1693
rect 1670 1693 1671 1697
rect 1675 1693 1676 1697
rect 1670 1692 1676 1693
rect 3190 1697 3196 1698
rect 3190 1693 3191 1697
rect 3195 1693 3196 1697
rect 3190 1692 3196 1693
rect 1630 1688 1636 1689
rect 1822 1683 1828 1684
rect 926 1679 932 1680
rect 926 1678 927 1679
rect 919 1676 927 1678
rect 110 1675 116 1676
rect 110 1671 111 1675
rect 115 1671 116 1675
rect 718 1675 725 1676
rect 110 1670 116 1671
rect 222 1671 228 1672
rect 222 1667 223 1671
rect 227 1667 228 1671
rect 222 1666 228 1667
rect 230 1671 237 1672
rect 230 1667 231 1671
rect 236 1667 237 1671
rect 230 1666 237 1667
rect 350 1671 356 1672
rect 350 1667 351 1671
rect 355 1667 356 1671
rect 350 1666 356 1667
rect 359 1671 365 1672
rect 359 1667 360 1671
rect 364 1667 365 1671
rect 359 1666 365 1667
rect 470 1671 476 1672
rect 470 1667 471 1671
rect 475 1667 476 1671
rect 470 1666 476 1667
rect 478 1671 485 1672
rect 478 1667 479 1671
rect 484 1667 485 1671
rect 478 1666 485 1667
rect 590 1671 596 1672
rect 590 1667 591 1671
rect 595 1667 596 1671
rect 590 1666 596 1667
rect 598 1671 605 1672
rect 598 1667 599 1671
rect 604 1667 605 1671
rect 598 1666 605 1667
rect 710 1671 716 1672
rect 710 1667 711 1671
rect 715 1667 716 1671
rect 718 1671 719 1675
rect 724 1671 725 1675
rect 830 1675 837 1676
rect 718 1670 725 1671
rect 822 1671 828 1672
rect 710 1666 716 1667
rect 822 1667 823 1671
rect 827 1667 828 1671
rect 830 1671 831 1675
rect 836 1674 837 1675
rect 919 1674 921 1676
rect 926 1675 927 1676
rect 931 1678 932 1679
rect 1670 1679 1676 1680
rect 931 1676 954 1678
rect 931 1675 932 1676
rect 926 1674 932 1675
rect 950 1675 957 1676
rect 836 1672 921 1674
rect 836 1671 837 1672
rect 830 1670 837 1671
rect 942 1671 948 1672
rect 822 1666 828 1667
rect 942 1667 943 1671
rect 947 1667 948 1671
rect 950 1671 951 1675
rect 956 1671 957 1675
rect 1630 1675 1636 1676
rect 950 1670 957 1671
rect 1062 1671 1068 1672
rect 942 1666 948 1667
rect 1062 1667 1063 1671
rect 1067 1667 1068 1671
rect 1062 1666 1068 1667
rect 1070 1671 1077 1672
rect 1070 1667 1071 1671
rect 1076 1667 1077 1671
rect 1630 1671 1631 1675
rect 1635 1671 1636 1675
rect 1670 1675 1671 1679
rect 1675 1675 1676 1679
rect 1822 1679 1823 1683
rect 1827 1682 1828 1683
rect 1827 1680 1890 1682
rect 1827 1679 1828 1680
rect 1822 1678 1828 1679
rect 1887 1679 1893 1680
rect 1670 1674 1676 1675
rect 1734 1675 1740 1676
rect 1630 1670 1636 1671
rect 1734 1671 1735 1675
rect 1739 1671 1740 1675
rect 1734 1670 1740 1671
rect 1743 1675 1749 1676
rect 1743 1671 1744 1675
rect 1748 1674 1749 1675
rect 1822 1675 1828 1676
rect 1822 1674 1823 1675
rect 1748 1672 1823 1674
rect 1748 1671 1749 1672
rect 1743 1670 1749 1671
rect 1822 1671 1823 1672
rect 1827 1671 1828 1675
rect 1822 1670 1828 1671
rect 1878 1675 1884 1676
rect 1878 1671 1879 1675
rect 1883 1671 1884 1675
rect 1887 1675 1888 1679
rect 1892 1678 1893 1679
rect 2030 1679 2037 1680
rect 1892 1676 1906 1678
rect 1892 1675 1893 1676
rect 1887 1674 1893 1675
rect 1878 1670 1884 1671
rect 1070 1666 1077 1667
rect 310 1663 316 1664
rect 310 1659 311 1663
rect 315 1662 316 1663
rect 334 1663 340 1664
rect 334 1662 335 1663
rect 315 1660 335 1662
rect 315 1659 316 1660
rect 310 1658 316 1659
rect 334 1659 335 1660
rect 339 1662 340 1663
rect 361 1662 363 1666
rect 1694 1665 1700 1666
rect 339 1660 363 1662
rect 339 1659 340 1660
rect 334 1658 340 1659
rect 361 1654 363 1660
rect 1670 1661 1676 1662
rect 1670 1657 1671 1661
rect 1675 1657 1676 1661
rect 1694 1661 1695 1665
rect 1699 1661 1700 1665
rect 1694 1660 1700 1661
rect 1703 1663 1709 1664
rect 1703 1659 1704 1663
rect 1708 1662 1709 1663
rect 1745 1662 1747 1670
rect 1708 1660 1747 1662
rect 1894 1665 1900 1666
rect 1894 1661 1895 1665
rect 1899 1661 1900 1665
rect 1904 1664 1906 1676
rect 2022 1675 2028 1676
rect 2022 1671 2023 1675
rect 2027 1671 2028 1675
rect 2030 1675 2031 1679
rect 2036 1678 2037 1679
rect 2106 1679 2112 1680
rect 2106 1678 2107 1679
rect 2036 1676 2107 1678
rect 2036 1675 2037 1676
rect 2030 1674 2037 1675
rect 2106 1675 2107 1676
rect 2111 1675 2112 1679
rect 2319 1679 2328 1680
rect 2106 1674 2112 1675
rect 2166 1675 2172 1676
rect 2022 1670 2028 1671
rect 2166 1671 2167 1675
rect 2171 1671 2172 1675
rect 2166 1670 2172 1671
rect 2175 1675 2181 1676
rect 2175 1671 2176 1675
rect 2180 1671 2181 1675
rect 2175 1670 2181 1671
rect 2310 1675 2316 1676
rect 2310 1671 2311 1675
rect 2315 1671 2316 1675
rect 2319 1675 2320 1679
rect 2327 1675 2328 1679
rect 2471 1679 2480 1680
rect 2319 1674 2328 1675
rect 2462 1675 2468 1676
rect 2310 1670 2316 1671
rect 2462 1671 2463 1675
rect 2467 1671 2468 1675
rect 2471 1675 2472 1679
rect 2479 1675 2480 1679
rect 2471 1674 2480 1675
rect 3190 1679 3196 1680
rect 3190 1675 3191 1679
rect 3195 1675 3196 1679
rect 3190 1674 3196 1675
rect 2462 1670 2468 1671
rect 2126 1665 2132 1666
rect 1894 1660 1900 1661
rect 1903 1663 1909 1664
rect 1708 1659 1709 1660
rect 1703 1658 1709 1659
rect 1903 1659 1904 1663
rect 1908 1659 1909 1663
rect 2126 1661 2127 1665
rect 2131 1661 2132 1665
rect 2126 1660 2132 1661
rect 1903 1658 1909 1659
rect 2106 1659 2112 1660
rect 1670 1656 1676 1657
rect 361 1652 395 1654
rect 134 1649 140 1650
rect 110 1645 116 1646
rect 110 1641 111 1645
rect 115 1641 116 1645
rect 134 1645 135 1649
rect 139 1645 140 1649
rect 134 1644 140 1645
rect 246 1649 252 1650
rect 246 1645 247 1649
rect 251 1645 252 1649
rect 246 1644 252 1645
rect 382 1649 388 1650
rect 382 1645 383 1649
rect 387 1645 388 1649
rect 393 1648 395 1652
rect 1705 1650 1707 1658
rect 2106 1655 2107 1659
rect 2111 1658 2112 1659
rect 2135 1659 2141 1660
rect 2135 1658 2136 1659
rect 2111 1656 2136 1658
rect 2111 1655 2112 1656
rect 2106 1654 2112 1655
rect 2135 1655 2136 1656
rect 2140 1658 2141 1659
rect 2177 1658 2179 1670
rect 2366 1665 2372 1666
rect 2366 1661 2367 1665
rect 2371 1661 2372 1665
rect 2366 1660 2372 1661
rect 2614 1665 2620 1666
rect 2614 1661 2615 1665
rect 2619 1661 2620 1665
rect 2614 1660 2620 1661
rect 2870 1665 2876 1666
rect 2870 1661 2871 1665
rect 2875 1661 2876 1665
rect 2870 1660 2876 1661
rect 3134 1665 3140 1666
rect 3134 1661 3135 1665
rect 3139 1661 3140 1665
rect 3134 1660 3140 1661
rect 3142 1663 3149 1664
rect 2140 1656 2179 1658
rect 2322 1659 2328 1660
rect 2140 1655 2141 1656
rect 2135 1654 2141 1655
rect 2322 1655 2323 1659
rect 2327 1658 2328 1659
rect 2375 1659 2381 1660
rect 2375 1658 2376 1659
rect 2327 1656 2376 1658
rect 2327 1655 2328 1656
rect 2322 1654 2328 1655
rect 2375 1655 2376 1656
rect 2380 1658 2381 1659
rect 2398 1659 2404 1660
rect 2398 1658 2399 1659
rect 2380 1656 2399 1658
rect 2380 1655 2381 1656
rect 2375 1654 2381 1655
rect 2398 1655 2399 1656
rect 2403 1655 2404 1659
rect 2398 1654 2404 1655
rect 2623 1659 2629 1660
rect 2623 1655 2624 1659
rect 2628 1658 2629 1659
rect 2718 1659 2724 1660
rect 2718 1658 2719 1659
rect 2628 1656 2719 1658
rect 2628 1655 2629 1656
rect 2623 1654 2629 1655
rect 2718 1655 2719 1656
rect 2723 1655 2724 1659
rect 2718 1654 2724 1655
rect 2879 1659 2885 1660
rect 2879 1655 2880 1659
rect 2884 1658 2885 1659
rect 2918 1659 2924 1660
rect 2918 1658 2919 1659
rect 2884 1656 2919 1658
rect 2884 1655 2885 1656
rect 2879 1654 2885 1655
rect 2918 1655 2919 1656
rect 2923 1655 2924 1659
rect 3142 1659 3143 1663
rect 3148 1662 3149 1663
rect 3166 1663 3172 1664
rect 3166 1662 3167 1663
rect 3148 1660 3167 1662
rect 3148 1659 3149 1660
rect 3142 1658 3149 1659
rect 3166 1659 3167 1660
rect 3171 1659 3172 1663
rect 3166 1658 3172 1659
rect 3190 1661 3196 1662
rect 3190 1657 3191 1661
rect 3195 1657 3196 1661
rect 3190 1656 3196 1657
rect 2918 1654 2924 1655
rect 534 1649 540 1650
rect 382 1644 388 1645
rect 391 1647 397 1648
rect 110 1640 116 1641
rect 142 1643 149 1644
rect 142 1639 143 1643
rect 148 1642 149 1643
rect 230 1643 236 1644
rect 230 1642 231 1643
rect 148 1640 231 1642
rect 148 1639 149 1640
rect 142 1638 149 1639
rect 230 1639 231 1640
rect 235 1642 236 1643
rect 255 1643 261 1644
rect 255 1642 256 1643
rect 235 1640 256 1642
rect 235 1639 236 1640
rect 230 1638 236 1639
rect 255 1639 256 1640
rect 260 1642 261 1643
rect 310 1643 316 1644
rect 310 1642 311 1643
rect 260 1640 311 1642
rect 260 1639 261 1640
rect 255 1638 261 1639
rect 310 1639 311 1640
rect 315 1639 316 1643
rect 391 1643 392 1647
rect 396 1646 397 1647
rect 478 1647 484 1648
rect 478 1646 479 1647
rect 396 1644 479 1646
rect 396 1643 397 1644
rect 391 1642 397 1643
rect 478 1643 479 1644
rect 483 1643 484 1647
rect 534 1645 535 1649
rect 539 1645 540 1649
rect 534 1644 540 1645
rect 710 1649 716 1650
rect 710 1645 711 1649
rect 715 1645 716 1649
rect 918 1649 924 1650
rect 710 1644 716 1645
rect 718 1647 725 1648
rect 478 1642 484 1643
rect 543 1643 549 1644
rect 543 1642 544 1643
rect 480 1640 544 1642
rect 310 1638 316 1639
rect 543 1639 544 1640
rect 548 1642 549 1643
rect 598 1643 604 1644
rect 598 1642 599 1643
rect 548 1640 599 1642
rect 548 1639 549 1640
rect 543 1638 549 1639
rect 598 1639 599 1640
rect 603 1639 604 1643
rect 718 1643 719 1647
rect 724 1643 725 1647
rect 918 1645 919 1649
rect 923 1645 924 1649
rect 1142 1649 1148 1650
rect 918 1644 924 1645
rect 926 1647 933 1648
rect 718 1642 725 1643
rect 926 1643 927 1647
rect 932 1643 933 1647
rect 1142 1645 1143 1649
rect 1147 1645 1148 1649
rect 1382 1649 1388 1650
rect 1142 1644 1148 1645
rect 1151 1647 1157 1648
rect 926 1642 933 1643
rect 1151 1643 1152 1647
rect 1156 1646 1157 1647
rect 1166 1647 1172 1648
rect 1166 1646 1167 1647
rect 1156 1644 1167 1646
rect 1156 1643 1157 1644
rect 1151 1642 1157 1643
rect 1166 1643 1167 1644
rect 1171 1643 1172 1647
rect 1382 1645 1383 1649
rect 1387 1645 1388 1649
rect 1382 1644 1388 1645
rect 1598 1649 1604 1650
rect 1598 1645 1599 1649
rect 1603 1645 1604 1649
rect 1609 1648 1707 1650
rect 1598 1644 1604 1645
rect 1606 1647 1613 1648
rect 1166 1642 1172 1643
rect 1391 1643 1397 1644
rect 598 1638 604 1639
rect 1391 1639 1392 1643
rect 1396 1642 1397 1643
rect 1422 1643 1428 1644
rect 1422 1642 1423 1643
rect 1396 1640 1423 1642
rect 1396 1639 1397 1640
rect 1391 1638 1397 1639
rect 1422 1639 1423 1640
rect 1427 1639 1428 1643
rect 1606 1643 1607 1647
rect 1612 1643 1613 1647
rect 1606 1642 1613 1643
rect 1630 1645 1636 1646
rect 1630 1641 1631 1645
rect 1635 1641 1636 1645
rect 1630 1640 1636 1641
rect 1670 1643 1676 1644
rect 1422 1638 1428 1639
rect 1670 1639 1671 1643
rect 1675 1639 1676 1643
rect 1670 1638 1676 1639
rect 3190 1643 3196 1644
rect 3190 1639 3191 1643
rect 3195 1639 3196 1643
rect 3190 1638 3196 1639
rect 1694 1636 1700 1637
rect 1694 1632 1695 1636
rect 1699 1632 1700 1636
rect 1694 1631 1700 1632
rect 1894 1636 1900 1637
rect 1894 1632 1895 1636
rect 1899 1632 1900 1636
rect 1894 1631 1900 1632
rect 2126 1636 2132 1637
rect 2126 1632 2127 1636
rect 2131 1632 2132 1636
rect 2126 1631 2132 1632
rect 2366 1636 2372 1637
rect 2366 1632 2367 1636
rect 2371 1632 2372 1636
rect 2366 1631 2372 1632
rect 2614 1636 2620 1637
rect 2614 1632 2615 1636
rect 2619 1632 2620 1636
rect 2614 1631 2620 1632
rect 2870 1636 2876 1637
rect 2870 1632 2871 1636
rect 2875 1632 2876 1636
rect 2870 1631 2876 1632
rect 3134 1636 3140 1637
rect 3134 1632 3135 1636
rect 3139 1632 3140 1636
rect 3134 1631 3140 1632
rect 110 1627 116 1628
rect 110 1623 111 1627
rect 115 1623 116 1627
rect 110 1622 116 1623
rect 1630 1627 1636 1628
rect 1630 1623 1631 1627
rect 1635 1623 1636 1627
rect 1630 1622 1636 1623
rect 134 1620 140 1621
rect 134 1616 135 1620
rect 139 1616 140 1620
rect 134 1615 140 1616
rect 246 1620 252 1621
rect 246 1616 247 1620
rect 251 1616 252 1620
rect 246 1615 252 1616
rect 382 1620 388 1621
rect 382 1616 383 1620
rect 387 1616 388 1620
rect 382 1615 388 1616
rect 534 1620 540 1621
rect 534 1616 535 1620
rect 539 1616 540 1620
rect 534 1615 540 1616
rect 710 1620 716 1621
rect 710 1616 711 1620
rect 715 1616 716 1620
rect 710 1615 716 1616
rect 918 1620 924 1621
rect 918 1616 919 1620
rect 923 1616 924 1620
rect 918 1615 924 1616
rect 1142 1620 1148 1621
rect 1142 1616 1143 1620
rect 1147 1616 1148 1620
rect 1142 1615 1148 1616
rect 1382 1620 1388 1621
rect 1382 1616 1383 1620
rect 1387 1616 1388 1620
rect 1382 1615 1388 1616
rect 1598 1620 1604 1621
rect 1598 1616 1599 1620
rect 1603 1616 1604 1620
rect 1598 1615 1604 1616
rect 2318 1620 2324 1621
rect 2318 1616 2319 1620
rect 2323 1616 2324 1620
rect 2318 1615 2324 1616
rect 2518 1620 2524 1621
rect 2518 1616 2519 1620
rect 2523 1616 2524 1620
rect 2518 1615 2524 1616
rect 2710 1620 2716 1621
rect 2710 1616 2711 1620
rect 2715 1616 2716 1620
rect 2710 1615 2716 1616
rect 2910 1620 2916 1621
rect 2910 1616 2911 1620
rect 2915 1616 2916 1620
rect 2910 1615 2916 1616
rect 3110 1620 3116 1621
rect 3110 1616 3111 1620
rect 3115 1616 3116 1620
rect 3110 1615 3116 1616
rect 1670 1613 1676 1614
rect 1670 1609 1671 1613
rect 1675 1609 1676 1613
rect 1670 1608 1676 1609
rect 3190 1613 3196 1614
rect 3190 1609 3191 1613
rect 3195 1609 3196 1613
rect 3190 1608 3196 1609
rect 134 1600 140 1601
rect 134 1596 135 1600
rect 139 1596 140 1600
rect 134 1595 140 1596
rect 302 1600 308 1601
rect 302 1596 303 1600
rect 307 1596 308 1600
rect 302 1595 308 1596
rect 502 1600 508 1601
rect 502 1596 503 1600
rect 507 1596 508 1600
rect 502 1595 508 1596
rect 694 1600 700 1601
rect 694 1596 695 1600
rect 699 1596 700 1600
rect 694 1595 700 1596
rect 886 1600 892 1601
rect 886 1596 887 1600
rect 891 1596 892 1600
rect 886 1595 892 1596
rect 1062 1600 1068 1601
rect 1062 1596 1063 1600
rect 1067 1596 1068 1600
rect 1062 1595 1068 1596
rect 1238 1600 1244 1601
rect 1238 1596 1239 1600
rect 1243 1596 1244 1600
rect 1238 1595 1244 1596
rect 1414 1600 1420 1601
rect 1414 1596 1415 1600
rect 1419 1596 1420 1600
rect 1414 1595 1420 1596
rect 1590 1600 1596 1601
rect 1590 1596 1591 1600
rect 1595 1596 1596 1600
rect 1590 1595 1596 1596
rect 1670 1595 1676 1596
rect 110 1593 116 1594
rect 110 1589 111 1593
rect 115 1589 116 1593
rect 110 1588 116 1589
rect 1630 1593 1636 1594
rect 1630 1589 1631 1593
rect 1635 1589 1636 1593
rect 1670 1591 1671 1595
rect 1675 1591 1676 1595
rect 3118 1595 3125 1596
rect 1670 1590 1676 1591
rect 2318 1591 2324 1592
rect 1630 1588 1636 1589
rect 2318 1587 2319 1591
rect 2323 1587 2324 1591
rect 2318 1586 2324 1587
rect 2327 1591 2333 1592
rect 2327 1587 2328 1591
rect 2332 1587 2333 1591
rect 2327 1586 2333 1587
rect 2518 1591 2524 1592
rect 2518 1587 2519 1591
rect 2523 1587 2524 1591
rect 2518 1586 2524 1587
rect 2526 1591 2533 1592
rect 2526 1587 2527 1591
rect 2532 1587 2533 1591
rect 2526 1586 2533 1587
rect 2710 1591 2716 1592
rect 2710 1587 2711 1591
rect 2715 1587 2716 1591
rect 2710 1586 2716 1587
rect 2718 1591 2725 1592
rect 2718 1587 2719 1591
rect 2724 1587 2725 1591
rect 2718 1586 2725 1587
rect 2910 1591 2916 1592
rect 2910 1587 2911 1591
rect 2915 1587 2916 1591
rect 2910 1586 2916 1587
rect 2918 1591 2925 1592
rect 2918 1587 2919 1591
rect 2924 1590 2925 1591
rect 3006 1591 3012 1592
rect 3006 1590 3007 1591
rect 2924 1588 3007 1590
rect 2924 1587 2925 1588
rect 2918 1586 2925 1587
rect 3006 1587 3007 1588
rect 3011 1587 3012 1591
rect 3006 1586 3012 1587
rect 3110 1591 3116 1592
rect 3110 1587 3111 1591
rect 3115 1587 3116 1591
rect 3118 1591 3119 1595
rect 3124 1594 3125 1595
rect 3142 1595 3148 1596
rect 3142 1594 3143 1595
rect 3124 1592 3143 1594
rect 3124 1591 3125 1592
rect 3118 1590 3125 1591
rect 3142 1591 3143 1592
rect 3147 1591 3148 1595
rect 3142 1590 3148 1591
rect 3190 1595 3196 1596
rect 3190 1591 3191 1595
rect 3195 1591 3196 1595
rect 3190 1590 3196 1591
rect 3110 1586 3116 1587
rect 2290 1583 2296 1584
rect 2270 1581 2276 1582
rect 478 1579 484 1580
rect 110 1575 116 1576
rect 110 1571 111 1575
rect 115 1571 116 1575
rect 142 1575 149 1576
rect 110 1570 116 1571
rect 134 1571 140 1572
rect 134 1567 135 1571
rect 139 1567 140 1571
rect 142 1571 143 1575
rect 148 1571 149 1575
rect 310 1575 317 1576
rect 142 1570 149 1571
rect 302 1571 308 1572
rect 134 1566 140 1567
rect 302 1567 303 1571
rect 307 1567 308 1571
rect 310 1571 311 1575
rect 316 1571 317 1575
rect 478 1575 479 1579
rect 483 1578 484 1579
rect 1166 1579 1172 1580
rect 483 1576 514 1578
rect 483 1575 484 1576
rect 478 1574 484 1575
rect 511 1575 517 1576
rect 310 1570 317 1571
rect 502 1571 508 1572
rect 302 1566 308 1567
rect 502 1567 503 1571
rect 507 1567 508 1571
rect 511 1571 512 1575
rect 516 1571 517 1575
rect 703 1575 709 1576
rect 511 1570 517 1571
rect 694 1571 700 1572
rect 502 1566 508 1567
rect 694 1567 695 1571
rect 699 1567 700 1571
rect 703 1571 704 1575
rect 708 1574 709 1575
rect 718 1575 724 1576
rect 718 1574 719 1575
rect 708 1572 719 1574
rect 708 1571 709 1572
rect 703 1570 709 1571
rect 718 1571 719 1572
rect 723 1571 724 1575
rect 1070 1575 1077 1576
rect 718 1570 724 1571
rect 886 1571 892 1572
rect 694 1566 700 1567
rect 886 1567 887 1571
rect 891 1567 892 1571
rect 886 1566 892 1567
rect 894 1571 901 1572
rect 894 1567 895 1571
rect 900 1570 901 1571
rect 926 1571 932 1572
rect 926 1570 927 1571
rect 900 1568 927 1570
rect 900 1567 901 1568
rect 894 1566 901 1567
rect 926 1567 927 1568
rect 931 1567 932 1571
rect 926 1566 932 1567
rect 1062 1571 1068 1572
rect 1062 1567 1063 1571
rect 1067 1567 1068 1571
rect 1070 1571 1071 1575
rect 1076 1571 1077 1575
rect 1166 1575 1167 1579
rect 1171 1578 1172 1579
rect 1171 1576 1250 1578
rect 1670 1577 1676 1578
rect 1171 1575 1172 1576
rect 1166 1574 1172 1575
rect 1247 1575 1253 1576
rect 1070 1570 1077 1571
rect 1238 1571 1244 1572
rect 1062 1566 1068 1567
rect 1238 1567 1239 1571
rect 1243 1567 1244 1571
rect 1247 1571 1248 1575
rect 1252 1574 1253 1575
rect 1286 1575 1292 1576
rect 1286 1574 1287 1575
rect 1252 1572 1287 1574
rect 1252 1571 1253 1572
rect 1247 1570 1253 1571
rect 1286 1571 1287 1572
rect 1291 1571 1292 1575
rect 1630 1575 1636 1576
rect 1286 1570 1292 1571
rect 1414 1571 1420 1572
rect 1238 1566 1244 1567
rect 1414 1567 1415 1571
rect 1419 1567 1420 1571
rect 1414 1566 1420 1567
rect 1422 1571 1429 1572
rect 1422 1567 1423 1571
rect 1428 1567 1429 1571
rect 1422 1566 1429 1567
rect 1590 1571 1596 1572
rect 1590 1567 1591 1571
rect 1595 1567 1596 1571
rect 1590 1566 1596 1567
rect 1599 1571 1605 1572
rect 1599 1567 1600 1571
rect 1604 1567 1605 1571
rect 1630 1571 1631 1575
rect 1635 1571 1636 1575
rect 1670 1573 1671 1577
rect 1675 1573 1676 1577
rect 2270 1577 2271 1581
rect 2275 1577 2276 1581
rect 2290 1580 2291 1583
rect 2270 1576 2276 1577
rect 2279 1579 2291 1580
rect 2295 1582 2296 1583
rect 2328 1582 2330 1586
rect 2295 1580 2330 1582
rect 2414 1581 2420 1582
rect 2295 1579 2296 1580
rect 2279 1575 2280 1579
rect 2284 1578 2296 1579
rect 2284 1575 2285 1578
rect 2414 1577 2415 1581
rect 2419 1577 2420 1581
rect 2414 1576 2420 1577
rect 2558 1581 2564 1582
rect 2558 1577 2559 1581
rect 2563 1577 2564 1581
rect 2558 1576 2564 1577
rect 2694 1581 2700 1582
rect 2694 1577 2695 1581
rect 2699 1577 2700 1581
rect 2694 1576 2700 1577
rect 2838 1581 2844 1582
rect 2838 1577 2839 1581
rect 2843 1577 2844 1581
rect 2838 1576 2844 1577
rect 2982 1581 2988 1582
rect 2982 1577 2983 1581
rect 2987 1577 2988 1581
rect 2982 1576 2988 1577
rect 3190 1577 3196 1578
rect 2279 1574 2285 1575
rect 2398 1575 2404 1576
rect 1670 1572 1676 1573
rect 1630 1570 1636 1571
rect 2398 1571 2399 1575
rect 2403 1574 2404 1575
rect 2423 1575 2429 1576
rect 2423 1574 2424 1575
rect 2403 1572 2424 1574
rect 2403 1571 2404 1572
rect 2398 1570 2404 1571
rect 2423 1571 2424 1572
rect 2428 1571 2429 1575
rect 2423 1570 2429 1571
rect 2526 1575 2532 1576
rect 2526 1571 2527 1575
rect 2531 1574 2532 1575
rect 2567 1575 2573 1576
rect 2567 1574 2568 1575
rect 2531 1572 2568 1574
rect 2531 1571 2532 1572
rect 2526 1570 2532 1571
rect 2567 1571 2568 1572
rect 2572 1571 2573 1575
rect 2567 1570 2573 1571
rect 2662 1575 2668 1576
rect 2662 1571 2663 1575
rect 2667 1574 2668 1575
rect 2703 1575 2709 1576
rect 2703 1574 2704 1575
rect 2667 1572 2704 1574
rect 2667 1571 2668 1572
rect 2662 1570 2668 1571
rect 2703 1571 2704 1572
rect 2708 1574 2709 1575
rect 2718 1575 2724 1576
rect 2718 1574 2719 1575
rect 2708 1572 2719 1574
rect 2708 1571 2709 1572
rect 2703 1570 2709 1571
rect 2718 1571 2719 1572
rect 2723 1571 2724 1575
rect 2718 1570 2724 1571
rect 2847 1575 2853 1576
rect 2847 1571 2848 1575
rect 2852 1574 2853 1575
rect 2918 1575 2924 1576
rect 2918 1574 2919 1575
rect 2852 1572 2919 1574
rect 2852 1571 2853 1572
rect 2847 1570 2853 1571
rect 2918 1571 2919 1572
rect 2923 1571 2924 1575
rect 2918 1570 2924 1571
rect 2991 1575 2997 1576
rect 2991 1571 2992 1575
rect 2996 1574 2997 1575
rect 3006 1575 3012 1576
rect 3006 1574 3007 1575
rect 2996 1572 3007 1574
rect 2996 1571 2997 1572
rect 2991 1570 2997 1571
rect 3006 1571 3007 1572
rect 3011 1571 3012 1575
rect 3190 1573 3191 1577
rect 3195 1573 3196 1577
rect 3190 1572 3196 1573
rect 3006 1570 3012 1571
rect 1599 1566 1605 1567
rect 1670 1559 1676 1560
rect 1670 1555 1671 1559
rect 1675 1555 1676 1559
rect 1670 1554 1676 1555
rect 3190 1559 3196 1560
rect 3190 1555 3191 1559
rect 3195 1555 3196 1559
rect 3190 1554 3196 1555
rect 2270 1552 2276 1553
rect 678 1549 684 1550
rect 110 1545 116 1546
rect 110 1541 111 1545
rect 115 1541 116 1545
rect 678 1545 679 1549
rect 683 1545 684 1549
rect 806 1549 812 1550
rect 678 1544 684 1545
rect 687 1547 693 1548
rect 687 1543 688 1547
rect 692 1546 693 1547
rect 718 1547 724 1548
rect 718 1546 719 1547
rect 692 1544 719 1546
rect 692 1543 693 1544
rect 687 1542 693 1543
rect 718 1543 719 1544
rect 723 1543 724 1547
rect 806 1545 807 1549
rect 811 1545 812 1549
rect 806 1544 812 1545
rect 926 1549 932 1550
rect 926 1545 927 1549
rect 931 1545 932 1549
rect 926 1544 932 1545
rect 1046 1549 1052 1550
rect 1046 1545 1047 1549
rect 1051 1545 1052 1549
rect 1166 1549 1172 1550
rect 1046 1544 1052 1545
rect 1055 1547 1061 1548
rect 718 1542 724 1543
rect 815 1543 821 1544
rect 110 1540 116 1541
rect 815 1539 816 1543
rect 820 1542 821 1543
rect 838 1543 844 1544
rect 838 1542 839 1543
rect 820 1540 839 1542
rect 820 1539 821 1540
rect 815 1538 821 1539
rect 838 1539 839 1540
rect 843 1542 844 1543
rect 894 1543 900 1544
rect 894 1542 895 1543
rect 843 1540 895 1542
rect 843 1539 844 1540
rect 838 1538 844 1539
rect 894 1539 895 1540
rect 899 1542 900 1543
rect 935 1543 941 1544
rect 935 1542 936 1543
rect 899 1540 936 1542
rect 899 1539 900 1540
rect 894 1538 900 1539
rect 935 1539 936 1540
rect 940 1542 941 1543
rect 1055 1543 1056 1547
rect 1060 1546 1061 1547
rect 1070 1547 1076 1548
rect 1070 1546 1071 1547
rect 1060 1544 1071 1546
rect 1060 1543 1061 1544
rect 1055 1542 1061 1543
rect 1070 1543 1071 1544
rect 1075 1543 1076 1547
rect 1166 1545 1167 1549
rect 1171 1545 1172 1549
rect 1278 1549 1284 1550
rect 1166 1544 1172 1545
rect 1174 1547 1181 1548
rect 1070 1542 1076 1543
rect 1174 1543 1175 1547
rect 1180 1546 1181 1547
rect 1190 1547 1196 1548
rect 1190 1546 1191 1547
rect 1180 1544 1191 1546
rect 1180 1543 1181 1544
rect 1174 1542 1181 1543
rect 1190 1543 1191 1544
rect 1195 1543 1196 1547
rect 1278 1545 1279 1549
rect 1283 1545 1284 1549
rect 1398 1549 1404 1550
rect 1278 1544 1284 1545
rect 1286 1547 1293 1548
rect 1190 1542 1196 1543
rect 1286 1543 1287 1547
rect 1292 1543 1293 1547
rect 1398 1545 1399 1549
rect 1403 1545 1404 1549
rect 1398 1544 1404 1545
rect 1518 1549 1524 1550
rect 1518 1545 1519 1549
rect 1523 1545 1524 1549
rect 2270 1548 2271 1552
rect 2275 1548 2276 1552
rect 2270 1547 2276 1548
rect 2414 1552 2420 1553
rect 2414 1548 2415 1552
rect 2419 1548 2420 1552
rect 2414 1547 2420 1548
rect 2558 1552 2564 1553
rect 2558 1548 2559 1552
rect 2563 1548 2564 1552
rect 2558 1547 2564 1548
rect 2694 1552 2700 1553
rect 2694 1548 2695 1552
rect 2699 1548 2700 1552
rect 2694 1547 2700 1548
rect 2838 1552 2844 1553
rect 2838 1548 2839 1552
rect 2843 1548 2844 1552
rect 2838 1547 2844 1548
rect 2982 1552 2988 1553
rect 2982 1548 2983 1552
rect 2987 1548 2988 1552
rect 2982 1547 2988 1548
rect 1518 1544 1524 1545
rect 1630 1545 1636 1546
rect 1286 1542 1293 1543
rect 1406 1543 1413 1544
rect 940 1540 1058 1542
rect 940 1539 941 1540
rect 935 1538 941 1539
rect 1406 1539 1407 1543
rect 1412 1542 1413 1543
rect 1422 1543 1428 1544
rect 1422 1542 1423 1543
rect 1412 1540 1423 1542
rect 1412 1539 1413 1540
rect 1406 1538 1413 1539
rect 1422 1539 1423 1540
rect 1427 1542 1428 1543
rect 1527 1543 1533 1544
rect 1527 1542 1528 1543
rect 1427 1540 1528 1542
rect 1427 1539 1428 1540
rect 1422 1538 1428 1539
rect 1527 1539 1528 1540
rect 1532 1542 1533 1543
rect 1598 1543 1604 1544
rect 1598 1542 1599 1543
rect 1532 1540 1599 1542
rect 1532 1539 1533 1540
rect 1527 1538 1533 1539
rect 1598 1539 1599 1540
rect 1603 1539 1604 1543
rect 1630 1541 1631 1545
rect 1635 1541 1636 1545
rect 1630 1540 1636 1541
rect 1598 1538 1604 1539
rect 2166 1532 2172 1533
rect 2166 1528 2167 1532
rect 2171 1528 2172 1532
rect 110 1527 116 1528
rect 110 1523 111 1527
rect 115 1523 116 1527
rect 110 1522 116 1523
rect 1630 1527 1636 1528
rect 2166 1527 2172 1528
rect 2278 1532 2284 1533
rect 2278 1528 2279 1532
rect 2283 1528 2284 1532
rect 2278 1527 2284 1528
rect 2390 1532 2396 1533
rect 2390 1528 2391 1532
rect 2395 1528 2396 1532
rect 2390 1527 2396 1528
rect 2502 1532 2508 1533
rect 2502 1528 2503 1532
rect 2507 1528 2508 1532
rect 2502 1527 2508 1528
rect 2614 1532 2620 1533
rect 2614 1528 2615 1532
rect 2619 1528 2620 1532
rect 2614 1527 2620 1528
rect 2734 1532 2740 1533
rect 2734 1528 2735 1532
rect 2739 1528 2740 1532
rect 2734 1527 2740 1528
rect 2854 1532 2860 1533
rect 2854 1528 2855 1532
rect 2859 1528 2860 1532
rect 2854 1527 2860 1528
rect 2982 1532 2988 1533
rect 2982 1528 2983 1532
rect 2987 1528 2988 1532
rect 2982 1527 2988 1528
rect 3110 1532 3116 1533
rect 3110 1528 3111 1532
rect 3115 1528 3116 1532
rect 3110 1527 3116 1528
rect 1630 1523 1631 1527
rect 1635 1523 1636 1527
rect 1630 1522 1636 1523
rect 1670 1525 1676 1526
rect 1670 1521 1671 1525
rect 1675 1521 1676 1525
rect 678 1520 684 1521
rect 678 1516 679 1520
rect 683 1516 684 1520
rect 678 1515 684 1516
rect 806 1520 812 1521
rect 806 1516 807 1520
rect 811 1516 812 1520
rect 806 1515 812 1516
rect 926 1520 932 1521
rect 926 1516 927 1520
rect 931 1516 932 1520
rect 926 1515 932 1516
rect 1046 1520 1052 1521
rect 1046 1516 1047 1520
rect 1051 1516 1052 1520
rect 1046 1515 1052 1516
rect 1166 1520 1172 1521
rect 1166 1516 1167 1520
rect 1171 1516 1172 1520
rect 1166 1515 1172 1516
rect 1278 1520 1284 1521
rect 1278 1516 1279 1520
rect 1283 1516 1284 1520
rect 1278 1515 1284 1516
rect 1398 1520 1404 1521
rect 1398 1516 1399 1520
rect 1403 1516 1404 1520
rect 1398 1515 1404 1516
rect 1518 1520 1524 1521
rect 1670 1520 1676 1521
rect 3190 1525 3196 1526
rect 3190 1521 3191 1525
rect 3195 1521 3196 1525
rect 3190 1520 3196 1521
rect 1518 1516 1519 1520
rect 1523 1516 1524 1520
rect 1518 1515 1524 1516
rect 2526 1511 2532 1512
rect 1670 1507 1676 1508
rect 1670 1503 1671 1507
rect 1675 1503 1676 1507
rect 2287 1507 2296 1508
rect 1670 1502 1676 1503
rect 2166 1503 2172 1504
rect 574 1500 580 1501
rect 574 1496 575 1500
rect 579 1496 580 1500
rect 574 1495 580 1496
rect 702 1500 708 1501
rect 702 1496 703 1500
rect 707 1496 708 1500
rect 702 1495 708 1496
rect 830 1500 836 1501
rect 830 1496 831 1500
rect 835 1496 836 1500
rect 830 1495 836 1496
rect 950 1500 956 1501
rect 950 1496 951 1500
rect 955 1496 956 1500
rect 950 1495 956 1496
rect 1070 1500 1076 1501
rect 1070 1496 1071 1500
rect 1075 1496 1076 1500
rect 1070 1495 1076 1496
rect 1182 1500 1188 1501
rect 1182 1496 1183 1500
rect 1187 1496 1188 1500
rect 1182 1495 1188 1496
rect 1294 1500 1300 1501
rect 1294 1496 1295 1500
rect 1299 1496 1300 1500
rect 1294 1495 1300 1496
rect 1414 1500 1420 1501
rect 1414 1496 1415 1500
rect 1419 1496 1420 1500
rect 2166 1499 2167 1503
rect 2171 1499 2172 1503
rect 2166 1498 2172 1499
rect 2175 1503 2181 1504
rect 2175 1499 2176 1503
rect 2180 1499 2181 1503
rect 2175 1498 2181 1499
rect 2278 1503 2284 1504
rect 2278 1499 2279 1503
rect 2283 1499 2284 1503
rect 2287 1503 2288 1507
rect 2295 1503 2296 1507
rect 2398 1507 2405 1508
rect 2287 1502 2296 1503
rect 2390 1503 2396 1504
rect 2278 1498 2284 1499
rect 2390 1499 2391 1503
rect 2395 1499 2396 1503
rect 2398 1503 2399 1507
rect 2404 1503 2405 1507
rect 2526 1507 2527 1511
rect 2531 1510 2532 1511
rect 2531 1508 2627 1510
rect 2664 1508 2746 1510
rect 2531 1507 2532 1508
rect 2526 1506 2532 1507
rect 2623 1507 2629 1508
rect 2398 1502 2405 1503
rect 2502 1503 2508 1504
rect 2390 1498 2396 1499
rect 2502 1499 2503 1503
rect 2507 1499 2508 1503
rect 2502 1498 2508 1499
rect 2511 1503 2517 1504
rect 2511 1499 2512 1503
rect 2516 1502 2517 1503
rect 2526 1503 2532 1504
rect 2526 1502 2527 1503
rect 2516 1500 2527 1502
rect 2516 1499 2517 1500
rect 2511 1498 2517 1499
rect 2526 1499 2527 1500
rect 2531 1499 2532 1503
rect 2526 1498 2532 1499
rect 2614 1503 2620 1504
rect 2614 1499 2615 1503
rect 2619 1499 2620 1503
rect 2623 1503 2624 1507
rect 2628 1506 2629 1507
rect 2662 1507 2668 1508
rect 2662 1506 2663 1507
rect 2628 1504 2663 1506
rect 2628 1503 2629 1504
rect 2623 1502 2629 1503
rect 2662 1503 2663 1504
rect 2667 1503 2668 1507
rect 2743 1507 2749 1508
rect 2662 1502 2668 1503
rect 2734 1503 2740 1504
rect 2614 1498 2620 1499
rect 2734 1499 2735 1503
rect 2739 1499 2740 1503
rect 2743 1503 2744 1507
rect 2748 1506 2749 1507
rect 2806 1507 2812 1508
rect 2806 1506 2807 1507
rect 2748 1504 2807 1506
rect 2748 1503 2749 1504
rect 2743 1502 2749 1503
rect 2806 1503 2807 1504
rect 2811 1503 2812 1507
rect 2862 1507 2869 1508
rect 2806 1502 2812 1503
rect 2854 1503 2860 1504
rect 2734 1498 2740 1499
rect 2854 1499 2855 1503
rect 2859 1499 2860 1503
rect 2862 1503 2863 1507
rect 2868 1506 2869 1507
rect 2918 1507 2924 1508
rect 2918 1506 2919 1507
rect 2868 1504 2919 1506
rect 2868 1503 2869 1504
rect 2862 1502 2869 1503
rect 2918 1503 2919 1504
rect 2923 1503 2924 1507
rect 3118 1507 3125 1508
rect 2918 1502 2924 1503
rect 2982 1503 2988 1504
rect 2854 1498 2860 1499
rect 2982 1499 2983 1503
rect 2987 1499 2988 1503
rect 2982 1498 2988 1499
rect 2991 1503 2997 1504
rect 2991 1499 2992 1503
rect 2996 1502 2997 1503
rect 3006 1503 3012 1504
rect 3006 1502 3007 1503
rect 2996 1500 3007 1502
rect 2996 1499 2997 1500
rect 2991 1498 2997 1499
rect 3006 1499 3007 1500
rect 3011 1499 3012 1503
rect 3006 1498 3012 1499
rect 3110 1503 3116 1504
rect 3110 1499 3111 1503
rect 3115 1499 3116 1503
rect 3118 1503 3119 1507
rect 3124 1503 3125 1507
rect 3118 1502 3125 1503
rect 3190 1507 3196 1508
rect 3190 1503 3191 1507
rect 3195 1503 3196 1507
rect 3190 1502 3196 1503
rect 3110 1498 3116 1499
rect 1414 1495 1420 1496
rect 2106 1495 2112 1496
rect 110 1493 116 1494
rect 110 1489 111 1493
rect 115 1489 116 1493
rect 110 1488 116 1489
rect 1630 1493 1636 1494
rect 1630 1489 1631 1493
rect 1635 1489 1636 1493
rect 2106 1491 2107 1495
rect 2111 1494 2112 1495
rect 2177 1494 2179 1498
rect 2111 1492 2179 1494
rect 2398 1495 2404 1496
rect 2111 1491 2112 1492
rect 2106 1490 2112 1491
rect 2398 1491 2399 1495
rect 2403 1494 2404 1495
rect 2486 1495 2492 1496
rect 2486 1494 2487 1495
rect 2403 1492 2487 1494
rect 2403 1491 2404 1492
rect 2398 1490 2404 1491
rect 2486 1491 2487 1492
rect 2491 1494 2492 1495
rect 2512 1494 2514 1498
rect 2491 1492 2522 1494
rect 2491 1491 2492 1492
rect 2486 1490 2492 1491
rect 1630 1488 1636 1489
rect 2086 1489 2092 1490
rect 1670 1485 1676 1486
rect 1670 1481 1671 1485
rect 1675 1481 1676 1485
rect 2086 1485 2087 1489
rect 2091 1485 2092 1489
rect 2086 1484 2092 1485
rect 2230 1489 2236 1490
rect 2230 1485 2231 1489
rect 2235 1485 2236 1489
rect 2374 1489 2380 1490
rect 2230 1484 2236 1485
rect 2238 1487 2245 1488
rect 1670 1480 1676 1481
rect 2095 1483 2101 1484
rect 1286 1479 1292 1480
rect 110 1475 116 1476
rect 110 1471 111 1475
rect 115 1471 116 1475
rect 1286 1475 1287 1479
rect 1291 1478 1292 1479
rect 1406 1479 1412 1480
rect 1406 1478 1407 1479
rect 1291 1476 1306 1478
rect 1399 1476 1407 1478
rect 1291 1475 1292 1476
rect 1286 1474 1292 1475
rect 1303 1475 1309 1476
rect 110 1470 116 1471
rect 574 1471 580 1472
rect 574 1467 575 1471
rect 579 1467 580 1471
rect 574 1466 580 1467
rect 583 1471 592 1472
rect 583 1467 584 1471
rect 591 1467 592 1471
rect 583 1466 592 1467
rect 702 1471 708 1472
rect 702 1467 703 1471
rect 707 1467 708 1471
rect 702 1466 708 1467
rect 711 1471 717 1472
rect 711 1467 712 1471
rect 716 1470 717 1471
rect 734 1471 740 1472
rect 734 1470 735 1471
rect 716 1468 735 1470
rect 716 1467 717 1468
rect 711 1466 717 1467
rect 734 1467 735 1468
rect 739 1467 740 1471
rect 734 1466 740 1467
rect 830 1471 836 1472
rect 830 1467 831 1471
rect 835 1467 836 1471
rect 830 1466 836 1467
rect 838 1471 845 1472
rect 838 1467 839 1471
rect 844 1467 845 1471
rect 838 1466 845 1467
rect 950 1471 956 1472
rect 950 1467 951 1471
rect 955 1467 956 1471
rect 950 1466 956 1467
rect 958 1471 965 1472
rect 958 1467 959 1471
rect 964 1467 965 1471
rect 958 1466 965 1467
rect 1070 1471 1076 1472
rect 1070 1467 1071 1471
rect 1075 1467 1076 1471
rect 1070 1466 1076 1467
rect 1078 1471 1085 1472
rect 1078 1467 1079 1471
rect 1084 1467 1085 1471
rect 1078 1466 1085 1467
rect 1182 1471 1188 1472
rect 1182 1467 1183 1471
rect 1187 1467 1188 1471
rect 1182 1466 1188 1467
rect 1190 1471 1197 1472
rect 1190 1467 1191 1471
rect 1196 1467 1197 1471
rect 1190 1466 1197 1467
rect 1294 1471 1300 1472
rect 1294 1467 1295 1471
rect 1299 1467 1300 1471
rect 1303 1471 1304 1475
rect 1308 1474 1309 1475
rect 1318 1475 1324 1476
rect 1318 1474 1319 1475
rect 1308 1472 1319 1474
rect 1308 1471 1309 1472
rect 1303 1470 1309 1471
rect 1318 1471 1319 1472
rect 1323 1474 1324 1475
rect 1399 1474 1401 1476
rect 1406 1475 1407 1476
rect 1411 1478 1412 1479
rect 2095 1479 2096 1483
rect 2100 1482 2101 1483
rect 2106 1483 2112 1484
rect 2106 1482 2107 1483
rect 2100 1480 2107 1482
rect 2100 1479 2101 1480
rect 2095 1478 2101 1479
rect 2106 1479 2107 1480
rect 2111 1479 2112 1483
rect 2238 1483 2239 1487
rect 2244 1486 2245 1487
rect 2290 1487 2296 1488
rect 2290 1486 2291 1487
rect 2244 1484 2291 1486
rect 2244 1483 2245 1484
rect 2238 1482 2245 1483
rect 2290 1483 2291 1484
rect 2295 1483 2296 1487
rect 2374 1485 2375 1489
rect 2379 1485 2380 1489
rect 2510 1489 2516 1490
rect 2374 1484 2380 1485
rect 2383 1487 2389 1488
rect 2290 1482 2296 1483
rect 2383 1483 2384 1487
rect 2388 1486 2389 1487
rect 2398 1487 2404 1488
rect 2398 1486 2399 1487
rect 2388 1484 2399 1486
rect 2388 1483 2389 1484
rect 2383 1482 2389 1483
rect 2398 1483 2399 1484
rect 2403 1483 2404 1487
rect 2510 1485 2511 1489
rect 2515 1485 2516 1489
rect 2520 1488 2522 1492
rect 2654 1489 2660 1490
rect 2510 1484 2516 1485
rect 2519 1487 2525 1488
rect 2398 1482 2404 1483
rect 2519 1483 2520 1487
rect 2524 1483 2525 1487
rect 2654 1485 2655 1489
rect 2659 1485 2660 1489
rect 2798 1489 2804 1490
rect 2654 1484 2660 1485
rect 2662 1487 2669 1488
rect 2519 1482 2525 1483
rect 2662 1483 2663 1487
rect 2668 1483 2669 1487
rect 2798 1485 2799 1489
rect 2803 1485 2804 1489
rect 2798 1484 2804 1485
rect 2806 1487 2813 1488
rect 2662 1482 2669 1483
rect 2806 1483 2807 1487
rect 2812 1486 2813 1487
rect 2812 1484 2841 1486
rect 3190 1485 3196 1486
rect 2812 1483 2813 1484
rect 2806 1482 2813 1483
rect 2839 1482 2841 1484
rect 2862 1483 2868 1484
rect 2862 1482 2863 1483
rect 2839 1480 2863 1482
rect 2106 1478 2112 1479
rect 2862 1479 2863 1480
rect 2867 1479 2868 1483
rect 3190 1481 3191 1485
rect 3195 1481 3196 1485
rect 3190 1480 3196 1481
rect 2862 1478 2868 1479
rect 1411 1476 1427 1478
rect 1411 1475 1412 1476
rect 1406 1474 1412 1475
rect 1423 1475 1429 1476
rect 1323 1472 1401 1474
rect 1323 1471 1324 1472
rect 1318 1470 1324 1471
rect 1414 1471 1420 1472
rect 1294 1466 1300 1467
rect 1414 1467 1415 1471
rect 1419 1467 1420 1471
rect 1423 1471 1424 1475
rect 1428 1471 1429 1475
rect 1423 1470 1429 1471
rect 1630 1475 1636 1476
rect 1630 1471 1631 1475
rect 1635 1471 1636 1475
rect 1630 1470 1636 1471
rect 1414 1466 1420 1467
rect 1670 1467 1676 1468
rect 1670 1463 1671 1467
rect 1675 1463 1676 1467
rect 1670 1462 1676 1463
rect 3190 1467 3196 1468
rect 3190 1463 3191 1467
rect 3195 1463 3196 1467
rect 3190 1462 3196 1463
rect 2086 1460 2092 1461
rect 2086 1456 2087 1460
rect 2091 1456 2092 1460
rect 2086 1455 2092 1456
rect 2230 1460 2236 1461
rect 2230 1456 2231 1460
rect 2235 1456 2236 1460
rect 2230 1455 2236 1456
rect 2374 1460 2380 1461
rect 2374 1456 2375 1460
rect 2379 1456 2380 1460
rect 2374 1455 2380 1456
rect 2510 1460 2516 1461
rect 2510 1456 2511 1460
rect 2515 1456 2516 1460
rect 2510 1455 2516 1456
rect 2654 1460 2660 1461
rect 2654 1456 2655 1460
rect 2659 1456 2660 1460
rect 2654 1455 2660 1456
rect 2798 1460 2804 1461
rect 2798 1456 2799 1460
rect 2803 1456 2804 1460
rect 2798 1455 2804 1456
rect 478 1449 484 1450
rect 110 1445 116 1446
rect 110 1441 111 1445
rect 115 1441 116 1445
rect 478 1445 479 1449
rect 483 1445 484 1449
rect 478 1444 484 1445
rect 606 1449 612 1450
rect 606 1445 607 1449
rect 611 1445 612 1449
rect 606 1444 612 1445
rect 726 1449 732 1450
rect 726 1445 727 1449
rect 731 1445 732 1449
rect 726 1444 732 1445
rect 846 1449 852 1450
rect 846 1445 847 1449
rect 851 1445 852 1449
rect 846 1444 852 1445
rect 966 1449 972 1450
rect 966 1445 967 1449
rect 971 1445 972 1449
rect 1078 1449 1084 1450
rect 966 1444 972 1445
rect 975 1447 981 1448
rect 110 1440 116 1441
rect 487 1443 493 1444
rect 487 1439 488 1443
rect 492 1442 493 1443
rect 586 1443 592 1444
rect 586 1442 587 1443
rect 492 1440 587 1442
rect 492 1439 493 1440
rect 487 1438 493 1439
rect 586 1439 587 1440
rect 591 1442 592 1443
rect 615 1443 621 1444
rect 615 1442 616 1443
rect 591 1440 616 1442
rect 591 1439 592 1440
rect 586 1438 592 1439
rect 615 1439 616 1440
rect 620 1442 621 1443
rect 634 1443 640 1444
rect 634 1442 635 1443
rect 620 1440 635 1442
rect 620 1439 621 1440
rect 615 1438 621 1439
rect 634 1439 635 1440
rect 639 1439 640 1443
rect 634 1438 640 1439
rect 734 1443 741 1444
rect 734 1439 735 1443
rect 740 1442 741 1443
rect 838 1443 844 1444
rect 838 1442 839 1443
rect 740 1440 839 1442
rect 740 1439 741 1440
rect 734 1438 741 1439
rect 838 1439 839 1440
rect 843 1442 844 1443
rect 855 1443 861 1444
rect 855 1442 856 1443
rect 843 1440 856 1442
rect 843 1439 844 1440
rect 838 1438 844 1439
rect 855 1439 856 1440
rect 860 1442 861 1443
rect 886 1443 892 1444
rect 886 1442 887 1443
rect 860 1440 887 1442
rect 860 1439 861 1440
rect 855 1438 861 1439
rect 886 1439 887 1440
rect 891 1442 892 1443
rect 958 1443 964 1444
rect 958 1442 959 1443
rect 891 1440 959 1442
rect 891 1439 892 1440
rect 886 1438 892 1439
rect 958 1439 959 1440
rect 963 1442 964 1443
rect 975 1443 976 1447
rect 980 1443 981 1447
rect 1078 1445 1079 1449
rect 1083 1445 1084 1449
rect 1078 1444 1084 1445
rect 1190 1449 1196 1450
rect 1190 1445 1191 1449
rect 1195 1445 1196 1449
rect 1310 1449 1316 1450
rect 1190 1444 1196 1445
rect 1198 1447 1205 1448
rect 975 1442 981 1443
rect 1086 1443 1093 1444
rect 963 1440 978 1442
rect 963 1439 964 1440
rect 958 1438 964 1439
rect 1086 1439 1087 1443
rect 1092 1442 1093 1443
rect 1102 1443 1108 1444
rect 1102 1442 1103 1443
rect 1092 1440 1103 1442
rect 1092 1439 1093 1440
rect 1086 1438 1093 1439
rect 1102 1439 1103 1440
rect 1107 1442 1108 1443
rect 1198 1443 1199 1447
rect 1204 1443 1205 1447
rect 1310 1445 1311 1449
rect 1315 1445 1316 1449
rect 1310 1444 1316 1445
rect 1318 1447 1325 1448
rect 1198 1442 1205 1443
rect 1318 1443 1319 1447
rect 1324 1443 1325 1447
rect 1318 1442 1325 1443
rect 1630 1445 1636 1446
rect 1107 1440 1202 1442
rect 1630 1441 1631 1445
rect 1635 1441 1636 1445
rect 1630 1440 1636 1441
rect 1982 1444 1988 1445
rect 1982 1440 1983 1444
rect 1987 1440 1988 1444
rect 1107 1439 1108 1440
rect 1982 1439 1988 1440
rect 2094 1444 2100 1445
rect 2094 1440 2095 1444
rect 2099 1440 2100 1444
rect 2094 1439 2100 1440
rect 2206 1444 2212 1445
rect 2206 1440 2207 1444
rect 2211 1440 2212 1444
rect 2206 1439 2212 1440
rect 2334 1444 2340 1445
rect 2334 1440 2335 1444
rect 2339 1440 2340 1444
rect 2334 1439 2340 1440
rect 2478 1444 2484 1445
rect 2478 1440 2479 1444
rect 2483 1440 2484 1444
rect 2478 1439 2484 1440
rect 2638 1444 2644 1445
rect 2638 1440 2639 1444
rect 2643 1440 2644 1444
rect 2638 1439 2644 1440
rect 2814 1444 2820 1445
rect 2814 1440 2815 1444
rect 2819 1440 2820 1444
rect 2814 1439 2820 1440
rect 2998 1444 3004 1445
rect 2998 1440 2999 1444
rect 3003 1440 3004 1444
rect 2998 1439 3004 1440
rect 3158 1444 3164 1445
rect 3158 1440 3159 1444
rect 3163 1440 3164 1444
rect 3158 1439 3164 1440
rect 1102 1438 1108 1439
rect 1670 1437 1676 1438
rect 1670 1433 1671 1437
rect 1675 1433 1676 1437
rect 1670 1432 1676 1433
rect 3190 1437 3196 1438
rect 3190 1433 3191 1437
rect 3195 1433 3196 1437
rect 3190 1432 3196 1433
rect 110 1427 116 1428
rect 110 1423 111 1427
rect 115 1423 116 1427
rect 110 1422 116 1423
rect 1630 1427 1636 1428
rect 1630 1423 1631 1427
rect 1635 1423 1636 1427
rect 1630 1422 1636 1423
rect 2238 1423 2244 1424
rect 2238 1422 2239 1423
rect 2103 1421 2109 1422
rect 478 1420 484 1421
rect 478 1416 479 1420
rect 483 1416 484 1420
rect 478 1415 484 1416
rect 606 1420 612 1421
rect 606 1416 607 1420
rect 611 1416 612 1420
rect 606 1415 612 1416
rect 726 1420 732 1421
rect 726 1416 727 1420
rect 731 1416 732 1420
rect 726 1415 732 1416
rect 846 1420 852 1421
rect 846 1416 847 1420
rect 851 1416 852 1420
rect 846 1415 852 1416
rect 966 1420 972 1421
rect 966 1416 967 1420
rect 971 1416 972 1420
rect 966 1415 972 1416
rect 1078 1420 1084 1421
rect 1078 1416 1079 1420
rect 1083 1416 1084 1420
rect 1078 1415 1084 1416
rect 1190 1420 1196 1421
rect 1190 1416 1191 1420
rect 1195 1416 1196 1420
rect 1190 1415 1196 1416
rect 1310 1420 1316 1421
rect 1310 1416 1311 1420
rect 1315 1416 1316 1420
rect 1310 1415 1316 1416
rect 1670 1419 1676 1420
rect 1670 1415 1671 1419
rect 1675 1415 1676 1419
rect 2103 1417 2104 1421
rect 2108 1420 2109 1421
rect 2116 1420 2239 1422
rect 2108 1419 2118 1420
rect 2111 1418 2118 1419
rect 2215 1419 2221 1420
rect 2103 1416 2107 1417
rect 1670 1414 1676 1415
rect 1982 1415 1988 1416
rect 1982 1411 1983 1415
rect 1987 1411 1988 1415
rect 1982 1410 1988 1411
rect 1990 1415 1997 1416
rect 1990 1411 1991 1415
rect 1996 1411 1997 1415
rect 1990 1410 1997 1411
rect 2094 1415 2100 1416
rect 2094 1411 2095 1415
rect 2099 1411 2100 1415
rect 2106 1415 2107 1416
rect 2111 1415 2112 1418
rect 2106 1414 2112 1415
rect 2206 1415 2212 1416
rect 2094 1410 2100 1411
rect 2206 1411 2207 1415
rect 2211 1411 2212 1415
rect 2215 1415 2216 1419
rect 2220 1415 2221 1419
rect 2238 1419 2239 1420
rect 2243 1419 2244 1423
rect 3006 1423 3012 1424
rect 2238 1418 2244 1419
rect 2343 1419 2349 1420
rect 2215 1414 2221 1415
rect 2334 1415 2340 1416
rect 2206 1410 2212 1411
rect 2334 1411 2335 1415
rect 2339 1411 2340 1415
rect 2343 1415 2344 1419
rect 2348 1418 2349 1419
rect 2398 1419 2404 1420
rect 2398 1418 2399 1419
rect 2348 1416 2399 1418
rect 2348 1415 2349 1416
rect 2343 1414 2349 1415
rect 2398 1415 2399 1416
rect 2403 1415 2404 1419
rect 2486 1419 2493 1420
rect 2398 1414 2404 1415
rect 2478 1415 2484 1416
rect 2334 1410 2340 1411
rect 2478 1411 2479 1415
rect 2483 1411 2484 1415
rect 2486 1415 2487 1419
rect 2492 1415 2493 1419
rect 2647 1419 2653 1420
rect 2486 1414 2493 1415
rect 2638 1415 2644 1416
rect 2478 1410 2484 1411
rect 2638 1411 2639 1415
rect 2643 1411 2644 1415
rect 2647 1415 2648 1419
rect 2652 1418 2653 1419
rect 2662 1419 2668 1420
rect 2662 1418 2663 1419
rect 2652 1416 2663 1418
rect 2652 1415 2653 1416
rect 2647 1414 2653 1415
rect 2662 1415 2663 1416
rect 2667 1415 2668 1419
rect 2862 1419 2868 1420
rect 2862 1418 2863 1419
rect 2839 1416 2863 1418
rect 2662 1414 2668 1415
rect 2814 1415 2820 1416
rect 2638 1410 2644 1411
rect 2814 1411 2815 1415
rect 2819 1411 2820 1415
rect 2814 1410 2820 1411
rect 2822 1415 2829 1416
rect 2822 1411 2823 1415
rect 2828 1414 2829 1415
rect 2839 1414 2841 1416
rect 2862 1415 2863 1416
rect 2867 1415 2868 1419
rect 3006 1419 3007 1423
rect 3011 1422 3012 1423
rect 3118 1423 3124 1424
rect 3118 1422 3119 1423
rect 3011 1420 3119 1422
rect 3011 1419 3013 1420
rect 3006 1418 3008 1419
rect 2862 1414 2868 1415
rect 2998 1415 3004 1416
rect 2828 1412 2841 1414
rect 2828 1411 2829 1412
rect 2822 1410 2829 1411
rect 2998 1411 2999 1415
rect 3003 1411 3004 1415
rect 3007 1415 3008 1418
rect 3012 1415 3013 1419
rect 3118 1419 3119 1420
rect 3123 1422 3124 1423
rect 3123 1420 3171 1422
rect 3123 1419 3124 1420
rect 3118 1418 3124 1419
rect 3166 1419 3173 1420
rect 3007 1414 3013 1415
rect 3158 1415 3164 1416
rect 2998 1410 3004 1411
rect 3158 1411 3159 1415
rect 3163 1411 3164 1415
rect 3166 1415 3167 1419
rect 3172 1415 3173 1419
rect 3166 1414 3173 1415
rect 3190 1419 3196 1420
rect 3190 1415 3191 1419
rect 3195 1415 3196 1419
rect 3190 1414 3196 1415
rect 3158 1410 3164 1411
rect 374 1396 380 1397
rect 374 1392 375 1396
rect 379 1392 380 1396
rect 374 1391 380 1392
rect 502 1396 508 1397
rect 502 1392 503 1396
rect 507 1392 508 1396
rect 502 1391 508 1392
rect 622 1396 628 1397
rect 622 1392 623 1396
rect 627 1392 628 1396
rect 622 1391 628 1392
rect 742 1396 748 1397
rect 742 1392 743 1396
rect 747 1392 748 1396
rect 742 1391 748 1392
rect 862 1396 868 1397
rect 862 1392 863 1396
rect 867 1392 868 1396
rect 862 1391 868 1392
rect 974 1396 980 1397
rect 974 1392 975 1396
rect 979 1392 980 1396
rect 974 1391 980 1392
rect 1094 1396 1100 1397
rect 1094 1392 1095 1396
rect 1099 1392 1100 1396
rect 1094 1391 1100 1392
rect 1214 1396 1220 1397
rect 1214 1392 1215 1396
rect 1219 1392 1220 1396
rect 1214 1391 1220 1392
rect 110 1389 116 1390
rect 110 1385 111 1389
rect 115 1385 116 1389
rect 110 1384 116 1385
rect 1630 1389 1636 1390
rect 1630 1385 1631 1389
rect 1635 1385 1636 1389
rect 1878 1389 1884 1390
rect 1630 1384 1636 1385
rect 1670 1385 1676 1386
rect 1670 1381 1671 1385
rect 1675 1381 1676 1385
rect 1878 1385 1879 1389
rect 1883 1385 1884 1389
rect 1878 1384 1884 1385
rect 1990 1389 1996 1390
rect 1990 1385 1991 1389
rect 1995 1385 1996 1389
rect 1990 1384 1996 1385
rect 2102 1389 2108 1390
rect 2102 1385 2103 1389
rect 2107 1385 2108 1389
rect 2102 1384 2108 1385
rect 2238 1389 2244 1390
rect 2238 1385 2239 1389
rect 2243 1385 2244 1389
rect 2390 1389 2396 1390
rect 2238 1384 2244 1385
rect 2246 1387 2253 1388
rect 1670 1380 1676 1381
rect 1886 1383 1893 1384
rect 1886 1379 1887 1383
rect 1892 1379 1893 1383
rect 1886 1378 1893 1379
rect 1998 1383 2005 1384
rect 1998 1379 1999 1383
rect 2004 1382 2005 1383
rect 2110 1383 2117 1384
rect 2110 1382 2111 1383
rect 2004 1380 2111 1382
rect 2004 1379 2005 1380
rect 1998 1378 2005 1379
rect 2110 1379 2111 1380
rect 2116 1379 2117 1383
rect 2246 1383 2247 1387
rect 2252 1383 2253 1387
rect 2390 1385 2391 1389
rect 2395 1385 2396 1389
rect 2566 1389 2572 1390
rect 2390 1384 2396 1385
rect 2398 1387 2405 1388
rect 2246 1382 2253 1383
rect 2398 1383 2399 1387
rect 2404 1383 2405 1387
rect 2566 1385 2567 1389
rect 2571 1385 2572 1389
rect 2766 1389 2772 1390
rect 2566 1384 2572 1385
rect 2575 1387 2581 1388
rect 2398 1382 2405 1383
rect 2575 1383 2576 1387
rect 2580 1386 2581 1387
rect 2662 1387 2668 1388
rect 2662 1386 2663 1387
rect 2580 1384 2663 1386
rect 2580 1383 2581 1384
rect 2575 1382 2581 1383
rect 2662 1383 2663 1384
rect 2667 1383 2668 1387
rect 2766 1385 2767 1389
rect 2771 1385 2772 1389
rect 2974 1389 2980 1390
rect 2766 1384 2772 1385
rect 2775 1387 2781 1388
rect 2662 1382 2668 1383
rect 2775 1383 2776 1387
rect 2780 1386 2781 1387
rect 2822 1387 2828 1388
rect 2822 1386 2823 1387
rect 2780 1384 2823 1386
rect 2780 1383 2781 1384
rect 2775 1382 2781 1383
rect 2822 1383 2823 1384
rect 2827 1383 2828 1387
rect 2974 1385 2975 1389
rect 2979 1385 2980 1389
rect 3158 1389 3164 1390
rect 2974 1384 2980 1385
rect 2982 1387 2989 1388
rect 2822 1382 2828 1383
rect 2982 1383 2983 1387
rect 2988 1386 2989 1387
rect 3006 1387 3012 1388
rect 3006 1386 3007 1387
rect 2988 1384 3007 1386
rect 2988 1383 2989 1384
rect 2982 1382 2989 1383
rect 3006 1383 3007 1384
rect 3011 1383 3012 1387
rect 3158 1385 3159 1389
rect 3163 1385 3164 1389
rect 3158 1384 3164 1385
rect 3166 1387 3173 1388
rect 3006 1382 3012 1383
rect 3166 1383 3167 1387
rect 3172 1383 3173 1387
rect 3166 1382 3173 1383
rect 3190 1385 3196 1386
rect 3190 1381 3191 1385
rect 3195 1381 3196 1385
rect 3190 1380 3196 1381
rect 2110 1378 2117 1379
rect 1105 1372 1227 1374
rect 110 1371 116 1372
rect 110 1367 111 1371
rect 115 1367 116 1371
rect 1105 1368 1107 1372
rect 1223 1371 1229 1372
rect 110 1366 116 1367
rect 374 1367 380 1368
rect 374 1363 375 1367
rect 379 1363 380 1367
rect 374 1362 380 1363
rect 382 1367 389 1368
rect 382 1363 383 1367
rect 388 1363 389 1367
rect 382 1362 389 1363
rect 502 1367 508 1368
rect 502 1363 503 1367
rect 507 1363 508 1367
rect 502 1362 508 1363
rect 511 1367 517 1368
rect 511 1363 512 1367
rect 516 1366 517 1367
rect 534 1367 540 1368
rect 534 1366 535 1367
rect 516 1364 535 1366
rect 516 1363 517 1364
rect 511 1362 517 1363
rect 534 1363 535 1364
rect 539 1363 540 1367
rect 534 1362 540 1363
rect 622 1367 628 1368
rect 622 1363 623 1367
rect 627 1363 628 1367
rect 622 1362 628 1363
rect 631 1367 640 1368
rect 631 1363 632 1367
rect 639 1363 640 1367
rect 631 1362 640 1363
rect 742 1367 748 1368
rect 742 1363 743 1367
rect 747 1363 748 1367
rect 742 1362 748 1363
rect 751 1367 757 1368
rect 751 1363 752 1367
rect 756 1366 757 1367
rect 786 1367 792 1368
rect 786 1366 787 1367
rect 756 1364 787 1366
rect 756 1363 757 1364
rect 751 1362 757 1363
rect 786 1363 787 1364
rect 791 1363 792 1367
rect 786 1362 792 1363
rect 862 1367 868 1368
rect 862 1363 863 1367
rect 867 1363 868 1367
rect 862 1362 868 1363
rect 871 1367 877 1368
rect 871 1363 872 1367
rect 876 1366 877 1367
rect 886 1367 892 1368
rect 886 1366 887 1367
rect 876 1364 887 1366
rect 876 1363 877 1364
rect 871 1362 877 1363
rect 886 1363 887 1364
rect 891 1363 892 1367
rect 886 1362 892 1363
rect 974 1367 980 1368
rect 974 1363 975 1367
rect 979 1363 980 1367
rect 974 1362 980 1363
rect 983 1367 989 1368
rect 983 1363 984 1367
rect 988 1366 989 1367
rect 1014 1367 1020 1368
rect 1014 1366 1015 1367
rect 988 1364 1015 1366
rect 988 1363 989 1364
rect 983 1362 989 1363
rect 1014 1363 1015 1364
rect 1019 1363 1020 1367
rect 1014 1362 1020 1363
rect 1094 1367 1100 1368
rect 1094 1363 1095 1367
rect 1099 1363 1100 1367
rect 1094 1362 1100 1363
rect 1102 1367 1109 1368
rect 1102 1363 1103 1367
rect 1108 1363 1109 1367
rect 1102 1362 1109 1363
rect 1214 1367 1220 1368
rect 1214 1363 1215 1367
rect 1219 1363 1220 1367
rect 1223 1367 1224 1371
rect 1228 1367 1229 1371
rect 1223 1366 1229 1367
rect 1630 1371 1636 1372
rect 1630 1367 1631 1371
rect 1635 1367 1636 1371
rect 1630 1366 1636 1367
rect 1670 1367 1676 1368
rect 1214 1362 1220 1363
rect 1670 1363 1671 1367
rect 1675 1363 1676 1367
rect 1670 1362 1676 1363
rect 3190 1367 3196 1368
rect 3190 1363 3191 1367
rect 3195 1363 3196 1367
rect 3190 1362 3196 1363
rect 1878 1360 1884 1361
rect 1878 1356 1879 1360
rect 1883 1356 1884 1360
rect 1878 1355 1884 1356
rect 1990 1360 1996 1361
rect 1990 1356 1991 1360
rect 1995 1356 1996 1360
rect 1990 1355 1996 1356
rect 2102 1360 2108 1361
rect 2102 1356 2103 1360
rect 2107 1356 2108 1360
rect 2102 1355 2108 1356
rect 2238 1360 2244 1361
rect 2238 1356 2239 1360
rect 2243 1356 2244 1360
rect 2238 1355 2244 1356
rect 2390 1360 2396 1361
rect 2390 1356 2391 1360
rect 2395 1356 2396 1360
rect 2390 1355 2396 1356
rect 2566 1360 2572 1361
rect 2566 1356 2567 1360
rect 2571 1356 2572 1360
rect 2566 1355 2572 1356
rect 2766 1360 2772 1361
rect 2766 1356 2767 1360
rect 2771 1356 2772 1360
rect 2766 1355 2772 1356
rect 2974 1360 2980 1361
rect 2974 1356 2975 1360
rect 2979 1356 2980 1360
rect 2974 1355 2980 1356
rect 3158 1360 3164 1361
rect 3158 1356 3159 1360
rect 3163 1356 3164 1360
rect 3158 1355 3164 1356
rect 270 1349 276 1350
rect 110 1345 116 1346
rect 110 1341 111 1345
rect 115 1341 116 1345
rect 270 1345 271 1349
rect 275 1345 276 1349
rect 270 1344 276 1345
rect 398 1349 404 1350
rect 398 1345 399 1349
rect 403 1345 404 1349
rect 398 1344 404 1345
rect 526 1349 532 1350
rect 526 1345 527 1349
rect 531 1345 532 1349
rect 526 1344 532 1345
rect 646 1349 652 1350
rect 646 1345 647 1349
rect 651 1345 652 1349
rect 646 1344 652 1345
rect 766 1349 772 1350
rect 766 1345 767 1349
rect 771 1345 772 1349
rect 766 1344 772 1345
rect 878 1349 884 1350
rect 878 1345 879 1349
rect 883 1345 884 1349
rect 878 1344 884 1345
rect 990 1349 996 1350
rect 990 1345 991 1349
rect 995 1345 996 1349
rect 990 1344 996 1345
rect 1110 1349 1116 1350
rect 1110 1345 1111 1349
rect 1115 1345 1116 1349
rect 1110 1344 1116 1345
rect 1630 1345 1636 1346
rect 110 1340 116 1341
rect 279 1343 285 1344
rect 279 1339 280 1343
rect 284 1342 285 1343
rect 310 1343 316 1344
rect 310 1342 311 1343
rect 284 1340 311 1342
rect 284 1339 285 1340
rect 279 1338 285 1339
rect 310 1339 311 1340
rect 315 1342 316 1343
rect 382 1343 388 1344
rect 382 1342 383 1343
rect 315 1340 383 1342
rect 315 1339 316 1340
rect 310 1338 316 1339
rect 382 1339 383 1340
rect 387 1342 388 1343
rect 407 1343 413 1344
rect 407 1342 408 1343
rect 387 1340 408 1342
rect 387 1339 388 1340
rect 382 1338 388 1339
rect 407 1339 408 1340
rect 412 1339 413 1343
rect 407 1338 413 1339
rect 534 1343 541 1344
rect 534 1339 535 1343
rect 540 1342 541 1343
rect 634 1343 640 1344
rect 634 1342 635 1343
rect 540 1340 635 1342
rect 540 1339 541 1340
rect 534 1338 541 1339
rect 634 1339 635 1340
rect 639 1342 640 1343
rect 655 1343 661 1344
rect 655 1342 656 1343
rect 639 1340 656 1342
rect 639 1339 640 1340
rect 634 1338 640 1339
rect 655 1339 656 1340
rect 660 1342 661 1343
rect 775 1343 781 1344
rect 775 1342 776 1343
rect 660 1340 776 1342
rect 660 1339 661 1340
rect 655 1338 661 1339
rect 775 1339 776 1340
rect 780 1342 781 1343
rect 786 1343 792 1344
rect 786 1342 787 1343
rect 780 1340 787 1342
rect 780 1339 781 1340
rect 775 1338 781 1339
rect 786 1339 787 1340
rect 791 1339 792 1343
rect 786 1338 792 1339
rect 887 1343 893 1344
rect 887 1339 888 1343
rect 892 1339 893 1343
rect 887 1338 893 1339
rect 999 1343 1005 1344
rect 999 1339 1000 1343
rect 1004 1342 1005 1343
rect 1014 1343 1020 1344
rect 1014 1342 1015 1343
rect 1004 1340 1015 1342
rect 1004 1339 1005 1340
rect 999 1338 1005 1339
rect 1014 1339 1015 1340
rect 1019 1342 1020 1343
rect 1102 1343 1108 1344
rect 1102 1342 1103 1343
rect 1019 1340 1103 1342
rect 1019 1339 1020 1340
rect 1014 1338 1020 1339
rect 1102 1339 1103 1340
rect 1107 1342 1108 1343
rect 1119 1343 1125 1344
rect 1119 1342 1120 1343
rect 1107 1340 1120 1342
rect 1107 1339 1108 1340
rect 1102 1338 1108 1339
rect 1119 1339 1120 1340
rect 1124 1339 1125 1343
rect 1630 1341 1631 1345
rect 1635 1341 1636 1345
rect 1630 1340 1636 1341
rect 1119 1338 1125 1339
rect 1774 1336 1780 1337
rect 1774 1332 1775 1336
rect 1779 1332 1780 1336
rect 1774 1331 1780 1332
rect 1886 1336 1892 1337
rect 1886 1332 1887 1336
rect 1891 1332 1892 1336
rect 1886 1331 1892 1332
rect 1990 1336 1996 1337
rect 1990 1332 1991 1336
rect 1995 1332 1996 1336
rect 1990 1331 1996 1332
rect 2094 1336 2100 1337
rect 2094 1332 2095 1336
rect 2099 1332 2100 1336
rect 2094 1331 2100 1332
rect 2198 1336 2204 1337
rect 2198 1332 2199 1336
rect 2203 1332 2204 1336
rect 2198 1331 2204 1332
rect 2302 1336 2308 1337
rect 2302 1332 2303 1336
rect 2307 1332 2308 1336
rect 2302 1331 2308 1332
rect 2406 1336 2412 1337
rect 2406 1332 2407 1336
rect 2411 1332 2412 1336
rect 2406 1331 2412 1332
rect 2510 1336 2516 1337
rect 2510 1332 2511 1336
rect 2515 1332 2516 1336
rect 2510 1331 2516 1332
rect 1670 1329 1676 1330
rect 110 1327 116 1328
rect 110 1323 111 1327
rect 115 1323 116 1327
rect 110 1322 116 1323
rect 1630 1327 1636 1328
rect 1630 1323 1631 1327
rect 1635 1323 1636 1327
rect 1670 1325 1671 1329
rect 1675 1325 1676 1329
rect 1670 1324 1676 1325
rect 3190 1329 3196 1330
rect 3190 1325 3191 1329
rect 3195 1325 3196 1329
rect 3190 1324 3196 1325
rect 1630 1322 1636 1323
rect 270 1320 276 1321
rect 270 1316 271 1320
rect 275 1316 276 1320
rect 270 1315 276 1316
rect 398 1320 404 1321
rect 398 1316 399 1320
rect 403 1316 404 1320
rect 398 1315 404 1316
rect 526 1320 532 1321
rect 526 1316 527 1320
rect 531 1316 532 1320
rect 526 1315 532 1316
rect 646 1320 652 1321
rect 646 1316 647 1320
rect 651 1316 652 1320
rect 646 1315 652 1316
rect 766 1320 772 1321
rect 766 1316 767 1320
rect 771 1316 772 1320
rect 766 1315 772 1316
rect 878 1320 884 1321
rect 878 1316 879 1320
rect 883 1316 884 1320
rect 878 1315 884 1316
rect 990 1320 996 1321
rect 990 1316 991 1320
rect 995 1316 996 1320
rect 990 1315 996 1316
rect 1110 1320 1116 1321
rect 1110 1316 1111 1320
rect 1115 1316 1116 1320
rect 1110 1315 1116 1316
rect 1894 1315 1900 1316
rect 1894 1314 1895 1315
rect 1880 1312 1895 1314
rect 1670 1311 1676 1312
rect 1670 1307 1671 1311
rect 1675 1307 1676 1311
rect 1670 1306 1676 1307
rect 1774 1307 1780 1308
rect 1774 1303 1775 1307
rect 1779 1303 1780 1307
rect 1774 1302 1780 1303
rect 1782 1307 1789 1308
rect 1782 1303 1783 1307
rect 1788 1306 1789 1307
rect 1880 1306 1882 1312
rect 1894 1311 1895 1312
rect 1899 1312 1900 1315
rect 1998 1315 2004 1316
rect 1998 1314 1999 1315
rect 1944 1312 1999 1314
rect 1899 1311 1901 1312
rect 1894 1310 1896 1311
rect 1788 1304 1882 1306
rect 1886 1307 1892 1308
rect 1788 1303 1789 1304
rect 1782 1302 1789 1303
rect 1886 1303 1887 1307
rect 1891 1303 1892 1307
rect 1895 1307 1896 1310
rect 1900 1310 1901 1311
rect 1942 1311 1948 1312
rect 1942 1310 1943 1311
rect 1900 1308 1943 1310
rect 1900 1307 1901 1308
rect 1895 1306 1901 1307
rect 1942 1307 1943 1308
rect 1947 1307 1948 1311
rect 1998 1311 1999 1312
rect 2003 1314 2004 1315
rect 2102 1315 2108 1316
rect 2102 1314 2103 1315
rect 2003 1312 2103 1314
rect 2107 1314 2108 1315
rect 2398 1315 2404 1316
rect 2107 1313 2109 1314
rect 2003 1311 2005 1312
rect 1998 1310 2000 1311
rect 1942 1306 1948 1307
rect 1990 1307 1996 1308
rect 1886 1302 1892 1303
rect 1990 1303 1991 1307
rect 1995 1303 1996 1307
rect 1999 1307 2000 1310
rect 2004 1307 2005 1311
rect 2102 1311 2103 1312
rect 2102 1310 2104 1311
rect 2103 1309 2104 1310
rect 2108 1309 2109 1313
rect 2103 1308 2109 1309
rect 2239 1312 2314 1314
rect 1999 1306 2005 1307
rect 2094 1307 2100 1308
rect 1990 1302 1996 1303
rect 2094 1303 2095 1307
rect 2099 1303 2100 1307
rect 2094 1302 2100 1303
rect 2198 1307 2204 1308
rect 2198 1303 2199 1307
rect 2203 1303 2204 1307
rect 2198 1302 2204 1303
rect 2207 1307 2213 1308
rect 2207 1303 2208 1307
rect 2212 1306 2213 1307
rect 2239 1306 2241 1312
rect 2312 1308 2314 1312
rect 2398 1311 2399 1315
rect 2403 1314 2404 1315
rect 2502 1315 2508 1316
rect 2502 1314 2503 1315
rect 2403 1312 2503 1314
rect 2403 1311 2404 1312
rect 2398 1310 2404 1311
rect 2415 1311 2421 1312
rect 2212 1304 2241 1306
rect 2302 1307 2308 1308
rect 2212 1303 2213 1304
rect 2207 1302 2213 1303
rect 2302 1303 2303 1307
rect 2307 1303 2308 1307
rect 2302 1302 2308 1303
rect 2311 1307 2317 1308
rect 2311 1303 2312 1307
rect 2316 1306 2317 1307
rect 2351 1307 2357 1308
rect 2351 1306 2352 1307
rect 2316 1304 2352 1306
rect 2316 1303 2317 1304
rect 2311 1302 2317 1303
rect 2351 1303 2352 1304
rect 2356 1303 2357 1307
rect 2351 1302 2357 1303
rect 2406 1307 2412 1308
rect 2406 1303 2407 1307
rect 2411 1303 2412 1307
rect 2415 1307 2416 1311
rect 2420 1307 2421 1311
rect 2502 1311 2503 1312
rect 2507 1314 2508 1315
rect 2507 1312 2522 1314
rect 2507 1311 2508 1312
rect 2502 1310 2508 1311
rect 2519 1311 2525 1312
rect 2415 1306 2421 1307
rect 2510 1307 2516 1308
rect 2406 1302 2412 1303
rect 2510 1303 2511 1307
rect 2515 1303 2516 1307
rect 2519 1307 2520 1311
rect 2524 1307 2525 1311
rect 2519 1306 2525 1307
rect 3190 1311 3196 1312
rect 3190 1307 3191 1311
rect 3195 1307 3196 1311
rect 3190 1306 3196 1307
rect 2510 1302 2516 1303
rect 2110 1299 2116 1300
rect 174 1296 180 1297
rect 174 1292 175 1296
rect 179 1292 180 1296
rect 174 1291 180 1292
rect 302 1296 308 1297
rect 302 1292 303 1296
rect 307 1292 308 1296
rect 302 1291 308 1292
rect 422 1296 428 1297
rect 422 1292 423 1296
rect 427 1292 428 1296
rect 422 1291 428 1292
rect 542 1296 548 1297
rect 542 1292 543 1296
rect 547 1292 548 1296
rect 542 1291 548 1292
rect 662 1296 668 1297
rect 662 1292 663 1296
rect 667 1292 668 1296
rect 662 1291 668 1292
rect 774 1296 780 1297
rect 774 1292 775 1296
rect 779 1292 780 1296
rect 774 1291 780 1292
rect 886 1296 892 1297
rect 886 1292 887 1296
rect 891 1292 892 1296
rect 886 1291 892 1292
rect 1006 1296 1012 1297
rect 1006 1292 1007 1296
rect 1011 1292 1012 1296
rect 2110 1295 2111 1299
rect 2115 1298 2116 1299
rect 2209 1298 2211 1302
rect 2312 1298 2314 1302
rect 2115 1296 2211 1298
rect 2304 1296 2314 1298
rect 2115 1295 2116 1296
rect 2110 1294 2116 1295
rect 1006 1291 1012 1292
rect 2304 1290 2306 1296
rect 110 1289 116 1290
rect 110 1285 111 1289
rect 115 1285 116 1289
rect 110 1284 116 1285
rect 1630 1289 1636 1290
rect 1630 1285 1631 1289
rect 1635 1285 1636 1289
rect 1694 1289 1700 1290
rect 1630 1284 1636 1285
rect 1670 1285 1676 1286
rect 1670 1281 1671 1285
rect 1675 1281 1676 1285
rect 1694 1285 1695 1289
rect 1699 1285 1700 1289
rect 1694 1284 1700 1285
rect 1790 1289 1796 1290
rect 1790 1285 1791 1289
rect 1795 1285 1796 1289
rect 1790 1284 1796 1285
rect 1934 1289 1940 1290
rect 1934 1285 1935 1289
rect 1939 1285 1940 1289
rect 2102 1289 2108 1290
rect 1934 1284 1940 1285
rect 1942 1287 1949 1288
rect 1670 1280 1676 1281
rect 1702 1283 1709 1284
rect 1702 1279 1703 1283
rect 1708 1282 1709 1283
rect 1782 1283 1788 1284
rect 1782 1282 1783 1283
rect 1708 1280 1783 1282
rect 1708 1279 1709 1280
rect 1702 1278 1709 1279
rect 1782 1279 1783 1280
rect 1787 1282 1788 1283
rect 1799 1283 1805 1284
rect 1799 1282 1800 1283
rect 1787 1280 1800 1282
rect 1787 1279 1788 1280
rect 1782 1278 1788 1279
rect 1799 1279 1800 1280
rect 1804 1279 1805 1283
rect 1942 1283 1943 1287
rect 1948 1283 1949 1287
rect 2102 1285 2103 1289
rect 2107 1285 2108 1289
rect 2294 1289 2300 1290
rect 2102 1284 2108 1285
rect 2110 1287 2117 1288
rect 1942 1282 1949 1283
rect 2110 1283 2111 1287
rect 2116 1283 2117 1287
rect 2294 1285 2295 1289
rect 2299 1285 2300 1289
rect 2294 1284 2300 1285
rect 2303 1289 2309 1290
rect 2303 1285 2304 1289
rect 2308 1285 2309 1289
rect 2303 1284 2309 1285
rect 2494 1289 2500 1290
rect 2494 1285 2495 1289
rect 2499 1285 2500 1289
rect 2710 1289 2716 1290
rect 2494 1284 2500 1285
rect 2502 1287 2509 1288
rect 2110 1282 2117 1283
rect 2502 1283 2503 1287
rect 2508 1283 2509 1287
rect 2710 1285 2711 1289
rect 2715 1285 2716 1289
rect 2710 1284 2716 1285
rect 2934 1289 2940 1290
rect 2934 1285 2935 1289
rect 2939 1285 2940 1289
rect 3158 1289 3164 1290
rect 2934 1284 2940 1285
rect 2943 1287 2949 1288
rect 2502 1282 2509 1283
rect 2718 1283 2725 1284
rect 1799 1278 1805 1279
rect 2718 1279 2719 1283
rect 2724 1279 2725 1283
rect 2943 1283 2944 1287
rect 2948 1286 2949 1287
rect 2982 1287 2988 1288
rect 2982 1286 2983 1287
rect 2948 1284 2983 1286
rect 2948 1283 2949 1284
rect 2943 1282 2949 1283
rect 2982 1283 2983 1284
rect 2987 1283 2988 1287
rect 3158 1285 3159 1289
rect 3163 1285 3164 1289
rect 3158 1284 3164 1285
rect 3166 1287 3173 1288
rect 2982 1282 2988 1283
rect 3166 1283 3167 1287
rect 3172 1283 3173 1287
rect 3166 1282 3173 1283
rect 3190 1285 3196 1286
rect 3190 1281 3191 1285
rect 3195 1281 3196 1285
rect 3190 1280 3196 1281
rect 2718 1278 2725 1279
rect 110 1271 116 1272
rect 110 1267 111 1271
rect 115 1267 116 1271
rect 310 1271 317 1272
rect 110 1266 116 1267
rect 174 1267 180 1268
rect 174 1263 175 1267
rect 179 1263 180 1267
rect 174 1262 180 1263
rect 183 1267 192 1268
rect 183 1263 184 1267
rect 191 1263 192 1267
rect 183 1262 192 1263
rect 302 1267 308 1268
rect 302 1263 303 1267
rect 307 1263 308 1267
rect 310 1267 311 1271
rect 316 1267 317 1271
rect 550 1271 557 1272
rect 310 1266 317 1267
rect 422 1267 428 1268
rect 302 1262 308 1263
rect 422 1263 423 1267
rect 427 1263 428 1267
rect 422 1262 428 1263
rect 430 1267 437 1268
rect 430 1263 431 1267
rect 436 1263 437 1267
rect 430 1262 437 1263
rect 542 1267 548 1268
rect 542 1263 543 1267
rect 547 1263 548 1267
rect 550 1267 551 1271
rect 556 1270 557 1271
rect 634 1271 640 1272
rect 634 1270 635 1271
rect 556 1268 635 1270
rect 556 1267 557 1268
rect 550 1266 557 1267
rect 634 1267 635 1268
rect 639 1267 640 1271
rect 1630 1271 1636 1272
rect 634 1266 640 1267
rect 662 1267 668 1268
rect 542 1262 548 1263
rect 662 1263 663 1267
rect 667 1263 668 1267
rect 662 1262 668 1263
rect 670 1267 677 1268
rect 670 1263 671 1267
rect 676 1263 677 1267
rect 670 1262 677 1263
rect 774 1267 780 1268
rect 774 1263 775 1267
rect 779 1263 780 1267
rect 774 1262 780 1263
rect 783 1267 792 1268
rect 783 1263 784 1267
rect 791 1263 792 1267
rect 783 1262 792 1263
rect 886 1267 892 1268
rect 886 1263 887 1267
rect 891 1263 892 1267
rect 886 1262 892 1263
rect 894 1267 901 1268
rect 894 1263 895 1267
rect 900 1263 901 1267
rect 894 1262 901 1263
rect 1006 1267 1012 1268
rect 1006 1263 1007 1267
rect 1011 1263 1012 1267
rect 1006 1262 1012 1263
rect 1015 1267 1021 1268
rect 1015 1263 1016 1267
rect 1020 1263 1021 1267
rect 1630 1267 1631 1271
rect 1635 1267 1636 1271
rect 1630 1266 1636 1267
rect 1670 1267 1676 1268
rect 1015 1262 1021 1263
rect 1670 1263 1671 1267
rect 1675 1263 1676 1267
rect 1670 1262 1676 1263
rect 3190 1267 3196 1268
rect 3190 1263 3191 1267
rect 3195 1263 3196 1267
rect 3190 1262 3196 1263
rect 866 1259 872 1260
rect 866 1255 867 1259
rect 871 1258 872 1259
rect 897 1258 899 1262
rect 871 1256 899 1258
rect 1694 1260 1700 1261
rect 1694 1256 1695 1260
rect 1699 1256 1700 1260
rect 871 1255 872 1256
rect 1694 1255 1700 1256
rect 1790 1260 1796 1261
rect 1790 1256 1791 1260
rect 1795 1256 1796 1260
rect 1790 1255 1796 1256
rect 1934 1260 1940 1261
rect 1934 1256 1935 1260
rect 1939 1256 1940 1260
rect 1934 1255 1940 1256
rect 2102 1260 2108 1261
rect 2102 1256 2103 1260
rect 2107 1256 2108 1260
rect 2102 1255 2108 1256
rect 2294 1260 2300 1261
rect 2294 1256 2295 1260
rect 2299 1256 2300 1260
rect 2294 1255 2300 1256
rect 2494 1260 2500 1261
rect 2494 1256 2495 1260
rect 2499 1256 2500 1260
rect 2494 1255 2500 1256
rect 2710 1260 2716 1261
rect 2710 1256 2711 1260
rect 2715 1256 2716 1260
rect 2710 1255 2716 1256
rect 2934 1260 2940 1261
rect 2934 1256 2935 1260
rect 2939 1256 2940 1260
rect 2934 1255 2940 1256
rect 3158 1260 3164 1261
rect 3158 1256 3159 1260
rect 3163 1256 3164 1260
rect 3158 1255 3164 1256
rect 866 1254 872 1255
rect 134 1245 140 1246
rect 110 1241 116 1242
rect 110 1237 111 1241
rect 115 1237 116 1241
rect 134 1241 135 1245
rect 139 1241 140 1245
rect 134 1240 140 1241
rect 230 1245 236 1246
rect 230 1241 231 1245
rect 235 1241 236 1245
rect 230 1240 236 1241
rect 358 1245 364 1246
rect 358 1241 359 1245
rect 363 1241 364 1245
rect 358 1240 364 1241
rect 502 1245 508 1246
rect 502 1241 503 1245
rect 507 1241 508 1245
rect 662 1245 668 1246
rect 502 1240 508 1241
rect 511 1243 517 1244
rect 110 1236 116 1237
rect 143 1239 149 1240
rect 143 1235 144 1239
rect 148 1238 149 1239
rect 186 1239 192 1240
rect 186 1238 187 1239
rect 148 1236 187 1238
rect 148 1235 149 1236
rect 143 1234 149 1235
rect 186 1235 187 1236
rect 191 1238 192 1239
rect 239 1239 245 1240
rect 239 1238 240 1239
rect 191 1236 240 1238
rect 191 1235 192 1236
rect 186 1234 192 1235
rect 239 1235 240 1236
rect 244 1238 245 1239
rect 258 1239 264 1240
rect 258 1238 259 1239
rect 244 1236 259 1238
rect 244 1235 245 1236
rect 239 1234 245 1235
rect 258 1235 259 1236
rect 263 1238 264 1239
rect 310 1239 316 1240
rect 310 1238 311 1239
rect 263 1236 311 1238
rect 263 1235 264 1236
rect 258 1234 264 1235
rect 310 1235 311 1236
rect 315 1238 316 1239
rect 367 1239 373 1240
rect 367 1238 368 1239
rect 315 1236 368 1238
rect 315 1235 316 1236
rect 310 1234 316 1235
rect 367 1235 368 1236
rect 372 1238 373 1239
rect 430 1239 436 1240
rect 430 1238 431 1239
rect 372 1236 431 1238
rect 372 1235 373 1236
rect 367 1234 373 1235
rect 430 1235 431 1236
rect 435 1238 436 1239
rect 511 1239 512 1243
rect 516 1242 517 1243
rect 550 1243 556 1244
rect 550 1242 551 1243
rect 516 1240 551 1242
rect 516 1239 517 1240
rect 511 1238 517 1239
rect 550 1239 551 1240
rect 555 1239 556 1243
rect 662 1241 663 1245
rect 667 1241 668 1245
rect 662 1240 668 1241
rect 830 1245 836 1246
rect 830 1241 831 1245
rect 835 1241 836 1245
rect 830 1240 836 1241
rect 1014 1245 1020 1246
rect 1014 1241 1015 1245
rect 1019 1241 1020 1245
rect 1014 1240 1020 1241
rect 1206 1245 1212 1246
rect 1206 1241 1207 1245
rect 1211 1241 1212 1245
rect 1206 1240 1212 1241
rect 1406 1245 1412 1246
rect 1406 1241 1407 1245
rect 1411 1241 1412 1245
rect 1406 1240 1412 1241
rect 1598 1245 1604 1246
rect 1598 1241 1599 1245
rect 1603 1241 1604 1245
rect 1598 1240 1604 1241
rect 1630 1241 1636 1242
rect 550 1238 556 1239
rect 670 1239 677 1240
rect 435 1236 514 1238
rect 435 1235 436 1236
rect 430 1234 436 1235
rect 670 1235 671 1239
rect 676 1235 677 1239
rect 670 1234 677 1235
rect 786 1239 792 1240
rect 786 1235 787 1239
rect 791 1238 792 1239
rect 839 1239 845 1240
rect 839 1238 840 1239
rect 791 1236 840 1238
rect 791 1235 792 1236
rect 786 1234 792 1235
rect 839 1235 840 1236
rect 844 1238 845 1239
rect 866 1239 872 1240
rect 866 1238 867 1239
rect 844 1236 867 1238
rect 844 1235 845 1236
rect 839 1234 845 1235
rect 866 1235 867 1236
rect 871 1235 872 1239
rect 866 1234 872 1235
rect 1006 1239 1012 1240
rect 1006 1235 1007 1239
rect 1011 1238 1012 1239
rect 1022 1239 1029 1240
rect 1022 1238 1023 1239
rect 1011 1236 1023 1238
rect 1011 1235 1012 1236
rect 1006 1234 1012 1235
rect 1022 1235 1023 1236
rect 1028 1235 1029 1239
rect 1022 1234 1029 1235
rect 1215 1239 1221 1240
rect 1215 1235 1216 1239
rect 1220 1238 1221 1239
rect 1230 1239 1236 1240
rect 1230 1238 1231 1239
rect 1220 1236 1231 1238
rect 1220 1235 1221 1236
rect 1215 1234 1221 1235
rect 1230 1235 1231 1236
rect 1235 1235 1236 1239
rect 1230 1234 1236 1235
rect 1415 1239 1421 1240
rect 1415 1235 1416 1239
rect 1420 1238 1421 1239
rect 1454 1239 1460 1240
rect 1454 1238 1455 1239
rect 1420 1236 1455 1238
rect 1420 1235 1421 1236
rect 1415 1234 1421 1235
rect 1454 1235 1455 1236
rect 1459 1235 1460 1239
rect 1454 1234 1460 1235
rect 1606 1239 1613 1240
rect 1606 1235 1607 1239
rect 1612 1235 1613 1239
rect 1630 1237 1631 1241
rect 1635 1237 1636 1241
rect 1630 1236 1636 1237
rect 1606 1234 1613 1235
rect 1694 1232 1700 1233
rect 1694 1228 1695 1232
rect 1699 1228 1700 1232
rect 1694 1227 1700 1228
rect 1982 1232 1988 1233
rect 1982 1228 1983 1232
rect 1987 1228 1988 1232
rect 1982 1227 1988 1228
rect 2254 1232 2260 1233
rect 2254 1228 2255 1232
rect 2259 1228 2260 1232
rect 2254 1227 2260 1228
rect 2494 1232 2500 1233
rect 2494 1228 2495 1232
rect 2499 1228 2500 1232
rect 2494 1227 2500 1228
rect 2710 1232 2716 1233
rect 2710 1228 2711 1232
rect 2715 1228 2716 1232
rect 2710 1227 2716 1228
rect 2918 1232 2924 1233
rect 2918 1228 2919 1232
rect 2923 1228 2924 1232
rect 2918 1227 2924 1228
rect 3134 1232 3140 1233
rect 3134 1228 3135 1232
rect 3139 1228 3140 1232
rect 3134 1227 3140 1228
rect 1670 1225 1676 1226
rect 110 1223 116 1224
rect 110 1219 111 1223
rect 115 1219 116 1223
rect 110 1218 116 1219
rect 1630 1223 1636 1224
rect 1630 1219 1631 1223
rect 1635 1219 1636 1223
rect 1670 1221 1671 1225
rect 1675 1221 1676 1225
rect 1670 1220 1676 1221
rect 3190 1225 3196 1226
rect 3190 1221 3191 1225
rect 3195 1221 3196 1225
rect 3190 1220 3196 1221
rect 1630 1218 1636 1219
rect 134 1216 140 1217
rect 134 1212 135 1216
rect 139 1212 140 1216
rect 134 1211 140 1212
rect 230 1216 236 1217
rect 230 1212 231 1216
rect 235 1212 236 1216
rect 230 1211 236 1212
rect 358 1216 364 1217
rect 358 1212 359 1216
rect 363 1212 364 1216
rect 358 1211 364 1212
rect 502 1216 508 1217
rect 502 1212 503 1216
rect 507 1212 508 1216
rect 502 1211 508 1212
rect 662 1216 668 1217
rect 662 1212 663 1216
rect 667 1212 668 1216
rect 662 1211 668 1212
rect 830 1216 836 1217
rect 830 1212 831 1216
rect 835 1212 836 1216
rect 830 1211 836 1212
rect 1014 1216 1020 1217
rect 1014 1212 1015 1216
rect 1019 1212 1020 1216
rect 1014 1211 1020 1212
rect 1206 1216 1212 1217
rect 1206 1212 1207 1216
rect 1211 1212 1212 1216
rect 1206 1211 1212 1212
rect 1406 1216 1412 1217
rect 1406 1212 1407 1216
rect 1411 1212 1412 1216
rect 1406 1211 1412 1212
rect 1598 1216 1604 1217
rect 1598 1212 1599 1216
rect 1603 1212 1604 1216
rect 1598 1211 1604 1212
rect 1606 1215 1612 1216
rect 1606 1211 1607 1215
rect 1611 1214 1612 1215
rect 1702 1215 1708 1216
rect 1702 1214 1703 1215
rect 1611 1212 1703 1214
rect 1611 1211 1612 1212
rect 1606 1210 1612 1211
rect 1702 1211 1703 1212
rect 1707 1211 1708 1215
rect 1702 1210 1708 1211
rect 1942 1211 1948 1212
rect 1705 1208 1707 1210
rect 1670 1207 1676 1208
rect 1670 1203 1671 1207
rect 1675 1203 1676 1207
rect 1703 1207 1709 1208
rect 1670 1202 1676 1203
rect 1694 1203 1700 1204
rect 1694 1199 1695 1203
rect 1699 1199 1700 1203
rect 1703 1203 1704 1207
rect 1708 1203 1709 1207
rect 1942 1207 1943 1211
rect 1947 1210 1948 1211
rect 1947 1208 1994 1210
rect 1947 1207 1948 1208
rect 1942 1206 1948 1207
rect 1991 1207 1997 1208
rect 1703 1202 1709 1203
rect 1982 1203 1988 1204
rect 1694 1198 1700 1199
rect 1982 1199 1983 1203
rect 1987 1199 1988 1203
rect 1991 1203 1992 1207
rect 1996 1203 1997 1207
rect 3142 1207 3149 1208
rect 1991 1202 1997 1203
rect 2254 1203 2260 1204
rect 1982 1198 1988 1199
rect 2254 1199 2255 1203
rect 2259 1199 2260 1203
rect 2254 1198 2260 1199
rect 2263 1203 2269 1204
rect 2263 1199 2264 1203
rect 2268 1202 2269 1203
rect 2351 1203 2357 1204
rect 2351 1202 2352 1203
rect 2268 1200 2352 1202
rect 2268 1199 2269 1200
rect 2263 1198 2269 1199
rect 2351 1199 2352 1200
rect 2356 1199 2357 1203
rect 2351 1198 2357 1199
rect 2494 1203 2500 1204
rect 2494 1199 2495 1203
rect 2499 1199 2500 1203
rect 2494 1198 2500 1199
rect 2503 1203 2512 1204
rect 2503 1199 2504 1203
rect 2511 1199 2512 1203
rect 2503 1198 2512 1199
rect 2710 1203 2716 1204
rect 2710 1199 2711 1203
rect 2715 1199 2716 1203
rect 2710 1198 2716 1199
rect 2718 1203 2725 1204
rect 2718 1199 2719 1203
rect 2724 1202 2725 1203
rect 2854 1203 2860 1204
rect 2854 1202 2855 1203
rect 2724 1200 2855 1202
rect 2724 1199 2725 1200
rect 2718 1198 2725 1199
rect 2854 1199 2855 1200
rect 2859 1199 2860 1203
rect 2854 1198 2860 1199
rect 2918 1203 2924 1204
rect 2918 1199 2919 1203
rect 2923 1199 2924 1203
rect 2918 1198 2924 1199
rect 2927 1203 2933 1204
rect 2927 1199 2928 1203
rect 2932 1202 2933 1203
rect 3006 1203 3012 1204
rect 3006 1202 3007 1203
rect 2932 1200 3007 1202
rect 2932 1199 2933 1200
rect 2927 1198 2933 1199
rect 3006 1199 3007 1200
rect 3011 1199 3012 1203
rect 3006 1198 3012 1199
rect 3134 1203 3140 1204
rect 3134 1199 3135 1203
rect 3139 1199 3140 1203
rect 3142 1203 3143 1207
rect 3148 1206 3149 1207
rect 3166 1207 3172 1208
rect 3166 1206 3167 1207
rect 3148 1204 3167 1206
rect 3148 1203 3149 1204
rect 3142 1202 3149 1203
rect 3166 1203 3167 1204
rect 3171 1203 3172 1207
rect 3166 1202 3172 1203
rect 3190 1207 3196 1208
rect 3190 1203 3191 1207
rect 3195 1203 3196 1207
rect 3190 1202 3196 1203
rect 3134 1198 3140 1199
rect 726 1196 732 1197
rect 726 1192 727 1196
rect 731 1192 732 1196
rect 726 1191 732 1192
rect 854 1196 860 1197
rect 854 1192 855 1196
rect 859 1192 860 1196
rect 854 1191 860 1192
rect 982 1196 988 1197
rect 982 1192 983 1196
rect 987 1192 988 1196
rect 982 1191 988 1192
rect 1102 1196 1108 1197
rect 1102 1192 1103 1196
rect 1107 1192 1108 1196
rect 1102 1191 1108 1192
rect 1222 1196 1228 1197
rect 1222 1192 1223 1196
rect 1227 1192 1228 1196
rect 1222 1191 1228 1192
rect 1334 1196 1340 1197
rect 1334 1192 1335 1196
rect 1339 1192 1340 1196
rect 1334 1191 1340 1192
rect 1446 1196 1452 1197
rect 1446 1192 1447 1196
rect 1451 1192 1452 1196
rect 1446 1191 1452 1192
rect 1566 1196 1572 1197
rect 1566 1192 1567 1196
rect 1571 1192 1572 1196
rect 1566 1191 1572 1192
rect 2182 1195 2188 1196
rect 2182 1191 2183 1195
rect 2187 1194 2188 1195
rect 2264 1194 2266 1198
rect 2187 1192 2266 1194
rect 2187 1191 2188 1192
rect 2182 1190 2188 1191
rect 110 1189 116 1190
rect 110 1185 111 1189
rect 115 1185 116 1189
rect 110 1184 116 1185
rect 1630 1189 1636 1190
rect 1630 1185 1631 1189
rect 1635 1185 1636 1189
rect 2246 1189 2252 1190
rect 1630 1184 1636 1185
rect 1670 1185 1676 1186
rect 1670 1181 1671 1185
rect 1675 1181 1676 1185
rect 2246 1185 2247 1189
rect 2251 1185 2252 1189
rect 2246 1184 2252 1185
rect 2255 1187 2261 1188
rect 2255 1183 2256 1187
rect 2260 1186 2261 1187
rect 2264 1186 2266 1192
rect 2260 1184 2266 1186
rect 2398 1189 2404 1190
rect 2398 1185 2399 1189
rect 2403 1185 2404 1189
rect 2398 1184 2404 1185
rect 2550 1189 2556 1190
rect 2550 1185 2551 1189
rect 2555 1185 2556 1189
rect 2550 1184 2556 1185
rect 2694 1189 2700 1190
rect 2694 1185 2695 1189
rect 2699 1185 2700 1189
rect 2694 1184 2700 1185
rect 2702 1187 2709 1188
rect 2260 1183 2261 1184
rect 2255 1182 2261 1183
rect 2351 1183 2357 1184
rect 1670 1180 1676 1181
rect 2351 1179 2352 1183
rect 2356 1182 2357 1183
rect 2407 1183 2413 1184
rect 2407 1182 2408 1183
rect 2356 1180 2408 1182
rect 2356 1179 2357 1180
rect 2351 1178 2357 1179
rect 2407 1179 2408 1180
rect 2412 1182 2413 1183
rect 2506 1183 2512 1184
rect 2506 1182 2507 1183
rect 2412 1180 2507 1182
rect 2412 1179 2413 1180
rect 2407 1178 2413 1179
rect 2506 1179 2507 1180
rect 2511 1182 2512 1183
rect 2559 1183 2565 1184
rect 2559 1182 2560 1183
rect 2511 1180 2560 1182
rect 2511 1179 2512 1180
rect 2506 1178 2512 1179
rect 2559 1179 2560 1180
rect 2564 1182 2565 1183
rect 2702 1183 2703 1187
rect 2708 1186 2709 1187
rect 2720 1186 2722 1198
rect 2708 1184 2722 1186
rect 2846 1189 2852 1190
rect 2846 1185 2847 1189
rect 2851 1185 2852 1189
rect 2846 1184 2852 1185
rect 2854 1187 2861 1188
rect 2708 1183 2709 1184
rect 2702 1182 2709 1183
rect 2854 1183 2855 1187
rect 2860 1186 2861 1187
rect 2929 1186 2931 1198
rect 2860 1184 2931 1186
rect 2998 1189 3004 1190
rect 2998 1185 2999 1189
rect 3003 1185 3004 1189
rect 2998 1184 3004 1185
rect 3190 1185 3196 1186
rect 2860 1183 2861 1184
rect 2854 1182 2861 1183
rect 3006 1183 3013 1184
rect 2564 1180 2706 1182
rect 2564 1179 2565 1180
rect 2559 1178 2565 1179
rect 3006 1179 3007 1183
rect 3012 1179 3013 1183
rect 3190 1181 3191 1185
rect 3195 1181 3196 1185
rect 3190 1180 3196 1181
rect 3006 1178 3013 1179
rect 110 1171 116 1172
rect 110 1167 111 1171
rect 115 1167 116 1171
rect 1230 1171 1237 1172
rect 110 1166 116 1167
rect 726 1167 732 1168
rect 726 1163 727 1167
rect 731 1163 732 1167
rect 726 1162 732 1163
rect 734 1167 741 1168
rect 734 1163 735 1167
rect 740 1163 741 1167
rect 734 1162 741 1163
rect 854 1167 860 1168
rect 854 1163 855 1167
rect 859 1163 860 1167
rect 854 1162 860 1163
rect 863 1167 872 1168
rect 863 1163 864 1167
rect 871 1163 872 1167
rect 863 1162 872 1163
rect 982 1167 988 1168
rect 982 1163 983 1167
rect 987 1163 988 1167
rect 982 1162 988 1163
rect 991 1167 997 1168
rect 991 1163 992 1167
rect 996 1166 997 1167
rect 1006 1167 1012 1168
rect 1006 1166 1007 1167
rect 996 1164 1007 1166
rect 996 1163 997 1164
rect 991 1162 997 1163
rect 1006 1163 1007 1164
rect 1011 1163 1012 1167
rect 1006 1162 1012 1163
rect 1102 1167 1108 1168
rect 1102 1163 1103 1167
rect 1107 1163 1108 1167
rect 1102 1162 1108 1163
rect 1110 1167 1117 1168
rect 1110 1163 1111 1167
rect 1116 1163 1117 1167
rect 1110 1162 1117 1163
rect 1222 1167 1228 1168
rect 1222 1163 1223 1167
rect 1227 1163 1228 1167
rect 1230 1167 1231 1171
rect 1236 1170 1237 1171
rect 1254 1171 1260 1172
rect 1254 1170 1255 1171
rect 1236 1168 1255 1170
rect 1236 1167 1237 1168
rect 1230 1166 1237 1167
rect 1254 1167 1255 1168
rect 1259 1167 1260 1171
rect 1575 1171 1581 1172
rect 1254 1166 1260 1167
rect 1334 1167 1340 1168
rect 1222 1162 1228 1163
rect 1334 1163 1335 1167
rect 1339 1163 1340 1167
rect 1334 1162 1340 1163
rect 1343 1167 1349 1168
rect 1343 1163 1344 1167
rect 1348 1163 1349 1167
rect 1343 1162 1349 1163
rect 1446 1167 1452 1168
rect 1446 1163 1447 1167
rect 1451 1163 1452 1167
rect 1446 1162 1452 1163
rect 1454 1167 1461 1168
rect 1454 1163 1455 1167
rect 1460 1163 1461 1167
rect 1454 1162 1461 1163
rect 1566 1167 1572 1168
rect 1566 1163 1567 1167
rect 1571 1163 1572 1167
rect 1575 1167 1576 1171
rect 1580 1170 1581 1171
rect 1606 1171 1612 1172
rect 1606 1170 1607 1171
rect 1580 1168 1607 1170
rect 1580 1167 1581 1168
rect 1575 1166 1581 1167
rect 1606 1167 1607 1168
rect 1611 1167 1612 1171
rect 1606 1166 1612 1167
rect 1630 1171 1636 1172
rect 1630 1167 1631 1171
rect 1635 1167 1636 1171
rect 1630 1166 1636 1167
rect 1670 1167 1676 1168
rect 1566 1162 1572 1163
rect 1670 1163 1671 1167
rect 1675 1163 1676 1167
rect 1670 1162 1676 1163
rect 3190 1167 3196 1168
rect 3190 1163 3191 1167
rect 3195 1163 3196 1167
rect 3190 1162 3196 1163
rect 2246 1160 2252 1161
rect 2246 1156 2247 1160
rect 2251 1156 2252 1160
rect 2246 1155 2252 1156
rect 2398 1160 2404 1161
rect 2398 1156 2399 1160
rect 2403 1156 2404 1160
rect 2398 1155 2404 1156
rect 2550 1160 2556 1161
rect 2550 1156 2551 1160
rect 2555 1156 2556 1160
rect 2550 1155 2556 1156
rect 2694 1160 2700 1161
rect 2694 1156 2695 1160
rect 2699 1156 2700 1160
rect 2694 1155 2700 1156
rect 2846 1160 2852 1161
rect 2846 1156 2847 1160
rect 2851 1156 2852 1160
rect 2846 1155 2852 1156
rect 2998 1160 3004 1161
rect 2998 1156 2999 1160
rect 3003 1156 3004 1160
rect 2998 1155 3004 1156
rect 2174 1148 2180 1149
rect 630 1145 636 1146
rect 110 1141 116 1142
rect 110 1137 111 1141
rect 115 1137 116 1141
rect 630 1141 631 1145
rect 635 1141 636 1145
rect 630 1140 636 1141
rect 758 1145 764 1146
rect 758 1141 759 1145
rect 763 1141 764 1145
rect 758 1140 764 1141
rect 878 1145 884 1146
rect 878 1141 879 1145
rect 883 1141 884 1145
rect 878 1140 884 1141
rect 998 1145 1004 1146
rect 998 1141 999 1145
rect 1003 1141 1004 1145
rect 998 1140 1004 1141
rect 1118 1145 1124 1146
rect 1118 1141 1119 1145
rect 1123 1141 1124 1145
rect 1118 1140 1124 1141
rect 1230 1145 1236 1146
rect 1230 1141 1231 1145
rect 1235 1141 1236 1145
rect 1230 1140 1236 1141
rect 1342 1145 1348 1146
rect 1342 1141 1343 1145
rect 1347 1141 1348 1145
rect 1342 1140 1348 1141
rect 1462 1145 1468 1146
rect 1462 1141 1463 1145
rect 1467 1141 1468 1145
rect 2174 1144 2175 1148
rect 2179 1144 2180 1148
rect 2174 1143 2180 1144
rect 2334 1148 2340 1149
rect 2334 1144 2335 1148
rect 2339 1144 2340 1148
rect 2334 1143 2340 1144
rect 2494 1148 2500 1149
rect 2494 1144 2495 1148
rect 2499 1144 2500 1148
rect 2494 1143 2500 1144
rect 2654 1148 2660 1149
rect 2654 1144 2655 1148
rect 2659 1144 2660 1148
rect 2654 1143 2660 1144
rect 2814 1148 2820 1149
rect 2814 1144 2815 1148
rect 2819 1144 2820 1148
rect 2814 1143 2820 1144
rect 2974 1148 2980 1149
rect 2974 1144 2975 1148
rect 2979 1144 2980 1148
rect 2974 1143 2980 1144
rect 3134 1148 3140 1149
rect 3134 1144 3135 1148
rect 3139 1144 3140 1148
rect 3134 1143 3140 1144
rect 1462 1140 1468 1141
rect 1630 1141 1636 1142
rect 110 1136 116 1137
rect 638 1139 645 1140
rect 638 1135 639 1139
rect 644 1138 645 1139
rect 670 1139 676 1140
rect 670 1138 671 1139
rect 644 1136 671 1138
rect 644 1135 645 1136
rect 638 1134 645 1135
rect 670 1135 671 1136
rect 675 1138 676 1139
rect 734 1139 740 1140
rect 734 1138 735 1139
rect 675 1136 735 1138
rect 675 1135 676 1136
rect 670 1134 676 1135
rect 734 1135 735 1136
rect 739 1138 740 1139
rect 767 1139 773 1140
rect 767 1138 768 1139
rect 739 1136 768 1138
rect 739 1135 740 1136
rect 734 1134 740 1135
rect 767 1135 768 1136
rect 772 1138 773 1139
rect 782 1139 788 1140
rect 782 1138 783 1139
rect 772 1136 783 1138
rect 772 1135 773 1136
rect 767 1134 773 1135
rect 782 1135 783 1136
rect 787 1135 788 1139
rect 782 1134 788 1135
rect 866 1139 872 1140
rect 866 1135 867 1139
rect 871 1138 872 1139
rect 887 1139 893 1140
rect 887 1138 888 1139
rect 871 1136 888 1138
rect 871 1135 872 1136
rect 866 1134 872 1135
rect 887 1135 888 1136
rect 892 1138 893 1139
rect 906 1139 912 1140
rect 906 1138 907 1139
rect 892 1136 907 1138
rect 892 1135 893 1136
rect 887 1134 893 1135
rect 906 1135 907 1136
rect 911 1135 912 1139
rect 906 1134 912 1135
rect 1006 1139 1013 1140
rect 1006 1135 1007 1139
rect 1012 1138 1013 1139
rect 1110 1139 1116 1140
rect 1110 1138 1111 1139
rect 1012 1136 1111 1138
rect 1012 1135 1013 1136
rect 1006 1134 1013 1135
rect 1110 1135 1111 1136
rect 1115 1138 1116 1139
rect 1127 1139 1133 1140
rect 1127 1138 1128 1139
rect 1115 1136 1128 1138
rect 1115 1135 1116 1136
rect 1110 1134 1116 1135
rect 1127 1135 1128 1136
rect 1132 1135 1133 1139
rect 1127 1134 1133 1135
rect 1239 1139 1245 1140
rect 1239 1135 1240 1139
rect 1244 1138 1245 1139
rect 1254 1139 1260 1140
rect 1254 1138 1255 1139
rect 1244 1136 1255 1138
rect 1244 1135 1245 1136
rect 1239 1134 1245 1135
rect 1254 1135 1255 1136
rect 1259 1138 1260 1139
rect 1350 1139 1357 1140
rect 1350 1138 1351 1139
rect 1259 1136 1351 1138
rect 1259 1135 1260 1136
rect 1254 1134 1260 1135
rect 1350 1135 1351 1136
rect 1356 1138 1357 1139
rect 1454 1139 1460 1140
rect 1454 1138 1455 1139
rect 1356 1136 1455 1138
rect 1356 1135 1357 1136
rect 1350 1134 1357 1135
rect 1454 1135 1455 1136
rect 1459 1138 1460 1139
rect 1471 1139 1477 1140
rect 1471 1138 1472 1139
rect 1459 1136 1472 1138
rect 1459 1135 1460 1136
rect 1454 1134 1460 1135
rect 1471 1135 1472 1136
rect 1476 1135 1477 1139
rect 1630 1137 1631 1141
rect 1635 1137 1636 1141
rect 1630 1136 1636 1137
rect 1670 1141 1676 1142
rect 1670 1137 1671 1141
rect 1675 1137 1676 1141
rect 1670 1136 1676 1137
rect 3190 1141 3196 1142
rect 3190 1137 3191 1141
rect 3195 1137 3196 1141
rect 3190 1136 3196 1137
rect 1471 1134 1477 1135
rect 110 1123 116 1124
rect 110 1119 111 1123
rect 115 1119 116 1123
rect 110 1118 116 1119
rect 1630 1123 1636 1124
rect 1630 1119 1631 1123
rect 1635 1119 1636 1123
rect 1630 1118 1636 1119
rect 1670 1123 1676 1124
rect 1670 1119 1671 1123
rect 1675 1119 1676 1123
rect 2343 1123 2349 1124
rect 1670 1118 1676 1119
rect 2174 1119 2180 1120
rect 630 1116 636 1117
rect 630 1112 631 1116
rect 635 1112 636 1116
rect 630 1111 636 1112
rect 758 1116 764 1117
rect 758 1112 759 1116
rect 763 1112 764 1116
rect 758 1111 764 1112
rect 878 1116 884 1117
rect 878 1112 879 1116
rect 883 1112 884 1116
rect 878 1111 884 1112
rect 998 1116 1004 1117
rect 998 1112 999 1116
rect 1003 1112 1004 1116
rect 998 1111 1004 1112
rect 1118 1116 1124 1117
rect 1118 1112 1119 1116
rect 1123 1112 1124 1116
rect 1118 1111 1124 1112
rect 1230 1116 1236 1117
rect 1230 1112 1231 1116
rect 1235 1112 1236 1116
rect 1230 1111 1236 1112
rect 1342 1116 1348 1117
rect 1342 1112 1343 1116
rect 1347 1112 1348 1116
rect 1342 1111 1348 1112
rect 1462 1116 1468 1117
rect 1462 1112 1463 1116
rect 1467 1112 1468 1116
rect 2174 1115 2175 1119
rect 2179 1115 2180 1119
rect 2174 1114 2180 1115
rect 2182 1119 2189 1120
rect 2182 1115 2183 1119
rect 2188 1115 2189 1119
rect 2182 1114 2189 1115
rect 2334 1119 2340 1120
rect 2334 1115 2335 1119
rect 2339 1115 2340 1119
rect 2343 1119 2344 1123
rect 2348 1122 2349 1123
rect 2351 1123 2357 1124
rect 2351 1122 2352 1123
rect 2348 1120 2352 1122
rect 2348 1119 2349 1120
rect 2343 1118 2349 1119
rect 2351 1119 2352 1120
rect 2356 1119 2357 1123
rect 2503 1123 2512 1124
rect 2351 1118 2357 1119
rect 2494 1119 2500 1120
rect 2334 1114 2340 1115
rect 2494 1115 2495 1119
rect 2499 1115 2500 1119
rect 2503 1119 2504 1123
rect 2511 1119 2512 1123
rect 2662 1123 2669 1124
rect 2503 1118 2512 1119
rect 2654 1119 2660 1120
rect 2494 1114 2500 1115
rect 2654 1115 2655 1119
rect 2659 1115 2660 1119
rect 2662 1119 2663 1123
rect 2668 1122 2669 1123
rect 2702 1123 2708 1124
rect 2702 1122 2703 1123
rect 2668 1120 2703 1122
rect 2668 1119 2669 1120
rect 2662 1118 2669 1119
rect 2702 1119 2703 1120
rect 2707 1119 2708 1123
rect 2822 1123 2829 1124
rect 2702 1118 2708 1119
rect 2814 1119 2820 1120
rect 2654 1114 2660 1115
rect 2814 1115 2815 1119
rect 2819 1115 2820 1119
rect 2822 1119 2823 1123
rect 2828 1122 2829 1123
rect 2854 1123 2860 1124
rect 2854 1122 2855 1123
rect 2828 1120 2855 1122
rect 2828 1119 2829 1120
rect 2822 1118 2829 1119
rect 2854 1119 2855 1120
rect 2859 1119 2860 1123
rect 2983 1123 2989 1124
rect 2854 1118 2860 1119
rect 2974 1119 2980 1120
rect 2814 1114 2820 1115
rect 2974 1115 2975 1119
rect 2979 1115 2980 1119
rect 2983 1119 2984 1123
rect 2988 1122 2989 1123
rect 3006 1123 3012 1124
rect 3006 1122 3007 1123
rect 2988 1120 3007 1122
rect 2988 1119 2989 1120
rect 2983 1118 2989 1119
rect 3006 1119 3007 1120
rect 3011 1119 3012 1123
rect 3142 1123 3149 1124
rect 3006 1118 3012 1119
rect 3134 1119 3140 1120
rect 2974 1114 2980 1115
rect 3134 1115 3135 1119
rect 3139 1115 3140 1119
rect 3142 1119 3143 1123
rect 3148 1119 3149 1123
rect 3142 1118 3149 1119
rect 3190 1123 3196 1124
rect 3190 1119 3191 1123
rect 3195 1119 3196 1123
rect 3190 1118 3196 1119
rect 3134 1114 3140 1115
rect 1462 1111 1468 1112
rect 2070 1105 2076 1106
rect 1670 1101 1676 1102
rect 1670 1097 1671 1101
rect 1675 1097 1676 1101
rect 2070 1101 2071 1105
rect 2075 1101 2076 1105
rect 2070 1100 2076 1101
rect 2190 1105 2196 1106
rect 2190 1101 2191 1105
rect 2195 1101 2196 1105
rect 2190 1100 2196 1101
rect 2326 1105 2332 1106
rect 2326 1101 2327 1105
rect 2331 1101 2332 1105
rect 2478 1105 2484 1106
rect 2326 1100 2332 1101
rect 2335 1103 2341 1104
rect 1670 1096 1676 1097
rect 2078 1099 2085 1100
rect 2078 1095 2079 1099
rect 2084 1098 2085 1099
rect 2182 1099 2188 1100
rect 2182 1098 2183 1099
rect 2084 1096 2183 1098
rect 2084 1095 2085 1096
rect 2078 1094 2085 1095
rect 2182 1095 2183 1096
rect 2187 1098 2188 1099
rect 2199 1099 2205 1100
rect 2199 1098 2200 1099
rect 2187 1096 2200 1098
rect 2187 1095 2188 1096
rect 2182 1094 2188 1095
rect 2199 1095 2200 1096
rect 2204 1095 2205 1099
rect 2335 1099 2336 1103
rect 2340 1102 2341 1103
rect 2350 1103 2357 1104
rect 2350 1102 2351 1103
rect 2340 1100 2351 1102
rect 2340 1099 2341 1100
rect 2335 1098 2341 1099
rect 2350 1099 2351 1100
rect 2356 1099 2357 1103
rect 2478 1101 2479 1105
rect 2483 1101 2484 1105
rect 2638 1105 2644 1106
rect 2478 1100 2484 1101
rect 2487 1103 2493 1104
rect 2350 1098 2357 1099
rect 2487 1099 2488 1103
rect 2492 1102 2493 1103
rect 2506 1103 2512 1104
rect 2506 1102 2507 1103
rect 2492 1100 2507 1102
rect 2492 1099 2493 1100
rect 2487 1098 2493 1099
rect 2506 1099 2507 1100
rect 2511 1099 2512 1103
rect 2638 1101 2639 1105
rect 2643 1101 2644 1105
rect 2814 1105 2820 1106
rect 2638 1100 2644 1101
rect 2647 1103 2653 1104
rect 2506 1098 2512 1099
rect 2647 1099 2648 1103
rect 2652 1102 2653 1103
rect 2662 1103 2668 1104
rect 2662 1102 2663 1103
rect 2652 1100 2663 1102
rect 2652 1099 2653 1100
rect 2647 1098 2653 1099
rect 2662 1099 2663 1100
rect 2667 1099 2668 1103
rect 2814 1101 2815 1105
rect 2819 1101 2820 1105
rect 2998 1105 3004 1106
rect 2814 1100 2820 1101
rect 2822 1103 2829 1104
rect 2662 1098 2668 1099
rect 2822 1099 2823 1103
rect 2828 1099 2829 1103
rect 2998 1101 2999 1105
rect 3003 1101 3004 1105
rect 2998 1100 3004 1101
rect 3158 1105 3164 1106
rect 3158 1101 3159 1105
rect 3163 1101 3164 1105
rect 3158 1100 3164 1101
rect 3190 1101 3196 1102
rect 2822 1098 2829 1099
rect 3006 1099 3013 1100
rect 2199 1094 2205 1095
rect 3006 1095 3007 1099
rect 3012 1095 3013 1099
rect 3006 1094 3013 1095
rect 3142 1099 3148 1100
rect 3142 1095 3143 1099
rect 3147 1098 3148 1099
rect 3166 1099 3173 1100
rect 3166 1098 3167 1099
rect 3147 1096 3167 1098
rect 3147 1095 3148 1096
rect 3142 1094 3148 1095
rect 3166 1095 3167 1096
rect 3172 1095 3173 1099
rect 3190 1097 3191 1101
rect 3195 1097 3196 1101
rect 3190 1096 3196 1097
rect 3166 1094 3173 1095
rect 526 1092 532 1093
rect 526 1088 527 1092
rect 531 1088 532 1092
rect 526 1087 532 1088
rect 654 1092 660 1093
rect 654 1088 655 1092
rect 659 1088 660 1092
rect 654 1087 660 1088
rect 774 1092 780 1093
rect 774 1088 775 1092
rect 779 1088 780 1092
rect 774 1087 780 1088
rect 894 1092 900 1093
rect 894 1088 895 1092
rect 899 1088 900 1092
rect 894 1087 900 1088
rect 1014 1092 1020 1093
rect 1014 1088 1015 1092
rect 1019 1088 1020 1092
rect 1014 1087 1020 1088
rect 1126 1092 1132 1093
rect 1126 1088 1127 1092
rect 1131 1088 1132 1092
rect 1126 1087 1132 1088
rect 1246 1092 1252 1093
rect 1246 1088 1247 1092
rect 1251 1088 1252 1092
rect 1246 1087 1252 1088
rect 1366 1092 1372 1093
rect 1366 1088 1367 1092
rect 1371 1088 1372 1092
rect 1366 1087 1372 1088
rect 110 1085 116 1086
rect 110 1081 111 1085
rect 115 1081 116 1085
rect 110 1080 116 1081
rect 1630 1085 1636 1086
rect 1630 1081 1631 1085
rect 1635 1081 1636 1085
rect 1630 1080 1636 1081
rect 1670 1083 1676 1084
rect 1670 1079 1671 1083
rect 1675 1079 1676 1083
rect 1670 1078 1676 1079
rect 3190 1083 3196 1084
rect 3190 1079 3191 1083
rect 3195 1079 3196 1083
rect 3190 1078 3196 1079
rect 2070 1076 2076 1077
rect 2070 1072 2071 1076
rect 2075 1072 2076 1076
rect 2070 1071 2076 1072
rect 2190 1076 2196 1077
rect 2190 1072 2191 1076
rect 2195 1072 2196 1076
rect 2190 1071 2196 1072
rect 2326 1076 2332 1077
rect 2326 1072 2327 1076
rect 2331 1072 2332 1076
rect 2326 1071 2332 1072
rect 2478 1076 2484 1077
rect 2478 1072 2479 1076
rect 2483 1072 2484 1076
rect 2478 1071 2484 1072
rect 2638 1076 2644 1077
rect 2638 1072 2639 1076
rect 2643 1072 2644 1076
rect 2638 1071 2644 1072
rect 2814 1076 2820 1077
rect 2814 1072 2815 1076
rect 2819 1072 2820 1076
rect 2814 1071 2820 1072
rect 2998 1076 3004 1077
rect 2998 1072 2999 1076
rect 3003 1072 3004 1076
rect 2998 1071 3004 1072
rect 3158 1076 3164 1077
rect 3158 1072 3159 1076
rect 3163 1072 3164 1076
rect 3158 1071 3164 1072
rect 1257 1068 1379 1070
rect 110 1067 116 1068
rect 110 1063 111 1067
rect 115 1063 116 1067
rect 782 1067 789 1068
rect 110 1062 116 1063
rect 526 1063 532 1064
rect 526 1059 527 1063
rect 531 1059 532 1063
rect 526 1058 532 1059
rect 534 1063 541 1064
rect 534 1059 535 1063
rect 540 1059 541 1063
rect 534 1058 541 1059
rect 654 1063 660 1064
rect 654 1059 655 1063
rect 659 1059 660 1063
rect 654 1058 660 1059
rect 663 1063 669 1064
rect 663 1059 664 1063
rect 668 1059 669 1063
rect 663 1058 669 1059
rect 774 1063 780 1064
rect 774 1059 775 1063
rect 779 1059 780 1063
rect 782 1063 783 1067
rect 788 1063 789 1067
rect 1257 1064 1259 1068
rect 1375 1067 1381 1068
rect 782 1062 789 1063
rect 894 1063 900 1064
rect 774 1058 780 1059
rect 894 1059 895 1063
rect 899 1059 900 1063
rect 894 1058 900 1059
rect 903 1063 912 1064
rect 903 1059 904 1063
rect 911 1059 912 1063
rect 903 1058 912 1059
rect 1014 1063 1020 1064
rect 1014 1059 1015 1063
rect 1019 1059 1020 1063
rect 1014 1058 1020 1059
rect 1023 1063 1029 1064
rect 1023 1059 1024 1063
rect 1028 1062 1029 1063
rect 1038 1063 1044 1064
rect 1038 1062 1039 1063
rect 1028 1060 1039 1062
rect 1028 1059 1029 1060
rect 1023 1058 1029 1059
rect 1038 1059 1039 1060
rect 1043 1059 1044 1063
rect 1038 1058 1044 1059
rect 1126 1063 1132 1064
rect 1126 1059 1127 1063
rect 1131 1059 1132 1063
rect 1126 1058 1132 1059
rect 1134 1063 1141 1064
rect 1134 1059 1135 1063
rect 1140 1059 1141 1063
rect 1134 1058 1141 1059
rect 1246 1063 1252 1064
rect 1246 1059 1247 1063
rect 1251 1059 1252 1063
rect 1246 1058 1252 1059
rect 1254 1063 1261 1064
rect 1254 1059 1255 1063
rect 1260 1059 1261 1063
rect 1254 1058 1261 1059
rect 1366 1063 1372 1064
rect 1366 1059 1367 1063
rect 1371 1059 1372 1063
rect 1375 1063 1376 1067
rect 1380 1063 1381 1067
rect 1375 1062 1381 1063
rect 1630 1067 1636 1068
rect 1630 1063 1631 1067
rect 1635 1063 1636 1067
rect 1630 1062 1636 1063
rect 1366 1058 1372 1059
rect 582 1055 588 1056
rect 582 1051 583 1055
rect 587 1054 588 1055
rect 638 1055 644 1056
rect 638 1054 639 1055
rect 587 1052 639 1054
rect 587 1051 588 1052
rect 582 1050 588 1051
rect 638 1051 639 1052
rect 643 1054 644 1055
rect 664 1054 666 1058
rect 643 1052 666 1054
rect 643 1051 644 1052
rect 638 1050 644 1051
rect 664 1050 666 1052
rect 1974 1052 1980 1053
rect 664 1048 690 1050
rect 422 1045 428 1046
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 422 1041 423 1045
rect 427 1041 428 1045
rect 422 1040 428 1041
rect 550 1045 556 1046
rect 550 1041 551 1045
rect 555 1041 556 1045
rect 550 1040 556 1041
rect 678 1045 684 1046
rect 678 1041 679 1045
rect 683 1041 684 1045
rect 688 1044 690 1048
rect 1974 1048 1975 1052
rect 1979 1048 1980 1052
rect 1974 1047 1980 1048
rect 2094 1052 2100 1053
rect 2094 1048 2095 1052
rect 2099 1048 2100 1052
rect 2094 1047 2100 1048
rect 2214 1052 2220 1053
rect 2214 1048 2215 1052
rect 2219 1048 2220 1052
rect 2214 1047 2220 1048
rect 2342 1052 2348 1053
rect 2342 1048 2343 1052
rect 2347 1048 2348 1052
rect 2342 1047 2348 1048
rect 2486 1052 2492 1053
rect 2486 1048 2487 1052
rect 2491 1048 2492 1052
rect 2486 1047 2492 1048
rect 2646 1052 2652 1053
rect 2646 1048 2647 1052
rect 2651 1048 2652 1052
rect 2646 1047 2652 1048
rect 2822 1052 2828 1053
rect 2822 1048 2823 1052
rect 2827 1048 2828 1052
rect 2822 1047 2828 1048
rect 2998 1052 3004 1053
rect 2998 1048 2999 1052
rect 3003 1048 3004 1052
rect 2998 1047 3004 1048
rect 3158 1052 3164 1053
rect 3158 1048 3159 1052
rect 3163 1048 3164 1052
rect 3158 1047 3164 1048
rect 798 1045 804 1046
rect 678 1040 684 1041
rect 687 1043 693 1044
rect 110 1036 116 1037
rect 431 1039 437 1040
rect 431 1035 432 1039
rect 436 1038 437 1039
rect 462 1039 468 1040
rect 462 1038 463 1039
rect 436 1036 463 1038
rect 436 1035 437 1036
rect 431 1034 437 1035
rect 462 1035 463 1036
rect 467 1038 468 1039
rect 534 1039 540 1040
rect 534 1038 535 1039
rect 467 1036 535 1038
rect 467 1035 468 1036
rect 462 1034 468 1035
rect 534 1035 535 1036
rect 539 1038 540 1039
rect 559 1039 565 1040
rect 559 1038 560 1039
rect 539 1036 560 1038
rect 539 1035 540 1036
rect 534 1034 540 1035
rect 559 1035 560 1036
rect 564 1038 565 1039
rect 582 1039 588 1040
rect 582 1038 583 1039
rect 564 1036 583 1038
rect 564 1035 565 1036
rect 559 1034 565 1035
rect 582 1035 583 1036
rect 587 1035 588 1039
rect 687 1039 688 1043
rect 692 1042 693 1043
rect 702 1043 708 1044
rect 702 1042 703 1043
rect 692 1040 703 1042
rect 692 1039 693 1040
rect 687 1038 693 1039
rect 702 1039 703 1040
rect 707 1039 708 1043
rect 798 1041 799 1045
rect 803 1041 804 1045
rect 798 1040 804 1041
rect 918 1045 924 1046
rect 918 1041 919 1045
rect 923 1041 924 1045
rect 918 1040 924 1041
rect 1030 1045 1036 1046
rect 1030 1041 1031 1045
rect 1035 1041 1036 1045
rect 1030 1040 1036 1041
rect 1142 1045 1148 1046
rect 1142 1041 1143 1045
rect 1147 1041 1148 1045
rect 1142 1040 1148 1041
rect 1262 1045 1268 1046
rect 1262 1041 1263 1045
rect 1267 1041 1268 1045
rect 1670 1045 1676 1046
rect 1262 1040 1268 1041
rect 1630 1041 1636 1042
rect 702 1038 708 1039
rect 782 1039 788 1040
rect 582 1034 588 1035
rect 782 1035 783 1039
rect 787 1038 788 1039
rect 807 1039 813 1040
rect 807 1038 808 1039
rect 787 1036 808 1038
rect 787 1035 788 1036
rect 782 1034 788 1035
rect 807 1035 808 1036
rect 812 1035 813 1039
rect 807 1034 813 1035
rect 906 1039 912 1040
rect 906 1035 907 1039
rect 911 1038 912 1039
rect 927 1039 933 1040
rect 927 1038 928 1039
rect 911 1036 928 1038
rect 911 1035 912 1036
rect 906 1034 912 1035
rect 927 1035 928 1036
rect 932 1038 933 1039
rect 1038 1039 1045 1040
rect 1038 1038 1039 1039
rect 932 1036 1039 1038
rect 932 1035 933 1036
rect 927 1034 933 1035
rect 1038 1035 1039 1036
rect 1044 1038 1045 1039
rect 1134 1039 1140 1040
rect 1134 1038 1135 1039
rect 1044 1036 1135 1038
rect 1044 1035 1045 1036
rect 1038 1034 1045 1035
rect 1134 1035 1135 1036
rect 1139 1038 1140 1039
rect 1151 1039 1157 1040
rect 1151 1038 1152 1039
rect 1139 1036 1152 1038
rect 1139 1035 1140 1036
rect 1134 1034 1140 1035
rect 1151 1035 1152 1036
rect 1156 1038 1157 1039
rect 1166 1039 1172 1040
rect 1166 1038 1167 1039
rect 1156 1036 1167 1038
rect 1156 1035 1157 1036
rect 1151 1034 1157 1035
rect 1166 1035 1167 1036
rect 1171 1038 1172 1039
rect 1254 1039 1260 1040
rect 1254 1038 1255 1039
rect 1171 1036 1255 1038
rect 1171 1035 1172 1036
rect 1166 1034 1172 1035
rect 1254 1035 1255 1036
rect 1259 1038 1260 1039
rect 1271 1039 1277 1040
rect 1271 1038 1272 1039
rect 1259 1036 1272 1038
rect 1259 1035 1260 1036
rect 1254 1034 1260 1035
rect 1271 1035 1272 1036
rect 1276 1035 1277 1039
rect 1630 1037 1631 1041
rect 1635 1037 1636 1041
rect 1670 1041 1671 1045
rect 1675 1041 1676 1045
rect 1670 1040 1676 1041
rect 3190 1045 3196 1046
rect 3190 1041 3191 1045
rect 3195 1041 3196 1045
rect 3190 1040 3196 1041
rect 1630 1036 1636 1037
rect 1271 1034 1277 1035
rect 3006 1031 3012 1032
rect 3006 1030 3007 1031
rect 2833 1028 3007 1030
rect 1670 1027 1676 1028
rect 110 1023 116 1024
rect 110 1019 111 1023
rect 115 1019 116 1023
rect 110 1018 116 1019
rect 1630 1023 1636 1024
rect 1630 1019 1631 1023
rect 1635 1019 1636 1023
rect 1670 1023 1671 1027
rect 1675 1023 1676 1027
rect 2350 1027 2357 1028
rect 1670 1022 1676 1023
rect 1974 1023 1980 1024
rect 1630 1018 1636 1019
rect 1974 1019 1975 1023
rect 1979 1019 1980 1023
rect 1974 1018 1980 1019
rect 1983 1023 1989 1024
rect 1983 1019 1984 1023
rect 1988 1019 1989 1023
rect 1983 1018 1989 1019
rect 2094 1023 2100 1024
rect 2094 1019 2095 1023
rect 2099 1019 2100 1023
rect 2094 1018 2100 1019
rect 2103 1023 2109 1024
rect 2103 1019 2104 1023
rect 2108 1019 2109 1023
rect 2103 1018 2109 1019
rect 2214 1023 2220 1024
rect 2214 1019 2215 1023
rect 2219 1019 2220 1023
rect 2214 1018 2220 1019
rect 2223 1023 2229 1024
rect 2223 1019 2224 1023
rect 2228 1019 2229 1023
rect 2223 1018 2229 1019
rect 2342 1023 2348 1024
rect 2342 1019 2343 1023
rect 2347 1019 2348 1023
rect 2350 1023 2351 1027
rect 2356 1023 2357 1027
rect 2830 1027 2837 1028
rect 2350 1022 2357 1023
rect 2486 1023 2492 1024
rect 2342 1018 2348 1019
rect 2486 1019 2487 1023
rect 2491 1019 2492 1023
rect 2486 1018 2492 1019
rect 2495 1023 2501 1024
rect 2495 1019 2496 1023
rect 2500 1019 2501 1023
rect 2495 1018 2501 1019
rect 2646 1023 2652 1024
rect 2646 1019 2647 1023
rect 2651 1019 2652 1023
rect 2646 1018 2652 1019
rect 2654 1023 2661 1024
rect 2654 1019 2655 1023
rect 2660 1019 2661 1023
rect 2654 1018 2661 1019
rect 2822 1023 2828 1024
rect 2822 1019 2823 1023
rect 2827 1019 2828 1023
rect 2830 1023 2831 1027
rect 2836 1023 2837 1027
rect 3006 1027 3007 1028
rect 3011 1030 3012 1031
rect 3011 1028 3170 1030
rect 3011 1027 3013 1028
rect 3006 1026 3008 1027
rect 2830 1022 2837 1023
rect 2998 1023 3004 1024
rect 2822 1018 2828 1019
rect 2998 1019 2999 1023
rect 3003 1019 3004 1023
rect 3007 1023 3008 1026
rect 3012 1023 3013 1027
rect 3166 1027 3173 1028
rect 3007 1022 3013 1023
rect 3158 1023 3164 1024
rect 2998 1018 3004 1019
rect 3158 1019 3159 1023
rect 3163 1019 3164 1023
rect 3166 1023 3167 1027
rect 3172 1023 3173 1027
rect 3166 1022 3173 1023
rect 3190 1027 3196 1028
rect 3190 1023 3191 1027
rect 3195 1023 3196 1027
rect 3190 1022 3196 1023
rect 3158 1018 3164 1019
rect 422 1016 428 1017
rect 422 1012 423 1016
rect 427 1012 428 1016
rect 422 1011 428 1012
rect 550 1016 556 1017
rect 550 1012 551 1016
rect 555 1012 556 1016
rect 550 1011 556 1012
rect 678 1016 684 1017
rect 678 1012 679 1016
rect 683 1012 684 1016
rect 678 1011 684 1012
rect 798 1016 804 1017
rect 798 1012 799 1016
rect 803 1012 804 1016
rect 798 1011 804 1012
rect 918 1016 924 1017
rect 918 1012 919 1016
rect 923 1012 924 1016
rect 918 1011 924 1012
rect 1030 1016 1036 1017
rect 1030 1012 1031 1016
rect 1035 1012 1036 1016
rect 1030 1011 1036 1012
rect 1142 1016 1148 1017
rect 1142 1012 1143 1016
rect 1147 1012 1148 1016
rect 1142 1011 1148 1012
rect 1262 1016 1268 1017
rect 1262 1012 1263 1016
rect 1267 1012 1268 1016
rect 1262 1011 1268 1012
rect 1926 1015 1932 1016
rect 1926 1011 1927 1015
rect 1931 1014 1932 1015
rect 1985 1014 1987 1018
rect 2078 1015 2084 1016
rect 2078 1014 2079 1015
rect 1931 1012 2079 1014
rect 1931 1011 1932 1012
rect 1926 1010 1932 1011
rect 1894 1009 1900 1010
rect 1670 1005 1676 1006
rect 1670 1001 1671 1005
rect 1675 1001 1676 1005
rect 1894 1005 1895 1009
rect 1899 1005 1900 1009
rect 1894 1004 1900 1005
rect 2046 1009 2052 1010
rect 2046 1005 2047 1009
rect 2051 1005 2052 1009
rect 2057 1008 2059 1012
rect 2078 1011 2079 1012
rect 2083 1014 2084 1015
rect 2105 1014 2107 1018
rect 2225 1014 2227 1018
rect 2230 1015 2236 1016
rect 2230 1014 2231 1015
rect 2083 1012 2231 1014
rect 2083 1011 2084 1012
rect 2078 1010 2084 1011
rect 2198 1009 2204 1010
rect 2046 1004 2052 1005
rect 2055 1007 2061 1008
rect 1670 1000 1676 1001
rect 1903 1003 1909 1004
rect 1903 999 1904 1003
rect 1908 1002 1909 1003
rect 1926 1003 1932 1004
rect 1926 1002 1927 1003
rect 1908 1000 1927 1002
rect 1908 999 1909 1000
rect 1903 998 1909 999
rect 1926 999 1927 1000
rect 1931 999 1932 1003
rect 2055 1003 2056 1007
rect 2060 1003 2061 1007
rect 2198 1005 2199 1009
rect 2203 1005 2204 1009
rect 2209 1008 2211 1012
rect 2230 1011 2231 1012
rect 2235 1011 2236 1015
rect 2496 1014 2498 1018
rect 2496 1012 2507 1014
rect 2230 1010 2236 1011
rect 2342 1009 2348 1010
rect 2198 1004 2204 1005
rect 2207 1007 2213 1008
rect 2055 1002 2061 1003
rect 2207 1003 2208 1007
rect 2212 1003 2213 1007
rect 2342 1005 2343 1009
rect 2347 1005 2348 1009
rect 2494 1009 2500 1010
rect 2342 1004 2348 1005
rect 2350 1007 2357 1008
rect 2207 1002 2213 1003
rect 2350 1003 2351 1007
rect 2356 1003 2357 1007
rect 2494 1005 2495 1009
rect 2499 1005 2500 1009
rect 2494 1004 2500 1005
rect 2505 1004 2507 1012
rect 2646 1009 2652 1010
rect 2646 1005 2647 1009
rect 2651 1005 2652 1009
rect 2646 1004 2652 1005
rect 3190 1005 3196 1006
rect 2350 1002 2357 1003
rect 2503 1003 2509 1004
rect 1926 998 1932 999
rect 2503 999 2504 1003
rect 2508 1002 2509 1003
rect 2654 1003 2661 1004
rect 2654 1002 2655 1003
rect 2508 1000 2655 1002
rect 2508 999 2509 1000
rect 2503 998 2509 999
rect 2654 999 2655 1000
rect 2660 1002 2661 1003
rect 2702 1003 2708 1004
rect 2702 1002 2703 1003
rect 2660 1000 2703 1002
rect 2660 999 2661 1000
rect 2654 998 2661 999
rect 2702 999 2703 1000
rect 2707 999 2708 1003
rect 3190 1001 3191 1005
rect 3195 1001 3196 1005
rect 3190 1000 3196 1001
rect 2702 998 2708 999
rect 326 992 332 993
rect 326 988 327 992
rect 331 988 332 992
rect 326 987 332 988
rect 454 992 460 993
rect 454 988 455 992
rect 459 988 460 992
rect 454 987 460 988
rect 574 992 580 993
rect 574 988 575 992
rect 579 988 580 992
rect 574 987 580 988
rect 694 992 700 993
rect 694 988 695 992
rect 699 988 700 992
rect 694 987 700 988
rect 814 992 820 993
rect 814 988 815 992
rect 819 988 820 992
rect 814 987 820 988
rect 926 992 932 993
rect 926 988 927 992
rect 931 988 932 992
rect 926 987 932 988
rect 1038 992 1044 993
rect 1038 988 1039 992
rect 1043 988 1044 992
rect 1038 987 1044 988
rect 1158 992 1164 993
rect 1158 988 1159 992
rect 1163 988 1164 992
rect 1158 987 1164 988
rect 1670 987 1676 988
rect 110 985 116 986
rect 110 981 111 985
rect 115 981 116 985
rect 110 980 116 981
rect 1630 985 1636 986
rect 1630 981 1631 985
rect 1635 981 1636 985
rect 1670 983 1671 987
rect 1675 983 1676 987
rect 1670 982 1676 983
rect 3190 987 3196 988
rect 3190 983 3191 987
rect 3195 983 3196 987
rect 3190 982 3196 983
rect 1630 980 1636 981
rect 1894 980 1900 981
rect 1894 976 1895 980
rect 1899 976 1900 980
rect 1894 975 1900 976
rect 2046 980 2052 981
rect 2046 976 2047 980
rect 2051 976 2052 980
rect 2046 975 2052 976
rect 2198 980 2204 981
rect 2198 976 2199 980
rect 2203 976 2204 980
rect 2198 975 2204 976
rect 2342 980 2348 981
rect 2342 976 2343 980
rect 2347 976 2348 980
rect 2342 975 2348 976
rect 2494 980 2500 981
rect 2494 976 2495 980
rect 2499 976 2500 980
rect 2494 975 2500 976
rect 2646 980 2652 981
rect 2646 976 2647 980
rect 2651 976 2652 980
rect 2646 975 2652 976
rect 1790 968 1796 969
rect 110 967 116 968
rect 110 963 111 967
rect 115 963 116 967
rect 582 967 589 968
rect 110 962 116 963
rect 326 963 332 964
rect 326 959 327 963
rect 331 959 332 963
rect 326 958 332 959
rect 334 963 341 964
rect 334 959 335 963
rect 340 959 341 963
rect 334 958 341 959
rect 454 963 460 964
rect 454 959 455 963
rect 459 959 460 963
rect 454 958 460 959
rect 462 963 469 964
rect 462 959 463 963
rect 468 959 469 963
rect 462 958 469 959
rect 574 963 580 964
rect 574 959 575 963
rect 579 959 580 963
rect 582 963 583 967
rect 588 963 589 967
rect 702 967 709 968
rect 582 962 589 963
rect 694 963 700 964
rect 574 958 580 959
rect 694 959 695 963
rect 699 959 700 963
rect 702 963 703 967
rect 708 963 709 967
rect 1630 967 1636 968
rect 702 962 709 963
rect 814 963 820 964
rect 694 958 700 959
rect 814 959 815 963
rect 819 959 820 963
rect 814 958 820 959
rect 823 963 829 964
rect 823 959 824 963
rect 828 959 829 963
rect 823 958 829 959
rect 926 963 932 964
rect 926 959 927 963
rect 931 959 932 963
rect 926 958 932 959
rect 935 963 941 964
rect 935 959 936 963
rect 940 962 941 963
rect 950 963 956 964
rect 950 962 951 963
rect 940 960 951 962
rect 940 959 941 960
rect 935 958 941 959
rect 950 959 951 960
rect 955 959 956 963
rect 950 958 956 959
rect 1038 963 1044 964
rect 1038 959 1039 963
rect 1043 959 1044 963
rect 1038 958 1044 959
rect 1047 963 1053 964
rect 1047 959 1048 963
rect 1052 962 1053 963
rect 1070 963 1076 964
rect 1070 962 1071 963
rect 1052 960 1071 962
rect 1052 959 1053 960
rect 1047 958 1053 959
rect 1070 959 1071 960
rect 1075 959 1076 963
rect 1070 958 1076 959
rect 1158 963 1164 964
rect 1158 959 1159 963
rect 1163 959 1164 963
rect 1158 958 1164 959
rect 1166 963 1173 964
rect 1166 959 1167 963
rect 1172 959 1173 963
rect 1630 963 1631 967
rect 1635 963 1636 967
rect 1790 964 1791 968
rect 1795 964 1796 968
rect 1790 963 1796 964
rect 1918 968 1924 969
rect 1918 964 1919 968
rect 1923 964 1924 968
rect 1918 963 1924 964
rect 2070 968 2076 969
rect 2070 964 2071 968
rect 2075 964 2076 968
rect 2070 963 2076 964
rect 2254 968 2260 969
rect 2254 964 2255 968
rect 2259 964 2260 968
rect 2254 963 2260 964
rect 2462 968 2468 969
rect 2462 964 2463 968
rect 2467 964 2468 968
rect 2462 963 2468 964
rect 2694 968 2700 969
rect 2694 964 2695 968
rect 2699 964 2700 968
rect 2694 963 2700 964
rect 2934 968 2940 969
rect 2934 964 2935 968
rect 2939 964 2940 968
rect 2934 963 2940 964
rect 3158 968 3164 969
rect 3158 964 3159 968
rect 3163 964 3164 968
rect 3158 963 3164 964
rect 1630 962 1636 963
rect 1166 958 1173 959
rect 1670 961 1676 962
rect 1670 957 1671 961
rect 1675 957 1676 961
rect 1670 956 1676 957
rect 3190 961 3196 962
rect 3190 957 3191 961
rect 3195 957 3196 961
rect 3190 956 3196 957
rect 2230 947 2236 948
rect 1670 943 1676 944
rect 222 941 228 942
rect 110 937 116 938
rect 110 933 111 937
rect 115 933 116 937
rect 222 937 223 941
rect 227 937 228 941
rect 350 941 356 942
rect 222 936 228 937
rect 231 939 237 940
rect 231 935 232 939
rect 236 938 237 939
rect 258 939 264 940
rect 258 938 259 939
rect 236 936 259 938
rect 236 935 237 936
rect 231 934 237 935
rect 258 935 259 936
rect 263 938 264 939
rect 334 939 340 940
rect 334 938 335 939
rect 263 936 335 938
rect 263 935 264 936
rect 258 934 264 935
rect 334 935 335 936
rect 339 935 340 939
rect 350 937 351 941
rect 355 937 356 941
rect 350 936 356 937
rect 470 941 476 942
rect 470 937 471 941
rect 475 937 476 941
rect 470 936 476 937
rect 590 941 596 942
rect 590 937 591 941
rect 595 937 596 941
rect 590 936 596 937
rect 710 941 716 942
rect 710 937 711 941
rect 715 937 716 941
rect 710 936 716 937
rect 822 941 828 942
rect 822 937 823 941
rect 827 937 828 941
rect 822 936 828 937
rect 942 941 948 942
rect 942 937 943 941
rect 947 937 948 941
rect 942 936 948 937
rect 1062 941 1068 942
rect 1062 937 1063 941
rect 1067 937 1068 941
rect 1670 939 1671 943
rect 1675 939 1676 943
rect 2230 943 2231 947
rect 2235 946 2236 947
rect 2235 944 2267 946
rect 2235 943 2236 944
rect 2230 942 2236 943
rect 2263 943 2269 944
rect 1670 938 1676 939
rect 1790 939 1796 940
rect 1062 936 1068 937
rect 1630 937 1636 938
rect 334 934 340 935
rect 359 935 365 936
rect 359 934 360 935
rect 110 932 116 933
rect 336 932 360 934
rect 359 931 360 932
rect 364 934 365 935
rect 462 935 468 936
rect 462 934 463 935
rect 364 932 463 934
rect 364 931 365 932
rect 359 930 365 931
rect 462 931 463 932
rect 467 934 468 935
rect 479 935 485 936
rect 479 934 480 935
rect 467 932 480 934
rect 467 931 468 932
rect 462 930 468 931
rect 479 931 480 932
rect 484 931 485 935
rect 479 930 485 931
rect 582 935 588 936
rect 582 931 583 935
rect 587 934 588 935
rect 599 935 605 936
rect 599 934 600 935
rect 587 932 600 934
rect 587 931 588 932
rect 582 930 588 931
rect 599 931 600 932
rect 604 931 605 935
rect 599 930 605 931
rect 702 935 708 936
rect 702 931 703 935
rect 707 934 708 935
rect 719 935 725 936
rect 719 934 720 935
rect 707 932 720 934
rect 707 931 708 932
rect 702 930 708 931
rect 719 931 720 932
rect 724 931 725 935
rect 719 930 725 931
rect 830 935 837 936
rect 830 931 831 935
rect 836 934 837 935
rect 950 935 957 936
rect 950 934 951 935
rect 836 932 951 934
rect 836 931 837 932
rect 830 930 837 931
rect 950 931 951 932
rect 956 934 957 935
rect 1070 935 1077 936
rect 1070 934 1071 935
rect 956 932 1071 934
rect 956 931 957 932
rect 950 930 957 931
rect 1070 931 1071 932
rect 1076 931 1077 935
rect 1630 933 1631 937
rect 1635 933 1636 937
rect 1790 935 1791 939
rect 1795 935 1796 939
rect 1790 934 1796 935
rect 1799 939 1808 940
rect 1799 935 1800 939
rect 1807 935 1808 939
rect 1799 934 1808 935
rect 1918 939 1924 940
rect 1918 935 1919 939
rect 1923 935 1924 939
rect 1918 934 1924 935
rect 1926 939 1933 940
rect 1926 935 1927 939
rect 1932 935 1933 939
rect 1926 934 1933 935
rect 2070 939 2076 940
rect 2070 935 2071 939
rect 2075 935 2076 939
rect 2070 934 2076 935
rect 2078 939 2085 940
rect 2078 935 2079 939
rect 2084 935 2085 939
rect 2078 934 2085 935
rect 2254 939 2260 940
rect 2254 935 2255 939
rect 2259 935 2260 939
rect 2263 939 2264 943
rect 2268 939 2269 943
rect 2702 943 2709 944
rect 2263 938 2269 939
rect 2462 939 2468 940
rect 2254 934 2260 935
rect 2462 935 2463 939
rect 2467 935 2468 939
rect 2462 934 2468 935
rect 2470 939 2477 940
rect 2470 935 2471 939
rect 2476 935 2477 939
rect 2470 934 2477 935
rect 2694 939 2700 940
rect 2694 935 2695 939
rect 2699 935 2700 939
rect 2702 939 2703 943
rect 2708 942 2709 943
rect 2830 943 2836 944
rect 2830 942 2831 943
rect 2708 940 2831 942
rect 2708 939 2709 940
rect 2702 938 2709 939
rect 2830 939 2831 940
rect 2835 939 2836 943
rect 2942 943 2949 944
rect 2830 938 2836 939
rect 2934 939 2940 940
rect 2694 934 2700 935
rect 2934 935 2935 939
rect 2939 935 2940 939
rect 2942 939 2943 943
rect 2948 942 2949 943
rect 3006 943 3012 944
rect 3006 942 3007 943
rect 2948 940 3007 942
rect 2948 939 2949 940
rect 2942 938 2949 939
rect 3006 939 3007 940
rect 3011 939 3012 943
rect 3166 943 3173 944
rect 3006 938 3012 939
rect 3158 939 3164 940
rect 2934 934 2940 935
rect 3158 935 3159 939
rect 3163 935 3164 939
rect 3166 939 3167 943
rect 3172 939 3173 943
rect 3166 938 3173 939
rect 3190 943 3196 944
rect 3190 939 3191 943
rect 3195 939 3196 943
rect 3190 938 3196 939
rect 3158 934 3164 935
rect 1630 932 1636 933
rect 1070 930 1077 931
rect 1718 921 1724 922
rect 110 919 116 920
rect 110 915 111 919
rect 115 915 116 919
rect 110 914 116 915
rect 1630 919 1636 920
rect 1630 915 1631 919
rect 1635 915 1636 919
rect 1630 914 1636 915
rect 1670 917 1676 918
rect 1670 913 1671 917
rect 1675 913 1676 917
rect 1718 917 1719 921
rect 1723 917 1724 921
rect 1718 916 1724 917
rect 1870 921 1876 922
rect 1870 917 1871 921
rect 1875 917 1876 921
rect 1870 916 1876 917
rect 2038 921 2044 922
rect 2038 917 2039 921
rect 2043 917 2044 921
rect 2038 916 2044 917
rect 2222 921 2228 922
rect 2222 917 2223 921
rect 2227 917 2228 921
rect 2438 921 2444 922
rect 2222 916 2228 917
rect 2230 919 2237 920
rect 222 912 228 913
rect 222 908 223 912
rect 227 908 228 912
rect 222 907 228 908
rect 350 912 356 913
rect 350 908 351 912
rect 355 908 356 912
rect 350 907 356 908
rect 470 912 476 913
rect 470 908 471 912
rect 475 908 476 912
rect 470 907 476 908
rect 590 912 596 913
rect 590 908 591 912
rect 595 908 596 912
rect 590 907 596 908
rect 710 912 716 913
rect 710 908 711 912
rect 715 908 716 912
rect 710 907 716 908
rect 822 912 828 913
rect 822 908 823 912
rect 827 908 828 912
rect 822 907 828 908
rect 942 912 948 913
rect 942 908 943 912
rect 947 908 948 912
rect 942 907 948 908
rect 1062 912 1068 913
rect 1670 912 1676 913
rect 1727 915 1733 916
rect 1062 908 1063 912
rect 1067 908 1068 912
rect 1727 911 1728 915
rect 1732 914 1733 915
rect 1802 915 1808 916
rect 1802 914 1803 915
rect 1732 912 1803 914
rect 1732 911 1733 912
rect 1727 910 1733 911
rect 1802 911 1803 912
rect 1807 914 1808 915
rect 1879 915 1885 916
rect 1879 914 1880 915
rect 1807 912 1880 914
rect 1807 911 1808 912
rect 1802 910 1808 911
rect 1879 911 1880 912
rect 1884 914 1885 915
rect 1926 915 1932 916
rect 1926 914 1927 915
rect 1884 912 1927 914
rect 1884 911 1885 912
rect 1879 910 1885 911
rect 1926 911 1927 912
rect 1931 914 1932 915
rect 2022 915 2028 916
rect 2022 914 2023 915
rect 1931 912 2023 914
rect 1931 911 1932 912
rect 1926 910 1932 911
rect 2022 911 2023 912
rect 2027 914 2028 915
rect 2047 915 2053 916
rect 2047 914 2048 915
rect 2027 912 2048 914
rect 2027 911 2028 912
rect 2022 910 2028 911
rect 2047 911 2048 912
rect 2052 914 2053 915
rect 2078 915 2084 916
rect 2078 914 2079 915
rect 2052 912 2079 914
rect 2052 911 2053 912
rect 2047 910 2053 911
rect 2078 911 2079 912
rect 2083 911 2084 915
rect 2230 915 2231 919
rect 2236 915 2237 919
rect 2438 917 2439 921
rect 2443 917 2444 921
rect 2670 921 2676 922
rect 2438 916 2444 917
rect 2446 919 2453 920
rect 2230 914 2237 915
rect 2446 915 2447 919
rect 2452 918 2453 919
rect 2470 919 2476 920
rect 2470 918 2471 919
rect 2452 916 2471 918
rect 2452 915 2453 916
rect 2446 914 2453 915
rect 2470 915 2471 916
rect 2475 915 2476 919
rect 2670 917 2671 921
rect 2675 917 2676 921
rect 2910 921 2916 922
rect 2670 916 2676 917
rect 2679 919 2685 920
rect 2470 914 2476 915
rect 2679 915 2680 919
rect 2684 918 2685 919
rect 2702 919 2708 920
rect 2702 918 2703 919
rect 2684 916 2703 918
rect 2684 915 2685 916
rect 2679 914 2685 915
rect 2702 915 2703 916
rect 2707 915 2708 919
rect 2910 917 2911 921
rect 2915 917 2916 921
rect 3158 921 3164 922
rect 2910 916 2916 917
rect 2919 919 2925 920
rect 2702 914 2708 915
rect 2919 915 2920 919
rect 2924 918 2925 919
rect 2942 919 2948 920
rect 2942 918 2943 919
rect 2924 916 2943 918
rect 2924 915 2925 916
rect 2919 914 2925 915
rect 2942 915 2943 916
rect 2947 915 2948 919
rect 3158 917 3159 921
rect 3163 917 3164 921
rect 3158 916 3164 917
rect 3166 919 3173 920
rect 2942 914 2948 915
rect 3166 915 3167 919
rect 3172 915 3173 919
rect 3166 914 3173 915
rect 3190 917 3196 918
rect 3190 913 3191 917
rect 3195 913 3196 917
rect 3190 912 3196 913
rect 2078 910 2084 911
rect 1062 907 1068 908
rect 1670 899 1676 900
rect 1670 895 1671 899
rect 1675 895 1676 899
rect 1670 894 1676 895
rect 3190 899 3196 900
rect 3190 895 3191 899
rect 3195 895 3196 899
rect 3190 894 3196 895
rect 1718 892 1724 893
rect 134 888 140 889
rect 134 884 135 888
rect 139 884 140 888
rect 134 883 140 884
rect 246 888 252 889
rect 246 884 247 888
rect 251 884 252 888
rect 246 883 252 884
rect 382 888 388 889
rect 382 884 383 888
rect 387 884 388 888
rect 382 883 388 884
rect 534 888 540 889
rect 534 884 535 888
rect 539 884 540 888
rect 534 883 540 884
rect 710 888 716 889
rect 710 884 711 888
rect 715 884 716 888
rect 710 883 716 884
rect 918 888 924 889
rect 918 884 919 888
rect 923 884 924 888
rect 918 883 924 884
rect 1142 888 1148 889
rect 1142 884 1143 888
rect 1147 884 1148 888
rect 1142 883 1148 884
rect 1382 888 1388 889
rect 1382 884 1383 888
rect 1387 884 1388 888
rect 1382 883 1388 884
rect 1598 888 1604 889
rect 1598 884 1599 888
rect 1603 884 1604 888
rect 1718 888 1719 892
rect 1723 888 1724 892
rect 1718 887 1724 888
rect 1870 892 1876 893
rect 1870 888 1871 892
rect 1875 888 1876 892
rect 1870 887 1876 888
rect 2038 892 2044 893
rect 2038 888 2039 892
rect 2043 888 2044 892
rect 2038 887 2044 888
rect 2222 892 2228 893
rect 2222 888 2223 892
rect 2227 888 2228 892
rect 2222 887 2228 888
rect 2438 892 2444 893
rect 2438 888 2439 892
rect 2443 888 2444 892
rect 2438 887 2444 888
rect 2670 892 2676 893
rect 2670 888 2671 892
rect 2675 888 2676 892
rect 2670 887 2676 888
rect 2910 892 2916 893
rect 2910 888 2911 892
rect 2915 888 2916 892
rect 2910 887 2916 888
rect 3158 892 3164 893
rect 3158 888 3159 892
rect 3163 888 3164 892
rect 3158 887 3164 888
rect 1598 883 1604 884
rect 110 881 116 882
rect 110 877 111 881
rect 115 877 116 881
rect 110 876 116 877
rect 1630 881 1636 882
rect 1630 877 1631 881
rect 1635 877 1636 881
rect 1630 876 1636 877
rect 1694 880 1700 881
rect 1694 876 1695 880
rect 1699 876 1700 880
rect 1694 875 1700 876
rect 2014 880 2020 881
rect 2014 876 2015 880
rect 2019 876 2020 880
rect 2014 875 2020 876
rect 2366 880 2372 881
rect 2366 876 2367 880
rect 2371 876 2372 880
rect 2366 875 2372 876
rect 2726 880 2732 881
rect 2726 876 2727 880
rect 2731 876 2732 880
rect 2726 875 2732 876
rect 3086 880 3092 881
rect 3086 876 3087 880
rect 3091 876 3092 880
rect 3086 875 3092 876
rect 1670 873 1676 874
rect 1670 869 1671 873
rect 1675 869 1676 873
rect 1670 868 1676 869
rect 3190 873 3196 874
rect 3190 869 3191 873
rect 3195 869 3196 873
rect 3190 868 3196 869
rect 110 863 116 864
rect 110 859 111 863
rect 115 859 116 863
rect 255 863 264 864
rect 110 858 116 859
rect 134 859 140 860
rect 134 855 135 859
rect 139 855 140 859
rect 134 854 140 855
rect 143 859 149 860
rect 143 855 144 859
rect 148 855 149 859
rect 143 854 149 855
rect 246 859 252 860
rect 246 855 247 859
rect 251 855 252 859
rect 255 859 256 863
rect 263 859 264 863
rect 1630 863 1636 864
rect 255 858 264 859
rect 382 859 388 860
rect 246 854 252 855
rect 382 855 383 859
rect 387 855 388 859
rect 382 854 388 855
rect 391 859 397 860
rect 391 855 392 859
rect 396 855 397 859
rect 391 854 397 855
rect 534 859 540 860
rect 534 855 535 859
rect 539 855 540 859
rect 534 854 540 855
rect 543 859 549 860
rect 543 855 544 859
rect 548 855 549 859
rect 543 854 549 855
rect 710 859 716 860
rect 710 855 711 859
rect 715 855 716 859
rect 710 854 716 855
rect 718 859 725 860
rect 718 855 719 859
rect 724 855 725 859
rect 718 854 725 855
rect 918 859 924 860
rect 918 855 919 859
rect 923 855 924 859
rect 918 854 924 855
rect 926 859 933 860
rect 926 855 927 859
rect 932 855 933 859
rect 926 854 933 855
rect 1142 859 1148 860
rect 1142 855 1143 859
rect 1147 855 1148 859
rect 1142 854 1148 855
rect 1151 859 1160 860
rect 1151 855 1152 859
rect 1159 858 1160 859
rect 1166 859 1172 860
rect 1166 858 1167 859
rect 1159 856 1167 858
rect 1159 855 1160 856
rect 1151 854 1160 855
rect 1166 855 1167 856
rect 1171 855 1172 859
rect 1166 854 1172 855
rect 1382 859 1388 860
rect 1382 855 1383 859
rect 1387 855 1388 859
rect 1382 854 1388 855
rect 1391 859 1400 860
rect 1391 855 1392 859
rect 1399 855 1400 859
rect 1391 854 1400 855
rect 1598 859 1604 860
rect 1598 855 1599 859
rect 1603 855 1604 859
rect 1598 854 1604 855
rect 1607 859 1613 860
rect 1607 855 1608 859
rect 1612 855 1613 859
rect 1630 859 1631 863
rect 1635 859 1636 863
rect 1630 858 1636 859
rect 1639 860 1707 862
rect 1607 854 1613 855
rect 1639 854 1641 860
rect 1705 856 1707 860
rect 134 845 140 846
rect 110 841 116 842
rect 110 837 111 841
rect 115 837 116 841
rect 134 841 135 845
rect 139 841 140 845
rect 144 844 146 854
rect 258 851 264 852
rect 258 847 259 851
rect 263 850 264 851
rect 392 850 394 854
rect 544 850 546 854
rect 1609 852 1641 854
rect 1670 855 1676 856
rect 582 851 588 852
rect 582 850 583 851
rect 263 848 583 850
rect 263 847 264 848
rect 258 846 264 847
rect 134 840 140 841
rect 143 843 149 844
rect 143 839 144 843
rect 148 842 149 843
rect 260 842 262 846
rect 148 840 262 842
rect 302 845 308 846
rect 302 841 303 845
rect 307 841 308 845
rect 312 844 314 848
rect 502 845 508 846
rect 302 840 308 841
rect 311 843 317 844
rect 148 839 149 840
rect 143 838 149 839
rect 311 839 312 843
rect 316 839 317 843
rect 502 841 503 845
rect 507 841 508 845
rect 512 844 514 848
rect 582 847 583 848
rect 587 847 588 851
rect 582 846 588 847
rect 694 845 700 846
rect 502 840 508 841
rect 511 843 517 844
rect 311 838 317 839
rect 511 839 512 843
rect 516 839 517 843
rect 694 841 695 845
rect 699 841 700 845
rect 694 840 700 841
rect 878 845 884 846
rect 878 841 879 845
rect 883 841 884 845
rect 878 840 884 841
rect 1046 845 1052 846
rect 1046 841 1047 845
rect 1051 841 1052 845
rect 1046 840 1052 841
rect 1198 845 1204 846
rect 1198 841 1199 845
rect 1203 841 1204 845
rect 1198 840 1204 841
rect 1334 845 1340 846
rect 1334 841 1335 845
rect 1339 841 1340 845
rect 1334 840 1340 841
rect 1470 845 1476 846
rect 1470 841 1471 845
rect 1475 841 1476 845
rect 1470 840 1476 841
rect 1598 845 1604 846
rect 1598 841 1599 845
rect 1603 841 1604 845
rect 1609 844 1611 852
rect 1670 851 1671 855
rect 1675 851 1676 855
rect 1703 855 1709 856
rect 1670 850 1676 851
rect 1694 851 1700 852
rect 1694 847 1695 851
rect 1699 847 1700 851
rect 1703 851 1704 855
rect 1708 851 1709 855
rect 2022 855 2029 856
rect 1703 850 1709 851
rect 2014 851 2020 852
rect 1694 846 1700 847
rect 2014 847 2015 851
rect 2019 847 2020 851
rect 2022 851 2023 855
rect 2028 851 2029 855
rect 2375 855 2381 856
rect 2022 850 2029 851
rect 2366 851 2372 852
rect 2014 846 2020 847
rect 2366 847 2367 851
rect 2371 847 2372 851
rect 2375 851 2376 855
rect 2380 854 2381 855
rect 2446 855 2452 856
rect 2446 854 2447 855
rect 2380 852 2447 854
rect 2380 851 2381 852
rect 2375 850 2381 851
rect 2446 851 2447 852
rect 2451 851 2452 855
rect 3095 855 3101 856
rect 2446 850 2452 851
rect 2726 851 2732 852
rect 2366 846 2372 847
rect 2726 847 2727 851
rect 2731 847 2732 851
rect 2726 846 2732 847
rect 2735 851 2744 852
rect 2735 847 2736 851
rect 2743 847 2744 851
rect 2735 846 2744 847
rect 3086 851 3092 852
rect 3086 847 3087 851
rect 3091 847 3092 851
rect 3095 851 3096 855
rect 3100 854 3101 855
rect 3118 855 3124 856
rect 3118 854 3119 855
rect 3100 852 3119 854
rect 3100 851 3101 852
rect 3095 850 3101 851
rect 3118 851 3119 852
rect 3123 854 3124 855
rect 3166 855 3172 856
rect 3166 854 3167 855
rect 3123 852 3167 854
rect 3123 851 3124 852
rect 3118 850 3124 851
rect 3166 851 3167 852
rect 3171 851 3172 855
rect 3166 850 3172 851
rect 3190 855 3196 856
rect 3190 851 3191 855
rect 3195 851 3196 855
rect 3190 850 3196 851
rect 3086 846 3092 847
rect 1598 840 1604 841
rect 1607 843 1613 844
rect 511 838 517 839
rect 686 839 692 840
rect 110 836 116 837
rect 686 835 687 839
rect 691 838 692 839
rect 703 839 709 840
rect 703 838 704 839
rect 691 836 704 838
rect 691 835 692 836
rect 686 834 692 835
rect 703 835 704 836
rect 708 838 709 839
rect 718 839 724 840
rect 718 838 719 839
rect 708 836 719 838
rect 708 835 709 836
rect 703 834 709 835
rect 718 835 719 836
rect 723 835 724 839
rect 718 834 724 835
rect 886 839 893 840
rect 886 835 887 839
rect 892 838 893 839
rect 926 839 932 840
rect 926 838 927 839
rect 892 836 927 838
rect 892 835 893 836
rect 886 834 893 835
rect 926 835 927 836
rect 931 835 932 839
rect 926 834 932 835
rect 1055 839 1061 840
rect 1055 835 1056 839
rect 1060 838 1061 839
rect 1070 839 1076 840
rect 1070 838 1071 839
rect 1060 836 1071 838
rect 1060 835 1061 836
rect 1055 834 1061 835
rect 1070 835 1071 836
rect 1075 838 1076 839
rect 1154 839 1160 840
rect 1154 838 1155 839
rect 1075 836 1155 838
rect 1075 835 1076 836
rect 1070 834 1076 835
rect 1154 835 1155 836
rect 1159 838 1160 839
rect 1207 839 1213 840
rect 1207 838 1208 839
rect 1159 836 1208 838
rect 1159 835 1160 836
rect 1154 834 1160 835
rect 1207 835 1208 836
rect 1212 838 1213 839
rect 1343 839 1349 840
rect 1343 838 1344 839
rect 1212 836 1344 838
rect 1212 835 1213 836
rect 1207 834 1213 835
rect 1343 835 1344 836
rect 1348 838 1349 839
rect 1394 839 1400 840
rect 1394 838 1395 839
rect 1348 836 1395 838
rect 1348 835 1349 836
rect 1343 834 1349 835
rect 1394 835 1395 836
rect 1399 838 1400 839
rect 1479 839 1485 840
rect 1479 838 1480 839
rect 1399 836 1480 838
rect 1399 835 1400 836
rect 1394 834 1400 835
rect 1479 835 1480 836
rect 1484 838 1485 839
rect 1526 839 1532 840
rect 1526 838 1527 839
rect 1484 836 1527 838
rect 1484 835 1485 836
rect 1479 834 1485 835
rect 1526 835 1527 836
rect 1531 838 1532 839
rect 1607 839 1608 843
rect 1612 839 1613 843
rect 1607 838 1613 839
rect 1630 841 1636 842
rect 1531 836 1611 838
rect 1630 837 1631 841
rect 1635 837 1636 841
rect 1630 836 1636 837
rect 1531 835 1532 836
rect 1526 834 1532 835
rect 2278 829 2284 830
rect 1670 825 1676 826
rect 110 823 116 824
rect 110 819 111 823
rect 115 819 116 823
rect 110 818 116 819
rect 1630 823 1636 824
rect 1630 819 1631 823
rect 1635 819 1636 823
rect 1670 821 1671 825
rect 1675 821 1676 825
rect 2278 825 2279 829
rect 2283 825 2284 829
rect 2278 824 2284 825
rect 2438 829 2444 830
rect 2438 825 2439 829
rect 2443 825 2444 829
rect 2582 829 2588 830
rect 2438 824 2444 825
rect 2446 827 2453 828
rect 1670 820 1676 821
rect 2230 823 2236 824
rect 1630 818 1636 819
rect 2230 819 2231 823
rect 2235 822 2236 823
rect 2287 823 2293 824
rect 2287 822 2288 823
rect 2235 820 2288 822
rect 2235 819 2236 820
rect 2230 818 2236 819
rect 2287 819 2288 820
rect 2292 822 2293 823
rect 2306 823 2312 824
rect 2306 822 2307 823
rect 2292 820 2307 822
rect 2292 819 2293 820
rect 2287 818 2293 819
rect 2306 819 2307 820
rect 2311 819 2312 823
rect 2446 823 2447 827
rect 2452 826 2453 827
rect 2458 827 2464 828
rect 2458 826 2459 827
rect 2452 824 2459 826
rect 2452 823 2453 824
rect 2446 822 2453 823
rect 2458 823 2459 824
rect 2463 823 2464 827
rect 2582 825 2583 829
rect 2587 825 2588 829
rect 2582 824 2588 825
rect 2718 829 2724 830
rect 2718 825 2719 829
rect 2723 825 2724 829
rect 2846 829 2852 830
rect 2718 824 2724 825
rect 2727 825 2733 826
rect 2458 822 2464 823
rect 2591 823 2597 824
rect 2306 818 2312 819
rect 2591 819 2592 823
rect 2596 822 2597 823
rect 2622 823 2628 824
rect 2622 822 2623 823
rect 2596 820 2623 822
rect 2596 819 2597 820
rect 2591 818 2597 819
rect 2622 819 2623 820
rect 2627 819 2628 823
rect 2727 821 2728 825
rect 2732 824 2733 825
rect 2846 825 2847 829
rect 2851 825 2852 829
rect 2846 824 2852 825
rect 2974 829 2980 830
rect 2974 825 2975 829
rect 2979 825 2980 829
rect 2974 824 2980 825
rect 3110 829 3116 830
rect 3110 825 3111 829
rect 3115 825 3116 829
rect 3110 824 3116 825
rect 3118 827 3125 828
rect 2732 823 2744 824
rect 2732 822 2739 823
rect 2732 821 2733 822
rect 2727 820 2733 821
rect 2622 818 2628 819
rect 2738 819 2739 822
rect 2743 822 2744 823
rect 2798 823 2804 824
rect 2798 822 2799 823
rect 2743 820 2799 822
rect 2743 819 2744 820
rect 2738 818 2744 819
rect 2798 819 2799 820
rect 2803 822 2804 823
rect 2855 823 2861 824
rect 2855 822 2856 823
rect 2803 820 2856 822
rect 2803 819 2804 820
rect 2798 818 2804 819
rect 2855 819 2856 820
rect 2860 819 2861 823
rect 2855 818 2861 819
rect 2930 823 2936 824
rect 2930 819 2931 823
rect 2935 822 2936 823
rect 2983 823 2989 824
rect 2983 822 2984 823
rect 2935 820 2984 822
rect 2935 819 2936 820
rect 2930 818 2936 819
rect 2983 819 2984 820
rect 2988 822 2989 823
rect 3054 823 3060 824
rect 3054 822 3055 823
rect 2988 820 3055 822
rect 2988 819 2989 820
rect 2983 818 2989 819
rect 3054 819 3055 820
rect 3059 822 3060 823
rect 3118 823 3119 827
rect 3124 823 3125 827
rect 3118 822 3125 823
rect 3190 825 3196 826
rect 3059 820 3122 822
rect 3190 821 3191 825
rect 3195 821 3196 825
rect 3190 820 3196 821
rect 3059 819 3060 820
rect 3054 818 3060 819
rect 134 816 140 817
rect 134 812 135 816
rect 139 812 140 816
rect 134 811 140 812
rect 302 816 308 817
rect 302 812 303 816
rect 307 812 308 816
rect 302 811 308 812
rect 502 816 508 817
rect 502 812 503 816
rect 507 812 508 816
rect 502 811 508 812
rect 694 816 700 817
rect 694 812 695 816
rect 699 812 700 816
rect 694 811 700 812
rect 878 816 884 817
rect 878 812 879 816
rect 883 812 884 816
rect 878 811 884 812
rect 1046 816 1052 817
rect 1046 812 1047 816
rect 1051 812 1052 816
rect 1046 811 1052 812
rect 1198 816 1204 817
rect 1198 812 1199 816
rect 1203 812 1204 816
rect 1198 811 1204 812
rect 1334 816 1340 817
rect 1334 812 1335 816
rect 1339 812 1340 816
rect 1334 811 1340 812
rect 1470 816 1476 817
rect 1470 812 1471 816
rect 1475 812 1476 816
rect 1470 811 1476 812
rect 1598 816 1604 817
rect 1598 812 1599 816
rect 1603 812 1604 816
rect 1598 811 1604 812
rect 1670 807 1676 808
rect 1670 803 1671 807
rect 1675 803 1676 807
rect 1670 802 1676 803
rect 3190 807 3196 808
rect 3190 803 3191 807
rect 3195 803 3196 807
rect 3190 802 3196 803
rect 2278 800 2284 801
rect 2278 796 2279 800
rect 2283 796 2284 800
rect 2278 795 2284 796
rect 2438 800 2444 801
rect 2438 796 2439 800
rect 2443 796 2444 800
rect 2438 795 2444 796
rect 2582 800 2588 801
rect 2582 796 2583 800
rect 2587 796 2588 800
rect 2582 795 2588 796
rect 2718 800 2724 801
rect 2718 796 2719 800
rect 2723 796 2724 800
rect 2718 795 2724 796
rect 2846 800 2852 801
rect 2846 796 2847 800
rect 2851 796 2852 800
rect 2846 795 2852 796
rect 2974 800 2980 801
rect 2974 796 2975 800
rect 2979 796 2980 800
rect 2974 795 2980 796
rect 3110 800 3116 801
rect 3110 796 3111 800
rect 3115 796 3116 800
rect 3110 795 3116 796
rect 678 788 684 789
rect 678 784 679 788
rect 683 784 684 788
rect 678 783 684 784
rect 806 788 812 789
rect 806 784 807 788
rect 811 784 812 788
rect 806 783 812 784
rect 926 788 932 789
rect 926 784 927 788
rect 931 784 932 788
rect 926 783 932 784
rect 1046 788 1052 789
rect 1046 784 1047 788
rect 1051 784 1052 788
rect 1046 783 1052 784
rect 1166 788 1172 789
rect 1166 784 1167 788
rect 1171 784 1172 788
rect 1166 783 1172 784
rect 1278 788 1284 789
rect 1278 784 1279 788
rect 1283 784 1284 788
rect 1278 783 1284 784
rect 1398 788 1404 789
rect 1398 784 1399 788
rect 1403 784 1404 788
rect 1398 783 1404 784
rect 1518 788 1524 789
rect 1518 784 1519 788
rect 1523 784 1524 788
rect 1518 783 1524 784
rect 2198 784 2204 785
rect 110 781 116 782
rect 110 777 111 781
rect 115 777 116 781
rect 110 776 116 777
rect 1630 781 1636 782
rect 1630 777 1631 781
rect 1635 777 1636 781
rect 2198 780 2199 784
rect 2203 780 2204 784
rect 2198 779 2204 780
rect 2358 784 2364 785
rect 2358 780 2359 784
rect 2363 780 2364 784
rect 2358 779 2364 780
rect 2510 784 2516 785
rect 2510 780 2511 784
rect 2515 780 2516 784
rect 2510 779 2516 780
rect 2654 784 2660 785
rect 2654 780 2655 784
rect 2659 780 2660 784
rect 2654 779 2660 780
rect 2790 784 2796 785
rect 2790 780 2791 784
rect 2795 780 2796 784
rect 2790 779 2796 780
rect 2918 784 2924 785
rect 2918 780 2919 784
rect 2923 780 2924 784
rect 2918 779 2924 780
rect 3046 784 3052 785
rect 3046 780 3047 784
rect 3051 780 3052 784
rect 3046 779 3052 780
rect 3158 784 3164 785
rect 3158 780 3159 784
rect 3163 780 3164 784
rect 3158 779 3164 780
rect 1630 776 1636 777
rect 1670 777 1676 778
rect 1670 773 1671 777
rect 1675 773 1676 777
rect 1670 772 1676 773
rect 3190 777 3196 778
rect 3190 773 3191 777
rect 3195 773 3196 777
rect 3190 772 3196 773
rect 1422 767 1428 768
rect 1422 766 1423 767
rect 1412 764 1423 766
rect 110 763 116 764
rect 110 759 111 763
rect 115 759 116 763
rect 1407 763 1414 764
rect 110 758 116 759
rect 678 759 684 760
rect 678 755 679 759
rect 683 755 684 759
rect 678 754 684 755
rect 686 759 693 760
rect 686 755 687 759
rect 692 755 693 759
rect 686 754 693 755
rect 806 759 812 760
rect 806 755 807 759
rect 811 755 812 759
rect 806 754 812 755
rect 814 759 821 760
rect 814 755 815 759
rect 820 755 821 759
rect 814 754 821 755
rect 926 759 932 760
rect 926 755 927 759
rect 931 755 932 759
rect 926 754 932 755
rect 934 759 941 760
rect 934 755 935 759
rect 940 755 941 759
rect 934 754 941 755
rect 1046 759 1052 760
rect 1046 755 1047 759
rect 1051 755 1052 759
rect 1046 754 1052 755
rect 1055 759 1064 760
rect 1055 755 1056 759
rect 1063 755 1064 759
rect 1055 754 1064 755
rect 1166 759 1172 760
rect 1166 755 1167 759
rect 1171 755 1172 759
rect 1166 754 1172 755
rect 1175 759 1181 760
rect 1175 755 1176 759
rect 1180 758 1181 759
rect 1190 759 1196 760
rect 1190 758 1191 759
rect 1180 756 1191 758
rect 1180 755 1181 756
rect 1175 754 1181 755
rect 1190 755 1191 756
rect 1195 755 1196 759
rect 1190 754 1196 755
rect 1278 759 1284 760
rect 1278 755 1279 759
rect 1283 755 1284 759
rect 1278 754 1284 755
rect 1287 759 1293 760
rect 1287 755 1288 759
rect 1292 758 1293 759
rect 1302 759 1308 760
rect 1302 758 1303 759
rect 1292 756 1303 758
rect 1292 755 1293 756
rect 1287 754 1293 755
rect 1302 755 1303 756
rect 1307 755 1308 759
rect 1302 754 1308 755
rect 1398 759 1404 760
rect 1398 755 1399 759
rect 1403 755 1404 759
rect 1407 759 1408 763
rect 1412 760 1414 763
rect 1422 763 1423 764
rect 1427 766 1428 767
rect 1427 764 1530 766
rect 1427 763 1428 764
rect 1422 762 1428 763
rect 1526 763 1533 764
rect 1412 759 1413 760
rect 1407 758 1413 759
rect 1518 759 1524 760
rect 1398 754 1404 755
rect 1518 755 1519 759
rect 1523 755 1524 759
rect 1526 759 1527 763
rect 1532 759 1533 763
rect 1526 758 1533 759
rect 1630 763 1636 764
rect 1630 759 1631 763
rect 1635 759 1636 763
rect 1630 758 1636 759
rect 1670 759 1676 760
rect 1518 754 1524 755
rect 1670 755 1671 759
rect 1675 755 1676 759
rect 2367 759 2373 760
rect 1670 754 1676 755
rect 2198 755 2204 756
rect 614 751 620 752
rect 614 747 615 751
rect 619 750 620 751
rect 689 750 691 754
rect 2198 751 2199 755
rect 2203 751 2204 755
rect 2198 750 2204 751
rect 2207 755 2213 756
rect 2207 751 2208 755
rect 2212 751 2213 755
rect 2207 750 2213 751
rect 2358 755 2364 756
rect 2358 751 2359 755
rect 2363 751 2364 755
rect 2367 755 2368 759
rect 2372 758 2373 759
rect 2458 759 2464 760
rect 2458 758 2459 759
rect 2372 756 2459 758
rect 2372 755 2373 756
rect 2367 754 2373 755
rect 2458 755 2459 756
rect 2463 755 2464 759
rect 2519 759 2525 760
rect 2458 754 2464 755
rect 2510 755 2516 756
rect 2358 750 2364 751
rect 2510 751 2511 755
rect 2515 751 2516 755
rect 2519 755 2520 759
rect 2524 758 2525 759
rect 2622 759 2628 760
rect 2622 758 2623 759
rect 2524 756 2623 758
rect 2524 755 2525 756
rect 2519 754 2525 755
rect 2622 755 2623 756
rect 2627 755 2628 759
rect 2927 759 2936 760
rect 2622 754 2628 755
rect 2654 755 2660 756
rect 2510 750 2516 751
rect 2654 751 2655 755
rect 2659 751 2660 755
rect 2654 750 2660 751
rect 2663 755 2669 756
rect 2663 751 2664 755
rect 2668 754 2669 755
rect 2766 755 2772 756
rect 2766 754 2767 755
rect 2668 752 2767 754
rect 2668 751 2669 752
rect 2663 750 2669 751
rect 2766 751 2767 752
rect 2771 751 2772 755
rect 2766 750 2772 751
rect 2790 755 2796 756
rect 2790 751 2791 755
rect 2795 751 2796 755
rect 2790 750 2796 751
rect 2798 755 2805 756
rect 2798 751 2799 755
rect 2804 751 2805 755
rect 2798 750 2805 751
rect 2918 755 2924 756
rect 2918 751 2919 755
rect 2923 751 2924 755
rect 2927 755 2928 759
rect 2935 755 2936 759
rect 3054 759 3061 760
rect 2927 754 2936 755
rect 3046 755 3052 756
rect 2918 750 2924 751
rect 3046 751 3047 755
rect 3051 751 3052 755
rect 3054 755 3055 759
rect 3060 755 3061 759
rect 3190 759 3196 760
rect 3054 754 3061 755
rect 3158 755 3164 756
rect 3046 750 3052 751
rect 3158 751 3159 755
rect 3163 751 3164 755
rect 3158 750 3164 751
rect 3166 755 3173 756
rect 3166 751 3167 755
rect 3172 751 3173 755
rect 3190 755 3191 759
rect 3195 755 3196 759
rect 3190 754 3196 755
rect 3166 750 3173 751
rect 619 748 691 750
rect 619 747 620 748
rect 614 746 620 747
rect 2158 747 2164 748
rect 2158 743 2159 747
rect 2163 746 2164 747
rect 2209 746 2211 750
rect 2163 744 2211 746
rect 2163 743 2164 744
rect 2158 742 2164 743
rect 574 741 580 742
rect 110 737 116 738
rect 110 733 111 737
rect 115 733 116 737
rect 574 737 575 741
rect 579 737 580 741
rect 574 736 580 737
rect 702 741 708 742
rect 702 737 703 741
rect 707 737 708 741
rect 702 736 708 737
rect 830 741 836 742
rect 830 737 831 741
rect 835 737 836 741
rect 830 736 836 737
rect 950 741 956 742
rect 950 737 951 741
rect 955 737 956 741
rect 950 736 956 737
rect 1070 741 1076 742
rect 1070 737 1071 741
rect 1075 737 1076 741
rect 1070 736 1076 737
rect 1182 741 1188 742
rect 1182 737 1183 741
rect 1187 737 1188 741
rect 1182 736 1188 737
rect 1294 741 1300 742
rect 1294 737 1295 741
rect 1299 737 1300 741
rect 1294 736 1300 737
rect 1414 741 1420 742
rect 1414 737 1415 741
rect 1419 737 1420 741
rect 2126 741 2132 742
rect 1414 736 1420 737
rect 1422 739 1429 740
rect 110 732 116 733
rect 582 735 589 736
rect 582 731 583 735
rect 588 734 589 735
rect 614 735 620 736
rect 614 734 615 735
rect 588 732 615 734
rect 588 731 589 732
rect 582 730 589 731
rect 614 731 615 732
rect 619 731 620 735
rect 614 730 620 731
rect 711 735 717 736
rect 711 731 712 735
rect 716 734 717 735
rect 814 735 820 736
rect 814 734 815 735
rect 716 732 815 734
rect 716 731 717 732
rect 711 730 717 731
rect 814 731 815 732
rect 819 734 820 735
rect 839 735 845 736
rect 839 734 840 735
rect 819 732 840 734
rect 819 731 820 732
rect 814 730 820 731
rect 839 731 840 732
rect 844 734 845 735
rect 854 735 860 736
rect 854 734 855 735
rect 844 732 855 734
rect 844 731 845 732
rect 839 730 845 731
rect 854 731 855 732
rect 859 734 860 735
rect 886 735 892 736
rect 886 734 887 735
rect 859 732 887 734
rect 859 731 860 732
rect 854 730 860 731
rect 886 731 887 732
rect 891 734 892 735
rect 934 735 940 736
rect 934 734 935 735
rect 891 732 935 734
rect 891 731 892 732
rect 886 730 892 731
rect 934 731 935 732
rect 939 734 940 735
rect 959 735 965 736
rect 959 734 960 735
rect 939 732 960 734
rect 939 731 940 732
rect 934 730 940 731
rect 959 731 960 732
rect 964 731 965 735
rect 959 730 965 731
rect 1058 735 1064 736
rect 1058 731 1059 735
rect 1063 734 1064 735
rect 1079 735 1085 736
rect 1079 734 1080 735
rect 1063 732 1080 734
rect 1063 731 1064 732
rect 1058 730 1064 731
rect 1079 731 1080 732
rect 1084 734 1085 735
rect 1190 735 1197 736
rect 1190 734 1191 735
rect 1084 732 1191 734
rect 1084 731 1085 732
rect 1079 730 1085 731
rect 1190 731 1191 732
rect 1196 734 1197 735
rect 1302 735 1309 736
rect 1302 734 1303 735
rect 1196 732 1303 734
rect 1196 731 1197 732
rect 1190 730 1197 731
rect 1302 731 1303 732
rect 1308 734 1309 735
rect 1318 735 1324 736
rect 1318 734 1319 735
rect 1308 732 1319 734
rect 1308 731 1309 732
rect 1302 730 1309 731
rect 1318 731 1319 732
rect 1323 734 1324 735
rect 1422 735 1423 739
rect 1428 735 1429 739
rect 1422 734 1429 735
rect 1630 737 1636 738
rect 1323 732 1426 734
rect 1630 733 1631 737
rect 1635 733 1636 737
rect 1630 732 1636 733
rect 1670 737 1676 738
rect 1670 733 1671 737
rect 1675 733 1676 737
rect 2126 737 2127 741
rect 2131 737 2132 741
rect 2126 736 2132 737
rect 2286 741 2292 742
rect 2286 737 2287 741
rect 2291 737 2292 741
rect 2286 736 2292 737
rect 2446 741 2452 742
rect 2446 737 2447 741
rect 2451 737 2452 741
rect 2446 736 2452 737
rect 2598 741 2604 742
rect 2598 737 2599 741
rect 2603 737 2604 741
rect 2598 736 2604 737
rect 2758 741 2764 742
rect 2758 737 2759 741
rect 2763 737 2764 741
rect 2758 736 2764 737
rect 2918 741 2924 742
rect 2918 737 2919 741
rect 2923 737 2924 741
rect 2918 736 2924 737
rect 2927 739 2936 740
rect 1670 732 1676 733
rect 2135 735 2141 736
rect 1323 731 1324 732
rect 1318 730 1324 731
rect 2135 731 2136 735
rect 2140 734 2141 735
rect 2158 735 2164 736
rect 2158 734 2159 735
rect 2140 732 2159 734
rect 2140 731 2141 732
rect 2135 730 2141 731
rect 2158 731 2159 732
rect 2163 731 2164 735
rect 2158 730 2164 731
rect 2295 735 2301 736
rect 2295 731 2296 735
rect 2300 734 2301 735
rect 2306 735 2312 736
rect 2306 734 2307 735
rect 2300 732 2307 734
rect 2300 731 2301 732
rect 2295 730 2301 731
rect 2306 731 2307 732
rect 2311 731 2312 735
rect 2306 730 2312 731
rect 2455 735 2464 736
rect 2455 731 2456 735
rect 2463 731 2464 735
rect 2455 730 2464 731
rect 2607 735 2613 736
rect 2607 731 2608 735
rect 2612 734 2613 735
rect 2622 735 2628 736
rect 2622 734 2623 735
rect 2612 732 2623 734
rect 2612 731 2613 732
rect 2607 730 2613 731
rect 2622 731 2623 732
rect 2627 731 2628 735
rect 2622 730 2628 731
rect 2766 735 2773 736
rect 2766 731 2767 735
rect 2772 734 2773 735
rect 2798 735 2804 736
rect 2798 734 2799 735
rect 2772 732 2799 734
rect 2772 731 2773 732
rect 2766 730 2773 731
rect 2798 731 2799 732
rect 2803 731 2804 735
rect 2927 735 2928 739
rect 2935 735 2936 739
rect 2927 734 2936 735
rect 3190 737 3196 738
rect 3190 733 3191 737
rect 3195 733 3196 737
rect 3190 732 3196 733
rect 2798 730 2804 731
rect 110 719 116 720
rect 110 715 111 719
rect 115 715 116 719
rect 110 714 116 715
rect 1630 719 1636 720
rect 1630 715 1631 719
rect 1635 715 1636 719
rect 1630 714 1636 715
rect 1670 719 1676 720
rect 1670 715 1671 719
rect 1675 715 1676 719
rect 1670 714 1676 715
rect 3190 719 3196 720
rect 3190 715 3191 719
rect 3195 715 3196 719
rect 3190 714 3196 715
rect 574 712 580 713
rect 574 708 575 712
rect 579 708 580 712
rect 574 707 580 708
rect 702 712 708 713
rect 702 708 703 712
rect 707 708 708 712
rect 702 707 708 708
rect 830 712 836 713
rect 830 708 831 712
rect 835 708 836 712
rect 830 707 836 708
rect 950 712 956 713
rect 950 708 951 712
rect 955 708 956 712
rect 950 707 956 708
rect 1070 712 1076 713
rect 1070 708 1071 712
rect 1075 708 1076 712
rect 1070 707 1076 708
rect 1182 712 1188 713
rect 1182 708 1183 712
rect 1187 708 1188 712
rect 1182 707 1188 708
rect 1294 712 1300 713
rect 1294 708 1295 712
rect 1299 708 1300 712
rect 1294 707 1300 708
rect 1414 712 1420 713
rect 1414 708 1415 712
rect 1419 708 1420 712
rect 1414 707 1420 708
rect 2126 712 2132 713
rect 2126 708 2127 712
rect 2131 708 2132 712
rect 2126 707 2132 708
rect 2286 712 2292 713
rect 2286 708 2287 712
rect 2291 708 2292 712
rect 2286 707 2292 708
rect 2446 712 2452 713
rect 2446 708 2447 712
rect 2451 708 2452 712
rect 2446 707 2452 708
rect 2598 712 2604 713
rect 2598 708 2599 712
rect 2603 708 2604 712
rect 2598 707 2604 708
rect 2758 712 2764 713
rect 2758 708 2759 712
rect 2763 708 2764 712
rect 2758 707 2764 708
rect 2918 712 2924 713
rect 2918 708 2919 712
rect 2923 708 2924 712
rect 2918 707 2924 708
rect 2022 700 2028 701
rect 2022 696 2023 700
rect 2027 696 2028 700
rect 2022 695 2028 696
rect 2150 700 2156 701
rect 2150 696 2151 700
rect 2155 696 2156 700
rect 2150 695 2156 696
rect 2294 700 2300 701
rect 2294 696 2295 700
rect 2299 696 2300 700
rect 2294 695 2300 696
rect 2446 700 2452 701
rect 2446 696 2447 700
rect 2451 696 2452 700
rect 2446 695 2452 696
rect 2614 700 2620 701
rect 2614 696 2615 700
rect 2619 696 2620 700
rect 2614 695 2620 696
rect 2798 700 2804 701
rect 2798 696 2799 700
rect 2803 696 2804 700
rect 2798 695 2804 696
rect 2990 700 2996 701
rect 2990 696 2991 700
rect 2995 696 2996 700
rect 2990 695 2996 696
rect 3158 700 3164 701
rect 3158 696 3159 700
rect 3163 696 3164 700
rect 3158 695 3164 696
rect 1670 693 1676 694
rect 1670 689 1671 693
rect 1675 689 1676 693
rect 478 688 484 689
rect 478 684 479 688
rect 483 684 484 688
rect 478 683 484 684
rect 606 688 612 689
rect 606 684 607 688
rect 611 684 612 688
rect 606 683 612 684
rect 726 688 732 689
rect 726 684 727 688
rect 731 684 732 688
rect 726 683 732 684
rect 846 688 852 689
rect 846 684 847 688
rect 851 684 852 688
rect 846 683 852 684
rect 966 688 972 689
rect 966 684 967 688
rect 971 684 972 688
rect 966 683 972 684
rect 1078 688 1084 689
rect 1078 684 1079 688
rect 1083 684 1084 688
rect 1078 683 1084 684
rect 1190 688 1196 689
rect 1190 684 1191 688
rect 1195 684 1196 688
rect 1190 683 1196 684
rect 1310 688 1316 689
rect 1670 688 1676 689
rect 3190 693 3196 694
rect 3190 689 3191 693
rect 3195 689 3196 693
rect 3190 688 3196 689
rect 1310 684 1311 688
rect 1315 684 1316 688
rect 1310 683 1316 684
rect 110 681 116 682
rect 110 677 111 681
rect 115 677 116 681
rect 110 676 116 677
rect 1630 681 1636 682
rect 1630 677 1631 681
rect 1635 677 1636 681
rect 1630 676 1636 677
rect 2930 679 2936 680
rect 1670 675 1676 676
rect 1670 671 1671 675
rect 1675 671 1676 675
rect 2930 675 2931 679
rect 2935 678 2936 679
rect 2935 676 3002 678
rect 2935 675 2936 676
rect 2930 674 2936 675
rect 2999 675 3005 676
rect 1670 670 1676 671
rect 2022 671 2028 672
rect 2022 667 2023 671
rect 2027 667 2028 671
rect 2022 666 2028 667
rect 2030 671 2037 672
rect 2030 667 2031 671
rect 2036 667 2037 671
rect 2030 666 2037 667
rect 2150 671 2156 672
rect 2150 667 2151 671
rect 2155 667 2156 671
rect 2150 666 2156 667
rect 2158 671 2165 672
rect 2158 667 2159 671
rect 2164 667 2165 671
rect 2158 666 2165 667
rect 2294 671 2300 672
rect 2294 667 2295 671
rect 2299 667 2300 671
rect 2294 666 2300 667
rect 2303 671 2312 672
rect 2303 667 2304 671
rect 2311 667 2312 671
rect 2303 666 2312 667
rect 2446 671 2452 672
rect 2446 667 2447 671
rect 2451 667 2452 671
rect 2446 666 2452 667
rect 2455 671 2464 672
rect 2455 667 2456 671
rect 2463 667 2464 671
rect 2455 666 2464 667
rect 2614 671 2620 672
rect 2614 667 2615 671
rect 2619 667 2620 671
rect 2614 666 2620 667
rect 2622 671 2629 672
rect 2622 667 2623 671
rect 2628 667 2629 671
rect 2622 666 2629 667
rect 2798 671 2804 672
rect 2798 667 2799 671
rect 2803 667 2804 671
rect 2798 666 2804 667
rect 2806 671 2813 672
rect 2806 667 2807 671
rect 2812 670 2813 671
rect 2870 671 2876 672
rect 2870 670 2871 671
rect 2812 668 2871 670
rect 2812 667 2813 668
rect 2806 666 2813 667
rect 2870 667 2871 668
rect 2875 667 2876 671
rect 2870 666 2876 667
rect 2990 671 2996 672
rect 2990 667 2991 671
rect 2995 667 2996 671
rect 2999 671 3000 675
rect 3004 671 3005 675
rect 3166 675 3173 676
rect 2999 670 3005 671
rect 3158 671 3164 672
rect 2990 666 2996 667
rect 3158 667 3159 671
rect 3163 667 3164 671
rect 3166 671 3167 675
rect 3172 671 3173 675
rect 3166 670 3173 671
rect 3190 675 3196 676
rect 3190 671 3191 675
rect 3195 671 3196 675
rect 3190 670 3196 671
rect 3158 666 3164 667
rect 1240 664 1322 666
rect 110 663 116 664
rect 110 659 111 663
rect 115 659 116 663
rect 1199 663 1205 664
rect 110 658 116 659
rect 478 659 484 660
rect 478 655 479 659
rect 483 655 484 659
rect 478 654 484 655
rect 486 659 493 660
rect 486 655 487 659
rect 492 655 493 659
rect 486 654 493 655
rect 606 659 612 660
rect 606 655 607 659
rect 611 655 612 659
rect 606 654 612 655
rect 614 659 621 660
rect 614 655 615 659
rect 620 658 621 659
rect 630 659 636 660
rect 630 658 631 659
rect 620 656 631 658
rect 620 655 621 656
rect 614 654 621 655
rect 630 655 631 656
rect 635 655 636 659
rect 630 654 636 655
rect 726 659 732 660
rect 726 655 727 659
rect 731 655 732 659
rect 726 654 732 655
rect 735 659 741 660
rect 735 655 736 659
rect 740 658 741 659
rect 750 659 756 660
rect 750 658 751 659
rect 740 656 751 658
rect 740 655 741 656
rect 735 654 741 655
rect 750 655 751 656
rect 755 655 756 659
rect 750 654 756 655
rect 846 659 852 660
rect 846 655 847 659
rect 851 655 852 659
rect 846 654 852 655
rect 854 659 861 660
rect 854 655 855 659
rect 860 655 861 659
rect 854 654 861 655
rect 966 659 972 660
rect 966 655 967 659
rect 971 655 972 659
rect 966 654 972 655
rect 975 659 981 660
rect 975 655 976 659
rect 980 658 981 659
rect 998 659 1004 660
rect 998 658 999 659
rect 980 656 999 658
rect 980 655 981 656
rect 975 654 981 655
rect 998 655 999 656
rect 1003 655 1004 659
rect 998 654 1004 655
rect 1078 659 1084 660
rect 1078 655 1079 659
rect 1083 655 1084 659
rect 1078 654 1084 655
rect 1087 659 1093 660
rect 1087 655 1088 659
rect 1092 658 1093 659
rect 1102 659 1108 660
rect 1102 658 1103 659
rect 1092 656 1103 658
rect 1092 655 1093 656
rect 1087 654 1093 655
rect 1102 655 1103 656
rect 1107 655 1108 659
rect 1102 654 1108 655
rect 1190 659 1196 660
rect 1190 655 1191 659
rect 1195 655 1196 659
rect 1199 659 1200 663
rect 1204 662 1205 663
rect 1222 663 1228 664
rect 1222 662 1223 663
rect 1204 660 1223 662
rect 1204 659 1205 660
rect 1199 658 1205 659
rect 1222 659 1223 660
rect 1227 662 1228 663
rect 1240 662 1242 664
rect 1227 660 1242 662
rect 1318 663 1325 664
rect 1227 659 1228 660
rect 1222 658 1228 659
rect 1310 659 1316 660
rect 1190 654 1196 655
rect 1310 655 1311 659
rect 1315 655 1316 659
rect 1318 659 1319 663
rect 1324 659 1325 663
rect 1318 658 1325 659
rect 1630 663 1636 664
rect 1630 659 1631 663
rect 1635 659 1636 663
rect 1630 658 1636 659
rect 1310 654 1316 655
rect 1918 653 1924 654
rect 1670 649 1676 650
rect 1670 645 1671 649
rect 1675 645 1676 649
rect 1918 649 1919 653
rect 1923 649 1924 653
rect 1918 648 1924 649
rect 2046 653 2052 654
rect 2046 649 2047 653
rect 2051 649 2052 653
rect 2046 648 2052 649
rect 2182 653 2188 654
rect 2182 649 2183 653
rect 2187 649 2188 653
rect 2182 648 2188 649
rect 2326 653 2332 654
rect 2326 649 2327 653
rect 2331 649 2332 653
rect 2326 648 2332 649
rect 2470 653 2476 654
rect 2470 649 2471 653
rect 2475 649 2476 653
rect 2470 648 2476 649
rect 2614 653 2620 654
rect 2614 649 2615 653
rect 2619 649 2620 653
rect 2614 648 2620 649
rect 2758 653 2764 654
rect 2758 649 2759 653
rect 2763 649 2764 653
rect 2758 648 2764 649
rect 2766 651 2773 652
rect 1670 644 1676 645
rect 1894 647 1900 648
rect 1894 643 1895 647
rect 1899 646 1900 647
rect 1927 647 1933 648
rect 1927 646 1928 647
rect 1899 644 1928 646
rect 1899 643 1900 644
rect 1894 642 1900 643
rect 1927 643 1928 644
rect 1932 643 1933 647
rect 1927 642 1933 643
rect 2030 647 2036 648
rect 2030 643 2031 647
rect 2035 646 2036 647
rect 2055 647 2061 648
rect 2055 646 2056 647
rect 2035 644 2056 646
rect 2035 643 2036 644
rect 2030 642 2036 643
rect 2055 643 2056 644
rect 2060 646 2061 647
rect 2158 647 2164 648
rect 2158 646 2159 647
rect 2060 644 2159 646
rect 2060 643 2061 644
rect 2055 642 2061 643
rect 2158 643 2159 644
rect 2163 646 2164 647
rect 2190 647 2197 648
rect 2190 646 2191 647
rect 2163 644 2191 646
rect 2163 643 2164 644
rect 2158 642 2164 643
rect 2190 643 2191 644
rect 2196 643 2197 647
rect 2190 642 2197 643
rect 2306 647 2312 648
rect 2306 643 2307 647
rect 2311 646 2312 647
rect 2335 647 2341 648
rect 2335 646 2336 647
rect 2311 644 2336 646
rect 2311 643 2312 644
rect 2306 642 2312 643
rect 2335 643 2336 644
rect 2340 646 2341 647
rect 2458 647 2464 648
rect 2458 646 2459 647
rect 2340 644 2459 646
rect 2340 643 2341 644
rect 2335 642 2341 643
rect 2458 643 2459 644
rect 2463 646 2464 647
rect 2479 647 2485 648
rect 2479 646 2480 647
rect 2463 644 2480 646
rect 2463 643 2464 644
rect 2458 642 2464 643
rect 2479 643 2480 644
rect 2484 646 2485 647
rect 2622 647 2629 648
rect 2622 646 2623 647
rect 2484 644 2623 646
rect 2484 643 2485 644
rect 2479 642 2485 643
rect 2622 643 2623 644
rect 2628 646 2629 647
rect 2766 647 2767 651
rect 2772 650 2773 651
rect 2806 651 2812 652
rect 2806 650 2807 651
rect 2772 648 2807 650
rect 2772 647 2773 648
rect 2766 646 2773 647
rect 2806 647 2807 648
rect 2811 647 2812 651
rect 2806 646 2812 647
rect 3190 649 3196 650
rect 2628 644 2770 646
rect 3190 645 3191 649
rect 3195 645 3196 649
rect 3190 644 3196 645
rect 2628 643 2629 644
rect 2622 642 2629 643
rect 374 637 380 638
rect 110 633 116 634
rect 110 629 111 633
rect 115 629 116 633
rect 374 633 375 637
rect 379 633 380 637
rect 374 632 380 633
rect 502 637 508 638
rect 502 633 503 637
rect 507 633 508 637
rect 502 632 508 633
rect 622 637 628 638
rect 622 633 623 637
rect 627 633 628 637
rect 622 632 628 633
rect 742 637 748 638
rect 742 633 743 637
rect 747 633 748 637
rect 862 637 868 638
rect 742 632 748 633
rect 750 635 757 636
rect 110 628 116 629
rect 383 631 389 632
rect 383 627 384 631
rect 388 630 389 631
rect 406 631 412 632
rect 406 630 407 631
rect 388 628 407 630
rect 388 627 389 628
rect 383 626 389 627
rect 406 627 407 628
rect 411 630 412 631
rect 486 631 492 632
rect 486 630 487 631
rect 411 628 487 630
rect 411 627 412 628
rect 406 626 412 627
rect 486 627 487 628
rect 491 630 492 631
rect 511 631 517 632
rect 511 630 512 631
rect 491 628 512 630
rect 491 627 492 628
rect 486 626 492 627
rect 511 627 512 628
rect 516 627 517 631
rect 511 626 517 627
rect 630 631 637 632
rect 630 627 631 631
rect 636 630 637 631
rect 670 631 676 632
rect 670 630 671 631
rect 636 628 671 630
rect 636 627 637 628
rect 630 626 637 627
rect 670 627 671 628
rect 675 627 676 631
rect 750 631 751 635
rect 756 634 757 635
rect 774 635 780 636
rect 774 634 775 635
rect 756 632 775 634
rect 756 631 757 632
rect 750 630 757 631
rect 774 631 775 632
rect 779 634 780 635
rect 779 632 801 634
rect 862 633 863 637
rect 867 633 868 637
rect 862 632 868 633
rect 974 637 980 638
rect 974 633 975 637
rect 979 633 980 637
rect 974 632 980 633
rect 1094 637 1100 638
rect 1094 633 1095 637
rect 1099 633 1100 637
rect 1094 632 1100 633
rect 1214 637 1220 638
rect 1214 633 1215 637
rect 1219 633 1220 637
rect 1214 632 1220 633
rect 1222 635 1229 636
rect 779 631 780 632
rect 774 630 780 631
rect 799 630 801 632
rect 854 631 860 632
rect 854 630 855 631
rect 799 628 855 630
rect 670 626 676 627
rect 854 627 855 628
rect 859 630 860 631
rect 871 631 877 632
rect 871 630 872 631
rect 859 628 872 630
rect 859 627 860 628
rect 854 626 860 627
rect 871 627 872 628
rect 876 627 877 631
rect 871 626 877 627
rect 983 631 989 632
rect 983 627 984 631
rect 988 630 989 631
rect 998 631 1004 632
rect 998 630 999 631
rect 988 628 999 630
rect 988 627 989 628
rect 983 626 989 627
rect 998 627 999 628
rect 1003 630 1004 631
rect 1102 631 1109 632
rect 1102 630 1103 631
rect 1003 628 1103 630
rect 1003 627 1004 628
rect 998 626 1004 627
rect 1102 627 1103 628
rect 1108 630 1109 631
rect 1222 631 1223 635
rect 1228 631 1229 635
rect 1222 630 1229 631
rect 1630 633 1636 634
rect 1108 628 1226 630
rect 1630 629 1631 633
rect 1635 629 1636 633
rect 1630 628 1636 629
rect 1670 631 1676 632
rect 1108 627 1109 628
rect 1102 626 1109 627
rect 1670 627 1671 631
rect 1675 627 1676 631
rect 1670 626 1676 627
rect 3190 631 3196 632
rect 3190 627 3191 631
rect 3195 627 3196 631
rect 3190 626 3196 627
rect 1918 624 1924 625
rect 1918 620 1919 624
rect 1923 620 1924 624
rect 1918 619 1924 620
rect 2046 624 2052 625
rect 2046 620 2047 624
rect 2051 620 2052 624
rect 2046 619 2052 620
rect 2182 624 2188 625
rect 2182 620 2183 624
rect 2187 620 2188 624
rect 2182 619 2188 620
rect 2326 624 2332 625
rect 2326 620 2327 624
rect 2331 620 2332 624
rect 2326 619 2332 620
rect 2470 624 2476 625
rect 2470 620 2471 624
rect 2475 620 2476 624
rect 2470 619 2476 620
rect 2614 624 2620 625
rect 2614 620 2615 624
rect 2619 620 2620 624
rect 2614 619 2620 620
rect 2758 624 2764 625
rect 2758 620 2759 624
rect 2763 620 2764 624
rect 2758 619 2764 620
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 110 610 116 611
rect 1630 615 1636 616
rect 1630 611 1631 615
rect 1635 611 1636 615
rect 1630 610 1636 611
rect 374 608 380 609
rect 374 604 375 608
rect 379 604 380 608
rect 374 603 380 604
rect 502 608 508 609
rect 502 604 503 608
rect 507 604 508 608
rect 502 603 508 604
rect 622 608 628 609
rect 622 604 623 608
rect 627 604 628 608
rect 622 603 628 604
rect 742 608 748 609
rect 742 604 743 608
rect 747 604 748 608
rect 742 603 748 604
rect 862 608 868 609
rect 862 604 863 608
rect 867 604 868 608
rect 862 603 868 604
rect 974 608 980 609
rect 974 604 975 608
rect 979 604 980 608
rect 974 603 980 604
rect 1094 608 1100 609
rect 1094 604 1095 608
rect 1099 604 1100 608
rect 1094 603 1100 604
rect 1214 608 1220 609
rect 1214 604 1215 608
rect 1219 604 1220 608
rect 1214 603 1220 604
rect 1846 608 1852 609
rect 1846 604 1847 608
rect 1851 604 1852 608
rect 1846 603 1852 604
rect 2014 608 2020 609
rect 2014 604 2015 608
rect 2019 604 2020 608
rect 2014 603 2020 604
rect 2182 608 2188 609
rect 2182 604 2183 608
rect 2187 604 2188 608
rect 2182 603 2188 604
rect 2358 608 2364 609
rect 2358 604 2359 608
rect 2363 604 2364 608
rect 2358 603 2364 604
rect 2550 608 2556 609
rect 2550 604 2551 608
rect 2555 604 2556 608
rect 2550 603 2556 604
rect 2750 608 2756 609
rect 2750 604 2751 608
rect 2755 604 2756 608
rect 2750 603 2756 604
rect 2958 608 2964 609
rect 2958 604 2959 608
rect 2963 604 2964 608
rect 2958 603 2964 604
rect 3158 608 3164 609
rect 3158 604 3159 608
rect 3163 604 3164 608
rect 3158 603 3164 604
rect 1670 601 1676 602
rect 1670 597 1671 601
rect 1675 597 1676 601
rect 1670 596 1676 597
rect 3190 601 3196 602
rect 3190 597 3191 601
rect 3195 597 3196 601
rect 3190 596 3196 597
rect 270 588 276 589
rect 270 584 271 588
rect 275 584 276 588
rect 270 583 276 584
rect 398 588 404 589
rect 398 584 399 588
rect 403 584 404 588
rect 398 583 404 584
rect 526 588 532 589
rect 526 584 527 588
rect 531 584 532 588
rect 526 583 532 584
rect 646 588 652 589
rect 646 584 647 588
rect 651 584 652 588
rect 646 583 652 584
rect 766 588 772 589
rect 766 584 767 588
rect 771 584 772 588
rect 766 583 772 584
rect 878 588 884 589
rect 878 584 879 588
rect 883 584 884 588
rect 878 583 884 584
rect 990 588 996 589
rect 990 584 991 588
rect 995 584 996 588
rect 990 583 996 584
rect 1110 588 1116 589
rect 1110 584 1111 588
rect 1115 584 1116 588
rect 2967 585 3170 586
rect 1110 583 1116 584
rect 1670 583 1676 584
rect 110 581 116 582
rect 110 577 111 581
rect 115 577 116 581
rect 110 576 116 577
rect 1630 581 1636 582
rect 1630 577 1631 581
rect 1635 577 1636 581
rect 1670 579 1671 583
rect 1675 579 1676 583
rect 2190 583 2197 584
rect 1670 578 1676 579
rect 1846 579 1852 580
rect 1630 576 1636 577
rect 1846 575 1847 579
rect 1851 575 1852 579
rect 1846 574 1852 575
rect 1855 579 1861 580
rect 1855 575 1856 579
rect 1860 575 1861 579
rect 1855 574 1861 575
rect 2014 579 2020 580
rect 2014 575 2015 579
rect 2019 575 2020 579
rect 2014 574 2020 575
rect 2023 579 2029 580
rect 2023 575 2024 579
rect 2028 575 2029 579
rect 2023 574 2029 575
rect 2182 579 2188 580
rect 2182 575 2183 579
rect 2187 575 2188 579
rect 2190 579 2191 583
rect 2196 582 2197 583
rect 2759 583 2765 584
rect 2196 580 2241 582
rect 2196 579 2197 580
rect 2190 578 2197 579
rect 2239 578 2241 580
rect 2358 579 2364 580
rect 2239 576 2259 578
rect 2182 574 2188 575
rect 1766 569 1772 570
rect 1670 565 1676 566
rect 110 563 116 564
rect 110 559 111 563
rect 115 559 116 563
rect 775 563 781 564
rect 110 558 116 559
rect 270 559 276 560
rect 270 555 271 559
rect 275 555 276 559
rect 270 554 276 555
rect 279 559 285 560
rect 279 555 280 559
rect 284 558 285 559
rect 310 559 316 560
rect 310 558 311 559
rect 284 556 311 558
rect 284 555 285 556
rect 279 554 285 555
rect 310 555 311 556
rect 315 555 316 559
rect 310 554 316 555
rect 398 559 404 560
rect 398 555 399 559
rect 403 555 404 559
rect 398 554 404 555
rect 406 559 413 560
rect 406 555 407 559
rect 412 558 413 559
rect 430 559 436 560
rect 430 558 431 559
rect 412 556 431 558
rect 412 555 413 556
rect 406 554 413 555
rect 430 555 431 556
rect 435 555 436 559
rect 430 554 436 555
rect 526 559 532 560
rect 526 555 527 559
rect 531 555 532 559
rect 526 554 532 555
rect 535 559 541 560
rect 535 555 536 559
rect 540 558 541 559
rect 550 559 556 560
rect 550 558 551 559
rect 540 556 551 558
rect 540 555 541 556
rect 535 554 541 555
rect 550 555 551 556
rect 555 555 556 559
rect 550 554 556 555
rect 646 559 652 560
rect 646 555 647 559
rect 651 555 652 559
rect 646 554 652 555
rect 655 559 661 560
rect 655 555 656 559
rect 660 558 661 559
rect 670 559 676 560
rect 670 558 671 559
rect 660 556 671 558
rect 660 555 661 556
rect 655 554 661 555
rect 670 555 671 556
rect 675 555 676 559
rect 670 554 676 555
rect 766 559 772 560
rect 766 555 767 559
rect 771 555 772 559
rect 775 559 776 563
rect 780 559 781 563
rect 1630 563 1636 564
rect 775 558 781 559
rect 878 559 884 560
rect 766 554 772 555
rect 878 555 879 559
rect 883 555 884 559
rect 878 554 884 555
rect 886 559 893 560
rect 886 555 887 559
rect 892 555 893 559
rect 886 554 893 555
rect 990 559 996 560
rect 990 555 991 559
rect 995 555 996 559
rect 990 554 996 555
rect 998 559 1005 560
rect 998 555 999 559
rect 1004 555 1005 559
rect 998 554 1005 555
rect 1110 559 1116 560
rect 1110 555 1111 559
rect 1115 555 1116 559
rect 1110 554 1116 555
rect 1119 559 1125 560
rect 1119 555 1120 559
rect 1124 558 1125 559
rect 1142 559 1148 560
rect 1142 558 1143 559
rect 1124 556 1143 558
rect 1124 555 1125 556
rect 1119 554 1125 555
rect 1142 555 1143 556
rect 1147 555 1148 559
rect 1630 559 1631 563
rect 1635 559 1636 563
rect 1670 561 1671 565
rect 1675 561 1676 565
rect 1766 565 1767 569
rect 1771 565 1772 569
rect 1766 564 1772 565
rect 1775 567 1781 568
rect 1775 563 1776 567
rect 1780 566 1781 567
rect 1857 566 1859 574
rect 1926 569 1932 570
rect 1894 567 1900 568
rect 1894 566 1895 567
rect 1780 564 1895 566
rect 1780 563 1781 564
rect 1775 562 1781 563
rect 1894 563 1895 564
rect 1899 563 1900 567
rect 1926 565 1927 569
rect 1931 565 1932 569
rect 1926 564 1932 565
rect 1894 562 1900 563
rect 1935 563 1941 564
rect 1935 562 1936 563
rect 1670 560 1676 561
rect 1896 560 1936 562
rect 1630 558 1636 559
rect 1935 559 1936 560
rect 1940 562 1941 563
rect 2025 562 2027 574
rect 2086 569 2092 570
rect 2086 565 2087 569
rect 2091 565 2092 569
rect 2086 564 2092 565
rect 2246 569 2252 570
rect 2246 565 2247 569
rect 2251 565 2252 569
rect 2257 568 2259 576
rect 2358 575 2359 579
rect 2363 575 2364 579
rect 2358 574 2364 575
rect 2367 579 2373 580
rect 2367 575 2368 579
rect 2372 578 2373 579
rect 2414 579 2420 580
rect 2414 578 2415 579
rect 2372 576 2415 578
rect 2372 575 2373 576
rect 2367 574 2373 575
rect 2414 575 2415 576
rect 2419 575 2420 579
rect 2414 574 2420 575
rect 2550 579 2556 580
rect 2550 575 2551 579
rect 2555 575 2556 579
rect 2550 574 2556 575
rect 2559 579 2565 580
rect 2559 575 2560 579
rect 2564 578 2565 579
rect 2750 579 2756 580
rect 2564 576 2579 578
rect 2564 575 2565 576
rect 2559 574 2565 575
rect 2406 569 2412 570
rect 2246 564 2252 565
rect 2255 567 2261 568
rect 2030 563 2036 564
rect 2030 562 2031 563
rect 1940 560 2031 562
rect 1940 559 1941 560
rect 1935 558 1941 559
rect 2030 559 2031 560
rect 2035 562 2036 563
rect 2095 563 2101 564
rect 2095 562 2096 563
rect 2035 560 2096 562
rect 2035 559 2036 560
rect 2030 558 2036 559
rect 2095 559 2096 560
rect 2100 562 2101 563
rect 2110 563 2116 564
rect 2110 562 2111 563
rect 2100 560 2111 562
rect 2100 559 2101 560
rect 2095 558 2101 559
rect 2110 559 2111 560
rect 2115 559 2116 563
rect 2255 563 2256 567
rect 2260 563 2261 567
rect 2406 565 2407 569
rect 2411 565 2412 569
rect 2566 569 2572 570
rect 2406 564 2412 565
rect 2414 567 2421 568
rect 2255 562 2261 563
rect 2414 563 2415 567
rect 2420 566 2421 567
rect 2458 567 2464 568
rect 2458 566 2459 567
rect 2420 564 2459 566
rect 2420 563 2421 564
rect 2414 562 2421 563
rect 2458 563 2459 564
rect 2463 563 2464 567
rect 2566 565 2567 569
rect 2571 565 2572 569
rect 2566 564 2572 565
rect 2577 564 2579 576
rect 2750 575 2751 579
rect 2755 575 2756 579
rect 2759 579 2760 583
rect 2764 579 2765 583
rect 2967 581 2968 585
rect 2972 584 3170 585
rect 2972 581 2973 584
rect 2967 580 2973 581
rect 3166 583 3173 584
rect 2759 578 2765 579
rect 2958 579 2964 580
rect 2750 574 2756 575
rect 2958 575 2959 579
rect 2963 575 2964 579
rect 2958 574 2964 575
rect 3158 579 3164 580
rect 3158 575 3159 579
rect 3163 575 3164 579
rect 3166 579 3167 583
rect 3172 579 3173 583
rect 3166 578 3173 579
rect 3190 583 3196 584
rect 3190 579 3191 583
rect 3195 579 3196 583
rect 3190 578 3196 579
rect 3158 574 3164 575
rect 3190 565 3196 566
rect 2458 562 2464 563
rect 2575 563 2581 564
rect 2110 558 2116 559
rect 2575 559 2576 563
rect 2580 562 2581 563
rect 2606 563 2612 564
rect 2606 562 2607 563
rect 2580 560 2607 562
rect 2580 559 2581 560
rect 2575 558 2581 559
rect 2606 559 2607 560
rect 2611 559 2612 563
rect 3190 561 3191 565
rect 3195 561 3196 565
rect 3190 560 3196 561
rect 2606 558 2612 559
rect 1142 554 1148 555
rect 310 551 316 552
rect 310 547 311 551
rect 315 550 316 551
rect 430 551 436 552
rect 430 550 431 551
rect 315 548 431 550
rect 315 547 316 548
rect 310 546 316 547
rect 430 547 431 548
rect 435 547 436 551
rect 430 546 436 547
rect 1670 547 1676 548
rect 1670 543 1671 547
rect 1675 543 1676 547
rect 1670 542 1676 543
rect 3190 547 3196 548
rect 3190 543 3191 547
rect 3195 543 3196 547
rect 3190 542 3196 543
rect 1766 540 1772 541
rect 174 537 180 538
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 174 533 175 537
rect 179 533 180 537
rect 174 532 180 533
rect 302 537 308 538
rect 302 533 303 537
rect 307 533 308 537
rect 302 532 308 533
rect 422 537 428 538
rect 422 533 423 537
rect 427 533 428 537
rect 542 537 548 538
rect 422 532 428 533
rect 430 535 437 536
rect 110 528 116 529
rect 146 531 152 532
rect 146 527 147 531
rect 151 530 152 531
rect 183 531 189 532
rect 183 530 184 531
rect 151 528 184 530
rect 151 527 152 528
rect 146 526 152 527
rect 183 527 184 528
rect 188 530 189 531
rect 310 531 317 532
rect 310 530 311 531
rect 188 528 311 530
rect 188 527 189 528
rect 183 526 189 527
rect 310 527 311 528
rect 316 527 317 531
rect 430 531 431 535
rect 436 531 437 535
rect 542 533 543 537
rect 547 533 548 537
rect 542 532 548 533
rect 662 537 668 538
rect 662 533 663 537
rect 667 533 668 537
rect 662 532 668 533
rect 774 537 780 538
rect 774 533 775 537
rect 779 533 780 537
rect 886 537 892 538
rect 774 532 780 533
rect 782 535 789 536
rect 430 530 437 531
rect 550 531 557 532
rect 310 526 317 527
rect 550 527 551 531
rect 556 530 557 531
rect 670 531 677 532
rect 670 530 671 531
rect 556 528 671 530
rect 556 527 557 528
rect 550 526 557 527
rect 670 527 671 528
rect 676 527 677 531
rect 782 531 783 535
rect 788 534 789 535
rect 788 532 801 534
rect 886 533 887 537
rect 891 533 892 537
rect 886 532 892 533
rect 1006 537 1012 538
rect 1006 533 1007 537
rect 1011 533 1012 537
rect 1766 536 1767 540
rect 1771 536 1772 540
rect 1766 535 1772 536
rect 1926 540 1932 541
rect 1926 536 1927 540
rect 1931 536 1932 540
rect 1926 535 1932 536
rect 2086 540 2092 541
rect 2086 536 2087 540
rect 2091 536 2092 540
rect 2086 535 2092 536
rect 2246 540 2252 541
rect 2246 536 2247 540
rect 2251 536 2252 540
rect 2246 535 2252 536
rect 2406 540 2412 541
rect 2406 536 2407 540
rect 2411 536 2412 540
rect 2406 535 2412 536
rect 2566 540 2572 541
rect 2566 536 2567 540
rect 2571 536 2572 540
rect 2566 535 2572 536
rect 1006 532 1012 533
rect 1630 533 1636 534
rect 788 531 789 532
rect 782 530 789 531
rect 799 530 801 532
rect 826 531 832 532
rect 826 530 827 531
rect 799 528 827 530
rect 670 526 677 527
rect 826 527 827 528
rect 831 530 832 531
rect 894 531 901 532
rect 894 530 895 531
rect 831 528 895 530
rect 831 527 832 528
rect 826 526 832 527
rect 894 527 895 528
rect 900 530 901 531
rect 998 531 1004 532
rect 998 530 999 531
rect 900 528 999 530
rect 900 527 901 528
rect 894 526 901 527
rect 998 527 999 528
rect 1003 530 1004 531
rect 1015 531 1021 532
rect 1015 530 1016 531
rect 1003 528 1016 530
rect 1003 527 1004 528
rect 998 526 1004 527
rect 1015 527 1016 528
rect 1020 527 1021 531
rect 1630 529 1631 533
rect 1635 529 1636 533
rect 1630 528 1636 529
rect 1694 528 1700 529
rect 1015 526 1021 527
rect 1694 524 1695 528
rect 1699 524 1700 528
rect 1694 523 1700 524
rect 1886 528 1892 529
rect 1886 524 1887 528
rect 1891 524 1892 528
rect 1886 523 1892 524
rect 2102 528 2108 529
rect 2102 524 2103 528
rect 2107 524 2108 528
rect 2102 523 2108 524
rect 2342 528 2348 529
rect 2342 524 2343 528
rect 2347 524 2348 528
rect 2342 523 2348 524
rect 2598 528 2604 529
rect 2598 524 2599 528
rect 2603 524 2604 528
rect 2598 523 2604 524
rect 2862 528 2868 529
rect 2862 524 2863 528
rect 2867 524 2868 528
rect 2862 523 2868 524
rect 3134 528 3140 529
rect 3134 524 3135 528
rect 3139 524 3140 528
rect 3134 523 3140 524
rect 1670 521 1676 522
rect 1670 517 1671 521
rect 1675 517 1676 521
rect 1670 516 1676 517
rect 3190 521 3196 522
rect 3190 517 3191 521
rect 3195 517 3196 521
rect 3190 516 3196 517
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 110 510 116 511
rect 1630 515 1636 516
rect 1630 511 1631 515
rect 1635 511 1636 515
rect 1630 510 1636 511
rect 174 508 180 509
rect 174 504 175 508
rect 179 504 180 508
rect 174 503 180 504
rect 302 508 308 509
rect 302 504 303 508
rect 307 504 308 508
rect 302 503 308 504
rect 422 508 428 509
rect 422 504 423 508
rect 427 504 428 508
rect 422 503 428 504
rect 542 508 548 509
rect 542 504 543 508
rect 547 504 548 508
rect 542 503 548 504
rect 662 508 668 509
rect 662 504 663 508
rect 667 504 668 508
rect 662 503 668 504
rect 774 508 780 509
rect 774 504 775 508
rect 779 504 780 508
rect 774 503 780 504
rect 886 508 892 509
rect 886 504 887 508
rect 891 504 892 508
rect 886 503 892 504
rect 1006 508 1012 509
rect 1006 504 1007 508
rect 1011 504 1012 508
rect 1006 503 1012 504
rect 1670 503 1676 504
rect 1670 499 1671 503
rect 1675 499 1676 503
rect 1894 503 1901 504
rect 1670 498 1676 499
rect 1694 499 1700 500
rect 1694 495 1695 499
rect 1699 495 1700 499
rect 1694 494 1700 495
rect 1702 499 1709 500
rect 1702 495 1703 499
rect 1708 495 1709 499
rect 1702 494 1709 495
rect 1886 499 1892 500
rect 1886 495 1887 499
rect 1891 495 1892 499
rect 1894 499 1895 503
rect 1900 499 1901 503
rect 2110 503 2117 504
rect 1894 498 1901 499
rect 2102 499 2108 500
rect 1886 494 1892 495
rect 2102 495 2103 499
rect 2107 495 2108 499
rect 2110 499 2111 503
rect 2116 499 2117 503
rect 2351 503 2357 504
rect 2110 498 2117 499
rect 2342 499 2348 500
rect 2102 494 2108 495
rect 2342 495 2343 499
rect 2347 495 2348 499
rect 2351 499 2352 503
rect 2356 502 2357 503
rect 2414 503 2420 504
rect 2414 502 2415 503
rect 2356 500 2415 502
rect 2356 499 2357 500
rect 2351 498 2357 499
rect 2414 499 2415 500
rect 2419 499 2420 503
rect 3142 503 3149 504
rect 2414 498 2420 499
rect 2598 499 2604 500
rect 2342 494 2348 495
rect 2598 495 2599 499
rect 2603 495 2604 499
rect 2598 494 2604 495
rect 2606 499 2613 500
rect 2606 495 2607 499
rect 2612 498 2613 499
rect 2630 499 2636 500
rect 2630 498 2631 499
rect 2612 496 2631 498
rect 2612 495 2613 496
rect 2606 494 2613 495
rect 2630 495 2631 496
rect 2635 495 2636 499
rect 2630 494 2636 495
rect 2862 499 2868 500
rect 2862 495 2863 499
rect 2867 495 2868 499
rect 2862 494 2868 495
rect 2870 499 2877 500
rect 2870 495 2871 499
rect 2876 498 2877 499
rect 2926 499 2932 500
rect 2926 498 2927 499
rect 2876 496 2927 498
rect 2876 495 2877 496
rect 2870 494 2877 495
rect 2926 495 2927 496
rect 2931 495 2932 499
rect 2926 494 2932 495
rect 3134 499 3140 500
rect 3134 495 3135 499
rect 3139 495 3140 499
rect 3142 499 3143 503
rect 3148 502 3149 503
rect 3166 503 3172 504
rect 3166 502 3167 503
rect 3148 500 3167 502
rect 3148 499 3149 500
rect 3142 498 3149 499
rect 3166 499 3167 500
rect 3171 499 3172 503
rect 3166 498 3172 499
rect 3190 503 3196 504
rect 3190 499 3191 503
rect 3195 499 3196 503
rect 3190 498 3196 499
rect 3134 494 3140 495
rect 134 484 140 485
rect 134 480 135 484
rect 139 480 140 484
rect 134 479 140 480
rect 230 484 236 485
rect 230 480 231 484
rect 235 480 236 484
rect 230 479 236 480
rect 358 484 364 485
rect 358 480 359 484
rect 363 480 364 484
rect 358 479 364 480
rect 502 484 508 485
rect 502 480 503 484
rect 507 480 508 484
rect 502 479 508 480
rect 654 484 660 485
rect 654 480 655 484
rect 659 480 660 484
rect 654 479 660 480
rect 814 484 820 485
rect 814 480 815 484
rect 819 480 820 484
rect 814 479 820 480
rect 974 484 980 485
rect 974 480 975 484
rect 979 480 980 484
rect 974 479 980 480
rect 1134 484 1140 485
rect 1134 480 1135 484
rect 1139 480 1140 484
rect 1134 479 1140 480
rect 1294 484 1300 485
rect 1294 480 1295 484
rect 1299 480 1300 484
rect 1294 479 1300 480
rect 1454 484 1460 485
rect 1454 480 1455 484
rect 1459 480 1460 484
rect 1454 479 1460 480
rect 1598 484 1604 485
rect 1598 480 1599 484
rect 1603 480 1604 484
rect 1598 479 1604 480
rect 1694 481 1700 482
rect 110 477 116 478
rect 110 473 111 477
rect 115 473 116 477
rect 110 472 116 473
rect 1630 477 1636 478
rect 1630 473 1631 477
rect 1635 473 1636 477
rect 1630 472 1636 473
rect 1670 477 1676 478
rect 1670 473 1671 477
rect 1675 473 1676 477
rect 1694 477 1695 481
rect 1699 477 1700 481
rect 2022 481 2028 482
rect 1694 476 1700 477
rect 1702 479 1709 480
rect 1702 475 1703 479
rect 1708 475 1709 479
rect 2022 477 2023 481
rect 2027 477 2028 481
rect 2382 481 2388 482
rect 2022 476 2028 477
rect 2030 479 2037 480
rect 1702 474 1709 475
rect 2030 475 2031 479
rect 2036 478 2037 479
rect 2058 479 2064 480
rect 2058 478 2059 479
rect 2036 476 2059 478
rect 2036 475 2037 476
rect 2030 474 2037 475
rect 2058 475 2059 476
rect 2063 475 2064 479
rect 2382 477 2383 481
rect 2387 477 2388 481
rect 2742 481 2748 482
rect 2382 476 2388 477
rect 2391 479 2397 480
rect 2058 474 2064 475
rect 2391 475 2392 479
rect 2396 478 2397 479
rect 2414 479 2420 480
rect 2414 478 2415 479
rect 2396 476 2415 478
rect 2396 475 2397 476
rect 2391 474 2397 475
rect 2414 475 2415 476
rect 2419 475 2420 479
rect 2742 477 2743 481
rect 2747 477 2748 481
rect 2742 476 2748 477
rect 3110 481 3116 482
rect 3110 477 3111 481
rect 3115 477 3116 481
rect 3110 476 3116 477
rect 3118 479 3125 480
rect 2414 474 2420 475
rect 2750 475 2757 476
rect 1670 472 1676 473
rect 2750 471 2751 475
rect 2756 471 2757 475
rect 3118 475 3119 479
rect 3124 478 3125 479
rect 3142 479 3148 480
rect 3142 478 3143 479
rect 3124 476 3143 478
rect 3124 475 3125 476
rect 3118 474 3125 475
rect 3142 475 3143 476
rect 3147 475 3148 479
rect 3142 474 3148 475
rect 3190 477 3196 478
rect 3190 473 3191 477
rect 3195 473 3196 477
rect 3190 472 3196 473
rect 2750 470 2757 471
rect 1606 467 1612 468
rect 470 463 476 464
rect 470 462 471 463
rect 148 460 471 462
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 143 459 152 460
rect 110 454 116 455
rect 134 455 140 456
rect 134 451 135 455
rect 139 451 140 455
rect 143 455 144 459
rect 151 455 152 459
rect 239 459 245 460
rect 143 454 152 455
rect 230 455 236 456
rect 134 450 140 451
rect 230 451 231 455
rect 235 451 236 455
rect 239 455 240 459
rect 244 455 245 459
rect 367 459 373 460
rect 239 454 245 455
rect 358 455 364 456
rect 230 450 236 451
rect 358 451 359 455
rect 363 451 364 455
rect 367 455 368 459
rect 372 455 373 459
rect 470 459 471 460
rect 475 462 476 463
rect 1606 463 1607 467
rect 1611 466 1612 467
rect 1702 467 1708 468
rect 1702 466 1703 467
rect 1611 464 1703 466
rect 1611 463 1612 464
rect 1606 462 1612 463
rect 1702 463 1703 464
rect 1707 463 1708 467
rect 1702 462 1708 463
rect 475 460 515 462
rect 475 459 476 460
rect 470 458 476 459
rect 511 459 517 460
rect 367 454 373 455
rect 502 455 508 456
rect 358 450 364 451
rect 502 451 503 455
rect 507 451 508 455
rect 511 455 512 459
rect 516 455 517 459
rect 1142 459 1149 460
rect 663 457 669 458
rect 663 456 664 457
rect 511 454 517 455
rect 654 455 660 456
rect 502 450 508 451
rect 654 451 655 455
rect 659 451 660 455
rect 654 450 660 451
rect 662 455 664 456
rect 662 451 663 455
rect 668 453 669 457
rect 667 452 669 453
rect 814 455 820 456
rect 667 451 668 452
rect 662 450 668 451
rect 814 451 815 455
rect 819 451 820 455
rect 814 450 820 451
rect 823 455 832 456
rect 823 451 824 455
rect 831 451 832 455
rect 823 450 832 451
rect 974 455 980 456
rect 974 451 975 455
rect 979 451 980 455
rect 974 450 980 451
rect 982 455 989 456
rect 982 451 983 455
rect 988 451 989 455
rect 982 450 989 451
rect 1134 455 1140 456
rect 1134 451 1135 455
rect 1139 451 1140 455
rect 1142 455 1143 459
rect 1148 455 1149 459
rect 1630 459 1636 460
rect 1142 454 1149 455
rect 1294 455 1300 456
rect 1134 450 1140 451
rect 1294 451 1295 455
rect 1299 451 1300 455
rect 1294 450 1300 451
rect 1303 455 1309 456
rect 1303 451 1304 455
rect 1308 454 1309 455
rect 1342 455 1348 456
rect 1342 454 1343 455
rect 1308 452 1343 454
rect 1308 451 1309 452
rect 1303 450 1309 451
rect 1342 451 1343 452
rect 1347 451 1348 455
rect 1342 450 1348 451
rect 1454 455 1460 456
rect 1454 451 1455 455
rect 1459 451 1460 455
rect 1454 450 1460 451
rect 1463 455 1472 456
rect 1463 451 1464 455
rect 1471 451 1472 455
rect 1463 450 1472 451
rect 1598 455 1604 456
rect 1598 451 1599 455
rect 1603 451 1604 455
rect 1598 450 1604 451
rect 1606 455 1613 456
rect 1606 451 1607 455
rect 1612 451 1613 455
rect 1630 455 1631 459
rect 1635 455 1636 459
rect 1630 454 1636 455
rect 1670 459 1676 460
rect 1670 455 1671 459
rect 1675 455 1676 459
rect 1670 454 1676 455
rect 3190 459 3196 460
rect 3190 455 3191 459
rect 3195 455 3196 459
rect 3190 454 3196 455
rect 1606 450 1613 451
rect 1694 452 1700 453
rect 1694 448 1695 452
rect 1699 448 1700 452
rect 1694 447 1700 448
rect 2022 452 2028 453
rect 2022 448 2023 452
rect 2027 448 2028 452
rect 2022 447 2028 448
rect 2382 452 2388 453
rect 2382 448 2383 452
rect 2387 448 2388 452
rect 2382 447 2388 448
rect 2742 452 2748 453
rect 2742 448 2743 452
rect 2747 448 2748 452
rect 2742 447 2748 448
rect 3110 452 3116 453
rect 3110 448 3111 452
rect 3115 448 3116 452
rect 3110 447 3116 448
rect 1142 439 1148 440
rect 1142 435 1143 439
rect 1147 438 1148 439
rect 1230 439 1236 440
rect 1230 438 1231 439
rect 1147 436 1231 438
rect 1147 435 1148 436
rect 1142 434 1148 435
rect 1230 435 1231 436
rect 1235 435 1236 439
rect 1230 434 1236 435
rect 1466 439 1472 440
rect 1466 435 1467 439
rect 1471 438 1472 439
rect 1606 439 1612 440
rect 1606 438 1607 439
rect 1471 436 1607 438
rect 1471 435 1472 436
rect 1466 434 1472 435
rect 1606 435 1607 436
rect 1611 435 1612 439
rect 1606 434 1612 435
rect 2246 436 2252 437
rect 726 433 732 434
rect 110 429 116 430
rect 110 425 111 429
rect 115 425 116 429
rect 726 429 727 433
rect 731 429 732 433
rect 726 428 732 429
rect 854 433 860 434
rect 854 429 855 433
rect 859 429 860 433
rect 854 428 860 429
rect 982 433 988 434
rect 982 429 983 433
rect 987 429 988 433
rect 982 428 988 429
rect 1102 433 1108 434
rect 1102 429 1103 433
rect 1107 429 1108 433
rect 1222 433 1228 434
rect 1102 428 1108 429
rect 1111 431 1117 432
rect 110 424 116 425
rect 735 427 741 428
rect 735 423 736 427
rect 740 426 741 427
rect 814 427 820 428
rect 814 426 815 427
rect 740 424 815 426
rect 740 423 741 424
rect 735 422 741 423
rect 814 423 815 424
rect 819 426 820 427
rect 826 427 832 428
rect 826 426 827 427
rect 819 424 827 426
rect 819 423 820 424
rect 814 422 820 423
rect 826 423 827 424
rect 831 426 832 427
rect 863 427 869 428
rect 863 426 864 427
rect 831 424 864 426
rect 831 423 832 424
rect 826 422 832 423
rect 863 423 864 424
rect 868 423 869 427
rect 863 422 869 423
rect 990 427 997 428
rect 990 423 991 427
rect 996 426 997 427
rect 1111 427 1112 431
rect 1116 430 1117 431
rect 1142 431 1148 432
rect 1142 430 1143 431
rect 1116 428 1143 430
rect 1116 427 1117 428
rect 1111 426 1117 427
rect 1142 427 1143 428
rect 1147 427 1148 431
rect 1222 429 1223 433
rect 1227 429 1228 433
rect 1334 433 1340 434
rect 1222 428 1228 429
rect 1230 431 1237 432
rect 1142 426 1148 427
rect 1230 427 1231 431
rect 1236 427 1237 431
rect 1334 429 1335 433
rect 1339 429 1340 433
rect 1334 428 1340 429
rect 1446 433 1452 434
rect 1446 429 1447 433
rect 1451 429 1452 433
rect 1446 428 1452 429
rect 1455 433 1461 434
rect 1455 429 1456 433
rect 1460 432 1461 433
rect 1566 433 1572 434
rect 1460 431 1472 432
rect 1460 430 1467 431
rect 1460 429 1461 430
rect 1455 428 1461 429
rect 1465 428 1467 430
rect 1230 426 1237 427
rect 1342 427 1349 428
rect 996 424 1114 426
rect 996 423 997 424
rect 990 422 997 423
rect 1342 423 1343 427
rect 1348 423 1349 427
rect 1466 427 1467 428
rect 1471 427 1472 431
rect 1566 429 1567 433
rect 1571 429 1572 433
rect 2246 432 2247 436
rect 2251 432 2252 436
rect 1566 428 1572 429
rect 1575 431 1581 432
rect 1466 426 1472 427
rect 1575 427 1576 431
rect 1580 430 1581 431
rect 1606 431 1612 432
rect 2246 431 2252 432
rect 2374 436 2380 437
rect 2374 432 2375 436
rect 2379 432 2380 436
rect 2374 431 2380 432
rect 2502 436 2508 437
rect 2502 432 2503 436
rect 2507 432 2508 436
rect 2502 431 2508 432
rect 2622 436 2628 437
rect 2622 432 2623 436
rect 2627 432 2628 436
rect 2622 431 2628 432
rect 2742 436 2748 437
rect 2742 432 2743 436
rect 2747 432 2748 436
rect 2742 431 2748 432
rect 2854 436 2860 437
rect 2854 432 2855 436
rect 2859 432 2860 436
rect 2854 431 2860 432
rect 2966 436 2972 437
rect 2966 432 2967 436
rect 2971 432 2972 436
rect 2966 431 2972 432
rect 3086 436 3092 437
rect 3086 432 3087 436
rect 3091 432 3092 436
rect 3086 431 3092 432
rect 1606 430 1607 431
rect 1580 428 1607 430
rect 1580 427 1581 428
rect 1575 426 1581 427
rect 1606 427 1607 428
rect 1611 427 1612 431
rect 1606 426 1612 427
rect 1630 429 1636 430
rect 1630 425 1631 429
rect 1635 425 1636 429
rect 1630 424 1636 425
rect 1670 429 1676 430
rect 1670 425 1671 429
rect 1675 425 1676 429
rect 1670 424 1676 425
rect 3190 429 3196 430
rect 3190 425 3191 429
rect 3195 425 3196 429
rect 3190 424 3196 425
rect 1342 422 1349 423
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 110 406 116 407
rect 1630 411 1636 412
rect 1630 407 1631 411
rect 1635 407 1636 411
rect 1630 406 1636 407
rect 1670 411 1676 412
rect 1670 407 1671 411
rect 1675 407 1676 411
rect 2862 411 2869 412
rect 1670 406 1676 407
rect 2246 407 2252 408
rect 726 404 732 405
rect 726 400 727 404
rect 731 400 732 404
rect 726 399 732 400
rect 854 404 860 405
rect 854 400 855 404
rect 859 400 860 404
rect 854 399 860 400
rect 982 404 988 405
rect 982 400 983 404
rect 987 400 988 404
rect 982 399 988 400
rect 1102 404 1108 405
rect 1102 400 1103 404
rect 1107 400 1108 404
rect 1102 399 1108 400
rect 1222 404 1228 405
rect 1222 400 1223 404
rect 1227 400 1228 404
rect 1222 399 1228 400
rect 1334 404 1340 405
rect 1334 400 1335 404
rect 1339 400 1340 404
rect 1334 399 1340 400
rect 1446 404 1452 405
rect 1446 400 1447 404
rect 1451 400 1452 404
rect 1446 399 1452 400
rect 1566 404 1572 405
rect 1566 400 1567 404
rect 1571 400 1572 404
rect 2246 403 2247 407
rect 2251 403 2252 407
rect 2246 402 2252 403
rect 2255 407 2264 408
rect 2255 403 2256 407
rect 2263 403 2264 407
rect 2255 402 2264 403
rect 2374 407 2380 408
rect 2374 403 2375 407
rect 2379 403 2380 407
rect 2374 402 2380 403
rect 2383 407 2392 408
rect 2383 403 2384 407
rect 2391 403 2392 407
rect 2383 402 2392 403
rect 2502 407 2508 408
rect 2502 403 2503 407
rect 2507 403 2508 407
rect 2502 402 2508 403
rect 2511 407 2520 408
rect 2511 403 2512 407
rect 2519 403 2520 407
rect 2511 402 2520 403
rect 2622 407 2628 408
rect 2622 403 2623 407
rect 2627 403 2628 407
rect 2622 402 2628 403
rect 2630 407 2637 408
rect 2630 403 2631 407
rect 2636 406 2637 407
rect 2670 407 2676 408
rect 2670 406 2671 407
rect 2636 404 2671 406
rect 2636 403 2637 404
rect 2630 402 2637 403
rect 2670 403 2671 404
rect 2675 403 2676 407
rect 2670 402 2676 403
rect 2742 407 2748 408
rect 2742 403 2743 407
rect 2747 403 2748 407
rect 2742 402 2748 403
rect 2750 407 2757 408
rect 2750 403 2751 407
rect 2756 406 2757 407
rect 2798 407 2804 408
rect 2798 406 2799 407
rect 2756 404 2799 406
rect 2756 403 2757 404
rect 2750 402 2757 403
rect 2798 403 2799 404
rect 2803 403 2804 407
rect 2798 402 2804 403
rect 2854 407 2860 408
rect 2854 403 2855 407
rect 2859 403 2860 407
rect 2862 407 2863 411
rect 2868 410 2869 411
rect 2926 411 2932 412
rect 2926 410 2927 411
rect 2868 408 2927 410
rect 2868 407 2869 408
rect 2862 406 2869 407
rect 2926 407 2927 408
rect 2931 407 2932 411
rect 3095 411 3101 412
rect 2926 406 2932 407
rect 2966 407 2972 408
rect 2854 402 2860 403
rect 2966 403 2967 407
rect 2971 403 2972 407
rect 2966 402 2972 403
rect 2974 407 2981 408
rect 2974 403 2975 407
rect 2980 406 2981 407
rect 3034 407 3040 408
rect 3034 406 3035 407
rect 2980 404 3035 406
rect 2980 403 2981 404
rect 2974 402 2981 403
rect 3034 403 3035 404
rect 3039 403 3040 407
rect 3034 402 3040 403
rect 3086 407 3092 408
rect 3086 403 3087 407
rect 3091 403 3092 407
rect 3095 407 3096 411
rect 3100 410 3101 411
rect 3118 411 3124 412
rect 3118 410 3119 411
rect 3100 408 3119 410
rect 3100 407 3101 408
rect 3095 406 3101 407
rect 3118 407 3119 408
rect 3123 407 3124 411
rect 3118 406 3124 407
rect 3190 411 3196 412
rect 3190 407 3191 411
rect 3195 407 3196 411
rect 3190 406 3196 407
rect 3086 402 3092 403
rect 1566 399 1572 400
rect 2150 385 2156 386
rect 646 384 652 385
rect 646 380 647 384
rect 651 380 652 384
rect 646 379 652 380
rect 806 384 812 385
rect 806 380 807 384
rect 811 380 812 384
rect 806 379 812 380
rect 950 384 956 385
rect 950 380 951 384
rect 955 380 956 384
rect 950 379 956 380
rect 1086 384 1092 385
rect 1086 380 1087 384
rect 1091 380 1092 384
rect 1086 379 1092 380
rect 1214 384 1220 385
rect 1214 380 1215 384
rect 1219 380 1220 384
rect 1214 379 1220 380
rect 1334 384 1340 385
rect 1334 380 1335 384
rect 1339 380 1340 384
rect 1334 379 1340 380
rect 1462 384 1468 385
rect 1462 380 1463 384
rect 1467 380 1468 384
rect 1462 379 1468 380
rect 1670 381 1676 382
rect 110 377 116 378
rect 110 373 111 377
rect 115 373 116 377
rect 110 372 116 373
rect 1630 377 1636 378
rect 1630 373 1631 377
rect 1635 373 1636 377
rect 1670 377 1671 381
rect 1675 377 1676 381
rect 2150 381 2151 385
rect 2155 381 2156 385
rect 2150 380 2156 381
rect 2278 385 2284 386
rect 2278 381 2279 385
rect 2283 381 2284 385
rect 2278 380 2284 381
rect 2406 385 2412 386
rect 2406 381 2407 385
rect 2411 381 2412 385
rect 2406 380 2412 381
rect 2534 385 2540 386
rect 2534 381 2535 385
rect 2539 381 2540 385
rect 2534 380 2540 381
rect 2662 385 2668 386
rect 2662 381 2663 385
rect 2667 381 2668 385
rect 2790 385 2796 386
rect 2662 380 2668 381
rect 2670 383 2677 384
rect 1670 376 1676 377
rect 2159 379 2165 380
rect 2159 375 2160 379
rect 2164 378 2165 379
rect 2258 379 2264 380
rect 2258 378 2259 379
rect 2164 376 2259 378
rect 2164 375 2165 376
rect 2159 374 2165 375
rect 2258 375 2259 376
rect 2263 378 2264 379
rect 2287 379 2293 380
rect 2287 378 2288 379
rect 2263 376 2288 378
rect 2263 375 2264 376
rect 2258 374 2264 375
rect 2287 375 2288 376
rect 2292 378 2293 379
rect 2386 379 2392 380
rect 2386 378 2387 379
rect 2292 376 2387 378
rect 2292 375 2293 376
rect 2287 374 2293 375
rect 2386 375 2387 376
rect 2391 378 2392 379
rect 2415 379 2421 380
rect 2415 378 2416 379
rect 2391 376 2416 378
rect 2391 375 2392 376
rect 2386 374 2392 375
rect 2415 375 2416 376
rect 2420 378 2421 379
rect 2514 379 2520 380
rect 2514 378 2515 379
rect 2420 376 2515 378
rect 2420 375 2421 376
rect 2415 374 2421 375
rect 2514 375 2515 376
rect 2519 378 2520 379
rect 2543 379 2549 380
rect 2543 378 2544 379
rect 2519 376 2544 378
rect 2519 375 2520 376
rect 2514 374 2520 375
rect 2543 375 2544 376
rect 2548 378 2549 379
rect 2574 379 2580 380
rect 2574 378 2575 379
rect 2548 376 2575 378
rect 2548 375 2549 376
rect 2543 374 2549 375
rect 2574 375 2575 376
rect 2579 375 2580 379
rect 2670 379 2671 383
rect 2676 382 2677 383
rect 2750 383 2756 384
rect 2750 382 2751 383
rect 2676 380 2751 382
rect 2676 379 2677 380
rect 2670 378 2677 379
rect 2750 379 2751 380
rect 2755 379 2756 383
rect 2790 381 2791 385
rect 2795 381 2796 385
rect 2918 385 2924 386
rect 2790 380 2796 381
rect 2798 383 2805 384
rect 2750 378 2756 379
rect 2798 379 2799 383
rect 2804 382 2805 383
rect 2862 383 2868 384
rect 2862 382 2863 383
rect 2804 380 2863 382
rect 2804 379 2805 380
rect 2798 378 2805 379
rect 2862 379 2863 380
rect 2867 379 2868 383
rect 2918 381 2919 385
rect 2923 381 2924 385
rect 3046 385 3052 386
rect 2918 380 2924 381
rect 2926 383 2933 384
rect 2862 378 2868 379
rect 2926 379 2927 383
rect 2932 382 2933 383
rect 2974 383 2980 384
rect 2974 382 2975 383
rect 2932 380 2975 382
rect 2932 379 2933 380
rect 2926 378 2933 379
rect 2974 379 2975 380
rect 2979 379 2980 383
rect 3046 381 3047 385
rect 3051 381 3052 385
rect 3046 380 3052 381
rect 3158 385 3164 386
rect 3158 381 3159 385
rect 3163 381 3164 385
rect 3158 380 3164 381
rect 3190 381 3196 382
rect 2974 378 2980 379
rect 3034 379 3040 380
rect 2574 374 2580 375
rect 3034 375 3035 379
rect 3039 378 3040 379
rect 3055 379 3061 380
rect 3055 378 3056 379
rect 3039 376 3056 378
rect 3039 375 3040 376
rect 3034 374 3040 375
rect 3055 375 3056 376
rect 3060 378 3061 379
rect 3118 379 3124 380
rect 3118 378 3119 379
rect 3060 376 3119 378
rect 3060 375 3061 376
rect 3055 374 3061 375
rect 3118 375 3119 376
rect 3123 378 3124 379
rect 3166 379 3173 380
rect 3166 378 3167 379
rect 3123 376 3167 378
rect 3123 375 3124 376
rect 3118 374 3124 375
rect 3166 375 3167 376
rect 3172 375 3173 379
rect 3190 377 3191 381
rect 3195 377 3196 381
rect 3190 376 3196 377
rect 3166 374 3173 375
rect 1630 372 1636 373
rect 1670 363 1676 364
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 654 359 661 360
rect 110 354 116 355
rect 646 355 652 356
rect 646 351 647 355
rect 651 351 652 355
rect 654 355 655 359
rect 660 355 661 359
rect 1470 359 1477 360
rect 654 354 661 355
rect 806 355 812 356
rect 646 350 652 351
rect 806 351 807 355
rect 811 351 812 355
rect 806 350 812 351
rect 814 355 821 356
rect 814 351 815 355
rect 820 351 821 355
rect 814 350 821 351
rect 950 355 956 356
rect 950 351 951 355
rect 955 351 956 355
rect 950 350 956 351
rect 959 355 965 356
rect 959 351 960 355
rect 964 354 965 355
rect 990 355 996 356
rect 990 354 991 355
rect 964 352 991 354
rect 964 351 965 352
rect 959 350 965 351
rect 990 351 991 352
rect 995 351 996 355
rect 990 350 996 351
rect 1086 355 1092 356
rect 1086 351 1087 355
rect 1091 351 1092 355
rect 1086 350 1092 351
rect 1095 355 1101 356
rect 1095 351 1096 355
rect 1100 354 1101 355
rect 1214 355 1220 356
rect 1100 352 1186 354
rect 1100 351 1101 352
rect 1095 350 1101 351
rect 542 341 548 342
rect 110 337 116 338
rect 110 333 111 337
rect 115 333 116 337
rect 542 337 543 341
rect 547 337 548 341
rect 542 336 548 337
rect 670 341 676 342
rect 670 337 671 341
rect 675 337 676 341
rect 670 336 676 337
rect 806 341 812 342
rect 806 337 807 341
rect 811 337 812 341
rect 806 336 812 337
rect 942 341 948 342
rect 942 337 943 341
rect 947 337 948 341
rect 942 336 948 337
rect 951 339 957 340
rect 110 332 116 333
rect 551 335 557 336
rect 551 331 552 335
rect 556 334 557 335
rect 630 335 636 336
rect 630 334 631 335
rect 556 332 631 334
rect 556 331 557 332
rect 551 330 557 331
rect 630 331 631 332
rect 635 334 636 335
rect 654 335 660 336
rect 654 334 655 335
rect 635 332 655 334
rect 635 331 636 332
rect 630 330 636 331
rect 654 331 655 332
rect 659 334 660 335
rect 679 335 685 336
rect 679 334 680 335
rect 659 332 680 334
rect 659 331 660 332
rect 654 330 660 331
rect 679 331 680 332
rect 684 331 685 335
rect 679 330 685 331
rect 814 335 821 336
rect 814 331 815 335
rect 820 334 821 335
rect 951 335 952 339
rect 956 338 957 339
rect 960 338 962 350
rect 956 336 962 338
rect 1078 341 1084 342
rect 1078 337 1079 341
rect 1083 337 1084 341
rect 1078 336 1084 337
rect 1087 339 1093 340
rect 956 335 957 336
rect 951 334 957 335
rect 1087 335 1088 339
rect 1092 338 1093 339
rect 1096 338 1098 350
rect 1184 346 1186 352
rect 1214 351 1215 355
rect 1219 351 1220 355
rect 1214 350 1220 351
rect 1223 355 1229 356
rect 1223 351 1224 355
rect 1228 354 1229 355
rect 1334 355 1340 356
rect 1228 352 1234 354
rect 1228 351 1229 352
rect 1223 350 1229 351
rect 1232 346 1234 352
rect 1334 351 1335 355
rect 1339 351 1340 355
rect 1334 350 1340 351
rect 1342 355 1349 356
rect 1342 351 1343 355
rect 1348 354 1349 355
rect 1462 355 1468 356
rect 1348 352 1378 354
rect 1348 351 1349 352
rect 1342 350 1349 351
rect 1184 344 1234 346
rect 1092 336 1098 338
rect 1222 341 1228 342
rect 1222 337 1223 341
rect 1227 337 1228 341
rect 1232 340 1234 344
rect 1366 341 1372 342
rect 1222 336 1228 337
rect 1231 339 1237 340
rect 1092 335 1093 336
rect 1087 334 1093 335
rect 1231 335 1232 339
rect 1236 338 1237 339
rect 1294 339 1300 340
rect 1294 338 1295 339
rect 1236 336 1295 338
rect 1236 335 1237 336
rect 1231 334 1237 335
rect 1294 335 1295 336
rect 1299 338 1300 339
rect 1342 339 1348 340
rect 1342 338 1343 339
rect 1299 336 1343 338
rect 1299 335 1300 336
rect 1294 334 1300 335
rect 1342 335 1343 336
rect 1347 335 1348 339
rect 1366 337 1367 341
rect 1371 337 1372 341
rect 1376 340 1378 352
rect 1462 351 1463 355
rect 1467 351 1468 355
rect 1470 355 1471 359
rect 1476 355 1477 359
rect 1470 354 1477 355
rect 1630 359 1636 360
rect 1630 355 1631 359
rect 1635 355 1636 359
rect 1670 359 1671 363
rect 1675 359 1676 363
rect 1670 358 1676 359
rect 3190 363 3196 364
rect 3190 359 3191 363
rect 3195 359 3196 363
rect 3190 358 3196 359
rect 1630 354 1636 355
rect 2150 356 2156 357
rect 2150 352 2151 356
rect 2155 352 2156 356
rect 2150 351 2156 352
rect 2278 356 2284 357
rect 2278 352 2279 356
rect 2283 352 2284 356
rect 2278 351 2284 352
rect 2406 356 2412 357
rect 2406 352 2407 356
rect 2411 352 2412 356
rect 2406 351 2412 352
rect 2534 356 2540 357
rect 2534 352 2535 356
rect 2539 352 2540 356
rect 2534 351 2540 352
rect 2662 356 2668 357
rect 2662 352 2663 356
rect 2667 352 2668 356
rect 2662 351 2668 352
rect 2790 356 2796 357
rect 2790 352 2791 356
rect 2795 352 2796 356
rect 2790 351 2796 352
rect 2918 356 2924 357
rect 2918 352 2919 356
rect 2923 352 2924 356
rect 2918 351 2924 352
rect 3046 356 3052 357
rect 3046 352 3047 356
rect 3051 352 3052 356
rect 3046 351 3052 352
rect 3158 356 3164 357
rect 3158 352 3159 356
rect 3163 352 3164 356
rect 3158 351 3164 352
rect 1462 350 1468 351
rect 1366 336 1372 337
rect 1375 339 1381 340
rect 1342 334 1348 335
rect 1375 335 1376 339
rect 1380 338 1381 339
rect 1470 339 1476 340
rect 1470 338 1471 339
rect 1380 336 1471 338
rect 1380 335 1381 336
rect 1375 334 1381 335
rect 1470 335 1471 336
rect 1475 335 1476 339
rect 1470 334 1476 335
rect 1630 337 1636 338
rect 820 332 954 334
rect 1630 333 1631 337
rect 1635 333 1636 337
rect 1630 332 1636 333
rect 2046 332 2052 333
rect 820 331 821 332
rect 814 330 821 331
rect 2046 328 2047 332
rect 2051 328 2052 332
rect 2046 327 2052 328
rect 2174 332 2180 333
rect 2174 328 2175 332
rect 2179 328 2180 332
rect 2174 327 2180 328
rect 2302 332 2308 333
rect 2302 328 2303 332
rect 2307 328 2308 332
rect 2302 327 2308 328
rect 2430 332 2436 333
rect 2430 328 2431 332
rect 2435 328 2436 332
rect 2430 327 2436 328
rect 2566 332 2572 333
rect 2566 328 2567 332
rect 2571 328 2572 332
rect 2566 327 2572 328
rect 2710 332 2716 333
rect 2710 328 2711 332
rect 2715 328 2716 332
rect 2710 327 2716 328
rect 2862 332 2868 333
rect 2862 328 2863 332
rect 2867 328 2868 332
rect 2862 327 2868 328
rect 3022 332 3028 333
rect 3022 328 3023 332
rect 3027 328 3028 332
rect 3022 327 3028 328
rect 3158 332 3164 333
rect 3158 328 3159 332
rect 3163 328 3164 332
rect 3158 327 3164 328
rect 1670 325 1676 326
rect 1670 321 1671 325
rect 1675 321 1676 325
rect 1670 320 1676 321
rect 3190 325 3196 326
rect 3190 321 3191 325
rect 3195 321 3196 325
rect 3190 320 3196 321
rect 110 319 116 320
rect 110 315 111 319
rect 115 315 116 319
rect 110 314 116 315
rect 1630 319 1636 320
rect 1630 315 1631 319
rect 1635 315 1636 319
rect 1630 314 1636 315
rect 542 312 548 313
rect 542 308 543 312
rect 547 308 548 312
rect 542 307 548 308
rect 670 312 676 313
rect 670 308 671 312
rect 675 308 676 312
rect 670 307 676 308
rect 806 312 812 313
rect 806 308 807 312
rect 811 308 812 312
rect 806 307 812 308
rect 942 312 948 313
rect 942 308 943 312
rect 947 308 948 312
rect 942 307 948 308
rect 1078 312 1084 313
rect 1078 308 1079 312
rect 1083 308 1084 312
rect 1078 307 1084 308
rect 1222 312 1228 313
rect 1222 308 1223 312
rect 1227 308 1228 312
rect 1222 307 1228 308
rect 1366 312 1372 313
rect 1366 308 1367 312
rect 1371 308 1372 312
rect 1366 307 1372 308
rect 1670 307 1676 308
rect 1670 303 1671 307
rect 1675 303 1676 307
rect 2439 307 2445 308
rect 1670 302 1676 303
rect 2046 303 2052 304
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 2046 298 2052 299
rect 2055 303 2064 304
rect 2055 299 2056 303
rect 2063 299 2064 303
rect 2055 298 2064 299
rect 2174 303 2180 304
rect 2174 299 2175 303
rect 2179 299 2180 303
rect 2174 298 2180 299
rect 2183 303 2192 304
rect 2183 299 2184 303
rect 2191 299 2192 303
rect 2183 298 2192 299
rect 2302 303 2308 304
rect 2302 299 2303 303
rect 2307 299 2308 303
rect 2302 298 2308 299
rect 2311 303 2317 304
rect 2311 299 2312 303
rect 2316 302 2317 303
rect 2326 303 2332 304
rect 2326 302 2327 303
rect 2316 300 2327 302
rect 2316 299 2317 300
rect 2311 298 2317 299
rect 2326 299 2327 300
rect 2331 299 2332 303
rect 2326 298 2332 299
rect 2430 303 2436 304
rect 2430 299 2431 303
rect 2435 299 2436 303
rect 2439 303 2440 307
rect 2444 303 2445 307
rect 2870 307 2877 308
rect 2439 302 2445 303
rect 2566 303 2572 304
rect 2430 298 2436 299
rect 2566 299 2567 303
rect 2571 299 2572 303
rect 2566 298 2572 299
rect 2574 303 2581 304
rect 2574 299 2575 303
rect 2580 302 2581 303
rect 2670 303 2676 304
rect 2670 302 2671 303
rect 2580 300 2671 302
rect 2580 299 2581 300
rect 2574 298 2581 299
rect 2670 299 2671 300
rect 2675 299 2676 303
rect 2670 298 2676 299
rect 2710 303 2716 304
rect 2710 299 2711 303
rect 2715 299 2716 303
rect 2710 298 2716 299
rect 2718 303 2725 304
rect 2718 299 2719 303
rect 2724 302 2725 303
rect 2790 303 2796 304
rect 2790 302 2791 303
rect 2724 300 2791 302
rect 2724 299 2725 300
rect 2718 298 2725 299
rect 2790 299 2791 300
rect 2795 299 2796 303
rect 2790 298 2796 299
rect 2862 303 2868 304
rect 2862 299 2863 303
rect 2867 299 2868 303
rect 2870 303 2871 307
rect 2876 306 2877 307
rect 2926 307 2932 308
rect 2926 306 2927 307
rect 2876 304 2927 306
rect 2876 303 2877 304
rect 2870 302 2877 303
rect 2926 303 2927 304
rect 2931 303 2932 307
rect 3031 307 3040 308
rect 2926 302 2932 303
rect 3022 303 3028 304
rect 2862 298 2868 299
rect 3022 299 3023 303
rect 3027 299 3028 303
rect 3031 303 3032 307
rect 3039 303 3040 307
rect 3166 307 3173 308
rect 3031 302 3040 303
rect 3158 303 3164 304
rect 3022 298 3028 299
rect 3158 299 3159 303
rect 3163 299 3164 303
rect 3166 303 3167 307
rect 3172 303 3173 307
rect 3166 302 3173 303
rect 3190 307 3196 308
rect 3190 303 3191 307
rect 3195 303 3196 307
rect 3190 302 3196 303
rect 3158 298 3164 299
rect 462 296 468 297
rect 462 292 463 296
rect 467 292 468 296
rect 462 291 468 292
rect 622 296 628 297
rect 622 292 623 296
rect 627 292 628 296
rect 622 291 628 292
rect 766 296 772 297
rect 766 292 767 296
rect 771 292 772 296
rect 766 291 772 292
rect 902 296 908 297
rect 902 292 903 296
rect 907 292 908 296
rect 902 291 908 292
rect 1030 296 1036 297
rect 1030 292 1031 296
rect 1035 292 1036 296
rect 1030 291 1036 292
rect 1158 296 1164 297
rect 1158 292 1159 296
rect 1163 292 1164 296
rect 1158 291 1164 292
rect 1286 296 1292 297
rect 1286 292 1287 296
rect 1291 292 1292 296
rect 1286 291 1292 292
rect 110 289 116 290
rect 110 285 111 289
rect 115 285 116 289
rect 110 284 116 285
rect 1630 289 1636 290
rect 1630 285 1631 289
rect 1635 285 1636 289
rect 1630 284 1636 285
rect 1942 285 1948 286
rect 1670 281 1676 282
rect 1670 277 1671 281
rect 1675 277 1676 281
rect 1942 281 1943 285
rect 1947 281 1948 285
rect 1942 280 1948 281
rect 2070 285 2076 286
rect 2070 281 2071 285
rect 2075 281 2076 285
rect 2070 280 2076 281
rect 2198 285 2204 286
rect 2198 281 2199 285
rect 2203 281 2204 285
rect 2198 280 2204 281
rect 2318 285 2324 286
rect 2318 281 2319 285
rect 2323 281 2324 285
rect 2318 280 2324 281
rect 2438 285 2444 286
rect 2438 281 2439 285
rect 2443 281 2444 285
rect 2438 280 2444 281
rect 2550 285 2556 286
rect 2550 281 2551 285
rect 2555 281 2556 285
rect 2662 285 2668 286
rect 2550 280 2556 281
rect 2559 283 2565 284
rect 1670 276 1676 277
rect 1951 279 1957 280
rect 1951 275 1952 279
rect 1956 278 1957 279
rect 2058 279 2064 280
rect 2058 278 2059 279
rect 1956 276 2059 278
rect 1956 275 1957 276
rect 1951 274 1957 275
rect 2058 275 2059 276
rect 2063 278 2064 279
rect 2079 279 2085 280
rect 2079 278 2080 279
rect 2063 276 2080 278
rect 2063 275 2064 276
rect 2058 274 2064 275
rect 2079 275 2080 276
rect 2084 278 2085 279
rect 2186 279 2192 280
rect 2186 278 2187 279
rect 2084 276 2187 278
rect 2084 275 2085 276
rect 2079 274 2085 275
rect 2186 275 2187 276
rect 2191 278 2192 279
rect 2207 279 2213 280
rect 2207 278 2208 279
rect 2191 276 2208 278
rect 2191 275 2192 276
rect 2186 274 2192 275
rect 2207 275 2208 276
rect 2212 278 2213 279
rect 2326 279 2333 280
rect 2326 278 2327 279
rect 2212 276 2327 278
rect 2212 275 2213 276
rect 2207 274 2213 275
rect 2326 275 2327 276
rect 2332 278 2333 279
rect 2446 279 2453 280
rect 2446 278 2447 279
rect 2332 276 2447 278
rect 2332 275 2333 276
rect 2326 274 2333 275
rect 2446 275 2447 276
rect 2452 278 2453 279
rect 2526 279 2532 280
rect 2526 278 2527 279
rect 2452 276 2527 278
rect 2452 275 2453 276
rect 2446 274 2453 275
rect 2526 275 2527 276
rect 2531 278 2532 279
rect 2559 279 2560 283
rect 2564 282 2565 283
rect 2574 283 2580 284
rect 2574 282 2575 283
rect 2564 280 2575 282
rect 2564 279 2565 280
rect 2559 278 2565 279
rect 2574 279 2575 280
rect 2579 279 2580 283
rect 2662 281 2663 285
rect 2667 281 2668 285
rect 2782 285 2788 286
rect 2662 280 2668 281
rect 2670 283 2677 284
rect 2574 278 2580 279
rect 2670 279 2671 283
rect 2676 282 2677 283
rect 2718 283 2724 284
rect 2718 282 2719 283
rect 2676 280 2719 282
rect 2676 279 2677 280
rect 2670 278 2677 279
rect 2718 279 2719 280
rect 2723 279 2724 283
rect 2782 281 2783 285
rect 2787 281 2788 285
rect 2782 280 2788 281
rect 2790 283 2797 284
rect 2718 278 2724 279
rect 2790 279 2791 283
rect 2796 282 2797 283
rect 2870 283 2876 284
rect 2870 282 2871 283
rect 2796 280 2871 282
rect 2796 279 2797 280
rect 2790 278 2797 279
rect 2870 279 2871 280
rect 2875 279 2876 283
rect 2870 278 2876 279
rect 3190 281 3196 282
rect 2531 276 2563 278
rect 3190 277 3191 281
rect 3195 277 3196 281
rect 3190 276 3196 277
rect 2531 275 2532 276
rect 2526 274 2532 275
rect 110 271 116 272
rect 110 267 111 271
rect 115 267 116 271
rect 470 271 477 272
rect 110 266 116 267
rect 462 267 468 268
rect 462 263 463 267
rect 467 263 468 267
rect 470 267 471 271
rect 476 267 477 271
rect 774 271 781 272
rect 470 266 477 267
rect 622 267 628 268
rect 462 262 468 263
rect 622 263 623 267
rect 627 263 628 267
rect 622 262 628 263
rect 630 267 637 268
rect 630 263 631 267
rect 636 263 637 267
rect 630 262 637 263
rect 766 267 772 268
rect 766 263 767 267
rect 771 263 772 267
rect 774 267 775 271
rect 780 270 781 271
rect 814 271 820 272
rect 814 270 815 271
rect 780 268 815 270
rect 780 267 781 268
rect 774 266 781 267
rect 814 267 815 268
rect 819 267 820 271
rect 1294 271 1301 272
rect 814 266 820 267
rect 902 267 908 268
rect 766 262 772 263
rect 902 263 903 267
rect 907 263 908 267
rect 902 262 908 263
rect 911 267 917 268
rect 911 263 912 267
rect 916 263 917 267
rect 911 262 917 263
rect 1030 267 1036 268
rect 1030 263 1031 267
rect 1035 263 1036 267
rect 1030 262 1036 263
rect 1039 267 1045 268
rect 1039 263 1040 267
rect 1044 263 1045 267
rect 1039 262 1045 263
rect 1158 267 1164 268
rect 1158 263 1159 267
rect 1163 263 1164 267
rect 1158 262 1164 263
rect 1167 267 1173 268
rect 1167 263 1168 267
rect 1172 266 1173 267
rect 1286 267 1292 268
rect 1172 264 1194 266
rect 1172 263 1173 264
rect 1167 262 1173 263
rect 912 258 914 262
rect 1040 258 1042 262
rect 912 256 1050 258
rect 358 253 364 254
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 358 249 359 253
rect 363 249 364 253
rect 486 253 492 254
rect 358 248 364 249
rect 366 251 373 252
rect 366 247 367 251
rect 372 250 373 251
rect 470 251 476 252
rect 470 250 471 251
rect 372 248 471 250
rect 372 247 373 248
rect 366 246 373 247
rect 470 247 471 248
rect 475 247 476 251
rect 486 249 487 253
rect 491 249 492 253
rect 486 248 492 249
rect 622 253 628 254
rect 622 249 623 253
rect 627 249 628 253
rect 622 248 628 249
rect 758 253 764 254
rect 758 249 759 253
rect 763 249 764 253
rect 894 253 900 254
rect 758 248 764 249
rect 767 249 773 250
rect 470 246 476 247
rect 495 247 501 248
rect 495 246 496 247
rect 110 244 116 245
rect 472 244 496 246
rect 495 243 496 244
rect 500 246 501 247
rect 630 247 637 248
rect 630 246 631 247
rect 500 244 631 246
rect 500 243 501 244
rect 495 242 501 243
rect 630 243 631 244
rect 636 243 637 247
rect 767 245 768 249
rect 772 245 773 249
rect 894 249 895 253
rect 899 249 900 253
rect 894 248 900 249
rect 903 251 909 252
rect 903 248 904 251
rect 767 244 773 245
rect 902 247 904 248
rect 908 250 909 251
rect 912 250 914 256
rect 908 248 914 250
rect 1038 253 1044 254
rect 1038 249 1039 253
rect 1043 249 1044 253
rect 1038 248 1044 249
rect 1048 248 1050 256
rect 1182 253 1188 254
rect 1182 249 1183 253
rect 1187 249 1188 253
rect 1192 252 1194 264
rect 1286 263 1287 267
rect 1291 263 1292 267
rect 1294 267 1295 271
rect 1300 267 1301 271
rect 1294 266 1301 267
rect 1630 271 1636 272
rect 1630 267 1631 271
rect 1635 267 1636 271
rect 1630 266 1636 267
rect 1286 262 1292 263
rect 1670 263 1676 264
rect 1670 259 1671 263
rect 1675 259 1676 263
rect 1670 258 1676 259
rect 3190 263 3196 264
rect 3190 259 3191 263
rect 3195 259 3196 263
rect 3190 258 3196 259
rect 1942 256 1948 257
rect 1942 252 1943 256
rect 1947 252 1948 256
rect 1182 248 1188 249
rect 1191 251 1197 252
rect 908 247 909 248
rect 630 242 637 243
rect 766 243 772 244
rect 766 239 767 243
rect 771 239 772 243
rect 902 243 903 247
rect 907 246 909 247
rect 1047 247 1053 248
rect 907 243 908 246
rect 902 242 908 243
rect 1047 243 1048 247
rect 1052 246 1053 247
rect 1191 247 1192 251
rect 1196 250 1197 251
rect 1294 251 1300 252
rect 1942 251 1948 252
rect 2070 256 2076 257
rect 2070 252 2071 256
rect 2075 252 2076 256
rect 2070 251 2076 252
rect 2198 256 2204 257
rect 2198 252 2199 256
rect 2203 252 2204 256
rect 2198 251 2204 252
rect 2318 256 2324 257
rect 2318 252 2319 256
rect 2323 252 2324 256
rect 2318 251 2324 252
rect 2438 256 2444 257
rect 2438 252 2439 256
rect 2443 252 2444 256
rect 2438 251 2444 252
rect 2550 256 2556 257
rect 2550 252 2551 256
rect 2555 252 2556 256
rect 2550 251 2556 252
rect 2662 256 2668 257
rect 2662 252 2663 256
rect 2667 252 2668 256
rect 2662 251 2668 252
rect 2782 256 2788 257
rect 2782 252 2783 256
rect 2787 252 2788 256
rect 2782 251 2788 252
rect 1294 250 1295 251
rect 1196 248 1295 250
rect 1196 247 1197 248
rect 1191 246 1197 247
rect 1294 247 1295 248
rect 1299 247 1300 251
rect 1294 246 1300 247
rect 1630 249 1636 250
rect 1052 244 1194 246
rect 1630 245 1631 249
rect 1635 245 1636 249
rect 1630 244 1636 245
rect 1052 243 1053 244
rect 1047 242 1053 243
rect 766 238 772 239
rect 1846 232 1852 233
rect 110 231 116 232
rect 110 227 111 231
rect 115 227 116 231
rect 110 226 116 227
rect 1630 231 1636 232
rect 1630 227 1631 231
rect 1635 227 1636 231
rect 1846 228 1847 232
rect 1851 228 1852 232
rect 1846 227 1852 228
rect 1974 232 1980 233
rect 1974 228 1975 232
rect 1979 228 1980 232
rect 1974 227 1980 228
rect 2102 232 2108 233
rect 2102 228 2103 232
rect 2107 228 2108 232
rect 2102 227 2108 228
rect 2246 232 2252 233
rect 2246 228 2247 232
rect 2251 228 2252 232
rect 2246 227 2252 228
rect 2406 232 2412 233
rect 2406 228 2407 232
rect 2411 228 2412 232
rect 2406 227 2412 228
rect 2582 232 2588 233
rect 2582 228 2583 232
rect 2587 228 2588 232
rect 2582 227 2588 228
rect 2766 232 2772 233
rect 2766 228 2767 232
rect 2771 228 2772 232
rect 2766 227 2772 228
rect 2966 232 2972 233
rect 2966 228 2967 232
rect 2971 228 2972 232
rect 2966 227 2972 228
rect 3158 232 3164 233
rect 3158 228 3159 232
rect 3163 228 3164 232
rect 3158 227 3164 228
rect 1630 226 1636 227
rect 1670 225 1676 226
rect 358 224 364 225
rect 358 220 359 224
rect 363 220 364 224
rect 358 219 364 220
rect 486 224 492 225
rect 486 220 487 224
rect 491 220 492 224
rect 486 219 492 220
rect 622 224 628 225
rect 622 220 623 224
rect 627 220 628 224
rect 622 219 628 220
rect 758 224 764 225
rect 758 220 759 224
rect 763 220 764 224
rect 758 219 764 220
rect 894 224 900 225
rect 894 220 895 224
rect 899 220 900 224
rect 894 219 900 220
rect 1038 224 1044 225
rect 1038 220 1039 224
rect 1043 220 1044 224
rect 1038 219 1044 220
rect 1182 224 1188 225
rect 1182 220 1183 224
rect 1187 220 1188 224
rect 1670 221 1671 225
rect 1675 221 1676 225
rect 1670 220 1676 221
rect 3190 225 3196 226
rect 3190 221 3191 225
rect 3195 221 3196 225
rect 3190 220 3196 221
rect 1182 219 1188 220
rect 2926 211 2932 212
rect 278 208 284 209
rect 278 204 279 208
rect 283 204 284 208
rect 278 203 284 204
rect 446 208 452 209
rect 446 204 447 208
rect 451 204 452 208
rect 446 203 452 204
rect 614 208 620 209
rect 614 204 615 208
rect 619 204 620 208
rect 614 203 620 204
rect 774 208 780 209
rect 774 204 775 208
rect 779 204 780 208
rect 774 203 780 204
rect 942 208 948 209
rect 942 204 943 208
rect 947 204 948 208
rect 942 203 948 204
rect 1110 208 1116 209
rect 1110 204 1111 208
rect 1115 204 1116 208
rect 1110 203 1116 204
rect 1670 207 1676 208
rect 1670 203 1671 207
rect 1675 203 1676 207
rect 2775 207 2781 208
rect 1670 202 1676 203
rect 1846 203 1852 204
rect 110 201 116 202
rect 110 197 111 201
rect 115 197 116 201
rect 110 196 116 197
rect 1630 201 1636 202
rect 1630 197 1631 201
rect 1635 197 1636 201
rect 1846 199 1847 203
rect 1851 199 1852 203
rect 1846 198 1852 199
rect 1854 203 1861 204
rect 1854 199 1855 203
rect 1860 199 1861 203
rect 1854 198 1861 199
rect 1974 203 1980 204
rect 1974 199 1975 203
rect 1979 199 1980 203
rect 1974 198 1980 199
rect 1982 203 1989 204
rect 1982 199 1983 203
rect 1988 199 1989 203
rect 1982 198 1989 199
rect 2102 203 2108 204
rect 2102 199 2103 203
rect 2107 199 2108 203
rect 2102 198 2108 199
rect 2110 203 2117 204
rect 2110 199 2111 203
rect 2116 199 2117 203
rect 2110 198 2117 199
rect 2246 203 2252 204
rect 2246 199 2247 203
rect 2251 199 2252 203
rect 2246 198 2252 199
rect 2254 203 2261 204
rect 2254 199 2255 203
rect 2260 202 2261 203
rect 2318 203 2324 204
rect 2318 202 2319 203
rect 2260 200 2319 202
rect 2260 199 2261 200
rect 2254 198 2261 199
rect 2318 199 2319 200
rect 2323 199 2324 203
rect 2318 198 2324 199
rect 2406 203 2412 204
rect 2406 199 2407 203
rect 2411 199 2412 203
rect 2406 198 2412 199
rect 2414 203 2421 204
rect 2414 199 2415 203
rect 2420 202 2421 203
rect 2502 203 2508 204
rect 2502 202 2503 203
rect 2420 200 2503 202
rect 2420 199 2421 200
rect 2414 198 2421 199
rect 2502 199 2503 200
rect 2507 199 2508 203
rect 2502 198 2508 199
rect 2582 203 2588 204
rect 2582 199 2583 203
rect 2587 199 2588 203
rect 2582 198 2588 199
rect 2590 203 2597 204
rect 2590 199 2591 203
rect 2596 199 2597 203
rect 2590 198 2597 199
rect 2766 203 2772 204
rect 2766 199 2767 203
rect 2771 199 2772 203
rect 2775 203 2776 207
rect 2780 206 2781 207
rect 2790 207 2796 208
rect 2790 206 2791 207
rect 2780 204 2791 206
rect 2780 203 2781 204
rect 2775 202 2781 203
rect 2790 203 2791 204
rect 2795 203 2796 207
rect 2926 207 2927 211
rect 2931 210 2932 211
rect 2931 208 2979 210
rect 2931 207 2932 208
rect 2926 206 2932 207
rect 2975 207 2981 208
rect 2790 202 2796 203
rect 2966 203 2972 204
rect 2766 198 2772 199
rect 2966 199 2967 203
rect 2971 199 2972 203
rect 2975 203 2976 207
rect 2980 203 2981 207
rect 3166 207 3173 208
rect 2975 202 2981 203
rect 3158 203 3164 204
rect 2966 198 2972 199
rect 3158 199 3159 203
rect 3163 199 3164 203
rect 3166 203 3167 207
rect 3172 203 3173 207
rect 3166 202 3173 203
rect 3190 207 3196 208
rect 3190 203 3191 207
rect 3195 203 3196 207
rect 3190 202 3196 203
rect 3158 198 3164 199
rect 1630 196 1636 197
rect 902 187 908 188
rect 110 183 116 184
rect 110 179 111 183
rect 115 179 116 183
rect 287 183 293 184
rect 110 178 116 179
rect 278 179 284 180
rect 278 175 279 179
rect 283 175 284 179
rect 287 179 288 183
rect 292 182 293 183
rect 366 183 372 184
rect 366 182 367 183
rect 292 180 367 182
rect 292 179 293 180
rect 287 178 293 179
rect 366 179 367 180
rect 371 179 372 183
rect 455 183 461 184
rect 366 178 372 179
rect 446 179 452 180
rect 278 174 284 175
rect 198 169 204 170
rect 110 165 116 166
rect 110 161 111 165
rect 115 161 116 165
rect 198 165 199 169
rect 203 165 204 169
rect 198 164 204 165
rect 207 167 213 168
rect 110 160 116 161
rect 146 163 152 164
rect 146 159 147 163
rect 151 162 152 163
rect 207 163 208 167
rect 212 166 213 167
rect 289 166 291 178
rect 368 176 379 178
rect 212 164 291 166
rect 366 169 372 170
rect 366 165 367 169
rect 371 165 372 169
rect 377 168 379 176
rect 446 175 447 179
rect 451 175 452 179
rect 455 179 456 183
rect 460 182 461 183
rect 470 183 476 184
rect 470 182 471 183
rect 460 180 471 182
rect 460 179 461 180
rect 455 178 461 179
rect 470 179 471 180
rect 475 179 476 183
rect 902 183 903 187
rect 907 186 908 187
rect 907 184 955 186
rect 907 183 908 184
rect 902 182 908 183
rect 951 183 957 184
rect 470 178 476 179
rect 614 179 620 180
rect 446 174 452 175
rect 614 175 615 179
rect 619 175 620 179
rect 614 174 620 175
rect 623 179 629 180
rect 623 175 624 179
rect 628 175 629 179
rect 623 174 629 175
rect 774 179 780 180
rect 774 175 775 179
rect 779 175 780 179
rect 774 174 780 175
rect 783 179 789 180
rect 783 175 784 179
rect 788 175 789 179
rect 783 174 789 175
rect 942 179 948 180
rect 942 175 943 179
rect 947 175 948 179
rect 951 179 952 183
rect 956 179 957 183
rect 1630 183 1636 184
rect 951 178 957 179
rect 1110 179 1116 180
rect 942 174 948 175
rect 1110 175 1111 179
rect 1115 175 1116 179
rect 1110 174 1116 175
rect 1119 179 1125 180
rect 1119 175 1120 179
rect 1124 175 1125 179
rect 1630 179 1631 183
rect 1635 179 1636 183
rect 1630 178 1636 179
rect 1742 181 1748 182
rect 1119 174 1125 175
rect 1670 177 1676 178
rect 534 169 540 170
rect 366 164 372 165
rect 375 167 381 168
rect 212 163 213 164
rect 207 162 213 163
rect 375 163 376 167
rect 380 163 381 167
rect 534 165 535 169
rect 539 165 540 169
rect 534 164 540 165
rect 694 169 700 170
rect 694 165 695 169
rect 699 165 700 169
rect 694 164 700 165
rect 375 162 381 163
rect 470 163 476 164
rect 151 160 211 162
rect 151 159 152 160
rect 146 158 152 159
rect 470 159 471 163
rect 475 162 476 163
rect 543 163 552 164
rect 543 162 544 163
rect 475 160 544 162
rect 475 159 476 160
rect 470 158 476 159
rect 543 159 544 160
rect 551 159 552 163
rect 543 158 552 159
rect 702 163 709 164
rect 702 159 703 163
rect 708 162 709 163
rect 766 163 772 164
rect 766 162 767 163
rect 708 160 767 162
rect 708 159 709 160
rect 702 158 709 159
rect 766 159 767 160
rect 771 162 772 163
rect 784 162 786 174
rect 862 169 868 170
rect 862 165 863 169
rect 867 165 868 169
rect 862 164 868 165
rect 1030 169 1036 170
rect 1030 165 1031 169
rect 1035 165 1036 169
rect 1030 164 1036 165
rect 1039 167 1045 168
rect 871 163 877 164
rect 871 162 872 163
rect 771 160 872 162
rect 771 159 772 160
rect 766 158 772 159
rect 871 159 872 160
rect 876 162 877 163
rect 902 163 908 164
rect 902 162 903 163
rect 876 160 903 162
rect 876 159 877 160
rect 871 158 877 159
rect 902 159 903 160
rect 907 159 908 163
rect 902 158 908 159
rect 1022 163 1028 164
rect 1022 159 1023 163
rect 1027 162 1028 163
rect 1039 163 1040 167
rect 1044 166 1045 167
rect 1120 166 1122 174
rect 1670 173 1671 177
rect 1675 173 1676 177
rect 1742 177 1743 181
rect 1747 177 1748 181
rect 1742 176 1748 177
rect 1870 181 1876 182
rect 1870 177 1871 181
rect 1875 177 1876 181
rect 1870 176 1876 177
rect 1998 181 2004 182
rect 1998 177 1999 181
rect 2003 177 2004 181
rect 1998 176 2004 177
rect 2142 181 2148 182
rect 2142 177 2143 181
rect 2147 177 2148 181
rect 2310 181 2316 182
rect 2142 176 2148 177
rect 2151 179 2157 180
rect 1670 172 1676 173
rect 1750 175 1757 176
rect 1750 171 1751 175
rect 1756 174 1757 175
rect 1854 175 1860 176
rect 1854 174 1855 175
rect 1756 172 1855 174
rect 1756 171 1757 172
rect 1750 170 1757 171
rect 1854 171 1855 172
rect 1859 174 1860 175
rect 1879 175 1885 176
rect 1879 174 1880 175
rect 1859 172 1880 174
rect 1859 171 1860 172
rect 1854 170 1860 171
rect 1879 171 1880 172
rect 1884 174 1885 175
rect 1982 175 1988 176
rect 1982 174 1983 175
rect 1884 172 1983 174
rect 1884 171 1885 172
rect 1879 170 1885 171
rect 1982 171 1983 172
rect 1987 174 1988 175
rect 2007 175 2013 176
rect 2007 174 2008 175
rect 1987 172 2008 174
rect 1987 171 1988 172
rect 1982 170 1988 171
rect 2007 171 2008 172
rect 2012 174 2013 175
rect 2110 175 2116 176
rect 2110 174 2111 175
rect 2012 172 2111 174
rect 2012 171 2013 172
rect 2007 170 2013 171
rect 2110 171 2111 172
rect 2115 174 2116 175
rect 2151 175 2152 179
rect 2156 178 2157 179
rect 2254 179 2260 180
rect 2254 178 2255 179
rect 2156 176 2255 178
rect 2156 175 2157 176
rect 2151 174 2157 175
rect 2254 175 2255 176
rect 2259 175 2260 179
rect 2310 177 2311 181
rect 2315 177 2316 181
rect 2494 181 2500 182
rect 2310 176 2316 177
rect 2318 179 2325 180
rect 2254 174 2260 175
rect 2318 175 2319 179
rect 2324 178 2325 179
rect 2358 179 2364 180
rect 2358 178 2359 179
rect 2324 176 2359 178
rect 2324 175 2325 176
rect 2318 174 2325 175
rect 2358 175 2359 176
rect 2363 178 2364 179
rect 2414 179 2420 180
rect 2414 178 2415 179
rect 2363 176 2415 178
rect 2363 175 2364 176
rect 2358 174 2364 175
rect 2414 175 2415 176
rect 2419 175 2420 179
rect 2494 177 2495 181
rect 2499 177 2500 181
rect 2702 181 2708 182
rect 2494 176 2500 177
rect 2502 179 2509 180
rect 2414 174 2420 175
rect 2502 175 2503 179
rect 2508 178 2509 179
rect 2590 179 2596 180
rect 2590 178 2591 179
rect 2508 176 2591 178
rect 2508 175 2509 176
rect 2502 174 2509 175
rect 2590 175 2591 176
rect 2595 175 2596 179
rect 2702 177 2703 181
rect 2707 177 2708 181
rect 2918 181 2924 182
rect 2714 179 2720 180
rect 2714 178 2715 179
rect 2702 176 2708 177
rect 2711 177 2715 178
rect 2590 174 2596 175
rect 2115 172 2155 174
rect 2711 173 2712 177
rect 2719 175 2720 179
rect 2918 177 2919 181
rect 2923 177 2924 181
rect 3134 181 3140 182
rect 2918 176 2924 177
rect 2926 179 2933 180
rect 2716 174 2720 175
rect 2926 175 2927 179
rect 2932 175 2933 179
rect 3134 177 3135 181
rect 3139 177 3140 181
rect 3134 176 3140 177
rect 3142 179 3149 180
rect 2926 174 2933 175
rect 3142 175 3143 179
rect 3148 178 3149 179
rect 3166 179 3172 180
rect 3166 178 3167 179
rect 3148 176 3167 178
rect 3148 175 3149 176
rect 3142 174 3149 175
rect 3166 175 3167 176
rect 3171 175 3172 179
rect 3166 174 3172 175
rect 3190 177 3196 178
rect 2716 173 2717 174
rect 2711 172 2717 173
rect 3190 173 3191 177
rect 3195 173 3196 177
rect 3190 172 3196 173
rect 2115 171 2116 172
rect 2110 170 2116 171
rect 1044 164 1122 166
rect 1630 165 1636 166
rect 1044 163 1045 164
rect 1039 162 1045 163
rect 1027 160 1041 162
rect 1630 161 1631 165
rect 1635 161 1636 165
rect 1630 160 1636 161
rect 1027 159 1028 160
rect 1022 158 1028 159
rect 1670 159 1676 160
rect 1670 155 1671 159
rect 1675 155 1676 159
rect 1670 154 1676 155
rect 3190 159 3196 160
rect 3190 155 3191 159
rect 3195 155 3196 159
rect 3190 154 3196 155
rect 1742 152 1748 153
rect 1742 148 1743 152
rect 1747 148 1748 152
rect 110 147 116 148
rect 110 143 111 147
rect 115 143 116 147
rect 110 142 116 143
rect 1630 147 1636 148
rect 1742 147 1748 148
rect 1870 152 1876 153
rect 1870 148 1871 152
rect 1875 148 1876 152
rect 1870 147 1876 148
rect 1998 152 2004 153
rect 1998 148 1999 152
rect 2003 148 2004 152
rect 1998 147 2004 148
rect 2142 152 2148 153
rect 2142 148 2143 152
rect 2147 148 2148 152
rect 2142 147 2148 148
rect 2310 152 2316 153
rect 2310 148 2311 152
rect 2315 148 2316 152
rect 2310 147 2316 148
rect 2494 152 2500 153
rect 2494 148 2495 152
rect 2499 148 2500 152
rect 2494 147 2500 148
rect 2702 152 2708 153
rect 2702 148 2703 152
rect 2707 148 2708 152
rect 2702 147 2708 148
rect 2918 152 2924 153
rect 2918 148 2919 152
rect 2923 148 2924 152
rect 2918 147 2924 148
rect 3134 152 3140 153
rect 3134 148 3135 152
rect 3139 148 3140 152
rect 3134 147 3140 148
rect 1630 143 1631 147
rect 1635 143 1636 147
rect 1630 142 1636 143
rect 198 140 204 141
rect 198 136 199 140
rect 203 136 204 140
rect 198 135 204 136
rect 366 140 372 141
rect 366 136 367 140
rect 371 136 372 140
rect 366 135 372 136
rect 534 140 540 141
rect 534 136 535 140
rect 539 136 540 140
rect 534 135 540 136
rect 694 140 700 141
rect 694 136 695 140
rect 699 136 700 140
rect 694 135 700 136
rect 862 140 868 141
rect 862 136 863 140
rect 867 136 868 140
rect 862 135 868 136
rect 1030 140 1036 141
rect 1030 136 1031 140
rect 1035 136 1036 140
rect 1030 135 1036 136
rect 1694 124 1700 125
rect 1694 120 1695 124
rect 1699 120 1700 124
rect 1694 119 1700 120
rect 1814 124 1820 125
rect 1814 120 1815 124
rect 1819 120 1820 124
rect 1814 119 1820 120
rect 1942 124 1948 125
rect 1942 120 1943 124
rect 1947 120 1948 124
rect 1942 119 1948 120
rect 2070 124 2076 125
rect 2070 120 2071 124
rect 2075 120 2076 124
rect 2070 119 2076 120
rect 2198 124 2204 125
rect 2198 120 2199 124
rect 2203 120 2204 124
rect 2198 119 2204 120
rect 2350 124 2356 125
rect 2350 120 2351 124
rect 2355 120 2356 124
rect 2350 119 2356 120
rect 2518 124 2524 125
rect 2518 120 2519 124
rect 2523 120 2524 124
rect 2518 119 2524 120
rect 2710 124 2716 125
rect 2710 120 2711 124
rect 2715 120 2716 124
rect 2710 119 2716 120
rect 2910 124 2916 125
rect 2910 120 2911 124
rect 2915 120 2916 124
rect 2910 119 2916 120
rect 3110 124 3116 125
rect 3110 120 3111 124
rect 3115 120 3116 124
rect 3110 119 3116 120
rect 1670 117 1676 118
rect 134 116 140 117
rect 134 112 135 116
rect 139 112 140 116
rect 134 111 140 112
rect 190 116 196 117
rect 190 112 191 116
rect 195 112 196 116
rect 190 111 196 112
rect 286 116 292 117
rect 286 112 287 116
rect 291 112 292 116
rect 286 111 292 112
rect 382 116 388 117
rect 382 112 383 116
rect 387 112 388 116
rect 382 111 388 112
rect 478 116 484 117
rect 478 112 479 116
rect 483 112 484 116
rect 478 111 484 112
rect 582 116 588 117
rect 582 112 583 116
rect 587 112 588 116
rect 582 111 588 112
rect 694 116 700 117
rect 694 112 695 116
rect 699 112 700 116
rect 694 111 700 112
rect 814 116 820 117
rect 814 112 815 116
rect 819 112 820 116
rect 814 111 820 112
rect 942 116 948 117
rect 942 112 943 116
rect 947 112 948 116
rect 942 111 948 112
rect 1078 116 1084 117
rect 1078 112 1079 116
rect 1083 112 1084 116
rect 1078 111 1084 112
rect 1214 116 1220 117
rect 1214 112 1215 116
rect 1219 112 1220 116
rect 1214 111 1220 112
rect 1350 116 1356 117
rect 1350 112 1351 116
rect 1355 112 1356 116
rect 1350 111 1356 112
rect 1486 116 1492 117
rect 1486 112 1487 116
rect 1491 112 1492 116
rect 1486 111 1492 112
rect 1598 116 1604 117
rect 1598 112 1599 116
rect 1603 112 1604 116
rect 1670 113 1671 117
rect 1675 113 1676 117
rect 1670 112 1676 113
rect 3190 117 3196 118
rect 3190 113 3191 117
rect 3195 113 3196 117
rect 3190 112 3196 113
rect 1598 111 1604 112
rect 110 109 116 110
rect 110 105 111 109
rect 115 105 116 109
rect 110 104 116 105
rect 1630 109 1636 110
rect 1630 105 1631 109
rect 1635 105 1636 109
rect 1630 104 1636 105
rect 1670 99 1676 100
rect 546 95 552 96
rect 546 94 547 95
rect 148 92 395 94
rect 489 92 547 94
rect 110 91 116 92
rect 110 87 111 91
rect 115 87 116 91
rect 143 91 152 92
rect 110 86 116 87
rect 134 87 140 88
rect 134 83 135 87
rect 139 83 140 87
rect 143 87 144 91
rect 151 87 152 91
rect 199 91 205 92
rect 143 86 152 87
rect 190 87 196 88
rect 134 82 140 83
rect 190 83 191 87
rect 195 83 196 87
rect 199 87 200 91
rect 204 87 205 91
rect 295 91 301 92
rect 199 86 205 87
rect 286 87 292 88
rect 190 82 196 83
rect 286 83 287 87
rect 291 83 292 87
rect 295 87 296 91
rect 300 87 301 91
rect 391 91 397 92
rect 295 86 301 87
rect 382 87 388 88
rect 286 82 292 83
rect 382 83 383 87
rect 387 83 388 87
rect 391 87 392 91
rect 396 87 397 91
rect 487 91 493 92
rect 391 86 397 87
rect 478 87 484 88
rect 382 82 388 83
rect 478 83 479 87
rect 483 83 484 87
rect 487 87 488 91
rect 492 87 493 91
rect 546 91 547 92
rect 551 94 552 95
rect 1022 95 1028 96
rect 1022 94 1023 95
rect 551 92 595 94
rect 808 92 1023 94
rect 551 91 552 92
rect 546 90 552 91
rect 591 91 597 92
rect 487 86 493 87
rect 582 87 588 88
rect 478 82 484 83
rect 582 83 583 87
rect 587 83 588 87
rect 591 87 592 91
rect 596 87 597 91
rect 702 91 709 92
rect 591 86 597 87
rect 694 87 700 88
rect 582 82 588 83
rect 694 83 695 87
rect 699 83 700 87
rect 702 87 703 91
rect 708 90 709 91
rect 808 90 810 92
rect 708 88 810 90
rect 823 91 829 92
rect 708 87 709 88
rect 702 86 709 87
rect 814 87 820 88
rect 694 82 700 83
rect 814 83 815 87
rect 819 83 820 87
rect 823 87 824 91
rect 828 87 829 91
rect 951 91 957 92
rect 823 86 829 87
rect 942 87 948 88
rect 814 82 820 83
rect 942 83 943 87
rect 947 83 948 87
rect 951 87 952 91
rect 956 87 957 91
rect 1022 91 1023 92
rect 1027 94 1028 95
rect 1670 95 1671 99
rect 1675 95 1676 99
rect 2358 99 2365 100
rect 1670 94 1676 95
rect 1694 95 1700 96
rect 1027 92 1611 94
rect 1027 91 1028 92
rect 1022 90 1028 91
rect 1087 91 1093 92
rect 951 86 957 87
rect 1078 87 1084 88
rect 942 82 948 83
rect 1078 83 1079 87
rect 1083 83 1084 87
rect 1087 87 1088 91
rect 1092 87 1093 91
rect 1223 91 1229 92
rect 1087 86 1093 87
rect 1214 87 1220 88
rect 1078 82 1084 83
rect 1214 83 1215 87
rect 1219 83 1220 87
rect 1223 87 1224 91
rect 1228 87 1229 91
rect 1359 91 1365 92
rect 1223 86 1229 87
rect 1350 87 1356 88
rect 1214 82 1220 83
rect 1350 83 1351 87
rect 1355 83 1356 87
rect 1359 87 1360 91
rect 1364 87 1365 91
rect 1495 91 1501 92
rect 1359 86 1365 87
rect 1486 87 1492 88
rect 1350 82 1356 83
rect 1486 83 1487 87
rect 1491 83 1492 87
rect 1495 87 1496 91
rect 1500 87 1501 91
rect 1607 91 1613 92
rect 1495 86 1501 87
rect 1598 87 1604 88
rect 1486 82 1492 83
rect 1598 83 1599 87
rect 1603 83 1604 87
rect 1607 87 1608 91
rect 1612 87 1613 91
rect 1607 86 1613 87
rect 1630 91 1636 92
rect 1630 87 1631 91
rect 1635 87 1636 91
rect 1694 91 1695 95
rect 1699 91 1700 95
rect 1694 90 1700 91
rect 1703 95 1709 96
rect 1703 91 1704 95
rect 1708 91 1709 95
rect 1703 90 1709 91
rect 1814 95 1820 96
rect 1814 91 1815 95
rect 1819 91 1820 95
rect 1814 90 1820 91
rect 1823 95 1829 96
rect 1823 91 1824 95
rect 1828 91 1829 95
rect 1823 90 1829 91
rect 1942 95 1948 96
rect 1942 91 1943 95
rect 1947 91 1948 95
rect 1942 90 1948 91
rect 1951 95 1957 96
rect 1951 91 1952 95
rect 1956 91 1957 95
rect 1951 90 1957 91
rect 2070 95 2076 96
rect 2070 91 2071 95
rect 2075 91 2076 95
rect 2070 90 2076 91
rect 2079 95 2085 96
rect 2079 91 2080 95
rect 2084 91 2085 95
rect 2079 90 2085 91
rect 2198 95 2204 96
rect 2198 91 2199 95
rect 2203 91 2204 95
rect 2198 90 2204 91
rect 2207 95 2213 96
rect 2207 91 2208 95
rect 2212 91 2213 95
rect 2207 90 2213 91
rect 2350 95 2356 96
rect 2350 91 2351 95
rect 2355 91 2356 95
rect 2358 95 2359 99
rect 2364 95 2365 99
rect 2526 99 2533 100
rect 2358 94 2365 95
rect 2518 95 2524 96
rect 2350 90 2356 91
rect 2518 91 2519 95
rect 2523 91 2524 95
rect 2526 95 2527 99
rect 2532 95 2533 99
rect 2718 99 2725 100
rect 2526 94 2533 95
rect 2710 95 2716 96
rect 2518 90 2524 91
rect 2710 91 2711 95
rect 2715 91 2716 95
rect 2718 95 2719 99
rect 2724 95 2725 99
rect 2919 99 2925 100
rect 2718 94 2725 95
rect 2910 95 2916 96
rect 2710 90 2716 91
rect 2910 91 2911 95
rect 2915 91 2916 95
rect 2919 95 2920 99
rect 2924 95 2925 99
rect 3119 99 3125 100
rect 2919 94 2925 95
rect 3110 95 3116 96
rect 2910 90 2916 91
rect 3110 91 3111 95
rect 3115 91 3116 95
rect 3119 95 3120 99
rect 3124 98 3125 99
rect 3142 99 3148 100
rect 3142 98 3143 99
rect 3124 96 3143 98
rect 3124 95 3125 96
rect 3119 94 3125 95
rect 3142 95 3143 96
rect 3147 95 3148 99
rect 3142 94 3148 95
rect 3190 99 3196 100
rect 3190 95 3191 99
rect 3195 95 3196 99
rect 3190 94 3196 95
rect 3110 90 3116 91
rect 1630 86 1636 87
rect 1704 86 1706 90
rect 1750 87 1756 88
rect 1750 86 1751 87
rect 1598 82 1604 83
rect 1609 82 1611 86
rect 1704 84 1751 86
rect 1704 82 1706 84
rect 1750 83 1751 84
rect 1755 86 1756 87
rect 1824 86 1826 90
rect 1952 86 1954 90
rect 2080 86 2082 90
rect 2209 86 2211 90
rect 1755 84 2211 86
rect 1755 83 1756 84
rect 1750 82 1756 83
rect 1609 80 1706 82
<< m3c >>
rect 3055 3300 3059 3304
rect 1671 3293 1675 3297
rect 3191 3293 3195 3297
rect 1671 3275 1675 3279
rect 3055 3271 3059 3275
rect 3119 3271 3123 3275
rect 3191 3275 3195 3279
rect 1671 3257 1675 3261
rect 2151 3261 2155 3265
rect 2287 3261 2291 3265
rect 2423 3261 2427 3265
rect 2567 3261 2571 3265
rect 2711 3261 2715 3265
rect 2855 3261 2859 3265
rect 2999 3261 3003 3265
rect 2183 3255 2187 3259
rect 2555 3255 2559 3259
rect 2735 3255 2739 3259
rect 3191 3257 3195 3261
rect 1671 3239 1675 3243
rect 3191 3239 3195 3243
rect 2151 3232 2155 3236
rect 2287 3232 2291 3236
rect 2423 3232 2427 3236
rect 2567 3232 2571 3236
rect 2711 3232 2715 3236
rect 2855 3232 2859 3236
rect 2999 3232 3003 3236
rect 1999 3220 2003 3224
rect 2175 3220 2179 3224
rect 2359 3220 2363 3224
rect 2543 3220 2547 3224
rect 2727 3220 2731 3224
rect 2919 3220 2923 3224
rect 3111 3220 3115 3224
rect 1671 3213 1675 3217
rect 3191 3213 3195 3217
rect 1671 3195 1675 3199
rect 1999 3191 2003 3195
rect 2047 3191 2051 3195
rect 2175 3191 2179 3195
rect 2183 3191 2184 3195
rect 2184 3191 2187 3195
rect 2235 3191 2239 3195
rect 2359 3191 2363 3195
rect 1671 3177 1675 3181
rect 1847 3181 1851 3185
rect 2039 3181 2043 3185
rect 1855 3175 1856 3179
rect 1856 3175 1859 3179
rect 2047 3179 2048 3183
rect 2048 3179 2051 3183
rect 2183 3179 2187 3183
rect 2247 3181 2251 3185
rect 2235 3175 2239 3179
rect 2543 3191 2547 3195
rect 2555 3195 2556 3199
rect 2556 3195 2559 3199
rect 2727 3191 2731 3195
rect 2735 3195 2736 3199
rect 2736 3195 2739 3199
rect 2919 3191 2923 3195
rect 2927 3191 2928 3195
rect 2928 3191 2931 3195
rect 3111 3191 3115 3195
rect 3119 3191 3120 3195
rect 3120 3191 3123 3195
rect 3191 3195 3195 3199
rect 2463 3181 2467 3185
rect 2695 3181 2699 3185
rect 2555 3175 2559 3179
rect 2703 3179 2704 3183
rect 2704 3179 2707 3183
rect 2735 3179 2739 3183
rect 2935 3181 2939 3185
rect 3159 3181 3163 3185
rect 2927 3175 2931 3179
rect 3191 3177 3195 3181
rect 1671 3159 1675 3163
rect 3191 3159 3195 3163
rect 1847 3152 1851 3156
rect 2039 3152 2043 3156
rect 2247 3152 2251 3156
rect 2463 3152 2467 3156
rect 2695 3152 2699 3156
rect 2935 3152 2939 3156
rect 3159 3152 3163 3156
rect 1695 3140 1699 3144
rect 1863 3140 1867 3144
rect 2023 3140 2027 3144
rect 2183 3140 2187 3144
rect 2343 3140 2347 3144
rect 2511 3140 2515 3144
rect 1671 3133 1675 3137
rect 3191 3133 3195 3137
rect 111 3117 115 3121
rect 807 3121 811 3125
rect 1079 3121 1083 3125
rect 1351 3121 1355 3125
rect 1599 3121 1603 3125
rect 839 3115 843 3119
rect 1087 3115 1088 3119
rect 1088 3115 1091 3119
rect 1343 3115 1347 3119
rect 1631 3117 1635 3121
rect 1855 3123 1859 3127
rect 1671 3115 1675 3119
rect 1695 3111 1699 3115
rect 1704 3115 1708 3119
rect 1863 3111 1867 3115
rect 2023 3111 2027 3115
rect 2047 3115 2051 3119
rect 2183 3111 2187 3115
rect 2235 3111 2239 3115
rect 2343 3111 2347 3115
rect 111 3099 115 3103
rect 1631 3099 1635 3103
rect 1879 3103 1883 3107
rect 1671 3097 1675 3101
rect 1959 3101 1963 3105
rect 2183 3101 2187 3105
rect 807 3092 811 3096
rect 1079 3092 1083 3096
rect 1351 3092 1355 3096
rect 1599 3092 1603 3096
rect 1879 3095 1883 3099
rect 2047 3095 2051 3099
rect 2415 3101 2419 3105
rect 2511 3111 2515 3115
rect 2555 3115 2559 3119
rect 3191 3115 3195 3119
rect 2655 3101 2659 3105
rect 2663 3099 2664 3103
rect 2664 3099 2667 3103
rect 2703 3099 2707 3103
rect 2903 3101 2907 3105
rect 3159 3101 3163 3105
rect 2911 3095 2912 3099
rect 2912 3095 2915 3099
rect 2927 3095 2931 3099
rect 3167 3095 3168 3099
rect 3168 3095 3171 3099
rect 3191 3097 3195 3101
rect 703 3076 707 3080
rect 831 3076 835 3080
rect 959 3076 963 3080
rect 1079 3076 1083 3080
rect 1199 3076 1203 3080
rect 1311 3076 1315 3080
rect 1423 3076 1427 3080
rect 1543 3076 1547 3080
rect 1671 3079 1675 3083
rect 3191 3079 3195 3083
rect 111 3069 115 3073
rect 1631 3069 1635 3073
rect 1959 3072 1963 3076
rect 2183 3072 2187 3076
rect 2415 3072 2419 3076
rect 2655 3072 2659 3076
rect 2903 3072 2907 3076
rect 3159 3072 3163 3076
rect 1871 3060 1875 3064
rect 2111 3060 2115 3064
rect 2367 3060 2371 3064
rect 2631 3060 2635 3064
rect 2903 3060 2907 3064
rect 3159 3060 3163 3064
rect 111 3051 115 3055
rect 703 3047 707 3051
rect 711 3047 712 3051
rect 712 3047 715 3051
rect 831 3047 835 3051
rect 839 3051 840 3055
rect 840 3051 843 3055
rect 959 3047 963 3051
rect 967 3047 968 3051
rect 968 3047 971 3051
rect 1079 3047 1083 3051
rect 1087 3051 1088 3055
rect 1088 3051 1091 3055
rect 1199 3047 1203 3051
rect 1207 3047 1208 3051
rect 1208 3047 1211 3051
rect 1311 3047 1315 3051
rect 1319 3047 1320 3051
rect 1320 3047 1323 3051
rect 1423 3047 1427 3051
rect 1447 3051 1451 3055
rect 1543 3047 1547 3051
rect 1631 3051 1635 3055
rect 1671 3053 1675 3057
rect 3191 3053 3195 3057
rect 1671 3035 1675 3039
rect 111 3025 115 3029
rect 623 3029 627 3033
rect 631 3027 632 3031
rect 632 3027 635 3031
rect 711 3027 715 3031
rect 783 3029 787 3033
rect 791 3027 792 3031
rect 792 3027 795 3031
rect 839 3027 843 3031
rect 927 3029 931 3033
rect 935 3027 936 3031
rect 936 3027 939 3031
rect 967 3027 971 3031
rect 1063 3029 1067 3033
rect 1087 3027 1091 3031
rect 1191 3029 1195 3033
rect 1199 3025 1200 3027
rect 1200 3025 1203 3027
rect 1311 3029 1315 3033
rect 1439 3029 1443 3033
rect 1199 3023 1203 3025
rect 1319 3023 1320 3027
rect 1320 3023 1323 3027
rect 1343 3023 1347 3027
rect 1447 3027 1448 3031
rect 1448 3027 1451 3031
rect 1871 3031 1875 3035
rect 1879 3035 1880 3039
rect 1880 3035 1883 3039
rect 2111 3031 2115 3035
rect 2135 3031 2139 3035
rect 2367 3031 2371 3035
rect 2631 3031 2635 3035
rect 2663 3035 2667 3039
rect 1631 3025 1635 3029
rect 1671 3017 1675 3021
rect 1791 3021 1795 3025
rect 1959 3021 1963 3025
rect 2127 3021 2131 3025
rect 2287 3021 2291 3025
rect 1715 3015 1719 3019
rect 1879 3015 1883 3019
rect 1911 3015 1915 3019
rect 2135 3015 2136 3019
rect 2136 3015 2139 3019
rect 2295 3019 2296 3023
rect 2296 3019 2299 3023
rect 2455 3021 2459 3025
rect 2623 3021 2627 3025
rect 2379 3015 2383 3019
rect 2527 3015 2531 3019
rect 2903 3031 2907 3035
rect 2911 3031 2912 3035
rect 2912 3031 2915 3035
rect 3159 3031 3163 3035
rect 3167 3035 3168 3039
rect 3168 3035 3171 3039
rect 3191 3035 3195 3039
rect 2631 3015 2635 3019
rect 3191 3017 3195 3021
rect 111 3007 115 3011
rect 1631 3007 1635 3011
rect 623 3000 627 3004
rect 783 3000 787 3004
rect 927 3000 931 3004
rect 1063 3000 1067 3004
rect 1191 3000 1195 3004
rect 1311 3000 1315 3004
rect 1439 3000 1443 3004
rect 1671 2999 1675 3003
rect 3191 2999 3195 3003
rect 1791 2992 1795 2996
rect 1959 2992 1963 2996
rect 2127 2992 2131 2996
rect 2287 2992 2291 2996
rect 2455 2992 2459 2996
rect 2623 2992 2627 2996
rect 519 2984 523 2988
rect 647 2984 651 2988
rect 783 2984 787 2988
rect 919 2984 923 2988
rect 1055 2984 1059 2988
rect 1191 2984 1195 2988
rect 1335 2984 1339 2988
rect 111 2977 115 2981
rect 1631 2977 1635 2981
rect 1703 2980 1707 2984
rect 1903 2980 1907 2984
rect 2127 2980 2131 2984
rect 2367 2980 2371 2984
rect 2623 2980 2627 2984
rect 2887 2980 2891 2984
rect 3159 2980 3163 2984
rect 1671 2973 1675 2977
rect 3191 2973 3195 2977
rect 111 2959 115 2963
rect 519 2955 523 2959
rect 647 2955 651 2959
rect 783 2955 787 2959
rect 791 2959 792 2963
rect 792 2959 795 2963
rect 803 2959 807 2963
rect 919 2955 923 2959
rect 928 2959 932 2963
rect 1055 2955 1059 2959
rect 1087 2959 1091 2963
rect 1103 2959 1107 2963
rect 1199 2963 1203 2967
rect 1191 2955 1195 2959
rect 1335 2955 1339 2959
rect 1343 2955 1344 2959
rect 1344 2955 1347 2959
rect 1631 2959 1635 2963
rect 1671 2955 1675 2959
rect 479 2947 483 2951
rect 111 2933 115 2937
rect 439 2937 443 2941
rect 599 2937 603 2941
rect 631 2947 635 2951
rect 1703 2951 1707 2955
rect 1715 2955 1716 2959
rect 1716 2955 1719 2959
rect 1903 2951 1907 2955
rect 1911 2955 1912 2959
rect 1912 2955 1915 2959
rect 2127 2951 2131 2955
rect 2135 2951 2136 2955
rect 2136 2951 2139 2955
rect 2231 2951 2235 2955
rect 2367 2951 2371 2955
rect 2379 2955 2380 2959
rect 2380 2955 2383 2959
rect 2623 2951 2627 2955
rect 2631 2955 2632 2959
rect 2632 2955 2635 2959
rect 2887 2951 2891 2955
rect 2911 2951 2915 2955
rect 3159 2951 3163 2955
rect 3167 2955 3168 2959
rect 3168 2955 3171 2959
rect 3191 2955 3195 2959
rect 479 2931 483 2935
rect 759 2937 763 2941
rect 927 2937 931 2941
rect 1095 2937 1099 2941
rect 1263 2937 1267 2941
rect 1439 2937 1443 2941
rect 803 2931 807 2935
rect 935 2931 936 2935
rect 936 2931 939 2935
rect 1103 2931 1104 2935
rect 1104 2931 1107 2935
rect 1343 2931 1347 2935
rect 1447 2935 1448 2939
rect 1448 2935 1451 2939
rect 1599 2937 1603 2941
rect 1631 2933 1635 2937
rect 1671 2937 1675 2941
rect 1695 2941 1699 2945
rect 1715 2939 1719 2943
rect 1935 2941 1939 2945
rect 2223 2941 2227 2945
rect 1611 2927 1615 2931
rect 1911 2935 1915 2939
rect 2231 2935 2232 2939
rect 2232 2935 2235 2939
rect 2295 2939 2299 2943
rect 2519 2941 2523 2945
rect 2527 2939 2528 2943
rect 2528 2939 2531 2943
rect 2823 2941 2827 2945
rect 3135 2941 3139 2945
rect 2835 2935 2836 2939
rect 2836 2935 2839 2939
rect 3143 2939 3144 2943
rect 3144 2939 3147 2943
rect 3167 2939 3171 2943
rect 3191 2937 3195 2941
rect 111 2915 115 2919
rect 1631 2915 1635 2919
rect 1671 2919 1675 2923
rect 3191 2919 3195 2923
rect 439 2908 443 2912
rect 599 2908 603 2912
rect 759 2908 763 2912
rect 927 2908 931 2912
rect 1095 2908 1099 2912
rect 1263 2908 1267 2912
rect 1439 2908 1443 2912
rect 1599 2908 1603 2912
rect 1695 2912 1699 2916
rect 1935 2912 1939 2916
rect 2223 2912 2227 2916
rect 2519 2912 2523 2916
rect 2823 2912 2827 2916
rect 3135 2912 3139 2916
rect 335 2896 339 2900
rect 471 2896 475 2900
rect 623 2896 627 2900
rect 791 2896 795 2900
rect 975 2896 979 2900
rect 1175 2896 1179 2900
rect 1383 2896 1387 2900
rect 1591 2896 1595 2900
rect 2295 2900 2299 2904
rect 2551 2900 2555 2904
rect 2815 2900 2819 2904
rect 3079 2900 3083 2904
rect 111 2889 115 2893
rect 1631 2889 1635 2893
rect 1671 2893 1675 2897
rect 3191 2893 3195 2897
rect 111 2871 115 2875
rect 335 2867 339 2871
rect 471 2867 475 2871
rect 479 2867 480 2871
rect 480 2867 483 2871
rect 623 2867 627 2871
rect 703 2867 707 2871
rect 791 2867 795 2871
rect 803 2867 804 2871
rect 804 2867 807 2871
rect 975 2867 979 2871
rect 983 2867 984 2871
rect 984 2867 987 2871
rect 1175 2867 1179 2871
rect 1383 2867 1387 2871
rect 1591 2867 1595 2871
rect 1611 2871 1615 2875
rect 1631 2871 1635 2875
rect 1671 2875 1675 2879
rect 2295 2871 2299 2875
rect 2303 2875 2304 2879
rect 2304 2875 2307 2879
rect 2527 2879 2531 2883
rect 2543 2879 2547 2883
rect 2551 2871 2555 2875
rect 2815 2871 2819 2875
rect 2835 2871 2839 2875
rect 3079 2871 3083 2875
rect 3191 2875 3195 2879
rect 287 2859 291 2863
rect 1095 2859 1099 2863
rect 1103 2859 1107 2863
rect 1343 2859 1347 2863
rect 1671 2857 1675 2861
rect 2207 2861 2211 2865
rect 2303 2859 2307 2863
rect 2375 2861 2379 2865
rect 2535 2861 2539 2865
rect 2383 2855 2384 2859
rect 2384 2855 2387 2859
rect 2543 2859 2544 2863
rect 2544 2859 2547 2863
rect 2679 2861 2683 2865
rect 2823 2861 2827 2865
rect 2967 2861 2971 2865
rect 3111 2861 3115 2865
rect 2687 2855 2688 2859
rect 2688 2855 2691 2859
rect 2835 2855 2836 2859
rect 2836 2855 2839 2859
rect 2975 2855 2976 2859
rect 2976 2855 2979 2859
rect 3143 2859 3147 2863
rect 3167 2859 3171 2863
rect 3191 2857 3195 2861
rect 111 2845 115 2849
rect 255 2849 259 2853
rect 415 2849 419 2853
rect 559 2849 563 2853
rect 695 2849 699 2853
rect 823 2849 827 2853
rect 951 2849 955 2853
rect 1087 2849 1091 2853
rect 287 2843 291 2847
rect 423 2843 424 2847
rect 424 2843 427 2847
rect 479 2843 483 2847
rect 703 2843 704 2847
rect 704 2843 707 2847
rect 803 2843 807 2847
rect 871 2843 875 2847
rect 935 2843 939 2847
rect 983 2843 987 2847
rect 1095 2843 1096 2847
rect 1096 2843 1099 2847
rect 1631 2845 1635 2849
rect 1671 2839 1675 2843
rect 3191 2839 3195 2843
rect 2207 2832 2211 2836
rect 111 2827 115 2831
rect 2375 2832 2379 2836
rect 2535 2832 2539 2836
rect 2679 2832 2683 2836
rect 2823 2832 2827 2836
rect 2967 2832 2971 2836
rect 3111 2832 3115 2836
rect 1631 2827 1635 2831
rect 255 2820 259 2824
rect 415 2820 419 2824
rect 559 2820 563 2824
rect 695 2820 699 2824
rect 823 2820 827 2824
rect 951 2820 955 2824
rect 1087 2820 1091 2824
rect 2127 2812 2131 2816
rect 2303 2812 2307 2816
rect 2479 2812 2483 2816
rect 2655 2812 2659 2816
rect 2831 2812 2835 2816
rect 3007 2812 3011 2816
rect 3159 2812 3163 2816
rect 1671 2805 1675 2809
rect 151 2800 155 2804
rect 279 2800 283 2804
rect 399 2800 403 2804
rect 519 2800 523 2804
rect 639 2800 643 2804
rect 751 2800 755 2804
rect 863 2800 867 2804
rect 3191 2805 3195 2809
rect 983 2800 987 2804
rect 111 2793 115 2797
rect 1631 2793 1635 2797
rect 1671 2787 1675 2791
rect 111 2775 115 2779
rect 287 2779 291 2783
rect 151 2771 155 2775
rect 159 2771 160 2775
rect 160 2771 163 2775
rect 279 2771 283 2775
rect 287 2771 288 2775
rect 288 2771 291 2775
rect 399 2771 403 2775
rect 423 2779 427 2783
rect 519 2771 523 2775
rect 631 2779 635 2783
rect 639 2771 643 2775
rect 703 2779 707 2783
rect 2127 2783 2131 2787
rect 2303 2783 2307 2787
rect 2311 2787 2312 2791
rect 2312 2787 2315 2791
rect 2351 2787 2355 2791
rect 2383 2787 2387 2791
rect 2479 2783 2483 2787
rect 2975 2791 2979 2795
rect 2655 2783 2659 2787
rect 2687 2783 2691 2787
rect 751 2771 755 2775
rect 863 2771 867 2775
rect 871 2775 872 2779
rect 872 2775 875 2779
rect 967 2775 971 2779
rect 983 2771 987 2775
rect 1631 2775 1635 2779
rect 1671 2769 1675 2773
rect 2039 2773 2043 2777
rect 2023 2767 2027 2771
rect 2207 2773 2211 2777
rect 2375 2773 2379 2777
rect 2231 2767 2235 2771
rect 2383 2771 2384 2775
rect 2384 2771 2387 2775
rect 2535 2773 2539 2777
rect 2559 2771 2563 2775
rect 2703 2773 2707 2777
rect 2831 2783 2835 2787
rect 2839 2783 2840 2787
rect 2840 2783 2843 2787
rect 3007 2783 3011 2787
rect 3015 2783 3016 2787
rect 3016 2783 3019 2787
rect 3159 2783 3163 2787
rect 3167 2783 3168 2787
rect 3168 2783 3171 2787
rect 3191 2787 3195 2791
rect 2871 2773 2875 2777
rect 2839 2767 2843 2771
rect 3191 2769 3195 2773
rect 111 2745 115 2749
rect 135 2749 139 2753
rect 159 2747 163 2751
rect 263 2749 267 2753
rect 431 2749 435 2753
rect 623 2749 627 2753
rect 287 2743 291 2747
rect 423 2743 427 2747
rect 631 2747 632 2751
rect 632 2747 635 2751
rect 839 2749 843 2753
rect 871 2747 875 2751
rect 1071 2749 1075 2753
rect 1319 2749 1323 2753
rect 1567 2749 1571 2753
rect 1103 2743 1107 2747
rect 1343 2743 1347 2747
rect 1575 2747 1576 2751
rect 1576 2747 1579 2751
rect 1611 2747 1615 2751
rect 1671 2751 1675 2755
rect 3191 2751 3195 2755
rect 1631 2745 1635 2749
rect 2039 2744 2043 2748
rect 2207 2744 2211 2748
rect 2375 2744 2379 2748
rect 2535 2744 2539 2748
rect 2703 2744 2707 2748
rect 2871 2744 2875 2748
rect 111 2727 115 2731
rect 1631 2727 1635 2731
rect 2015 2728 2019 2732
rect 2199 2728 2203 2732
rect 2383 2728 2387 2732
rect 2575 2728 2579 2732
rect 2775 2728 2779 2732
rect 2975 2728 2979 2732
rect 3159 2728 3163 2732
rect 135 2720 139 2724
rect 263 2720 267 2724
rect 431 2720 435 2724
rect 623 2720 627 2724
rect 839 2720 843 2724
rect 1071 2720 1075 2724
rect 1319 2720 1323 2724
rect 1567 2720 1571 2724
rect 1671 2721 1675 2725
rect 3191 2721 3195 2725
rect 1671 2703 1675 2707
rect 2559 2707 2563 2711
rect 703 2696 707 2700
rect 831 2696 835 2700
rect 959 2696 963 2700
rect 1079 2696 1083 2700
rect 1199 2696 1203 2700
rect 1311 2696 1315 2700
rect 1423 2696 1427 2700
rect 1543 2696 1547 2700
rect 2015 2699 2019 2703
rect 2023 2699 2024 2703
rect 2024 2699 2027 2703
rect 2199 2699 2203 2703
rect 2207 2699 2208 2703
rect 2208 2699 2211 2703
rect 2383 2699 2387 2703
rect 2391 2699 2392 2703
rect 2392 2699 2395 2703
rect 2447 2699 2451 2703
rect 2575 2699 2579 2703
rect 2775 2699 2779 2703
rect 2783 2703 2784 2707
rect 2784 2703 2787 2707
rect 2839 2703 2843 2707
rect 2927 2703 2931 2707
rect 2975 2699 2979 2703
rect 3015 2699 3019 2703
rect 3159 2699 3163 2703
rect 3167 2699 3168 2703
rect 3168 2699 3171 2703
rect 3191 2703 3195 2707
rect 111 2689 115 2693
rect 1631 2689 1635 2693
rect 111 2671 115 2675
rect 631 2675 635 2679
rect 703 2667 707 2671
rect 743 2671 747 2675
rect 831 2667 835 2671
rect 863 2667 867 2671
rect 959 2667 963 2671
rect 967 2671 968 2675
rect 968 2671 971 2675
rect 1079 2667 1083 2671
rect 1103 2667 1107 2671
rect 1199 2667 1203 2671
rect 1207 2667 1208 2671
rect 1208 2667 1211 2671
rect 1311 2667 1315 2671
rect 1343 2675 1347 2679
rect 1423 2667 1427 2671
rect 1447 2675 1451 2679
rect 1671 2677 1675 2681
rect 1999 2681 2003 2685
rect 2175 2681 2179 2685
rect 2359 2681 2363 2685
rect 1543 2667 1547 2671
rect 1575 2671 1579 2675
rect 1631 2671 1635 2675
rect 2007 2675 2008 2679
rect 2008 2675 2011 2679
rect 2023 2675 2027 2679
rect 2207 2675 2211 2679
rect 2351 2675 2355 2679
rect 2391 2679 2395 2683
rect 2551 2681 2555 2685
rect 2559 2679 2560 2683
rect 2560 2679 2563 2683
rect 2759 2681 2763 2685
rect 2783 2679 2787 2683
rect 2967 2681 2971 2685
rect 2927 2675 2931 2679
rect 3159 2681 3163 2685
rect 3167 2675 3168 2679
rect 3168 2675 3171 2679
rect 3191 2677 3195 2681
rect 1671 2659 1675 2663
rect 3191 2659 3195 2663
rect 111 2645 115 2649
rect 607 2649 611 2653
rect 631 2647 635 2651
rect 735 2649 739 2653
rect 743 2647 744 2651
rect 744 2647 747 2651
rect 855 2649 859 2653
rect 975 2649 979 2653
rect 1095 2649 1099 2653
rect 1207 2649 1211 2653
rect 1319 2649 1323 2653
rect 863 2643 864 2647
rect 864 2643 867 2647
rect 967 2643 971 2647
rect 1103 2643 1104 2647
rect 1104 2643 1107 2647
rect 1215 2643 1216 2647
rect 1216 2643 1219 2647
rect 1343 2647 1347 2651
rect 1439 2649 1443 2653
rect 1999 2652 2003 2656
rect 2175 2652 2179 2656
rect 2359 2652 2363 2656
rect 2551 2652 2555 2656
rect 2759 2652 2763 2656
rect 2967 2652 2971 2656
rect 3159 2652 3163 2656
rect 1447 2647 1448 2651
rect 1448 2647 1451 2651
rect 1631 2645 1635 2649
rect 1911 2640 1915 2644
rect 2103 2640 2107 2644
rect 2295 2640 2299 2644
rect 2487 2640 2491 2644
rect 2687 2640 2691 2644
rect 1671 2633 1675 2637
rect 3191 2633 3195 2637
rect 111 2627 115 2631
rect 1631 2627 1635 2631
rect 607 2620 611 2624
rect 735 2620 739 2624
rect 855 2620 859 2624
rect 975 2620 979 2624
rect 1095 2620 1099 2624
rect 1207 2620 1211 2624
rect 1319 2620 1323 2624
rect 1439 2620 1443 2624
rect 1671 2615 1675 2619
rect 1911 2611 1915 2615
rect 1919 2611 1920 2615
rect 1920 2611 1923 2615
rect 2103 2611 2107 2615
rect 2295 2611 2299 2615
rect 2327 2615 2331 2619
rect 2351 2615 2355 2619
rect 2487 2611 2491 2615
rect 503 2596 507 2600
rect 631 2596 635 2600
rect 751 2596 755 2600
rect 871 2596 875 2600
rect 991 2596 995 2600
rect 1103 2596 1107 2600
rect 1215 2596 1219 2600
rect 1335 2596 1339 2600
rect 1671 2597 1675 2601
rect 1823 2601 1827 2605
rect 2015 2601 2019 2605
rect 2215 2601 2219 2605
rect 2439 2601 2443 2605
rect 1831 2595 1832 2599
rect 1832 2595 1835 2599
rect 1919 2595 1923 2599
rect 2007 2595 2011 2599
rect 2063 2595 2067 2599
rect 2207 2595 2211 2599
rect 2223 2595 2224 2599
rect 2224 2595 2227 2599
rect 2447 2599 2448 2603
rect 2448 2599 2451 2603
rect 2671 2601 2675 2605
rect 2687 2611 2691 2615
rect 2783 2615 2787 2619
rect 3191 2615 3195 2619
rect 2919 2601 2923 2605
rect 3159 2601 3163 2605
rect 2927 2595 2928 2599
rect 2928 2595 2931 2599
rect 3143 2595 3147 2599
rect 3167 2595 3168 2599
rect 3168 2595 3171 2599
rect 3191 2597 3195 2601
rect 111 2589 115 2593
rect 1631 2589 1635 2593
rect 111 2571 115 2575
rect 863 2575 867 2579
rect 503 2567 507 2571
rect 511 2567 512 2571
rect 512 2567 515 2571
rect 631 2567 635 2571
rect 639 2567 640 2571
rect 640 2567 643 2571
rect 751 2567 755 2571
rect 783 2567 787 2571
rect 871 2567 875 2571
rect 903 2575 907 2579
rect 1671 2579 1675 2583
rect 3191 2579 3195 2583
rect 991 2567 995 2571
rect 1015 2571 1019 2575
rect 1103 2567 1107 2571
rect 1127 2567 1131 2571
rect 1215 2567 1219 2571
rect 1223 2571 1224 2575
rect 1224 2571 1227 2575
rect 1247 2571 1251 2575
rect 1335 2567 1339 2571
rect 1343 2571 1344 2575
rect 1344 2571 1347 2575
rect 1631 2571 1635 2575
rect 1823 2572 1827 2576
rect 2015 2572 2019 2576
rect 2215 2572 2219 2576
rect 2439 2572 2443 2576
rect 2671 2572 2675 2576
rect 2919 2572 2923 2576
rect 3159 2572 3163 2576
rect 1735 2556 1739 2560
rect 1895 2556 1899 2560
rect 2055 2556 2059 2560
rect 2215 2556 2219 2560
rect 2375 2556 2379 2560
rect 2535 2556 2539 2560
rect 111 2541 115 2545
rect 399 2545 403 2549
rect 527 2545 531 2549
rect 655 2545 659 2549
rect 775 2545 779 2549
rect 443 2539 447 2543
rect 511 2539 515 2543
rect 639 2539 643 2543
rect 783 2543 784 2547
rect 784 2543 787 2547
rect 863 2543 867 2547
rect 895 2545 899 2549
rect 903 2543 904 2547
rect 904 2543 907 2547
rect 1007 2545 1011 2549
rect 1015 2543 1016 2547
rect 1016 2543 1019 2547
rect 1119 2545 1123 2549
rect 1239 2545 1243 2549
rect 1671 2549 1675 2553
rect 3191 2549 3195 2553
rect 1127 2539 1128 2543
rect 1128 2539 1131 2543
rect 1247 2543 1248 2547
rect 1248 2543 1251 2547
rect 1631 2541 1635 2545
rect 1671 2531 1675 2535
rect 111 2523 115 2527
rect 1631 2523 1635 2527
rect 1735 2527 1739 2531
rect 1895 2527 1899 2531
rect 1903 2527 1904 2531
rect 1904 2527 1907 2531
rect 1919 2527 1923 2531
rect 2055 2527 2059 2531
rect 2063 2531 2064 2535
rect 2064 2531 2067 2535
rect 2215 2527 2219 2531
rect 2223 2531 2224 2535
rect 2224 2531 2227 2535
rect 2375 2527 2379 2531
rect 2535 2527 2539 2531
rect 3191 2531 3195 2535
rect 399 2516 403 2520
rect 527 2516 531 2520
rect 655 2516 659 2520
rect 775 2516 779 2520
rect 895 2516 899 2520
rect 1007 2516 1011 2520
rect 1119 2516 1123 2520
rect 1239 2516 1243 2520
rect 1671 2509 1675 2513
rect 1695 2513 1699 2517
rect 1863 2513 1867 2517
rect 2079 2513 2083 2517
rect 2319 2513 2323 2517
rect 1831 2507 1835 2511
rect 1903 2507 1907 2511
rect 2063 2507 2067 2511
rect 2327 2511 2328 2515
rect 2328 2511 2331 2515
rect 2575 2519 2579 2523
rect 2583 2513 2587 2517
rect 2855 2513 2859 2517
rect 3135 2513 3139 2517
rect 2863 2507 2864 2511
rect 2864 2507 2867 2511
rect 2927 2507 2931 2511
rect 2975 2507 2979 2511
rect 3143 2507 3144 2511
rect 3144 2507 3147 2511
rect 3191 2509 3195 2513
rect 303 2492 307 2496
rect 431 2492 435 2496
rect 559 2492 563 2496
rect 703 2492 707 2496
rect 863 2492 867 2496
rect 1039 2492 1043 2496
rect 1223 2492 1227 2496
rect 1423 2492 1427 2496
rect 1599 2492 1603 2496
rect 1671 2491 1675 2495
rect 3191 2491 3195 2495
rect 111 2485 115 2489
rect 1631 2485 1635 2489
rect 1695 2484 1699 2488
rect 1863 2484 1867 2488
rect 2079 2484 2083 2488
rect 2319 2484 2323 2488
rect 2583 2484 2587 2488
rect 2855 2484 2859 2488
rect 3135 2484 3139 2488
rect 111 2467 115 2471
rect 303 2463 307 2467
rect 311 2463 312 2467
rect 312 2463 315 2467
rect 431 2463 435 2467
rect 439 2463 440 2467
rect 440 2463 443 2467
rect 559 2463 563 2467
rect 611 2463 615 2467
rect 703 2463 707 2467
rect 775 2463 779 2467
rect 863 2463 867 2467
rect 903 2467 907 2471
rect 1039 2463 1043 2467
rect 1047 2467 1048 2471
rect 1048 2467 1051 2471
rect 1127 2467 1131 2471
rect 1383 2471 1387 2475
rect 1223 2463 1227 2467
rect 1247 2463 1251 2467
rect 1423 2463 1427 2467
rect 1575 2471 1579 2475
rect 1599 2463 1603 2467
rect 1631 2467 1635 2471
rect 2319 2464 2323 2468
rect 2567 2464 2571 2468
rect 2823 2464 2827 2468
rect 3079 2464 3083 2468
rect 1671 2457 1675 2461
rect 3191 2457 3195 2461
rect 111 2445 115 2449
rect 199 2449 203 2453
rect 327 2449 331 2453
rect 455 2449 459 2453
rect 599 2449 603 2453
rect 767 2449 771 2453
rect 951 2449 955 2453
rect 247 2443 251 2447
rect 311 2443 315 2447
rect 439 2443 443 2447
rect 611 2443 612 2447
rect 612 2443 615 2447
rect 775 2443 776 2447
rect 776 2443 779 2447
rect 1047 2447 1051 2451
rect 1159 2449 1163 2453
rect 1183 2447 1187 2451
rect 1247 2447 1251 2451
rect 1375 2449 1379 2453
rect 1383 2447 1384 2451
rect 1384 2447 1387 2451
rect 1591 2449 1595 2453
rect 1631 2445 1635 2449
rect 1671 2439 1675 2443
rect 2319 2435 2323 2439
rect 2327 2439 2328 2443
rect 2328 2439 2331 2443
rect 2567 2435 2571 2439
rect 2575 2439 2576 2443
rect 2576 2439 2579 2443
rect 2823 2435 2827 2439
rect 2863 2439 2867 2443
rect 111 2427 115 2431
rect 1631 2427 1635 2431
rect 199 2420 203 2424
rect 327 2420 331 2424
rect 455 2420 459 2424
rect 599 2420 603 2424
rect 767 2420 771 2424
rect 951 2420 955 2424
rect 1159 2420 1163 2424
rect 1375 2420 1379 2424
rect 1591 2420 1595 2424
rect 1671 2421 1675 2425
rect 2231 2425 2235 2429
rect 2239 2423 2240 2427
rect 2240 2423 2243 2427
rect 2327 2423 2331 2427
rect 2343 2423 2347 2427
rect 2391 2425 2395 2429
rect 2543 2425 2547 2429
rect 2575 2423 2579 2427
rect 2687 2425 2691 2429
rect 2823 2425 2827 2429
rect 3079 2435 3083 2439
rect 3191 2439 3195 2443
rect 2667 2419 2671 2423
rect 2967 2425 2971 2429
rect 3111 2425 3115 2429
rect 2975 2419 2976 2423
rect 2976 2419 2979 2423
rect 3015 2419 3019 2423
rect 3143 2419 3147 2423
rect 3167 2419 3171 2423
rect 3191 2421 3195 2425
rect 1671 2403 1675 2407
rect 3191 2403 3195 2407
rect 135 2392 139 2396
rect 239 2392 243 2396
rect 359 2392 363 2396
rect 479 2392 483 2396
rect 591 2392 595 2396
rect 703 2392 707 2396
rect 815 2392 819 2396
rect 935 2392 939 2396
rect 2231 2396 2235 2400
rect 2391 2396 2395 2400
rect 2543 2396 2547 2400
rect 2687 2396 2691 2400
rect 2823 2396 2827 2400
rect 2967 2396 2971 2400
rect 3111 2396 3115 2400
rect 111 2385 115 2389
rect 1631 2385 1635 2389
rect 611 2375 615 2379
rect 2143 2376 2147 2380
rect 2311 2376 2315 2380
rect 2479 2376 2483 2380
rect 2655 2376 2659 2380
rect 2831 2376 2835 2380
rect 3007 2376 3011 2380
rect 3159 2376 3163 2380
rect 111 2367 115 2371
rect 135 2363 139 2367
rect 143 2363 144 2367
rect 144 2363 147 2367
rect 239 2363 243 2367
rect 247 2363 248 2367
rect 248 2363 251 2367
rect 359 2363 363 2367
rect 367 2363 368 2367
rect 368 2363 371 2367
rect 479 2363 483 2367
rect 575 2363 579 2367
rect 591 2363 595 2367
rect 703 2363 707 2367
rect 775 2363 779 2367
rect 815 2363 819 2367
rect 935 2363 939 2367
rect 943 2363 944 2367
rect 944 2363 947 2367
rect 983 2363 987 2367
rect 1631 2367 1635 2371
rect 1671 2369 1675 2373
rect 3191 2369 3195 2373
rect 791 2355 795 2359
rect 1671 2351 1675 2355
rect 111 2341 115 2345
rect 135 2345 139 2349
rect 343 2345 347 2349
rect 567 2345 571 2349
rect 775 2345 779 2349
rect 975 2345 979 2349
rect 143 2339 144 2343
rect 144 2339 147 2343
rect 183 2339 187 2343
rect 247 2339 251 2343
rect 367 2339 371 2343
rect 575 2339 576 2343
rect 576 2339 579 2343
rect 783 2339 784 2343
rect 784 2339 787 2343
rect 983 2343 984 2347
rect 984 2343 987 2347
rect 1175 2345 1179 2349
rect 1367 2345 1371 2349
rect 1167 2339 1171 2343
rect 1183 2339 1184 2343
rect 1184 2339 1187 2343
rect 1375 2343 1376 2347
rect 1376 2343 1379 2347
rect 1567 2345 1571 2349
rect 1575 2343 1576 2347
rect 1576 2343 1579 2347
rect 2143 2347 2147 2351
rect 2175 2347 2179 2351
rect 2239 2351 2243 2355
rect 2311 2347 2315 2351
rect 2343 2351 2347 2355
rect 2479 2347 2483 2351
rect 2655 2347 2659 2351
rect 2667 2351 2668 2355
rect 2668 2351 2671 2355
rect 2831 2347 2835 2351
rect 1631 2341 1635 2345
rect 1671 2333 1675 2337
rect 2183 2337 2187 2341
rect 2335 2337 2339 2341
rect 2175 2331 2179 2335
rect 2343 2335 2344 2339
rect 2344 2335 2347 2339
rect 2479 2337 2483 2341
rect 2623 2337 2627 2341
rect 2487 2331 2488 2335
rect 2488 2331 2491 2335
rect 2631 2335 2632 2339
rect 2632 2335 2635 2339
rect 2667 2335 2671 2339
rect 2767 2337 2771 2341
rect 2799 2335 2803 2339
rect 2919 2337 2923 2341
rect 3007 2347 3011 2351
rect 3015 2351 3016 2355
rect 3016 2351 3019 2355
rect 3167 2355 3171 2359
rect 3159 2347 3163 2351
rect 3167 2347 3168 2351
rect 3168 2347 3171 2351
rect 3191 2351 3195 2355
rect 3015 2335 3019 2339
rect 3191 2333 3195 2337
rect 111 2323 115 2327
rect 1631 2323 1635 2327
rect 135 2316 139 2320
rect 343 2316 347 2320
rect 567 2316 571 2320
rect 775 2316 779 2320
rect 975 2316 979 2320
rect 1175 2316 1179 2320
rect 1367 2316 1371 2320
rect 1567 2316 1571 2320
rect 1671 2315 1675 2319
rect 3191 2315 3195 2319
rect 2183 2308 2187 2312
rect 2335 2308 2339 2312
rect 2479 2308 2483 2312
rect 2623 2308 2627 2312
rect 2767 2308 2771 2312
rect 2919 2308 2923 2312
rect 655 2292 659 2296
rect 783 2292 787 2296
rect 903 2292 907 2296
rect 1023 2292 1027 2296
rect 1143 2292 1147 2296
rect 1255 2292 1259 2296
rect 1367 2292 1371 2296
rect 1487 2292 1491 2296
rect 2095 2292 2099 2296
rect 2263 2292 2267 2296
rect 2431 2292 2435 2296
rect 2607 2292 2611 2296
rect 2791 2292 2795 2296
rect 2983 2292 2987 2296
rect 3159 2292 3163 2296
rect 111 2285 115 2289
rect 1631 2285 1635 2289
rect 1671 2285 1675 2289
rect 3191 2285 3195 2289
rect 111 2267 115 2271
rect 655 2263 659 2267
rect 663 2263 664 2267
rect 664 2263 667 2267
rect 783 2263 787 2267
rect 791 2263 792 2267
rect 792 2263 795 2267
rect 815 2263 819 2267
rect 903 2263 907 2267
rect 943 2267 947 2271
rect 951 2267 955 2271
rect 1023 2263 1027 2267
rect 1055 2267 1059 2271
rect 1143 2263 1147 2267
rect 1167 2267 1171 2271
rect 1255 2263 1259 2267
rect 1279 2267 1283 2271
rect 1399 2271 1403 2275
rect 1367 2263 1371 2267
rect 1375 2263 1376 2267
rect 1376 2263 1379 2267
rect 1487 2263 1491 2267
rect 1631 2267 1635 2271
rect 1671 2267 1675 2271
rect 2023 2271 2027 2275
rect 2095 2263 2099 2267
rect 2263 2263 2267 2267
rect 2303 2263 2307 2267
rect 2431 2263 2435 2267
rect 2487 2263 2491 2267
rect 2607 2263 2611 2267
rect 2631 2263 2635 2267
rect 2791 2263 2795 2267
rect 2799 2267 2800 2271
rect 2800 2267 2803 2271
rect 2983 2263 2987 2267
rect 2991 2267 2992 2271
rect 2992 2267 2995 2271
rect 3015 2267 3019 2271
rect 3159 2263 3163 2267
rect 3167 2263 3168 2267
rect 3168 2263 3171 2267
rect 3191 2267 3195 2271
rect 1671 2249 1675 2253
rect 2015 2253 2019 2257
rect 2167 2253 2171 2257
rect 2319 2253 2323 2257
rect 2463 2253 2467 2257
rect 111 2237 115 2241
rect 551 2241 555 2245
rect 679 2241 683 2245
rect 807 2241 811 2245
rect 575 2235 579 2239
rect 607 2235 611 2239
rect 663 2235 667 2239
rect 815 2239 816 2243
rect 816 2239 819 2243
rect 927 2241 931 2245
rect 1047 2241 1051 2245
rect 1055 2245 1059 2247
rect 1055 2243 1056 2245
rect 1056 2243 1059 2245
rect 1159 2241 1163 2245
rect 1167 2245 1171 2247
rect 2023 2247 2024 2251
rect 2024 2247 2027 2251
rect 2175 2247 2176 2251
rect 2176 2247 2179 2251
rect 2303 2247 2307 2251
rect 2487 2251 2491 2255
rect 2607 2253 2611 2257
rect 2615 2251 2616 2255
rect 2616 2251 2619 2255
rect 2759 2253 2763 2257
rect 2767 2251 2768 2255
rect 2768 2251 2771 2255
rect 2799 2251 2803 2255
rect 3191 2249 3195 2253
rect 1167 2243 1168 2245
rect 1168 2243 1171 2245
rect 1271 2241 1275 2245
rect 951 2235 955 2239
rect 1279 2239 1280 2243
rect 1280 2239 1283 2243
rect 1391 2241 1395 2245
rect 1399 2239 1400 2243
rect 1400 2239 1403 2243
rect 1631 2237 1635 2241
rect 1671 2231 1675 2235
rect 3191 2231 3195 2235
rect 2015 2224 2019 2228
rect 111 2219 115 2223
rect 2167 2224 2171 2228
rect 2319 2224 2323 2228
rect 2463 2224 2467 2228
rect 2607 2224 2611 2228
rect 2759 2224 2763 2228
rect 1631 2219 1635 2223
rect 551 2212 555 2216
rect 679 2212 683 2216
rect 807 2212 811 2216
rect 927 2212 931 2216
rect 1047 2212 1051 2216
rect 1159 2212 1163 2216
rect 1271 2212 1275 2216
rect 1391 2212 1395 2216
rect 1927 2208 1931 2212
rect 2103 2208 2107 2212
rect 2295 2208 2299 2212
rect 2503 2208 2507 2212
rect 2719 2208 2723 2212
rect 2951 2208 2955 2212
rect 3159 2208 3163 2212
rect 1671 2201 1675 2205
rect 3191 2201 3195 2205
rect 455 2192 459 2196
rect 583 2192 587 2196
rect 703 2192 707 2196
rect 823 2192 827 2196
rect 943 2192 947 2196
rect 1055 2192 1059 2196
rect 1167 2192 1171 2196
rect 1287 2192 1291 2196
rect 2023 2191 2027 2195
rect 111 2185 115 2189
rect 1631 2185 1635 2189
rect 1671 2183 1675 2187
rect 2119 2187 2123 2191
rect 2175 2187 2179 2191
rect 1927 2179 1931 2183
rect 2023 2179 2027 2183
rect 2103 2179 2107 2183
rect 2295 2179 2299 2183
rect 2303 2179 2304 2183
rect 2304 2179 2307 2183
rect 2503 2179 2507 2183
rect 111 2167 115 2171
rect 455 2163 459 2167
rect 463 2163 464 2167
rect 464 2163 467 2167
rect 583 2163 587 2167
rect 607 2163 611 2167
rect 703 2163 707 2167
rect 711 2163 712 2167
rect 712 2163 715 2167
rect 823 2163 827 2167
rect 863 2163 867 2167
rect 943 2163 947 2167
rect 951 2163 952 2167
rect 952 2163 955 2167
rect 975 2163 979 2167
rect 1055 2163 1059 2167
rect 1063 2167 1064 2171
rect 1064 2167 1067 2171
rect 1167 2163 1171 2167
rect 1175 2167 1176 2171
rect 1176 2167 1179 2171
rect 1279 2171 1283 2175
rect 1287 2163 1291 2167
rect 1631 2167 1635 2171
rect 1671 2165 1675 2169
rect 1847 2169 1851 2173
rect 1999 2169 2003 2173
rect 2023 2167 2027 2171
rect 2151 2169 2155 2173
rect 2175 2167 2179 2171
rect 2295 2169 2299 2173
rect 2447 2169 2451 2173
rect 2303 2163 2304 2167
rect 2304 2163 2307 2167
rect 2471 2167 2475 2171
rect 2599 2169 2603 2173
rect 2615 2179 2619 2183
rect 2719 2179 2723 2183
rect 2727 2183 2728 2187
rect 2728 2183 2731 2187
rect 2767 2183 2771 2187
rect 2951 2179 2955 2183
rect 2959 2183 2960 2187
rect 2960 2183 2963 2187
rect 2991 2183 2995 2187
rect 3159 2179 3163 2183
rect 3167 2179 3168 2183
rect 3168 2179 3171 2183
rect 3191 2183 3195 2187
rect 3191 2165 3195 2169
rect 1671 2147 1675 2151
rect 3191 2147 3195 2151
rect 111 2137 115 2141
rect 351 2141 355 2145
rect 479 2141 483 2145
rect 599 2141 603 2145
rect 719 2141 723 2145
rect 839 2141 843 2145
rect 951 2141 955 2145
rect 1063 2141 1067 2145
rect 1183 2141 1187 2145
rect 383 2135 387 2139
rect 463 2135 467 2139
rect 607 2135 608 2139
rect 608 2135 611 2139
rect 711 2135 715 2139
rect 863 2135 867 2139
rect 975 2135 979 2139
rect 1071 2135 1072 2139
rect 1072 2135 1075 2139
rect 1175 2135 1179 2139
rect 1631 2137 1635 2141
rect 1847 2140 1851 2144
rect 1999 2140 2003 2144
rect 2151 2140 2155 2144
rect 2295 2140 2299 2144
rect 2447 2140 2451 2144
rect 2599 2140 2603 2144
rect 1759 2124 1763 2128
rect 111 2119 115 2123
rect 1911 2124 1915 2128
rect 2071 2124 2075 2128
rect 2255 2124 2259 2128
rect 2463 2124 2467 2128
rect 2687 2124 2691 2128
rect 2927 2124 2931 2128
rect 3159 2124 3163 2128
rect 1631 2119 1635 2123
rect 1671 2117 1675 2121
rect 351 2112 355 2116
rect 479 2112 483 2116
rect 599 2112 603 2116
rect 719 2112 723 2116
rect 839 2112 843 2116
rect 951 2112 955 2116
rect 1063 2112 1067 2116
rect 3191 2117 3195 2121
rect 1183 2112 1187 2116
rect 1671 2099 1675 2103
rect 1759 2095 1763 2099
rect 247 2088 251 2092
rect 375 2088 379 2092
rect 503 2088 507 2092
rect 623 2088 627 2092
rect 743 2088 747 2092
rect 855 2088 859 2092
rect 967 2088 971 2092
rect 1087 2088 1091 2092
rect 111 2081 115 2085
rect 1631 2081 1635 2085
rect 1671 2081 1675 2085
rect 1695 2085 1699 2089
rect 1823 2085 1827 2089
rect 1911 2095 1915 2099
rect 1703 2079 1704 2083
rect 1704 2079 1707 2083
rect 1967 2085 1971 2089
rect 2071 2095 2075 2099
rect 2119 2099 2123 2103
rect 2255 2095 2259 2099
rect 2303 2095 2307 2099
rect 2463 2095 2467 2099
rect 2471 2099 2472 2103
rect 2472 2099 2475 2103
rect 2687 2095 2691 2099
rect 2727 2099 2731 2103
rect 2927 2095 2931 2099
rect 2959 2099 2963 2103
rect 3159 2095 3163 2099
rect 3167 2095 3168 2099
rect 3168 2095 3171 2099
rect 3191 2099 3195 2103
rect 2023 2083 2027 2087
rect 2111 2085 2115 2089
rect 2119 2083 2120 2087
rect 2120 2083 2123 2087
rect 2255 2085 2259 2089
rect 2407 2085 2411 2089
rect 2247 2079 2251 2083
rect 2415 2083 2416 2087
rect 2416 2083 2419 2087
rect 2471 2083 2475 2087
rect 3191 2081 3195 2085
rect 111 2063 115 2067
rect 607 2067 611 2071
rect 247 2059 251 2063
rect 255 2059 256 2063
rect 256 2059 259 2063
rect 375 2059 379 2063
rect 383 2059 384 2063
rect 384 2059 387 2063
rect 503 2059 507 2063
rect 567 2059 571 2063
rect 623 2059 627 2063
rect 1071 2067 1075 2071
rect 743 2059 747 2063
rect 767 2059 771 2063
rect 855 2059 859 2063
rect 863 2059 864 2063
rect 864 2059 867 2063
rect 967 2059 971 2063
rect 975 2059 976 2063
rect 976 2059 979 2063
rect 1087 2059 1091 2063
rect 1191 2063 1195 2067
rect 1631 2063 1635 2067
rect 1671 2063 1675 2067
rect 3191 2063 3195 2067
rect 1695 2056 1699 2060
rect 1823 2056 1827 2060
rect 1967 2056 1971 2060
rect 2111 2056 2115 2060
rect 2255 2056 2259 2060
rect 2407 2056 2411 2060
rect 111 2037 115 2041
rect 175 2041 179 2045
rect 367 2041 371 2045
rect 559 2041 563 2045
rect 759 2041 763 2045
rect 967 2041 971 2045
rect 1183 2041 1187 2045
rect 183 2035 184 2039
rect 184 2035 187 2039
rect 376 2035 380 2039
rect 567 2035 568 2039
rect 568 2035 571 2039
rect 767 2035 768 2039
rect 768 2035 771 2039
rect 919 2035 923 2039
rect 975 2035 976 2039
rect 976 2035 979 2039
rect 1191 2039 1192 2043
rect 1192 2039 1195 2043
rect 1399 2041 1403 2045
rect 1599 2041 1603 2045
rect 1695 2044 1699 2048
rect 2039 2044 2043 2048
rect 2407 2044 2411 2048
rect 2767 2044 2771 2048
rect 3135 2044 3139 2048
rect 1411 2035 1412 2039
rect 1412 2035 1415 2039
rect 1631 2037 1635 2041
rect 1671 2037 1675 2041
rect 3191 2037 3195 2041
rect 1611 2031 1615 2035
rect 1703 2031 1707 2035
rect 111 2019 115 2023
rect 1631 2019 1635 2023
rect 1671 2019 1675 2023
rect 175 2012 179 2016
rect 367 2012 371 2016
rect 559 2012 563 2016
rect 759 2012 763 2016
rect 967 2012 971 2016
rect 1183 2012 1187 2016
rect 1399 2012 1403 2016
rect 1599 2012 1603 2016
rect 1695 2015 1699 2019
rect 1703 2019 1704 2023
rect 1704 2019 1707 2023
rect 2023 2023 2027 2027
rect 2039 2015 2043 2019
rect 2407 2015 2411 2019
rect 2415 2019 2416 2023
rect 2416 2019 2419 2023
rect 2727 2023 2731 2027
rect 2767 2015 2771 2019
rect 2855 2019 2859 2023
rect 3135 2015 3139 2019
rect 3143 2015 3144 2019
rect 3144 2015 3147 2019
rect 3191 2019 3195 2023
rect 135 2000 139 2004
rect 231 2000 235 2004
rect 351 2000 355 2004
rect 463 2000 467 2004
rect 575 2000 579 2004
rect 687 2000 691 2004
rect 799 2000 803 2004
rect 911 2000 915 2004
rect 111 1993 115 1997
rect 1631 1993 1635 1997
rect 1671 1993 1675 1997
rect 2263 1997 2267 2001
rect 2415 1997 2419 2001
rect 2247 1991 2251 1995
rect 2423 1995 2424 1999
rect 2424 1995 2427 1999
rect 2559 1997 2563 2001
rect 2703 1997 2707 2001
rect 2551 1991 2555 1995
rect 2727 1995 2731 1999
rect 2839 1997 2843 2001
rect 2975 1997 2979 2001
rect 3111 1997 3115 2001
rect 2859 1991 2863 1995
rect 3007 1991 3011 1995
rect 3143 1991 3147 1995
rect 3167 1991 3171 1995
rect 3191 1993 3195 1997
rect 111 1975 115 1979
rect 183 1979 187 1983
rect 135 1971 139 1975
rect 143 1971 144 1975
rect 144 1971 147 1975
rect 231 1971 235 1975
rect 255 1979 259 1983
rect 351 1971 355 1975
rect 375 1979 379 1983
rect 463 1971 467 1975
rect 567 1979 571 1983
rect 575 1971 579 1975
rect 687 1971 691 1975
rect 799 1971 803 1975
rect 911 1971 915 1975
rect 919 1971 920 1975
rect 920 1971 923 1975
rect 1631 1975 1635 1979
rect 1671 1975 1675 1979
rect 3191 1975 3195 1979
rect 767 1963 771 1967
rect 2263 1968 2267 1972
rect 2415 1968 2419 1972
rect 2559 1968 2563 1972
rect 2703 1968 2707 1972
rect 2839 1968 2843 1972
rect 2975 1968 2979 1972
rect 3111 1968 3115 1972
rect 863 1959 867 1963
rect 111 1949 115 1953
rect 727 1953 731 1957
rect 855 1953 859 1957
rect 767 1947 771 1951
rect 887 1951 891 1955
rect 983 1953 987 1957
rect 1103 1953 1107 1957
rect 1223 1953 1227 1957
rect 1335 1953 1339 1957
rect 1447 1953 1451 1957
rect 1567 1953 1571 1957
rect 2239 1956 2243 1960
rect 919 1947 923 1951
rect 1007 1947 1011 1951
rect 1127 1947 1131 1951
rect 1243 1943 1247 1947
rect 1355 1943 1359 1947
rect 1411 1947 1415 1951
rect 1471 1947 1475 1951
rect 2391 1956 2395 1960
rect 2543 1956 2547 1960
rect 2695 1956 2699 1960
rect 2847 1956 2851 1960
rect 2999 1956 3003 1960
rect 1611 1951 1615 1955
rect 1631 1949 1635 1953
rect 1671 1949 1675 1953
rect 3191 1949 3195 1953
rect 111 1931 115 1935
rect 1631 1931 1635 1935
rect 1671 1931 1675 1935
rect 727 1924 731 1928
rect 855 1924 859 1928
rect 983 1924 987 1928
rect 1103 1924 1107 1928
rect 1223 1924 1227 1928
rect 1335 1924 1339 1928
rect 1447 1924 1451 1928
rect 1567 1924 1571 1928
rect 2239 1927 2243 1931
rect 2247 1927 2248 1931
rect 2248 1927 2251 1931
rect 2391 1927 2395 1931
rect 2423 1931 2427 1935
rect 2543 1927 2547 1931
rect 2551 1931 2552 1935
rect 2552 1931 2555 1935
rect 2695 1927 2699 1931
rect 2703 1931 2704 1935
rect 2704 1931 2707 1935
rect 2727 1931 2731 1935
rect 2847 1927 2851 1931
rect 2855 1931 2856 1935
rect 2856 1931 2859 1935
rect 2999 1927 3003 1931
rect 3007 1931 3008 1935
rect 3008 1931 3011 1935
rect 3191 1931 3195 1935
rect 1671 1909 1675 1913
rect 2151 1913 2155 1917
rect 2311 1913 2315 1917
rect 2471 1913 2475 1917
rect 2639 1913 2643 1917
rect 2159 1907 2160 1911
rect 2160 1907 2163 1911
rect 2247 1907 2251 1911
rect 2423 1907 2427 1911
rect 2703 1911 2707 1915
rect 2815 1913 2819 1917
rect 2823 1911 2824 1915
rect 2824 1911 2827 1915
rect 2855 1911 2859 1915
rect 2999 1913 3003 1917
rect 3007 1911 3008 1915
rect 3008 1911 3011 1915
rect 3159 1913 3163 1917
rect 3167 1911 3168 1915
rect 3168 1911 3171 1915
rect 3191 1909 3195 1913
rect 631 1900 635 1904
rect 759 1900 763 1904
rect 879 1900 883 1904
rect 999 1900 1003 1904
rect 1119 1900 1123 1904
rect 1231 1900 1235 1904
rect 1343 1900 1347 1904
rect 1463 1900 1467 1904
rect 111 1893 115 1897
rect 1631 1893 1635 1897
rect 1671 1891 1675 1895
rect 3191 1891 3195 1895
rect 2151 1884 2155 1888
rect 2311 1884 2315 1888
rect 2471 1884 2475 1888
rect 2639 1884 2643 1888
rect 2815 1884 2819 1888
rect 2999 1884 3003 1888
rect 3159 1884 3163 1888
rect 111 1875 115 1879
rect 631 1871 635 1875
rect 639 1871 640 1875
rect 640 1871 643 1875
rect 759 1871 763 1875
rect 767 1871 768 1875
rect 768 1871 771 1875
rect 879 1871 883 1875
rect 887 1875 888 1879
rect 888 1875 891 1879
rect 999 1871 1003 1875
rect 1007 1875 1008 1879
rect 1008 1875 1011 1879
rect 1119 1871 1123 1875
rect 1127 1875 1128 1879
rect 1128 1875 1131 1879
rect 1231 1871 1235 1875
rect 1243 1875 1244 1879
rect 1244 1875 1247 1879
rect 1255 1875 1259 1879
rect 1343 1871 1347 1875
rect 1355 1875 1356 1879
rect 1356 1875 1359 1879
rect 1463 1871 1467 1875
rect 1471 1875 1472 1879
rect 1472 1875 1475 1879
rect 1631 1875 1635 1879
rect 2071 1868 2075 1872
rect 2239 1868 2243 1872
rect 2415 1868 2419 1872
rect 2599 1868 2603 1872
rect 2791 1868 2795 1872
rect 2983 1868 2987 1872
rect 3159 1868 3163 1872
rect 1671 1861 1675 1865
rect 3191 1861 3195 1865
rect 111 1845 115 1849
rect 527 1849 531 1853
rect 639 1847 643 1851
rect 655 1849 659 1853
rect 775 1849 779 1853
rect 895 1849 899 1853
rect 1015 1849 1019 1853
rect 1127 1849 1131 1853
rect 687 1843 691 1847
rect 767 1843 771 1847
rect 807 1843 811 1847
rect 887 1843 891 1847
rect 927 1843 931 1847
rect 1007 1843 1011 1847
rect 1039 1843 1043 1847
rect 1135 1847 1136 1851
rect 1136 1847 1139 1851
rect 1247 1849 1251 1853
rect 1255 1847 1256 1851
rect 1256 1847 1259 1851
rect 1367 1849 1371 1853
rect 1355 1843 1359 1847
rect 1631 1845 1635 1849
rect 1671 1843 1675 1847
rect 2159 1847 2163 1851
rect 2247 1847 2251 1851
rect 2071 1839 2075 1843
rect 2079 1839 2080 1843
rect 2080 1839 2083 1843
rect 2239 1839 2243 1843
rect 2415 1839 2419 1843
rect 2423 1843 2424 1847
rect 2424 1843 2427 1847
rect 2551 1847 2555 1851
rect 2591 1847 2595 1851
rect 2599 1839 2603 1843
rect 2791 1839 2795 1843
rect 2823 1843 2827 1847
rect 111 1827 115 1831
rect 1631 1827 1635 1831
rect 1671 1825 1675 1829
rect 1983 1829 1987 1833
rect 2135 1829 2139 1833
rect 2287 1829 2291 1833
rect 2431 1829 2435 1833
rect 2583 1829 2587 1833
rect 527 1820 531 1824
rect 655 1820 659 1824
rect 775 1820 779 1824
rect 895 1820 899 1824
rect 1015 1820 1019 1824
rect 1127 1820 1131 1824
rect 1247 1820 1251 1824
rect 1367 1820 1371 1824
rect 1991 1823 1992 1827
rect 1992 1823 1995 1827
rect 2087 1823 2091 1827
rect 2159 1823 2163 1827
rect 2247 1823 2251 1827
rect 2423 1823 2427 1827
rect 2495 1823 2499 1827
rect 2591 1827 2592 1831
rect 2592 1827 2595 1831
rect 2735 1829 2739 1833
rect 2743 1827 2744 1831
rect 2744 1827 2747 1831
rect 2983 1839 2987 1843
rect 3007 1843 3011 1847
rect 3159 1839 3163 1843
rect 3167 1843 3168 1847
rect 3168 1843 3171 1847
rect 3191 1843 3195 1847
rect 3191 1825 3195 1829
rect 1671 1807 1675 1811
rect 3191 1807 3195 1811
rect 423 1800 427 1804
rect 551 1800 555 1804
rect 679 1800 683 1804
rect 799 1800 803 1804
rect 919 1800 923 1804
rect 1031 1800 1035 1804
rect 1143 1800 1147 1804
rect 1263 1800 1267 1804
rect 1983 1800 1987 1804
rect 2135 1800 2139 1804
rect 2287 1800 2291 1804
rect 2431 1800 2435 1804
rect 2583 1800 2587 1804
rect 2735 1800 2739 1804
rect 111 1793 115 1797
rect 1631 1793 1635 1797
rect 1903 1788 1907 1792
rect 2079 1788 2083 1792
rect 2271 1788 2275 1792
rect 2487 1788 2491 1792
rect 2711 1788 2715 1792
rect 2943 1788 2947 1792
rect 3159 1788 3163 1792
rect 111 1775 115 1779
rect 423 1771 427 1775
rect 431 1771 432 1775
rect 432 1771 435 1775
rect 551 1771 555 1775
rect 559 1771 560 1775
rect 560 1771 563 1775
rect 679 1771 683 1775
rect 687 1775 688 1779
rect 688 1775 691 1779
rect 799 1771 803 1775
rect 807 1775 808 1779
rect 808 1775 811 1779
rect 919 1771 923 1775
rect 927 1775 928 1779
rect 928 1775 931 1779
rect 1031 1771 1035 1775
rect 1039 1775 1040 1779
rect 1040 1775 1043 1779
rect 1135 1779 1139 1783
rect 1143 1771 1147 1775
rect 1255 1779 1259 1783
rect 1671 1781 1675 1785
rect 3191 1781 3195 1785
rect 1263 1771 1267 1775
rect 1631 1775 1635 1779
rect 1671 1763 1675 1767
rect 1903 1759 1907 1763
rect 1991 1763 1995 1767
rect 2087 1767 2091 1771
rect 2079 1759 2083 1763
rect 2247 1767 2251 1771
rect 2271 1759 2275 1763
rect 2487 1759 2491 1763
rect 2495 1763 2496 1767
rect 2496 1763 2499 1767
rect 2711 1759 2715 1763
rect 2743 1763 2747 1767
rect 2943 1759 2947 1763
rect 2951 1763 2952 1767
rect 2952 1763 2955 1767
rect 3007 1763 3011 1767
rect 3159 1759 3163 1763
rect 3167 1763 3168 1767
rect 3168 1763 3171 1767
rect 3191 1763 3195 1767
rect 111 1745 115 1749
rect 327 1749 331 1753
rect 455 1749 459 1753
rect 575 1749 579 1753
rect 695 1749 699 1753
rect 815 1749 819 1753
rect 335 1743 336 1747
rect 336 1743 339 1747
rect 431 1743 435 1747
rect 559 1743 563 1747
rect 719 1743 723 1747
rect 823 1745 824 1747
rect 824 1745 827 1747
rect 927 1749 931 1753
rect 1039 1749 1043 1753
rect 1159 1749 1163 1753
rect 823 1743 827 1745
rect 951 1743 955 1747
rect 1167 1743 1168 1747
rect 1168 1743 1171 1747
rect 1631 1745 1635 1749
rect 1671 1737 1675 1741
rect 1815 1741 1819 1745
rect 1967 1741 1971 1745
rect 2127 1741 2131 1745
rect 2303 1741 2307 1745
rect 2503 1741 2507 1745
rect 2711 1741 2715 1745
rect 2935 1741 2939 1745
rect 3159 1741 3163 1745
rect 1823 1735 1824 1739
rect 1824 1735 1827 1739
rect 2031 1735 2035 1739
rect 2323 1735 2327 1739
rect 2475 1735 2479 1739
rect 2719 1735 2720 1739
rect 2720 1735 2723 1739
rect 2944 1735 2948 1739
rect 3167 1739 3168 1743
rect 3168 1739 3171 1743
rect 3191 1737 3195 1741
rect 111 1727 115 1731
rect 1631 1727 1635 1731
rect 327 1720 331 1724
rect 455 1720 459 1724
rect 575 1720 579 1724
rect 695 1720 699 1724
rect 815 1720 819 1724
rect 927 1720 931 1724
rect 1039 1720 1043 1724
rect 1159 1720 1163 1724
rect 1671 1719 1675 1723
rect 3191 1719 3195 1723
rect 1815 1712 1819 1716
rect 1967 1712 1971 1716
rect 2127 1712 2131 1716
rect 2303 1712 2307 1716
rect 2503 1712 2507 1716
rect 2711 1712 2715 1716
rect 2935 1712 2939 1716
rect 3159 1712 3163 1716
rect 223 1696 227 1700
rect 351 1696 355 1700
rect 471 1696 475 1700
rect 591 1696 595 1700
rect 711 1696 715 1700
rect 823 1696 827 1700
rect 943 1696 947 1700
rect 1063 1696 1067 1700
rect 1735 1700 1739 1704
rect 1879 1700 1883 1704
rect 2023 1700 2027 1704
rect 2167 1700 2171 1704
rect 2311 1700 2315 1704
rect 2463 1700 2467 1704
rect 111 1689 115 1693
rect 1631 1689 1635 1693
rect 1671 1693 1675 1697
rect 3191 1693 3195 1697
rect 111 1671 115 1675
rect 223 1667 227 1671
rect 231 1667 232 1671
rect 232 1667 235 1671
rect 351 1667 355 1671
rect 471 1667 475 1671
rect 479 1667 480 1671
rect 480 1667 483 1671
rect 591 1667 595 1671
rect 599 1667 600 1671
rect 600 1667 603 1671
rect 711 1667 715 1671
rect 719 1671 720 1675
rect 720 1671 723 1675
rect 823 1667 827 1671
rect 831 1671 832 1675
rect 832 1671 835 1675
rect 927 1675 931 1679
rect 943 1667 947 1671
rect 951 1671 952 1675
rect 952 1671 955 1675
rect 1063 1667 1067 1671
rect 1071 1667 1072 1671
rect 1072 1667 1075 1671
rect 1631 1671 1635 1675
rect 1671 1675 1675 1679
rect 1823 1679 1827 1683
rect 1735 1671 1739 1675
rect 1823 1671 1827 1675
rect 1879 1671 1883 1675
rect 311 1659 315 1663
rect 335 1659 339 1663
rect 1671 1657 1675 1661
rect 1695 1661 1699 1665
rect 1895 1661 1899 1665
rect 2023 1671 2027 1675
rect 2031 1675 2032 1679
rect 2032 1675 2035 1679
rect 2107 1675 2111 1679
rect 2167 1671 2171 1675
rect 2311 1671 2315 1675
rect 2323 1675 2324 1679
rect 2324 1675 2327 1679
rect 2463 1671 2467 1675
rect 2475 1675 2476 1679
rect 2476 1675 2479 1679
rect 3191 1675 3195 1679
rect 2127 1661 2131 1665
rect 111 1641 115 1645
rect 135 1645 139 1649
rect 247 1645 251 1649
rect 383 1645 387 1649
rect 2107 1655 2111 1659
rect 2367 1661 2371 1665
rect 2615 1661 2619 1665
rect 2871 1661 2875 1665
rect 3135 1661 3139 1665
rect 2323 1655 2327 1659
rect 2399 1655 2403 1659
rect 2719 1655 2723 1659
rect 2919 1655 2923 1659
rect 3143 1659 3144 1663
rect 3144 1659 3147 1663
rect 3167 1659 3171 1663
rect 3191 1657 3195 1661
rect 143 1639 144 1643
rect 144 1639 147 1643
rect 231 1639 235 1643
rect 311 1639 315 1643
rect 479 1643 483 1647
rect 535 1645 539 1649
rect 711 1645 715 1649
rect 599 1639 603 1643
rect 719 1643 720 1647
rect 720 1643 723 1647
rect 919 1645 923 1649
rect 927 1643 928 1647
rect 928 1643 931 1647
rect 1143 1645 1147 1649
rect 1167 1643 1171 1647
rect 1383 1645 1387 1649
rect 1599 1645 1603 1649
rect 1423 1639 1427 1643
rect 1607 1643 1608 1647
rect 1608 1643 1611 1647
rect 1631 1641 1635 1645
rect 1671 1639 1675 1643
rect 3191 1639 3195 1643
rect 1695 1632 1699 1636
rect 1895 1632 1899 1636
rect 2127 1632 2131 1636
rect 2367 1632 2371 1636
rect 2615 1632 2619 1636
rect 2871 1632 2875 1636
rect 3135 1632 3139 1636
rect 111 1623 115 1627
rect 1631 1623 1635 1627
rect 135 1616 139 1620
rect 247 1616 251 1620
rect 383 1616 387 1620
rect 535 1616 539 1620
rect 711 1616 715 1620
rect 919 1616 923 1620
rect 1143 1616 1147 1620
rect 1383 1616 1387 1620
rect 1599 1616 1603 1620
rect 2319 1616 2323 1620
rect 2519 1616 2523 1620
rect 2711 1616 2715 1620
rect 2911 1616 2915 1620
rect 3111 1616 3115 1620
rect 1671 1609 1675 1613
rect 3191 1609 3195 1613
rect 135 1596 139 1600
rect 303 1596 307 1600
rect 503 1596 507 1600
rect 695 1596 699 1600
rect 887 1596 891 1600
rect 1063 1596 1067 1600
rect 1239 1596 1243 1600
rect 1415 1596 1419 1600
rect 1591 1596 1595 1600
rect 111 1589 115 1593
rect 1631 1589 1635 1593
rect 1671 1591 1675 1595
rect 2319 1587 2323 1591
rect 2519 1587 2523 1591
rect 2527 1587 2528 1591
rect 2528 1587 2531 1591
rect 2711 1587 2715 1591
rect 2719 1587 2720 1591
rect 2720 1587 2723 1591
rect 2911 1587 2915 1591
rect 2919 1587 2920 1591
rect 2920 1587 2923 1591
rect 3007 1587 3011 1591
rect 3111 1587 3115 1591
rect 3119 1591 3120 1595
rect 3120 1591 3123 1595
rect 3143 1591 3147 1595
rect 3191 1591 3195 1595
rect 111 1571 115 1575
rect 135 1567 139 1571
rect 143 1571 144 1575
rect 144 1571 147 1575
rect 303 1567 307 1571
rect 311 1571 312 1575
rect 312 1571 315 1575
rect 479 1575 483 1579
rect 503 1567 507 1571
rect 695 1567 699 1571
rect 719 1571 723 1575
rect 887 1567 891 1571
rect 895 1567 896 1571
rect 896 1567 899 1571
rect 927 1567 931 1571
rect 1063 1567 1067 1571
rect 1071 1571 1072 1575
rect 1072 1571 1075 1575
rect 1167 1575 1171 1579
rect 1239 1567 1243 1571
rect 1287 1571 1291 1575
rect 1415 1567 1419 1571
rect 1423 1567 1424 1571
rect 1424 1567 1427 1571
rect 1591 1567 1595 1571
rect 1600 1567 1604 1571
rect 1631 1571 1635 1575
rect 1671 1573 1675 1577
rect 2271 1577 2275 1581
rect 2291 1579 2295 1583
rect 2415 1577 2419 1581
rect 2559 1577 2563 1581
rect 2695 1577 2699 1581
rect 2839 1577 2843 1581
rect 2983 1577 2987 1581
rect 2399 1571 2403 1575
rect 2527 1571 2531 1575
rect 2663 1571 2667 1575
rect 2719 1571 2723 1575
rect 2919 1571 2923 1575
rect 3007 1571 3011 1575
rect 3191 1573 3195 1577
rect 1671 1555 1675 1559
rect 3191 1555 3195 1559
rect 111 1541 115 1545
rect 679 1545 683 1549
rect 719 1543 723 1547
rect 807 1545 811 1549
rect 927 1545 931 1549
rect 1047 1545 1051 1549
rect 839 1539 843 1543
rect 895 1539 899 1543
rect 1071 1543 1075 1547
rect 1167 1545 1171 1549
rect 1175 1543 1176 1547
rect 1176 1543 1179 1547
rect 1191 1543 1195 1547
rect 1279 1545 1283 1549
rect 1287 1543 1288 1547
rect 1288 1543 1291 1547
rect 1399 1545 1403 1549
rect 1519 1545 1523 1549
rect 2271 1548 2275 1552
rect 2415 1548 2419 1552
rect 2559 1548 2563 1552
rect 2695 1548 2699 1552
rect 2839 1548 2843 1552
rect 2983 1548 2987 1552
rect 1407 1539 1408 1543
rect 1408 1539 1411 1543
rect 1423 1539 1427 1543
rect 1599 1539 1603 1543
rect 1631 1541 1635 1545
rect 2167 1528 2171 1532
rect 111 1523 115 1527
rect 2279 1528 2283 1532
rect 2391 1528 2395 1532
rect 2503 1528 2507 1532
rect 2615 1528 2619 1532
rect 2735 1528 2739 1532
rect 2855 1528 2859 1532
rect 2983 1528 2987 1532
rect 3111 1528 3115 1532
rect 1631 1523 1635 1527
rect 1671 1521 1675 1525
rect 679 1516 683 1520
rect 807 1516 811 1520
rect 927 1516 931 1520
rect 1047 1516 1051 1520
rect 1167 1516 1171 1520
rect 1279 1516 1283 1520
rect 1399 1516 1403 1520
rect 3191 1521 3195 1525
rect 1519 1516 1523 1520
rect 1671 1503 1675 1507
rect 575 1496 579 1500
rect 703 1496 707 1500
rect 831 1496 835 1500
rect 951 1496 955 1500
rect 1071 1496 1075 1500
rect 1183 1496 1187 1500
rect 1295 1496 1299 1500
rect 1415 1496 1419 1500
rect 2167 1499 2171 1503
rect 2279 1499 2283 1503
rect 2291 1503 2292 1507
rect 2292 1503 2295 1507
rect 2391 1499 2395 1503
rect 2399 1503 2400 1507
rect 2400 1503 2403 1507
rect 2527 1507 2531 1511
rect 2503 1499 2507 1503
rect 2527 1499 2531 1503
rect 2615 1499 2619 1503
rect 2663 1503 2667 1507
rect 2735 1499 2739 1503
rect 2807 1503 2811 1507
rect 2855 1499 2859 1503
rect 2863 1503 2864 1507
rect 2864 1503 2867 1507
rect 2919 1503 2923 1507
rect 2983 1499 2987 1503
rect 3007 1499 3011 1503
rect 3111 1499 3115 1503
rect 3119 1503 3120 1507
rect 3120 1503 3123 1507
rect 3191 1503 3195 1507
rect 111 1489 115 1493
rect 1631 1489 1635 1493
rect 2107 1491 2111 1495
rect 2399 1491 2403 1495
rect 2487 1491 2491 1495
rect 1671 1481 1675 1485
rect 2087 1485 2091 1489
rect 2231 1485 2235 1489
rect 111 1471 115 1475
rect 1287 1475 1291 1479
rect 575 1467 579 1471
rect 587 1467 588 1471
rect 588 1467 591 1471
rect 703 1467 707 1471
rect 735 1467 739 1471
rect 831 1467 835 1471
rect 839 1467 840 1471
rect 840 1467 843 1471
rect 951 1467 955 1471
rect 959 1467 960 1471
rect 960 1467 963 1471
rect 1071 1467 1075 1471
rect 1079 1467 1080 1471
rect 1080 1467 1083 1471
rect 1183 1467 1187 1471
rect 1191 1467 1192 1471
rect 1192 1467 1195 1471
rect 1295 1467 1299 1471
rect 1319 1471 1323 1475
rect 1407 1475 1411 1479
rect 2107 1479 2111 1483
rect 2239 1483 2240 1487
rect 2240 1483 2243 1487
rect 2291 1483 2295 1487
rect 2375 1485 2379 1489
rect 2399 1483 2403 1487
rect 2511 1485 2515 1489
rect 2655 1485 2659 1489
rect 2663 1483 2664 1487
rect 2664 1483 2667 1487
rect 2799 1485 2803 1489
rect 2807 1483 2808 1487
rect 2808 1483 2811 1487
rect 2863 1479 2867 1483
rect 3191 1481 3195 1485
rect 1415 1467 1419 1471
rect 1631 1471 1635 1475
rect 1671 1463 1675 1467
rect 3191 1463 3195 1467
rect 2087 1456 2091 1460
rect 2231 1456 2235 1460
rect 2375 1456 2379 1460
rect 2511 1456 2515 1460
rect 2655 1456 2659 1460
rect 2799 1456 2803 1460
rect 111 1441 115 1445
rect 479 1445 483 1449
rect 607 1445 611 1449
rect 727 1445 731 1449
rect 847 1445 851 1449
rect 967 1445 971 1449
rect 587 1439 591 1443
rect 635 1439 639 1443
rect 735 1439 736 1443
rect 736 1439 739 1443
rect 839 1439 843 1443
rect 887 1439 891 1443
rect 959 1439 963 1443
rect 1079 1445 1083 1449
rect 1191 1445 1195 1449
rect 1087 1439 1088 1443
rect 1088 1439 1091 1443
rect 1103 1439 1107 1443
rect 1199 1443 1200 1447
rect 1200 1443 1203 1447
rect 1311 1445 1315 1449
rect 1319 1443 1320 1447
rect 1320 1443 1323 1447
rect 1631 1441 1635 1445
rect 1983 1440 1987 1444
rect 2095 1440 2099 1444
rect 2207 1440 2211 1444
rect 2335 1440 2339 1444
rect 2479 1440 2483 1444
rect 2639 1440 2643 1444
rect 2815 1440 2819 1444
rect 2999 1440 3003 1444
rect 3159 1440 3163 1444
rect 1671 1433 1675 1437
rect 3191 1433 3195 1437
rect 111 1423 115 1427
rect 1631 1423 1635 1427
rect 479 1416 483 1420
rect 607 1416 611 1420
rect 727 1416 731 1420
rect 847 1416 851 1420
rect 967 1416 971 1420
rect 1079 1416 1083 1420
rect 1191 1416 1195 1420
rect 1311 1416 1315 1420
rect 1671 1415 1675 1419
rect 2107 1417 2108 1419
rect 2108 1417 2111 1419
rect 1983 1411 1987 1415
rect 1991 1411 1992 1415
rect 1992 1411 1995 1415
rect 2095 1411 2099 1415
rect 2107 1415 2111 1417
rect 2207 1411 2211 1415
rect 2239 1419 2243 1423
rect 2335 1411 2339 1415
rect 2399 1415 2403 1419
rect 2479 1411 2483 1415
rect 2487 1415 2488 1419
rect 2488 1415 2491 1419
rect 2639 1411 2643 1415
rect 2663 1415 2667 1419
rect 2815 1411 2819 1415
rect 2823 1411 2824 1415
rect 2824 1411 2827 1415
rect 2863 1415 2867 1419
rect 3007 1419 3011 1423
rect 2999 1411 3003 1415
rect 3119 1419 3123 1423
rect 3159 1411 3163 1415
rect 3167 1415 3168 1419
rect 3168 1415 3171 1419
rect 3191 1415 3195 1419
rect 375 1392 379 1396
rect 503 1392 507 1396
rect 623 1392 627 1396
rect 743 1392 747 1396
rect 863 1392 867 1396
rect 975 1392 979 1396
rect 1095 1392 1099 1396
rect 1215 1392 1219 1396
rect 111 1385 115 1389
rect 1631 1385 1635 1389
rect 1671 1381 1675 1385
rect 1879 1385 1883 1389
rect 1991 1385 1995 1389
rect 2103 1385 2107 1389
rect 2239 1385 2243 1389
rect 1887 1379 1888 1383
rect 1888 1379 1891 1383
rect 1999 1379 2000 1383
rect 2000 1379 2003 1383
rect 2111 1379 2112 1383
rect 2112 1379 2115 1383
rect 2247 1383 2248 1387
rect 2248 1383 2251 1387
rect 2391 1385 2395 1389
rect 2399 1383 2400 1387
rect 2400 1383 2403 1387
rect 2567 1385 2571 1389
rect 2663 1383 2667 1387
rect 2767 1385 2771 1389
rect 2823 1383 2827 1387
rect 2975 1385 2979 1389
rect 2983 1383 2984 1387
rect 2984 1383 2987 1387
rect 3007 1383 3011 1387
rect 3159 1385 3163 1389
rect 3167 1383 3168 1387
rect 3168 1383 3171 1387
rect 3191 1381 3195 1385
rect 111 1367 115 1371
rect 375 1363 379 1367
rect 383 1363 384 1367
rect 384 1363 387 1367
rect 503 1363 507 1367
rect 535 1363 539 1367
rect 623 1363 627 1367
rect 635 1363 636 1367
rect 636 1363 639 1367
rect 743 1363 747 1367
rect 787 1363 791 1367
rect 863 1363 867 1367
rect 887 1363 891 1367
rect 975 1363 979 1367
rect 1015 1363 1019 1367
rect 1095 1363 1099 1367
rect 1103 1363 1104 1367
rect 1104 1363 1107 1367
rect 1215 1363 1219 1367
rect 1631 1367 1635 1371
rect 1671 1363 1675 1367
rect 3191 1363 3195 1367
rect 1879 1356 1883 1360
rect 1991 1356 1995 1360
rect 2103 1356 2107 1360
rect 2239 1356 2243 1360
rect 2391 1356 2395 1360
rect 2567 1356 2571 1360
rect 2767 1356 2771 1360
rect 2975 1356 2979 1360
rect 3159 1356 3163 1360
rect 111 1341 115 1345
rect 271 1345 275 1349
rect 399 1345 403 1349
rect 527 1345 531 1349
rect 647 1345 651 1349
rect 767 1345 771 1349
rect 879 1345 883 1349
rect 991 1345 995 1349
rect 1111 1345 1115 1349
rect 311 1339 315 1343
rect 383 1339 387 1343
rect 535 1339 536 1343
rect 536 1339 539 1343
rect 635 1339 639 1343
rect 787 1339 791 1343
rect 888 1339 892 1343
rect 1015 1339 1019 1343
rect 1103 1339 1107 1343
rect 1631 1341 1635 1345
rect 1775 1332 1779 1336
rect 1887 1332 1891 1336
rect 1991 1332 1995 1336
rect 2095 1332 2099 1336
rect 2199 1332 2203 1336
rect 2303 1332 2307 1336
rect 2407 1332 2411 1336
rect 2511 1332 2515 1336
rect 111 1323 115 1327
rect 1631 1323 1635 1327
rect 1671 1325 1675 1329
rect 3191 1325 3195 1329
rect 271 1316 275 1320
rect 399 1316 403 1320
rect 527 1316 531 1320
rect 647 1316 651 1320
rect 767 1316 771 1320
rect 879 1316 883 1320
rect 991 1316 995 1320
rect 1111 1316 1115 1320
rect 1671 1307 1675 1311
rect 1775 1303 1779 1307
rect 1783 1303 1784 1307
rect 1784 1303 1787 1307
rect 1895 1311 1899 1315
rect 1887 1303 1891 1307
rect 1943 1307 1947 1311
rect 1999 1311 2003 1315
rect 2103 1313 2107 1315
rect 1991 1303 1995 1307
rect 2103 1311 2104 1313
rect 2104 1311 2107 1313
rect 2095 1303 2099 1307
rect 2199 1303 2203 1307
rect 2399 1311 2403 1315
rect 2303 1303 2307 1307
rect 2407 1303 2411 1307
rect 2503 1311 2507 1315
rect 2511 1303 2515 1307
rect 3191 1307 3195 1311
rect 175 1292 179 1296
rect 303 1292 307 1296
rect 423 1292 427 1296
rect 543 1292 547 1296
rect 663 1292 667 1296
rect 775 1292 779 1296
rect 887 1292 891 1296
rect 1007 1292 1011 1296
rect 2111 1295 2115 1299
rect 111 1285 115 1289
rect 1631 1285 1635 1289
rect 1671 1281 1675 1285
rect 1695 1285 1699 1289
rect 1791 1285 1795 1289
rect 1935 1285 1939 1289
rect 1703 1279 1704 1283
rect 1704 1279 1707 1283
rect 1783 1279 1787 1283
rect 1943 1283 1944 1287
rect 1944 1283 1947 1287
rect 2103 1285 2107 1289
rect 2111 1283 2112 1287
rect 2112 1283 2115 1287
rect 2295 1285 2299 1289
rect 2495 1285 2499 1289
rect 2503 1283 2504 1287
rect 2504 1283 2507 1287
rect 2711 1285 2715 1289
rect 2935 1285 2939 1289
rect 2719 1279 2720 1283
rect 2720 1279 2723 1283
rect 2983 1283 2987 1287
rect 3159 1285 3163 1289
rect 3167 1283 3168 1287
rect 3168 1283 3171 1287
rect 3191 1281 3195 1285
rect 111 1267 115 1271
rect 175 1263 179 1267
rect 187 1263 188 1267
rect 188 1263 191 1267
rect 303 1263 307 1267
rect 311 1267 312 1271
rect 312 1267 315 1271
rect 423 1263 427 1267
rect 431 1263 432 1267
rect 432 1263 435 1267
rect 543 1263 547 1267
rect 551 1267 552 1271
rect 552 1267 555 1271
rect 635 1267 639 1271
rect 663 1263 667 1267
rect 671 1263 672 1267
rect 672 1263 675 1267
rect 775 1263 779 1267
rect 787 1263 788 1267
rect 788 1263 791 1267
rect 887 1263 891 1267
rect 895 1263 896 1267
rect 896 1263 899 1267
rect 1007 1263 1011 1267
rect 1016 1263 1020 1267
rect 1631 1267 1635 1271
rect 1671 1263 1675 1267
rect 3191 1263 3195 1267
rect 867 1255 871 1259
rect 1695 1256 1699 1260
rect 1791 1256 1795 1260
rect 1935 1256 1939 1260
rect 2103 1256 2107 1260
rect 2295 1256 2299 1260
rect 2495 1256 2499 1260
rect 2711 1256 2715 1260
rect 2935 1256 2939 1260
rect 3159 1256 3163 1260
rect 111 1237 115 1241
rect 135 1241 139 1245
rect 231 1241 235 1245
rect 359 1241 363 1245
rect 503 1241 507 1245
rect 187 1235 191 1239
rect 259 1235 263 1239
rect 311 1235 315 1239
rect 431 1235 435 1239
rect 551 1239 555 1243
rect 663 1241 667 1245
rect 831 1241 835 1245
rect 1015 1241 1019 1245
rect 1207 1241 1211 1245
rect 1407 1241 1411 1245
rect 1599 1241 1603 1245
rect 671 1235 672 1239
rect 672 1235 675 1239
rect 787 1235 791 1239
rect 867 1235 871 1239
rect 1007 1235 1011 1239
rect 1023 1235 1024 1239
rect 1024 1235 1027 1239
rect 1231 1235 1235 1239
rect 1455 1235 1459 1239
rect 1607 1235 1608 1239
rect 1608 1235 1611 1239
rect 1631 1237 1635 1241
rect 1695 1228 1699 1232
rect 1983 1228 1987 1232
rect 2255 1228 2259 1232
rect 2495 1228 2499 1232
rect 2711 1228 2715 1232
rect 2919 1228 2923 1232
rect 3135 1228 3139 1232
rect 111 1219 115 1223
rect 1631 1219 1635 1223
rect 1671 1221 1675 1225
rect 3191 1221 3195 1225
rect 135 1212 139 1216
rect 231 1212 235 1216
rect 359 1212 363 1216
rect 503 1212 507 1216
rect 663 1212 667 1216
rect 831 1212 835 1216
rect 1015 1212 1019 1216
rect 1207 1212 1211 1216
rect 1407 1212 1411 1216
rect 1599 1212 1603 1216
rect 1607 1211 1611 1215
rect 1703 1211 1707 1215
rect 1671 1203 1675 1207
rect 1695 1199 1699 1203
rect 1943 1207 1947 1211
rect 1983 1199 1987 1203
rect 2255 1199 2259 1203
rect 2495 1199 2499 1203
rect 2507 1199 2508 1203
rect 2508 1199 2511 1203
rect 2711 1199 2715 1203
rect 2719 1199 2720 1203
rect 2720 1199 2723 1203
rect 2855 1199 2859 1203
rect 2919 1199 2923 1203
rect 3007 1199 3011 1203
rect 3135 1199 3139 1203
rect 3143 1203 3144 1207
rect 3144 1203 3147 1207
rect 3167 1203 3171 1207
rect 3191 1203 3195 1207
rect 727 1192 731 1196
rect 855 1192 859 1196
rect 983 1192 987 1196
rect 1103 1192 1107 1196
rect 1223 1192 1227 1196
rect 1335 1192 1339 1196
rect 1447 1192 1451 1196
rect 1567 1192 1571 1196
rect 2183 1191 2187 1195
rect 111 1185 115 1189
rect 1631 1185 1635 1189
rect 1671 1181 1675 1185
rect 2247 1185 2251 1189
rect 2399 1185 2403 1189
rect 2551 1185 2555 1189
rect 2695 1185 2699 1189
rect 2507 1179 2511 1183
rect 2703 1183 2704 1187
rect 2704 1183 2707 1187
rect 2847 1185 2851 1189
rect 2855 1183 2856 1187
rect 2856 1183 2859 1187
rect 2999 1185 3003 1189
rect 3007 1179 3008 1183
rect 3008 1179 3011 1183
rect 3191 1181 3195 1185
rect 111 1167 115 1171
rect 727 1163 731 1167
rect 735 1163 736 1167
rect 736 1163 739 1167
rect 855 1163 859 1167
rect 867 1163 868 1167
rect 868 1163 871 1167
rect 983 1163 987 1167
rect 1007 1163 1011 1167
rect 1103 1163 1107 1167
rect 1111 1163 1112 1167
rect 1112 1163 1115 1167
rect 1223 1163 1227 1167
rect 1231 1167 1232 1171
rect 1232 1167 1235 1171
rect 1255 1167 1259 1171
rect 1335 1163 1339 1167
rect 1344 1163 1348 1167
rect 1447 1163 1451 1167
rect 1455 1163 1456 1167
rect 1456 1163 1459 1167
rect 1567 1163 1571 1167
rect 1607 1167 1611 1171
rect 1631 1167 1635 1171
rect 1671 1163 1675 1167
rect 3191 1163 3195 1167
rect 2247 1156 2251 1160
rect 2399 1156 2403 1160
rect 2551 1156 2555 1160
rect 2695 1156 2699 1160
rect 2847 1156 2851 1160
rect 2999 1156 3003 1160
rect 111 1137 115 1141
rect 631 1141 635 1145
rect 759 1141 763 1145
rect 879 1141 883 1145
rect 999 1141 1003 1145
rect 1119 1141 1123 1145
rect 1231 1141 1235 1145
rect 1343 1141 1347 1145
rect 1463 1141 1467 1145
rect 2175 1144 2179 1148
rect 2335 1144 2339 1148
rect 2495 1144 2499 1148
rect 2655 1144 2659 1148
rect 2815 1144 2819 1148
rect 2975 1144 2979 1148
rect 3135 1144 3139 1148
rect 639 1135 640 1139
rect 640 1135 643 1139
rect 671 1135 675 1139
rect 735 1135 739 1139
rect 783 1135 787 1139
rect 867 1135 871 1139
rect 907 1135 911 1139
rect 1007 1135 1008 1139
rect 1008 1135 1011 1139
rect 1111 1135 1115 1139
rect 1128 1135 1132 1139
rect 1255 1135 1259 1139
rect 1351 1135 1352 1139
rect 1352 1135 1355 1139
rect 1455 1135 1459 1139
rect 1631 1137 1635 1141
rect 1671 1137 1675 1141
rect 3191 1137 3195 1141
rect 111 1119 115 1123
rect 1631 1119 1635 1123
rect 1671 1119 1675 1123
rect 631 1112 635 1116
rect 759 1112 763 1116
rect 879 1112 883 1116
rect 999 1112 1003 1116
rect 1119 1112 1123 1116
rect 1231 1112 1235 1116
rect 1343 1112 1347 1116
rect 1463 1112 1467 1116
rect 2175 1115 2179 1119
rect 2183 1115 2184 1119
rect 2184 1115 2187 1119
rect 2335 1115 2339 1119
rect 2495 1115 2499 1119
rect 2507 1119 2508 1123
rect 2508 1119 2511 1123
rect 2655 1115 2659 1119
rect 2663 1119 2664 1123
rect 2664 1119 2667 1123
rect 2703 1119 2707 1123
rect 2815 1115 2819 1119
rect 2823 1119 2824 1123
rect 2824 1119 2827 1123
rect 2855 1119 2859 1123
rect 2975 1115 2979 1119
rect 3007 1119 3011 1123
rect 3135 1115 3139 1119
rect 3143 1119 3144 1123
rect 3144 1119 3147 1123
rect 3191 1119 3195 1123
rect 1671 1097 1675 1101
rect 2071 1101 2075 1105
rect 2191 1101 2195 1105
rect 2327 1101 2331 1105
rect 2079 1095 2080 1099
rect 2080 1095 2083 1099
rect 2183 1095 2187 1099
rect 2351 1099 2352 1103
rect 2352 1099 2355 1103
rect 2479 1101 2483 1105
rect 2507 1099 2511 1103
rect 2639 1101 2643 1105
rect 2663 1099 2667 1103
rect 2815 1101 2819 1105
rect 2823 1099 2824 1103
rect 2824 1099 2827 1103
rect 2999 1101 3003 1105
rect 3159 1101 3163 1105
rect 3007 1095 3008 1099
rect 3008 1095 3011 1099
rect 3143 1095 3147 1099
rect 3167 1095 3168 1099
rect 3168 1095 3171 1099
rect 3191 1097 3195 1101
rect 527 1088 531 1092
rect 655 1088 659 1092
rect 775 1088 779 1092
rect 895 1088 899 1092
rect 1015 1088 1019 1092
rect 1127 1088 1131 1092
rect 1247 1088 1251 1092
rect 1367 1088 1371 1092
rect 111 1081 115 1085
rect 1631 1081 1635 1085
rect 1671 1079 1675 1083
rect 3191 1079 3195 1083
rect 2071 1072 2075 1076
rect 2191 1072 2195 1076
rect 2327 1072 2331 1076
rect 2479 1072 2483 1076
rect 2639 1072 2643 1076
rect 2815 1072 2819 1076
rect 2999 1072 3003 1076
rect 3159 1072 3163 1076
rect 111 1063 115 1067
rect 527 1059 531 1063
rect 535 1059 536 1063
rect 536 1059 539 1063
rect 655 1059 659 1063
rect 775 1059 779 1063
rect 783 1063 784 1067
rect 784 1063 787 1067
rect 895 1059 899 1063
rect 907 1059 908 1063
rect 908 1059 911 1063
rect 1015 1059 1019 1063
rect 1039 1059 1043 1063
rect 1127 1059 1131 1063
rect 1135 1059 1136 1063
rect 1136 1059 1139 1063
rect 1247 1059 1251 1063
rect 1255 1059 1256 1063
rect 1256 1059 1259 1063
rect 1367 1059 1371 1063
rect 1631 1063 1635 1067
rect 583 1051 587 1055
rect 639 1051 643 1055
rect 111 1037 115 1041
rect 423 1041 427 1045
rect 551 1041 555 1045
rect 679 1041 683 1045
rect 1975 1048 1979 1052
rect 2095 1048 2099 1052
rect 2215 1048 2219 1052
rect 2343 1048 2347 1052
rect 2487 1048 2491 1052
rect 2647 1048 2651 1052
rect 2823 1048 2827 1052
rect 2999 1048 3003 1052
rect 3159 1048 3163 1052
rect 463 1035 467 1039
rect 535 1035 539 1039
rect 583 1035 587 1039
rect 703 1039 707 1043
rect 799 1041 803 1045
rect 919 1041 923 1045
rect 1031 1041 1035 1045
rect 1143 1041 1147 1045
rect 1263 1041 1267 1045
rect 783 1035 787 1039
rect 907 1035 911 1039
rect 1039 1035 1040 1039
rect 1040 1035 1043 1039
rect 1135 1035 1139 1039
rect 1167 1035 1171 1039
rect 1255 1035 1259 1039
rect 1631 1037 1635 1041
rect 1671 1041 1675 1045
rect 3191 1041 3195 1045
rect 111 1019 115 1023
rect 1631 1019 1635 1023
rect 1671 1023 1675 1027
rect 1975 1019 1979 1023
rect 2095 1019 2099 1023
rect 2215 1019 2219 1023
rect 2343 1019 2347 1023
rect 2351 1023 2352 1027
rect 2352 1023 2355 1027
rect 2487 1019 2491 1023
rect 2647 1019 2651 1023
rect 2655 1019 2656 1023
rect 2656 1019 2659 1023
rect 2823 1019 2827 1023
rect 2831 1023 2832 1027
rect 2832 1023 2835 1027
rect 3007 1027 3011 1031
rect 2999 1019 3003 1023
rect 3159 1019 3163 1023
rect 3167 1023 3168 1027
rect 3168 1023 3171 1027
rect 3191 1023 3195 1027
rect 423 1012 427 1016
rect 551 1012 555 1016
rect 679 1012 683 1016
rect 799 1012 803 1016
rect 919 1012 923 1016
rect 1031 1012 1035 1016
rect 1143 1012 1147 1016
rect 1263 1012 1267 1016
rect 1927 1011 1931 1015
rect 1671 1001 1675 1005
rect 1895 1005 1899 1009
rect 2047 1005 2051 1009
rect 2079 1011 2083 1015
rect 1927 999 1931 1003
rect 2199 1005 2203 1009
rect 2231 1011 2235 1015
rect 2343 1005 2347 1009
rect 2351 1003 2352 1007
rect 2352 1003 2355 1007
rect 2495 1005 2499 1009
rect 2647 1005 2651 1009
rect 2655 999 2656 1003
rect 2656 999 2659 1003
rect 2703 999 2707 1003
rect 3191 1001 3195 1005
rect 327 988 331 992
rect 455 988 459 992
rect 575 988 579 992
rect 695 988 699 992
rect 815 988 819 992
rect 927 988 931 992
rect 1039 988 1043 992
rect 1159 988 1163 992
rect 111 981 115 985
rect 1631 981 1635 985
rect 1671 983 1675 987
rect 3191 983 3195 987
rect 1895 976 1899 980
rect 2047 976 2051 980
rect 2199 976 2203 980
rect 2343 976 2347 980
rect 2495 976 2499 980
rect 2647 976 2651 980
rect 111 963 115 967
rect 327 959 331 963
rect 335 959 336 963
rect 336 959 339 963
rect 455 959 459 963
rect 463 959 464 963
rect 464 959 467 963
rect 575 959 579 963
rect 583 963 584 967
rect 584 963 587 967
rect 695 959 699 963
rect 703 963 704 967
rect 704 963 707 967
rect 815 959 819 963
rect 824 959 828 963
rect 927 959 931 963
rect 951 959 955 963
rect 1039 959 1043 963
rect 1071 959 1075 963
rect 1159 959 1163 963
rect 1167 959 1168 963
rect 1168 959 1171 963
rect 1631 963 1635 967
rect 1791 964 1795 968
rect 1919 964 1923 968
rect 2071 964 2075 968
rect 2255 964 2259 968
rect 2463 964 2467 968
rect 2695 964 2699 968
rect 2935 964 2939 968
rect 3159 964 3163 968
rect 1671 957 1675 961
rect 3191 957 3195 961
rect 111 933 115 937
rect 223 937 227 941
rect 259 935 263 939
rect 335 935 339 939
rect 351 937 355 941
rect 471 937 475 941
rect 591 937 595 941
rect 711 937 715 941
rect 823 937 827 941
rect 943 937 947 941
rect 1063 937 1067 941
rect 1671 939 1675 943
rect 2231 943 2235 947
rect 463 931 467 935
rect 583 931 587 935
rect 703 931 707 935
rect 831 931 832 935
rect 832 931 835 935
rect 951 931 952 935
rect 952 931 955 935
rect 1071 931 1072 935
rect 1072 931 1075 935
rect 1631 933 1635 937
rect 1791 935 1795 939
rect 1803 935 1804 939
rect 1804 935 1807 939
rect 1919 935 1923 939
rect 1927 935 1928 939
rect 1928 935 1931 939
rect 2071 935 2075 939
rect 2079 935 2080 939
rect 2080 935 2083 939
rect 2255 935 2259 939
rect 2463 935 2467 939
rect 2471 935 2472 939
rect 2472 935 2475 939
rect 2695 935 2699 939
rect 2703 939 2704 943
rect 2704 939 2707 943
rect 2831 939 2835 943
rect 2935 935 2939 939
rect 2943 939 2944 943
rect 2944 939 2947 943
rect 3007 939 3011 943
rect 3159 935 3163 939
rect 3167 939 3168 943
rect 3168 939 3171 943
rect 3191 939 3195 943
rect 111 915 115 919
rect 1631 915 1635 919
rect 1671 913 1675 917
rect 1719 917 1723 921
rect 1871 917 1875 921
rect 2039 917 2043 921
rect 2223 917 2227 921
rect 223 908 227 912
rect 351 908 355 912
rect 471 908 475 912
rect 591 908 595 912
rect 711 908 715 912
rect 823 908 827 912
rect 943 908 947 912
rect 1063 908 1067 912
rect 1803 911 1807 915
rect 1927 911 1931 915
rect 2023 911 2027 915
rect 2079 911 2083 915
rect 2231 915 2232 919
rect 2232 915 2235 919
rect 2439 917 2443 921
rect 2447 915 2448 919
rect 2448 915 2451 919
rect 2471 915 2475 919
rect 2671 917 2675 921
rect 2703 915 2707 919
rect 2911 917 2915 921
rect 2943 915 2947 919
rect 3159 917 3163 921
rect 3167 915 3168 919
rect 3168 915 3171 919
rect 3191 913 3195 917
rect 1671 895 1675 899
rect 3191 895 3195 899
rect 135 884 139 888
rect 247 884 251 888
rect 383 884 387 888
rect 535 884 539 888
rect 711 884 715 888
rect 919 884 923 888
rect 1143 884 1147 888
rect 1383 884 1387 888
rect 1599 884 1603 888
rect 1719 888 1723 892
rect 1871 888 1875 892
rect 2039 888 2043 892
rect 2223 888 2227 892
rect 2439 888 2443 892
rect 2671 888 2675 892
rect 2911 888 2915 892
rect 3159 888 3163 892
rect 111 877 115 881
rect 1631 877 1635 881
rect 1695 876 1699 880
rect 2015 876 2019 880
rect 2367 876 2371 880
rect 2727 876 2731 880
rect 3087 876 3091 880
rect 1671 869 1675 873
rect 3191 869 3195 873
rect 111 859 115 863
rect 135 855 139 859
rect 247 855 251 859
rect 259 859 260 863
rect 260 859 263 863
rect 383 855 387 859
rect 535 855 539 859
rect 711 855 715 859
rect 719 855 720 859
rect 720 855 723 859
rect 919 855 923 859
rect 927 855 928 859
rect 928 855 931 859
rect 1143 855 1147 859
rect 1155 855 1156 859
rect 1156 855 1159 859
rect 1167 855 1171 859
rect 1383 855 1387 859
rect 1395 855 1396 859
rect 1396 855 1399 859
rect 1599 855 1603 859
rect 1631 859 1635 863
rect 111 837 115 841
rect 135 841 139 845
rect 259 847 263 851
rect 303 841 307 845
rect 503 841 507 845
rect 583 847 587 851
rect 695 841 699 845
rect 879 841 883 845
rect 1047 841 1051 845
rect 1199 841 1203 845
rect 1335 841 1339 845
rect 1471 841 1475 845
rect 1599 841 1603 845
rect 1671 851 1675 855
rect 1695 847 1699 851
rect 2015 847 2019 851
rect 2023 851 2024 855
rect 2024 851 2027 855
rect 2367 847 2371 851
rect 2447 851 2451 855
rect 2727 847 2731 851
rect 2739 847 2740 851
rect 2740 847 2743 851
rect 3087 847 3091 851
rect 3119 851 3123 855
rect 3167 851 3171 855
rect 3191 851 3195 855
rect 687 835 691 839
rect 719 835 723 839
rect 887 835 888 839
rect 888 835 891 839
rect 927 835 931 839
rect 1071 835 1075 839
rect 1155 835 1159 839
rect 1395 835 1399 839
rect 1527 835 1531 839
rect 1631 837 1635 841
rect 111 819 115 823
rect 1631 819 1635 823
rect 1671 821 1675 825
rect 2279 825 2283 829
rect 2439 825 2443 829
rect 2231 819 2235 823
rect 2307 819 2311 823
rect 2447 823 2448 827
rect 2448 823 2451 827
rect 2459 823 2463 827
rect 2583 825 2587 829
rect 2719 825 2723 829
rect 2623 819 2627 823
rect 2847 825 2851 829
rect 2975 825 2979 829
rect 3111 825 3115 829
rect 2739 819 2743 823
rect 2799 819 2803 823
rect 2931 819 2935 823
rect 3055 819 3059 823
rect 3119 823 3120 827
rect 3120 823 3123 827
rect 3191 821 3195 825
rect 135 812 139 816
rect 303 812 307 816
rect 503 812 507 816
rect 695 812 699 816
rect 879 812 883 816
rect 1047 812 1051 816
rect 1199 812 1203 816
rect 1335 812 1339 816
rect 1471 812 1475 816
rect 1599 812 1603 816
rect 1671 803 1675 807
rect 3191 803 3195 807
rect 2279 796 2283 800
rect 2439 796 2443 800
rect 2583 796 2587 800
rect 2719 796 2723 800
rect 2847 796 2851 800
rect 2975 796 2979 800
rect 3111 796 3115 800
rect 679 784 683 788
rect 807 784 811 788
rect 927 784 931 788
rect 1047 784 1051 788
rect 1167 784 1171 788
rect 1279 784 1283 788
rect 1399 784 1403 788
rect 1519 784 1523 788
rect 111 777 115 781
rect 1631 777 1635 781
rect 2199 780 2203 784
rect 2359 780 2363 784
rect 2511 780 2515 784
rect 2655 780 2659 784
rect 2791 780 2795 784
rect 2919 780 2923 784
rect 3047 780 3051 784
rect 3159 780 3163 784
rect 1671 773 1675 777
rect 3191 773 3195 777
rect 111 759 115 763
rect 679 755 683 759
rect 687 755 688 759
rect 688 755 691 759
rect 807 755 811 759
rect 815 755 816 759
rect 816 755 819 759
rect 927 755 931 759
rect 935 755 936 759
rect 936 755 939 759
rect 1047 755 1051 759
rect 1059 755 1060 759
rect 1060 755 1063 759
rect 1167 755 1171 759
rect 1191 755 1195 759
rect 1279 755 1283 759
rect 1303 755 1307 759
rect 1399 755 1403 759
rect 1423 763 1427 767
rect 1519 755 1523 759
rect 1527 759 1528 763
rect 1528 759 1531 763
rect 1631 759 1635 763
rect 1671 755 1675 759
rect 615 747 619 751
rect 2199 751 2203 755
rect 2359 751 2363 755
rect 2459 755 2463 759
rect 2511 751 2515 755
rect 2623 755 2627 759
rect 2655 751 2659 755
rect 2767 751 2771 755
rect 2791 751 2795 755
rect 2799 751 2800 755
rect 2800 751 2803 755
rect 2919 751 2923 755
rect 2931 755 2932 759
rect 2932 755 2935 759
rect 3047 751 3051 755
rect 3055 755 3056 759
rect 3056 755 3059 759
rect 3159 751 3163 755
rect 3167 751 3168 755
rect 3168 751 3171 755
rect 3191 755 3195 759
rect 2159 743 2163 747
rect 111 733 115 737
rect 575 737 579 741
rect 703 737 707 741
rect 831 737 835 741
rect 951 737 955 741
rect 1071 737 1075 741
rect 1183 737 1187 741
rect 1295 737 1299 741
rect 1415 737 1419 741
rect 583 731 584 735
rect 584 731 587 735
rect 615 731 619 735
rect 815 731 819 735
rect 855 731 859 735
rect 887 731 891 735
rect 935 731 939 735
rect 1059 731 1063 735
rect 1191 731 1192 735
rect 1192 731 1195 735
rect 1303 731 1304 735
rect 1304 731 1307 735
rect 1319 731 1323 735
rect 1423 735 1424 739
rect 1424 735 1427 739
rect 1631 733 1635 737
rect 1671 733 1675 737
rect 2127 737 2131 741
rect 2287 737 2291 741
rect 2447 737 2451 741
rect 2599 737 2603 741
rect 2759 737 2763 741
rect 2919 737 2923 741
rect 2159 731 2163 735
rect 2307 731 2311 735
rect 2459 731 2460 735
rect 2460 731 2463 735
rect 2623 731 2627 735
rect 2767 731 2768 735
rect 2768 731 2771 735
rect 2799 731 2803 735
rect 2931 735 2932 739
rect 2932 735 2935 739
rect 3191 733 3195 737
rect 111 715 115 719
rect 1631 715 1635 719
rect 1671 715 1675 719
rect 3191 715 3195 719
rect 575 708 579 712
rect 703 708 707 712
rect 831 708 835 712
rect 951 708 955 712
rect 1071 708 1075 712
rect 1183 708 1187 712
rect 1295 708 1299 712
rect 1415 708 1419 712
rect 2127 708 2131 712
rect 2287 708 2291 712
rect 2447 708 2451 712
rect 2599 708 2603 712
rect 2759 708 2763 712
rect 2919 708 2923 712
rect 2023 696 2027 700
rect 2151 696 2155 700
rect 2295 696 2299 700
rect 2447 696 2451 700
rect 2615 696 2619 700
rect 2799 696 2803 700
rect 2991 696 2995 700
rect 3159 696 3163 700
rect 1671 689 1675 693
rect 479 684 483 688
rect 607 684 611 688
rect 727 684 731 688
rect 847 684 851 688
rect 967 684 971 688
rect 1079 684 1083 688
rect 1191 684 1195 688
rect 3191 689 3195 693
rect 1311 684 1315 688
rect 111 677 115 681
rect 1631 677 1635 681
rect 1671 671 1675 675
rect 2931 675 2935 679
rect 2023 667 2027 671
rect 2031 667 2032 671
rect 2032 667 2035 671
rect 2151 667 2155 671
rect 2159 667 2160 671
rect 2160 667 2163 671
rect 2295 667 2299 671
rect 2307 667 2308 671
rect 2308 667 2311 671
rect 2447 667 2451 671
rect 2459 667 2460 671
rect 2460 667 2463 671
rect 2615 667 2619 671
rect 2623 667 2624 671
rect 2624 667 2627 671
rect 2799 667 2803 671
rect 2807 667 2808 671
rect 2808 667 2811 671
rect 2871 667 2875 671
rect 2991 667 2995 671
rect 3159 667 3163 671
rect 3167 671 3168 675
rect 3168 671 3171 675
rect 3191 671 3195 675
rect 111 659 115 663
rect 479 655 483 659
rect 487 655 488 659
rect 488 655 491 659
rect 607 655 611 659
rect 615 655 616 659
rect 616 655 619 659
rect 631 655 635 659
rect 727 655 731 659
rect 751 655 755 659
rect 847 655 851 659
rect 855 655 856 659
rect 856 655 859 659
rect 967 655 971 659
rect 999 655 1003 659
rect 1079 655 1083 659
rect 1103 655 1107 659
rect 1191 655 1195 659
rect 1223 659 1227 663
rect 1311 655 1315 659
rect 1319 659 1320 663
rect 1320 659 1323 663
rect 1631 659 1635 663
rect 1671 645 1675 649
rect 1919 649 1923 653
rect 2047 649 2051 653
rect 2183 649 2187 653
rect 2327 649 2331 653
rect 2471 649 2475 653
rect 2615 649 2619 653
rect 2759 649 2763 653
rect 1895 643 1899 647
rect 2031 643 2035 647
rect 2159 643 2163 647
rect 2191 643 2192 647
rect 2192 643 2195 647
rect 2307 643 2311 647
rect 2459 643 2463 647
rect 2623 643 2624 647
rect 2624 643 2627 647
rect 2767 647 2768 651
rect 2768 647 2771 651
rect 2807 647 2811 651
rect 3191 645 3195 649
rect 111 629 115 633
rect 375 633 379 637
rect 503 633 507 637
rect 623 633 627 637
rect 743 633 747 637
rect 407 627 411 631
rect 487 627 491 631
rect 631 627 632 631
rect 632 627 635 631
rect 671 627 675 631
rect 751 631 752 635
rect 752 631 755 635
rect 775 631 779 635
rect 863 633 867 637
rect 975 633 979 637
rect 1095 633 1099 637
rect 1215 633 1219 637
rect 855 627 859 631
rect 999 627 1003 631
rect 1103 627 1104 631
rect 1104 627 1107 631
rect 1223 631 1224 635
rect 1224 631 1227 635
rect 1631 629 1635 633
rect 1671 627 1675 631
rect 3191 627 3195 631
rect 1919 620 1923 624
rect 2047 620 2051 624
rect 2183 620 2187 624
rect 2327 620 2331 624
rect 2471 620 2475 624
rect 2615 620 2619 624
rect 2759 620 2763 624
rect 111 611 115 615
rect 1631 611 1635 615
rect 375 604 379 608
rect 503 604 507 608
rect 623 604 627 608
rect 743 604 747 608
rect 863 604 867 608
rect 975 604 979 608
rect 1095 604 1099 608
rect 1215 604 1219 608
rect 1847 604 1851 608
rect 2015 604 2019 608
rect 2183 604 2187 608
rect 2359 604 2363 608
rect 2551 604 2555 608
rect 2751 604 2755 608
rect 2959 604 2963 608
rect 3159 604 3163 608
rect 1671 597 1675 601
rect 3191 597 3195 601
rect 271 584 275 588
rect 399 584 403 588
rect 527 584 531 588
rect 647 584 651 588
rect 767 584 771 588
rect 879 584 883 588
rect 991 584 995 588
rect 1111 584 1115 588
rect 111 577 115 581
rect 1631 577 1635 581
rect 1671 579 1675 583
rect 1847 575 1851 579
rect 2015 575 2019 579
rect 2183 575 2187 579
rect 2191 579 2192 583
rect 2192 579 2195 583
rect 111 559 115 563
rect 271 555 275 559
rect 311 555 315 559
rect 399 555 403 559
rect 407 555 408 559
rect 408 555 411 559
rect 431 555 435 559
rect 527 555 531 559
rect 551 555 555 559
rect 647 555 651 559
rect 671 555 675 559
rect 767 555 771 559
rect 776 559 780 563
rect 879 555 883 559
rect 887 555 888 559
rect 888 555 891 559
rect 991 555 995 559
rect 999 555 1000 559
rect 1000 555 1003 559
rect 1111 555 1115 559
rect 1143 555 1147 559
rect 1631 559 1635 563
rect 1671 561 1675 565
rect 1767 565 1771 569
rect 1895 563 1899 567
rect 1927 565 1931 569
rect 2087 565 2091 569
rect 2247 565 2251 569
rect 2359 575 2363 579
rect 2415 575 2419 579
rect 2551 575 2555 579
rect 2031 559 2035 563
rect 2111 559 2115 563
rect 2407 565 2411 569
rect 2415 563 2416 567
rect 2416 563 2419 567
rect 2459 563 2463 567
rect 2567 565 2571 569
rect 2751 575 2755 579
rect 2760 579 2764 583
rect 2959 575 2963 579
rect 3159 575 3163 579
rect 3167 579 3168 583
rect 3168 579 3171 583
rect 3191 579 3195 583
rect 2607 559 2611 563
rect 3191 561 3195 565
rect 311 547 315 551
rect 431 547 435 551
rect 1671 543 1675 547
rect 3191 543 3195 547
rect 111 529 115 533
rect 175 533 179 537
rect 303 533 307 537
rect 423 533 427 537
rect 147 527 151 531
rect 311 527 312 531
rect 312 527 315 531
rect 431 531 432 535
rect 432 531 435 535
rect 543 533 547 537
rect 663 533 667 537
rect 775 533 779 537
rect 551 527 552 531
rect 552 527 555 531
rect 671 527 672 531
rect 672 527 675 531
rect 783 531 784 535
rect 784 531 787 535
rect 887 533 891 537
rect 1007 533 1011 537
rect 1767 536 1771 540
rect 1927 536 1931 540
rect 2087 536 2091 540
rect 2247 536 2251 540
rect 2407 536 2411 540
rect 2567 536 2571 540
rect 827 527 831 531
rect 895 527 896 531
rect 896 527 899 531
rect 999 527 1003 531
rect 1631 529 1635 533
rect 1695 524 1699 528
rect 1887 524 1891 528
rect 2103 524 2107 528
rect 2343 524 2347 528
rect 2599 524 2603 528
rect 2863 524 2867 528
rect 3135 524 3139 528
rect 1671 517 1675 521
rect 3191 517 3195 521
rect 111 511 115 515
rect 1631 511 1635 515
rect 175 504 179 508
rect 303 504 307 508
rect 423 504 427 508
rect 543 504 547 508
rect 663 504 667 508
rect 775 504 779 508
rect 887 504 891 508
rect 1007 504 1011 508
rect 1671 499 1675 503
rect 1695 495 1699 499
rect 1703 495 1704 499
rect 1704 495 1707 499
rect 1887 495 1891 499
rect 1895 499 1896 503
rect 1896 499 1899 503
rect 2103 495 2107 499
rect 2111 499 2112 503
rect 2112 499 2115 503
rect 2343 495 2347 499
rect 2415 499 2419 503
rect 2599 495 2603 499
rect 2607 495 2608 499
rect 2608 495 2611 499
rect 2631 495 2635 499
rect 2863 495 2867 499
rect 2871 495 2872 499
rect 2872 495 2875 499
rect 2927 495 2931 499
rect 3135 495 3139 499
rect 3143 499 3144 503
rect 3144 499 3147 503
rect 3167 499 3171 503
rect 3191 499 3195 503
rect 135 480 139 484
rect 231 480 235 484
rect 359 480 363 484
rect 503 480 507 484
rect 655 480 659 484
rect 815 480 819 484
rect 975 480 979 484
rect 1135 480 1139 484
rect 1295 480 1299 484
rect 1455 480 1459 484
rect 1599 480 1603 484
rect 111 473 115 477
rect 1631 473 1635 477
rect 1671 473 1675 477
rect 1695 477 1699 481
rect 1703 475 1704 479
rect 1704 475 1707 479
rect 2023 477 2027 481
rect 2031 475 2032 479
rect 2032 475 2035 479
rect 2059 475 2063 479
rect 2383 477 2387 481
rect 2415 475 2419 479
rect 2743 477 2747 481
rect 3111 477 3115 481
rect 2751 471 2752 475
rect 2752 471 2755 475
rect 3119 475 3120 479
rect 3120 475 3123 479
rect 3143 475 3147 479
rect 3191 473 3195 477
rect 111 455 115 459
rect 135 451 139 455
rect 147 455 148 459
rect 148 455 151 459
rect 231 451 235 455
rect 359 451 363 455
rect 471 459 475 463
rect 1607 463 1611 467
rect 1703 463 1707 467
rect 503 451 507 455
rect 655 451 659 455
rect 663 453 664 455
rect 664 453 667 455
rect 663 451 667 453
rect 815 451 819 455
rect 827 451 828 455
rect 828 451 831 455
rect 975 451 979 455
rect 983 451 984 455
rect 984 451 987 455
rect 1135 451 1139 455
rect 1143 455 1144 459
rect 1144 455 1147 459
rect 1295 451 1299 455
rect 1343 451 1347 455
rect 1455 451 1459 455
rect 1467 451 1468 455
rect 1468 451 1471 455
rect 1599 451 1603 455
rect 1607 451 1608 455
rect 1608 451 1611 455
rect 1631 455 1635 459
rect 1671 455 1675 459
rect 3191 455 3195 459
rect 1695 448 1699 452
rect 2023 448 2027 452
rect 2383 448 2387 452
rect 2743 448 2747 452
rect 3111 448 3115 452
rect 1143 435 1147 439
rect 1231 435 1235 439
rect 1467 435 1471 439
rect 1607 435 1611 439
rect 111 425 115 429
rect 727 429 731 433
rect 855 429 859 433
rect 983 429 987 433
rect 1103 429 1107 433
rect 815 423 819 427
rect 827 423 831 427
rect 991 423 992 427
rect 992 423 995 427
rect 1143 427 1147 431
rect 1223 429 1227 433
rect 1231 427 1232 431
rect 1232 427 1235 431
rect 1335 429 1339 433
rect 1447 429 1451 433
rect 1343 423 1344 427
rect 1344 423 1347 427
rect 1467 427 1471 431
rect 1567 429 1571 433
rect 2247 432 2251 436
rect 2375 432 2379 436
rect 2503 432 2507 436
rect 2623 432 2627 436
rect 2743 432 2747 436
rect 2855 432 2859 436
rect 2967 432 2971 436
rect 3087 432 3091 436
rect 1607 427 1611 431
rect 1631 425 1635 429
rect 1671 425 1675 429
rect 3191 425 3195 429
rect 111 407 115 411
rect 1631 407 1635 411
rect 1671 407 1675 411
rect 727 400 731 404
rect 855 400 859 404
rect 983 400 987 404
rect 1103 400 1107 404
rect 1223 400 1227 404
rect 1335 400 1339 404
rect 1447 400 1451 404
rect 1567 400 1571 404
rect 2247 403 2251 407
rect 2259 403 2260 407
rect 2260 403 2263 407
rect 2375 403 2379 407
rect 2387 403 2388 407
rect 2388 403 2391 407
rect 2503 403 2507 407
rect 2515 403 2516 407
rect 2516 403 2519 407
rect 2623 403 2627 407
rect 2631 403 2632 407
rect 2632 403 2635 407
rect 2671 403 2675 407
rect 2743 403 2747 407
rect 2751 403 2752 407
rect 2752 403 2755 407
rect 2799 403 2803 407
rect 2855 403 2859 407
rect 2863 407 2864 411
rect 2864 407 2867 411
rect 2927 407 2931 411
rect 2967 403 2971 407
rect 2975 403 2976 407
rect 2976 403 2979 407
rect 3035 403 3039 407
rect 3087 403 3091 407
rect 3119 407 3123 411
rect 3191 407 3195 411
rect 647 380 651 384
rect 807 380 811 384
rect 951 380 955 384
rect 1087 380 1091 384
rect 1215 380 1219 384
rect 1335 380 1339 384
rect 1463 380 1467 384
rect 111 373 115 377
rect 1631 373 1635 377
rect 1671 377 1675 381
rect 2151 381 2155 385
rect 2279 381 2283 385
rect 2407 381 2411 385
rect 2535 381 2539 385
rect 2663 381 2667 385
rect 2259 375 2263 379
rect 2387 375 2391 379
rect 2515 375 2519 379
rect 2575 375 2579 379
rect 2671 379 2672 383
rect 2672 379 2675 383
rect 2751 379 2755 383
rect 2791 381 2795 385
rect 2799 379 2800 383
rect 2800 379 2803 383
rect 2863 379 2867 383
rect 2919 381 2923 385
rect 2927 379 2928 383
rect 2928 379 2931 383
rect 2975 379 2979 383
rect 3047 381 3051 385
rect 3159 381 3163 385
rect 3035 375 3039 379
rect 3119 375 3123 379
rect 3167 375 3168 379
rect 3168 375 3171 379
rect 3191 377 3195 381
rect 111 355 115 359
rect 647 351 651 355
rect 655 355 656 359
rect 656 355 659 359
rect 807 351 811 355
rect 815 351 816 355
rect 816 351 819 355
rect 951 351 955 355
rect 991 351 995 355
rect 1087 351 1091 355
rect 111 333 115 337
rect 543 337 547 341
rect 671 337 675 341
rect 807 337 811 341
rect 943 337 947 341
rect 631 331 635 335
rect 655 331 659 335
rect 815 331 816 335
rect 816 331 819 335
rect 1079 337 1083 341
rect 1215 351 1219 355
rect 1335 351 1339 355
rect 1343 351 1344 355
rect 1344 351 1347 355
rect 1223 337 1227 341
rect 1295 335 1299 339
rect 1343 335 1347 339
rect 1367 337 1371 341
rect 1463 351 1467 355
rect 1471 355 1472 359
rect 1472 355 1475 359
rect 1631 355 1635 359
rect 1671 359 1675 363
rect 3191 359 3195 363
rect 2151 352 2155 356
rect 2279 352 2283 356
rect 2407 352 2411 356
rect 2535 352 2539 356
rect 2663 352 2667 356
rect 2791 352 2795 356
rect 2919 352 2923 356
rect 3047 352 3051 356
rect 3159 352 3163 356
rect 1471 335 1475 339
rect 1631 333 1635 337
rect 2047 328 2051 332
rect 2175 328 2179 332
rect 2303 328 2307 332
rect 2431 328 2435 332
rect 2567 328 2571 332
rect 2711 328 2715 332
rect 2863 328 2867 332
rect 3023 328 3027 332
rect 3159 328 3163 332
rect 1671 321 1675 325
rect 3191 321 3195 325
rect 111 315 115 319
rect 1631 315 1635 319
rect 543 308 547 312
rect 671 308 675 312
rect 807 308 811 312
rect 943 308 947 312
rect 1079 308 1083 312
rect 1223 308 1227 312
rect 1367 308 1371 312
rect 1671 303 1675 307
rect 2047 299 2051 303
rect 2059 299 2060 303
rect 2060 299 2063 303
rect 2175 299 2179 303
rect 2187 299 2188 303
rect 2188 299 2191 303
rect 2303 299 2307 303
rect 2327 299 2331 303
rect 2431 299 2435 303
rect 2440 303 2444 307
rect 2567 299 2571 303
rect 2575 299 2576 303
rect 2576 299 2579 303
rect 2671 299 2675 303
rect 2711 299 2715 303
rect 2719 299 2720 303
rect 2720 299 2723 303
rect 2791 299 2795 303
rect 2863 299 2867 303
rect 2871 303 2872 307
rect 2872 303 2875 307
rect 2927 303 2931 307
rect 3023 299 3027 303
rect 3035 303 3036 307
rect 3036 303 3039 307
rect 3159 299 3163 303
rect 3167 303 3168 307
rect 3168 303 3171 307
rect 3191 303 3195 307
rect 463 292 467 296
rect 623 292 627 296
rect 767 292 771 296
rect 903 292 907 296
rect 1031 292 1035 296
rect 1159 292 1163 296
rect 1287 292 1291 296
rect 111 285 115 289
rect 1631 285 1635 289
rect 1671 277 1675 281
rect 1943 281 1947 285
rect 2071 281 2075 285
rect 2199 281 2203 285
rect 2319 281 2323 285
rect 2439 281 2443 285
rect 2551 281 2555 285
rect 2059 275 2063 279
rect 2187 275 2191 279
rect 2327 275 2328 279
rect 2328 275 2331 279
rect 2447 275 2448 279
rect 2448 275 2451 279
rect 2527 275 2531 279
rect 2575 279 2579 283
rect 2663 281 2667 285
rect 2671 279 2672 283
rect 2672 279 2675 283
rect 2719 279 2723 283
rect 2783 281 2787 285
rect 2791 279 2792 283
rect 2792 279 2795 283
rect 2871 279 2875 283
rect 3191 277 3195 281
rect 111 267 115 271
rect 463 263 467 267
rect 471 267 472 271
rect 472 267 475 271
rect 623 263 627 267
rect 631 263 632 267
rect 632 263 635 267
rect 767 263 771 267
rect 775 267 776 271
rect 776 267 779 271
rect 815 267 819 271
rect 903 263 907 267
rect 1031 263 1035 267
rect 1159 263 1163 267
rect 111 245 115 249
rect 359 249 363 253
rect 367 247 368 251
rect 368 247 371 251
rect 471 247 475 251
rect 487 249 491 253
rect 623 249 627 253
rect 759 249 763 253
rect 631 243 632 247
rect 632 243 635 247
rect 895 249 899 253
rect 1039 249 1043 253
rect 1183 249 1187 253
rect 1287 263 1291 267
rect 1295 267 1296 271
rect 1296 267 1299 271
rect 1631 267 1635 271
rect 1671 259 1675 263
rect 3191 259 3195 263
rect 1943 252 1947 256
rect 767 239 771 243
rect 903 243 907 247
rect 2071 252 2075 256
rect 2199 252 2203 256
rect 2319 252 2323 256
rect 2439 252 2443 256
rect 2551 252 2555 256
rect 2663 252 2667 256
rect 2783 252 2787 256
rect 1295 247 1299 251
rect 1631 245 1635 249
rect 111 227 115 231
rect 1631 227 1635 231
rect 1847 228 1851 232
rect 1975 228 1979 232
rect 2103 228 2107 232
rect 2247 228 2251 232
rect 2407 228 2411 232
rect 2583 228 2587 232
rect 2767 228 2771 232
rect 2967 228 2971 232
rect 3159 228 3163 232
rect 359 220 363 224
rect 487 220 491 224
rect 623 220 627 224
rect 759 220 763 224
rect 895 220 899 224
rect 1039 220 1043 224
rect 1183 220 1187 224
rect 1671 221 1675 225
rect 3191 221 3195 225
rect 279 204 283 208
rect 447 204 451 208
rect 615 204 619 208
rect 775 204 779 208
rect 943 204 947 208
rect 1111 204 1115 208
rect 1671 203 1675 207
rect 111 197 115 201
rect 1631 197 1635 201
rect 1847 199 1851 203
rect 1855 199 1856 203
rect 1856 199 1859 203
rect 1975 199 1979 203
rect 1983 199 1984 203
rect 1984 199 1987 203
rect 2103 199 2107 203
rect 2111 199 2112 203
rect 2112 199 2115 203
rect 2247 199 2251 203
rect 2255 199 2256 203
rect 2256 199 2259 203
rect 2319 199 2323 203
rect 2407 199 2411 203
rect 2415 199 2416 203
rect 2416 199 2419 203
rect 2503 199 2507 203
rect 2583 199 2587 203
rect 2591 199 2592 203
rect 2592 199 2595 203
rect 2767 199 2771 203
rect 2791 203 2795 207
rect 2927 207 2931 211
rect 2967 199 2971 203
rect 3159 199 3163 203
rect 3167 203 3168 207
rect 3168 203 3171 207
rect 3191 203 3195 207
rect 111 179 115 183
rect 279 175 283 179
rect 367 179 371 183
rect 111 161 115 165
rect 199 165 203 169
rect 147 159 151 163
rect 367 165 371 169
rect 447 175 451 179
rect 471 179 475 183
rect 903 183 907 187
rect 615 175 619 179
rect 624 175 628 179
rect 775 175 779 179
rect 943 175 947 179
rect 1111 175 1115 179
rect 1631 179 1635 183
rect 535 165 539 169
rect 695 165 699 169
rect 471 159 475 163
rect 547 159 548 163
rect 548 159 551 163
rect 703 159 704 163
rect 704 159 707 163
rect 767 159 771 163
rect 863 165 867 169
rect 1031 165 1035 169
rect 903 159 907 163
rect 1023 159 1027 163
rect 1671 173 1675 177
rect 1743 177 1747 181
rect 1871 177 1875 181
rect 1999 177 2003 181
rect 2143 177 2147 181
rect 1751 171 1752 175
rect 1752 171 1755 175
rect 1855 171 1859 175
rect 1983 171 1987 175
rect 2111 171 2115 175
rect 2255 175 2259 179
rect 2311 177 2315 181
rect 2319 175 2320 179
rect 2320 175 2323 179
rect 2359 175 2363 179
rect 2415 175 2419 179
rect 2495 177 2499 181
rect 2503 175 2504 179
rect 2504 175 2507 179
rect 2591 175 2595 179
rect 2703 177 2707 181
rect 2715 177 2719 179
rect 2715 175 2716 177
rect 2716 175 2719 177
rect 2919 177 2923 181
rect 2927 175 2928 179
rect 2928 175 2931 179
rect 3135 177 3139 181
rect 3143 175 3144 179
rect 3144 175 3147 179
rect 3167 175 3171 179
rect 3191 173 3195 177
rect 1631 161 1635 165
rect 1671 155 1675 159
rect 3191 155 3195 159
rect 1743 148 1747 152
rect 111 143 115 147
rect 1871 148 1875 152
rect 1999 148 2003 152
rect 2143 148 2147 152
rect 2311 148 2315 152
rect 2495 148 2499 152
rect 2703 148 2707 152
rect 2919 148 2923 152
rect 3135 148 3139 152
rect 1631 143 1635 147
rect 199 136 203 140
rect 367 136 371 140
rect 535 136 539 140
rect 695 136 699 140
rect 863 136 867 140
rect 1031 136 1035 140
rect 1695 120 1699 124
rect 1815 120 1819 124
rect 1943 120 1947 124
rect 2071 120 2075 124
rect 2199 120 2203 124
rect 2351 120 2355 124
rect 2519 120 2523 124
rect 2711 120 2715 124
rect 2911 120 2915 124
rect 3111 120 3115 124
rect 135 112 139 116
rect 191 112 195 116
rect 287 112 291 116
rect 383 112 387 116
rect 479 112 483 116
rect 583 112 587 116
rect 695 112 699 116
rect 815 112 819 116
rect 943 112 947 116
rect 1079 112 1083 116
rect 1215 112 1219 116
rect 1351 112 1355 116
rect 1487 112 1491 116
rect 1599 112 1603 116
rect 1671 113 1675 117
rect 3191 113 3195 117
rect 111 105 115 109
rect 1631 105 1635 109
rect 111 87 115 91
rect 135 83 139 87
rect 147 87 148 91
rect 148 87 151 91
rect 191 83 195 87
rect 287 83 291 87
rect 383 83 387 87
rect 479 83 483 87
rect 547 91 551 95
rect 583 83 587 87
rect 695 83 699 87
rect 703 87 704 91
rect 704 87 707 91
rect 815 83 819 87
rect 943 83 947 87
rect 1023 91 1027 95
rect 1671 95 1675 99
rect 1079 83 1083 87
rect 1215 83 1219 87
rect 1351 83 1355 87
rect 1487 83 1491 87
rect 1599 83 1603 87
rect 1631 87 1635 91
rect 1695 91 1699 95
rect 1815 91 1819 95
rect 1943 91 1947 95
rect 2071 91 2075 95
rect 2199 91 2203 95
rect 2351 91 2355 95
rect 2359 95 2360 99
rect 2360 95 2363 99
rect 2519 91 2523 95
rect 2527 95 2528 99
rect 2528 95 2531 99
rect 2711 91 2715 95
rect 2719 95 2720 99
rect 2720 95 2723 99
rect 2911 91 2915 95
rect 2920 95 2924 99
rect 3111 91 3115 95
rect 3143 95 3147 99
rect 3191 95 3195 99
rect 1751 83 1755 87
<< m3 >>
rect 1671 3310 1675 3311
rect 1671 3305 1675 3306
rect 3055 3310 3059 3311
rect 3055 3305 3059 3306
rect 3191 3310 3195 3311
rect 3191 3305 3195 3306
rect 1672 3298 1674 3305
rect 3054 3304 3060 3305
rect 3054 3300 3055 3304
rect 3059 3300 3060 3304
rect 3054 3299 3060 3300
rect 3192 3298 3194 3305
rect 1670 3297 1676 3298
rect 1670 3293 1671 3297
rect 1675 3293 1676 3297
rect 1670 3292 1676 3293
rect 3190 3297 3196 3298
rect 3190 3293 3191 3297
rect 3195 3293 3196 3297
rect 3190 3292 3196 3293
rect 1670 3279 1676 3280
rect 1670 3275 1671 3279
rect 1675 3275 1676 3279
rect 3190 3279 3196 3280
rect 1670 3274 1676 3275
rect 3054 3275 3060 3276
rect 1672 3271 1674 3274
rect 3054 3271 3055 3275
rect 3059 3271 3060 3275
rect 1671 3270 1675 3271
rect 2151 3270 2155 3271
rect 2287 3270 2291 3271
rect 2423 3270 2427 3271
rect 2567 3270 2571 3271
rect 2711 3270 2715 3271
rect 2855 3270 2859 3271
rect 2999 3270 3003 3271
rect 3054 3270 3060 3271
rect 3118 3275 3124 3276
rect 3118 3271 3119 3275
rect 3123 3271 3124 3275
rect 3190 3275 3191 3279
rect 3195 3275 3196 3279
rect 3190 3274 3196 3275
rect 3192 3271 3194 3274
rect 3118 3270 3124 3271
rect 3191 3270 3195 3271
rect 1671 3265 1675 3266
rect 2150 3265 2156 3266
rect 1672 3262 1674 3265
rect 1670 3261 1676 3262
rect 1670 3257 1671 3261
rect 1675 3257 1676 3261
rect 2150 3261 2151 3265
rect 2155 3261 2156 3265
rect 2150 3260 2156 3261
rect 2286 3265 2292 3266
rect 2286 3261 2287 3265
rect 2291 3261 2292 3265
rect 2286 3260 2292 3261
rect 2422 3265 2428 3266
rect 2422 3261 2423 3265
rect 2427 3261 2428 3265
rect 2422 3260 2428 3261
rect 2566 3265 2572 3266
rect 2566 3261 2567 3265
rect 2571 3261 2572 3265
rect 2566 3260 2572 3261
rect 2710 3265 2716 3266
rect 2710 3261 2711 3265
rect 2715 3261 2716 3265
rect 2710 3260 2716 3261
rect 2854 3265 2860 3266
rect 2854 3261 2855 3265
rect 2859 3261 2860 3265
rect 2854 3260 2860 3261
rect 2998 3265 3004 3266
rect 3055 3265 3059 3266
rect 2998 3261 2999 3265
rect 3003 3261 3004 3265
rect 2998 3260 3004 3261
rect 1670 3256 1676 3257
rect 2182 3259 2188 3260
rect 2182 3255 2183 3259
rect 2187 3255 2188 3259
rect 2182 3254 2188 3255
rect 2554 3259 2560 3260
rect 2554 3255 2555 3259
rect 2559 3255 2560 3259
rect 2554 3254 2560 3255
rect 2734 3259 2740 3260
rect 2734 3255 2735 3259
rect 2739 3255 2740 3259
rect 2734 3254 2740 3255
rect 1670 3243 1676 3244
rect 1670 3239 1671 3243
rect 1675 3239 1676 3243
rect 1670 3238 1676 3239
rect 1672 3231 1674 3238
rect 2150 3236 2156 3237
rect 2150 3232 2151 3236
rect 2155 3232 2156 3236
rect 2150 3231 2156 3232
rect 1671 3230 1675 3231
rect 1671 3225 1675 3226
rect 1999 3230 2003 3231
rect 1999 3225 2003 3226
rect 2151 3230 2155 3231
rect 2151 3225 2155 3226
rect 2175 3230 2179 3231
rect 2175 3225 2179 3226
rect 1672 3218 1674 3225
rect 1998 3224 2004 3225
rect 1998 3220 1999 3224
rect 2003 3220 2004 3224
rect 1998 3219 2004 3220
rect 2174 3224 2180 3225
rect 2174 3220 2175 3224
rect 2179 3220 2180 3224
rect 2174 3219 2180 3220
rect 1670 3217 1676 3218
rect 1670 3213 1671 3217
rect 1675 3213 1676 3217
rect 1670 3212 1676 3213
rect 1670 3199 1676 3200
rect 1670 3195 1671 3199
rect 1675 3195 1676 3199
rect 2184 3196 2186 3254
rect 2286 3236 2292 3237
rect 2286 3232 2287 3236
rect 2291 3232 2292 3236
rect 2286 3231 2292 3232
rect 2422 3236 2428 3237
rect 2422 3232 2423 3236
rect 2427 3232 2428 3236
rect 2422 3231 2428 3232
rect 2287 3230 2291 3231
rect 2287 3225 2291 3226
rect 2359 3230 2363 3231
rect 2359 3225 2363 3226
rect 2423 3230 2427 3231
rect 2423 3225 2427 3226
rect 2543 3230 2547 3231
rect 2543 3225 2547 3226
rect 2358 3224 2364 3225
rect 2358 3220 2359 3224
rect 2363 3220 2364 3224
rect 2358 3219 2364 3220
rect 2542 3224 2548 3225
rect 2542 3220 2543 3224
rect 2547 3220 2548 3224
rect 2542 3219 2548 3220
rect 2556 3200 2558 3254
rect 2566 3236 2572 3237
rect 2566 3232 2567 3236
rect 2571 3232 2572 3236
rect 2566 3231 2572 3232
rect 2710 3236 2716 3237
rect 2710 3232 2711 3236
rect 2715 3232 2716 3236
rect 2710 3231 2716 3232
rect 2567 3230 2571 3231
rect 2567 3225 2571 3226
rect 2711 3230 2715 3231
rect 2711 3225 2715 3226
rect 2727 3230 2731 3231
rect 2727 3225 2731 3226
rect 2726 3224 2732 3225
rect 2726 3220 2727 3224
rect 2731 3220 2732 3224
rect 2726 3219 2732 3220
rect 2736 3200 2738 3254
rect 2854 3236 2860 3237
rect 2854 3232 2855 3236
rect 2859 3232 2860 3236
rect 2854 3231 2860 3232
rect 2998 3236 3004 3237
rect 2998 3232 2999 3236
rect 3003 3232 3004 3236
rect 2998 3231 3004 3232
rect 2855 3230 2859 3231
rect 2855 3225 2859 3226
rect 2919 3230 2923 3231
rect 2919 3225 2923 3226
rect 2999 3230 3003 3231
rect 2999 3225 3003 3226
rect 3111 3230 3115 3231
rect 3111 3225 3115 3226
rect 2918 3224 2924 3225
rect 2918 3220 2919 3224
rect 2923 3220 2924 3224
rect 2918 3219 2924 3220
rect 3110 3224 3116 3225
rect 3110 3220 3111 3224
rect 3115 3220 3116 3224
rect 3110 3219 3116 3220
rect 2554 3199 2560 3200
rect 1670 3194 1676 3195
rect 1998 3195 2004 3196
rect 1672 3191 1674 3194
rect 1998 3191 1999 3195
rect 2003 3191 2004 3195
rect 2046 3195 2052 3196
rect 2046 3191 2047 3195
rect 2051 3191 2052 3195
rect 1671 3190 1675 3191
rect 1847 3190 1851 3191
rect 1998 3190 2004 3191
rect 2039 3190 2043 3191
rect 2046 3190 2052 3191
rect 2174 3195 2180 3196
rect 2174 3191 2175 3195
rect 2179 3191 2180 3195
rect 2174 3190 2180 3191
rect 2182 3195 2188 3196
rect 2182 3191 2183 3195
rect 2187 3191 2188 3195
rect 2182 3190 2188 3191
rect 2234 3195 2240 3196
rect 2234 3191 2235 3195
rect 2239 3191 2240 3195
rect 2358 3195 2364 3196
rect 2358 3191 2359 3195
rect 2363 3191 2364 3195
rect 2542 3195 2548 3196
rect 2542 3191 2543 3195
rect 2547 3191 2548 3195
rect 2554 3195 2555 3199
rect 2559 3195 2560 3199
rect 2734 3199 2740 3200
rect 2554 3194 2560 3195
rect 2726 3195 2732 3196
rect 2234 3190 2240 3191
rect 2247 3190 2251 3191
rect 2358 3190 2364 3191
rect 2463 3190 2467 3191
rect 2542 3190 2548 3191
rect 1671 3185 1675 3186
rect 1846 3185 1852 3186
rect 1999 3185 2003 3186
rect 2038 3185 2044 3186
rect 1672 3182 1674 3185
rect 1670 3181 1676 3182
rect 1670 3177 1671 3181
rect 1675 3177 1676 3181
rect 1846 3181 1847 3185
rect 1851 3181 1852 3185
rect 1846 3180 1852 3181
rect 2038 3181 2039 3185
rect 2043 3181 2044 3185
rect 2048 3184 2050 3190
rect 2175 3185 2179 3186
rect 2184 3184 2186 3190
rect 2038 3180 2044 3181
rect 2046 3183 2052 3184
rect 1670 3176 1676 3177
rect 1854 3179 1860 3180
rect 1854 3175 1855 3179
rect 1859 3175 1860 3179
rect 2046 3179 2047 3183
rect 2051 3179 2052 3183
rect 2046 3178 2052 3179
rect 2182 3183 2188 3184
rect 2182 3179 2183 3183
rect 2187 3179 2188 3183
rect 2236 3180 2238 3190
rect 2246 3185 2252 3186
rect 2359 3185 2363 3186
rect 2462 3185 2468 3186
rect 2543 3185 2547 3186
rect 2246 3181 2247 3185
rect 2251 3181 2252 3185
rect 2246 3180 2252 3181
rect 2462 3181 2463 3185
rect 2467 3181 2468 3185
rect 2462 3180 2468 3181
rect 2556 3180 2558 3194
rect 2726 3191 2727 3195
rect 2731 3191 2732 3195
rect 2734 3195 2735 3199
rect 2739 3195 2740 3199
rect 3120 3196 3122 3270
rect 3191 3265 3195 3266
rect 3192 3262 3194 3265
rect 3190 3261 3196 3262
rect 3190 3257 3191 3261
rect 3195 3257 3196 3261
rect 3190 3256 3196 3257
rect 3190 3243 3196 3244
rect 3190 3239 3191 3243
rect 3195 3239 3196 3243
rect 3190 3238 3196 3239
rect 3192 3231 3194 3238
rect 3191 3230 3195 3231
rect 3191 3225 3195 3226
rect 3192 3218 3194 3225
rect 3190 3217 3196 3218
rect 3190 3213 3191 3217
rect 3195 3213 3196 3217
rect 3190 3212 3196 3213
rect 3190 3199 3196 3200
rect 2734 3194 2740 3195
rect 2918 3195 2924 3196
rect 2695 3190 2699 3191
rect 2726 3190 2732 3191
rect 2694 3185 2700 3186
rect 2727 3185 2731 3186
rect 2694 3181 2695 3185
rect 2699 3181 2700 3185
rect 2736 3184 2738 3194
rect 2918 3191 2919 3195
rect 2923 3191 2924 3195
rect 2918 3190 2924 3191
rect 2926 3195 2932 3196
rect 2926 3191 2927 3195
rect 2931 3191 2932 3195
rect 3110 3195 3116 3196
rect 3110 3191 3111 3195
rect 3115 3191 3116 3195
rect 2926 3190 2932 3191
rect 2935 3190 2939 3191
rect 3110 3190 3116 3191
rect 3118 3195 3124 3196
rect 3118 3191 3119 3195
rect 3123 3191 3124 3195
rect 3190 3195 3191 3199
rect 3195 3195 3196 3199
rect 3190 3194 3196 3195
rect 3192 3191 3194 3194
rect 3118 3190 3124 3191
rect 3159 3190 3163 3191
rect 2919 3185 2923 3186
rect 2694 3180 2700 3181
rect 2702 3183 2708 3184
rect 2182 3178 2188 3179
rect 2234 3179 2240 3180
rect 1854 3174 1860 3175
rect 1670 3163 1676 3164
rect 1670 3159 1671 3163
rect 1675 3159 1676 3163
rect 1670 3158 1676 3159
rect 1672 3151 1674 3158
rect 1846 3156 1852 3157
rect 1846 3152 1847 3156
rect 1851 3152 1852 3156
rect 1846 3151 1852 3152
rect 1671 3150 1675 3151
rect 1671 3145 1675 3146
rect 1695 3150 1699 3151
rect 1695 3145 1699 3146
rect 1847 3150 1851 3151
rect 1847 3145 1851 3146
rect 1672 3138 1674 3145
rect 1694 3144 1700 3145
rect 1694 3140 1695 3144
rect 1699 3140 1700 3144
rect 1694 3139 1700 3140
rect 1670 3137 1676 3138
rect 1670 3133 1671 3137
rect 1675 3133 1676 3137
rect 1670 3132 1676 3133
rect 111 3130 115 3131
rect 807 3130 811 3131
rect 1079 3130 1083 3131
rect 1351 3130 1355 3131
rect 1599 3130 1603 3131
rect 1631 3130 1635 3131
rect 1856 3128 1858 3174
rect 2038 3156 2044 3157
rect 2038 3152 2039 3156
rect 2043 3152 2044 3156
rect 2038 3151 2044 3152
rect 1863 3150 1867 3151
rect 1863 3145 1867 3146
rect 2023 3150 2027 3151
rect 2023 3145 2027 3146
rect 2039 3150 2043 3151
rect 2039 3145 2043 3146
rect 1862 3144 1868 3145
rect 1862 3140 1863 3144
rect 1867 3140 1868 3144
rect 1862 3139 1868 3140
rect 2022 3144 2028 3145
rect 2022 3140 2023 3144
rect 2027 3140 2028 3144
rect 2022 3139 2028 3140
rect 111 3125 115 3126
rect 806 3125 812 3126
rect 112 3122 114 3125
rect 110 3121 116 3122
rect 110 3117 111 3121
rect 115 3117 116 3121
rect 806 3121 807 3125
rect 811 3121 812 3125
rect 806 3120 812 3121
rect 1078 3125 1084 3126
rect 1078 3121 1079 3125
rect 1083 3121 1084 3125
rect 1078 3120 1084 3121
rect 1350 3125 1356 3126
rect 1350 3121 1351 3125
rect 1355 3121 1356 3125
rect 1350 3120 1356 3121
rect 1598 3125 1604 3126
rect 1631 3125 1635 3126
rect 1854 3127 1860 3128
rect 1598 3121 1599 3125
rect 1603 3121 1604 3125
rect 1632 3122 1634 3125
rect 1854 3123 1855 3127
rect 1859 3123 1860 3127
rect 1854 3122 1860 3123
rect 1598 3120 1604 3121
rect 1630 3121 1636 3122
rect 110 3116 116 3117
rect 838 3119 844 3120
rect 838 3115 839 3119
rect 843 3115 844 3119
rect 838 3114 844 3115
rect 1086 3119 1092 3120
rect 1086 3115 1087 3119
rect 1091 3115 1092 3119
rect 1086 3114 1092 3115
rect 1342 3119 1348 3120
rect 1342 3115 1343 3119
rect 1347 3115 1348 3119
rect 1630 3117 1631 3121
rect 1635 3117 1636 3121
rect 2048 3120 2050 3178
rect 2234 3175 2235 3179
rect 2239 3175 2240 3179
rect 2234 3174 2240 3175
rect 2554 3179 2560 3180
rect 2554 3175 2555 3179
rect 2559 3175 2560 3179
rect 2702 3179 2703 3183
rect 2707 3179 2708 3183
rect 2702 3178 2708 3179
rect 2734 3183 2740 3184
rect 2734 3179 2735 3183
rect 2739 3179 2740 3183
rect 2928 3180 2930 3190
rect 3191 3190 3195 3191
rect 2934 3185 2940 3186
rect 3111 3185 3115 3186
rect 3158 3185 3164 3186
rect 3191 3185 3195 3186
rect 2934 3181 2935 3185
rect 2939 3181 2940 3185
rect 2934 3180 2940 3181
rect 3158 3181 3159 3185
rect 3163 3181 3164 3185
rect 3192 3182 3194 3185
rect 3158 3180 3164 3181
rect 3190 3181 3196 3182
rect 2734 3178 2740 3179
rect 2926 3179 2932 3180
rect 2554 3174 2560 3175
rect 2183 3150 2187 3151
rect 2183 3145 2187 3146
rect 2182 3144 2188 3145
rect 2182 3140 2183 3144
rect 2187 3140 2188 3144
rect 2182 3139 2188 3140
rect 1630 3116 1636 3117
rect 1670 3119 1676 3120
rect 1342 3114 1348 3115
rect 1670 3115 1671 3119
rect 1675 3115 1676 3119
rect 1703 3119 1709 3120
rect 1670 3114 1676 3115
rect 1694 3115 1700 3116
rect 110 3103 116 3104
rect 110 3099 111 3103
rect 115 3099 116 3103
rect 110 3098 116 3099
rect 112 3087 114 3098
rect 806 3096 812 3097
rect 806 3092 807 3096
rect 811 3092 812 3096
rect 806 3091 812 3092
rect 808 3087 810 3091
rect 111 3086 115 3087
rect 111 3081 115 3082
rect 703 3086 707 3087
rect 703 3081 707 3082
rect 807 3086 811 3087
rect 807 3081 811 3082
rect 831 3086 835 3087
rect 831 3081 835 3082
rect 112 3074 114 3081
rect 702 3080 708 3081
rect 702 3076 703 3080
rect 707 3076 708 3080
rect 702 3075 708 3076
rect 830 3080 836 3081
rect 830 3076 831 3080
rect 835 3076 836 3080
rect 830 3075 836 3076
rect 110 3073 116 3074
rect 110 3069 111 3073
rect 115 3069 116 3073
rect 110 3068 116 3069
rect 840 3056 842 3114
rect 1078 3096 1084 3097
rect 1078 3092 1079 3096
rect 1083 3092 1084 3096
rect 1078 3091 1084 3092
rect 1080 3087 1082 3091
rect 959 3086 963 3087
rect 959 3081 963 3082
rect 1079 3086 1083 3087
rect 1079 3081 1083 3082
rect 958 3080 964 3081
rect 958 3076 959 3080
rect 963 3076 964 3080
rect 958 3075 964 3076
rect 1078 3080 1084 3081
rect 1078 3076 1079 3080
rect 1083 3076 1084 3080
rect 1078 3075 1084 3076
rect 1088 3056 1090 3114
rect 1199 3086 1203 3087
rect 1199 3081 1203 3082
rect 1311 3086 1315 3087
rect 1311 3081 1315 3082
rect 1198 3080 1204 3081
rect 1198 3076 1199 3080
rect 1203 3076 1204 3080
rect 1198 3075 1204 3076
rect 1310 3080 1316 3081
rect 1310 3076 1311 3080
rect 1315 3076 1316 3080
rect 1310 3075 1316 3076
rect 110 3055 116 3056
rect 110 3051 111 3055
rect 115 3051 116 3055
rect 838 3055 844 3056
rect 110 3050 116 3051
rect 702 3051 708 3052
rect 112 3039 114 3050
rect 702 3047 703 3051
rect 707 3047 708 3051
rect 702 3046 708 3047
rect 710 3051 716 3052
rect 710 3047 711 3051
rect 715 3047 716 3051
rect 710 3046 716 3047
rect 830 3051 836 3052
rect 830 3047 831 3051
rect 835 3047 836 3051
rect 838 3051 839 3055
rect 843 3051 844 3055
rect 1086 3055 1092 3056
rect 838 3050 844 3051
rect 958 3051 964 3052
rect 830 3046 836 3047
rect 704 3039 706 3046
rect 111 3038 115 3039
rect 623 3038 627 3039
rect 703 3038 707 3039
rect 111 3033 115 3034
rect 622 3033 628 3034
rect 703 3033 707 3034
rect 112 3030 114 3033
rect 110 3029 116 3030
rect 110 3025 111 3029
rect 115 3025 116 3029
rect 622 3029 623 3033
rect 627 3029 628 3033
rect 712 3032 714 3046
rect 832 3039 834 3046
rect 783 3038 787 3039
rect 831 3038 835 3039
rect 782 3033 788 3034
rect 831 3033 835 3034
rect 622 3028 628 3029
rect 630 3031 636 3032
rect 630 3027 631 3031
rect 635 3027 636 3031
rect 630 3026 636 3027
rect 710 3031 716 3032
rect 710 3027 711 3031
rect 715 3027 716 3031
rect 782 3029 783 3033
rect 787 3029 788 3033
rect 840 3032 842 3050
rect 958 3047 959 3051
rect 963 3047 964 3051
rect 958 3046 964 3047
rect 966 3051 972 3052
rect 966 3047 967 3051
rect 971 3047 972 3051
rect 966 3046 972 3047
rect 1078 3051 1084 3052
rect 1078 3047 1079 3051
rect 1083 3047 1084 3051
rect 1086 3051 1087 3055
rect 1091 3051 1092 3055
rect 1086 3050 1092 3051
rect 1198 3051 1204 3052
rect 1078 3046 1084 3047
rect 960 3039 962 3046
rect 927 3038 931 3039
rect 959 3038 963 3039
rect 926 3033 932 3034
rect 959 3033 963 3034
rect 782 3028 788 3029
rect 790 3031 796 3032
rect 710 3026 716 3027
rect 790 3027 791 3031
rect 795 3027 796 3031
rect 790 3026 796 3027
rect 838 3031 844 3032
rect 838 3027 839 3031
rect 843 3027 844 3031
rect 926 3029 927 3033
rect 931 3029 932 3033
rect 968 3032 970 3046
rect 1080 3039 1082 3046
rect 1063 3038 1067 3039
rect 1079 3038 1083 3039
rect 1062 3033 1068 3034
rect 1079 3033 1083 3034
rect 926 3028 932 3029
rect 934 3031 940 3032
rect 838 3026 844 3027
rect 934 3027 935 3031
rect 939 3027 940 3031
rect 934 3026 940 3027
rect 966 3031 972 3032
rect 966 3027 967 3031
rect 971 3027 972 3031
rect 1062 3029 1063 3033
rect 1067 3029 1068 3033
rect 1088 3032 1090 3050
rect 1198 3047 1199 3051
rect 1203 3047 1204 3051
rect 1198 3046 1204 3047
rect 1206 3051 1212 3052
rect 1206 3047 1207 3051
rect 1211 3047 1212 3051
rect 1206 3046 1212 3047
rect 1310 3051 1316 3052
rect 1310 3047 1311 3051
rect 1315 3047 1316 3051
rect 1310 3046 1316 3047
rect 1318 3051 1324 3052
rect 1318 3047 1319 3051
rect 1323 3047 1324 3051
rect 1318 3046 1324 3047
rect 1200 3039 1202 3046
rect 1191 3038 1195 3039
rect 1199 3038 1203 3039
rect 1190 3033 1196 3034
rect 1199 3033 1203 3034
rect 1062 3028 1068 3029
rect 1086 3031 1092 3032
rect 966 3026 972 3027
rect 1086 3027 1087 3031
rect 1091 3027 1092 3031
rect 1190 3029 1191 3033
rect 1195 3029 1196 3033
rect 1190 3028 1196 3029
rect 1086 3026 1092 3027
rect 1198 3027 1204 3028
rect 110 3024 116 3025
rect 110 3011 116 3012
rect 110 3007 111 3011
rect 115 3007 116 3011
rect 110 3006 116 3007
rect 112 2995 114 3006
rect 622 3004 628 3005
rect 622 3000 623 3004
rect 627 3000 628 3004
rect 622 2999 628 3000
rect 624 2995 626 2999
rect 111 2994 115 2995
rect 111 2989 115 2990
rect 519 2994 523 2995
rect 519 2989 523 2990
rect 623 2994 627 2995
rect 623 2989 627 2990
rect 112 2982 114 2989
rect 518 2988 524 2989
rect 518 2984 519 2988
rect 523 2984 524 2988
rect 518 2983 524 2984
rect 110 2981 116 2982
rect 110 2977 111 2981
rect 115 2977 116 2981
rect 110 2976 116 2977
rect 110 2963 116 2964
rect 110 2959 111 2963
rect 115 2959 116 2963
rect 110 2958 116 2959
rect 518 2959 524 2960
rect 112 2947 114 2958
rect 518 2955 519 2959
rect 523 2955 524 2959
rect 518 2954 524 2955
rect 478 2951 484 2952
rect 478 2947 479 2951
rect 483 2947 484 2951
rect 520 2947 522 2954
rect 632 2952 634 3026
rect 782 3004 788 3005
rect 782 3000 783 3004
rect 787 3000 788 3004
rect 782 2999 788 3000
rect 784 2995 786 2999
rect 647 2994 651 2995
rect 647 2989 651 2990
rect 783 2994 787 2995
rect 783 2989 787 2990
rect 646 2988 652 2989
rect 646 2984 647 2988
rect 651 2984 652 2988
rect 646 2983 652 2984
rect 782 2988 788 2989
rect 782 2984 783 2988
rect 787 2984 788 2988
rect 782 2983 788 2984
rect 792 2964 794 3026
rect 926 3004 932 3005
rect 926 3000 927 3004
rect 931 3000 932 3004
rect 926 2999 932 3000
rect 928 2995 930 2999
rect 919 2994 923 2995
rect 919 2989 923 2990
rect 927 2994 931 2995
rect 927 2989 931 2990
rect 918 2988 924 2989
rect 918 2984 919 2988
rect 923 2984 924 2988
rect 918 2983 924 2984
rect 790 2963 796 2964
rect 646 2959 652 2960
rect 646 2955 647 2959
rect 651 2955 652 2959
rect 646 2954 652 2955
rect 782 2959 788 2960
rect 782 2955 783 2959
rect 787 2955 788 2959
rect 790 2959 791 2963
rect 795 2959 796 2963
rect 790 2958 796 2959
rect 802 2963 808 2964
rect 802 2959 803 2963
rect 807 2959 808 2963
rect 927 2963 933 2964
rect 802 2958 808 2959
rect 918 2959 924 2960
rect 782 2954 788 2955
rect 630 2951 636 2952
rect 630 2947 631 2951
rect 635 2947 636 2951
rect 648 2947 650 2954
rect 784 2947 786 2954
rect 111 2946 115 2947
rect 439 2946 443 2947
rect 478 2946 484 2947
rect 519 2946 523 2947
rect 111 2941 115 2942
rect 438 2941 444 2942
rect 112 2938 114 2941
rect 110 2937 116 2938
rect 110 2933 111 2937
rect 115 2933 116 2937
rect 438 2937 439 2941
rect 443 2937 444 2941
rect 438 2936 444 2937
rect 480 2936 482 2946
rect 599 2946 603 2947
rect 630 2946 636 2947
rect 647 2946 651 2947
rect 759 2946 763 2947
rect 783 2946 787 2947
rect 519 2941 523 2942
rect 598 2941 604 2942
rect 647 2941 651 2942
rect 758 2941 764 2942
rect 783 2941 787 2942
rect 598 2937 599 2941
rect 603 2937 604 2941
rect 598 2936 604 2937
rect 758 2937 759 2941
rect 763 2937 764 2941
rect 758 2936 764 2937
rect 804 2936 806 2958
rect 918 2955 919 2959
rect 923 2955 924 2959
rect 927 2959 928 2963
rect 932 2962 933 2963
rect 936 2962 938 3026
rect 1062 3004 1068 3005
rect 1062 3000 1063 3004
rect 1067 3000 1068 3004
rect 1062 2999 1068 3000
rect 1064 2995 1066 2999
rect 1055 2994 1059 2995
rect 1055 2989 1059 2990
rect 1063 2994 1067 2995
rect 1063 2989 1067 2990
rect 1054 2988 1060 2989
rect 1054 2984 1055 2988
rect 1059 2984 1060 2988
rect 1054 2983 1060 2984
rect 1088 2964 1090 3026
rect 1198 3023 1199 3027
rect 1203 3026 1204 3027
rect 1208 3026 1210 3046
rect 1312 3039 1314 3046
rect 1311 3038 1315 3039
rect 1310 3033 1316 3034
rect 1310 3029 1311 3033
rect 1315 3029 1316 3033
rect 1310 3028 1316 3029
rect 1320 3028 1322 3046
rect 1344 3028 1346 3114
rect 1672 3111 1674 3114
rect 1694 3111 1695 3115
rect 1699 3111 1700 3115
rect 1703 3115 1704 3119
rect 1708 3118 1709 3119
rect 2046 3119 2052 3120
rect 1708 3116 1714 3118
rect 1708 3115 1709 3116
rect 1703 3114 1709 3115
rect 1671 3110 1675 3111
rect 1694 3110 1700 3111
rect 1671 3105 1675 3106
rect 1695 3105 1699 3106
rect 1630 3103 1636 3104
rect 1630 3099 1631 3103
rect 1635 3099 1636 3103
rect 1672 3102 1674 3105
rect 1630 3098 1636 3099
rect 1670 3101 1676 3102
rect 1350 3096 1356 3097
rect 1350 3092 1351 3096
rect 1355 3092 1356 3096
rect 1350 3091 1356 3092
rect 1598 3096 1604 3097
rect 1598 3092 1599 3096
rect 1603 3092 1604 3096
rect 1598 3091 1604 3092
rect 1352 3087 1354 3091
rect 1600 3087 1602 3091
rect 1632 3087 1634 3098
rect 1670 3097 1671 3101
rect 1675 3097 1676 3101
rect 1670 3096 1676 3097
rect 1351 3086 1355 3087
rect 1351 3081 1355 3082
rect 1423 3086 1427 3087
rect 1423 3081 1427 3082
rect 1543 3086 1547 3087
rect 1543 3081 1547 3082
rect 1599 3086 1603 3087
rect 1599 3081 1603 3082
rect 1631 3086 1635 3087
rect 1631 3081 1635 3082
rect 1670 3083 1676 3084
rect 1422 3080 1428 3081
rect 1422 3076 1423 3080
rect 1427 3076 1428 3080
rect 1422 3075 1428 3076
rect 1542 3080 1548 3081
rect 1542 3076 1543 3080
rect 1547 3076 1548 3080
rect 1542 3075 1548 3076
rect 1632 3074 1634 3081
rect 1670 3079 1671 3083
rect 1675 3079 1676 3083
rect 1670 3078 1676 3079
rect 1630 3073 1636 3074
rect 1630 3069 1631 3073
rect 1635 3069 1636 3073
rect 1672 3071 1674 3078
rect 1712 3073 1714 3116
rect 1862 3115 1868 3116
rect 1862 3111 1863 3115
rect 1867 3111 1868 3115
rect 2022 3115 2028 3116
rect 2022 3111 2023 3115
rect 2027 3111 2028 3115
rect 2046 3115 2047 3119
rect 2051 3115 2052 3119
rect 2236 3116 2238 3174
rect 2246 3156 2252 3157
rect 2246 3152 2247 3156
rect 2251 3152 2252 3156
rect 2246 3151 2252 3152
rect 2462 3156 2468 3157
rect 2462 3152 2463 3156
rect 2467 3152 2468 3156
rect 2462 3151 2468 3152
rect 2247 3150 2251 3151
rect 2247 3145 2251 3146
rect 2343 3150 2347 3151
rect 2343 3145 2347 3146
rect 2463 3150 2467 3151
rect 2463 3145 2467 3146
rect 2511 3150 2515 3151
rect 2511 3145 2515 3146
rect 2342 3144 2348 3145
rect 2342 3140 2343 3144
rect 2347 3140 2348 3144
rect 2342 3139 2348 3140
rect 2510 3144 2516 3145
rect 2510 3140 2511 3144
rect 2515 3140 2516 3144
rect 2510 3139 2516 3140
rect 2556 3120 2558 3174
rect 2694 3156 2700 3157
rect 2694 3152 2695 3156
rect 2699 3152 2700 3156
rect 2694 3151 2700 3152
rect 2695 3150 2699 3151
rect 2695 3145 2699 3146
rect 2554 3119 2560 3120
rect 2046 3114 2052 3115
rect 2182 3115 2188 3116
rect 1862 3110 1868 3111
rect 1959 3110 1963 3111
rect 2022 3110 2028 3111
rect 1863 3105 1867 3106
rect 1878 3107 1884 3108
rect 1878 3103 1879 3107
rect 1883 3103 1884 3107
rect 1878 3102 1884 3103
rect 1958 3105 1964 3106
rect 2023 3105 2027 3106
rect 1880 3100 1882 3102
rect 1958 3101 1959 3105
rect 1963 3101 1964 3105
rect 1958 3100 1964 3101
rect 2048 3100 2050 3114
rect 2182 3111 2183 3115
rect 2187 3111 2188 3115
rect 2182 3110 2188 3111
rect 2234 3115 2240 3116
rect 2234 3111 2235 3115
rect 2239 3111 2240 3115
rect 2234 3110 2240 3111
rect 2342 3115 2348 3116
rect 2342 3111 2343 3115
rect 2347 3111 2348 3115
rect 2510 3115 2516 3116
rect 2510 3111 2511 3115
rect 2515 3111 2516 3115
rect 2554 3115 2555 3119
rect 2559 3115 2560 3119
rect 2554 3114 2560 3115
rect 2342 3110 2348 3111
rect 2415 3110 2419 3111
rect 2510 3110 2516 3111
rect 2655 3110 2659 3111
rect 2182 3105 2188 3106
rect 2343 3105 2347 3106
rect 2414 3105 2420 3106
rect 2511 3105 2515 3106
rect 2654 3105 2660 3106
rect 2182 3101 2183 3105
rect 2187 3101 2188 3105
rect 2182 3100 2188 3101
rect 2414 3101 2415 3105
rect 2419 3101 2420 3105
rect 2414 3100 2420 3101
rect 2654 3101 2655 3105
rect 2659 3101 2660 3105
rect 2704 3104 2706 3178
rect 2926 3175 2927 3179
rect 2931 3175 2932 3179
rect 3190 3177 3191 3181
rect 3195 3177 3196 3181
rect 3190 3176 3196 3177
rect 2926 3174 2932 3175
rect 2903 3110 2907 3111
rect 2902 3105 2908 3106
rect 2654 3100 2660 3101
rect 2662 3103 2668 3104
rect 1878 3099 1884 3100
rect 1878 3095 1879 3099
rect 1883 3095 1884 3099
rect 1878 3094 1884 3095
rect 2046 3099 2052 3100
rect 2046 3095 2047 3099
rect 2051 3095 2052 3099
rect 2662 3099 2663 3103
rect 2667 3099 2668 3103
rect 2662 3098 2668 3099
rect 2702 3103 2708 3104
rect 2702 3099 2703 3103
rect 2707 3099 2708 3103
rect 2902 3101 2903 3105
rect 2907 3101 2908 3105
rect 2902 3100 2908 3101
rect 2928 3100 2930 3174
rect 3190 3163 3196 3164
rect 3190 3159 3191 3163
rect 3195 3159 3196 3163
rect 3190 3158 3196 3159
rect 2934 3156 2940 3157
rect 2934 3152 2935 3156
rect 2939 3152 2940 3156
rect 2934 3151 2940 3152
rect 3158 3156 3164 3157
rect 3158 3152 3159 3156
rect 3163 3152 3164 3156
rect 3158 3151 3164 3152
rect 3192 3151 3194 3158
rect 2935 3150 2939 3151
rect 2935 3145 2939 3146
rect 3159 3150 3163 3151
rect 3159 3145 3163 3146
rect 3191 3150 3195 3151
rect 3191 3145 3195 3146
rect 3192 3138 3194 3145
rect 3190 3137 3196 3138
rect 3190 3133 3191 3137
rect 3195 3133 3196 3137
rect 3190 3132 3196 3133
rect 3190 3119 3196 3120
rect 3190 3115 3191 3119
rect 3195 3115 3196 3119
rect 3190 3114 3196 3115
rect 3192 3111 3194 3114
rect 3159 3110 3163 3111
rect 3191 3110 3195 3111
rect 3158 3105 3164 3106
rect 3191 3105 3195 3106
rect 3158 3101 3159 3105
rect 3163 3101 3164 3105
rect 3192 3102 3194 3105
rect 3158 3100 3164 3101
rect 3190 3101 3196 3102
rect 2702 3098 2708 3099
rect 2910 3099 2916 3100
rect 2046 3094 2052 3095
rect 1712 3071 1718 3073
rect 1630 3068 1636 3069
rect 1671 3070 1675 3071
rect 1671 3065 1675 3066
rect 1672 3058 1674 3065
rect 1670 3057 1676 3058
rect 1446 3055 1452 3056
rect 1422 3051 1428 3052
rect 1422 3047 1423 3051
rect 1427 3047 1428 3051
rect 1446 3051 1447 3055
rect 1451 3051 1452 3055
rect 1630 3055 1636 3056
rect 1446 3050 1452 3051
rect 1542 3051 1548 3052
rect 1422 3046 1428 3047
rect 1424 3039 1426 3046
rect 1423 3038 1427 3039
rect 1439 3038 1443 3039
rect 1423 3033 1427 3034
rect 1438 3033 1444 3034
rect 1438 3029 1439 3033
rect 1443 3029 1444 3033
rect 1448 3032 1450 3050
rect 1542 3047 1543 3051
rect 1547 3047 1548 3051
rect 1630 3051 1631 3055
rect 1635 3051 1636 3055
rect 1670 3053 1671 3057
rect 1675 3053 1676 3057
rect 1670 3052 1676 3053
rect 1630 3050 1636 3051
rect 1542 3046 1548 3047
rect 1544 3039 1546 3046
rect 1632 3039 1634 3050
rect 1670 3039 1676 3040
rect 1543 3038 1547 3039
rect 1543 3033 1547 3034
rect 1631 3038 1635 3039
rect 1670 3035 1671 3039
rect 1675 3035 1676 3039
rect 1670 3034 1676 3035
rect 1631 3033 1635 3034
rect 1438 3028 1444 3029
rect 1446 3031 1452 3032
rect 1203 3024 1210 3026
rect 1318 3027 1324 3028
rect 1203 3023 1204 3024
rect 1198 3022 1204 3023
rect 1318 3023 1319 3027
rect 1323 3023 1324 3027
rect 1318 3022 1324 3023
rect 1342 3027 1348 3028
rect 1342 3023 1343 3027
rect 1347 3023 1348 3027
rect 1446 3027 1447 3031
rect 1451 3027 1452 3031
rect 1632 3030 1634 3033
rect 1672 3031 1674 3034
rect 1671 3030 1675 3031
rect 1446 3026 1452 3027
rect 1630 3029 1636 3030
rect 1342 3022 1348 3023
rect 1190 3004 1196 3005
rect 1190 3000 1191 3004
rect 1195 3000 1196 3004
rect 1190 2999 1196 3000
rect 1192 2995 1194 2999
rect 1191 2994 1195 2995
rect 1191 2989 1195 2990
rect 1190 2988 1196 2989
rect 1190 2984 1191 2988
rect 1195 2984 1196 2988
rect 1190 2983 1196 2984
rect 1200 2968 1202 3022
rect 1310 3004 1316 3005
rect 1310 3000 1311 3004
rect 1315 3000 1316 3004
rect 1310 2999 1316 3000
rect 1312 2995 1314 2999
rect 1311 2994 1315 2995
rect 1311 2989 1315 2990
rect 1335 2994 1339 2995
rect 1335 2989 1339 2990
rect 1334 2988 1340 2989
rect 1334 2984 1335 2988
rect 1339 2984 1340 2988
rect 1334 2983 1340 2984
rect 1198 2967 1204 2968
rect 932 2960 938 2962
rect 1086 2963 1092 2964
rect 932 2959 933 2960
rect 927 2958 933 2959
rect 918 2954 924 2955
rect 920 2947 922 2954
rect 919 2946 923 2947
rect 927 2946 931 2947
rect 919 2941 923 2942
rect 926 2941 932 2942
rect 926 2937 927 2941
rect 931 2937 932 2941
rect 926 2936 932 2937
rect 936 2936 938 2960
rect 1054 2959 1060 2960
rect 1054 2955 1055 2959
rect 1059 2955 1060 2959
rect 1086 2959 1087 2963
rect 1091 2959 1092 2963
rect 1086 2958 1092 2959
rect 1102 2963 1108 2964
rect 1102 2959 1103 2963
rect 1107 2959 1108 2963
rect 1198 2963 1199 2967
rect 1203 2963 1204 2967
rect 1198 2962 1204 2963
rect 1344 2960 1346 3022
rect 1438 3004 1444 3005
rect 1438 3000 1439 3004
rect 1443 3000 1444 3004
rect 1438 2999 1444 3000
rect 1440 2995 1442 2999
rect 1439 2994 1443 2995
rect 1439 2989 1443 2990
rect 1102 2958 1108 2959
rect 1190 2959 1196 2960
rect 1054 2954 1060 2955
rect 1056 2947 1058 2954
rect 1055 2946 1059 2947
rect 1095 2946 1099 2947
rect 1055 2941 1059 2942
rect 1094 2941 1100 2942
rect 1094 2937 1095 2941
rect 1099 2937 1100 2941
rect 1094 2936 1100 2937
rect 1104 2936 1106 2958
rect 1190 2955 1191 2959
rect 1195 2955 1196 2959
rect 1190 2954 1196 2955
rect 1334 2959 1340 2960
rect 1334 2955 1335 2959
rect 1339 2955 1340 2959
rect 1334 2954 1340 2955
rect 1342 2959 1348 2960
rect 1342 2955 1343 2959
rect 1347 2955 1348 2959
rect 1342 2954 1348 2955
rect 1192 2947 1194 2954
rect 1336 2947 1338 2954
rect 1191 2946 1195 2947
rect 1263 2946 1267 2947
rect 1335 2946 1339 2947
rect 1191 2941 1195 2942
rect 1262 2941 1268 2942
rect 1335 2941 1339 2942
rect 1262 2937 1263 2941
rect 1267 2937 1268 2941
rect 1262 2936 1268 2937
rect 1344 2936 1346 2954
rect 1439 2946 1443 2947
rect 1438 2941 1444 2942
rect 1438 2937 1439 2941
rect 1443 2937 1444 2941
rect 1448 2940 1450 3026
rect 1630 3025 1631 3029
rect 1635 3025 1636 3029
rect 1671 3025 1675 3026
rect 1630 3024 1636 3025
rect 1672 3022 1674 3025
rect 1670 3021 1676 3022
rect 1670 3017 1671 3021
rect 1675 3017 1676 3021
rect 1716 3020 1718 3071
rect 1871 3070 1875 3071
rect 1871 3065 1875 3066
rect 1870 3064 1876 3065
rect 1870 3060 1871 3064
rect 1875 3060 1876 3064
rect 1870 3059 1876 3060
rect 1880 3040 1882 3094
rect 1958 3076 1964 3077
rect 1958 3072 1959 3076
rect 1963 3072 1964 3076
rect 1958 3071 1964 3072
rect 2182 3076 2188 3077
rect 2182 3072 2183 3076
rect 2187 3072 2188 3076
rect 2182 3071 2188 3072
rect 2414 3076 2420 3077
rect 2414 3072 2415 3076
rect 2419 3072 2420 3076
rect 2414 3071 2420 3072
rect 2654 3076 2660 3077
rect 2654 3072 2655 3076
rect 2659 3072 2660 3076
rect 2654 3071 2660 3072
rect 1959 3070 1963 3071
rect 1959 3065 1963 3066
rect 2111 3070 2115 3071
rect 2111 3065 2115 3066
rect 2183 3070 2187 3071
rect 2183 3065 2187 3066
rect 2367 3070 2371 3071
rect 2367 3065 2371 3066
rect 2415 3070 2419 3071
rect 2415 3065 2419 3066
rect 2631 3070 2635 3071
rect 2631 3065 2635 3066
rect 2655 3070 2659 3071
rect 2655 3065 2659 3066
rect 2110 3064 2116 3065
rect 2110 3060 2111 3064
rect 2115 3060 2116 3064
rect 2110 3059 2116 3060
rect 2366 3064 2372 3065
rect 2366 3060 2367 3064
rect 2371 3060 2372 3064
rect 2366 3059 2372 3060
rect 2630 3064 2636 3065
rect 2630 3060 2631 3064
rect 2635 3060 2636 3064
rect 2630 3059 2636 3060
rect 2664 3040 2666 3098
rect 2910 3095 2911 3099
rect 2915 3095 2916 3099
rect 2910 3094 2916 3095
rect 2926 3099 2932 3100
rect 2926 3095 2927 3099
rect 2931 3095 2932 3099
rect 2926 3094 2932 3095
rect 3166 3099 3172 3100
rect 3166 3095 3167 3099
rect 3171 3095 3172 3099
rect 3190 3097 3191 3101
rect 3195 3097 3196 3101
rect 3190 3096 3196 3097
rect 3166 3094 3172 3095
rect 2902 3076 2908 3077
rect 2902 3072 2903 3076
rect 2907 3072 2908 3076
rect 2902 3071 2908 3072
rect 2903 3070 2907 3071
rect 2903 3065 2907 3066
rect 2902 3064 2908 3065
rect 2902 3060 2903 3064
rect 2907 3060 2908 3064
rect 2902 3059 2908 3060
rect 1878 3039 1884 3040
rect 1870 3035 1876 3036
rect 1870 3031 1871 3035
rect 1875 3031 1876 3035
rect 1878 3035 1879 3039
rect 1883 3035 1884 3039
rect 2662 3039 2668 3040
rect 1878 3034 1884 3035
rect 2110 3035 2116 3036
rect 1791 3030 1795 3031
rect 1870 3030 1876 3031
rect 1790 3025 1796 3026
rect 1871 3025 1875 3026
rect 1790 3021 1791 3025
rect 1795 3021 1796 3025
rect 1790 3020 1796 3021
rect 1880 3020 1882 3034
rect 2110 3031 2111 3035
rect 2115 3031 2116 3035
rect 2134 3035 2140 3036
rect 2134 3031 2135 3035
rect 2139 3031 2140 3035
rect 2366 3035 2372 3036
rect 2366 3031 2367 3035
rect 2371 3031 2372 3035
rect 2630 3035 2636 3036
rect 2630 3031 2631 3035
rect 2635 3031 2636 3035
rect 2662 3035 2663 3039
rect 2667 3035 2668 3039
rect 2912 3036 2914 3094
rect 3158 3076 3164 3077
rect 3158 3072 3159 3076
rect 3163 3072 3164 3076
rect 3158 3071 3164 3072
rect 3159 3070 3163 3071
rect 3159 3065 3163 3066
rect 3158 3064 3164 3065
rect 3158 3060 3159 3064
rect 3163 3060 3164 3064
rect 3158 3059 3164 3060
rect 3168 3040 3170 3094
rect 3190 3083 3196 3084
rect 3190 3079 3191 3083
rect 3195 3079 3196 3083
rect 3190 3078 3196 3079
rect 3192 3071 3194 3078
rect 3191 3070 3195 3071
rect 3191 3065 3195 3066
rect 3192 3058 3194 3065
rect 3190 3057 3196 3058
rect 3190 3053 3191 3057
rect 3195 3053 3196 3057
rect 3190 3052 3196 3053
rect 3166 3039 3172 3040
rect 2662 3034 2668 3035
rect 2902 3035 2908 3036
rect 1959 3030 1963 3031
rect 2110 3030 2116 3031
rect 2127 3030 2131 3031
rect 2134 3030 2140 3031
rect 2287 3030 2291 3031
rect 2366 3030 2372 3031
rect 2455 3030 2459 3031
rect 1958 3025 1964 3026
rect 2111 3025 2115 3026
rect 2126 3025 2132 3026
rect 1958 3021 1959 3025
rect 1963 3021 1964 3025
rect 1958 3020 1964 3021
rect 2126 3021 2127 3025
rect 2131 3021 2132 3025
rect 2126 3020 2132 3021
rect 2136 3020 2138 3030
rect 2623 3030 2627 3031
rect 2630 3030 2636 3031
rect 2902 3031 2903 3035
rect 2907 3031 2908 3035
rect 2902 3030 2908 3031
rect 2910 3035 2916 3036
rect 2910 3031 2911 3035
rect 2915 3031 2916 3035
rect 2910 3030 2916 3031
rect 3158 3035 3164 3036
rect 3158 3031 3159 3035
rect 3163 3031 3164 3035
rect 3166 3035 3167 3039
rect 3171 3035 3172 3039
rect 3166 3034 3172 3035
rect 3190 3039 3196 3040
rect 3190 3035 3191 3039
rect 3195 3035 3196 3039
rect 3190 3034 3196 3035
rect 3158 3030 3164 3031
rect 2286 3025 2292 3026
rect 2367 3025 2371 3026
rect 2454 3025 2460 3026
rect 2286 3021 2287 3025
rect 2291 3021 2292 3025
rect 2286 3020 2292 3021
rect 2294 3023 2300 3024
rect 1670 3016 1676 3017
rect 1714 3019 1720 3020
rect 1714 3015 1715 3019
rect 1719 3015 1720 3019
rect 1714 3014 1720 3015
rect 1878 3019 1884 3020
rect 1878 3015 1879 3019
rect 1883 3015 1884 3019
rect 1878 3014 1884 3015
rect 1910 3019 1916 3020
rect 1910 3015 1911 3019
rect 1915 3015 1916 3019
rect 1910 3014 1916 3015
rect 2134 3019 2140 3020
rect 2134 3015 2135 3019
rect 2139 3015 2140 3019
rect 2294 3019 2295 3023
rect 2299 3019 2300 3023
rect 2454 3021 2455 3025
rect 2459 3021 2460 3025
rect 2454 3020 2460 3021
rect 2622 3025 2628 3026
rect 2631 3025 2635 3026
rect 2903 3025 2907 3026
rect 2622 3021 2623 3025
rect 2627 3021 2628 3025
rect 2622 3020 2628 3021
rect 2294 3018 2300 3019
rect 2378 3019 2384 3020
rect 2134 3014 2140 3015
rect 1630 3011 1636 3012
rect 1630 3007 1631 3011
rect 1635 3007 1636 3011
rect 1630 3006 1636 3007
rect 1632 2995 1634 3006
rect 1670 3003 1676 3004
rect 1670 2999 1671 3003
rect 1675 2999 1676 3003
rect 1670 2998 1676 2999
rect 1631 2994 1635 2995
rect 1672 2991 1674 2998
rect 1631 2989 1635 2990
rect 1671 2990 1675 2991
rect 1632 2982 1634 2989
rect 1671 2985 1675 2986
rect 1703 2990 1707 2991
rect 1703 2985 1707 2986
rect 1630 2981 1636 2982
rect 1630 2977 1631 2981
rect 1635 2977 1636 2981
rect 1672 2978 1674 2985
rect 1702 2984 1708 2985
rect 1702 2980 1703 2984
rect 1707 2980 1708 2984
rect 1702 2979 1708 2980
rect 1630 2976 1636 2977
rect 1670 2977 1676 2978
rect 1670 2973 1671 2977
rect 1675 2973 1676 2977
rect 1670 2972 1676 2973
rect 1630 2963 1636 2964
rect 1630 2959 1631 2963
rect 1635 2959 1636 2963
rect 1716 2960 1718 3014
rect 1790 2996 1796 2997
rect 1790 2992 1791 2996
rect 1795 2992 1796 2996
rect 1790 2991 1796 2992
rect 1791 2990 1795 2991
rect 1791 2985 1795 2986
rect 1903 2990 1907 2991
rect 1903 2985 1907 2986
rect 1902 2984 1908 2985
rect 1902 2980 1903 2984
rect 1907 2980 1908 2984
rect 1902 2979 1908 2980
rect 1912 2960 1914 3014
rect 1958 2996 1964 2997
rect 1958 2992 1959 2996
rect 1963 2992 1964 2996
rect 1958 2991 1964 2992
rect 2126 2996 2132 2997
rect 2126 2992 2127 2996
rect 2131 2992 2132 2996
rect 2126 2991 2132 2992
rect 1959 2990 1963 2991
rect 1959 2985 1963 2986
rect 2127 2990 2131 2991
rect 2127 2985 2131 2986
rect 2126 2984 2132 2985
rect 2126 2980 2127 2984
rect 2131 2980 2132 2984
rect 2126 2979 2132 2980
rect 1630 2958 1636 2959
rect 1670 2959 1676 2960
rect 1632 2947 1634 2958
rect 1670 2955 1671 2959
rect 1675 2955 1676 2959
rect 1714 2959 1720 2960
rect 1670 2954 1676 2955
rect 1702 2955 1708 2956
rect 1672 2951 1674 2954
rect 1702 2951 1703 2955
rect 1707 2951 1708 2955
rect 1714 2955 1715 2959
rect 1719 2955 1720 2959
rect 1910 2959 1916 2960
rect 1714 2954 1720 2955
rect 1902 2955 1908 2956
rect 1671 2950 1675 2951
rect 1599 2946 1603 2947
rect 1631 2946 1635 2947
rect 1695 2950 1699 2951
rect 1702 2950 1708 2951
rect 1671 2945 1675 2946
rect 1694 2945 1700 2946
rect 1703 2945 1707 2946
rect 1672 2942 1674 2945
rect 1598 2941 1604 2942
rect 1631 2941 1635 2942
rect 1670 2941 1676 2942
rect 1438 2936 1444 2937
rect 1446 2939 1452 2940
rect 110 2932 116 2933
rect 478 2935 484 2936
rect 478 2931 479 2935
rect 483 2931 484 2935
rect 478 2930 484 2931
rect 802 2935 808 2936
rect 802 2931 803 2935
rect 807 2931 808 2935
rect 802 2930 808 2931
rect 934 2935 940 2936
rect 934 2931 935 2935
rect 939 2931 940 2935
rect 934 2930 940 2931
rect 1102 2935 1108 2936
rect 1102 2931 1103 2935
rect 1107 2931 1108 2935
rect 1102 2930 1108 2931
rect 1342 2935 1348 2936
rect 1342 2931 1343 2935
rect 1347 2931 1348 2935
rect 1446 2935 1447 2939
rect 1451 2935 1452 2939
rect 1598 2937 1599 2941
rect 1603 2937 1604 2941
rect 1632 2938 1634 2941
rect 1598 2936 1604 2937
rect 1630 2937 1636 2938
rect 1446 2934 1452 2935
rect 1630 2933 1631 2937
rect 1635 2933 1636 2937
rect 1670 2937 1671 2941
rect 1675 2937 1676 2941
rect 1694 2941 1695 2945
rect 1699 2941 1700 2945
rect 1716 2944 1718 2954
rect 1902 2951 1903 2955
rect 1907 2951 1908 2955
rect 1910 2955 1911 2959
rect 1915 2955 1916 2959
rect 2136 2956 2138 3014
rect 2286 2996 2292 2997
rect 2286 2992 2287 2996
rect 2291 2992 2292 2996
rect 2286 2991 2292 2992
rect 2287 2990 2291 2991
rect 2287 2985 2291 2986
rect 1910 2954 1916 2955
rect 2126 2955 2132 2956
rect 1902 2950 1908 2951
rect 1903 2945 1907 2946
rect 1694 2940 1700 2941
rect 1714 2943 1720 2944
rect 1714 2939 1715 2943
rect 1719 2939 1720 2943
rect 1912 2940 1914 2954
rect 2126 2951 2127 2955
rect 2131 2951 2132 2955
rect 1935 2950 1939 2951
rect 2126 2950 2132 2951
rect 2134 2955 2140 2956
rect 2134 2951 2135 2955
rect 2139 2951 2140 2955
rect 2230 2955 2236 2956
rect 2230 2951 2231 2955
rect 2235 2951 2236 2955
rect 2134 2950 2140 2951
rect 2223 2950 2227 2951
rect 2230 2950 2236 2951
rect 1934 2945 1940 2946
rect 2127 2945 2131 2946
rect 2222 2945 2228 2946
rect 1934 2941 1935 2945
rect 1939 2941 1940 2945
rect 1934 2940 1940 2941
rect 2222 2941 2223 2945
rect 2227 2941 2228 2945
rect 2222 2940 2228 2941
rect 2232 2940 2234 2950
rect 2296 2944 2298 3018
rect 2378 3015 2379 3019
rect 2383 3015 2384 3019
rect 2378 3014 2384 3015
rect 2526 3019 2532 3020
rect 2526 3015 2527 3019
rect 2531 3015 2532 3019
rect 2526 3014 2532 3015
rect 2630 3019 2636 3020
rect 2630 3015 2631 3019
rect 2635 3015 2636 3019
rect 2630 3014 2636 3015
rect 2367 2990 2371 2991
rect 2367 2985 2371 2986
rect 2366 2984 2372 2985
rect 2366 2980 2367 2984
rect 2371 2980 2372 2984
rect 2366 2979 2372 2980
rect 2380 2960 2382 3014
rect 2454 2996 2460 2997
rect 2454 2992 2455 2996
rect 2459 2992 2460 2996
rect 2454 2991 2460 2992
rect 2455 2990 2459 2991
rect 2455 2985 2459 2986
rect 2378 2959 2384 2960
rect 2366 2955 2372 2956
rect 2366 2951 2367 2955
rect 2371 2951 2372 2955
rect 2378 2955 2379 2959
rect 2383 2955 2384 2959
rect 2378 2954 2384 2955
rect 2366 2950 2372 2951
rect 2519 2950 2523 2951
rect 2367 2945 2371 2946
rect 2518 2945 2524 2946
rect 2294 2943 2300 2944
rect 1714 2938 1720 2939
rect 1910 2939 1916 2940
rect 1670 2936 1676 2937
rect 1910 2935 1911 2939
rect 1915 2935 1916 2939
rect 1910 2934 1916 2935
rect 2230 2939 2236 2940
rect 2230 2935 2231 2939
rect 2235 2935 2236 2939
rect 2294 2939 2295 2943
rect 2299 2939 2300 2943
rect 2518 2941 2519 2945
rect 2523 2941 2524 2945
rect 2528 2944 2530 3014
rect 2622 2996 2628 2997
rect 2622 2992 2623 2996
rect 2627 2992 2628 2996
rect 2622 2991 2628 2992
rect 2623 2990 2627 2991
rect 2623 2985 2627 2986
rect 2622 2984 2628 2985
rect 2622 2980 2623 2984
rect 2627 2980 2628 2984
rect 2622 2979 2628 2980
rect 2632 2960 2634 3014
rect 2887 2990 2891 2991
rect 2887 2985 2891 2986
rect 2886 2984 2892 2985
rect 2886 2980 2887 2984
rect 2891 2980 2892 2984
rect 2886 2979 2892 2980
rect 2630 2959 2636 2960
rect 2622 2955 2628 2956
rect 2622 2951 2623 2955
rect 2627 2951 2628 2955
rect 2630 2955 2631 2959
rect 2635 2955 2636 2959
rect 2912 2956 2914 3030
rect 3159 3025 3163 3026
rect 3159 2990 3163 2991
rect 3159 2985 3163 2986
rect 3158 2984 3164 2985
rect 3158 2980 3159 2984
rect 3163 2980 3164 2984
rect 3158 2979 3164 2980
rect 3168 2960 3170 3034
rect 3192 3031 3194 3034
rect 3191 3030 3195 3031
rect 3191 3025 3195 3026
rect 3192 3022 3194 3025
rect 3190 3021 3196 3022
rect 3190 3017 3191 3021
rect 3195 3017 3196 3021
rect 3190 3016 3196 3017
rect 3190 3003 3196 3004
rect 3190 2999 3191 3003
rect 3195 2999 3196 3003
rect 3190 2998 3196 2999
rect 3192 2991 3194 2998
rect 3191 2990 3195 2991
rect 3191 2985 3195 2986
rect 3192 2978 3194 2985
rect 3190 2977 3196 2978
rect 3190 2973 3191 2977
rect 3195 2973 3196 2977
rect 3190 2972 3196 2973
rect 3166 2959 3172 2960
rect 2630 2954 2636 2955
rect 2886 2955 2892 2956
rect 2886 2951 2887 2955
rect 2891 2951 2892 2955
rect 2622 2950 2628 2951
rect 2823 2950 2827 2951
rect 2886 2950 2892 2951
rect 2910 2955 2916 2956
rect 2910 2951 2911 2955
rect 2915 2951 2916 2955
rect 3158 2955 3164 2956
rect 3158 2951 3159 2955
rect 3163 2951 3164 2955
rect 3166 2955 3167 2959
rect 3171 2955 3172 2959
rect 3166 2954 3172 2955
rect 3190 2959 3196 2960
rect 3190 2955 3191 2959
rect 3195 2955 3196 2959
rect 3190 2954 3196 2955
rect 2910 2950 2916 2951
rect 3135 2950 3139 2951
rect 3158 2950 3164 2951
rect 2623 2945 2627 2946
rect 2822 2945 2828 2946
rect 2887 2945 2891 2946
rect 3134 2945 3140 2946
rect 3159 2945 3163 2946
rect 2518 2940 2524 2941
rect 2526 2943 2532 2944
rect 2294 2938 2300 2939
rect 2526 2939 2527 2943
rect 2531 2939 2532 2943
rect 2822 2941 2823 2945
rect 2827 2941 2828 2945
rect 2822 2940 2828 2941
rect 3134 2941 3135 2945
rect 3139 2941 3140 2945
rect 3168 2944 3170 2954
rect 3192 2951 3194 2954
rect 3191 2950 3195 2951
rect 3191 2945 3195 2946
rect 3134 2940 3140 2941
rect 3142 2943 3148 2944
rect 2526 2938 2532 2939
rect 2834 2939 2840 2940
rect 2230 2934 2236 2935
rect 1630 2932 1636 2933
rect 1342 2930 1348 2931
rect 1610 2931 1616 2932
rect 110 2919 116 2920
rect 110 2915 111 2919
rect 115 2915 116 2919
rect 110 2914 116 2915
rect 112 2907 114 2914
rect 438 2912 444 2913
rect 438 2908 439 2912
rect 443 2908 444 2912
rect 438 2907 444 2908
rect 111 2906 115 2907
rect 111 2901 115 2902
rect 335 2906 339 2907
rect 335 2901 339 2902
rect 439 2906 443 2907
rect 439 2901 443 2902
rect 471 2906 475 2907
rect 471 2901 475 2902
rect 112 2894 114 2901
rect 334 2900 340 2901
rect 334 2896 335 2900
rect 339 2896 340 2900
rect 334 2895 340 2896
rect 470 2900 476 2901
rect 470 2896 471 2900
rect 475 2896 476 2900
rect 470 2895 476 2896
rect 110 2893 116 2894
rect 110 2889 111 2893
rect 115 2889 116 2893
rect 110 2888 116 2889
rect 110 2875 116 2876
rect 110 2871 111 2875
rect 115 2871 116 2875
rect 480 2872 482 2930
rect 598 2912 604 2913
rect 598 2908 599 2912
rect 603 2908 604 2912
rect 598 2907 604 2908
rect 758 2912 764 2913
rect 758 2908 759 2912
rect 763 2908 764 2912
rect 758 2907 764 2908
rect 599 2906 603 2907
rect 599 2901 603 2902
rect 623 2906 627 2907
rect 623 2901 627 2902
rect 759 2906 763 2907
rect 759 2901 763 2902
rect 791 2906 795 2907
rect 791 2901 795 2902
rect 622 2900 628 2901
rect 622 2896 623 2900
rect 627 2896 628 2900
rect 622 2895 628 2896
rect 790 2900 796 2901
rect 790 2896 791 2900
rect 795 2896 796 2900
rect 790 2895 796 2896
rect 804 2872 806 2930
rect 926 2912 932 2913
rect 926 2908 927 2912
rect 931 2908 932 2912
rect 926 2907 932 2908
rect 927 2906 931 2907
rect 927 2901 931 2902
rect 110 2870 116 2871
rect 334 2871 340 2872
rect 112 2859 114 2870
rect 334 2867 335 2871
rect 339 2867 340 2871
rect 334 2866 340 2867
rect 470 2871 476 2872
rect 470 2867 471 2871
rect 475 2867 476 2871
rect 470 2866 476 2867
rect 478 2871 484 2872
rect 478 2867 479 2871
rect 483 2867 484 2871
rect 478 2866 484 2867
rect 622 2871 628 2872
rect 622 2867 623 2871
rect 627 2867 628 2871
rect 622 2866 628 2867
rect 702 2871 708 2872
rect 702 2867 703 2871
rect 707 2867 708 2871
rect 702 2866 708 2867
rect 790 2871 796 2872
rect 790 2867 791 2871
rect 795 2867 796 2871
rect 790 2866 796 2867
rect 802 2871 808 2872
rect 802 2867 803 2871
rect 807 2867 808 2871
rect 802 2866 808 2867
rect 286 2863 292 2864
rect 286 2859 287 2863
rect 291 2859 292 2863
rect 336 2859 338 2866
rect 472 2859 474 2866
rect 111 2858 115 2859
rect 255 2858 259 2859
rect 286 2858 292 2859
rect 335 2858 339 2859
rect 111 2853 115 2854
rect 254 2853 260 2854
rect 112 2850 114 2853
rect 110 2849 116 2850
rect 110 2845 111 2849
rect 115 2845 116 2849
rect 254 2849 255 2853
rect 259 2849 260 2853
rect 254 2848 260 2849
rect 288 2848 290 2858
rect 415 2858 419 2859
rect 471 2858 475 2859
rect 335 2853 339 2854
rect 414 2853 420 2854
rect 471 2853 475 2854
rect 414 2849 415 2853
rect 419 2849 420 2853
rect 414 2848 420 2849
rect 480 2848 482 2866
rect 624 2859 626 2866
rect 559 2858 563 2859
rect 623 2858 627 2859
rect 695 2858 699 2859
rect 558 2853 564 2854
rect 623 2853 627 2854
rect 694 2853 700 2854
rect 558 2849 559 2853
rect 563 2849 564 2853
rect 558 2848 564 2849
rect 694 2849 695 2853
rect 699 2849 700 2853
rect 694 2848 700 2849
rect 704 2848 706 2866
rect 792 2859 794 2866
rect 791 2858 795 2859
rect 791 2853 795 2854
rect 804 2848 806 2866
rect 823 2858 827 2859
rect 822 2853 828 2854
rect 822 2849 823 2853
rect 827 2849 828 2853
rect 822 2848 828 2849
rect 936 2848 938 2930
rect 1094 2912 1100 2913
rect 1094 2908 1095 2912
rect 1099 2908 1100 2912
rect 1094 2907 1100 2908
rect 975 2906 979 2907
rect 975 2901 979 2902
rect 1095 2906 1099 2907
rect 1095 2901 1099 2902
rect 974 2900 980 2901
rect 974 2896 975 2900
rect 979 2896 980 2900
rect 974 2895 980 2896
rect 974 2871 980 2872
rect 974 2867 975 2871
rect 979 2867 980 2871
rect 974 2866 980 2867
rect 982 2871 988 2872
rect 982 2867 983 2871
rect 987 2867 988 2871
rect 982 2866 988 2867
rect 976 2859 978 2866
rect 951 2858 955 2859
rect 975 2858 979 2859
rect 950 2853 956 2854
rect 975 2853 979 2854
rect 950 2849 951 2853
rect 955 2849 956 2853
rect 950 2848 956 2849
rect 984 2848 986 2866
rect 1104 2864 1106 2930
rect 1262 2912 1268 2913
rect 1262 2908 1263 2912
rect 1267 2908 1268 2912
rect 1262 2907 1268 2908
rect 1175 2906 1179 2907
rect 1175 2901 1179 2902
rect 1263 2906 1267 2907
rect 1263 2901 1267 2902
rect 1174 2900 1180 2901
rect 1174 2896 1175 2900
rect 1179 2896 1180 2900
rect 1174 2895 1180 2896
rect 1174 2871 1180 2872
rect 1174 2867 1175 2871
rect 1179 2867 1180 2871
rect 1174 2866 1180 2867
rect 1094 2863 1100 2864
rect 1094 2859 1095 2863
rect 1099 2859 1100 2863
rect 1087 2858 1091 2859
rect 1094 2858 1100 2859
rect 1102 2863 1108 2864
rect 1102 2859 1103 2863
rect 1107 2859 1108 2863
rect 1176 2859 1178 2866
rect 1344 2864 1346 2930
rect 1610 2927 1611 2931
rect 1615 2927 1616 2931
rect 1610 2926 1616 2927
rect 1438 2912 1444 2913
rect 1438 2908 1439 2912
rect 1443 2908 1444 2912
rect 1438 2907 1444 2908
rect 1598 2912 1604 2913
rect 1598 2908 1599 2912
rect 1603 2908 1604 2912
rect 1598 2907 1604 2908
rect 1383 2906 1387 2907
rect 1383 2901 1387 2902
rect 1439 2906 1443 2907
rect 1439 2901 1443 2902
rect 1591 2906 1595 2907
rect 1591 2901 1595 2902
rect 1599 2906 1603 2907
rect 1599 2901 1603 2902
rect 1382 2900 1388 2901
rect 1382 2896 1383 2900
rect 1387 2896 1388 2900
rect 1382 2895 1388 2896
rect 1590 2900 1596 2901
rect 1590 2896 1591 2900
rect 1595 2896 1596 2900
rect 1590 2895 1596 2896
rect 1612 2876 1614 2926
rect 1670 2923 1676 2924
rect 1630 2919 1636 2920
rect 1630 2915 1631 2919
rect 1635 2915 1636 2919
rect 1670 2919 1671 2923
rect 1675 2919 1676 2923
rect 1670 2918 1676 2919
rect 1630 2914 1636 2915
rect 1632 2907 1634 2914
rect 1672 2911 1674 2918
rect 1694 2916 1700 2917
rect 1694 2912 1695 2916
rect 1699 2912 1700 2916
rect 1694 2911 1700 2912
rect 1934 2916 1940 2917
rect 1934 2912 1935 2916
rect 1939 2912 1940 2916
rect 1934 2911 1940 2912
rect 2222 2916 2228 2917
rect 2222 2912 2223 2916
rect 2227 2912 2228 2916
rect 2222 2911 2228 2912
rect 1671 2910 1675 2911
rect 1631 2906 1635 2907
rect 1671 2905 1675 2906
rect 1695 2910 1699 2911
rect 1695 2905 1699 2906
rect 1935 2910 1939 2911
rect 1935 2905 1939 2906
rect 2223 2910 2227 2911
rect 2223 2905 2227 2906
rect 1631 2901 1635 2902
rect 1632 2894 1634 2901
rect 1672 2898 1674 2905
rect 1670 2897 1676 2898
rect 1630 2893 1636 2894
rect 1630 2889 1631 2893
rect 1635 2889 1636 2893
rect 1670 2893 1671 2897
rect 1675 2893 1676 2897
rect 1670 2892 1676 2893
rect 1630 2888 1636 2889
rect 1670 2879 1676 2880
rect 1610 2875 1616 2876
rect 1382 2871 1388 2872
rect 1382 2867 1383 2871
rect 1387 2867 1388 2871
rect 1382 2866 1388 2867
rect 1590 2871 1596 2872
rect 1590 2867 1591 2871
rect 1595 2867 1596 2871
rect 1610 2871 1611 2875
rect 1615 2871 1616 2875
rect 1610 2870 1616 2871
rect 1630 2875 1636 2876
rect 1630 2871 1631 2875
rect 1635 2871 1636 2875
rect 1670 2875 1671 2879
rect 1675 2875 1676 2879
rect 1670 2874 1676 2875
rect 1672 2871 1674 2874
rect 1630 2870 1636 2871
rect 1671 2870 1675 2871
rect 1590 2866 1596 2867
rect 1342 2863 1348 2864
rect 1342 2859 1343 2863
rect 1347 2859 1348 2863
rect 1384 2859 1386 2866
rect 1592 2859 1594 2866
rect 1102 2858 1108 2859
rect 1175 2858 1179 2859
rect 1342 2858 1348 2859
rect 1383 2858 1387 2859
rect 1086 2853 1092 2854
rect 1086 2849 1087 2853
rect 1091 2849 1092 2853
rect 1086 2848 1092 2849
rect 1096 2848 1098 2858
rect 1175 2853 1179 2854
rect 110 2844 116 2845
rect 286 2847 292 2848
rect 286 2843 287 2847
rect 291 2843 292 2847
rect 286 2842 292 2843
rect 422 2847 428 2848
rect 422 2843 423 2847
rect 427 2843 428 2847
rect 422 2842 428 2843
rect 478 2847 484 2848
rect 478 2843 479 2847
rect 483 2843 484 2847
rect 478 2842 484 2843
rect 702 2847 708 2848
rect 702 2843 703 2847
rect 707 2843 708 2847
rect 702 2842 708 2843
rect 802 2847 808 2848
rect 802 2843 803 2847
rect 807 2843 808 2847
rect 802 2842 808 2843
rect 870 2847 876 2848
rect 870 2843 871 2847
rect 875 2843 876 2847
rect 870 2842 876 2843
rect 934 2847 940 2848
rect 934 2843 935 2847
rect 939 2843 940 2847
rect 934 2842 940 2843
rect 982 2847 988 2848
rect 982 2843 983 2847
rect 987 2843 988 2847
rect 982 2842 988 2843
rect 1094 2847 1100 2848
rect 1094 2843 1095 2847
rect 1099 2843 1100 2847
rect 1094 2842 1100 2843
rect 110 2831 116 2832
rect 110 2827 111 2831
rect 115 2827 116 2831
rect 110 2826 116 2827
rect 112 2811 114 2826
rect 254 2824 260 2825
rect 254 2820 255 2824
rect 259 2820 260 2824
rect 254 2819 260 2820
rect 256 2811 258 2819
rect 111 2810 115 2811
rect 111 2805 115 2806
rect 151 2810 155 2811
rect 151 2805 155 2806
rect 255 2810 259 2811
rect 255 2805 259 2806
rect 279 2810 283 2811
rect 279 2805 283 2806
rect 112 2798 114 2805
rect 150 2804 156 2805
rect 150 2800 151 2804
rect 155 2800 156 2804
rect 150 2799 156 2800
rect 278 2804 284 2805
rect 278 2800 279 2804
rect 283 2800 284 2804
rect 278 2799 284 2800
rect 110 2797 116 2798
rect 110 2793 111 2797
rect 115 2793 116 2797
rect 110 2792 116 2793
rect 288 2784 290 2842
rect 414 2824 420 2825
rect 414 2820 415 2824
rect 419 2820 420 2824
rect 414 2819 420 2820
rect 416 2811 418 2819
rect 399 2810 403 2811
rect 399 2805 403 2806
rect 415 2810 419 2811
rect 415 2805 419 2806
rect 398 2804 404 2805
rect 398 2800 399 2804
rect 403 2800 404 2804
rect 398 2799 404 2800
rect 424 2784 426 2842
rect 558 2824 564 2825
rect 558 2820 559 2824
rect 563 2820 564 2824
rect 558 2819 564 2820
rect 694 2824 700 2825
rect 694 2820 695 2824
rect 699 2820 700 2824
rect 694 2819 700 2820
rect 560 2811 562 2819
rect 696 2811 698 2819
rect 519 2810 523 2811
rect 519 2805 523 2806
rect 559 2810 563 2811
rect 559 2805 563 2806
rect 639 2810 643 2811
rect 639 2805 643 2806
rect 695 2810 699 2811
rect 695 2805 699 2806
rect 518 2804 524 2805
rect 518 2800 519 2804
rect 523 2800 524 2804
rect 518 2799 524 2800
rect 638 2804 644 2805
rect 638 2800 639 2804
rect 643 2800 644 2804
rect 638 2799 644 2800
rect 704 2784 706 2842
rect 822 2824 828 2825
rect 822 2820 823 2824
rect 827 2820 828 2824
rect 822 2819 828 2820
rect 824 2811 826 2819
rect 751 2810 755 2811
rect 751 2805 755 2806
rect 823 2810 827 2811
rect 823 2805 827 2806
rect 863 2810 867 2811
rect 863 2805 867 2806
rect 750 2804 756 2805
rect 750 2800 751 2804
rect 755 2800 756 2804
rect 750 2799 756 2800
rect 862 2804 868 2805
rect 862 2800 863 2804
rect 867 2800 868 2804
rect 862 2799 868 2800
rect 286 2783 292 2784
rect 110 2779 116 2780
rect 110 2775 111 2779
rect 115 2775 116 2779
rect 286 2779 287 2783
rect 291 2779 292 2783
rect 286 2778 292 2779
rect 422 2783 428 2784
rect 422 2779 423 2783
rect 427 2779 428 2783
rect 422 2778 428 2779
rect 630 2783 636 2784
rect 630 2779 631 2783
rect 635 2779 636 2783
rect 630 2778 636 2779
rect 702 2783 708 2784
rect 702 2779 703 2783
rect 707 2779 708 2783
rect 872 2780 874 2842
rect 1096 2833 1098 2842
rect 1096 2831 1106 2833
rect 950 2824 956 2825
rect 950 2820 951 2824
rect 955 2820 956 2824
rect 950 2819 956 2820
rect 1086 2824 1092 2825
rect 1086 2820 1087 2824
rect 1091 2820 1092 2824
rect 1086 2819 1092 2820
rect 952 2811 954 2819
rect 1088 2811 1090 2819
rect 951 2810 955 2811
rect 951 2805 955 2806
rect 983 2810 987 2811
rect 983 2805 987 2806
rect 1087 2810 1091 2811
rect 1087 2805 1091 2806
rect 982 2804 988 2805
rect 982 2800 983 2804
rect 987 2800 988 2804
rect 982 2799 988 2800
rect 702 2778 708 2779
rect 870 2779 876 2780
rect 288 2776 290 2778
rect 110 2774 116 2775
rect 150 2775 156 2776
rect 112 2759 114 2774
rect 150 2771 151 2775
rect 155 2771 156 2775
rect 150 2770 156 2771
rect 158 2775 164 2776
rect 158 2771 159 2775
rect 163 2771 164 2775
rect 158 2770 164 2771
rect 278 2775 284 2776
rect 278 2771 279 2775
rect 283 2771 284 2775
rect 278 2770 284 2771
rect 286 2775 292 2776
rect 286 2771 287 2775
rect 291 2771 292 2775
rect 286 2770 292 2771
rect 398 2775 404 2776
rect 398 2771 399 2775
rect 403 2771 404 2775
rect 398 2770 404 2771
rect 152 2759 154 2770
rect 111 2758 115 2759
rect 135 2758 139 2759
rect 151 2758 155 2759
rect 111 2753 115 2754
rect 134 2753 140 2754
rect 151 2753 155 2754
rect 112 2750 114 2753
rect 110 2749 116 2750
rect 110 2745 111 2749
rect 115 2745 116 2749
rect 134 2749 135 2753
rect 139 2749 140 2753
rect 160 2752 162 2770
rect 280 2759 282 2770
rect 263 2758 267 2759
rect 279 2758 283 2759
rect 262 2753 268 2754
rect 279 2753 283 2754
rect 134 2748 140 2749
rect 158 2751 164 2752
rect 158 2747 159 2751
rect 163 2747 164 2751
rect 262 2749 263 2753
rect 267 2749 268 2753
rect 262 2748 268 2749
rect 288 2748 290 2770
rect 400 2759 402 2770
rect 399 2758 403 2759
rect 399 2753 403 2754
rect 424 2748 426 2778
rect 518 2775 524 2776
rect 518 2771 519 2775
rect 523 2771 524 2775
rect 518 2770 524 2771
rect 520 2759 522 2770
rect 431 2758 435 2759
rect 519 2758 523 2759
rect 623 2758 627 2759
rect 430 2753 436 2754
rect 519 2753 523 2754
rect 622 2753 628 2754
rect 430 2749 431 2753
rect 435 2749 436 2753
rect 430 2748 436 2749
rect 622 2749 623 2753
rect 627 2749 628 2753
rect 632 2752 634 2778
rect 638 2775 644 2776
rect 638 2771 639 2775
rect 643 2771 644 2775
rect 638 2770 644 2771
rect 750 2775 756 2776
rect 750 2771 751 2775
rect 755 2771 756 2775
rect 750 2770 756 2771
rect 862 2775 868 2776
rect 862 2771 863 2775
rect 867 2771 868 2775
rect 870 2775 871 2779
rect 875 2775 876 2779
rect 870 2774 876 2775
rect 966 2779 972 2780
rect 966 2775 967 2779
rect 971 2775 972 2779
rect 966 2774 972 2775
rect 982 2775 988 2776
rect 862 2770 868 2771
rect 640 2759 642 2770
rect 752 2759 754 2770
rect 864 2759 866 2770
rect 639 2758 643 2759
rect 639 2753 643 2754
rect 751 2758 755 2759
rect 839 2758 843 2759
rect 863 2758 867 2759
rect 751 2753 755 2754
rect 838 2753 844 2754
rect 863 2753 867 2754
rect 622 2748 628 2749
rect 630 2751 636 2752
rect 158 2746 164 2747
rect 286 2747 292 2748
rect 110 2744 116 2745
rect 286 2743 287 2747
rect 291 2743 292 2747
rect 286 2742 292 2743
rect 422 2747 428 2748
rect 422 2743 423 2747
rect 427 2743 428 2747
rect 630 2747 631 2751
rect 635 2747 636 2751
rect 838 2749 839 2753
rect 843 2749 844 2753
rect 872 2752 874 2774
rect 838 2748 844 2749
rect 870 2751 876 2752
rect 630 2746 636 2747
rect 870 2747 871 2751
rect 875 2747 876 2751
rect 870 2746 876 2747
rect 422 2742 428 2743
rect 110 2731 116 2732
rect 110 2727 111 2731
rect 115 2727 116 2731
rect 110 2726 116 2727
rect 112 2707 114 2726
rect 134 2724 140 2725
rect 134 2720 135 2724
rect 139 2720 140 2724
rect 134 2719 140 2720
rect 262 2724 268 2725
rect 262 2720 263 2724
rect 267 2720 268 2724
rect 262 2719 268 2720
rect 430 2724 436 2725
rect 430 2720 431 2724
rect 435 2720 436 2724
rect 430 2719 436 2720
rect 622 2724 628 2725
rect 622 2720 623 2724
rect 627 2720 628 2724
rect 622 2719 628 2720
rect 136 2707 138 2719
rect 264 2707 266 2719
rect 432 2707 434 2719
rect 624 2707 626 2719
rect 111 2706 115 2707
rect 111 2701 115 2702
rect 135 2706 139 2707
rect 135 2701 139 2702
rect 263 2706 267 2707
rect 263 2701 267 2702
rect 431 2706 435 2707
rect 431 2701 435 2702
rect 623 2706 627 2707
rect 623 2701 627 2702
rect 112 2694 114 2701
rect 110 2693 116 2694
rect 110 2689 111 2693
rect 115 2689 116 2693
rect 110 2688 116 2689
rect 632 2680 634 2746
rect 838 2724 844 2725
rect 838 2720 839 2724
rect 843 2720 844 2724
rect 838 2719 844 2720
rect 840 2707 842 2719
rect 703 2706 707 2707
rect 703 2701 707 2702
rect 831 2706 835 2707
rect 831 2701 835 2702
rect 839 2706 843 2707
rect 839 2701 843 2702
rect 959 2706 963 2707
rect 959 2701 963 2702
rect 702 2700 708 2701
rect 702 2696 703 2700
rect 707 2696 708 2700
rect 702 2695 708 2696
rect 830 2700 836 2701
rect 830 2696 831 2700
rect 835 2696 836 2700
rect 830 2695 836 2696
rect 958 2700 964 2701
rect 958 2696 959 2700
rect 963 2696 964 2700
rect 958 2695 964 2696
rect 630 2679 636 2680
rect 110 2675 116 2676
rect 110 2671 111 2675
rect 115 2671 116 2675
rect 630 2675 631 2679
rect 635 2675 636 2679
rect 968 2676 970 2774
rect 982 2771 983 2775
rect 987 2771 988 2775
rect 982 2770 988 2771
rect 984 2759 986 2770
rect 983 2758 987 2759
rect 1071 2758 1075 2759
rect 983 2753 987 2754
rect 1070 2753 1076 2754
rect 1070 2749 1071 2753
rect 1075 2749 1076 2753
rect 1070 2748 1076 2749
rect 1104 2748 1106 2831
rect 1319 2758 1323 2759
rect 1318 2753 1324 2754
rect 1318 2749 1319 2753
rect 1323 2749 1324 2753
rect 1318 2748 1324 2749
rect 1344 2748 1346 2858
rect 1383 2853 1387 2854
rect 1591 2858 1595 2859
rect 1591 2853 1595 2854
rect 1567 2758 1571 2759
rect 1566 2753 1572 2754
rect 1566 2749 1567 2753
rect 1571 2749 1572 2753
rect 1612 2752 1614 2870
rect 1632 2859 1634 2870
rect 2207 2870 2211 2871
rect 1671 2865 1675 2866
rect 2206 2865 2212 2866
rect 1672 2862 1674 2865
rect 1670 2861 1676 2862
rect 1631 2858 1635 2859
rect 1670 2857 1671 2861
rect 1675 2857 1676 2861
rect 2206 2861 2207 2865
rect 2211 2861 2212 2865
rect 2206 2860 2212 2861
rect 1670 2856 1676 2857
rect 1631 2853 1635 2854
rect 1632 2850 1634 2853
rect 1630 2849 1636 2850
rect 1630 2845 1631 2849
rect 1635 2845 1636 2849
rect 1630 2844 1636 2845
rect 1670 2843 1676 2844
rect 1670 2839 1671 2843
rect 1675 2839 1676 2843
rect 1670 2838 1676 2839
rect 1630 2831 1636 2832
rect 1630 2827 1631 2831
rect 1635 2827 1636 2831
rect 1630 2826 1636 2827
rect 1632 2811 1634 2826
rect 1672 2823 1674 2838
rect 2206 2836 2212 2837
rect 2206 2832 2207 2836
rect 2211 2832 2212 2836
rect 2206 2831 2212 2832
rect 2208 2823 2210 2831
rect 1671 2822 1675 2823
rect 1671 2817 1675 2818
rect 2127 2822 2131 2823
rect 2127 2817 2131 2818
rect 2207 2822 2211 2823
rect 2207 2817 2211 2818
rect 1631 2810 1635 2811
rect 1672 2810 1674 2817
rect 2126 2816 2132 2817
rect 2126 2812 2127 2816
rect 2131 2812 2132 2816
rect 2126 2811 2132 2812
rect 1631 2805 1635 2806
rect 1670 2809 1676 2810
rect 1670 2805 1671 2809
rect 1675 2805 1676 2809
rect 1632 2798 1634 2805
rect 1670 2804 1676 2805
rect 1630 2797 1636 2798
rect 1630 2793 1631 2797
rect 1635 2793 1636 2797
rect 1630 2792 1636 2793
rect 1670 2791 1676 2792
rect 1670 2787 1671 2791
rect 1675 2787 1676 2791
rect 1670 2786 1676 2787
rect 2126 2787 2132 2788
rect 1672 2783 1674 2786
rect 2126 2783 2127 2787
rect 2131 2783 2132 2787
rect 1671 2782 1675 2783
rect 1630 2779 1636 2780
rect 1630 2775 1631 2779
rect 1635 2775 1636 2779
rect 2039 2782 2043 2783
rect 2126 2782 2132 2783
rect 2207 2782 2211 2783
rect 1671 2777 1675 2778
rect 2038 2777 2044 2778
rect 2127 2777 2131 2778
rect 2206 2777 2212 2778
rect 1630 2774 1636 2775
rect 1672 2774 1674 2777
rect 1632 2759 1634 2774
rect 1670 2773 1676 2774
rect 1670 2769 1671 2773
rect 1675 2769 1676 2773
rect 2038 2773 2039 2777
rect 2043 2773 2044 2777
rect 2038 2772 2044 2773
rect 2206 2773 2207 2777
rect 2211 2773 2212 2777
rect 2206 2772 2212 2773
rect 2232 2772 2234 2934
rect 2296 2915 2298 2938
rect 2518 2916 2524 2917
rect 2296 2913 2306 2915
rect 2295 2910 2299 2911
rect 2295 2905 2299 2906
rect 2294 2904 2300 2905
rect 2294 2900 2295 2904
rect 2299 2900 2300 2904
rect 2294 2899 2300 2900
rect 2304 2880 2306 2913
rect 2518 2912 2519 2916
rect 2523 2912 2524 2916
rect 2518 2911 2524 2912
rect 2519 2910 2523 2911
rect 2519 2905 2523 2906
rect 2528 2884 2530 2938
rect 2834 2935 2835 2939
rect 2839 2935 2840 2939
rect 3142 2939 3143 2943
rect 3147 2939 3148 2943
rect 3142 2938 3148 2939
rect 3166 2943 3172 2944
rect 3166 2939 3167 2943
rect 3171 2939 3172 2943
rect 3192 2942 3194 2945
rect 3166 2938 3172 2939
rect 3190 2941 3196 2942
rect 2834 2934 2840 2935
rect 2822 2916 2828 2917
rect 2822 2912 2823 2916
rect 2827 2912 2828 2916
rect 2822 2911 2828 2912
rect 2551 2910 2555 2911
rect 2551 2905 2555 2906
rect 2815 2910 2819 2911
rect 2815 2905 2819 2906
rect 2823 2910 2827 2911
rect 2823 2905 2827 2906
rect 2550 2904 2556 2905
rect 2550 2900 2551 2904
rect 2555 2900 2556 2904
rect 2550 2899 2556 2900
rect 2814 2904 2820 2905
rect 2814 2900 2815 2904
rect 2819 2900 2820 2904
rect 2814 2899 2820 2900
rect 2526 2883 2532 2884
rect 2302 2879 2308 2880
rect 2294 2875 2300 2876
rect 2294 2871 2295 2875
rect 2299 2871 2300 2875
rect 2302 2875 2303 2879
rect 2307 2875 2308 2879
rect 2526 2879 2527 2883
rect 2531 2879 2532 2883
rect 2526 2878 2532 2879
rect 2542 2883 2548 2884
rect 2542 2879 2543 2883
rect 2547 2879 2548 2883
rect 2542 2878 2548 2879
rect 2302 2874 2308 2875
rect 2294 2870 2300 2871
rect 2295 2865 2299 2866
rect 2304 2864 2306 2874
rect 2375 2870 2379 2871
rect 2535 2870 2539 2871
rect 2374 2865 2380 2866
rect 2302 2863 2308 2864
rect 2302 2859 2303 2863
rect 2307 2859 2308 2863
rect 2374 2861 2375 2865
rect 2379 2861 2380 2865
rect 2374 2860 2380 2861
rect 2534 2865 2540 2866
rect 2534 2861 2535 2865
rect 2539 2861 2540 2865
rect 2544 2864 2546 2878
rect 2836 2876 2838 2934
rect 3134 2916 3140 2917
rect 3134 2912 3135 2916
rect 3139 2912 3140 2916
rect 3134 2911 3140 2912
rect 3079 2910 3083 2911
rect 3079 2905 3083 2906
rect 3135 2910 3139 2911
rect 3135 2905 3139 2906
rect 3078 2904 3084 2905
rect 3078 2900 3079 2904
rect 3083 2900 3084 2904
rect 3078 2899 3084 2900
rect 2550 2875 2556 2876
rect 2550 2871 2551 2875
rect 2555 2871 2556 2875
rect 2814 2875 2820 2876
rect 2814 2871 2815 2875
rect 2819 2871 2820 2875
rect 2834 2875 2840 2876
rect 2834 2871 2835 2875
rect 2839 2871 2840 2875
rect 3078 2875 3084 2876
rect 3078 2871 3079 2875
rect 3083 2871 3084 2875
rect 2550 2870 2556 2871
rect 2679 2870 2683 2871
rect 2814 2870 2820 2871
rect 2823 2870 2827 2871
rect 2834 2870 2840 2871
rect 2967 2870 2971 2871
rect 3078 2870 3084 2871
rect 3111 2870 3115 2871
rect 2551 2865 2555 2866
rect 2678 2865 2684 2866
rect 2815 2865 2819 2866
rect 2822 2865 2828 2866
rect 2534 2860 2540 2861
rect 2542 2863 2548 2864
rect 2302 2858 2308 2859
rect 2382 2859 2388 2860
rect 2304 2833 2306 2858
rect 2382 2855 2383 2859
rect 2387 2855 2388 2859
rect 2542 2859 2543 2863
rect 2547 2859 2548 2863
rect 2678 2861 2679 2865
rect 2683 2861 2684 2865
rect 2678 2860 2684 2861
rect 2822 2861 2823 2865
rect 2827 2861 2828 2865
rect 2822 2860 2828 2861
rect 2836 2860 2838 2870
rect 2966 2865 2972 2866
rect 3079 2865 3083 2866
rect 3110 2865 3116 2866
rect 2966 2861 2967 2865
rect 2971 2861 2972 2865
rect 2966 2860 2972 2861
rect 3110 2861 3111 2865
rect 3115 2861 3116 2865
rect 3144 2864 3146 2938
rect 3190 2937 3191 2941
rect 3195 2937 3196 2941
rect 3190 2936 3196 2937
rect 3190 2923 3196 2924
rect 3190 2919 3191 2923
rect 3195 2919 3196 2923
rect 3190 2918 3196 2919
rect 3192 2911 3194 2918
rect 3191 2910 3195 2911
rect 3191 2905 3195 2906
rect 3192 2898 3194 2905
rect 3190 2897 3196 2898
rect 3190 2893 3191 2897
rect 3195 2893 3196 2897
rect 3190 2892 3196 2893
rect 3190 2879 3196 2880
rect 3190 2875 3191 2879
rect 3195 2875 3196 2879
rect 3190 2874 3196 2875
rect 3192 2871 3194 2874
rect 3191 2870 3195 2871
rect 3191 2865 3195 2866
rect 3110 2860 3116 2861
rect 3142 2863 3148 2864
rect 2542 2858 2548 2859
rect 2686 2859 2692 2860
rect 2382 2854 2388 2855
rect 2686 2855 2687 2859
rect 2691 2855 2692 2859
rect 2686 2854 2692 2855
rect 2834 2859 2840 2860
rect 2834 2855 2835 2859
rect 2839 2855 2840 2859
rect 2834 2854 2840 2855
rect 2974 2859 2980 2860
rect 2974 2855 2975 2859
rect 2979 2855 2980 2859
rect 3142 2859 3143 2863
rect 3147 2859 3148 2863
rect 3142 2858 3148 2859
rect 3166 2863 3172 2864
rect 3166 2859 3167 2863
rect 3171 2859 3172 2863
rect 3192 2862 3194 2865
rect 3166 2858 3172 2859
rect 3190 2861 3196 2862
rect 2974 2854 2980 2855
rect 2374 2836 2380 2837
rect 2304 2831 2314 2833
rect 2374 2832 2375 2836
rect 2379 2832 2380 2836
rect 2374 2831 2380 2832
rect 2303 2822 2307 2823
rect 2303 2817 2307 2818
rect 2302 2816 2308 2817
rect 2302 2812 2303 2816
rect 2307 2812 2308 2816
rect 2302 2811 2308 2812
rect 2312 2792 2314 2831
rect 2376 2823 2378 2831
rect 2375 2822 2379 2823
rect 2375 2817 2379 2818
rect 2384 2792 2386 2854
rect 2534 2836 2540 2837
rect 2534 2832 2535 2836
rect 2539 2832 2540 2836
rect 2534 2831 2540 2832
rect 2678 2836 2684 2837
rect 2678 2832 2679 2836
rect 2683 2832 2684 2836
rect 2678 2831 2684 2832
rect 2536 2823 2538 2831
rect 2680 2823 2682 2831
rect 2479 2822 2483 2823
rect 2479 2817 2483 2818
rect 2535 2822 2539 2823
rect 2535 2817 2539 2818
rect 2655 2822 2659 2823
rect 2655 2817 2659 2818
rect 2679 2822 2683 2823
rect 2679 2817 2683 2818
rect 2478 2816 2484 2817
rect 2478 2812 2479 2816
rect 2483 2812 2484 2816
rect 2478 2811 2484 2812
rect 2654 2816 2660 2817
rect 2654 2812 2655 2816
rect 2659 2812 2660 2816
rect 2654 2811 2660 2812
rect 2310 2791 2316 2792
rect 2302 2787 2308 2788
rect 2302 2783 2303 2787
rect 2307 2783 2308 2787
rect 2310 2787 2311 2791
rect 2315 2787 2316 2791
rect 2310 2786 2316 2787
rect 2350 2791 2356 2792
rect 2350 2787 2351 2791
rect 2355 2787 2356 2791
rect 2350 2786 2356 2787
rect 2382 2791 2388 2792
rect 2382 2787 2383 2791
rect 2387 2787 2388 2791
rect 2688 2788 2690 2854
rect 2836 2851 2838 2854
rect 2836 2849 2842 2851
rect 2822 2836 2828 2837
rect 2822 2832 2823 2836
rect 2827 2832 2828 2836
rect 2822 2831 2828 2832
rect 2824 2823 2826 2831
rect 2823 2822 2827 2823
rect 2823 2817 2827 2818
rect 2831 2822 2835 2823
rect 2831 2817 2835 2818
rect 2830 2816 2836 2817
rect 2830 2812 2831 2816
rect 2835 2812 2836 2816
rect 2830 2811 2836 2812
rect 2840 2788 2842 2849
rect 2966 2836 2972 2837
rect 2966 2832 2967 2836
rect 2971 2832 2972 2836
rect 2966 2831 2972 2832
rect 2968 2823 2970 2831
rect 2967 2822 2971 2823
rect 2967 2817 2971 2818
rect 2976 2796 2978 2854
rect 3110 2836 3116 2837
rect 3110 2832 3111 2836
rect 3115 2832 3116 2836
rect 3110 2831 3116 2832
rect 3112 2823 3114 2831
rect 3007 2822 3011 2823
rect 3007 2817 3011 2818
rect 3111 2822 3115 2823
rect 3111 2817 3115 2818
rect 3159 2822 3163 2823
rect 3159 2817 3163 2818
rect 3006 2816 3012 2817
rect 3006 2812 3007 2816
rect 3011 2812 3012 2816
rect 3006 2811 3012 2812
rect 3158 2816 3164 2817
rect 3158 2812 3159 2816
rect 3163 2812 3164 2816
rect 3158 2811 3164 2812
rect 2974 2795 2980 2796
rect 2974 2791 2975 2795
rect 2979 2791 2980 2795
rect 2974 2790 2980 2791
rect 3168 2788 3170 2858
rect 3190 2857 3191 2861
rect 3195 2857 3196 2861
rect 3190 2856 3196 2857
rect 3190 2843 3196 2844
rect 3190 2839 3191 2843
rect 3195 2839 3196 2843
rect 3190 2838 3196 2839
rect 3192 2823 3194 2838
rect 3191 2822 3195 2823
rect 3191 2817 3195 2818
rect 3192 2810 3194 2817
rect 3190 2809 3196 2810
rect 3190 2805 3191 2809
rect 3195 2805 3196 2809
rect 3190 2804 3196 2805
rect 3190 2791 3196 2792
rect 2382 2786 2388 2787
rect 2478 2787 2484 2788
rect 2302 2782 2308 2783
rect 2303 2777 2307 2778
rect 1670 2768 1676 2769
rect 2022 2771 2028 2772
rect 2022 2767 2023 2771
rect 2027 2767 2028 2771
rect 2022 2766 2028 2767
rect 2230 2771 2236 2772
rect 2230 2767 2231 2771
rect 2235 2767 2236 2771
rect 2230 2766 2236 2767
rect 1631 2758 1635 2759
rect 1631 2753 1635 2754
rect 1670 2755 1676 2756
rect 1566 2748 1572 2749
rect 1574 2751 1580 2752
rect 1102 2747 1108 2748
rect 1102 2743 1103 2747
rect 1107 2743 1108 2747
rect 1102 2742 1108 2743
rect 1342 2747 1348 2748
rect 1342 2743 1343 2747
rect 1347 2743 1348 2747
rect 1574 2747 1575 2751
rect 1579 2747 1580 2751
rect 1574 2746 1580 2747
rect 1610 2751 1616 2752
rect 1610 2747 1611 2751
rect 1615 2747 1616 2751
rect 1632 2750 1634 2753
rect 1670 2751 1671 2755
rect 1675 2751 1676 2755
rect 1670 2750 1676 2751
rect 1610 2746 1616 2747
rect 1630 2749 1636 2750
rect 1342 2742 1348 2743
rect 1070 2724 1076 2725
rect 1070 2720 1071 2724
rect 1075 2720 1076 2724
rect 1070 2719 1076 2720
rect 1072 2707 1074 2719
rect 1071 2706 1075 2707
rect 1071 2701 1075 2702
rect 1079 2706 1083 2707
rect 1079 2701 1083 2702
rect 1078 2700 1084 2701
rect 1078 2696 1079 2700
rect 1083 2696 1084 2700
rect 1078 2695 1084 2696
rect 630 2674 636 2675
rect 742 2675 748 2676
rect 110 2670 116 2671
rect 112 2659 114 2670
rect 111 2658 115 2659
rect 607 2658 611 2659
rect 111 2653 115 2654
rect 606 2653 612 2654
rect 112 2650 114 2653
rect 110 2649 116 2650
rect 110 2645 111 2649
rect 115 2645 116 2649
rect 606 2649 607 2653
rect 611 2649 612 2653
rect 632 2652 634 2674
rect 702 2671 708 2672
rect 702 2667 703 2671
rect 707 2667 708 2671
rect 742 2671 743 2675
rect 747 2671 748 2675
rect 966 2675 972 2676
rect 742 2670 748 2671
rect 830 2671 836 2672
rect 702 2666 708 2667
rect 704 2659 706 2666
rect 703 2658 707 2659
rect 735 2658 739 2659
rect 703 2653 707 2654
rect 734 2653 740 2654
rect 606 2648 612 2649
rect 630 2651 636 2652
rect 630 2647 631 2651
rect 635 2647 636 2651
rect 734 2649 735 2653
rect 739 2649 740 2653
rect 744 2652 746 2670
rect 830 2667 831 2671
rect 835 2667 836 2671
rect 830 2666 836 2667
rect 862 2671 868 2672
rect 862 2667 863 2671
rect 867 2667 868 2671
rect 862 2666 868 2667
rect 958 2671 964 2672
rect 958 2667 959 2671
rect 963 2667 964 2671
rect 966 2671 967 2675
rect 971 2671 972 2675
rect 1104 2672 1106 2742
rect 1318 2724 1324 2725
rect 1318 2720 1319 2724
rect 1323 2720 1324 2724
rect 1318 2719 1324 2720
rect 1320 2707 1322 2719
rect 1199 2706 1203 2707
rect 1199 2701 1203 2702
rect 1311 2706 1315 2707
rect 1311 2701 1315 2702
rect 1319 2706 1323 2707
rect 1319 2701 1323 2702
rect 1198 2700 1204 2701
rect 1198 2696 1199 2700
rect 1203 2696 1204 2700
rect 1198 2695 1204 2696
rect 1310 2700 1316 2701
rect 1310 2696 1311 2700
rect 1315 2696 1316 2700
rect 1310 2695 1316 2696
rect 1344 2680 1346 2742
rect 1566 2724 1572 2725
rect 1566 2720 1567 2724
rect 1571 2720 1572 2724
rect 1566 2719 1572 2720
rect 1568 2707 1570 2719
rect 1423 2706 1427 2707
rect 1423 2701 1427 2702
rect 1543 2706 1547 2707
rect 1543 2701 1547 2702
rect 1567 2706 1571 2707
rect 1567 2701 1571 2702
rect 1422 2700 1428 2701
rect 1422 2696 1423 2700
rect 1427 2696 1428 2700
rect 1422 2695 1428 2696
rect 1542 2700 1548 2701
rect 1542 2696 1543 2700
rect 1547 2696 1548 2700
rect 1542 2695 1548 2696
rect 1342 2679 1348 2680
rect 1342 2675 1343 2679
rect 1347 2675 1348 2679
rect 1342 2674 1348 2675
rect 1446 2679 1452 2680
rect 1446 2675 1447 2679
rect 1451 2675 1452 2679
rect 1576 2676 1578 2746
rect 1630 2745 1631 2749
rect 1635 2745 1636 2749
rect 1630 2744 1636 2745
rect 1672 2739 1674 2750
rect 1671 2738 1675 2739
rect 1671 2733 1675 2734
rect 2015 2738 2019 2739
rect 2015 2733 2019 2734
rect 1630 2731 1636 2732
rect 1630 2727 1631 2731
rect 1635 2727 1636 2731
rect 1630 2726 1636 2727
rect 1672 2726 1674 2733
rect 2014 2732 2020 2733
rect 2014 2728 2015 2732
rect 2019 2728 2020 2732
rect 2014 2727 2020 2728
rect 1632 2707 1634 2726
rect 1670 2725 1676 2726
rect 1670 2721 1671 2725
rect 1675 2721 1676 2725
rect 1670 2720 1676 2721
rect 1670 2707 1676 2708
rect 1631 2706 1635 2707
rect 1670 2703 1671 2707
rect 1675 2703 1676 2707
rect 2024 2704 2026 2766
rect 2038 2748 2044 2749
rect 2038 2744 2039 2748
rect 2043 2744 2044 2748
rect 2038 2743 2044 2744
rect 2206 2748 2212 2749
rect 2206 2744 2207 2748
rect 2211 2744 2212 2748
rect 2206 2743 2212 2744
rect 2040 2739 2042 2743
rect 2208 2739 2210 2743
rect 2039 2738 2043 2739
rect 2039 2733 2043 2734
rect 2199 2738 2203 2739
rect 2199 2733 2203 2734
rect 2207 2738 2211 2739
rect 2207 2733 2211 2734
rect 2198 2732 2204 2733
rect 2198 2728 2199 2732
rect 2203 2728 2204 2732
rect 2198 2727 2204 2728
rect 1670 2702 1676 2703
rect 2014 2703 2020 2704
rect 1631 2701 1635 2702
rect 1632 2694 1634 2701
rect 1630 2693 1636 2694
rect 1630 2689 1631 2693
rect 1635 2689 1636 2693
rect 1672 2691 1674 2702
rect 2014 2699 2015 2703
rect 2019 2699 2020 2703
rect 2014 2698 2020 2699
rect 2022 2703 2028 2704
rect 2022 2699 2023 2703
rect 2027 2699 2028 2703
rect 2022 2698 2028 2699
rect 2198 2703 2204 2704
rect 2198 2699 2199 2703
rect 2203 2699 2204 2703
rect 2198 2698 2204 2699
rect 2206 2703 2212 2704
rect 2206 2699 2207 2703
rect 2211 2699 2212 2703
rect 2206 2698 2212 2699
rect 2016 2691 2018 2698
rect 1630 2688 1636 2689
rect 1671 2690 1675 2691
rect 1999 2690 2003 2691
rect 2015 2690 2019 2691
rect 1671 2685 1675 2686
rect 1998 2685 2004 2686
rect 2015 2685 2019 2686
rect 1672 2682 1674 2685
rect 1670 2681 1676 2682
rect 1670 2677 1671 2681
rect 1675 2677 1676 2681
rect 1998 2681 1999 2685
rect 2003 2681 2004 2685
rect 1998 2680 2004 2681
rect 2024 2680 2026 2698
rect 2200 2691 2202 2698
rect 2175 2690 2179 2691
rect 2199 2690 2203 2691
rect 2174 2685 2180 2686
rect 2199 2685 2203 2686
rect 2174 2681 2175 2685
rect 2179 2681 2180 2685
rect 2174 2680 2180 2681
rect 2208 2680 2210 2698
rect 2352 2680 2354 2786
rect 2375 2782 2379 2783
rect 2374 2777 2380 2778
rect 2374 2773 2375 2777
rect 2379 2773 2380 2777
rect 2384 2776 2386 2786
rect 2478 2783 2479 2787
rect 2483 2783 2484 2787
rect 2654 2787 2660 2788
rect 2654 2783 2655 2787
rect 2659 2783 2660 2787
rect 2478 2782 2484 2783
rect 2535 2782 2539 2783
rect 2654 2782 2660 2783
rect 2686 2787 2692 2788
rect 2686 2783 2687 2787
rect 2691 2783 2692 2787
rect 2830 2787 2836 2788
rect 2830 2783 2831 2787
rect 2835 2783 2836 2787
rect 2686 2782 2692 2783
rect 2703 2782 2707 2783
rect 2830 2782 2836 2783
rect 2838 2787 2844 2788
rect 2838 2783 2839 2787
rect 2843 2783 2844 2787
rect 3006 2787 3012 2788
rect 3006 2783 3007 2787
rect 3011 2783 3012 2787
rect 2838 2782 2844 2783
rect 2871 2782 2875 2783
rect 3006 2782 3012 2783
rect 3014 2787 3020 2788
rect 3014 2783 3015 2787
rect 3019 2783 3020 2787
rect 3014 2782 3020 2783
rect 3158 2787 3164 2788
rect 3158 2783 3159 2787
rect 3163 2783 3164 2787
rect 3158 2782 3164 2783
rect 3166 2787 3172 2788
rect 3166 2783 3167 2787
rect 3171 2783 3172 2787
rect 3190 2787 3191 2791
rect 3195 2787 3196 2791
rect 3190 2786 3196 2787
rect 3192 2783 3194 2786
rect 3166 2782 3172 2783
rect 3191 2782 3195 2783
rect 2479 2777 2483 2778
rect 2534 2777 2540 2778
rect 2655 2777 2659 2778
rect 2702 2777 2708 2778
rect 2831 2777 2835 2778
rect 2374 2772 2380 2773
rect 2382 2775 2388 2776
rect 2382 2771 2383 2775
rect 2387 2771 2388 2775
rect 2534 2773 2535 2777
rect 2539 2773 2540 2777
rect 2534 2772 2540 2773
rect 2558 2775 2564 2776
rect 2382 2770 2388 2771
rect 2558 2771 2559 2775
rect 2563 2771 2564 2775
rect 2702 2773 2703 2777
rect 2707 2773 2708 2777
rect 2702 2772 2708 2773
rect 2840 2772 2842 2782
rect 2870 2777 2876 2778
rect 3007 2777 3011 2778
rect 2870 2773 2871 2777
rect 2875 2773 2876 2777
rect 2870 2772 2876 2773
rect 2558 2770 2564 2771
rect 2838 2771 2844 2772
rect 2374 2748 2380 2749
rect 2374 2744 2375 2748
rect 2379 2744 2380 2748
rect 2374 2743 2380 2744
rect 2534 2748 2540 2749
rect 2534 2744 2535 2748
rect 2539 2744 2540 2748
rect 2534 2743 2540 2744
rect 2376 2739 2378 2743
rect 2536 2739 2538 2743
rect 2375 2738 2379 2739
rect 2375 2733 2379 2734
rect 2383 2738 2387 2739
rect 2383 2733 2387 2734
rect 2535 2738 2539 2739
rect 2535 2733 2539 2734
rect 2382 2732 2388 2733
rect 2382 2728 2383 2732
rect 2387 2728 2388 2732
rect 2382 2727 2388 2728
rect 2560 2712 2562 2770
rect 2838 2767 2839 2771
rect 2843 2767 2844 2771
rect 2838 2766 2844 2767
rect 2702 2748 2708 2749
rect 2702 2744 2703 2748
rect 2707 2744 2708 2748
rect 2702 2743 2708 2744
rect 2704 2739 2706 2743
rect 2575 2738 2579 2739
rect 2575 2733 2579 2734
rect 2703 2738 2707 2739
rect 2703 2733 2707 2734
rect 2775 2738 2779 2739
rect 2775 2733 2779 2734
rect 2574 2732 2580 2733
rect 2574 2728 2575 2732
rect 2579 2728 2580 2732
rect 2574 2727 2580 2728
rect 2774 2732 2780 2733
rect 2774 2728 2775 2732
rect 2779 2728 2780 2732
rect 2774 2727 2780 2728
rect 2558 2711 2564 2712
rect 2558 2707 2559 2711
rect 2563 2707 2564 2711
rect 2840 2708 2842 2766
rect 2870 2748 2876 2749
rect 2870 2744 2871 2748
rect 2875 2744 2876 2748
rect 2870 2743 2876 2744
rect 2872 2739 2874 2743
rect 2871 2738 2875 2739
rect 2871 2733 2875 2734
rect 2975 2738 2979 2739
rect 2975 2733 2979 2734
rect 2974 2732 2980 2733
rect 2974 2728 2975 2732
rect 2979 2728 2980 2732
rect 2974 2727 2980 2728
rect 2558 2706 2564 2707
rect 2782 2707 2788 2708
rect 2382 2703 2388 2704
rect 2382 2699 2383 2703
rect 2387 2699 2388 2703
rect 2382 2698 2388 2699
rect 2390 2703 2396 2704
rect 2390 2699 2391 2703
rect 2395 2699 2396 2703
rect 2390 2698 2396 2699
rect 2446 2703 2452 2704
rect 2446 2699 2447 2703
rect 2451 2699 2452 2703
rect 2446 2698 2452 2699
rect 2384 2691 2386 2698
rect 2359 2690 2363 2691
rect 2383 2690 2387 2691
rect 2358 2685 2364 2686
rect 2383 2685 2387 2686
rect 2358 2681 2359 2685
rect 2363 2681 2364 2685
rect 2392 2684 2394 2698
rect 2358 2680 2364 2681
rect 2390 2683 2396 2684
rect 1670 2676 1676 2677
rect 2006 2679 2012 2680
rect 1446 2674 1452 2675
rect 1574 2675 1580 2676
rect 966 2670 972 2671
rect 1078 2671 1084 2672
rect 958 2666 964 2667
rect 832 2659 834 2666
rect 831 2658 835 2659
rect 855 2658 859 2659
rect 831 2653 835 2654
rect 854 2653 860 2654
rect 734 2648 740 2649
rect 742 2651 748 2652
rect 630 2646 636 2647
rect 742 2647 743 2651
rect 747 2647 748 2651
rect 854 2649 855 2653
rect 859 2649 860 2653
rect 854 2648 860 2649
rect 864 2648 866 2666
rect 960 2659 962 2666
rect 959 2658 963 2659
rect 959 2653 963 2654
rect 968 2648 970 2670
rect 1078 2667 1079 2671
rect 1083 2667 1084 2671
rect 1078 2666 1084 2667
rect 1102 2671 1108 2672
rect 1102 2667 1103 2671
rect 1107 2667 1108 2671
rect 1102 2666 1108 2667
rect 1198 2671 1204 2672
rect 1198 2667 1199 2671
rect 1203 2667 1204 2671
rect 1198 2666 1204 2667
rect 1206 2671 1212 2672
rect 1206 2667 1207 2671
rect 1211 2667 1212 2671
rect 1310 2671 1316 2672
rect 1310 2667 1311 2671
rect 1315 2667 1316 2671
rect 1206 2666 1218 2667
rect 1310 2666 1316 2667
rect 1080 2659 1082 2666
rect 975 2658 979 2659
rect 1079 2658 1083 2659
rect 1095 2658 1099 2659
rect 974 2653 980 2654
rect 1079 2653 1083 2654
rect 1094 2653 1100 2654
rect 974 2649 975 2653
rect 979 2649 980 2653
rect 974 2648 980 2649
rect 1094 2649 1095 2653
rect 1099 2649 1100 2653
rect 1094 2648 1100 2649
rect 1104 2648 1106 2666
rect 1200 2659 1202 2666
rect 1208 2665 1218 2666
rect 1199 2658 1203 2659
rect 1207 2658 1211 2659
rect 1199 2653 1203 2654
rect 1206 2653 1212 2654
rect 1206 2649 1207 2653
rect 1211 2649 1212 2653
rect 1206 2648 1212 2649
rect 1216 2648 1218 2665
rect 1312 2659 1314 2666
rect 1311 2658 1315 2659
rect 1319 2658 1323 2659
rect 1311 2653 1315 2654
rect 1318 2653 1324 2654
rect 1318 2649 1319 2653
rect 1323 2649 1324 2653
rect 1344 2652 1346 2674
rect 1422 2671 1428 2672
rect 1422 2667 1423 2671
rect 1427 2667 1428 2671
rect 1422 2666 1428 2667
rect 1424 2659 1426 2666
rect 1423 2658 1427 2659
rect 1439 2658 1443 2659
rect 1423 2653 1427 2654
rect 1438 2653 1444 2654
rect 1318 2648 1324 2649
rect 1342 2651 1348 2652
rect 742 2646 748 2647
rect 862 2647 868 2648
rect 110 2644 116 2645
rect 862 2643 863 2647
rect 867 2643 868 2647
rect 862 2642 868 2643
rect 966 2647 972 2648
rect 966 2643 967 2647
rect 971 2643 972 2647
rect 966 2642 972 2643
rect 1102 2647 1108 2648
rect 1102 2643 1103 2647
rect 1107 2643 1108 2647
rect 1102 2642 1108 2643
rect 1214 2647 1220 2648
rect 1214 2643 1215 2647
rect 1219 2643 1220 2647
rect 1342 2647 1343 2651
rect 1347 2647 1348 2651
rect 1438 2649 1439 2653
rect 1443 2649 1444 2653
rect 1448 2652 1450 2674
rect 1542 2671 1548 2672
rect 1542 2667 1543 2671
rect 1547 2667 1548 2671
rect 1574 2671 1575 2675
rect 1579 2671 1580 2675
rect 1574 2670 1580 2671
rect 1630 2675 1636 2676
rect 1630 2671 1631 2675
rect 1635 2671 1636 2675
rect 2006 2675 2007 2679
rect 2011 2675 2012 2679
rect 2006 2674 2012 2675
rect 2022 2679 2028 2680
rect 2022 2675 2023 2679
rect 2027 2675 2028 2679
rect 2022 2674 2028 2675
rect 2206 2679 2212 2680
rect 2206 2675 2207 2679
rect 2211 2675 2212 2679
rect 2206 2674 2212 2675
rect 2350 2679 2356 2680
rect 2350 2675 2351 2679
rect 2355 2675 2356 2679
rect 2390 2679 2391 2683
rect 2395 2679 2396 2683
rect 2390 2678 2396 2679
rect 2350 2674 2356 2675
rect 1630 2670 1636 2671
rect 1542 2666 1548 2667
rect 1544 2659 1546 2666
rect 1632 2659 1634 2670
rect 1670 2663 1676 2664
rect 1670 2659 1671 2663
rect 1675 2659 1676 2663
rect 1543 2658 1547 2659
rect 1543 2653 1547 2654
rect 1631 2658 1635 2659
rect 1670 2658 1676 2659
rect 1631 2653 1635 2654
rect 1438 2648 1444 2649
rect 1446 2651 1452 2652
rect 1342 2646 1348 2647
rect 1446 2647 1447 2651
rect 1451 2647 1452 2651
rect 1632 2650 1634 2653
rect 1672 2651 1674 2658
rect 1998 2656 2004 2657
rect 1998 2652 1999 2656
rect 2003 2652 2004 2656
rect 1998 2651 2004 2652
rect 1671 2650 1675 2651
rect 1446 2646 1452 2647
rect 1630 2649 1636 2650
rect 1214 2642 1226 2643
rect 110 2631 116 2632
rect 110 2627 111 2631
rect 115 2627 116 2631
rect 110 2626 116 2627
rect 112 2607 114 2626
rect 606 2624 612 2625
rect 606 2620 607 2624
rect 611 2620 612 2624
rect 606 2619 612 2620
rect 734 2624 740 2625
rect 734 2620 735 2624
rect 739 2620 740 2624
rect 734 2619 740 2620
rect 854 2624 860 2625
rect 854 2620 855 2624
rect 859 2620 860 2624
rect 854 2619 860 2620
rect 608 2607 610 2619
rect 736 2607 738 2619
rect 856 2607 858 2619
rect 111 2606 115 2607
rect 111 2601 115 2602
rect 503 2606 507 2607
rect 503 2601 507 2602
rect 607 2606 611 2607
rect 607 2601 611 2602
rect 631 2606 635 2607
rect 631 2601 635 2602
rect 735 2606 739 2607
rect 735 2601 739 2602
rect 751 2606 755 2607
rect 751 2601 755 2602
rect 855 2606 859 2607
rect 855 2601 859 2602
rect 112 2594 114 2601
rect 502 2600 508 2601
rect 502 2596 503 2600
rect 507 2596 508 2600
rect 502 2595 508 2596
rect 630 2600 636 2601
rect 630 2596 631 2600
rect 635 2596 636 2600
rect 630 2595 636 2596
rect 750 2600 756 2601
rect 750 2596 751 2600
rect 755 2596 756 2600
rect 750 2595 756 2596
rect 110 2593 116 2594
rect 110 2589 111 2593
rect 115 2589 116 2593
rect 110 2588 116 2589
rect 864 2580 866 2642
rect 1216 2641 1226 2642
rect 974 2624 980 2625
rect 974 2620 975 2624
rect 979 2620 980 2624
rect 974 2619 980 2620
rect 1094 2624 1100 2625
rect 1094 2620 1095 2624
rect 1099 2620 1100 2624
rect 1094 2619 1100 2620
rect 1206 2624 1212 2625
rect 1206 2620 1207 2624
rect 1211 2620 1212 2624
rect 1206 2619 1212 2620
rect 976 2607 978 2619
rect 1096 2607 1098 2619
rect 1208 2607 1210 2619
rect 871 2606 875 2607
rect 871 2601 875 2602
rect 975 2606 979 2607
rect 975 2601 979 2602
rect 991 2606 995 2607
rect 991 2601 995 2602
rect 1095 2606 1099 2607
rect 1095 2601 1099 2602
rect 1103 2606 1107 2607
rect 1103 2601 1107 2602
rect 1207 2606 1211 2607
rect 1207 2601 1211 2602
rect 1215 2606 1219 2607
rect 1215 2601 1219 2602
rect 870 2600 876 2601
rect 870 2596 871 2600
rect 875 2596 876 2600
rect 870 2595 876 2596
rect 990 2600 996 2601
rect 990 2596 991 2600
rect 995 2596 996 2600
rect 990 2595 996 2596
rect 1102 2600 1108 2601
rect 1102 2596 1103 2600
rect 1107 2596 1108 2600
rect 1102 2595 1108 2596
rect 1214 2600 1220 2601
rect 1214 2596 1215 2600
rect 1219 2596 1220 2600
rect 1214 2595 1220 2596
rect 862 2579 868 2580
rect 110 2575 116 2576
rect 110 2571 111 2575
rect 115 2571 116 2575
rect 862 2575 863 2579
rect 867 2575 868 2579
rect 862 2574 868 2575
rect 902 2579 908 2580
rect 902 2575 903 2579
rect 907 2575 908 2579
rect 1224 2576 1226 2641
rect 1318 2624 1324 2625
rect 1318 2620 1319 2624
rect 1323 2620 1324 2624
rect 1318 2619 1324 2620
rect 1320 2607 1322 2619
rect 1319 2606 1323 2607
rect 1319 2601 1323 2602
rect 1335 2606 1339 2607
rect 1335 2601 1339 2602
rect 1334 2600 1340 2601
rect 1334 2596 1335 2600
rect 1339 2596 1340 2600
rect 1334 2595 1340 2596
rect 1344 2576 1346 2646
rect 1630 2645 1631 2649
rect 1635 2645 1636 2649
rect 1671 2645 1675 2646
rect 1911 2650 1915 2651
rect 1911 2645 1915 2646
rect 1999 2650 2003 2651
rect 1999 2645 2003 2646
rect 1630 2644 1636 2645
rect 1672 2638 1674 2645
rect 1910 2644 1916 2645
rect 1910 2640 1911 2644
rect 1915 2640 1916 2644
rect 1910 2639 1916 2640
rect 1670 2637 1676 2638
rect 1670 2633 1671 2637
rect 1675 2633 1676 2637
rect 1670 2632 1676 2633
rect 1630 2631 1636 2632
rect 1630 2627 1631 2631
rect 1635 2627 1636 2631
rect 1630 2626 1636 2627
rect 1438 2624 1444 2625
rect 1438 2620 1439 2624
rect 1443 2620 1444 2624
rect 1438 2619 1444 2620
rect 1440 2607 1442 2619
rect 1632 2607 1634 2626
rect 1670 2619 1676 2620
rect 1670 2615 1671 2619
rect 1675 2615 1676 2619
rect 1670 2614 1676 2615
rect 1910 2615 1916 2616
rect 1672 2611 1674 2614
rect 1910 2611 1911 2615
rect 1915 2611 1916 2615
rect 1671 2610 1675 2611
rect 1439 2606 1443 2607
rect 1439 2601 1443 2602
rect 1631 2606 1635 2607
rect 1823 2610 1827 2611
rect 1910 2610 1916 2611
rect 1918 2615 1924 2616
rect 1918 2611 1919 2615
rect 1923 2611 1924 2615
rect 1918 2610 1924 2611
rect 1671 2605 1675 2606
rect 1822 2605 1828 2606
rect 1911 2605 1915 2606
rect 1672 2602 1674 2605
rect 1631 2601 1635 2602
rect 1670 2601 1676 2602
rect 1632 2594 1634 2601
rect 1670 2597 1671 2601
rect 1675 2597 1676 2601
rect 1822 2601 1823 2605
rect 1827 2601 1828 2605
rect 1822 2600 1828 2601
rect 1920 2600 1922 2610
rect 2008 2600 2010 2674
rect 2174 2656 2180 2657
rect 2174 2652 2175 2656
rect 2179 2652 2180 2656
rect 2174 2651 2180 2652
rect 2103 2650 2107 2651
rect 2103 2645 2107 2646
rect 2175 2650 2179 2651
rect 2175 2645 2179 2646
rect 2102 2644 2108 2645
rect 2102 2640 2103 2644
rect 2107 2640 2108 2644
rect 2102 2639 2108 2640
rect 2102 2615 2108 2616
rect 2102 2611 2103 2615
rect 2107 2611 2108 2615
rect 2015 2610 2019 2611
rect 2102 2610 2108 2611
rect 2014 2605 2020 2606
rect 2103 2605 2107 2606
rect 2014 2601 2015 2605
rect 2019 2601 2020 2605
rect 2014 2600 2020 2601
rect 2208 2600 2210 2674
rect 2295 2650 2299 2651
rect 2295 2645 2299 2646
rect 2294 2644 2300 2645
rect 2294 2640 2295 2644
rect 2299 2640 2300 2644
rect 2294 2639 2300 2640
rect 2352 2620 2354 2674
rect 2358 2656 2364 2657
rect 2358 2652 2359 2656
rect 2363 2652 2364 2656
rect 2358 2651 2364 2652
rect 2359 2650 2363 2651
rect 2359 2645 2363 2646
rect 2326 2619 2332 2620
rect 2294 2615 2300 2616
rect 2294 2611 2295 2615
rect 2299 2611 2300 2615
rect 2326 2615 2327 2619
rect 2331 2615 2332 2619
rect 2326 2614 2332 2615
rect 2350 2619 2356 2620
rect 2350 2615 2351 2619
rect 2355 2615 2356 2619
rect 2350 2614 2356 2615
rect 2215 2610 2219 2611
rect 2294 2610 2300 2611
rect 2214 2605 2220 2606
rect 2295 2605 2299 2606
rect 2214 2601 2215 2605
rect 2219 2601 2220 2605
rect 2214 2600 2220 2601
rect 1670 2596 1676 2597
rect 1830 2599 1836 2600
rect 1830 2595 1831 2599
rect 1835 2595 1836 2599
rect 1830 2594 1836 2595
rect 1918 2599 1924 2600
rect 1918 2595 1919 2599
rect 1923 2595 1924 2599
rect 1918 2594 1924 2595
rect 2006 2599 2012 2600
rect 2006 2595 2007 2599
rect 2011 2595 2012 2599
rect 2006 2594 2012 2595
rect 2062 2599 2068 2600
rect 2062 2595 2063 2599
rect 2067 2595 2068 2599
rect 2062 2594 2068 2595
rect 2206 2599 2212 2600
rect 2206 2595 2207 2599
rect 2211 2595 2212 2599
rect 2206 2594 2212 2595
rect 2222 2599 2228 2600
rect 2222 2595 2223 2599
rect 2227 2595 2228 2599
rect 2222 2594 2228 2595
rect 1630 2593 1636 2594
rect 1630 2589 1631 2593
rect 1635 2589 1636 2593
rect 1630 2588 1636 2589
rect 1670 2583 1676 2584
rect 1670 2579 1671 2583
rect 1675 2579 1676 2583
rect 1670 2578 1676 2579
rect 902 2574 908 2575
rect 1014 2575 1020 2576
rect 110 2570 116 2571
rect 502 2571 508 2572
rect 112 2555 114 2570
rect 502 2567 503 2571
rect 507 2567 508 2571
rect 502 2566 508 2567
rect 510 2571 516 2572
rect 510 2567 511 2571
rect 515 2567 516 2571
rect 510 2566 516 2567
rect 630 2571 636 2572
rect 630 2567 631 2571
rect 635 2567 636 2571
rect 630 2566 636 2567
rect 638 2571 644 2572
rect 638 2567 639 2571
rect 643 2567 644 2571
rect 638 2566 644 2567
rect 750 2571 756 2572
rect 750 2567 751 2571
rect 755 2567 756 2571
rect 750 2566 756 2567
rect 782 2571 788 2572
rect 782 2567 783 2571
rect 787 2567 788 2571
rect 782 2566 788 2567
rect 504 2555 506 2566
rect 111 2554 115 2555
rect 399 2554 403 2555
rect 503 2554 507 2555
rect 111 2549 115 2550
rect 398 2549 404 2550
rect 503 2549 507 2550
rect 112 2546 114 2549
rect 110 2545 116 2546
rect 110 2541 111 2545
rect 115 2541 116 2545
rect 398 2545 399 2549
rect 403 2545 404 2549
rect 398 2544 404 2545
rect 512 2544 514 2566
rect 632 2555 634 2566
rect 527 2554 531 2555
rect 631 2554 635 2555
rect 526 2549 532 2550
rect 631 2549 635 2550
rect 526 2545 527 2549
rect 531 2545 532 2549
rect 526 2544 532 2545
rect 640 2544 642 2566
rect 752 2555 754 2566
rect 655 2554 659 2555
rect 751 2554 755 2555
rect 775 2554 779 2555
rect 654 2549 660 2550
rect 751 2549 755 2550
rect 774 2549 780 2550
rect 654 2545 655 2549
rect 659 2545 660 2549
rect 654 2544 660 2545
rect 774 2545 775 2549
rect 779 2545 780 2549
rect 784 2548 786 2566
rect 864 2548 866 2574
rect 870 2571 876 2572
rect 870 2567 871 2571
rect 875 2567 876 2571
rect 870 2566 876 2567
rect 872 2555 874 2566
rect 871 2554 875 2555
rect 895 2554 899 2555
rect 871 2549 875 2550
rect 894 2549 900 2550
rect 774 2544 780 2545
rect 782 2547 788 2548
rect 110 2540 116 2541
rect 442 2543 448 2544
rect 442 2539 443 2543
rect 447 2539 448 2543
rect 442 2538 448 2539
rect 510 2543 516 2544
rect 510 2539 511 2543
rect 515 2539 516 2543
rect 510 2538 516 2539
rect 638 2543 644 2544
rect 638 2539 639 2543
rect 643 2539 644 2543
rect 782 2543 783 2547
rect 787 2543 788 2547
rect 782 2542 788 2543
rect 862 2547 868 2548
rect 862 2543 863 2547
rect 867 2543 868 2547
rect 894 2545 895 2549
rect 899 2545 900 2549
rect 904 2548 906 2574
rect 990 2571 996 2572
rect 990 2567 991 2571
rect 995 2567 996 2571
rect 1014 2571 1015 2575
rect 1019 2571 1020 2575
rect 1222 2575 1228 2576
rect 1014 2570 1020 2571
rect 1102 2571 1108 2572
rect 990 2566 996 2567
rect 992 2555 994 2566
rect 991 2554 995 2555
rect 1007 2554 1011 2555
rect 991 2549 995 2550
rect 1006 2549 1012 2550
rect 894 2544 900 2545
rect 902 2547 908 2548
rect 862 2542 868 2543
rect 902 2543 903 2547
rect 907 2543 908 2547
rect 1006 2545 1007 2549
rect 1011 2545 1012 2549
rect 1016 2548 1018 2570
rect 1102 2567 1103 2571
rect 1107 2567 1108 2571
rect 1102 2566 1108 2567
rect 1126 2571 1132 2572
rect 1126 2567 1127 2571
rect 1131 2567 1132 2571
rect 1126 2566 1132 2567
rect 1214 2571 1220 2572
rect 1214 2567 1215 2571
rect 1219 2567 1220 2571
rect 1222 2571 1223 2575
rect 1227 2571 1228 2575
rect 1222 2570 1228 2571
rect 1246 2575 1252 2576
rect 1246 2571 1247 2575
rect 1251 2571 1252 2575
rect 1342 2575 1348 2576
rect 1246 2570 1252 2571
rect 1334 2571 1340 2572
rect 1214 2566 1220 2567
rect 1104 2555 1106 2566
rect 1103 2554 1107 2555
rect 1119 2554 1123 2555
rect 1103 2549 1107 2550
rect 1118 2549 1124 2550
rect 1006 2544 1012 2545
rect 1014 2547 1020 2548
rect 902 2542 908 2543
rect 1014 2543 1015 2547
rect 1019 2543 1020 2547
rect 1118 2545 1119 2549
rect 1123 2545 1124 2549
rect 1118 2544 1124 2545
rect 1128 2544 1130 2566
rect 1216 2555 1218 2566
rect 1215 2554 1219 2555
rect 1239 2554 1243 2555
rect 1215 2549 1219 2550
rect 1238 2549 1244 2550
rect 1238 2545 1239 2549
rect 1243 2545 1244 2549
rect 1248 2548 1250 2570
rect 1334 2567 1335 2571
rect 1339 2567 1340 2571
rect 1342 2571 1343 2575
rect 1347 2571 1348 2575
rect 1342 2570 1348 2571
rect 1630 2575 1636 2576
rect 1630 2571 1631 2575
rect 1635 2571 1636 2575
rect 1630 2570 1636 2571
rect 1334 2566 1340 2567
rect 1336 2555 1338 2566
rect 1632 2555 1634 2570
rect 1672 2567 1674 2578
rect 1822 2576 1828 2577
rect 1822 2572 1823 2576
rect 1827 2572 1828 2576
rect 1822 2571 1828 2572
rect 1824 2567 1826 2571
rect 1671 2566 1675 2567
rect 1671 2561 1675 2562
rect 1735 2566 1739 2567
rect 1735 2561 1739 2562
rect 1823 2566 1827 2567
rect 1823 2561 1827 2562
rect 1335 2554 1339 2555
rect 1335 2549 1339 2550
rect 1631 2554 1635 2555
rect 1672 2554 1674 2561
rect 1734 2560 1740 2561
rect 1734 2556 1735 2560
rect 1739 2556 1740 2560
rect 1734 2555 1740 2556
rect 1631 2549 1635 2550
rect 1670 2553 1676 2554
rect 1670 2549 1671 2553
rect 1675 2549 1676 2553
rect 1238 2544 1244 2545
rect 1246 2547 1252 2548
rect 1014 2542 1020 2543
rect 1126 2543 1132 2544
rect 638 2538 644 2539
rect 110 2527 116 2528
rect 110 2523 111 2527
rect 115 2523 116 2527
rect 110 2522 116 2523
rect 112 2503 114 2522
rect 398 2520 404 2521
rect 398 2516 399 2520
rect 403 2516 404 2520
rect 398 2515 404 2516
rect 400 2503 402 2515
rect 111 2502 115 2503
rect 111 2497 115 2498
rect 303 2502 307 2503
rect 303 2497 307 2498
rect 399 2502 403 2503
rect 399 2497 403 2498
rect 431 2502 435 2503
rect 431 2497 435 2498
rect 112 2490 114 2497
rect 302 2496 308 2497
rect 302 2492 303 2496
rect 307 2492 308 2496
rect 302 2491 308 2492
rect 430 2496 436 2497
rect 430 2492 431 2496
rect 435 2492 436 2496
rect 430 2491 436 2492
rect 110 2489 116 2490
rect 110 2485 111 2489
rect 115 2485 116 2489
rect 110 2484 116 2485
rect 444 2473 446 2538
rect 526 2520 532 2521
rect 526 2516 527 2520
rect 531 2516 532 2520
rect 526 2515 532 2516
rect 654 2520 660 2521
rect 654 2516 655 2520
rect 659 2516 660 2520
rect 654 2515 660 2516
rect 774 2520 780 2521
rect 774 2516 775 2520
rect 779 2516 780 2520
rect 774 2515 780 2516
rect 528 2503 530 2515
rect 656 2503 658 2515
rect 776 2503 778 2515
rect 527 2502 531 2503
rect 527 2497 531 2498
rect 559 2502 563 2503
rect 559 2497 563 2498
rect 655 2502 659 2503
rect 655 2497 659 2498
rect 703 2502 707 2503
rect 703 2497 707 2498
rect 775 2502 779 2503
rect 775 2497 779 2498
rect 558 2496 564 2497
rect 558 2492 559 2496
rect 563 2492 564 2496
rect 558 2491 564 2492
rect 702 2496 708 2497
rect 702 2492 703 2496
rect 707 2492 708 2496
rect 702 2491 708 2492
rect 784 2473 786 2542
rect 894 2520 900 2521
rect 894 2516 895 2520
rect 899 2516 900 2520
rect 894 2515 900 2516
rect 896 2503 898 2515
rect 863 2502 867 2503
rect 863 2497 867 2498
rect 895 2502 899 2503
rect 895 2497 899 2498
rect 862 2496 868 2497
rect 862 2492 863 2496
rect 867 2492 868 2496
rect 862 2491 868 2492
rect 110 2471 116 2472
rect 110 2467 111 2471
rect 115 2467 116 2471
rect 440 2471 446 2473
rect 776 2471 786 2473
rect 904 2472 906 2542
rect 1126 2539 1127 2543
rect 1131 2539 1132 2543
rect 1246 2543 1247 2547
rect 1251 2543 1252 2547
rect 1632 2546 1634 2549
rect 1670 2548 1676 2549
rect 1246 2542 1252 2543
rect 1630 2545 1636 2546
rect 1126 2538 1132 2539
rect 1006 2520 1012 2521
rect 1006 2516 1007 2520
rect 1011 2516 1012 2520
rect 1006 2515 1012 2516
rect 1118 2520 1124 2521
rect 1118 2516 1119 2520
rect 1123 2516 1124 2520
rect 1118 2515 1124 2516
rect 1008 2503 1010 2515
rect 1120 2503 1122 2515
rect 1007 2502 1011 2503
rect 1007 2497 1011 2498
rect 1039 2502 1043 2503
rect 1039 2497 1043 2498
rect 1119 2502 1123 2503
rect 1119 2497 1123 2498
rect 1038 2496 1044 2497
rect 1038 2492 1039 2496
rect 1043 2492 1044 2496
rect 1038 2491 1044 2492
rect 1128 2472 1130 2538
rect 1238 2520 1244 2521
rect 1238 2516 1239 2520
rect 1243 2516 1244 2520
rect 1238 2515 1244 2516
rect 1240 2503 1242 2515
rect 1223 2502 1227 2503
rect 1223 2497 1227 2498
rect 1239 2502 1243 2503
rect 1239 2497 1243 2498
rect 1222 2496 1228 2497
rect 1222 2492 1223 2496
rect 1227 2492 1228 2496
rect 1222 2491 1228 2492
rect 902 2471 908 2472
rect 440 2468 442 2471
rect 776 2468 778 2471
rect 110 2466 116 2467
rect 302 2467 308 2468
rect 112 2459 114 2466
rect 302 2463 303 2467
rect 307 2463 308 2467
rect 302 2462 308 2463
rect 310 2467 316 2468
rect 310 2463 311 2467
rect 315 2463 316 2467
rect 310 2462 316 2463
rect 430 2467 436 2468
rect 430 2463 431 2467
rect 435 2463 436 2467
rect 430 2462 436 2463
rect 438 2467 444 2468
rect 438 2463 439 2467
rect 443 2463 444 2467
rect 438 2462 444 2463
rect 558 2467 564 2468
rect 558 2463 559 2467
rect 563 2463 564 2467
rect 558 2462 564 2463
rect 610 2467 616 2468
rect 610 2463 611 2467
rect 615 2463 616 2467
rect 610 2462 616 2463
rect 702 2467 708 2468
rect 702 2463 703 2467
rect 707 2463 708 2467
rect 702 2462 708 2463
rect 774 2467 780 2468
rect 774 2463 775 2467
rect 779 2463 780 2467
rect 774 2462 780 2463
rect 862 2467 868 2468
rect 862 2463 863 2467
rect 867 2463 868 2467
rect 902 2467 903 2471
rect 907 2467 908 2471
rect 1046 2471 1052 2472
rect 902 2466 908 2467
rect 1038 2467 1044 2468
rect 862 2462 868 2463
rect 1038 2463 1039 2467
rect 1043 2463 1044 2467
rect 1046 2467 1047 2471
rect 1051 2467 1052 2471
rect 1046 2466 1052 2467
rect 1126 2471 1132 2472
rect 1126 2467 1127 2471
rect 1131 2467 1132 2471
rect 1248 2468 1250 2542
rect 1630 2541 1631 2545
rect 1635 2541 1636 2545
rect 1630 2540 1636 2541
rect 1670 2535 1676 2536
rect 1670 2531 1671 2535
rect 1675 2531 1676 2535
rect 1670 2530 1676 2531
rect 1734 2531 1740 2532
rect 1630 2527 1636 2528
rect 1630 2523 1631 2527
rect 1635 2523 1636 2527
rect 1672 2523 1674 2530
rect 1734 2527 1735 2531
rect 1739 2527 1740 2531
rect 1734 2526 1740 2527
rect 1736 2523 1738 2526
rect 1630 2522 1636 2523
rect 1671 2522 1675 2523
rect 1632 2503 1634 2522
rect 1695 2522 1699 2523
rect 1735 2522 1739 2523
rect 1671 2517 1675 2518
rect 1694 2517 1700 2518
rect 1735 2517 1739 2518
rect 1672 2514 1674 2517
rect 1670 2513 1676 2514
rect 1670 2509 1671 2513
rect 1675 2509 1676 2513
rect 1694 2513 1695 2517
rect 1699 2513 1700 2517
rect 1694 2512 1700 2513
rect 1832 2512 1834 2594
rect 1895 2566 1899 2567
rect 1895 2561 1899 2562
rect 1894 2560 1900 2561
rect 1894 2556 1895 2560
rect 1899 2556 1900 2560
rect 1894 2555 1900 2556
rect 1920 2532 1922 2594
rect 2014 2576 2020 2577
rect 2014 2572 2015 2576
rect 2019 2572 2020 2576
rect 2014 2571 2020 2572
rect 2016 2567 2018 2571
rect 2015 2566 2019 2567
rect 2015 2561 2019 2562
rect 2055 2566 2059 2567
rect 2055 2561 2059 2562
rect 2054 2560 2060 2561
rect 2054 2556 2055 2560
rect 2059 2556 2060 2560
rect 2054 2555 2060 2556
rect 2064 2536 2066 2594
rect 2214 2576 2220 2577
rect 2214 2572 2215 2576
rect 2219 2572 2220 2576
rect 2214 2571 2220 2572
rect 2216 2567 2218 2571
rect 2215 2566 2219 2567
rect 2215 2561 2219 2562
rect 2214 2560 2220 2561
rect 2214 2556 2215 2560
rect 2219 2556 2220 2560
rect 2214 2555 2220 2556
rect 2224 2536 2226 2594
rect 2062 2535 2068 2536
rect 1894 2531 1900 2532
rect 1894 2527 1895 2531
rect 1899 2527 1900 2531
rect 1894 2526 1900 2527
rect 1902 2531 1908 2532
rect 1902 2527 1903 2531
rect 1907 2527 1908 2531
rect 1902 2526 1908 2527
rect 1918 2531 1924 2532
rect 1918 2527 1919 2531
rect 1923 2527 1924 2531
rect 1918 2526 1924 2527
rect 2054 2531 2060 2532
rect 2054 2527 2055 2531
rect 2059 2527 2060 2531
rect 2062 2531 2063 2535
rect 2067 2531 2068 2535
rect 2222 2535 2228 2536
rect 2062 2530 2068 2531
rect 2214 2531 2220 2532
rect 2054 2526 2060 2527
rect 1896 2523 1898 2526
rect 1863 2522 1867 2523
rect 1895 2522 1899 2523
rect 1862 2517 1868 2518
rect 1895 2517 1899 2518
rect 1862 2513 1863 2517
rect 1867 2513 1868 2517
rect 1862 2512 1868 2513
rect 1904 2512 1906 2526
rect 2056 2523 2058 2526
rect 2055 2522 2059 2523
rect 2055 2517 2059 2518
rect 2064 2512 2066 2530
rect 2214 2527 2215 2531
rect 2219 2527 2220 2531
rect 2222 2531 2223 2535
rect 2227 2531 2228 2535
rect 2222 2530 2228 2531
rect 2214 2526 2220 2527
rect 2216 2523 2218 2526
rect 2079 2522 2083 2523
rect 2215 2522 2219 2523
rect 2319 2522 2323 2523
rect 2078 2517 2084 2518
rect 2215 2517 2219 2518
rect 2318 2517 2324 2518
rect 2078 2513 2079 2517
rect 2083 2513 2084 2517
rect 2078 2512 2084 2513
rect 2318 2513 2319 2517
rect 2323 2513 2324 2517
rect 2328 2516 2330 2614
rect 2439 2610 2443 2611
rect 2438 2605 2444 2606
rect 2438 2601 2439 2605
rect 2443 2601 2444 2605
rect 2448 2604 2450 2698
rect 2551 2690 2555 2691
rect 2550 2685 2556 2686
rect 2550 2681 2551 2685
rect 2555 2681 2556 2685
rect 2560 2684 2562 2706
rect 2574 2703 2580 2704
rect 2574 2699 2575 2703
rect 2579 2699 2580 2703
rect 2574 2698 2580 2699
rect 2774 2703 2780 2704
rect 2774 2699 2775 2703
rect 2779 2699 2780 2703
rect 2782 2703 2783 2707
rect 2787 2703 2788 2707
rect 2782 2702 2788 2703
rect 2838 2707 2844 2708
rect 2838 2703 2839 2707
rect 2843 2703 2844 2707
rect 2838 2702 2844 2703
rect 2926 2707 2932 2708
rect 2926 2703 2927 2707
rect 2931 2703 2932 2707
rect 3016 2704 3018 2782
rect 3159 2777 3163 2778
rect 3159 2738 3163 2739
rect 3159 2733 3163 2734
rect 3158 2732 3164 2733
rect 3158 2728 3159 2732
rect 3163 2728 3164 2732
rect 3158 2727 3164 2728
rect 3168 2704 3170 2782
rect 3191 2777 3195 2778
rect 3192 2774 3194 2777
rect 3190 2773 3196 2774
rect 3190 2769 3191 2773
rect 3195 2769 3196 2773
rect 3190 2768 3196 2769
rect 3190 2755 3196 2756
rect 3190 2751 3191 2755
rect 3195 2751 3196 2755
rect 3190 2750 3196 2751
rect 3192 2739 3194 2750
rect 3191 2738 3195 2739
rect 3191 2733 3195 2734
rect 3192 2726 3194 2733
rect 3190 2725 3196 2726
rect 3190 2721 3191 2725
rect 3195 2721 3196 2725
rect 3190 2720 3196 2721
rect 3190 2707 3196 2708
rect 2926 2702 2932 2703
rect 2974 2703 2980 2704
rect 2774 2698 2780 2699
rect 2576 2691 2578 2698
rect 2776 2691 2778 2698
rect 2575 2690 2579 2691
rect 2759 2690 2763 2691
rect 2775 2690 2779 2691
rect 2575 2685 2579 2686
rect 2758 2685 2764 2686
rect 2775 2685 2779 2686
rect 2550 2680 2556 2681
rect 2558 2683 2564 2684
rect 2558 2679 2559 2683
rect 2563 2679 2564 2683
rect 2758 2681 2759 2685
rect 2763 2681 2764 2685
rect 2784 2684 2786 2702
rect 2758 2680 2764 2681
rect 2782 2683 2788 2684
rect 2558 2678 2564 2679
rect 2782 2679 2783 2683
rect 2787 2679 2788 2683
rect 2928 2680 2930 2702
rect 2974 2699 2975 2703
rect 2979 2699 2980 2703
rect 2974 2698 2980 2699
rect 3014 2703 3020 2704
rect 3014 2699 3015 2703
rect 3019 2699 3020 2703
rect 3014 2698 3020 2699
rect 3158 2703 3164 2704
rect 3158 2699 3159 2703
rect 3163 2699 3164 2703
rect 3158 2698 3164 2699
rect 3166 2703 3172 2704
rect 3166 2699 3167 2703
rect 3171 2699 3172 2703
rect 3190 2703 3191 2707
rect 3195 2703 3196 2707
rect 3190 2702 3196 2703
rect 3166 2698 3172 2699
rect 2976 2691 2978 2698
rect 3160 2691 3162 2698
rect 2967 2690 2971 2691
rect 2975 2690 2979 2691
rect 3159 2690 3163 2691
rect 2966 2685 2972 2686
rect 2975 2685 2979 2686
rect 3158 2685 3164 2686
rect 2966 2681 2967 2685
rect 2971 2681 2972 2685
rect 2966 2680 2972 2681
rect 3158 2681 3159 2685
rect 3163 2681 3164 2685
rect 3158 2680 3164 2681
rect 3168 2680 3170 2698
rect 3192 2691 3194 2702
rect 3191 2690 3195 2691
rect 3191 2685 3195 2686
rect 3192 2682 3194 2685
rect 3190 2681 3196 2682
rect 2782 2678 2788 2679
rect 2926 2679 2932 2680
rect 2550 2656 2556 2657
rect 2550 2652 2551 2656
rect 2555 2652 2556 2656
rect 2550 2651 2556 2652
rect 2758 2656 2764 2657
rect 2758 2652 2759 2656
rect 2763 2652 2764 2656
rect 2758 2651 2764 2652
rect 2487 2650 2491 2651
rect 2487 2645 2491 2646
rect 2551 2650 2555 2651
rect 2551 2645 2555 2646
rect 2687 2650 2691 2651
rect 2687 2645 2691 2646
rect 2759 2650 2763 2651
rect 2759 2645 2763 2646
rect 2486 2644 2492 2645
rect 2486 2640 2487 2644
rect 2491 2640 2492 2644
rect 2486 2639 2492 2640
rect 2686 2644 2692 2645
rect 2686 2640 2687 2644
rect 2691 2640 2692 2644
rect 2686 2639 2692 2640
rect 2784 2620 2786 2678
rect 2926 2675 2927 2679
rect 2931 2675 2932 2679
rect 2926 2674 2932 2675
rect 3166 2679 3172 2680
rect 3166 2675 3167 2679
rect 3171 2675 3172 2679
rect 3190 2677 3191 2681
rect 3195 2677 3196 2681
rect 3190 2676 3196 2677
rect 3166 2674 3172 2675
rect 2782 2619 2788 2620
rect 2486 2615 2492 2616
rect 2486 2611 2487 2615
rect 2491 2611 2492 2615
rect 2686 2615 2692 2616
rect 2686 2611 2687 2615
rect 2691 2611 2692 2615
rect 2782 2615 2783 2619
rect 2787 2615 2788 2619
rect 2782 2614 2788 2615
rect 2486 2610 2492 2611
rect 2671 2610 2675 2611
rect 2686 2610 2692 2611
rect 2919 2610 2923 2611
rect 2487 2605 2491 2606
rect 2670 2605 2676 2606
rect 2687 2605 2691 2606
rect 2918 2605 2924 2606
rect 2438 2600 2444 2601
rect 2446 2603 2452 2604
rect 2446 2599 2447 2603
rect 2451 2599 2452 2603
rect 2670 2601 2671 2605
rect 2675 2601 2676 2605
rect 2670 2600 2676 2601
rect 2918 2601 2919 2605
rect 2923 2601 2924 2605
rect 2918 2600 2924 2601
rect 2928 2600 2930 2674
rect 2966 2656 2972 2657
rect 2966 2652 2967 2656
rect 2971 2652 2972 2656
rect 2966 2651 2972 2652
rect 3158 2656 3164 2657
rect 3158 2652 3159 2656
rect 3163 2652 3164 2656
rect 3158 2651 3164 2652
rect 2967 2650 2971 2651
rect 2967 2645 2971 2646
rect 3159 2650 3163 2651
rect 3159 2645 3163 2646
rect 3159 2610 3163 2611
rect 3158 2605 3164 2606
rect 3158 2601 3159 2605
rect 3163 2601 3164 2605
rect 3158 2600 3164 2601
rect 3168 2600 3170 2674
rect 3190 2663 3196 2664
rect 3190 2659 3191 2663
rect 3195 2659 3196 2663
rect 3190 2658 3196 2659
rect 3192 2651 3194 2658
rect 3191 2650 3195 2651
rect 3191 2645 3195 2646
rect 3192 2638 3194 2645
rect 3190 2637 3196 2638
rect 3190 2633 3191 2637
rect 3195 2633 3196 2637
rect 3190 2632 3196 2633
rect 3190 2619 3196 2620
rect 3190 2615 3191 2619
rect 3195 2615 3196 2619
rect 3190 2614 3196 2615
rect 3192 2611 3194 2614
rect 3191 2610 3195 2611
rect 3191 2605 3195 2606
rect 3192 2602 3194 2605
rect 3190 2601 3196 2602
rect 2446 2598 2452 2599
rect 2926 2599 2932 2600
rect 2926 2595 2927 2599
rect 2931 2595 2932 2599
rect 2926 2594 2932 2595
rect 3142 2599 3148 2600
rect 3142 2595 3143 2599
rect 3147 2595 3148 2599
rect 3142 2594 3148 2595
rect 3166 2599 3172 2600
rect 3166 2595 3167 2599
rect 3171 2595 3172 2599
rect 3190 2597 3191 2601
rect 3195 2597 3196 2601
rect 3190 2596 3196 2597
rect 3166 2594 3172 2595
rect 2438 2576 2444 2577
rect 2438 2572 2439 2576
rect 2443 2572 2444 2576
rect 2438 2571 2444 2572
rect 2670 2576 2676 2577
rect 2670 2572 2671 2576
rect 2675 2572 2676 2576
rect 2670 2571 2676 2572
rect 2918 2576 2924 2577
rect 2918 2572 2919 2576
rect 2923 2572 2924 2576
rect 2918 2571 2924 2572
rect 2440 2567 2442 2571
rect 2672 2567 2674 2571
rect 2920 2567 2922 2571
rect 2375 2566 2379 2567
rect 2375 2561 2379 2562
rect 2439 2566 2443 2567
rect 2439 2561 2443 2562
rect 2535 2566 2539 2567
rect 2535 2561 2539 2562
rect 2671 2566 2675 2567
rect 2671 2561 2675 2562
rect 2919 2566 2923 2567
rect 2919 2561 2923 2562
rect 2374 2560 2380 2561
rect 2374 2556 2375 2560
rect 2379 2556 2380 2560
rect 2374 2555 2380 2556
rect 2534 2560 2540 2561
rect 2534 2556 2535 2560
rect 2539 2556 2540 2560
rect 2534 2555 2540 2556
rect 2374 2531 2380 2532
rect 2374 2527 2375 2531
rect 2379 2527 2380 2531
rect 2374 2526 2380 2527
rect 2534 2531 2540 2532
rect 2534 2527 2535 2531
rect 2539 2527 2540 2531
rect 2534 2526 2540 2527
rect 2376 2523 2378 2526
rect 2536 2523 2538 2526
rect 2574 2523 2580 2524
rect 2375 2522 2379 2523
rect 2375 2517 2379 2518
rect 2535 2522 2539 2523
rect 2574 2519 2575 2523
rect 2579 2519 2580 2523
rect 2574 2518 2580 2519
rect 2583 2522 2587 2523
rect 2855 2522 2859 2523
rect 2535 2517 2539 2518
rect 2318 2512 2324 2513
rect 2326 2515 2332 2516
rect 1670 2508 1676 2509
rect 1830 2511 1836 2512
rect 1830 2507 1831 2511
rect 1835 2507 1836 2511
rect 1830 2506 1836 2507
rect 1902 2511 1908 2512
rect 1902 2507 1903 2511
rect 1907 2507 1908 2511
rect 1902 2506 1908 2507
rect 2062 2511 2068 2512
rect 2062 2507 2063 2511
rect 2067 2507 2068 2511
rect 2326 2511 2327 2515
rect 2331 2511 2332 2515
rect 2326 2510 2332 2511
rect 2062 2506 2068 2507
rect 1423 2502 1427 2503
rect 1423 2497 1427 2498
rect 1599 2502 1603 2503
rect 1599 2497 1603 2498
rect 1631 2502 1635 2503
rect 1631 2497 1635 2498
rect 1422 2496 1428 2497
rect 1422 2492 1423 2496
rect 1427 2492 1428 2496
rect 1422 2491 1428 2492
rect 1598 2496 1604 2497
rect 1598 2492 1599 2496
rect 1603 2492 1604 2496
rect 1598 2491 1604 2492
rect 1632 2490 1634 2497
rect 1670 2495 1676 2496
rect 1670 2491 1671 2495
rect 1675 2491 1676 2495
rect 1670 2490 1676 2491
rect 1630 2489 1636 2490
rect 1630 2485 1631 2489
rect 1635 2485 1636 2489
rect 1630 2484 1636 2485
rect 1382 2475 1388 2476
rect 1382 2471 1383 2475
rect 1387 2471 1388 2475
rect 1382 2470 1388 2471
rect 1574 2475 1580 2476
rect 1672 2475 1674 2490
rect 1694 2488 1700 2489
rect 1694 2484 1695 2488
rect 1699 2484 1700 2488
rect 1694 2483 1700 2484
rect 1862 2488 1868 2489
rect 1862 2484 1863 2488
rect 1867 2484 1868 2488
rect 1862 2483 1868 2484
rect 2078 2488 2084 2489
rect 2078 2484 2079 2488
rect 2083 2484 2084 2488
rect 2078 2483 2084 2484
rect 2318 2488 2324 2489
rect 2318 2484 2319 2488
rect 2323 2484 2324 2488
rect 2318 2483 2324 2484
rect 1696 2475 1698 2483
rect 1864 2475 1866 2483
rect 2080 2475 2082 2483
rect 2320 2475 2322 2483
rect 1574 2471 1575 2475
rect 1579 2471 1580 2475
rect 1671 2474 1675 2475
rect 1574 2470 1580 2471
rect 1630 2471 1636 2472
rect 1126 2466 1132 2467
rect 1222 2467 1228 2468
rect 1038 2462 1044 2463
rect 304 2459 306 2462
rect 111 2458 115 2459
rect 199 2458 203 2459
rect 303 2458 307 2459
rect 111 2453 115 2454
rect 198 2453 204 2454
rect 303 2453 307 2454
rect 112 2450 114 2453
rect 110 2449 116 2450
rect 110 2445 111 2449
rect 115 2445 116 2449
rect 198 2449 199 2453
rect 203 2449 204 2453
rect 198 2448 204 2449
rect 312 2448 314 2462
rect 432 2459 434 2462
rect 327 2458 331 2459
rect 431 2458 435 2459
rect 326 2453 332 2454
rect 431 2453 435 2454
rect 326 2449 327 2453
rect 331 2449 332 2453
rect 326 2448 332 2449
rect 440 2448 442 2462
rect 560 2459 562 2462
rect 455 2458 459 2459
rect 559 2458 563 2459
rect 599 2458 603 2459
rect 454 2453 460 2454
rect 559 2453 563 2454
rect 598 2453 604 2454
rect 454 2449 455 2453
rect 459 2449 460 2453
rect 454 2448 460 2449
rect 598 2449 599 2453
rect 603 2449 604 2453
rect 598 2448 604 2449
rect 612 2448 614 2462
rect 704 2459 706 2462
rect 703 2458 707 2459
rect 767 2458 771 2459
rect 703 2453 707 2454
rect 766 2453 772 2454
rect 766 2449 767 2453
rect 771 2449 772 2453
rect 766 2448 772 2449
rect 776 2448 778 2462
rect 864 2459 866 2462
rect 1040 2459 1042 2462
rect 863 2458 867 2459
rect 951 2458 955 2459
rect 1039 2458 1043 2459
rect 863 2453 867 2454
rect 950 2453 956 2454
rect 1039 2453 1043 2454
rect 950 2449 951 2453
rect 955 2449 956 2453
rect 1048 2452 1050 2466
rect 1222 2463 1223 2467
rect 1227 2463 1228 2467
rect 1222 2462 1228 2463
rect 1246 2467 1252 2468
rect 1246 2463 1247 2467
rect 1251 2463 1252 2467
rect 1246 2462 1252 2463
rect 1224 2459 1226 2462
rect 1159 2458 1163 2459
rect 1223 2458 1227 2459
rect 1158 2453 1164 2454
rect 1223 2453 1227 2454
rect 950 2448 956 2449
rect 1046 2451 1052 2452
rect 110 2444 116 2445
rect 246 2447 252 2448
rect 246 2443 247 2447
rect 251 2443 252 2447
rect 246 2442 252 2443
rect 310 2447 316 2448
rect 310 2443 311 2447
rect 315 2443 316 2447
rect 310 2442 316 2443
rect 438 2447 444 2448
rect 438 2443 439 2447
rect 443 2443 444 2447
rect 438 2442 444 2443
rect 610 2447 616 2448
rect 610 2443 611 2447
rect 615 2443 616 2447
rect 610 2442 616 2443
rect 774 2447 780 2448
rect 774 2443 775 2447
rect 779 2443 780 2447
rect 1046 2447 1047 2451
rect 1051 2447 1052 2451
rect 1158 2449 1159 2453
rect 1163 2449 1164 2453
rect 1248 2452 1250 2462
rect 1375 2458 1379 2459
rect 1374 2453 1380 2454
rect 1158 2448 1164 2449
rect 1182 2451 1188 2452
rect 1046 2446 1052 2447
rect 1182 2447 1183 2451
rect 1187 2447 1188 2451
rect 1182 2446 1188 2447
rect 1246 2451 1252 2452
rect 1246 2447 1247 2451
rect 1251 2447 1252 2451
rect 1374 2449 1375 2453
rect 1379 2449 1380 2453
rect 1384 2452 1386 2470
rect 1422 2467 1428 2468
rect 1422 2463 1423 2467
rect 1427 2463 1428 2467
rect 1422 2462 1428 2463
rect 1424 2459 1426 2462
rect 1423 2458 1427 2459
rect 1423 2453 1427 2454
rect 1374 2448 1380 2449
rect 1382 2451 1388 2452
rect 1246 2446 1252 2447
rect 1382 2447 1383 2451
rect 1387 2447 1388 2451
rect 1382 2446 1388 2447
rect 774 2442 780 2443
rect 110 2431 116 2432
rect 110 2427 111 2431
rect 115 2427 116 2431
rect 110 2426 116 2427
rect 112 2403 114 2426
rect 198 2424 204 2425
rect 198 2420 199 2424
rect 203 2420 204 2424
rect 198 2419 204 2420
rect 200 2403 202 2419
rect 111 2402 115 2403
rect 111 2397 115 2398
rect 135 2402 139 2403
rect 135 2397 139 2398
rect 199 2402 203 2403
rect 199 2397 203 2398
rect 239 2402 243 2403
rect 239 2397 243 2398
rect 112 2390 114 2397
rect 134 2396 140 2397
rect 134 2392 135 2396
rect 139 2392 140 2396
rect 134 2391 140 2392
rect 238 2396 244 2397
rect 238 2392 239 2396
rect 243 2392 244 2396
rect 238 2391 244 2392
rect 110 2389 116 2390
rect 110 2385 111 2389
rect 115 2385 116 2389
rect 110 2384 116 2385
rect 110 2371 116 2372
rect 110 2367 111 2371
rect 115 2367 116 2371
rect 248 2368 250 2442
rect 326 2424 332 2425
rect 326 2420 327 2424
rect 331 2420 332 2424
rect 326 2419 332 2420
rect 454 2424 460 2425
rect 454 2420 455 2424
rect 459 2420 460 2424
rect 454 2419 460 2420
rect 598 2424 604 2425
rect 598 2420 599 2424
rect 603 2420 604 2424
rect 598 2419 604 2420
rect 328 2403 330 2419
rect 456 2403 458 2419
rect 600 2403 602 2419
rect 327 2402 331 2403
rect 327 2397 331 2398
rect 359 2402 363 2403
rect 359 2397 363 2398
rect 455 2402 459 2403
rect 455 2397 459 2398
rect 479 2402 483 2403
rect 479 2397 483 2398
rect 591 2402 595 2403
rect 591 2397 595 2398
rect 599 2402 603 2403
rect 599 2397 603 2398
rect 358 2396 364 2397
rect 358 2392 359 2396
rect 363 2392 364 2396
rect 358 2391 364 2392
rect 478 2396 484 2397
rect 478 2392 479 2396
rect 483 2392 484 2396
rect 478 2391 484 2392
rect 590 2396 596 2397
rect 590 2392 591 2396
rect 595 2392 596 2396
rect 590 2391 596 2392
rect 612 2380 614 2442
rect 766 2424 772 2425
rect 766 2420 767 2424
rect 771 2420 772 2424
rect 766 2419 772 2420
rect 768 2403 770 2419
rect 703 2402 707 2403
rect 703 2397 707 2398
rect 767 2402 771 2403
rect 767 2397 771 2398
rect 702 2396 708 2397
rect 702 2392 703 2396
rect 707 2392 708 2396
rect 702 2391 708 2392
rect 610 2379 616 2380
rect 610 2375 611 2379
rect 615 2375 616 2379
rect 610 2374 616 2375
rect 776 2368 778 2442
rect 950 2424 956 2425
rect 950 2420 951 2424
rect 955 2420 956 2424
rect 950 2419 956 2420
rect 1158 2424 1164 2425
rect 1158 2420 1159 2424
rect 1163 2420 1164 2424
rect 1158 2419 1164 2420
rect 952 2403 954 2419
rect 1160 2403 1162 2419
rect 815 2402 819 2403
rect 815 2397 819 2398
rect 935 2402 939 2403
rect 935 2397 939 2398
rect 951 2402 955 2403
rect 951 2397 955 2398
rect 1159 2402 1163 2403
rect 1159 2397 1163 2398
rect 814 2396 820 2397
rect 814 2392 815 2396
rect 819 2392 820 2396
rect 814 2391 820 2392
rect 934 2396 940 2397
rect 934 2392 935 2396
rect 939 2392 940 2396
rect 934 2391 940 2392
rect 110 2366 116 2367
rect 134 2367 140 2368
rect 112 2355 114 2366
rect 134 2363 135 2367
rect 139 2363 140 2367
rect 134 2362 140 2363
rect 142 2367 148 2368
rect 142 2363 143 2367
rect 147 2363 148 2367
rect 142 2362 148 2363
rect 238 2367 244 2368
rect 238 2363 239 2367
rect 243 2363 244 2367
rect 238 2362 244 2363
rect 246 2367 252 2368
rect 246 2363 247 2367
rect 251 2363 252 2367
rect 246 2362 252 2363
rect 358 2367 364 2368
rect 358 2363 359 2367
rect 363 2363 364 2367
rect 358 2362 364 2363
rect 366 2367 372 2368
rect 366 2363 367 2367
rect 371 2363 372 2367
rect 366 2362 372 2363
rect 478 2367 484 2368
rect 478 2363 479 2367
rect 483 2363 484 2367
rect 478 2362 484 2363
rect 574 2367 580 2368
rect 574 2363 575 2367
rect 579 2363 580 2367
rect 574 2362 580 2363
rect 590 2367 596 2368
rect 590 2363 591 2367
rect 595 2363 596 2367
rect 590 2362 596 2363
rect 702 2367 708 2368
rect 702 2363 703 2367
rect 707 2363 708 2367
rect 702 2362 708 2363
rect 774 2367 780 2368
rect 774 2363 775 2367
rect 779 2363 780 2367
rect 774 2362 780 2363
rect 814 2367 820 2368
rect 814 2363 815 2367
rect 819 2363 820 2367
rect 814 2362 820 2363
rect 934 2367 940 2368
rect 934 2363 935 2367
rect 939 2363 940 2367
rect 934 2362 940 2363
rect 942 2367 948 2368
rect 942 2363 943 2367
rect 947 2363 948 2367
rect 942 2362 948 2363
rect 982 2367 988 2368
rect 982 2363 983 2367
rect 987 2363 988 2367
rect 982 2362 988 2363
rect 136 2355 138 2362
rect 111 2354 115 2355
rect 135 2354 139 2355
rect 111 2349 115 2350
rect 134 2349 140 2350
rect 112 2346 114 2349
rect 110 2345 116 2346
rect 110 2341 111 2345
rect 115 2341 116 2345
rect 134 2345 135 2349
rect 139 2345 140 2349
rect 134 2344 140 2345
rect 144 2344 146 2362
rect 240 2355 242 2362
rect 239 2354 243 2355
rect 239 2349 243 2350
rect 248 2344 250 2362
rect 360 2355 362 2362
rect 343 2354 347 2355
rect 359 2354 363 2355
rect 342 2349 348 2350
rect 359 2349 363 2350
rect 342 2345 343 2349
rect 347 2345 348 2349
rect 342 2344 348 2345
rect 368 2344 370 2362
rect 480 2355 482 2362
rect 479 2354 483 2355
rect 567 2354 571 2355
rect 479 2349 483 2350
rect 566 2349 572 2350
rect 566 2345 567 2349
rect 571 2345 572 2349
rect 566 2344 572 2345
rect 576 2344 578 2362
rect 592 2355 594 2362
rect 704 2355 706 2362
rect 790 2359 796 2360
rect 790 2355 791 2359
rect 795 2355 796 2359
rect 816 2355 818 2362
rect 936 2355 938 2362
rect 591 2354 595 2355
rect 591 2349 595 2350
rect 703 2354 707 2355
rect 775 2354 779 2355
rect 790 2354 796 2355
rect 815 2354 819 2355
rect 703 2349 707 2350
rect 774 2349 780 2350
rect 774 2345 775 2349
rect 779 2345 780 2349
rect 774 2344 780 2345
rect 110 2340 116 2341
rect 142 2343 148 2344
rect 142 2339 143 2343
rect 147 2339 148 2343
rect 142 2338 148 2339
rect 182 2343 188 2344
rect 182 2339 183 2343
rect 187 2339 188 2343
rect 182 2338 188 2339
rect 246 2343 252 2344
rect 246 2339 247 2343
rect 251 2339 252 2343
rect 246 2338 252 2339
rect 366 2343 372 2344
rect 366 2339 367 2343
rect 371 2339 372 2343
rect 366 2338 372 2339
rect 574 2343 580 2344
rect 574 2339 575 2343
rect 579 2339 580 2343
rect 574 2338 580 2339
rect 782 2343 788 2344
rect 782 2339 783 2343
rect 787 2339 788 2343
rect 792 2339 794 2354
rect 815 2349 819 2350
rect 935 2354 939 2355
rect 935 2349 939 2350
rect 782 2338 794 2339
rect 110 2327 116 2328
rect 110 2323 111 2327
rect 115 2323 116 2327
rect 110 2322 116 2323
rect 112 2303 114 2322
rect 134 2320 140 2321
rect 134 2316 135 2320
rect 139 2316 140 2320
rect 134 2315 140 2316
rect 136 2303 138 2315
rect 111 2302 115 2303
rect 111 2297 115 2298
rect 135 2302 139 2303
rect 135 2297 139 2298
rect 112 2290 114 2297
rect 110 2289 116 2290
rect 110 2285 111 2289
rect 115 2285 116 2289
rect 110 2284 116 2285
rect 110 2271 116 2272
rect 110 2267 111 2271
rect 115 2267 116 2271
rect 110 2266 116 2267
rect 112 2251 114 2266
rect 111 2250 115 2251
rect 111 2245 115 2246
rect 112 2242 114 2245
rect 110 2241 116 2242
rect 110 2237 111 2241
rect 115 2237 116 2241
rect 110 2236 116 2237
rect 110 2223 116 2224
rect 110 2219 111 2223
rect 115 2219 116 2223
rect 110 2218 116 2219
rect 112 2203 114 2218
rect 111 2202 115 2203
rect 111 2197 115 2198
rect 112 2190 114 2197
rect 110 2189 116 2190
rect 110 2185 111 2189
rect 115 2185 116 2189
rect 110 2184 116 2185
rect 110 2171 116 2172
rect 110 2167 111 2171
rect 115 2167 116 2171
rect 110 2166 116 2167
rect 112 2151 114 2166
rect 111 2150 115 2151
rect 111 2145 115 2146
rect 112 2142 114 2145
rect 110 2141 116 2142
rect 110 2137 111 2141
rect 115 2137 116 2141
rect 110 2136 116 2137
rect 110 2123 116 2124
rect 110 2119 111 2123
rect 115 2119 116 2123
rect 110 2118 116 2119
rect 112 2099 114 2118
rect 111 2098 115 2099
rect 111 2093 115 2094
rect 112 2086 114 2093
rect 110 2085 116 2086
rect 110 2081 111 2085
rect 115 2081 116 2085
rect 110 2080 116 2081
rect 110 2067 116 2068
rect 110 2063 111 2067
rect 115 2063 116 2067
rect 110 2062 116 2063
rect 112 2051 114 2062
rect 111 2050 115 2051
rect 175 2050 179 2051
rect 111 2045 115 2046
rect 174 2045 180 2046
rect 112 2042 114 2045
rect 110 2041 116 2042
rect 110 2037 111 2041
rect 115 2037 116 2041
rect 174 2041 175 2045
rect 179 2041 180 2045
rect 174 2040 180 2041
rect 184 2040 186 2338
rect 342 2320 348 2321
rect 342 2316 343 2320
rect 347 2316 348 2320
rect 342 2315 348 2316
rect 566 2320 572 2321
rect 566 2316 567 2320
rect 571 2316 572 2320
rect 566 2315 572 2316
rect 344 2303 346 2315
rect 568 2303 570 2315
rect 343 2302 347 2303
rect 343 2297 347 2298
rect 567 2302 571 2303
rect 567 2297 571 2298
rect 551 2250 555 2251
rect 550 2245 556 2246
rect 550 2241 551 2245
rect 555 2241 556 2245
rect 550 2240 556 2241
rect 576 2240 578 2338
rect 784 2337 794 2338
rect 774 2320 780 2321
rect 774 2316 775 2320
rect 779 2316 780 2320
rect 774 2315 780 2316
rect 776 2303 778 2315
rect 655 2302 659 2303
rect 655 2297 659 2298
rect 775 2302 779 2303
rect 775 2297 779 2298
rect 783 2302 787 2303
rect 783 2297 787 2298
rect 654 2296 660 2297
rect 654 2292 655 2296
rect 659 2292 660 2296
rect 654 2291 660 2292
rect 782 2296 788 2297
rect 782 2292 783 2296
rect 787 2292 788 2296
rect 782 2291 788 2292
rect 792 2268 794 2337
rect 903 2302 907 2303
rect 903 2297 907 2298
rect 902 2296 908 2297
rect 902 2292 903 2296
rect 907 2292 908 2296
rect 902 2291 908 2292
rect 944 2272 946 2362
rect 975 2354 979 2355
rect 974 2349 980 2350
rect 974 2345 975 2349
rect 979 2345 980 2349
rect 984 2348 986 2362
rect 1175 2354 1179 2355
rect 1174 2349 1180 2350
rect 974 2344 980 2345
rect 982 2347 988 2348
rect 982 2343 983 2347
rect 987 2343 988 2347
rect 1174 2345 1175 2349
rect 1179 2345 1180 2349
rect 1174 2344 1180 2345
rect 1184 2344 1186 2446
rect 1374 2424 1380 2425
rect 1374 2420 1375 2424
rect 1379 2420 1380 2424
rect 1374 2419 1380 2420
rect 1376 2403 1378 2419
rect 1375 2402 1379 2403
rect 1375 2397 1379 2398
rect 1384 2355 1386 2446
rect 1367 2354 1371 2355
rect 1376 2353 1386 2355
rect 1567 2354 1571 2355
rect 1366 2349 1372 2350
rect 1366 2345 1367 2349
rect 1371 2345 1372 2349
rect 1376 2348 1378 2353
rect 1566 2349 1572 2350
rect 1366 2344 1372 2345
rect 1374 2347 1380 2348
rect 982 2342 988 2343
rect 1166 2343 1172 2344
rect 1166 2339 1167 2343
rect 1171 2339 1172 2343
rect 1166 2338 1172 2339
rect 1182 2343 1188 2344
rect 1182 2339 1183 2343
rect 1187 2339 1188 2343
rect 1374 2343 1375 2347
rect 1379 2343 1380 2347
rect 1566 2345 1567 2349
rect 1571 2345 1572 2349
rect 1576 2348 1578 2470
rect 1598 2467 1604 2468
rect 1598 2463 1599 2467
rect 1603 2463 1604 2467
rect 1630 2467 1631 2471
rect 1635 2467 1636 2471
rect 1671 2469 1675 2470
rect 1695 2474 1699 2475
rect 1695 2469 1699 2470
rect 1863 2474 1867 2475
rect 1863 2469 1867 2470
rect 2079 2474 2083 2475
rect 2079 2469 2083 2470
rect 2319 2474 2323 2475
rect 2319 2469 2323 2470
rect 1630 2466 1636 2467
rect 1598 2462 1604 2463
rect 1600 2459 1602 2462
rect 1632 2459 1634 2466
rect 1672 2462 1674 2469
rect 2318 2468 2324 2469
rect 2318 2464 2319 2468
rect 2323 2464 2324 2468
rect 2318 2463 2324 2464
rect 1670 2461 1676 2462
rect 1591 2458 1595 2459
rect 1599 2458 1603 2459
rect 1590 2453 1596 2454
rect 1599 2453 1603 2454
rect 1631 2458 1635 2459
rect 1670 2457 1671 2461
rect 1675 2457 1676 2461
rect 1670 2456 1676 2457
rect 1631 2453 1635 2454
rect 1590 2449 1591 2453
rect 1595 2449 1596 2453
rect 1632 2450 1634 2453
rect 1590 2448 1596 2449
rect 1630 2449 1636 2450
rect 1630 2445 1631 2449
rect 1635 2445 1636 2449
rect 1630 2444 1636 2445
rect 2328 2444 2330 2510
rect 2567 2474 2571 2475
rect 2567 2469 2571 2470
rect 2566 2468 2572 2469
rect 2566 2464 2567 2468
rect 2571 2464 2572 2468
rect 2566 2463 2572 2464
rect 2576 2444 2578 2518
rect 2582 2517 2588 2518
rect 2582 2513 2583 2517
rect 2587 2513 2588 2517
rect 2582 2512 2588 2513
rect 2854 2517 2860 2518
rect 2854 2513 2855 2517
rect 2859 2513 2860 2517
rect 2854 2512 2860 2513
rect 2928 2512 2930 2594
rect 3135 2522 3139 2523
rect 3134 2517 3140 2518
rect 3134 2513 3135 2517
rect 3139 2513 3140 2517
rect 3134 2512 3140 2513
rect 3144 2512 3146 2594
rect 3190 2583 3196 2584
rect 3190 2579 3191 2583
rect 3195 2579 3196 2583
rect 3190 2578 3196 2579
rect 3158 2576 3164 2577
rect 3158 2572 3159 2576
rect 3163 2572 3164 2576
rect 3158 2571 3164 2572
rect 3160 2567 3162 2571
rect 3192 2567 3194 2578
rect 3159 2566 3163 2567
rect 3159 2561 3163 2562
rect 3191 2566 3195 2567
rect 3191 2561 3195 2562
rect 3192 2554 3194 2561
rect 3190 2553 3196 2554
rect 3190 2549 3191 2553
rect 3195 2549 3196 2553
rect 3190 2548 3196 2549
rect 3190 2535 3196 2536
rect 3190 2531 3191 2535
rect 3195 2531 3196 2535
rect 3190 2530 3196 2531
rect 3192 2523 3194 2530
rect 3191 2522 3195 2523
rect 3191 2517 3195 2518
rect 3192 2514 3194 2517
rect 3190 2513 3196 2514
rect 2862 2511 2868 2512
rect 2862 2507 2863 2511
rect 2867 2507 2868 2511
rect 2862 2506 2868 2507
rect 2926 2511 2932 2512
rect 2926 2507 2927 2511
rect 2931 2507 2932 2511
rect 2926 2506 2932 2507
rect 2974 2511 2980 2512
rect 2974 2507 2975 2511
rect 2979 2507 2980 2511
rect 2974 2506 2980 2507
rect 3142 2511 3148 2512
rect 3142 2507 3143 2511
rect 3147 2507 3148 2511
rect 3190 2509 3191 2513
rect 3195 2509 3196 2513
rect 3190 2508 3196 2509
rect 3142 2506 3148 2507
rect 2582 2488 2588 2489
rect 2582 2484 2583 2488
rect 2587 2484 2588 2488
rect 2582 2483 2588 2484
rect 2854 2488 2860 2489
rect 2854 2484 2855 2488
rect 2859 2484 2860 2488
rect 2854 2483 2860 2484
rect 2584 2475 2586 2483
rect 2856 2475 2858 2483
rect 2583 2474 2587 2475
rect 2583 2469 2587 2470
rect 2823 2474 2827 2475
rect 2823 2469 2827 2470
rect 2855 2474 2859 2475
rect 2855 2469 2859 2470
rect 2822 2468 2828 2469
rect 2822 2464 2823 2468
rect 2827 2464 2828 2468
rect 2822 2463 2828 2464
rect 2864 2444 2866 2506
rect 1670 2443 1676 2444
rect 1670 2439 1671 2443
rect 1675 2439 1676 2443
rect 2326 2443 2332 2444
rect 1670 2438 1676 2439
rect 2318 2439 2324 2440
rect 1672 2435 1674 2438
rect 2318 2435 2319 2439
rect 2323 2435 2324 2439
rect 2326 2439 2327 2443
rect 2331 2439 2332 2443
rect 2574 2443 2580 2444
rect 2326 2438 2332 2439
rect 2566 2439 2572 2440
rect 1671 2434 1675 2435
rect 1630 2431 1636 2432
rect 1630 2427 1631 2431
rect 1635 2427 1636 2431
rect 2231 2434 2235 2435
rect 2318 2434 2324 2435
rect 1671 2429 1675 2430
rect 2230 2429 2236 2430
rect 2319 2429 2323 2430
rect 1630 2426 1636 2427
rect 1672 2426 1674 2429
rect 1590 2424 1596 2425
rect 1590 2420 1591 2424
rect 1595 2420 1596 2424
rect 1590 2419 1596 2420
rect 1592 2403 1594 2419
rect 1632 2403 1634 2426
rect 1670 2425 1676 2426
rect 1670 2421 1671 2425
rect 1675 2421 1676 2425
rect 2230 2425 2231 2429
rect 2235 2425 2236 2429
rect 2328 2428 2330 2438
rect 2566 2435 2567 2439
rect 2571 2435 2572 2439
rect 2574 2439 2575 2443
rect 2579 2439 2580 2443
rect 2862 2443 2868 2444
rect 2574 2438 2580 2439
rect 2822 2439 2828 2440
rect 2391 2434 2395 2435
rect 2543 2434 2547 2435
rect 2566 2434 2572 2435
rect 2390 2429 2396 2430
rect 2230 2424 2236 2425
rect 2238 2427 2244 2428
rect 2238 2423 2239 2427
rect 2243 2423 2244 2427
rect 2238 2422 2244 2423
rect 2326 2427 2332 2428
rect 2326 2423 2327 2427
rect 2331 2423 2332 2427
rect 2326 2422 2332 2423
rect 2342 2427 2348 2428
rect 2342 2423 2343 2427
rect 2347 2423 2348 2427
rect 2390 2425 2391 2429
rect 2395 2425 2396 2429
rect 2390 2424 2396 2425
rect 2542 2429 2548 2430
rect 2567 2429 2571 2430
rect 2542 2425 2543 2429
rect 2547 2425 2548 2429
rect 2576 2428 2578 2438
rect 2822 2435 2823 2439
rect 2827 2435 2828 2439
rect 2862 2439 2863 2443
rect 2867 2439 2868 2443
rect 2862 2438 2868 2439
rect 2687 2434 2691 2435
rect 2822 2434 2828 2435
rect 2967 2434 2971 2435
rect 2686 2429 2692 2430
rect 2542 2424 2548 2425
rect 2574 2427 2580 2428
rect 2342 2422 2348 2423
rect 2574 2423 2575 2427
rect 2579 2423 2580 2427
rect 2686 2425 2687 2429
rect 2691 2425 2692 2429
rect 2686 2424 2692 2425
rect 2822 2429 2828 2430
rect 2822 2425 2823 2429
rect 2827 2425 2828 2429
rect 2822 2424 2828 2425
rect 2966 2429 2972 2430
rect 2966 2425 2967 2429
rect 2971 2425 2972 2429
rect 2966 2424 2972 2425
rect 2976 2424 2978 2506
rect 3134 2488 3140 2489
rect 3134 2484 3135 2488
rect 3139 2484 3140 2488
rect 3134 2483 3140 2484
rect 3136 2475 3138 2483
rect 3079 2474 3083 2475
rect 3079 2469 3083 2470
rect 3135 2474 3139 2475
rect 3135 2469 3139 2470
rect 3078 2468 3084 2469
rect 3078 2464 3079 2468
rect 3083 2464 3084 2468
rect 3078 2463 3084 2464
rect 3078 2439 3084 2440
rect 3078 2435 3079 2439
rect 3083 2435 3084 2439
rect 3078 2434 3084 2435
rect 3111 2434 3115 2435
rect 3079 2429 3083 2430
rect 3110 2429 3116 2430
rect 3110 2425 3111 2429
rect 3115 2425 3116 2429
rect 3110 2424 3116 2425
rect 3144 2424 3146 2506
rect 3190 2495 3196 2496
rect 3190 2491 3191 2495
rect 3195 2491 3196 2495
rect 3190 2490 3196 2491
rect 3192 2475 3194 2490
rect 3191 2474 3195 2475
rect 3191 2469 3195 2470
rect 3192 2462 3194 2469
rect 3190 2461 3196 2462
rect 3190 2457 3191 2461
rect 3195 2457 3196 2461
rect 3190 2456 3196 2457
rect 3190 2443 3196 2444
rect 3190 2439 3191 2443
rect 3195 2439 3196 2443
rect 3190 2438 3196 2439
rect 3192 2435 3194 2438
rect 3191 2434 3195 2435
rect 3191 2429 3195 2430
rect 3192 2426 3194 2429
rect 3190 2425 3196 2426
rect 2574 2422 2580 2423
rect 2666 2423 2672 2424
rect 1670 2420 1676 2421
rect 1670 2407 1676 2408
rect 1670 2403 1671 2407
rect 1675 2403 1676 2407
rect 1591 2402 1595 2403
rect 1591 2397 1595 2398
rect 1631 2402 1635 2403
rect 1670 2402 1676 2403
rect 1631 2397 1635 2398
rect 1632 2390 1634 2397
rect 1630 2389 1636 2390
rect 1630 2385 1631 2389
rect 1635 2385 1636 2389
rect 1672 2387 1674 2402
rect 2230 2400 2236 2401
rect 2230 2396 2231 2400
rect 2235 2396 2236 2400
rect 2230 2395 2236 2396
rect 2232 2387 2234 2395
rect 1630 2384 1636 2385
rect 1671 2386 1675 2387
rect 1671 2381 1675 2382
rect 2143 2386 2147 2387
rect 2143 2381 2147 2382
rect 2231 2386 2235 2387
rect 2231 2381 2235 2382
rect 1672 2374 1674 2381
rect 2142 2380 2148 2381
rect 2142 2376 2143 2380
rect 2147 2376 2148 2380
rect 2142 2375 2148 2376
rect 1670 2373 1676 2374
rect 1630 2371 1636 2372
rect 1630 2367 1631 2371
rect 1635 2367 1636 2371
rect 1670 2369 1671 2373
rect 1675 2369 1676 2373
rect 1670 2368 1676 2369
rect 1630 2366 1636 2367
rect 1632 2355 1634 2366
rect 2240 2356 2242 2422
rect 2311 2386 2315 2387
rect 2311 2381 2315 2382
rect 2310 2380 2316 2381
rect 2310 2376 2311 2380
rect 2315 2376 2316 2380
rect 2310 2375 2316 2376
rect 2344 2356 2346 2422
rect 2666 2419 2667 2423
rect 2671 2419 2672 2423
rect 2666 2418 2672 2419
rect 2974 2423 2980 2424
rect 2974 2419 2975 2423
rect 2979 2419 2980 2423
rect 2974 2418 2980 2419
rect 3014 2423 3020 2424
rect 3014 2419 3015 2423
rect 3019 2419 3020 2423
rect 3014 2418 3020 2419
rect 3142 2423 3148 2424
rect 3142 2419 3143 2423
rect 3147 2419 3148 2423
rect 3142 2418 3148 2419
rect 3166 2423 3172 2424
rect 3166 2419 3167 2423
rect 3171 2419 3172 2423
rect 3190 2421 3191 2425
rect 3195 2421 3196 2425
rect 3190 2420 3196 2421
rect 3166 2418 3172 2419
rect 2390 2400 2396 2401
rect 2390 2396 2391 2400
rect 2395 2396 2396 2400
rect 2390 2395 2396 2396
rect 2542 2400 2548 2401
rect 2542 2396 2543 2400
rect 2547 2396 2548 2400
rect 2542 2395 2548 2396
rect 2392 2387 2394 2395
rect 2544 2387 2546 2395
rect 2391 2386 2395 2387
rect 2391 2381 2395 2382
rect 2479 2386 2483 2387
rect 2479 2381 2483 2382
rect 2543 2386 2547 2387
rect 2543 2381 2547 2382
rect 2655 2386 2659 2387
rect 2655 2381 2659 2382
rect 2478 2380 2484 2381
rect 2478 2376 2479 2380
rect 2483 2376 2484 2380
rect 2478 2375 2484 2376
rect 2654 2380 2660 2381
rect 2654 2376 2655 2380
rect 2659 2376 2660 2380
rect 2654 2375 2660 2376
rect 2668 2356 2670 2418
rect 2686 2400 2692 2401
rect 2686 2396 2687 2400
rect 2691 2396 2692 2400
rect 2686 2395 2692 2396
rect 2822 2400 2828 2401
rect 2822 2396 2823 2400
rect 2827 2396 2828 2400
rect 2822 2395 2828 2396
rect 2966 2400 2972 2401
rect 2966 2396 2967 2400
rect 2971 2396 2972 2400
rect 2966 2395 2972 2396
rect 2688 2387 2690 2395
rect 2824 2387 2826 2395
rect 2968 2387 2970 2395
rect 2687 2386 2691 2387
rect 2687 2381 2691 2382
rect 2823 2386 2827 2387
rect 2823 2381 2827 2382
rect 2831 2386 2835 2387
rect 2831 2381 2835 2382
rect 2967 2386 2971 2387
rect 2967 2381 2971 2382
rect 3007 2386 3011 2387
rect 3007 2381 3011 2382
rect 2830 2380 2836 2381
rect 2830 2376 2831 2380
rect 2835 2376 2836 2380
rect 2830 2375 2836 2376
rect 3006 2380 3012 2381
rect 3006 2376 3007 2380
rect 3011 2376 3012 2380
rect 3006 2375 3012 2376
rect 3016 2356 3018 2418
rect 3110 2400 3116 2401
rect 3110 2396 3111 2400
rect 3115 2396 3116 2400
rect 3110 2395 3116 2396
rect 3112 2387 3114 2395
rect 3111 2386 3115 2387
rect 3111 2381 3115 2382
rect 3159 2386 3163 2387
rect 3159 2381 3163 2382
rect 3158 2380 3164 2381
rect 3158 2376 3159 2380
rect 3163 2376 3164 2380
rect 3158 2375 3164 2376
rect 3168 2360 3170 2418
rect 3190 2407 3196 2408
rect 3190 2403 3191 2407
rect 3195 2403 3196 2407
rect 3190 2402 3196 2403
rect 3192 2387 3194 2402
rect 3191 2386 3195 2387
rect 3191 2381 3195 2382
rect 3192 2374 3194 2381
rect 3190 2373 3196 2374
rect 3190 2369 3191 2373
rect 3195 2369 3196 2373
rect 3190 2368 3196 2369
rect 3166 2359 3172 2360
rect 1670 2355 1676 2356
rect 1631 2354 1635 2355
rect 1670 2351 1671 2355
rect 1675 2351 1676 2355
rect 2238 2355 2244 2356
rect 1670 2350 1676 2351
rect 2142 2351 2148 2352
rect 1631 2349 1635 2350
rect 1566 2344 1572 2345
rect 1574 2347 1580 2348
rect 1374 2342 1380 2343
rect 1574 2343 1575 2347
rect 1579 2343 1580 2347
rect 1632 2346 1634 2349
rect 1672 2347 1674 2350
rect 2142 2347 2143 2351
rect 2147 2347 2148 2351
rect 1671 2346 1675 2347
rect 2142 2346 2148 2347
rect 2174 2351 2180 2352
rect 2174 2347 2175 2351
rect 2179 2347 2180 2351
rect 2238 2351 2239 2355
rect 2243 2351 2244 2355
rect 2342 2355 2348 2356
rect 2238 2350 2244 2351
rect 2310 2351 2316 2352
rect 2310 2347 2311 2351
rect 2315 2347 2316 2351
rect 2342 2351 2343 2355
rect 2347 2351 2348 2355
rect 2666 2355 2672 2356
rect 2342 2350 2348 2351
rect 2478 2351 2484 2352
rect 2174 2346 2180 2347
rect 2183 2346 2187 2347
rect 2310 2346 2316 2347
rect 2335 2346 2339 2347
rect 1574 2342 1580 2343
rect 1630 2345 1636 2346
rect 1182 2338 1188 2339
rect 974 2320 980 2321
rect 974 2316 975 2320
rect 979 2316 980 2320
rect 974 2315 980 2316
rect 976 2303 978 2315
rect 975 2302 979 2303
rect 975 2297 979 2298
rect 1023 2302 1027 2303
rect 1023 2297 1027 2298
rect 1143 2302 1147 2303
rect 1143 2297 1147 2298
rect 1022 2296 1028 2297
rect 1022 2292 1023 2296
rect 1027 2292 1028 2296
rect 1022 2291 1028 2292
rect 1142 2296 1148 2297
rect 1142 2292 1143 2296
rect 1147 2292 1148 2296
rect 1142 2291 1148 2292
rect 1168 2272 1170 2338
rect 1174 2320 1180 2321
rect 1174 2316 1175 2320
rect 1179 2316 1180 2320
rect 1174 2315 1180 2316
rect 1366 2320 1372 2321
rect 1366 2316 1367 2320
rect 1371 2316 1372 2320
rect 1366 2315 1372 2316
rect 1176 2303 1178 2315
rect 1368 2303 1370 2315
rect 1175 2302 1179 2303
rect 1175 2297 1179 2298
rect 1255 2302 1259 2303
rect 1255 2297 1259 2298
rect 1367 2302 1371 2303
rect 1367 2297 1371 2298
rect 1254 2296 1260 2297
rect 1254 2292 1255 2296
rect 1259 2292 1260 2296
rect 1254 2291 1260 2292
rect 1366 2296 1372 2297
rect 1366 2292 1367 2296
rect 1371 2292 1372 2296
rect 1366 2291 1372 2292
rect 942 2271 948 2272
rect 654 2267 660 2268
rect 654 2263 655 2267
rect 659 2263 660 2267
rect 654 2262 660 2263
rect 662 2267 668 2268
rect 662 2263 663 2267
rect 667 2263 668 2267
rect 662 2262 668 2263
rect 782 2267 788 2268
rect 782 2263 783 2267
rect 787 2263 788 2267
rect 782 2262 788 2263
rect 790 2267 796 2268
rect 790 2263 791 2267
rect 795 2263 796 2267
rect 790 2262 796 2263
rect 814 2267 820 2268
rect 814 2263 815 2267
rect 819 2263 820 2267
rect 814 2262 820 2263
rect 902 2267 908 2268
rect 902 2263 903 2267
rect 907 2263 908 2267
rect 942 2267 943 2271
rect 947 2267 948 2271
rect 942 2266 948 2267
rect 950 2271 956 2272
rect 950 2267 951 2271
rect 955 2267 956 2271
rect 1054 2271 1060 2272
rect 950 2266 956 2267
rect 1022 2267 1028 2268
rect 902 2262 908 2263
rect 656 2251 658 2262
rect 655 2250 659 2251
rect 655 2245 659 2246
rect 664 2240 666 2262
rect 784 2251 786 2262
rect 679 2250 683 2251
rect 783 2250 787 2251
rect 807 2250 811 2251
rect 678 2245 684 2246
rect 783 2245 787 2246
rect 806 2245 812 2246
rect 678 2241 679 2245
rect 683 2241 684 2245
rect 678 2240 684 2241
rect 806 2241 807 2245
rect 811 2241 812 2245
rect 816 2244 818 2262
rect 904 2251 906 2262
rect 903 2250 907 2251
rect 927 2250 931 2251
rect 903 2245 907 2246
rect 926 2245 932 2246
rect 806 2240 812 2241
rect 814 2243 820 2244
rect 574 2239 580 2240
rect 574 2235 575 2239
rect 579 2235 580 2239
rect 574 2234 580 2235
rect 606 2239 612 2240
rect 606 2235 607 2239
rect 611 2235 612 2239
rect 606 2234 612 2235
rect 662 2239 668 2240
rect 662 2235 663 2239
rect 667 2235 668 2239
rect 814 2239 815 2243
rect 819 2239 820 2243
rect 926 2241 927 2245
rect 931 2241 932 2245
rect 926 2240 932 2241
rect 952 2240 954 2266
rect 1022 2263 1023 2267
rect 1027 2263 1028 2267
rect 1054 2267 1055 2271
rect 1059 2267 1060 2271
rect 1166 2271 1172 2272
rect 1054 2266 1060 2267
rect 1142 2267 1148 2268
rect 1022 2262 1028 2263
rect 1024 2251 1026 2262
rect 1023 2250 1027 2251
rect 1047 2250 1051 2251
rect 1056 2248 1058 2266
rect 1142 2263 1143 2267
rect 1147 2263 1148 2267
rect 1166 2267 1167 2271
rect 1171 2267 1172 2271
rect 1278 2271 1284 2272
rect 1166 2266 1172 2267
rect 1254 2267 1260 2268
rect 1142 2262 1148 2263
rect 1144 2251 1146 2262
rect 1143 2250 1147 2251
rect 1054 2247 1060 2248
rect 1023 2245 1027 2246
rect 1046 2245 1052 2246
rect 1046 2241 1047 2245
rect 1051 2241 1052 2245
rect 1054 2243 1055 2247
rect 1059 2243 1060 2247
rect 1159 2250 1163 2251
rect 1168 2248 1170 2266
rect 1254 2263 1255 2267
rect 1259 2263 1260 2267
rect 1278 2267 1279 2271
rect 1283 2267 1284 2271
rect 1376 2268 1378 2342
rect 1630 2341 1631 2345
rect 1635 2341 1636 2345
rect 1671 2341 1675 2342
rect 2143 2341 2147 2342
rect 1630 2340 1636 2341
rect 1672 2338 1674 2341
rect 1670 2337 1676 2338
rect 1670 2333 1671 2337
rect 1675 2333 1676 2337
rect 2176 2336 2178 2346
rect 2182 2341 2188 2342
rect 2311 2341 2315 2342
rect 2334 2341 2340 2342
rect 2182 2337 2183 2341
rect 2187 2337 2188 2341
rect 2182 2336 2188 2337
rect 2334 2337 2335 2341
rect 2339 2337 2340 2341
rect 2344 2340 2346 2350
rect 2478 2347 2479 2351
rect 2483 2347 2484 2351
rect 2654 2351 2660 2352
rect 2654 2347 2655 2351
rect 2659 2347 2660 2351
rect 2666 2351 2667 2355
rect 2671 2351 2672 2355
rect 3014 2355 3020 2356
rect 2666 2350 2672 2351
rect 2830 2351 2836 2352
rect 2478 2346 2484 2347
rect 2623 2346 2627 2347
rect 2654 2346 2660 2347
rect 2478 2341 2484 2342
rect 2334 2336 2340 2337
rect 2342 2339 2348 2340
rect 1670 2332 1676 2333
rect 2174 2335 2180 2336
rect 2174 2331 2175 2335
rect 2179 2331 2180 2335
rect 2342 2335 2343 2339
rect 2347 2335 2348 2339
rect 2478 2337 2479 2341
rect 2483 2337 2484 2341
rect 2478 2336 2484 2337
rect 2622 2341 2628 2342
rect 2655 2341 2659 2342
rect 2622 2337 2623 2341
rect 2627 2337 2628 2341
rect 2668 2340 2670 2350
rect 2830 2347 2831 2351
rect 2835 2347 2836 2351
rect 3006 2351 3012 2352
rect 3006 2347 3007 2351
rect 3011 2347 3012 2351
rect 3014 2351 3015 2355
rect 3019 2351 3020 2355
rect 3166 2355 3167 2359
rect 3171 2355 3172 2359
rect 3166 2354 3172 2355
rect 3190 2355 3196 2356
rect 3168 2352 3170 2354
rect 3014 2350 3020 2351
rect 3158 2351 3164 2352
rect 2767 2346 2771 2347
rect 2830 2346 2836 2347
rect 2919 2346 2923 2347
rect 3006 2346 3012 2347
rect 2766 2341 2772 2342
rect 2831 2341 2835 2342
rect 2918 2341 2924 2342
rect 3007 2341 3011 2342
rect 2622 2336 2628 2337
rect 2630 2339 2636 2340
rect 2342 2334 2348 2335
rect 2486 2335 2492 2336
rect 2174 2330 2180 2331
rect 2486 2331 2487 2335
rect 2491 2331 2492 2335
rect 2630 2335 2631 2339
rect 2635 2335 2636 2339
rect 2630 2334 2636 2335
rect 2666 2339 2672 2340
rect 2666 2335 2667 2339
rect 2671 2335 2672 2339
rect 2766 2337 2767 2341
rect 2771 2337 2772 2341
rect 2766 2336 2772 2337
rect 2798 2339 2804 2340
rect 2666 2334 2672 2335
rect 2798 2335 2799 2339
rect 2803 2335 2804 2339
rect 2918 2337 2919 2341
rect 2923 2337 2924 2341
rect 3016 2340 3018 2350
rect 3158 2347 3159 2351
rect 3163 2347 3164 2351
rect 3158 2346 3164 2347
rect 3166 2351 3172 2352
rect 3166 2347 3167 2351
rect 3171 2347 3172 2351
rect 3190 2351 3191 2355
rect 3195 2351 3196 2355
rect 3190 2350 3196 2351
rect 3192 2347 3194 2350
rect 3166 2346 3172 2347
rect 3191 2346 3195 2347
rect 3159 2341 3163 2342
rect 2918 2336 2924 2337
rect 3014 2339 3020 2340
rect 2798 2334 2804 2335
rect 3014 2335 3015 2339
rect 3019 2335 3020 2339
rect 3014 2334 3020 2335
rect 2486 2330 2492 2331
rect 1630 2327 1636 2328
rect 1630 2323 1631 2327
rect 1635 2323 1636 2327
rect 1630 2322 1636 2323
rect 1566 2320 1572 2321
rect 1566 2316 1567 2320
rect 1571 2316 1572 2320
rect 1566 2315 1572 2316
rect 1568 2303 1570 2315
rect 1632 2303 1634 2322
rect 1670 2319 1676 2320
rect 1670 2315 1671 2319
rect 1675 2315 1676 2319
rect 1670 2314 1676 2315
rect 1672 2303 1674 2314
rect 1487 2302 1491 2303
rect 1487 2297 1491 2298
rect 1567 2302 1571 2303
rect 1567 2297 1571 2298
rect 1631 2302 1635 2303
rect 1631 2297 1635 2298
rect 1671 2302 1675 2303
rect 1671 2297 1675 2298
rect 2095 2302 2099 2303
rect 2095 2297 2099 2298
rect 1486 2296 1492 2297
rect 1486 2292 1487 2296
rect 1491 2292 1492 2296
rect 1486 2291 1492 2292
rect 1632 2290 1634 2297
rect 1672 2290 1674 2297
rect 2094 2296 2100 2297
rect 2094 2292 2095 2296
rect 2099 2292 2100 2296
rect 2094 2291 2100 2292
rect 1630 2289 1636 2290
rect 1630 2285 1631 2289
rect 1635 2285 1636 2289
rect 1630 2284 1636 2285
rect 1670 2289 1676 2290
rect 1670 2285 1671 2289
rect 1675 2285 1676 2289
rect 1670 2284 1676 2285
rect 1398 2275 1404 2276
rect 1398 2271 1399 2275
rect 1403 2271 1404 2275
rect 2022 2275 2028 2276
rect 1398 2270 1404 2271
rect 1630 2271 1636 2272
rect 1278 2266 1284 2267
rect 1366 2267 1372 2268
rect 1254 2262 1260 2263
rect 1256 2251 1258 2262
rect 1255 2250 1259 2251
rect 1166 2247 1172 2248
rect 1143 2245 1147 2246
rect 1158 2245 1164 2246
rect 1054 2242 1060 2243
rect 1046 2240 1052 2241
rect 1158 2241 1159 2245
rect 1163 2241 1164 2245
rect 1166 2243 1167 2247
rect 1171 2243 1172 2247
rect 1271 2250 1275 2251
rect 1255 2245 1259 2246
rect 1270 2245 1276 2246
rect 1166 2242 1172 2243
rect 1158 2240 1164 2241
rect 814 2238 820 2239
rect 950 2239 956 2240
rect 662 2234 668 2235
rect 950 2235 951 2239
rect 955 2235 956 2239
rect 950 2234 956 2235
rect 550 2216 556 2217
rect 550 2212 551 2216
rect 555 2212 556 2216
rect 550 2211 556 2212
rect 552 2203 554 2211
rect 455 2202 459 2203
rect 455 2197 459 2198
rect 551 2202 555 2203
rect 551 2197 555 2198
rect 583 2202 587 2203
rect 583 2197 587 2198
rect 454 2196 460 2197
rect 454 2192 455 2196
rect 459 2192 460 2196
rect 454 2191 460 2192
rect 582 2196 588 2197
rect 582 2192 583 2196
rect 587 2192 588 2196
rect 582 2191 588 2192
rect 608 2168 610 2234
rect 678 2216 684 2217
rect 678 2212 679 2216
rect 683 2212 684 2216
rect 678 2211 684 2212
rect 806 2216 812 2217
rect 806 2212 807 2216
rect 811 2212 812 2216
rect 806 2211 812 2212
rect 926 2216 932 2217
rect 926 2212 927 2216
rect 931 2212 932 2216
rect 926 2211 932 2212
rect 680 2203 682 2211
rect 808 2203 810 2211
rect 928 2203 930 2211
rect 679 2202 683 2203
rect 679 2197 683 2198
rect 703 2202 707 2203
rect 703 2197 707 2198
rect 807 2202 811 2203
rect 807 2197 811 2198
rect 823 2202 827 2203
rect 823 2197 827 2198
rect 927 2202 931 2203
rect 927 2197 931 2198
rect 943 2202 947 2203
rect 943 2197 947 2198
rect 702 2196 708 2197
rect 702 2192 703 2196
rect 707 2192 708 2196
rect 702 2191 708 2192
rect 822 2196 828 2197
rect 822 2192 823 2196
rect 827 2192 828 2196
rect 822 2191 828 2192
rect 942 2196 948 2197
rect 942 2192 943 2196
rect 947 2192 948 2196
rect 942 2191 948 2192
rect 952 2168 954 2234
rect 1046 2216 1052 2217
rect 1046 2212 1047 2216
rect 1051 2212 1052 2216
rect 1046 2211 1052 2212
rect 1158 2216 1164 2217
rect 1158 2212 1159 2216
rect 1163 2212 1164 2216
rect 1158 2211 1164 2212
rect 1168 2211 1170 2242
rect 1270 2241 1271 2245
rect 1275 2241 1276 2245
rect 1280 2244 1282 2266
rect 1366 2263 1367 2267
rect 1371 2263 1372 2267
rect 1366 2262 1372 2263
rect 1374 2267 1380 2268
rect 1374 2263 1375 2267
rect 1379 2263 1380 2267
rect 1374 2262 1380 2263
rect 1368 2251 1370 2262
rect 1367 2250 1371 2251
rect 1391 2250 1395 2251
rect 1367 2245 1371 2246
rect 1390 2245 1396 2246
rect 1270 2240 1276 2241
rect 1278 2243 1284 2244
rect 1278 2239 1279 2243
rect 1283 2239 1284 2243
rect 1390 2241 1391 2245
rect 1395 2241 1396 2245
rect 1400 2244 1402 2270
rect 1486 2267 1492 2268
rect 1486 2263 1487 2267
rect 1491 2263 1492 2267
rect 1630 2267 1631 2271
rect 1635 2267 1636 2271
rect 1630 2266 1636 2267
rect 1670 2271 1676 2272
rect 1670 2267 1671 2271
rect 1675 2267 1676 2271
rect 2022 2271 2023 2275
rect 2027 2271 2028 2275
rect 2022 2270 2028 2271
rect 1670 2266 1676 2267
rect 1486 2262 1492 2263
rect 1488 2251 1490 2262
rect 1632 2251 1634 2266
rect 1672 2263 1674 2266
rect 1671 2262 1675 2263
rect 2015 2262 2019 2263
rect 1671 2257 1675 2258
rect 2014 2257 2020 2258
rect 1672 2254 1674 2257
rect 1670 2253 1676 2254
rect 1487 2250 1491 2251
rect 1487 2245 1491 2246
rect 1631 2250 1635 2251
rect 1670 2249 1671 2253
rect 1675 2249 1676 2253
rect 2014 2253 2015 2257
rect 2019 2253 2020 2257
rect 2014 2252 2020 2253
rect 2024 2252 2026 2270
rect 2094 2267 2100 2268
rect 2094 2263 2095 2267
rect 2099 2263 2100 2267
rect 2094 2262 2100 2263
rect 2167 2262 2171 2263
rect 2095 2257 2099 2258
rect 2166 2257 2172 2258
rect 2166 2253 2167 2257
rect 2171 2253 2172 2257
rect 2166 2252 2172 2253
rect 2176 2252 2178 2330
rect 2182 2312 2188 2313
rect 2182 2308 2183 2312
rect 2187 2308 2188 2312
rect 2182 2307 2188 2308
rect 2334 2312 2340 2313
rect 2334 2308 2335 2312
rect 2339 2308 2340 2312
rect 2334 2307 2340 2308
rect 2478 2312 2484 2313
rect 2478 2308 2479 2312
rect 2483 2308 2484 2312
rect 2478 2307 2484 2308
rect 2184 2303 2186 2307
rect 2336 2303 2338 2307
rect 2480 2303 2482 2307
rect 2183 2302 2187 2303
rect 2183 2297 2187 2298
rect 2263 2302 2267 2303
rect 2263 2297 2267 2298
rect 2335 2302 2339 2303
rect 2335 2297 2339 2298
rect 2431 2302 2435 2303
rect 2431 2297 2435 2298
rect 2479 2302 2483 2303
rect 2479 2297 2483 2298
rect 2262 2296 2268 2297
rect 2262 2292 2263 2296
rect 2267 2292 2268 2296
rect 2262 2291 2268 2292
rect 2430 2296 2436 2297
rect 2430 2292 2431 2296
rect 2435 2292 2436 2296
rect 2430 2291 2436 2292
rect 2488 2268 2490 2330
rect 2622 2312 2628 2313
rect 2622 2308 2623 2312
rect 2627 2308 2628 2312
rect 2622 2307 2628 2308
rect 2624 2303 2626 2307
rect 2607 2302 2611 2303
rect 2607 2297 2611 2298
rect 2623 2302 2627 2303
rect 2623 2297 2627 2298
rect 2606 2296 2612 2297
rect 2606 2292 2607 2296
rect 2611 2292 2612 2296
rect 2606 2291 2612 2292
rect 2632 2268 2634 2334
rect 2766 2312 2772 2313
rect 2766 2308 2767 2312
rect 2771 2308 2772 2312
rect 2766 2307 2772 2308
rect 2768 2303 2770 2307
rect 2767 2302 2771 2303
rect 2767 2297 2771 2298
rect 2791 2302 2795 2303
rect 2791 2297 2795 2298
rect 2790 2296 2796 2297
rect 2790 2292 2791 2296
rect 2795 2292 2796 2296
rect 2790 2291 2796 2292
rect 2800 2272 2802 2334
rect 2918 2312 2924 2313
rect 2918 2308 2919 2312
rect 2923 2308 2924 2312
rect 2918 2307 2924 2308
rect 2920 2303 2922 2307
rect 2919 2302 2923 2303
rect 2919 2297 2923 2298
rect 2983 2302 2987 2303
rect 2983 2297 2987 2298
rect 2982 2296 2988 2297
rect 2982 2292 2983 2296
rect 2987 2292 2988 2296
rect 2982 2291 2988 2292
rect 3016 2272 3018 2334
rect 3159 2302 3163 2303
rect 3159 2297 3163 2298
rect 3158 2296 3164 2297
rect 3158 2292 3159 2296
rect 3163 2292 3164 2296
rect 3158 2291 3164 2292
rect 2798 2271 2804 2272
rect 2262 2267 2268 2268
rect 2262 2263 2263 2267
rect 2267 2263 2268 2267
rect 2262 2262 2268 2263
rect 2302 2267 2308 2268
rect 2302 2263 2303 2267
rect 2307 2263 2308 2267
rect 2430 2267 2436 2268
rect 2430 2263 2431 2267
rect 2435 2263 2436 2267
rect 2486 2267 2492 2268
rect 2486 2263 2487 2267
rect 2491 2263 2492 2267
rect 2302 2262 2308 2263
rect 2319 2262 2323 2263
rect 2430 2262 2436 2263
rect 2463 2262 2467 2263
rect 2486 2262 2492 2263
rect 2606 2267 2612 2268
rect 2606 2263 2607 2267
rect 2611 2263 2612 2267
rect 2606 2262 2612 2263
rect 2630 2267 2636 2268
rect 2630 2263 2631 2267
rect 2635 2263 2636 2267
rect 2790 2267 2796 2268
rect 2790 2263 2791 2267
rect 2795 2263 2796 2267
rect 2798 2267 2799 2271
rect 2803 2267 2804 2271
rect 2990 2271 2996 2272
rect 2798 2266 2804 2267
rect 2982 2267 2988 2268
rect 2630 2262 2636 2263
rect 2759 2262 2763 2263
rect 2790 2262 2796 2263
rect 2263 2257 2267 2258
rect 2304 2252 2306 2262
rect 2318 2257 2324 2258
rect 2431 2257 2435 2258
rect 2462 2257 2468 2258
rect 2318 2253 2319 2257
rect 2323 2253 2324 2257
rect 2318 2252 2324 2253
rect 2462 2253 2463 2257
rect 2467 2253 2468 2257
rect 2488 2256 2490 2262
rect 2606 2257 2612 2258
rect 2462 2252 2468 2253
rect 2486 2255 2492 2256
rect 1670 2248 1676 2249
rect 2022 2251 2028 2252
rect 2022 2247 2023 2251
rect 2027 2247 2028 2251
rect 2022 2246 2028 2247
rect 2174 2251 2180 2252
rect 2174 2247 2175 2251
rect 2179 2247 2180 2251
rect 2174 2246 2180 2247
rect 2302 2251 2308 2252
rect 2302 2247 2303 2251
rect 2307 2247 2308 2251
rect 2486 2251 2487 2255
rect 2491 2251 2492 2255
rect 2606 2253 2607 2257
rect 2611 2253 2612 2257
rect 2758 2257 2764 2258
rect 2791 2257 2795 2258
rect 2606 2252 2612 2253
rect 2614 2255 2620 2256
rect 2486 2250 2492 2251
rect 2614 2251 2615 2255
rect 2619 2251 2620 2255
rect 2758 2253 2759 2257
rect 2763 2253 2764 2257
rect 2800 2256 2802 2266
rect 2982 2263 2983 2267
rect 2987 2263 2988 2267
rect 2990 2267 2991 2271
rect 2995 2267 2996 2271
rect 2990 2266 2996 2267
rect 3014 2271 3020 2272
rect 3014 2267 3015 2271
rect 3019 2267 3020 2271
rect 3168 2268 3170 2346
rect 3191 2341 3195 2342
rect 3192 2338 3194 2341
rect 3190 2337 3196 2338
rect 3190 2333 3191 2337
rect 3195 2333 3196 2337
rect 3190 2332 3196 2333
rect 3190 2319 3196 2320
rect 3190 2315 3191 2319
rect 3195 2315 3196 2319
rect 3190 2314 3196 2315
rect 3192 2303 3194 2314
rect 3191 2302 3195 2303
rect 3191 2297 3195 2298
rect 3192 2290 3194 2297
rect 3190 2289 3196 2290
rect 3190 2285 3191 2289
rect 3195 2285 3196 2289
rect 3190 2284 3196 2285
rect 3190 2271 3196 2272
rect 3014 2266 3020 2267
rect 3158 2267 3164 2268
rect 2982 2262 2988 2263
rect 2983 2257 2987 2258
rect 2758 2252 2764 2253
rect 2766 2255 2772 2256
rect 2614 2250 2620 2251
rect 2766 2251 2767 2255
rect 2771 2251 2772 2255
rect 2766 2250 2772 2251
rect 2798 2255 2804 2256
rect 2798 2251 2799 2255
rect 2803 2251 2804 2255
rect 2798 2250 2804 2251
rect 2302 2246 2308 2247
rect 1631 2245 1635 2246
rect 1390 2240 1396 2241
rect 1398 2243 1404 2244
rect 1278 2238 1284 2239
rect 1398 2239 1399 2243
rect 1403 2239 1404 2243
rect 1632 2242 1634 2245
rect 1398 2238 1404 2239
rect 1630 2241 1636 2242
rect 1270 2216 1276 2217
rect 1270 2212 1271 2216
rect 1275 2212 1276 2216
rect 1270 2211 1276 2212
rect 1048 2203 1050 2211
rect 1160 2203 1162 2211
rect 1168 2209 1178 2211
rect 1047 2202 1051 2203
rect 1047 2197 1051 2198
rect 1055 2202 1059 2203
rect 1055 2197 1059 2198
rect 1159 2202 1163 2203
rect 1159 2197 1163 2198
rect 1167 2202 1171 2203
rect 1167 2197 1171 2198
rect 1054 2196 1060 2197
rect 1054 2192 1055 2196
rect 1059 2192 1060 2196
rect 1054 2191 1060 2192
rect 1166 2196 1172 2197
rect 1166 2192 1167 2196
rect 1171 2192 1172 2196
rect 1166 2191 1172 2192
rect 1176 2172 1178 2209
rect 1272 2203 1274 2211
rect 1271 2202 1275 2203
rect 1271 2197 1275 2198
rect 1280 2176 1282 2238
rect 1630 2237 1631 2241
rect 1635 2237 1636 2241
rect 1630 2236 1636 2237
rect 1670 2235 1676 2236
rect 1670 2231 1671 2235
rect 1675 2231 1676 2235
rect 1670 2230 1676 2231
rect 1630 2223 1636 2224
rect 1630 2219 1631 2223
rect 1635 2219 1636 2223
rect 1672 2219 1674 2230
rect 2014 2228 2020 2229
rect 2014 2224 2015 2228
rect 2019 2224 2020 2228
rect 2014 2223 2020 2224
rect 2016 2219 2018 2223
rect 1630 2218 1636 2219
rect 1671 2218 1675 2219
rect 1390 2216 1396 2217
rect 1390 2212 1391 2216
rect 1395 2212 1396 2216
rect 1390 2211 1396 2212
rect 1392 2203 1394 2211
rect 1632 2203 1634 2218
rect 1671 2213 1675 2214
rect 1927 2218 1931 2219
rect 1927 2213 1931 2214
rect 2015 2218 2019 2219
rect 2015 2213 2019 2214
rect 1672 2206 1674 2213
rect 1926 2212 1932 2213
rect 1926 2208 1927 2212
rect 1931 2208 1932 2212
rect 1926 2207 1932 2208
rect 1670 2205 1676 2206
rect 1287 2202 1291 2203
rect 1287 2197 1291 2198
rect 1391 2202 1395 2203
rect 1391 2197 1395 2198
rect 1631 2202 1635 2203
rect 1670 2201 1671 2205
rect 1675 2201 1676 2205
rect 1670 2200 1676 2201
rect 1631 2197 1635 2198
rect 1286 2196 1292 2197
rect 1286 2192 1287 2196
rect 1291 2192 1292 2196
rect 1286 2191 1292 2192
rect 1632 2190 1634 2197
rect 2024 2196 2026 2246
rect 2166 2228 2172 2229
rect 2166 2224 2167 2228
rect 2171 2224 2172 2228
rect 2166 2223 2172 2224
rect 2168 2219 2170 2223
rect 2103 2218 2107 2219
rect 2103 2213 2107 2214
rect 2167 2218 2171 2219
rect 2167 2213 2171 2214
rect 2102 2212 2108 2213
rect 2102 2208 2103 2212
rect 2107 2208 2108 2212
rect 2102 2207 2108 2208
rect 2022 2195 2028 2196
rect 2022 2191 2023 2195
rect 2027 2191 2028 2195
rect 2176 2192 2178 2246
rect 2295 2218 2299 2219
rect 2295 2213 2299 2214
rect 2294 2212 2300 2213
rect 2294 2208 2295 2212
rect 2299 2208 2300 2212
rect 2294 2207 2300 2208
rect 2022 2190 2028 2191
rect 2118 2191 2124 2192
rect 1630 2189 1636 2190
rect 1630 2185 1631 2189
rect 1635 2185 1636 2189
rect 1630 2184 1636 2185
rect 1670 2187 1676 2188
rect 1670 2183 1671 2187
rect 1675 2183 1676 2187
rect 2024 2184 2026 2190
rect 2118 2187 2119 2191
rect 2123 2187 2124 2191
rect 2118 2186 2124 2187
rect 2174 2191 2180 2192
rect 2174 2187 2175 2191
rect 2179 2187 2180 2191
rect 2174 2186 2180 2187
rect 1670 2182 1676 2183
rect 1926 2183 1932 2184
rect 1672 2179 1674 2182
rect 1926 2179 1927 2183
rect 1931 2179 1932 2183
rect 2022 2183 2028 2184
rect 2022 2179 2023 2183
rect 2027 2179 2028 2183
rect 1671 2178 1675 2179
rect 1278 2175 1284 2176
rect 1062 2171 1068 2172
rect 454 2167 460 2168
rect 454 2163 455 2167
rect 459 2163 460 2167
rect 454 2162 460 2163
rect 462 2167 468 2168
rect 462 2163 463 2167
rect 467 2163 468 2167
rect 462 2162 468 2163
rect 582 2167 588 2168
rect 582 2163 583 2167
rect 587 2163 588 2167
rect 582 2162 588 2163
rect 606 2167 612 2168
rect 606 2163 607 2167
rect 611 2163 612 2167
rect 606 2162 612 2163
rect 702 2167 708 2168
rect 702 2163 703 2167
rect 707 2163 708 2167
rect 702 2162 708 2163
rect 710 2167 716 2168
rect 710 2163 711 2167
rect 715 2163 716 2167
rect 710 2162 716 2163
rect 822 2167 828 2168
rect 822 2163 823 2167
rect 827 2163 828 2167
rect 822 2162 828 2163
rect 862 2167 868 2168
rect 862 2163 863 2167
rect 867 2163 868 2167
rect 862 2162 868 2163
rect 942 2167 948 2168
rect 942 2163 943 2167
rect 947 2163 948 2167
rect 942 2162 948 2163
rect 950 2167 956 2168
rect 950 2163 951 2167
rect 955 2163 956 2167
rect 950 2162 956 2163
rect 974 2167 980 2168
rect 974 2163 975 2167
rect 979 2163 980 2167
rect 974 2162 980 2163
rect 1054 2167 1060 2168
rect 1054 2163 1055 2167
rect 1059 2163 1060 2167
rect 1062 2167 1063 2171
rect 1067 2167 1068 2171
rect 1174 2171 1180 2172
rect 1062 2166 1068 2167
rect 1166 2167 1172 2168
rect 1054 2162 1060 2163
rect 1064 2163 1066 2166
rect 1166 2163 1167 2167
rect 1171 2163 1172 2167
rect 1174 2167 1175 2171
rect 1179 2167 1180 2171
rect 1278 2171 1279 2175
rect 1283 2171 1284 2175
rect 1847 2178 1851 2179
rect 1926 2178 1932 2179
rect 1999 2178 2003 2179
rect 2022 2178 2028 2179
rect 2102 2183 2108 2184
rect 2102 2179 2103 2183
rect 2107 2179 2108 2183
rect 2102 2178 2108 2179
rect 1671 2173 1675 2174
rect 1846 2173 1852 2174
rect 1927 2173 1931 2174
rect 1998 2173 2004 2174
rect 1278 2170 1284 2171
rect 1630 2171 1636 2172
rect 1174 2166 1180 2167
rect 1286 2167 1292 2168
rect 456 2151 458 2162
rect 351 2150 355 2151
rect 455 2150 459 2151
rect 350 2145 356 2146
rect 455 2145 459 2146
rect 350 2141 351 2145
rect 355 2141 356 2145
rect 350 2140 356 2141
rect 464 2140 466 2162
rect 584 2151 586 2162
rect 479 2150 483 2151
rect 583 2150 587 2151
rect 599 2150 603 2151
rect 478 2145 484 2146
rect 583 2145 587 2146
rect 598 2145 604 2146
rect 478 2141 479 2145
rect 483 2141 484 2145
rect 478 2140 484 2141
rect 598 2141 599 2145
rect 603 2141 604 2145
rect 598 2140 604 2141
rect 608 2140 610 2162
rect 704 2151 706 2162
rect 703 2150 707 2151
rect 703 2145 707 2146
rect 712 2140 714 2162
rect 824 2151 826 2162
rect 719 2150 723 2151
rect 823 2150 827 2151
rect 839 2150 843 2151
rect 718 2145 724 2146
rect 823 2145 827 2146
rect 838 2145 844 2146
rect 718 2141 719 2145
rect 723 2141 724 2145
rect 718 2140 724 2141
rect 838 2141 839 2145
rect 843 2141 844 2145
rect 838 2140 844 2141
rect 864 2140 866 2162
rect 944 2151 946 2162
rect 943 2150 947 2151
rect 951 2150 955 2151
rect 943 2145 947 2146
rect 950 2145 956 2146
rect 950 2141 951 2145
rect 955 2141 956 2145
rect 950 2140 956 2141
rect 976 2140 978 2162
rect 1056 2151 1058 2162
rect 1064 2161 1074 2163
rect 1166 2162 1172 2163
rect 1055 2150 1059 2151
rect 1063 2150 1067 2151
rect 1055 2145 1059 2146
rect 1062 2145 1068 2146
rect 1062 2141 1063 2145
rect 1067 2141 1068 2145
rect 1062 2140 1068 2141
rect 1072 2140 1074 2161
rect 1168 2151 1170 2162
rect 1167 2150 1171 2151
rect 1167 2145 1171 2146
rect 1176 2140 1178 2166
rect 1286 2163 1287 2167
rect 1291 2163 1292 2167
rect 1630 2167 1631 2171
rect 1635 2167 1636 2171
rect 1672 2170 1674 2173
rect 1630 2166 1636 2167
rect 1670 2169 1676 2170
rect 1286 2162 1292 2163
rect 1288 2151 1290 2162
rect 1632 2151 1634 2166
rect 1670 2165 1671 2169
rect 1675 2165 1676 2169
rect 1846 2169 1847 2173
rect 1851 2169 1852 2173
rect 1846 2168 1852 2169
rect 1998 2169 1999 2173
rect 2003 2169 2004 2173
rect 2024 2172 2026 2178
rect 2103 2173 2107 2174
rect 1998 2168 2004 2169
rect 2022 2171 2028 2172
rect 2022 2167 2023 2171
rect 2027 2167 2028 2171
rect 2022 2166 2028 2167
rect 1670 2164 1676 2165
rect 1670 2151 1676 2152
rect 1183 2150 1187 2151
rect 1287 2150 1291 2151
rect 1182 2145 1188 2146
rect 1287 2145 1291 2146
rect 1631 2150 1635 2151
rect 1670 2147 1671 2151
rect 1675 2147 1676 2151
rect 1670 2146 1676 2147
rect 1631 2145 1635 2146
rect 1182 2141 1183 2145
rect 1187 2141 1188 2145
rect 1632 2142 1634 2145
rect 1182 2140 1188 2141
rect 1630 2141 1636 2142
rect 382 2139 388 2140
rect 382 2135 383 2139
rect 387 2135 388 2139
rect 382 2134 388 2135
rect 462 2139 468 2140
rect 462 2135 463 2139
rect 467 2135 468 2139
rect 462 2134 468 2135
rect 606 2139 612 2140
rect 606 2135 607 2139
rect 611 2135 612 2139
rect 606 2134 612 2135
rect 710 2139 716 2140
rect 710 2135 711 2139
rect 715 2135 716 2139
rect 710 2134 716 2135
rect 862 2139 868 2140
rect 862 2135 863 2139
rect 867 2135 868 2139
rect 862 2134 868 2135
rect 974 2139 980 2140
rect 974 2135 975 2139
rect 979 2135 980 2139
rect 974 2134 980 2135
rect 1070 2139 1076 2140
rect 1070 2135 1071 2139
rect 1075 2135 1076 2139
rect 1070 2134 1076 2135
rect 1174 2139 1180 2140
rect 1174 2135 1175 2139
rect 1179 2135 1180 2139
rect 1630 2137 1631 2141
rect 1635 2137 1636 2141
rect 1630 2136 1636 2137
rect 1672 2135 1674 2146
rect 1846 2144 1852 2145
rect 1846 2140 1847 2144
rect 1851 2140 1852 2144
rect 1846 2139 1852 2140
rect 1998 2144 2004 2145
rect 1998 2140 1999 2144
rect 2003 2140 2004 2144
rect 1998 2139 2004 2140
rect 1848 2135 1850 2139
rect 2000 2135 2002 2139
rect 1174 2134 1180 2135
rect 1671 2134 1675 2135
rect 350 2116 356 2117
rect 350 2112 351 2116
rect 355 2112 356 2116
rect 350 2111 356 2112
rect 352 2099 354 2111
rect 247 2098 251 2099
rect 247 2093 251 2094
rect 351 2098 355 2099
rect 351 2093 355 2094
rect 375 2098 379 2099
rect 375 2093 379 2094
rect 246 2092 252 2093
rect 246 2088 247 2092
rect 251 2088 252 2092
rect 246 2087 252 2088
rect 374 2092 380 2093
rect 374 2088 375 2092
rect 379 2088 380 2092
rect 374 2087 380 2088
rect 384 2064 386 2134
rect 478 2116 484 2117
rect 478 2112 479 2116
rect 483 2112 484 2116
rect 478 2111 484 2112
rect 598 2116 604 2117
rect 598 2112 599 2116
rect 603 2112 604 2116
rect 598 2111 604 2112
rect 480 2099 482 2111
rect 600 2099 602 2111
rect 479 2098 483 2099
rect 479 2093 483 2094
rect 503 2098 507 2099
rect 503 2093 507 2094
rect 599 2098 603 2099
rect 599 2093 603 2094
rect 502 2092 508 2093
rect 502 2088 503 2092
rect 507 2088 508 2092
rect 502 2087 508 2088
rect 608 2072 610 2134
rect 718 2116 724 2117
rect 718 2112 719 2116
rect 723 2112 724 2116
rect 718 2111 724 2112
rect 838 2116 844 2117
rect 838 2112 839 2116
rect 843 2112 844 2116
rect 838 2111 844 2112
rect 720 2099 722 2111
rect 840 2099 842 2111
rect 623 2098 627 2099
rect 623 2093 627 2094
rect 719 2098 723 2099
rect 719 2093 723 2094
rect 743 2098 747 2099
rect 743 2093 747 2094
rect 839 2098 843 2099
rect 839 2093 843 2094
rect 855 2098 859 2099
rect 855 2093 859 2094
rect 622 2092 628 2093
rect 622 2088 623 2092
rect 627 2088 628 2092
rect 622 2087 628 2088
rect 742 2092 748 2093
rect 742 2088 743 2092
rect 747 2088 748 2092
rect 742 2087 748 2088
rect 854 2092 860 2093
rect 854 2088 855 2092
rect 859 2088 860 2092
rect 854 2087 860 2088
rect 606 2071 612 2072
rect 606 2067 607 2071
rect 611 2067 612 2071
rect 606 2066 612 2067
rect 864 2064 866 2134
rect 950 2116 956 2117
rect 950 2112 951 2116
rect 955 2112 956 2116
rect 950 2111 956 2112
rect 952 2099 954 2111
rect 951 2098 955 2099
rect 951 2093 955 2094
rect 967 2098 971 2099
rect 967 2093 971 2094
rect 966 2092 972 2093
rect 966 2088 967 2092
rect 971 2088 972 2092
rect 966 2087 972 2088
rect 976 2064 978 2134
rect 1062 2116 1068 2117
rect 1062 2112 1063 2116
rect 1067 2112 1068 2116
rect 1062 2111 1068 2112
rect 1064 2099 1066 2111
rect 1063 2098 1067 2099
rect 1063 2093 1067 2094
rect 1072 2072 1074 2134
rect 1671 2129 1675 2130
rect 1759 2134 1763 2135
rect 1759 2129 1763 2130
rect 1847 2134 1851 2135
rect 1847 2129 1851 2130
rect 1911 2134 1915 2135
rect 1911 2129 1915 2130
rect 1999 2134 2003 2135
rect 1999 2129 2003 2130
rect 1630 2123 1636 2124
rect 1630 2119 1631 2123
rect 1635 2119 1636 2123
rect 1672 2122 1674 2129
rect 1758 2128 1764 2129
rect 1758 2124 1759 2128
rect 1763 2124 1764 2128
rect 1758 2123 1764 2124
rect 1910 2128 1916 2129
rect 1910 2124 1911 2128
rect 1915 2124 1916 2128
rect 1910 2123 1916 2124
rect 1630 2118 1636 2119
rect 1670 2121 1676 2122
rect 1182 2116 1188 2117
rect 1182 2112 1183 2116
rect 1187 2112 1188 2116
rect 1182 2111 1188 2112
rect 1184 2099 1186 2111
rect 1632 2099 1634 2118
rect 1670 2117 1671 2121
rect 1675 2117 1676 2121
rect 1670 2116 1676 2117
rect 1670 2103 1676 2104
rect 1670 2099 1671 2103
rect 1675 2099 1676 2103
rect 1087 2098 1091 2099
rect 1087 2093 1091 2094
rect 1183 2098 1187 2099
rect 1183 2093 1187 2094
rect 1631 2098 1635 2099
rect 1670 2098 1676 2099
rect 1758 2099 1764 2100
rect 1672 2095 1674 2098
rect 1758 2095 1759 2099
rect 1763 2095 1764 2099
rect 1910 2099 1916 2100
rect 1910 2095 1911 2099
rect 1915 2095 1916 2099
rect 1631 2093 1635 2094
rect 1671 2094 1675 2095
rect 1086 2092 1092 2093
rect 1086 2088 1087 2092
rect 1091 2088 1092 2092
rect 1086 2087 1092 2088
rect 1632 2086 1634 2093
rect 1695 2094 1699 2095
rect 1758 2094 1764 2095
rect 1823 2094 1827 2095
rect 1910 2094 1916 2095
rect 1967 2094 1971 2095
rect 1671 2089 1675 2090
rect 1694 2089 1700 2090
rect 1759 2089 1763 2090
rect 1822 2089 1828 2090
rect 1911 2089 1915 2090
rect 1966 2089 1972 2090
rect 1672 2086 1674 2089
rect 1630 2085 1636 2086
rect 1630 2081 1631 2085
rect 1635 2081 1636 2085
rect 1630 2080 1636 2081
rect 1670 2085 1676 2086
rect 1670 2081 1671 2085
rect 1675 2081 1676 2085
rect 1694 2085 1695 2089
rect 1699 2085 1700 2089
rect 1694 2084 1700 2085
rect 1822 2085 1823 2089
rect 1827 2085 1828 2089
rect 1822 2084 1828 2085
rect 1966 2085 1967 2089
rect 1971 2085 1972 2089
rect 2024 2088 2026 2166
rect 2071 2134 2075 2135
rect 2071 2129 2075 2130
rect 2070 2128 2076 2129
rect 2070 2124 2071 2128
rect 2075 2124 2076 2128
rect 2070 2123 2076 2124
rect 2120 2104 2122 2186
rect 2151 2178 2155 2179
rect 2150 2173 2156 2174
rect 2150 2169 2151 2173
rect 2155 2169 2156 2173
rect 2176 2172 2178 2186
rect 2304 2184 2306 2246
rect 2318 2228 2324 2229
rect 2318 2224 2319 2228
rect 2323 2224 2324 2228
rect 2318 2223 2324 2224
rect 2462 2228 2468 2229
rect 2462 2224 2463 2228
rect 2467 2224 2468 2228
rect 2462 2223 2468 2224
rect 2606 2228 2612 2229
rect 2606 2224 2607 2228
rect 2611 2224 2612 2228
rect 2606 2223 2612 2224
rect 2320 2219 2322 2223
rect 2464 2219 2466 2223
rect 2608 2219 2610 2223
rect 2319 2218 2323 2219
rect 2319 2213 2323 2214
rect 2463 2218 2467 2219
rect 2463 2213 2467 2214
rect 2503 2218 2507 2219
rect 2503 2213 2507 2214
rect 2607 2218 2611 2219
rect 2607 2213 2611 2214
rect 2502 2212 2508 2213
rect 2502 2208 2503 2212
rect 2507 2208 2508 2212
rect 2502 2207 2508 2208
rect 2616 2184 2618 2250
rect 2758 2228 2764 2229
rect 2758 2224 2759 2228
rect 2763 2224 2764 2228
rect 2758 2223 2764 2224
rect 2760 2219 2762 2223
rect 2719 2218 2723 2219
rect 2719 2213 2723 2214
rect 2759 2218 2763 2219
rect 2759 2213 2763 2214
rect 2718 2212 2724 2213
rect 2718 2208 2719 2212
rect 2723 2208 2724 2212
rect 2718 2207 2724 2208
rect 2768 2188 2770 2250
rect 2951 2218 2955 2219
rect 2951 2213 2955 2214
rect 2950 2212 2956 2213
rect 2950 2208 2951 2212
rect 2955 2208 2956 2212
rect 2950 2207 2956 2208
rect 2992 2188 2994 2266
rect 3158 2263 3159 2267
rect 3163 2263 3164 2267
rect 3158 2262 3164 2263
rect 3166 2267 3172 2268
rect 3166 2263 3167 2267
rect 3171 2263 3172 2267
rect 3190 2267 3191 2271
rect 3195 2267 3196 2271
rect 3190 2266 3196 2267
rect 3192 2263 3194 2266
rect 3166 2262 3172 2263
rect 3191 2262 3195 2263
rect 3159 2257 3163 2258
rect 3159 2218 3163 2219
rect 3159 2213 3163 2214
rect 3158 2212 3164 2213
rect 3158 2208 3159 2212
rect 3163 2208 3164 2212
rect 3158 2207 3164 2208
rect 2726 2187 2732 2188
rect 2294 2183 2300 2184
rect 2294 2179 2295 2183
rect 2299 2179 2300 2183
rect 2294 2178 2300 2179
rect 2302 2183 2308 2184
rect 2302 2179 2303 2183
rect 2307 2179 2308 2183
rect 2502 2183 2508 2184
rect 2502 2179 2503 2183
rect 2507 2179 2508 2183
rect 2614 2183 2620 2184
rect 2614 2179 2615 2183
rect 2619 2179 2620 2183
rect 2302 2178 2308 2179
rect 2447 2178 2451 2179
rect 2502 2178 2508 2179
rect 2599 2178 2603 2179
rect 2614 2178 2620 2179
rect 2718 2183 2724 2184
rect 2718 2179 2719 2183
rect 2723 2179 2724 2183
rect 2726 2183 2727 2187
rect 2731 2183 2732 2187
rect 2726 2182 2732 2183
rect 2766 2187 2772 2188
rect 2766 2183 2767 2187
rect 2771 2183 2772 2187
rect 2958 2187 2964 2188
rect 2766 2182 2772 2183
rect 2950 2183 2956 2184
rect 2718 2178 2724 2179
rect 2294 2173 2300 2174
rect 2150 2168 2156 2169
rect 2174 2171 2180 2172
rect 2174 2167 2175 2171
rect 2179 2167 2180 2171
rect 2294 2169 2295 2173
rect 2299 2169 2300 2173
rect 2294 2168 2300 2169
rect 2304 2168 2306 2178
rect 2446 2173 2452 2174
rect 2503 2173 2507 2174
rect 2598 2173 2604 2174
rect 2719 2173 2723 2174
rect 2446 2169 2447 2173
rect 2451 2169 2452 2173
rect 2446 2168 2452 2169
rect 2470 2171 2476 2172
rect 2174 2166 2180 2167
rect 2302 2167 2308 2168
rect 2302 2163 2303 2167
rect 2307 2163 2308 2167
rect 2470 2167 2471 2171
rect 2475 2167 2476 2171
rect 2598 2169 2599 2173
rect 2603 2169 2604 2173
rect 2598 2168 2604 2169
rect 2470 2166 2476 2167
rect 2302 2162 2308 2163
rect 2150 2144 2156 2145
rect 2150 2140 2151 2144
rect 2155 2140 2156 2144
rect 2150 2139 2156 2140
rect 2294 2144 2300 2145
rect 2294 2140 2295 2144
rect 2299 2140 2300 2144
rect 2294 2139 2300 2140
rect 2152 2135 2154 2139
rect 2296 2135 2298 2139
rect 2151 2134 2155 2135
rect 2151 2129 2155 2130
rect 2255 2134 2259 2135
rect 2255 2129 2259 2130
rect 2295 2134 2299 2135
rect 2295 2129 2299 2130
rect 2254 2128 2260 2129
rect 2254 2124 2255 2128
rect 2259 2124 2260 2128
rect 2254 2123 2260 2124
rect 2118 2103 2124 2104
rect 2070 2099 2076 2100
rect 2070 2095 2071 2099
rect 2075 2095 2076 2099
rect 2118 2099 2119 2103
rect 2123 2099 2124 2103
rect 2304 2100 2306 2162
rect 2446 2144 2452 2145
rect 2446 2140 2447 2144
rect 2451 2140 2452 2144
rect 2446 2139 2452 2140
rect 2448 2135 2450 2139
rect 2447 2134 2451 2135
rect 2447 2129 2451 2130
rect 2463 2134 2467 2135
rect 2463 2129 2467 2130
rect 2462 2128 2468 2129
rect 2462 2124 2463 2128
rect 2467 2124 2468 2128
rect 2462 2123 2468 2124
rect 2472 2104 2474 2166
rect 2598 2144 2604 2145
rect 2598 2140 2599 2144
rect 2603 2140 2604 2144
rect 2598 2139 2604 2140
rect 2600 2135 2602 2139
rect 2599 2134 2603 2135
rect 2599 2129 2603 2130
rect 2687 2134 2691 2135
rect 2687 2129 2691 2130
rect 2686 2128 2692 2129
rect 2686 2124 2687 2128
rect 2691 2124 2692 2128
rect 2686 2123 2692 2124
rect 2728 2104 2730 2182
rect 2950 2179 2951 2183
rect 2955 2179 2956 2183
rect 2958 2183 2959 2187
rect 2963 2183 2964 2187
rect 2958 2182 2964 2183
rect 2990 2187 2996 2188
rect 2990 2183 2991 2187
rect 2995 2183 2996 2187
rect 3168 2184 3170 2262
rect 3191 2257 3195 2258
rect 3192 2254 3194 2257
rect 3190 2253 3196 2254
rect 3190 2249 3191 2253
rect 3195 2249 3196 2253
rect 3190 2248 3196 2249
rect 3190 2235 3196 2236
rect 3190 2231 3191 2235
rect 3195 2231 3196 2235
rect 3190 2230 3196 2231
rect 3192 2219 3194 2230
rect 3191 2218 3195 2219
rect 3191 2213 3195 2214
rect 3192 2206 3194 2213
rect 3190 2205 3196 2206
rect 3190 2201 3191 2205
rect 3195 2201 3196 2205
rect 3190 2200 3196 2201
rect 3190 2187 3196 2188
rect 2990 2182 2996 2183
rect 3158 2183 3164 2184
rect 2950 2178 2956 2179
rect 2951 2173 2955 2174
rect 2927 2134 2931 2135
rect 2927 2129 2931 2130
rect 2926 2128 2932 2129
rect 2926 2124 2927 2128
rect 2931 2124 2932 2128
rect 2926 2123 2932 2124
rect 2960 2104 2962 2182
rect 3158 2179 3159 2183
rect 3163 2179 3164 2183
rect 3158 2178 3164 2179
rect 3166 2183 3172 2184
rect 3166 2179 3167 2183
rect 3171 2179 3172 2183
rect 3190 2183 3191 2187
rect 3195 2183 3196 2187
rect 3190 2182 3196 2183
rect 3192 2179 3194 2182
rect 3166 2178 3172 2179
rect 3191 2178 3195 2179
rect 3159 2173 3163 2174
rect 3159 2134 3163 2135
rect 3159 2129 3163 2130
rect 3158 2128 3164 2129
rect 3158 2124 3159 2128
rect 3163 2124 3164 2128
rect 3158 2123 3164 2124
rect 2470 2103 2476 2104
rect 2118 2098 2124 2099
rect 2254 2099 2260 2100
rect 2070 2094 2076 2095
rect 2111 2094 2115 2095
rect 2071 2089 2075 2090
rect 2110 2089 2116 2090
rect 1966 2084 1972 2085
rect 2022 2087 2028 2088
rect 1670 2080 1676 2081
rect 1702 2083 1708 2084
rect 1702 2079 1703 2083
rect 1707 2079 1708 2083
rect 2022 2083 2023 2087
rect 2027 2083 2028 2087
rect 2110 2085 2111 2089
rect 2115 2085 2116 2089
rect 2120 2088 2122 2098
rect 2254 2095 2255 2099
rect 2259 2095 2260 2099
rect 2254 2094 2260 2095
rect 2302 2099 2308 2100
rect 2302 2095 2303 2099
rect 2307 2095 2308 2099
rect 2462 2099 2468 2100
rect 2462 2095 2463 2099
rect 2467 2095 2468 2099
rect 2470 2099 2471 2103
rect 2475 2099 2476 2103
rect 2726 2103 2732 2104
rect 2470 2098 2476 2099
rect 2686 2099 2692 2100
rect 2302 2094 2308 2095
rect 2407 2094 2411 2095
rect 2462 2094 2468 2095
rect 2254 2089 2260 2090
rect 2110 2084 2116 2085
rect 2118 2087 2124 2088
rect 2022 2082 2028 2083
rect 2118 2083 2119 2087
rect 2123 2083 2124 2087
rect 2254 2085 2255 2089
rect 2259 2085 2260 2089
rect 2254 2084 2260 2085
rect 2406 2089 2412 2090
rect 2463 2089 2467 2090
rect 2406 2085 2407 2089
rect 2411 2085 2412 2089
rect 2472 2088 2474 2098
rect 2686 2095 2687 2099
rect 2691 2095 2692 2099
rect 2726 2099 2727 2103
rect 2731 2099 2732 2103
rect 2958 2103 2964 2104
rect 2726 2098 2732 2099
rect 2926 2099 2932 2100
rect 2686 2094 2692 2095
rect 2687 2089 2691 2090
rect 2406 2084 2412 2085
rect 2414 2087 2420 2088
rect 2118 2082 2124 2083
rect 2246 2083 2252 2084
rect 1702 2078 1708 2079
rect 1070 2071 1076 2072
rect 1070 2067 1071 2071
rect 1075 2067 1076 2071
rect 1070 2066 1076 2067
rect 1190 2067 1196 2068
rect 246 2063 252 2064
rect 246 2059 247 2063
rect 251 2059 252 2063
rect 246 2058 252 2059
rect 254 2063 260 2064
rect 254 2059 255 2063
rect 259 2059 260 2063
rect 254 2058 260 2059
rect 374 2063 380 2064
rect 374 2059 375 2063
rect 379 2059 380 2063
rect 374 2058 380 2059
rect 382 2063 388 2064
rect 382 2059 383 2063
rect 387 2059 388 2063
rect 382 2058 388 2059
rect 502 2063 508 2064
rect 502 2059 503 2063
rect 507 2059 508 2063
rect 502 2058 508 2059
rect 566 2063 572 2064
rect 566 2059 567 2063
rect 571 2059 572 2063
rect 566 2058 572 2059
rect 622 2063 628 2064
rect 622 2059 623 2063
rect 627 2059 628 2063
rect 622 2058 628 2059
rect 742 2063 748 2064
rect 742 2059 743 2063
rect 747 2059 748 2063
rect 742 2058 748 2059
rect 766 2063 772 2064
rect 766 2059 767 2063
rect 771 2059 772 2063
rect 766 2058 772 2059
rect 854 2063 860 2064
rect 854 2059 855 2063
rect 859 2059 860 2063
rect 854 2058 860 2059
rect 862 2063 868 2064
rect 862 2059 863 2063
rect 867 2059 868 2063
rect 862 2058 868 2059
rect 966 2063 972 2064
rect 966 2059 967 2063
rect 971 2059 972 2063
rect 966 2058 972 2059
rect 974 2063 980 2064
rect 974 2059 975 2063
rect 979 2059 980 2063
rect 974 2058 980 2059
rect 1086 2063 1092 2064
rect 1086 2059 1087 2063
rect 1091 2059 1092 2063
rect 1190 2063 1191 2067
rect 1195 2063 1196 2067
rect 1190 2062 1196 2063
rect 1630 2067 1636 2068
rect 1630 2063 1631 2067
rect 1635 2063 1636 2067
rect 1630 2062 1636 2063
rect 1670 2067 1676 2068
rect 1670 2063 1671 2067
rect 1675 2063 1676 2067
rect 1670 2062 1676 2063
rect 1086 2058 1092 2059
rect 248 2051 250 2058
rect 247 2050 251 2051
rect 247 2045 251 2046
rect 110 2036 116 2037
rect 182 2039 188 2040
rect 182 2035 183 2039
rect 187 2035 188 2039
rect 182 2034 188 2035
rect 110 2023 116 2024
rect 110 2019 111 2023
rect 115 2019 116 2023
rect 110 2018 116 2019
rect 112 2011 114 2018
rect 174 2016 180 2017
rect 174 2012 175 2016
rect 179 2012 180 2016
rect 174 2011 180 2012
rect 111 2010 115 2011
rect 111 2005 115 2006
rect 135 2010 139 2011
rect 135 2005 139 2006
rect 175 2010 179 2011
rect 175 2005 179 2006
rect 112 1998 114 2005
rect 134 2004 140 2005
rect 134 2000 135 2004
rect 139 2000 140 2004
rect 134 1999 140 2000
rect 110 1997 116 1998
rect 110 1993 111 1997
rect 115 1993 116 1997
rect 110 1992 116 1993
rect 184 1984 186 2034
rect 231 2010 235 2011
rect 231 2005 235 2006
rect 230 2004 236 2005
rect 230 2000 231 2004
rect 235 2000 236 2004
rect 230 1999 236 2000
rect 256 1984 258 2058
rect 376 2051 378 2058
rect 367 2050 371 2051
rect 375 2050 379 2051
rect 366 2045 372 2046
rect 375 2045 379 2046
rect 366 2041 367 2045
rect 371 2041 372 2045
rect 366 2040 372 2041
rect 375 2039 381 2040
rect 375 2035 376 2039
rect 380 2038 381 2039
rect 384 2038 386 2058
rect 504 2051 506 2058
rect 503 2050 507 2051
rect 559 2050 563 2051
rect 503 2045 507 2046
rect 558 2045 564 2046
rect 558 2041 559 2045
rect 563 2041 564 2045
rect 558 2040 564 2041
rect 568 2040 570 2058
rect 624 2051 626 2058
rect 744 2051 746 2058
rect 623 2050 627 2051
rect 623 2045 627 2046
rect 743 2050 747 2051
rect 759 2050 763 2051
rect 743 2045 747 2046
rect 758 2045 764 2046
rect 758 2041 759 2045
rect 763 2041 764 2045
rect 758 2040 764 2041
rect 768 2040 770 2058
rect 856 2051 858 2058
rect 855 2050 859 2051
rect 855 2045 859 2046
rect 380 2036 386 2038
rect 566 2039 572 2040
rect 380 2035 381 2036
rect 375 2034 381 2035
rect 566 2035 567 2039
rect 571 2035 572 2039
rect 566 2034 572 2035
rect 766 2039 772 2040
rect 766 2035 767 2039
rect 771 2035 772 2039
rect 766 2034 772 2035
rect 366 2016 372 2017
rect 366 2012 367 2016
rect 371 2012 372 2016
rect 366 2011 372 2012
rect 351 2010 355 2011
rect 351 2005 355 2006
rect 367 2010 371 2011
rect 367 2005 371 2006
rect 350 2004 356 2005
rect 350 2000 351 2004
rect 355 2000 356 2004
rect 350 1999 356 2000
rect 376 1984 378 2034
rect 558 2016 564 2017
rect 558 2012 559 2016
rect 563 2012 564 2016
rect 558 2011 564 2012
rect 463 2010 467 2011
rect 463 2005 467 2006
rect 559 2010 563 2011
rect 559 2005 563 2006
rect 462 2004 468 2005
rect 462 2000 463 2004
rect 467 2000 468 2004
rect 462 1999 468 2000
rect 568 1984 570 2034
rect 758 2016 764 2017
rect 758 2012 759 2016
rect 763 2012 764 2016
rect 758 2011 764 2012
rect 575 2010 579 2011
rect 575 2005 579 2006
rect 687 2010 691 2011
rect 687 2005 691 2006
rect 759 2010 763 2011
rect 759 2005 763 2006
rect 574 2004 580 2005
rect 574 2000 575 2004
rect 579 2000 580 2004
rect 574 1999 580 2000
rect 686 2004 692 2005
rect 686 2000 687 2004
rect 691 2000 692 2004
rect 686 1999 692 2000
rect 182 1983 188 1984
rect 110 1979 116 1980
rect 110 1975 111 1979
rect 115 1975 116 1979
rect 182 1979 183 1983
rect 187 1979 188 1983
rect 182 1978 188 1979
rect 254 1983 260 1984
rect 254 1979 255 1983
rect 259 1979 260 1983
rect 254 1978 260 1979
rect 374 1983 380 1984
rect 374 1979 375 1983
rect 379 1979 380 1983
rect 374 1978 380 1979
rect 566 1983 572 1984
rect 566 1979 567 1983
rect 571 1979 572 1983
rect 566 1978 572 1979
rect 110 1974 116 1975
rect 134 1975 140 1976
rect 112 1963 114 1974
rect 134 1971 135 1975
rect 139 1971 140 1975
rect 134 1970 140 1971
rect 142 1975 148 1976
rect 142 1971 143 1975
rect 147 1971 148 1975
rect 142 1970 148 1971
rect 230 1975 236 1976
rect 230 1971 231 1975
rect 235 1971 236 1975
rect 230 1970 236 1971
rect 350 1975 356 1976
rect 350 1971 351 1975
rect 355 1971 356 1975
rect 350 1970 356 1971
rect 462 1975 468 1976
rect 462 1971 463 1975
rect 467 1971 468 1975
rect 462 1970 468 1971
rect 574 1975 580 1976
rect 574 1971 575 1975
rect 579 1971 580 1975
rect 574 1970 580 1971
rect 686 1975 692 1976
rect 686 1971 687 1975
rect 691 1971 692 1975
rect 686 1970 692 1971
rect 136 1963 138 1970
rect 111 1962 115 1963
rect 111 1957 115 1958
rect 135 1962 139 1963
rect 135 1957 139 1958
rect 112 1954 114 1957
rect 110 1953 116 1954
rect 110 1949 111 1953
rect 115 1949 116 1953
rect 110 1948 116 1949
rect 110 1935 116 1936
rect 110 1931 111 1935
rect 115 1931 116 1935
rect 110 1930 116 1931
rect 112 1911 114 1930
rect 111 1910 115 1911
rect 111 1905 115 1906
rect 112 1898 114 1905
rect 110 1897 116 1898
rect 110 1893 111 1897
rect 115 1893 116 1897
rect 110 1892 116 1893
rect 110 1879 116 1880
rect 110 1875 111 1879
rect 115 1875 116 1879
rect 110 1874 116 1875
rect 112 1859 114 1874
rect 111 1858 115 1859
rect 111 1853 115 1854
rect 112 1850 114 1853
rect 110 1849 116 1850
rect 110 1845 111 1849
rect 115 1845 116 1849
rect 110 1844 116 1845
rect 110 1831 116 1832
rect 110 1827 111 1831
rect 115 1827 116 1831
rect 110 1826 116 1827
rect 112 1811 114 1826
rect 111 1810 115 1811
rect 111 1805 115 1806
rect 112 1798 114 1805
rect 110 1797 116 1798
rect 110 1793 111 1797
rect 115 1793 116 1797
rect 110 1792 116 1793
rect 110 1779 116 1780
rect 110 1775 111 1779
rect 115 1775 116 1779
rect 110 1774 116 1775
rect 112 1759 114 1774
rect 111 1758 115 1759
rect 111 1753 115 1754
rect 112 1750 114 1753
rect 110 1749 116 1750
rect 110 1745 111 1749
rect 115 1745 116 1749
rect 110 1744 116 1745
rect 110 1731 116 1732
rect 110 1727 111 1731
rect 115 1727 116 1731
rect 110 1726 116 1727
rect 112 1707 114 1726
rect 111 1706 115 1707
rect 111 1701 115 1702
rect 112 1694 114 1701
rect 110 1693 116 1694
rect 110 1689 111 1693
rect 115 1689 116 1693
rect 110 1688 116 1689
rect 110 1675 116 1676
rect 110 1671 111 1675
rect 115 1671 116 1675
rect 110 1670 116 1671
rect 112 1655 114 1670
rect 111 1654 115 1655
rect 135 1654 139 1655
rect 111 1649 115 1650
rect 134 1649 140 1650
rect 112 1646 114 1649
rect 110 1645 116 1646
rect 110 1641 111 1645
rect 115 1641 116 1645
rect 134 1645 135 1649
rect 139 1645 140 1649
rect 134 1644 140 1645
rect 144 1644 146 1970
rect 232 1963 234 1970
rect 352 1963 354 1970
rect 464 1963 466 1970
rect 576 1963 578 1970
rect 688 1963 690 1970
rect 768 1968 770 2034
rect 799 2010 803 2011
rect 799 2005 803 2006
rect 798 2004 804 2005
rect 798 2000 799 2004
rect 803 2000 804 2004
rect 798 1999 804 2000
rect 798 1975 804 1976
rect 798 1971 799 1975
rect 803 1971 804 1975
rect 798 1970 804 1971
rect 766 1967 772 1968
rect 766 1963 767 1967
rect 771 1963 772 1967
rect 800 1963 802 1970
rect 864 1964 866 2058
rect 968 2051 970 2058
rect 967 2050 971 2051
rect 966 2045 972 2046
rect 966 2041 967 2045
rect 971 2041 972 2045
rect 966 2040 972 2041
rect 976 2040 978 2058
rect 1088 2051 1090 2058
rect 1087 2050 1091 2051
rect 1183 2050 1187 2051
rect 1087 2045 1091 2046
rect 1182 2045 1188 2046
rect 1182 2041 1183 2045
rect 1187 2041 1188 2045
rect 1192 2044 1194 2062
rect 1632 2051 1634 2062
rect 1672 2055 1674 2062
rect 1694 2060 1700 2061
rect 1694 2056 1695 2060
rect 1699 2056 1700 2060
rect 1694 2055 1700 2056
rect 1671 2054 1675 2055
rect 1399 2050 1403 2051
rect 1599 2050 1603 2051
rect 1631 2050 1635 2051
rect 1671 2049 1675 2050
rect 1695 2054 1699 2055
rect 1695 2049 1699 2050
rect 1398 2045 1404 2046
rect 1182 2040 1188 2041
rect 1190 2043 1196 2044
rect 918 2039 924 2040
rect 918 2035 919 2039
rect 923 2035 924 2039
rect 918 2034 924 2035
rect 974 2039 980 2040
rect 974 2035 975 2039
rect 979 2035 980 2039
rect 1190 2039 1191 2043
rect 1195 2039 1196 2043
rect 1398 2041 1399 2045
rect 1403 2041 1404 2045
rect 1398 2040 1404 2041
rect 1598 2045 1604 2046
rect 1631 2045 1635 2046
rect 1598 2041 1599 2045
rect 1603 2041 1604 2045
rect 1632 2042 1634 2045
rect 1672 2042 1674 2049
rect 1694 2048 1700 2049
rect 1694 2044 1695 2048
rect 1699 2044 1700 2048
rect 1694 2043 1700 2044
rect 1598 2040 1604 2041
rect 1630 2041 1636 2042
rect 1190 2038 1196 2039
rect 1410 2039 1416 2040
rect 974 2034 980 2035
rect 1410 2035 1411 2039
rect 1415 2035 1416 2039
rect 1630 2037 1631 2041
rect 1635 2037 1636 2041
rect 1630 2036 1636 2037
rect 1670 2041 1676 2042
rect 1670 2037 1671 2041
rect 1675 2037 1676 2041
rect 1670 2036 1676 2037
rect 1704 2036 1706 2078
rect 1822 2060 1828 2061
rect 1822 2056 1823 2060
rect 1827 2056 1828 2060
rect 1822 2055 1828 2056
rect 1966 2060 1972 2061
rect 1966 2056 1967 2060
rect 1971 2056 1972 2060
rect 1966 2055 1972 2056
rect 1823 2054 1827 2055
rect 1823 2049 1827 2050
rect 1967 2054 1971 2055
rect 1967 2049 1971 2050
rect 1410 2034 1416 2035
rect 1610 2035 1616 2036
rect 911 2010 915 2011
rect 911 2005 915 2006
rect 910 2004 916 2005
rect 910 2000 911 2004
rect 915 2000 916 2004
rect 910 1999 916 2000
rect 920 1976 922 2034
rect 966 2016 972 2017
rect 966 2012 967 2016
rect 971 2012 972 2016
rect 966 2011 972 2012
rect 1182 2016 1188 2017
rect 1182 2012 1183 2016
rect 1187 2012 1188 2016
rect 1182 2011 1188 2012
rect 1398 2016 1404 2017
rect 1398 2012 1399 2016
rect 1403 2012 1404 2016
rect 1398 2011 1404 2012
rect 967 2010 971 2011
rect 967 2005 971 2006
rect 1183 2010 1187 2011
rect 1183 2005 1187 2006
rect 1399 2010 1403 2011
rect 1399 2005 1403 2006
rect 910 1975 916 1976
rect 910 1971 911 1975
rect 915 1971 916 1975
rect 910 1970 916 1971
rect 918 1975 924 1976
rect 918 1971 919 1975
rect 923 1971 924 1975
rect 918 1970 924 1971
rect 862 1963 868 1964
rect 912 1963 914 1970
rect 231 1962 235 1963
rect 231 1957 235 1958
rect 351 1962 355 1963
rect 351 1957 355 1958
rect 463 1962 467 1963
rect 463 1957 467 1958
rect 575 1962 579 1963
rect 575 1957 579 1958
rect 687 1962 691 1963
rect 727 1962 731 1963
rect 766 1962 772 1963
rect 799 1962 803 1963
rect 687 1957 691 1958
rect 726 1957 732 1958
rect 726 1953 727 1957
rect 731 1953 732 1957
rect 726 1952 732 1953
rect 768 1952 770 1962
rect 855 1962 859 1963
rect 862 1959 863 1963
rect 867 1959 868 1963
rect 862 1958 868 1959
rect 911 1962 915 1963
rect 799 1957 803 1958
rect 854 1957 860 1958
rect 911 1957 915 1958
rect 854 1953 855 1957
rect 859 1953 860 1957
rect 854 1952 860 1953
rect 886 1955 892 1956
rect 766 1951 772 1952
rect 766 1947 767 1951
rect 771 1947 772 1951
rect 886 1951 887 1955
rect 891 1951 892 1955
rect 920 1952 922 1970
rect 983 1962 987 1963
rect 1103 1962 1107 1963
rect 1223 1962 1227 1963
rect 1335 1962 1339 1963
rect 982 1957 988 1958
rect 982 1953 983 1957
rect 987 1953 988 1957
rect 982 1952 988 1953
rect 1102 1957 1108 1958
rect 1102 1953 1103 1957
rect 1107 1953 1108 1957
rect 1102 1952 1108 1953
rect 1222 1957 1228 1958
rect 1222 1953 1223 1957
rect 1227 1953 1228 1957
rect 1222 1952 1228 1953
rect 1334 1957 1340 1958
rect 1334 1953 1335 1957
rect 1339 1953 1340 1957
rect 1334 1952 1340 1953
rect 1412 1952 1414 2034
rect 1610 2031 1611 2035
rect 1615 2031 1616 2035
rect 1610 2030 1616 2031
rect 1702 2035 1708 2036
rect 1702 2031 1703 2035
rect 1707 2031 1708 2035
rect 1702 2030 1708 2031
rect 1598 2016 1604 2017
rect 1598 2012 1599 2016
rect 1603 2012 1604 2016
rect 1598 2011 1604 2012
rect 1599 2010 1603 2011
rect 1599 2005 1603 2006
rect 1447 1962 1451 1963
rect 1567 1962 1571 1963
rect 1446 1957 1452 1958
rect 1446 1953 1447 1957
rect 1451 1953 1452 1957
rect 1446 1952 1452 1953
rect 1566 1957 1572 1958
rect 1566 1953 1567 1957
rect 1571 1953 1572 1957
rect 1612 1956 1614 2030
rect 1704 2024 1706 2030
rect 2024 2028 2026 2082
rect 2246 2079 2247 2083
rect 2251 2079 2252 2083
rect 2414 2083 2415 2087
rect 2419 2083 2420 2087
rect 2414 2082 2420 2083
rect 2470 2087 2476 2088
rect 2470 2083 2471 2087
rect 2475 2083 2476 2087
rect 2470 2082 2476 2083
rect 2246 2078 2252 2079
rect 2110 2060 2116 2061
rect 2110 2056 2111 2060
rect 2115 2056 2116 2060
rect 2110 2055 2116 2056
rect 2039 2054 2043 2055
rect 2039 2049 2043 2050
rect 2111 2054 2115 2055
rect 2111 2049 2115 2050
rect 2038 2048 2044 2049
rect 2038 2044 2039 2048
rect 2043 2044 2044 2048
rect 2038 2043 2044 2044
rect 2022 2027 2028 2028
rect 1630 2023 1636 2024
rect 1630 2019 1631 2023
rect 1635 2019 1636 2023
rect 1630 2018 1636 2019
rect 1670 2023 1676 2024
rect 1670 2019 1671 2023
rect 1675 2019 1676 2023
rect 1702 2023 1708 2024
rect 1670 2018 1676 2019
rect 1694 2019 1700 2020
rect 1632 2011 1634 2018
rect 1631 2010 1635 2011
rect 1672 2007 1674 2018
rect 1694 2015 1695 2019
rect 1699 2015 1700 2019
rect 1702 2019 1703 2023
rect 1707 2019 1708 2023
rect 2022 2023 2023 2027
rect 2027 2023 2028 2027
rect 2022 2022 2028 2023
rect 1702 2018 1708 2019
rect 2038 2019 2044 2020
rect 1694 2014 1700 2015
rect 2038 2015 2039 2019
rect 2043 2015 2044 2019
rect 2038 2014 2044 2015
rect 1696 2007 1698 2014
rect 2040 2007 2042 2014
rect 1631 2005 1635 2006
rect 1671 2006 1675 2007
rect 1632 1998 1634 2005
rect 1671 2001 1675 2002
rect 1695 2006 1699 2007
rect 1695 2001 1699 2002
rect 2039 2006 2043 2007
rect 2039 2001 2043 2002
rect 1672 1998 1674 2001
rect 1630 1997 1636 1998
rect 1630 1993 1631 1997
rect 1635 1993 1636 1997
rect 1630 1992 1636 1993
rect 1670 1997 1676 1998
rect 1670 1993 1671 1997
rect 1675 1993 1676 1997
rect 2248 1996 2250 2078
rect 2254 2060 2260 2061
rect 2254 2056 2255 2060
rect 2259 2056 2260 2060
rect 2254 2055 2260 2056
rect 2406 2060 2412 2061
rect 2406 2056 2407 2060
rect 2411 2056 2412 2060
rect 2406 2055 2412 2056
rect 2255 2054 2259 2055
rect 2255 2049 2259 2050
rect 2407 2054 2411 2055
rect 2407 2049 2411 2050
rect 2406 2048 2412 2049
rect 2406 2044 2407 2048
rect 2411 2044 2412 2048
rect 2406 2043 2412 2044
rect 2416 2024 2418 2082
rect 2728 2028 2730 2098
rect 2926 2095 2927 2099
rect 2931 2095 2932 2099
rect 2958 2099 2959 2103
rect 2963 2099 2964 2103
rect 3168 2100 3170 2178
rect 3191 2173 3195 2174
rect 3192 2170 3194 2173
rect 3190 2169 3196 2170
rect 3190 2165 3191 2169
rect 3195 2165 3196 2169
rect 3190 2164 3196 2165
rect 3190 2151 3196 2152
rect 3190 2147 3191 2151
rect 3195 2147 3196 2151
rect 3190 2146 3196 2147
rect 3192 2135 3194 2146
rect 3191 2134 3195 2135
rect 3191 2129 3195 2130
rect 3192 2122 3194 2129
rect 3190 2121 3196 2122
rect 3190 2117 3191 2121
rect 3195 2117 3196 2121
rect 3190 2116 3196 2117
rect 3190 2103 3196 2104
rect 2958 2098 2964 2099
rect 3158 2099 3164 2100
rect 2926 2094 2932 2095
rect 3158 2095 3159 2099
rect 3163 2095 3164 2099
rect 3158 2094 3164 2095
rect 3166 2099 3172 2100
rect 3166 2095 3167 2099
rect 3171 2095 3172 2099
rect 3190 2099 3191 2103
rect 3195 2099 3196 2103
rect 3190 2098 3196 2099
rect 3192 2095 3194 2098
rect 3166 2094 3172 2095
rect 3191 2094 3195 2095
rect 2927 2089 2931 2090
rect 3159 2089 3163 2090
rect 2767 2054 2771 2055
rect 2767 2049 2771 2050
rect 3135 2054 3139 2055
rect 3135 2049 3139 2050
rect 2766 2048 2772 2049
rect 2766 2044 2767 2048
rect 2771 2044 2772 2048
rect 2766 2043 2772 2044
rect 3134 2048 3140 2049
rect 3134 2044 3135 2048
rect 3139 2044 3140 2048
rect 3134 2043 3140 2044
rect 2726 2027 2732 2028
rect 2414 2023 2420 2024
rect 2406 2019 2412 2020
rect 2406 2015 2407 2019
rect 2411 2015 2412 2019
rect 2414 2019 2415 2023
rect 2419 2019 2420 2023
rect 2726 2023 2727 2027
rect 2731 2023 2732 2027
rect 2726 2022 2732 2023
rect 2854 2023 2860 2024
rect 2414 2018 2420 2019
rect 2406 2014 2412 2015
rect 2408 2007 2410 2014
rect 2416 2011 2418 2018
rect 2416 2009 2426 2011
rect 2263 2006 2267 2007
rect 2407 2006 2411 2007
rect 2415 2006 2419 2007
rect 2262 2001 2268 2002
rect 2407 2001 2411 2002
rect 2414 2001 2420 2002
rect 2262 1997 2263 2001
rect 2267 1997 2268 2001
rect 2262 1996 2268 1997
rect 2414 1997 2415 2001
rect 2419 1997 2420 2001
rect 2424 2000 2426 2009
rect 2559 2006 2563 2007
rect 2703 2006 2707 2007
rect 2558 2001 2564 2002
rect 2414 1996 2420 1997
rect 2422 1999 2428 2000
rect 1670 1992 1676 1993
rect 2246 1995 2252 1996
rect 2246 1991 2247 1995
rect 2251 1991 2252 1995
rect 2422 1995 2423 1999
rect 2427 1995 2428 1999
rect 2558 1997 2559 2001
rect 2563 1997 2564 2001
rect 2558 1996 2564 1997
rect 2702 2001 2708 2002
rect 2702 1997 2703 2001
rect 2707 1997 2708 2001
rect 2728 2000 2730 2022
rect 2766 2019 2772 2020
rect 2766 2015 2767 2019
rect 2771 2015 2772 2019
rect 2854 2019 2855 2023
rect 2859 2019 2860 2023
rect 2854 2018 2860 2019
rect 3134 2019 3140 2020
rect 2766 2014 2772 2015
rect 2768 2007 2770 2014
rect 2767 2006 2771 2007
rect 2839 2006 2843 2007
rect 2767 2001 2771 2002
rect 2838 2001 2844 2002
rect 2702 1996 2708 1997
rect 2726 1999 2732 2000
rect 2422 1994 2428 1995
rect 2550 1995 2556 1996
rect 2246 1990 2252 1991
rect 1630 1979 1636 1980
rect 1630 1975 1631 1979
rect 1635 1975 1636 1979
rect 1630 1974 1636 1975
rect 1670 1979 1676 1980
rect 1670 1975 1671 1979
rect 1675 1975 1676 1979
rect 1670 1974 1676 1975
rect 1632 1963 1634 1974
rect 1672 1967 1674 1974
rect 1671 1966 1675 1967
rect 1631 1962 1635 1963
rect 1671 1961 1675 1962
rect 2239 1966 2243 1967
rect 2239 1961 2243 1962
rect 1631 1957 1635 1958
rect 1566 1952 1572 1953
rect 1610 1955 1616 1956
rect 886 1950 892 1951
rect 918 1951 924 1952
rect 766 1946 772 1947
rect 726 1928 732 1929
rect 726 1924 727 1928
rect 731 1924 732 1928
rect 726 1923 732 1924
rect 728 1911 730 1923
rect 631 1910 635 1911
rect 631 1905 635 1906
rect 727 1910 731 1911
rect 727 1905 731 1906
rect 759 1910 763 1911
rect 759 1905 763 1906
rect 630 1904 636 1905
rect 630 1900 631 1904
rect 635 1900 636 1904
rect 630 1899 636 1900
rect 758 1904 764 1905
rect 758 1900 759 1904
rect 763 1900 764 1904
rect 758 1899 764 1900
rect 768 1876 770 1946
rect 854 1928 860 1929
rect 854 1924 855 1928
rect 859 1924 860 1928
rect 854 1923 860 1924
rect 856 1911 858 1923
rect 855 1910 859 1911
rect 855 1905 859 1906
rect 879 1910 883 1911
rect 879 1905 883 1906
rect 878 1904 884 1905
rect 878 1900 879 1904
rect 883 1900 884 1904
rect 878 1899 884 1900
rect 888 1880 890 1950
rect 918 1947 919 1951
rect 923 1947 924 1951
rect 918 1946 924 1947
rect 1006 1951 1012 1952
rect 1006 1947 1007 1951
rect 1011 1947 1012 1951
rect 1006 1946 1012 1947
rect 1126 1951 1132 1952
rect 1126 1947 1127 1951
rect 1131 1947 1132 1951
rect 1410 1951 1416 1952
rect 1126 1946 1132 1947
rect 1242 1947 1248 1948
rect 982 1928 988 1929
rect 982 1924 983 1928
rect 987 1924 988 1928
rect 982 1923 988 1924
rect 984 1911 986 1923
rect 983 1910 987 1911
rect 983 1905 987 1906
rect 999 1910 1003 1911
rect 999 1905 1003 1906
rect 998 1904 1004 1905
rect 998 1900 999 1904
rect 1003 1900 1004 1904
rect 998 1899 1004 1900
rect 1008 1880 1010 1946
rect 1102 1928 1108 1929
rect 1102 1924 1103 1928
rect 1107 1924 1108 1928
rect 1102 1923 1108 1924
rect 1104 1911 1106 1923
rect 1103 1910 1107 1911
rect 1103 1905 1107 1906
rect 1119 1910 1123 1911
rect 1119 1905 1123 1906
rect 1118 1904 1124 1905
rect 1118 1900 1119 1904
rect 1123 1900 1124 1904
rect 1118 1899 1124 1900
rect 1128 1880 1130 1946
rect 1242 1943 1243 1947
rect 1247 1943 1248 1947
rect 1242 1942 1248 1943
rect 1354 1947 1360 1948
rect 1354 1943 1355 1947
rect 1359 1943 1360 1947
rect 1410 1947 1411 1951
rect 1415 1947 1416 1951
rect 1410 1946 1416 1947
rect 1470 1951 1476 1952
rect 1470 1947 1471 1951
rect 1475 1947 1476 1951
rect 1610 1951 1611 1955
rect 1615 1951 1616 1955
rect 1632 1954 1634 1957
rect 1672 1954 1674 1961
rect 2238 1960 2244 1961
rect 2238 1956 2239 1960
rect 2243 1956 2244 1960
rect 2238 1955 2244 1956
rect 1610 1950 1616 1951
rect 1630 1953 1636 1954
rect 1630 1949 1631 1953
rect 1635 1949 1636 1953
rect 1630 1948 1636 1949
rect 1670 1953 1676 1954
rect 1670 1949 1671 1953
rect 1675 1949 1676 1953
rect 1670 1948 1676 1949
rect 1470 1946 1476 1947
rect 1354 1942 1360 1943
rect 1222 1928 1228 1929
rect 1222 1924 1223 1928
rect 1227 1924 1228 1928
rect 1222 1923 1228 1924
rect 1224 1911 1226 1923
rect 1223 1910 1227 1911
rect 1223 1905 1227 1906
rect 1231 1910 1235 1911
rect 1231 1905 1235 1906
rect 1230 1904 1236 1905
rect 1230 1900 1231 1904
rect 1235 1900 1236 1904
rect 1230 1899 1236 1900
rect 1244 1880 1246 1942
rect 1334 1928 1340 1929
rect 1334 1924 1335 1928
rect 1339 1924 1340 1928
rect 1334 1923 1340 1924
rect 1336 1911 1338 1923
rect 1335 1910 1339 1911
rect 1335 1905 1339 1906
rect 1343 1910 1347 1911
rect 1343 1905 1347 1906
rect 1342 1904 1348 1905
rect 1342 1900 1343 1904
rect 1347 1900 1348 1904
rect 1342 1899 1348 1900
rect 1356 1880 1358 1942
rect 1446 1928 1452 1929
rect 1446 1924 1447 1928
rect 1451 1924 1452 1928
rect 1446 1923 1452 1924
rect 1448 1911 1450 1923
rect 1447 1910 1451 1911
rect 1447 1905 1451 1906
rect 1463 1910 1467 1911
rect 1463 1905 1467 1906
rect 1462 1904 1468 1905
rect 1462 1900 1463 1904
rect 1467 1900 1468 1904
rect 1462 1899 1468 1900
rect 1472 1880 1474 1946
rect 1630 1935 1636 1936
rect 1630 1931 1631 1935
rect 1635 1931 1636 1935
rect 1630 1930 1636 1931
rect 1670 1935 1676 1936
rect 1670 1931 1671 1935
rect 1675 1931 1676 1935
rect 2248 1932 2250 1990
rect 2262 1972 2268 1973
rect 2262 1968 2263 1972
rect 2267 1968 2268 1972
rect 2262 1967 2268 1968
rect 2414 1972 2420 1973
rect 2414 1968 2415 1972
rect 2419 1968 2420 1972
rect 2414 1967 2420 1968
rect 2263 1966 2267 1967
rect 2263 1961 2267 1962
rect 2391 1966 2395 1967
rect 2391 1961 2395 1962
rect 2415 1966 2419 1967
rect 2415 1961 2419 1962
rect 2390 1960 2396 1961
rect 2390 1956 2391 1960
rect 2395 1956 2396 1960
rect 2390 1955 2396 1956
rect 2424 1936 2426 1994
rect 2550 1991 2551 1995
rect 2555 1991 2556 1995
rect 2726 1995 2727 1999
rect 2731 1995 2732 1999
rect 2838 1997 2839 2001
rect 2843 1997 2844 2001
rect 2838 1996 2844 1997
rect 2856 1996 2858 2018
rect 3134 2015 3135 2019
rect 3139 2015 3140 2019
rect 3134 2014 3140 2015
rect 3142 2019 3148 2020
rect 3142 2015 3143 2019
rect 3147 2015 3148 2019
rect 3142 2014 3148 2015
rect 3136 2007 3138 2014
rect 2975 2006 2979 2007
rect 3111 2006 3115 2007
rect 3135 2006 3139 2007
rect 2974 2001 2980 2002
rect 2974 1997 2975 2001
rect 2979 1997 2980 2001
rect 2974 1996 2980 1997
rect 3110 2001 3116 2002
rect 3135 2001 3139 2002
rect 3110 1997 3111 2001
rect 3115 1997 3116 2001
rect 3110 1996 3116 1997
rect 3144 1996 3146 2014
rect 3168 1996 3170 2094
rect 3191 2089 3195 2090
rect 3192 2086 3194 2089
rect 3190 2085 3196 2086
rect 3190 2081 3191 2085
rect 3195 2081 3196 2085
rect 3190 2080 3196 2081
rect 3190 2067 3196 2068
rect 3190 2063 3191 2067
rect 3195 2063 3196 2067
rect 3190 2062 3196 2063
rect 3192 2055 3194 2062
rect 3191 2054 3195 2055
rect 3191 2049 3195 2050
rect 3192 2042 3194 2049
rect 3190 2041 3196 2042
rect 3190 2037 3191 2041
rect 3195 2037 3196 2041
rect 3190 2036 3196 2037
rect 3190 2023 3196 2024
rect 3190 2019 3191 2023
rect 3195 2019 3196 2023
rect 3190 2018 3196 2019
rect 3192 2007 3194 2018
rect 3191 2006 3195 2007
rect 3191 2001 3195 2002
rect 3192 1998 3194 2001
rect 3190 1997 3196 1998
rect 2726 1994 2732 1995
rect 2856 1995 2864 1996
rect 2550 1990 2556 1991
rect 2543 1966 2547 1967
rect 2543 1961 2547 1962
rect 2542 1960 2548 1961
rect 2542 1956 2543 1960
rect 2547 1956 2548 1960
rect 2542 1955 2548 1956
rect 2552 1936 2554 1990
rect 2558 1972 2564 1973
rect 2558 1968 2559 1972
rect 2563 1968 2564 1972
rect 2558 1967 2564 1968
rect 2702 1972 2708 1973
rect 2702 1968 2703 1972
rect 2707 1968 2708 1972
rect 2702 1967 2708 1968
rect 2559 1966 2563 1967
rect 2559 1961 2563 1962
rect 2695 1966 2699 1967
rect 2695 1961 2699 1962
rect 2703 1966 2707 1967
rect 2703 1961 2707 1962
rect 2694 1960 2700 1961
rect 2694 1956 2695 1960
rect 2699 1956 2700 1960
rect 2694 1955 2700 1956
rect 2728 1936 2730 1994
rect 2856 1991 2859 1995
rect 2863 1991 2864 1995
rect 2856 1990 2864 1991
rect 3006 1995 3012 1996
rect 3006 1991 3007 1995
rect 3011 1991 3012 1995
rect 3006 1990 3012 1991
rect 3142 1995 3148 1996
rect 3142 1991 3143 1995
rect 3147 1991 3148 1995
rect 3142 1990 3148 1991
rect 3166 1995 3172 1996
rect 3166 1991 3167 1995
rect 3171 1991 3172 1995
rect 3190 1993 3191 1997
rect 3195 1993 3196 1997
rect 3190 1992 3196 1993
rect 3166 1990 3172 1991
rect 2838 1972 2844 1973
rect 2838 1968 2839 1972
rect 2843 1968 2844 1972
rect 2838 1967 2844 1968
rect 2839 1966 2843 1967
rect 2839 1961 2843 1962
rect 2847 1966 2851 1967
rect 2847 1961 2851 1962
rect 2846 1960 2852 1961
rect 2846 1956 2847 1960
rect 2851 1956 2852 1960
rect 2846 1955 2852 1956
rect 2856 1936 2858 1990
rect 2974 1972 2980 1973
rect 2974 1968 2975 1972
rect 2979 1968 2980 1972
rect 2974 1967 2980 1968
rect 2975 1966 2979 1967
rect 2975 1961 2979 1962
rect 2999 1966 3003 1967
rect 2999 1961 3003 1962
rect 2998 1960 3004 1961
rect 2998 1956 2999 1960
rect 3003 1956 3004 1960
rect 2998 1955 3004 1956
rect 3008 1936 3010 1990
rect 3110 1972 3116 1973
rect 3110 1968 3111 1972
rect 3115 1968 3116 1972
rect 3110 1967 3116 1968
rect 3111 1966 3115 1967
rect 3111 1961 3115 1962
rect 2422 1935 2428 1936
rect 1670 1930 1676 1931
rect 2238 1931 2244 1932
rect 1566 1928 1572 1929
rect 1566 1924 1567 1928
rect 1571 1924 1572 1928
rect 1566 1923 1572 1924
rect 1568 1911 1570 1923
rect 1632 1911 1634 1930
rect 1672 1923 1674 1930
rect 2238 1927 2239 1931
rect 2243 1927 2244 1931
rect 2238 1926 2244 1927
rect 2246 1931 2252 1932
rect 2246 1927 2247 1931
rect 2251 1927 2252 1931
rect 2246 1926 2252 1927
rect 2390 1931 2396 1932
rect 2390 1927 2391 1931
rect 2395 1927 2396 1931
rect 2422 1931 2423 1935
rect 2427 1931 2428 1935
rect 2550 1935 2556 1936
rect 2422 1930 2428 1931
rect 2542 1931 2548 1932
rect 2390 1926 2396 1927
rect 2240 1923 2242 1926
rect 1671 1922 1675 1923
rect 2151 1922 2155 1923
rect 2239 1922 2243 1923
rect 1671 1917 1675 1918
rect 2150 1917 2156 1918
rect 2239 1917 2243 1918
rect 1672 1914 1674 1917
rect 1670 1913 1676 1914
rect 1567 1910 1571 1911
rect 1567 1905 1571 1906
rect 1631 1910 1635 1911
rect 1670 1909 1671 1913
rect 1675 1909 1676 1913
rect 2150 1913 2151 1917
rect 2155 1913 2156 1917
rect 2150 1912 2156 1913
rect 2248 1912 2250 1926
rect 2392 1923 2394 1926
rect 2311 1922 2315 1923
rect 2391 1922 2395 1923
rect 2310 1917 2316 1918
rect 2391 1917 2395 1918
rect 2310 1913 2311 1917
rect 2315 1913 2316 1917
rect 2310 1912 2316 1913
rect 2424 1912 2426 1930
rect 2542 1927 2543 1931
rect 2547 1927 2548 1931
rect 2550 1931 2551 1935
rect 2555 1931 2556 1935
rect 2702 1935 2708 1936
rect 2550 1930 2556 1931
rect 2694 1931 2700 1932
rect 2542 1926 2548 1927
rect 2544 1923 2546 1926
rect 2471 1922 2475 1923
rect 2543 1922 2547 1923
rect 2470 1917 2476 1918
rect 2543 1917 2547 1918
rect 2470 1913 2471 1917
rect 2475 1913 2476 1917
rect 2470 1912 2476 1913
rect 1670 1908 1676 1909
rect 2158 1911 2164 1912
rect 2158 1907 2159 1911
rect 2163 1907 2164 1911
rect 2158 1906 2164 1907
rect 2246 1911 2252 1912
rect 2246 1907 2247 1911
rect 2251 1907 2252 1911
rect 2246 1906 2252 1907
rect 2422 1911 2428 1912
rect 2422 1907 2423 1911
rect 2427 1907 2428 1911
rect 2422 1906 2428 1907
rect 1631 1905 1635 1906
rect 1632 1898 1634 1905
rect 1630 1897 1636 1898
rect 1630 1893 1631 1897
rect 1635 1893 1636 1897
rect 1630 1892 1636 1893
rect 1670 1895 1676 1896
rect 1670 1891 1671 1895
rect 1675 1891 1676 1895
rect 1670 1890 1676 1891
rect 886 1879 892 1880
rect 630 1875 636 1876
rect 630 1871 631 1875
rect 635 1871 636 1875
rect 630 1870 636 1871
rect 638 1875 644 1876
rect 638 1871 639 1875
rect 643 1871 644 1875
rect 638 1870 644 1871
rect 758 1875 764 1876
rect 758 1871 759 1875
rect 763 1871 764 1875
rect 758 1870 764 1871
rect 766 1875 772 1876
rect 766 1871 767 1875
rect 771 1871 772 1875
rect 766 1870 772 1871
rect 878 1875 884 1876
rect 878 1871 879 1875
rect 883 1871 884 1875
rect 886 1875 887 1879
rect 891 1875 892 1879
rect 1006 1879 1012 1880
rect 886 1874 892 1875
rect 998 1875 1004 1876
rect 878 1870 884 1871
rect 632 1859 634 1870
rect 527 1858 531 1859
rect 631 1858 635 1859
rect 526 1853 532 1854
rect 631 1853 635 1854
rect 526 1849 527 1853
rect 531 1849 532 1853
rect 640 1852 642 1870
rect 760 1859 762 1870
rect 655 1858 659 1859
rect 759 1858 763 1859
rect 654 1853 660 1854
rect 759 1853 763 1854
rect 526 1848 532 1849
rect 638 1851 644 1852
rect 638 1847 639 1851
rect 643 1847 644 1851
rect 654 1849 655 1853
rect 659 1849 660 1853
rect 654 1848 660 1849
rect 768 1848 770 1870
rect 880 1859 882 1870
rect 775 1858 779 1859
rect 879 1858 883 1859
rect 774 1853 780 1854
rect 879 1853 883 1854
rect 774 1849 775 1853
rect 779 1849 780 1853
rect 774 1848 780 1849
rect 888 1848 890 1874
rect 998 1871 999 1875
rect 1003 1871 1004 1875
rect 1006 1875 1007 1879
rect 1011 1875 1012 1879
rect 1126 1879 1132 1880
rect 1006 1874 1012 1875
rect 1118 1875 1124 1876
rect 998 1870 1004 1871
rect 1000 1859 1002 1870
rect 895 1858 899 1859
rect 999 1858 1003 1859
rect 894 1853 900 1854
rect 999 1853 1003 1854
rect 894 1849 895 1853
rect 899 1849 900 1853
rect 894 1848 900 1849
rect 1008 1848 1010 1874
rect 1118 1871 1119 1875
rect 1123 1871 1124 1875
rect 1126 1875 1127 1879
rect 1131 1875 1132 1879
rect 1242 1879 1248 1880
rect 1230 1875 1236 1876
rect 1126 1874 1138 1875
rect 1128 1873 1138 1874
rect 1118 1870 1124 1871
rect 1120 1859 1122 1870
rect 1015 1858 1019 1859
rect 1119 1858 1123 1859
rect 1127 1858 1131 1859
rect 1014 1853 1020 1854
rect 1119 1853 1123 1854
rect 1126 1853 1132 1854
rect 1014 1849 1015 1853
rect 1019 1849 1020 1853
rect 1014 1848 1020 1849
rect 1126 1849 1127 1853
rect 1131 1849 1132 1853
rect 1136 1852 1138 1873
rect 1230 1871 1231 1875
rect 1235 1871 1236 1875
rect 1242 1875 1243 1879
rect 1247 1875 1248 1879
rect 1242 1874 1248 1875
rect 1254 1879 1260 1880
rect 1254 1875 1255 1879
rect 1259 1875 1260 1879
rect 1354 1879 1360 1880
rect 1254 1874 1260 1875
rect 1342 1875 1348 1876
rect 1230 1870 1236 1871
rect 1232 1859 1234 1870
rect 1231 1858 1235 1859
rect 1247 1858 1251 1859
rect 1231 1853 1235 1854
rect 1246 1853 1252 1854
rect 1126 1848 1132 1849
rect 1134 1851 1140 1852
rect 638 1846 644 1847
rect 686 1847 692 1848
rect 686 1843 687 1847
rect 691 1843 692 1847
rect 686 1842 692 1843
rect 766 1847 772 1848
rect 766 1843 767 1847
rect 771 1843 772 1847
rect 766 1842 772 1843
rect 806 1847 812 1848
rect 806 1843 807 1847
rect 811 1843 812 1847
rect 806 1842 812 1843
rect 886 1847 892 1848
rect 886 1843 887 1847
rect 891 1843 892 1847
rect 886 1842 892 1843
rect 926 1847 932 1848
rect 926 1843 927 1847
rect 931 1843 932 1847
rect 926 1842 932 1843
rect 1006 1847 1012 1848
rect 1006 1843 1007 1847
rect 1011 1843 1012 1847
rect 1006 1842 1012 1843
rect 1038 1847 1044 1848
rect 1038 1843 1039 1847
rect 1043 1843 1044 1847
rect 1134 1847 1135 1851
rect 1139 1847 1140 1851
rect 1246 1849 1247 1853
rect 1251 1849 1252 1853
rect 1256 1852 1258 1874
rect 1342 1871 1343 1875
rect 1347 1871 1348 1875
rect 1354 1875 1355 1879
rect 1359 1875 1360 1879
rect 1470 1879 1476 1880
rect 1354 1874 1360 1875
rect 1462 1875 1468 1876
rect 1342 1870 1348 1871
rect 1344 1859 1346 1870
rect 1343 1858 1347 1859
rect 1343 1853 1347 1854
rect 1246 1848 1252 1849
rect 1254 1851 1260 1852
rect 1134 1846 1140 1847
rect 1254 1847 1255 1851
rect 1259 1847 1260 1851
rect 1356 1848 1358 1874
rect 1462 1871 1463 1875
rect 1467 1871 1468 1875
rect 1470 1875 1471 1879
rect 1475 1875 1476 1879
rect 1470 1874 1476 1875
rect 1630 1879 1636 1880
rect 1672 1879 1674 1890
rect 2150 1888 2156 1889
rect 2150 1884 2151 1888
rect 2155 1884 2156 1888
rect 2150 1883 2156 1884
rect 2152 1879 2154 1883
rect 1630 1875 1631 1879
rect 1635 1875 1636 1879
rect 1630 1874 1636 1875
rect 1671 1878 1675 1879
rect 1462 1870 1468 1871
rect 1464 1859 1466 1870
rect 1632 1859 1634 1874
rect 1671 1873 1675 1874
rect 2071 1878 2075 1879
rect 2071 1873 2075 1874
rect 2151 1878 2155 1879
rect 2151 1873 2155 1874
rect 1672 1866 1674 1873
rect 2070 1872 2076 1873
rect 2070 1868 2071 1872
rect 2075 1868 2076 1872
rect 2070 1867 2076 1868
rect 1670 1865 1676 1866
rect 1670 1861 1671 1865
rect 1675 1861 1676 1865
rect 1670 1860 1676 1861
rect 1367 1858 1371 1859
rect 1463 1858 1467 1859
rect 1366 1853 1372 1854
rect 1463 1853 1467 1854
rect 1631 1858 1635 1859
rect 1631 1853 1635 1854
rect 1366 1849 1367 1853
rect 1371 1849 1372 1853
rect 1632 1850 1634 1853
rect 2160 1852 2162 1906
rect 2239 1878 2243 1879
rect 2239 1873 2243 1874
rect 2238 1872 2244 1873
rect 2238 1868 2239 1872
rect 2243 1868 2244 1872
rect 2238 1867 2244 1868
rect 2248 1852 2250 1906
rect 2310 1888 2316 1889
rect 2310 1884 2311 1888
rect 2315 1884 2316 1888
rect 2310 1883 2316 1884
rect 2312 1879 2314 1883
rect 2311 1878 2315 1879
rect 2311 1873 2315 1874
rect 2415 1878 2419 1879
rect 2415 1873 2419 1874
rect 2414 1872 2420 1873
rect 2414 1868 2415 1872
rect 2419 1868 2420 1872
rect 2414 1867 2420 1868
rect 2158 1851 2164 1852
rect 1366 1848 1372 1849
rect 1630 1849 1636 1850
rect 1254 1846 1260 1847
rect 1354 1847 1360 1848
rect 1038 1842 1044 1843
rect 526 1824 532 1825
rect 526 1820 527 1824
rect 531 1820 532 1824
rect 526 1819 532 1820
rect 654 1824 660 1825
rect 654 1820 655 1824
rect 659 1820 660 1824
rect 654 1819 660 1820
rect 528 1811 530 1819
rect 656 1811 658 1819
rect 423 1810 427 1811
rect 423 1805 427 1806
rect 527 1810 531 1811
rect 527 1805 531 1806
rect 551 1810 555 1811
rect 551 1805 555 1806
rect 655 1810 659 1811
rect 655 1805 659 1806
rect 679 1810 683 1811
rect 679 1805 683 1806
rect 422 1804 428 1805
rect 422 1800 423 1804
rect 427 1800 428 1804
rect 422 1799 428 1800
rect 550 1804 556 1805
rect 550 1800 551 1804
rect 555 1800 556 1804
rect 550 1799 556 1800
rect 678 1804 684 1805
rect 678 1800 679 1804
rect 683 1800 684 1804
rect 678 1799 684 1800
rect 688 1780 690 1842
rect 774 1824 780 1825
rect 774 1820 775 1824
rect 779 1820 780 1824
rect 774 1819 780 1820
rect 776 1811 778 1819
rect 775 1810 779 1811
rect 775 1805 779 1806
rect 799 1810 803 1811
rect 799 1805 803 1806
rect 798 1804 804 1805
rect 798 1800 799 1804
rect 803 1800 804 1804
rect 798 1799 804 1800
rect 808 1780 810 1842
rect 894 1824 900 1825
rect 894 1820 895 1824
rect 899 1820 900 1824
rect 894 1819 900 1820
rect 896 1811 898 1819
rect 895 1810 899 1811
rect 895 1805 899 1806
rect 919 1810 923 1811
rect 919 1805 923 1806
rect 918 1804 924 1805
rect 918 1800 919 1804
rect 923 1800 924 1804
rect 918 1799 924 1800
rect 928 1780 930 1842
rect 1014 1824 1020 1825
rect 1014 1820 1015 1824
rect 1019 1820 1020 1824
rect 1014 1819 1020 1820
rect 1016 1811 1018 1819
rect 1015 1810 1019 1811
rect 1015 1805 1019 1806
rect 1031 1810 1035 1811
rect 1031 1805 1035 1806
rect 1030 1804 1036 1805
rect 1030 1800 1031 1804
rect 1035 1800 1036 1804
rect 1030 1799 1036 1800
rect 1040 1780 1042 1842
rect 1126 1824 1132 1825
rect 1126 1820 1127 1824
rect 1131 1820 1132 1824
rect 1126 1819 1132 1820
rect 1128 1811 1130 1819
rect 1127 1810 1131 1811
rect 1127 1805 1131 1806
rect 1136 1784 1138 1846
rect 1246 1824 1252 1825
rect 1246 1820 1247 1824
rect 1251 1820 1252 1824
rect 1246 1819 1252 1820
rect 1248 1811 1250 1819
rect 1143 1810 1147 1811
rect 1143 1805 1147 1806
rect 1247 1810 1251 1811
rect 1247 1805 1251 1806
rect 1142 1804 1148 1805
rect 1142 1800 1143 1804
rect 1147 1800 1148 1804
rect 1142 1799 1148 1800
rect 1256 1784 1258 1846
rect 1354 1843 1355 1847
rect 1359 1843 1360 1847
rect 1630 1845 1631 1849
rect 1635 1845 1636 1849
rect 1630 1844 1636 1845
rect 1670 1847 1676 1848
rect 1354 1842 1360 1843
rect 1670 1843 1671 1847
rect 1675 1843 1676 1847
rect 2158 1847 2159 1851
rect 2163 1847 2164 1851
rect 2158 1846 2164 1847
rect 2246 1851 2252 1852
rect 2246 1847 2247 1851
rect 2251 1847 2252 1851
rect 2424 1848 2426 1906
rect 2470 1888 2476 1889
rect 2470 1884 2471 1888
rect 2475 1884 2476 1888
rect 2470 1883 2476 1884
rect 2472 1879 2474 1883
rect 2471 1878 2475 1879
rect 2471 1873 2475 1874
rect 2552 1852 2554 1930
rect 2694 1927 2695 1931
rect 2699 1927 2700 1931
rect 2702 1931 2703 1935
rect 2707 1931 2708 1935
rect 2702 1930 2708 1931
rect 2726 1935 2732 1936
rect 2726 1931 2727 1935
rect 2731 1931 2732 1935
rect 2854 1935 2860 1936
rect 2726 1930 2732 1931
rect 2846 1931 2852 1932
rect 2694 1926 2700 1927
rect 2696 1923 2698 1926
rect 2639 1922 2643 1923
rect 2695 1922 2699 1923
rect 2638 1917 2644 1918
rect 2695 1917 2699 1918
rect 2638 1913 2639 1917
rect 2643 1913 2644 1917
rect 2704 1916 2706 1930
rect 2846 1927 2847 1931
rect 2851 1927 2852 1931
rect 2854 1931 2855 1935
rect 2859 1931 2860 1935
rect 3006 1935 3012 1936
rect 2854 1930 2860 1931
rect 2998 1931 3004 1932
rect 2846 1926 2852 1927
rect 2848 1923 2850 1926
rect 2815 1922 2819 1923
rect 2847 1922 2851 1923
rect 2814 1917 2820 1918
rect 2847 1917 2851 1918
rect 2638 1912 2644 1913
rect 2702 1915 2708 1916
rect 2702 1911 2703 1915
rect 2707 1911 2708 1915
rect 2814 1913 2815 1917
rect 2819 1913 2820 1917
rect 2856 1916 2858 1930
rect 2998 1927 2999 1931
rect 3003 1927 3004 1931
rect 3006 1931 3007 1935
rect 3011 1931 3012 1935
rect 3006 1930 3012 1931
rect 2998 1926 3004 1927
rect 3000 1923 3002 1926
rect 2999 1922 3003 1923
rect 2998 1917 3004 1918
rect 2814 1912 2820 1913
rect 2822 1915 2828 1916
rect 2702 1910 2708 1911
rect 2822 1911 2823 1915
rect 2827 1911 2828 1915
rect 2822 1910 2828 1911
rect 2854 1915 2860 1916
rect 2854 1911 2855 1915
rect 2859 1911 2860 1915
rect 2998 1913 2999 1917
rect 3003 1913 3004 1917
rect 3008 1916 3010 1930
rect 3159 1922 3163 1923
rect 3158 1917 3164 1918
rect 2998 1912 3004 1913
rect 3006 1915 3012 1916
rect 2854 1910 2860 1911
rect 3006 1911 3007 1915
rect 3011 1911 3012 1915
rect 3158 1913 3159 1917
rect 3163 1913 3164 1917
rect 3168 1916 3170 1990
rect 3190 1979 3196 1980
rect 3190 1975 3191 1979
rect 3195 1975 3196 1979
rect 3190 1974 3196 1975
rect 3192 1967 3194 1974
rect 3191 1966 3195 1967
rect 3191 1961 3195 1962
rect 3192 1954 3194 1961
rect 3190 1953 3196 1954
rect 3190 1949 3191 1953
rect 3195 1949 3196 1953
rect 3190 1948 3196 1949
rect 3190 1935 3196 1936
rect 3190 1931 3191 1935
rect 3195 1931 3196 1935
rect 3190 1930 3196 1931
rect 3192 1923 3194 1930
rect 3191 1922 3195 1923
rect 3191 1917 3195 1918
rect 3158 1912 3164 1913
rect 3166 1915 3172 1916
rect 3006 1910 3012 1911
rect 3166 1911 3167 1915
rect 3171 1911 3172 1915
rect 3192 1914 3194 1917
rect 3166 1910 3172 1911
rect 3190 1913 3196 1914
rect 2638 1888 2644 1889
rect 2638 1884 2639 1888
rect 2643 1884 2644 1888
rect 2638 1883 2644 1884
rect 2814 1888 2820 1889
rect 2814 1884 2815 1888
rect 2819 1884 2820 1888
rect 2814 1883 2820 1884
rect 2640 1879 2642 1883
rect 2816 1879 2818 1883
rect 2599 1878 2603 1879
rect 2599 1873 2603 1874
rect 2639 1878 2643 1879
rect 2639 1873 2643 1874
rect 2791 1878 2795 1879
rect 2791 1873 2795 1874
rect 2815 1878 2819 1879
rect 2815 1873 2819 1874
rect 2598 1872 2604 1873
rect 2598 1868 2599 1872
rect 2603 1868 2604 1872
rect 2598 1867 2604 1868
rect 2790 1872 2796 1873
rect 2790 1868 2791 1872
rect 2795 1868 2796 1872
rect 2790 1867 2796 1868
rect 2550 1851 2556 1852
rect 2246 1846 2252 1847
rect 2422 1847 2428 1848
rect 1670 1842 1676 1843
rect 2070 1843 2076 1844
rect 1672 1839 1674 1842
rect 2070 1839 2071 1843
rect 2075 1839 2076 1843
rect 1671 1838 1675 1839
rect 1983 1838 1987 1839
rect 2070 1838 2076 1839
rect 2078 1843 2084 1844
rect 2078 1839 2079 1843
rect 2083 1839 2084 1843
rect 2078 1838 2084 1839
rect 2135 1838 2139 1839
rect 1671 1833 1675 1834
rect 1982 1833 1988 1834
rect 2071 1833 2075 1834
rect 1630 1831 1636 1832
rect 1630 1827 1631 1831
rect 1635 1827 1636 1831
rect 1672 1830 1674 1833
rect 1630 1826 1636 1827
rect 1670 1829 1676 1830
rect 1366 1824 1372 1825
rect 1366 1820 1367 1824
rect 1371 1820 1372 1824
rect 1366 1819 1372 1820
rect 1368 1811 1370 1819
rect 1632 1811 1634 1826
rect 1670 1825 1671 1829
rect 1675 1825 1676 1829
rect 1982 1829 1983 1833
rect 1987 1829 1988 1833
rect 1982 1828 1988 1829
rect 1670 1824 1676 1825
rect 1990 1827 1996 1828
rect 1990 1823 1991 1827
rect 1995 1823 1996 1827
rect 2080 1827 2082 1838
rect 2134 1833 2140 1834
rect 2134 1829 2135 1833
rect 2139 1829 2140 1833
rect 2134 1828 2140 1829
rect 2160 1828 2162 1846
rect 2238 1843 2244 1844
rect 2238 1839 2239 1843
rect 2243 1839 2244 1843
rect 2238 1838 2244 1839
rect 2239 1833 2243 1834
rect 2248 1828 2250 1846
rect 2414 1843 2420 1844
rect 2414 1839 2415 1843
rect 2419 1839 2420 1843
rect 2422 1843 2423 1847
rect 2427 1843 2428 1847
rect 2550 1847 2551 1851
rect 2555 1847 2556 1851
rect 2550 1846 2556 1847
rect 2590 1851 2596 1852
rect 2590 1847 2591 1851
rect 2595 1847 2596 1851
rect 2824 1848 2826 1910
rect 2998 1888 3004 1889
rect 2998 1884 2999 1888
rect 3003 1884 3004 1888
rect 2998 1883 3004 1884
rect 3000 1879 3002 1883
rect 2983 1878 2987 1879
rect 2983 1873 2987 1874
rect 2999 1878 3003 1879
rect 2999 1873 3003 1874
rect 2982 1872 2988 1873
rect 2982 1868 2983 1872
rect 2987 1868 2988 1872
rect 2982 1867 2988 1868
rect 3008 1848 3010 1910
rect 3158 1888 3164 1889
rect 3158 1884 3159 1888
rect 3163 1884 3164 1888
rect 3158 1883 3164 1884
rect 3160 1879 3162 1883
rect 3159 1878 3163 1879
rect 3159 1873 3163 1874
rect 3158 1872 3164 1873
rect 3158 1868 3159 1872
rect 3163 1868 3164 1872
rect 3158 1867 3164 1868
rect 3168 1848 3170 1910
rect 3190 1909 3191 1913
rect 3195 1909 3196 1913
rect 3190 1908 3196 1909
rect 3190 1895 3196 1896
rect 3190 1891 3191 1895
rect 3195 1891 3196 1895
rect 3190 1890 3196 1891
rect 3192 1879 3194 1890
rect 3191 1878 3195 1879
rect 3191 1873 3195 1874
rect 3192 1866 3194 1873
rect 3190 1865 3196 1866
rect 3190 1861 3191 1865
rect 3195 1861 3196 1865
rect 3190 1860 3196 1861
rect 2590 1846 2596 1847
rect 2822 1847 2828 1848
rect 2422 1842 2428 1843
rect 2287 1838 2291 1839
rect 2414 1838 2420 1839
rect 2286 1833 2292 1834
rect 2415 1833 2419 1834
rect 2286 1829 2287 1833
rect 2291 1829 2292 1833
rect 2286 1828 2292 1829
rect 2424 1828 2426 1842
rect 2431 1838 2435 1839
rect 2583 1838 2587 1839
rect 2430 1833 2436 1834
rect 2430 1829 2431 1833
rect 2435 1829 2436 1833
rect 2430 1828 2436 1829
rect 2582 1833 2588 1834
rect 2582 1829 2583 1833
rect 2587 1829 2588 1833
rect 2592 1832 2594 1846
rect 2598 1843 2604 1844
rect 2598 1839 2599 1843
rect 2603 1839 2604 1843
rect 2790 1843 2796 1844
rect 2790 1839 2791 1843
rect 2795 1839 2796 1843
rect 2822 1843 2823 1847
rect 2827 1843 2828 1847
rect 3006 1847 3012 1848
rect 2822 1842 2828 1843
rect 2982 1843 2988 1844
rect 2598 1838 2604 1839
rect 2735 1838 2739 1839
rect 2790 1838 2796 1839
rect 2982 1839 2983 1843
rect 2987 1839 2988 1843
rect 3006 1843 3007 1847
rect 3011 1843 3012 1847
rect 3166 1847 3172 1848
rect 3006 1842 3012 1843
rect 3158 1843 3164 1844
rect 2982 1838 2988 1839
rect 2599 1833 2603 1834
rect 2734 1833 2740 1834
rect 2791 1833 2795 1834
rect 2983 1833 2987 1834
rect 2582 1828 2588 1829
rect 2590 1831 2596 1832
rect 2086 1827 2092 1828
rect 2080 1825 2087 1827
rect 1990 1822 1996 1823
rect 2086 1823 2087 1825
rect 2091 1823 2092 1827
rect 2086 1822 2092 1823
rect 2158 1827 2164 1828
rect 2158 1823 2159 1827
rect 2163 1823 2164 1827
rect 2158 1822 2164 1823
rect 2246 1827 2252 1828
rect 2246 1823 2247 1827
rect 2251 1823 2252 1827
rect 2246 1822 2252 1823
rect 2422 1827 2428 1828
rect 2422 1823 2423 1827
rect 2427 1823 2428 1827
rect 2422 1822 2428 1823
rect 2494 1827 2500 1828
rect 2494 1823 2495 1827
rect 2499 1823 2500 1827
rect 2590 1827 2591 1831
rect 2595 1827 2596 1831
rect 2734 1829 2735 1833
rect 2739 1829 2740 1833
rect 2734 1828 2740 1829
rect 2742 1831 2748 1832
rect 2590 1826 2596 1827
rect 2742 1827 2743 1831
rect 2747 1827 2748 1831
rect 2742 1826 2748 1827
rect 2494 1822 2500 1823
rect 1670 1811 1676 1812
rect 1263 1810 1267 1811
rect 1263 1805 1267 1806
rect 1367 1810 1371 1811
rect 1367 1805 1371 1806
rect 1631 1810 1635 1811
rect 1670 1807 1671 1811
rect 1675 1807 1676 1811
rect 1670 1806 1676 1807
rect 1631 1805 1635 1806
rect 1262 1804 1268 1805
rect 1262 1800 1263 1804
rect 1267 1800 1268 1804
rect 1262 1799 1268 1800
rect 1632 1798 1634 1805
rect 1672 1799 1674 1806
rect 1982 1804 1988 1805
rect 1982 1800 1983 1804
rect 1987 1800 1988 1804
rect 1982 1799 1988 1800
rect 1671 1798 1675 1799
rect 1630 1797 1636 1798
rect 1630 1793 1631 1797
rect 1635 1793 1636 1797
rect 1671 1793 1675 1794
rect 1903 1798 1907 1799
rect 1903 1793 1907 1794
rect 1983 1798 1987 1799
rect 1983 1793 1987 1794
rect 1630 1792 1636 1793
rect 1672 1786 1674 1793
rect 1902 1792 1908 1793
rect 1902 1788 1903 1792
rect 1907 1788 1908 1792
rect 1902 1787 1908 1788
rect 1670 1785 1676 1786
rect 1134 1783 1140 1784
rect 686 1779 692 1780
rect 422 1775 428 1776
rect 422 1771 423 1775
rect 427 1771 428 1775
rect 422 1770 428 1771
rect 430 1775 436 1776
rect 430 1771 431 1775
rect 435 1771 436 1775
rect 430 1770 436 1771
rect 550 1775 556 1776
rect 550 1771 551 1775
rect 555 1771 556 1775
rect 550 1770 556 1771
rect 558 1775 564 1776
rect 558 1771 559 1775
rect 563 1771 564 1775
rect 558 1770 564 1771
rect 678 1775 684 1776
rect 678 1771 679 1775
rect 683 1771 684 1775
rect 686 1775 687 1779
rect 691 1775 692 1779
rect 806 1779 812 1780
rect 686 1774 692 1775
rect 798 1775 804 1776
rect 678 1770 684 1771
rect 798 1771 799 1775
rect 803 1771 804 1775
rect 806 1775 807 1779
rect 811 1775 812 1779
rect 926 1779 932 1780
rect 806 1774 812 1775
rect 918 1775 924 1776
rect 798 1770 804 1771
rect 918 1771 919 1775
rect 923 1771 924 1775
rect 926 1775 927 1779
rect 931 1775 932 1779
rect 1038 1779 1044 1780
rect 926 1774 932 1775
rect 1030 1775 1036 1776
rect 918 1770 924 1771
rect 1030 1771 1031 1775
rect 1035 1771 1036 1775
rect 1038 1775 1039 1779
rect 1043 1775 1044 1779
rect 1134 1779 1135 1783
rect 1139 1779 1140 1783
rect 1134 1778 1140 1779
rect 1254 1783 1260 1784
rect 1254 1779 1255 1783
rect 1259 1779 1260 1783
rect 1670 1781 1671 1785
rect 1675 1781 1676 1785
rect 1670 1780 1676 1781
rect 1254 1778 1260 1779
rect 1630 1779 1636 1780
rect 1038 1774 1044 1775
rect 1142 1775 1148 1776
rect 1030 1770 1036 1771
rect 1142 1771 1143 1775
rect 1147 1771 1148 1775
rect 1142 1770 1148 1771
rect 1262 1775 1268 1776
rect 1262 1771 1263 1775
rect 1267 1771 1268 1775
rect 1630 1775 1631 1779
rect 1635 1775 1636 1779
rect 1630 1774 1636 1775
rect 1262 1770 1268 1771
rect 424 1759 426 1770
rect 327 1758 331 1759
rect 423 1758 427 1759
rect 326 1753 332 1754
rect 423 1753 427 1754
rect 326 1749 327 1753
rect 331 1749 332 1753
rect 326 1748 332 1749
rect 432 1748 434 1770
rect 552 1759 554 1770
rect 455 1758 459 1759
rect 551 1758 555 1759
rect 454 1753 460 1754
rect 551 1753 555 1754
rect 454 1749 455 1753
rect 459 1749 460 1753
rect 454 1748 460 1749
rect 560 1748 562 1770
rect 680 1759 682 1770
rect 800 1759 802 1770
rect 920 1759 922 1770
rect 1032 1759 1034 1770
rect 1144 1759 1146 1770
rect 1264 1759 1266 1770
rect 1632 1759 1634 1774
rect 1992 1768 1994 1822
rect 2079 1798 2083 1799
rect 2079 1793 2083 1794
rect 2078 1792 2084 1793
rect 2078 1788 2079 1792
rect 2083 1788 2084 1792
rect 2078 1787 2084 1788
rect 2088 1772 2090 1822
rect 2134 1804 2140 1805
rect 2134 1800 2135 1804
rect 2139 1800 2140 1804
rect 2134 1799 2140 1800
rect 2135 1798 2139 1799
rect 2135 1793 2139 1794
rect 2248 1772 2250 1822
rect 2286 1804 2292 1805
rect 2286 1800 2287 1804
rect 2291 1800 2292 1804
rect 2286 1799 2292 1800
rect 2430 1804 2436 1805
rect 2430 1800 2431 1804
rect 2435 1800 2436 1804
rect 2430 1799 2436 1800
rect 2271 1798 2275 1799
rect 2271 1793 2275 1794
rect 2287 1798 2291 1799
rect 2287 1793 2291 1794
rect 2431 1798 2435 1799
rect 2431 1793 2435 1794
rect 2487 1798 2491 1799
rect 2487 1793 2491 1794
rect 2270 1792 2276 1793
rect 2270 1788 2271 1792
rect 2275 1788 2276 1792
rect 2270 1787 2276 1788
rect 2486 1792 2492 1793
rect 2486 1788 2487 1792
rect 2491 1788 2492 1792
rect 2486 1787 2492 1788
rect 2086 1771 2092 1772
rect 1670 1767 1676 1768
rect 1670 1763 1671 1767
rect 1675 1763 1676 1767
rect 1990 1767 1996 1768
rect 1670 1762 1676 1763
rect 1902 1763 1908 1764
rect 575 1758 579 1759
rect 679 1758 683 1759
rect 695 1758 699 1759
rect 799 1758 803 1759
rect 815 1758 819 1759
rect 919 1758 923 1759
rect 927 1758 931 1759
rect 1031 1758 1035 1759
rect 1039 1758 1043 1759
rect 1143 1758 1147 1759
rect 1159 1758 1163 1759
rect 1263 1758 1267 1759
rect 574 1753 580 1754
rect 679 1753 683 1754
rect 694 1753 700 1754
rect 799 1753 803 1754
rect 814 1753 820 1754
rect 919 1753 923 1754
rect 926 1753 932 1754
rect 1031 1753 1035 1754
rect 1038 1753 1044 1754
rect 1143 1753 1147 1754
rect 1158 1753 1164 1754
rect 1263 1753 1267 1754
rect 1631 1758 1635 1759
rect 1631 1753 1635 1754
rect 574 1749 575 1753
rect 579 1749 580 1753
rect 574 1748 580 1749
rect 694 1749 695 1753
rect 699 1749 700 1753
rect 694 1748 700 1749
rect 814 1749 815 1753
rect 819 1749 820 1753
rect 814 1748 820 1749
rect 926 1749 927 1753
rect 931 1749 932 1753
rect 926 1748 932 1749
rect 1038 1749 1039 1753
rect 1043 1749 1044 1753
rect 1038 1748 1044 1749
rect 1158 1749 1159 1753
rect 1163 1749 1164 1753
rect 1632 1750 1634 1753
rect 1672 1751 1674 1762
rect 1902 1759 1903 1763
rect 1907 1759 1908 1763
rect 1990 1763 1991 1767
rect 1995 1763 1996 1767
rect 2086 1767 2087 1771
rect 2091 1767 2092 1771
rect 2086 1766 2092 1767
rect 2246 1771 2252 1772
rect 2246 1767 2247 1771
rect 2251 1767 2252 1771
rect 2496 1768 2498 1822
rect 2582 1804 2588 1805
rect 2582 1800 2583 1804
rect 2587 1800 2588 1804
rect 2582 1799 2588 1800
rect 2734 1804 2740 1805
rect 2734 1800 2735 1804
rect 2739 1800 2740 1804
rect 2734 1799 2740 1800
rect 2583 1798 2587 1799
rect 2583 1793 2587 1794
rect 2711 1798 2715 1799
rect 2711 1793 2715 1794
rect 2735 1798 2739 1799
rect 2735 1793 2739 1794
rect 2710 1792 2716 1793
rect 2710 1788 2711 1792
rect 2715 1788 2716 1792
rect 2710 1787 2716 1788
rect 2744 1768 2746 1826
rect 2943 1798 2947 1799
rect 2943 1793 2947 1794
rect 2942 1792 2948 1793
rect 2942 1788 2943 1792
rect 2947 1788 2948 1792
rect 2942 1787 2948 1788
rect 3008 1768 3010 1842
rect 3158 1839 3159 1843
rect 3163 1839 3164 1843
rect 3166 1843 3167 1847
rect 3171 1843 3172 1847
rect 3166 1842 3172 1843
rect 3190 1847 3196 1848
rect 3190 1843 3191 1847
rect 3195 1843 3196 1847
rect 3190 1842 3196 1843
rect 3158 1838 3164 1839
rect 3159 1833 3163 1834
rect 3159 1798 3163 1799
rect 3159 1793 3163 1794
rect 3158 1792 3164 1793
rect 3158 1788 3159 1792
rect 3163 1788 3164 1792
rect 3158 1787 3164 1788
rect 3168 1768 3170 1842
rect 3192 1839 3194 1842
rect 3191 1838 3195 1839
rect 3191 1833 3195 1834
rect 3192 1830 3194 1833
rect 3190 1829 3196 1830
rect 3190 1825 3191 1829
rect 3195 1825 3196 1829
rect 3190 1824 3196 1825
rect 3190 1811 3196 1812
rect 3190 1807 3191 1811
rect 3195 1807 3196 1811
rect 3190 1806 3196 1807
rect 3192 1799 3194 1806
rect 3191 1798 3195 1799
rect 3191 1793 3195 1794
rect 3192 1786 3194 1793
rect 3190 1785 3196 1786
rect 3190 1781 3191 1785
rect 3195 1781 3196 1785
rect 3190 1780 3196 1781
rect 2246 1766 2252 1767
rect 2494 1767 2500 1768
rect 1990 1762 1996 1763
rect 2078 1763 2084 1764
rect 1902 1758 1908 1759
rect 2078 1759 2079 1763
rect 2083 1759 2084 1763
rect 2078 1758 2084 1759
rect 2270 1763 2276 1764
rect 2270 1759 2271 1763
rect 2275 1759 2276 1763
rect 2270 1758 2276 1759
rect 2486 1763 2492 1764
rect 2486 1759 2487 1763
rect 2491 1759 2492 1763
rect 2494 1763 2495 1767
rect 2499 1763 2500 1767
rect 2742 1767 2748 1768
rect 2494 1762 2500 1763
rect 2710 1763 2716 1764
rect 2486 1758 2492 1759
rect 2710 1759 2711 1763
rect 2715 1759 2716 1763
rect 2742 1763 2743 1767
rect 2747 1763 2748 1767
rect 2950 1767 2956 1768
rect 2742 1762 2748 1763
rect 2942 1763 2948 1764
rect 2710 1758 2716 1759
rect 2942 1759 2943 1763
rect 2947 1759 2948 1763
rect 2950 1763 2951 1767
rect 2955 1763 2956 1767
rect 2950 1762 2956 1763
rect 3006 1767 3012 1768
rect 3006 1763 3007 1767
rect 3011 1763 3012 1767
rect 3166 1767 3172 1768
rect 3006 1762 3012 1763
rect 3158 1763 3164 1764
rect 2942 1758 2948 1759
rect 1904 1751 1906 1758
rect 2080 1751 2082 1758
rect 2272 1751 2274 1758
rect 2488 1751 2490 1758
rect 2712 1751 2714 1758
rect 2944 1751 2946 1758
rect 1671 1750 1675 1751
rect 1158 1748 1164 1749
rect 1630 1749 1636 1750
rect 334 1747 340 1748
rect 334 1743 335 1747
rect 339 1743 340 1747
rect 334 1742 340 1743
rect 430 1747 436 1748
rect 430 1743 431 1747
rect 435 1743 436 1747
rect 430 1742 436 1743
rect 558 1747 564 1748
rect 558 1743 559 1747
rect 563 1743 564 1747
rect 558 1742 564 1743
rect 718 1747 724 1748
rect 718 1743 719 1747
rect 723 1743 724 1747
rect 718 1742 724 1743
rect 822 1747 828 1748
rect 822 1743 823 1747
rect 827 1746 828 1747
rect 950 1747 956 1748
rect 827 1744 834 1746
rect 827 1743 828 1744
rect 822 1742 828 1743
rect 326 1724 332 1725
rect 326 1720 327 1724
rect 331 1720 332 1724
rect 326 1719 332 1720
rect 328 1707 330 1719
rect 223 1706 227 1707
rect 223 1701 227 1702
rect 327 1706 331 1707
rect 327 1701 331 1702
rect 222 1700 228 1701
rect 222 1696 223 1700
rect 227 1696 228 1700
rect 222 1695 228 1696
rect 222 1671 228 1672
rect 222 1667 223 1671
rect 227 1667 228 1671
rect 222 1666 228 1667
rect 230 1671 236 1672
rect 230 1667 231 1671
rect 235 1667 236 1671
rect 230 1666 236 1667
rect 224 1655 226 1666
rect 223 1654 227 1655
rect 223 1649 227 1650
rect 232 1644 234 1666
rect 336 1664 338 1742
rect 454 1724 460 1725
rect 454 1720 455 1724
rect 459 1720 460 1724
rect 454 1719 460 1720
rect 574 1724 580 1725
rect 574 1720 575 1724
rect 579 1720 580 1724
rect 574 1719 580 1720
rect 694 1724 700 1725
rect 694 1720 695 1724
rect 699 1720 700 1724
rect 694 1719 700 1720
rect 456 1707 458 1719
rect 576 1707 578 1719
rect 696 1707 698 1719
rect 351 1706 355 1707
rect 351 1701 355 1702
rect 455 1706 459 1707
rect 455 1701 459 1702
rect 471 1706 475 1707
rect 471 1701 475 1702
rect 575 1706 579 1707
rect 575 1701 579 1702
rect 591 1706 595 1707
rect 591 1701 595 1702
rect 695 1706 699 1707
rect 695 1701 699 1702
rect 711 1706 715 1707
rect 711 1701 715 1702
rect 350 1700 356 1701
rect 350 1696 351 1700
rect 355 1696 356 1700
rect 350 1695 356 1696
rect 470 1700 476 1701
rect 470 1696 471 1700
rect 475 1696 476 1700
rect 470 1695 476 1696
rect 590 1700 596 1701
rect 590 1696 591 1700
rect 595 1696 596 1700
rect 590 1695 596 1696
rect 710 1700 716 1701
rect 710 1696 711 1700
rect 715 1696 716 1700
rect 710 1695 716 1696
rect 720 1676 722 1742
rect 814 1724 820 1725
rect 814 1720 815 1724
rect 819 1720 820 1724
rect 814 1719 820 1720
rect 816 1707 818 1719
rect 815 1706 819 1707
rect 815 1701 819 1702
rect 823 1706 827 1707
rect 823 1701 827 1702
rect 822 1700 828 1701
rect 822 1696 823 1700
rect 827 1696 828 1700
rect 822 1695 828 1696
rect 832 1676 834 1744
rect 950 1743 951 1747
rect 955 1743 956 1747
rect 950 1742 956 1743
rect 1166 1747 1172 1748
rect 1166 1743 1167 1747
rect 1171 1743 1172 1747
rect 1630 1745 1631 1749
rect 1635 1745 1636 1749
rect 1815 1750 1819 1751
rect 1903 1750 1907 1751
rect 1967 1750 1971 1751
rect 2079 1750 2083 1751
rect 2127 1750 2131 1751
rect 2271 1750 2275 1751
rect 2303 1750 2307 1751
rect 2487 1750 2491 1751
rect 2503 1750 2507 1751
rect 2711 1750 2715 1751
rect 2935 1750 2939 1751
rect 2943 1750 2947 1751
rect 1671 1745 1675 1746
rect 1814 1745 1820 1746
rect 1903 1745 1907 1746
rect 1966 1745 1972 1746
rect 2079 1745 2083 1746
rect 2126 1745 2132 1746
rect 2271 1745 2275 1746
rect 2302 1745 2308 1746
rect 2487 1745 2491 1746
rect 2502 1745 2508 1746
rect 1630 1744 1636 1745
rect 1166 1742 1172 1743
rect 1672 1742 1674 1745
rect 926 1724 932 1725
rect 926 1720 927 1724
rect 931 1720 932 1724
rect 926 1719 932 1720
rect 928 1707 930 1719
rect 927 1706 931 1707
rect 927 1701 931 1702
rect 943 1706 947 1707
rect 943 1701 947 1702
rect 942 1700 948 1701
rect 942 1696 943 1700
rect 947 1696 948 1700
rect 942 1695 948 1696
rect 926 1679 932 1680
rect 718 1675 724 1676
rect 350 1671 356 1672
rect 350 1667 351 1671
rect 355 1667 356 1671
rect 350 1666 356 1667
rect 470 1671 476 1672
rect 470 1667 471 1671
rect 475 1667 476 1671
rect 470 1666 476 1667
rect 478 1671 484 1672
rect 478 1667 479 1671
rect 483 1667 484 1671
rect 478 1666 484 1667
rect 590 1671 596 1672
rect 590 1667 591 1671
rect 595 1667 596 1671
rect 590 1666 596 1667
rect 598 1671 604 1672
rect 598 1667 599 1671
rect 603 1667 604 1671
rect 598 1666 604 1667
rect 710 1671 716 1672
rect 710 1667 711 1671
rect 715 1667 716 1671
rect 718 1671 719 1675
rect 723 1671 724 1675
rect 830 1675 836 1676
rect 718 1670 724 1671
rect 822 1671 828 1672
rect 710 1666 716 1667
rect 310 1663 316 1664
rect 310 1659 311 1663
rect 315 1659 316 1663
rect 310 1658 316 1659
rect 334 1663 340 1664
rect 334 1659 335 1663
rect 339 1659 340 1663
rect 334 1658 340 1659
rect 247 1654 251 1655
rect 246 1649 252 1650
rect 246 1645 247 1649
rect 251 1645 252 1649
rect 246 1644 252 1645
rect 312 1644 314 1658
rect 352 1655 354 1666
rect 472 1655 474 1666
rect 351 1654 355 1655
rect 383 1654 387 1655
rect 471 1654 475 1655
rect 351 1649 355 1650
rect 382 1649 388 1650
rect 471 1649 475 1650
rect 382 1645 383 1649
rect 387 1645 388 1649
rect 480 1648 482 1666
rect 592 1655 594 1666
rect 535 1654 539 1655
rect 591 1654 595 1655
rect 534 1649 540 1650
rect 591 1649 595 1650
rect 382 1644 388 1645
rect 478 1647 484 1648
rect 110 1640 116 1641
rect 142 1643 148 1644
rect 142 1639 143 1643
rect 147 1639 148 1643
rect 142 1638 148 1639
rect 230 1643 236 1644
rect 230 1639 231 1643
rect 235 1639 236 1643
rect 230 1638 236 1639
rect 310 1643 316 1644
rect 310 1639 311 1643
rect 315 1639 316 1643
rect 478 1643 479 1647
rect 483 1643 484 1647
rect 534 1645 535 1649
rect 539 1645 540 1649
rect 534 1644 540 1645
rect 600 1644 602 1666
rect 712 1655 714 1666
rect 711 1654 715 1655
rect 710 1649 716 1650
rect 710 1645 711 1649
rect 715 1645 716 1649
rect 720 1648 722 1670
rect 822 1667 823 1671
rect 827 1667 828 1671
rect 830 1671 831 1675
rect 835 1671 836 1675
rect 926 1675 927 1679
rect 931 1675 932 1679
rect 952 1676 954 1742
rect 1038 1724 1044 1725
rect 1038 1720 1039 1724
rect 1043 1720 1044 1724
rect 1038 1719 1044 1720
rect 1158 1724 1164 1725
rect 1158 1720 1159 1724
rect 1163 1720 1164 1724
rect 1158 1719 1164 1720
rect 1040 1707 1042 1719
rect 1160 1707 1162 1719
rect 1039 1706 1043 1707
rect 1039 1701 1043 1702
rect 1063 1706 1067 1707
rect 1063 1701 1067 1702
rect 1159 1706 1163 1707
rect 1159 1701 1163 1702
rect 1062 1700 1068 1701
rect 1062 1696 1063 1700
rect 1067 1696 1068 1700
rect 1062 1695 1068 1696
rect 926 1674 932 1675
rect 950 1675 956 1676
rect 830 1670 836 1671
rect 822 1666 828 1667
rect 824 1655 826 1666
rect 823 1654 827 1655
rect 919 1654 923 1655
rect 823 1649 827 1650
rect 918 1649 924 1650
rect 710 1644 716 1645
rect 718 1647 724 1648
rect 478 1642 484 1643
rect 598 1643 604 1644
rect 310 1638 316 1639
rect 110 1627 116 1628
rect 110 1623 111 1627
rect 115 1623 116 1627
rect 110 1622 116 1623
rect 112 1607 114 1622
rect 134 1620 140 1621
rect 134 1616 135 1620
rect 139 1616 140 1620
rect 134 1615 140 1616
rect 136 1607 138 1615
rect 111 1606 115 1607
rect 111 1601 115 1602
rect 135 1606 139 1607
rect 135 1601 139 1602
rect 112 1594 114 1601
rect 134 1600 140 1601
rect 134 1596 135 1600
rect 139 1596 140 1600
rect 134 1595 140 1596
rect 110 1593 116 1594
rect 110 1589 111 1593
rect 115 1589 116 1593
rect 110 1588 116 1589
rect 144 1576 146 1638
rect 246 1620 252 1621
rect 246 1616 247 1620
rect 251 1616 252 1620
rect 246 1615 252 1616
rect 248 1607 250 1615
rect 247 1606 251 1607
rect 247 1601 251 1602
rect 303 1606 307 1607
rect 303 1601 307 1602
rect 302 1600 308 1601
rect 302 1596 303 1600
rect 307 1596 308 1600
rect 302 1595 308 1596
rect 312 1576 314 1638
rect 382 1620 388 1621
rect 382 1616 383 1620
rect 387 1616 388 1620
rect 382 1615 388 1616
rect 384 1607 386 1615
rect 383 1606 387 1607
rect 383 1601 387 1602
rect 480 1580 482 1642
rect 598 1639 599 1643
rect 603 1639 604 1643
rect 718 1643 719 1647
rect 723 1643 724 1647
rect 918 1645 919 1649
rect 923 1645 924 1649
rect 928 1648 930 1674
rect 942 1671 948 1672
rect 942 1667 943 1671
rect 947 1667 948 1671
rect 950 1671 951 1675
rect 955 1671 956 1675
rect 950 1670 956 1671
rect 1062 1671 1068 1672
rect 942 1666 948 1667
rect 1062 1667 1063 1671
rect 1067 1667 1068 1671
rect 1062 1666 1068 1667
rect 1070 1671 1076 1672
rect 1070 1667 1071 1671
rect 1075 1667 1076 1671
rect 1070 1666 1076 1667
rect 944 1655 946 1666
rect 1064 1655 1066 1666
rect 943 1654 947 1655
rect 943 1649 947 1650
rect 1063 1654 1067 1655
rect 1063 1649 1067 1650
rect 918 1644 924 1645
rect 926 1647 932 1648
rect 718 1642 724 1643
rect 926 1643 927 1647
rect 931 1643 932 1647
rect 926 1642 932 1643
rect 598 1638 604 1639
rect 534 1620 540 1621
rect 534 1616 535 1620
rect 539 1616 540 1620
rect 534 1615 540 1616
rect 710 1620 716 1621
rect 710 1616 711 1620
rect 715 1616 716 1620
rect 710 1615 716 1616
rect 536 1607 538 1615
rect 712 1607 714 1615
rect 503 1606 507 1607
rect 503 1601 507 1602
rect 535 1606 539 1607
rect 535 1601 539 1602
rect 695 1606 699 1607
rect 695 1601 699 1602
rect 711 1606 715 1607
rect 711 1601 715 1602
rect 502 1600 508 1601
rect 502 1596 503 1600
rect 507 1596 508 1600
rect 502 1595 508 1596
rect 694 1600 700 1601
rect 694 1596 695 1600
rect 699 1596 700 1600
rect 694 1595 700 1596
rect 478 1579 484 1580
rect 110 1575 116 1576
rect 110 1571 111 1575
rect 115 1571 116 1575
rect 142 1575 148 1576
rect 110 1570 116 1571
rect 134 1571 140 1572
rect 112 1555 114 1570
rect 134 1567 135 1571
rect 139 1567 140 1571
rect 142 1571 143 1575
rect 147 1571 148 1575
rect 310 1575 316 1576
rect 142 1570 148 1571
rect 302 1571 308 1572
rect 134 1566 140 1567
rect 302 1567 303 1571
rect 307 1567 308 1571
rect 310 1571 311 1575
rect 315 1571 316 1575
rect 478 1575 479 1579
rect 483 1575 484 1579
rect 720 1576 722 1642
rect 918 1620 924 1621
rect 918 1616 919 1620
rect 923 1616 924 1620
rect 918 1615 924 1616
rect 920 1607 922 1615
rect 887 1606 891 1607
rect 887 1601 891 1602
rect 919 1606 923 1607
rect 919 1601 923 1602
rect 886 1600 892 1601
rect 886 1596 887 1600
rect 891 1596 892 1600
rect 886 1595 892 1596
rect 478 1574 484 1575
rect 718 1575 724 1576
rect 310 1570 316 1571
rect 502 1571 508 1572
rect 302 1566 308 1567
rect 502 1567 503 1571
rect 507 1567 508 1571
rect 502 1566 508 1567
rect 694 1571 700 1572
rect 694 1567 695 1571
rect 699 1567 700 1571
rect 718 1571 719 1575
rect 723 1571 724 1575
rect 928 1572 930 1642
rect 1063 1606 1067 1607
rect 1063 1601 1067 1602
rect 1062 1600 1068 1601
rect 1062 1596 1063 1600
rect 1067 1596 1068 1600
rect 1062 1595 1068 1596
rect 1072 1576 1074 1666
rect 1143 1654 1147 1655
rect 1142 1649 1148 1650
rect 1142 1645 1143 1649
rect 1147 1645 1148 1649
rect 1168 1648 1170 1742
rect 1670 1741 1676 1742
rect 1670 1737 1671 1741
rect 1675 1737 1676 1741
rect 1814 1741 1815 1745
rect 1819 1741 1820 1745
rect 1814 1740 1820 1741
rect 1966 1741 1967 1745
rect 1971 1741 1972 1745
rect 1966 1740 1972 1741
rect 2126 1741 2127 1745
rect 2131 1741 2132 1745
rect 2126 1740 2132 1741
rect 2302 1741 2303 1745
rect 2307 1741 2308 1745
rect 2302 1740 2308 1741
rect 2502 1741 2503 1745
rect 2507 1741 2508 1745
rect 2502 1740 2508 1741
rect 2710 1745 2716 1746
rect 2710 1741 2711 1745
rect 2715 1741 2716 1745
rect 2710 1740 2716 1741
rect 2934 1745 2940 1746
rect 2943 1745 2947 1746
rect 2934 1741 2935 1745
rect 2939 1741 2940 1745
rect 2934 1740 2940 1741
rect 1670 1736 1676 1737
rect 1822 1739 1828 1740
rect 1822 1735 1823 1739
rect 1827 1735 1828 1739
rect 1822 1734 1828 1735
rect 2030 1739 2036 1740
rect 2030 1735 2031 1739
rect 2035 1735 2036 1739
rect 2030 1734 2036 1735
rect 2322 1739 2328 1740
rect 2322 1735 2323 1739
rect 2327 1735 2328 1739
rect 2322 1734 2328 1735
rect 2474 1739 2480 1740
rect 2474 1735 2475 1739
rect 2479 1735 2480 1739
rect 2474 1734 2480 1735
rect 2718 1739 2724 1740
rect 2718 1735 2719 1739
rect 2723 1735 2724 1739
rect 2718 1734 2724 1735
rect 2943 1739 2949 1740
rect 2943 1735 2944 1739
rect 2948 1738 2949 1739
rect 2952 1738 2954 1762
rect 3158 1759 3159 1763
rect 3163 1759 3164 1763
rect 3166 1763 3167 1767
rect 3171 1763 3172 1767
rect 3166 1762 3172 1763
rect 3190 1767 3196 1768
rect 3190 1763 3191 1767
rect 3195 1763 3196 1767
rect 3190 1762 3196 1763
rect 3158 1758 3164 1759
rect 3160 1751 3162 1758
rect 3159 1750 3163 1751
rect 3158 1745 3164 1746
rect 3158 1741 3159 1745
rect 3163 1741 3164 1745
rect 3168 1744 3170 1762
rect 3192 1751 3194 1762
rect 3191 1750 3195 1751
rect 3191 1745 3195 1746
rect 3158 1740 3164 1741
rect 3166 1743 3172 1744
rect 3166 1739 3167 1743
rect 3171 1739 3172 1743
rect 3192 1742 3194 1745
rect 3166 1738 3172 1739
rect 3190 1741 3196 1742
rect 2948 1736 2954 1738
rect 2948 1735 2949 1736
rect 2943 1734 2949 1735
rect 1630 1731 1636 1732
rect 1630 1727 1631 1731
rect 1635 1727 1636 1731
rect 1630 1726 1636 1727
rect 1632 1707 1634 1726
rect 1670 1723 1676 1724
rect 1670 1719 1671 1723
rect 1675 1719 1676 1723
rect 1670 1718 1676 1719
rect 1672 1711 1674 1718
rect 1814 1716 1820 1717
rect 1814 1712 1815 1716
rect 1819 1712 1820 1716
rect 1814 1711 1820 1712
rect 1671 1710 1675 1711
rect 1631 1706 1635 1707
rect 1671 1705 1675 1706
rect 1735 1710 1739 1711
rect 1735 1705 1739 1706
rect 1815 1710 1819 1711
rect 1815 1705 1819 1706
rect 1631 1701 1635 1702
rect 1632 1694 1634 1701
rect 1672 1698 1674 1705
rect 1734 1704 1740 1705
rect 1734 1700 1735 1704
rect 1739 1700 1740 1704
rect 1734 1699 1740 1700
rect 1670 1697 1676 1698
rect 1630 1693 1636 1694
rect 1630 1689 1631 1693
rect 1635 1689 1636 1693
rect 1670 1693 1671 1697
rect 1675 1693 1676 1697
rect 1670 1692 1676 1693
rect 1630 1688 1636 1689
rect 1824 1684 1826 1734
rect 1966 1716 1972 1717
rect 1966 1712 1967 1716
rect 1971 1712 1972 1716
rect 1966 1711 1972 1712
rect 1879 1710 1883 1711
rect 1879 1705 1883 1706
rect 1967 1710 1971 1711
rect 1967 1705 1971 1706
rect 2023 1710 2027 1711
rect 2023 1705 2027 1706
rect 1878 1704 1884 1705
rect 1878 1700 1879 1704
rect 1883 1700 1884 1704
rect 1878 1699 1884 1700
rect 2022 1704 2028 1705
rect 2022 1700 2023 1704
rect 2027 1700 2028 1704
rect 2022 1699 2028 1700
rect 1822 1683 1828 1684
rect 1670 1679 1676 1680
rect 1630 1675 1636 1676
rect 1630 1671 1631 1675
rect 1635 1671 1636 1675
rect 1670 1675 1671 1679
rect 1675 1675 1676 1679
rect 1822 1679 1823 1683
rect 1827 1679 1828 1683
rect 2032 1680 2034 1734
rect 2126 1716 2132 1717
rect 2126 1712 2127 1716
rect 2131 1712 2132 1716
rect 2126 1711 2132 1712
rect 2302 1716 2308 1717
rect 2302 1712 2303 1716
rect 2307 1712 2308 1716
rect 2302 1711 2308 1712
rect 2127 1710 2131 1711
rect 2127 1705 2131 1706
rect 2167 1710 2171 1711
rect 2167 1705 2171 1706
rect 2303 1710 2307 1711
rect 2303 1705 2307 1706
rect 2311 1710 2315 1711
rect 2311 1705 2315 1706
rect 2166 1704 2172 1705
rect 2166 1700 2167 1704
rect 2171 1700 2172 1704
rect 2166 1699 2172 1700
rect 2310 1704 2316 1705
rect 2310 1700 2311 1704
rect 2315 1700 2316 1704
rect 2310 1699 2316 1700
rect 2324 1680 2326 1734
rect 2463 1710 2467 1711
rect 2463 1705 2467 1706
rect 2462 1704 2468 1705
rect 2462 1700 2463 1704
rect 2467 1700 2468 1704
rect 2462 1699 2468 1700
rect 2476 1680 2478 1734
rect 2502 1716 2508 1717
rect 2502 1712 2503 1716
rect 2507 1712 2508 1716
rect 2502 1711 2508 1712
rect 2710 1716 2716 1717
rect 2710 1712 2711 1716
rect 2715 1712 2716 1716
rect 2710 1711 2716 1712
rect 2503 1710 2507 1711
rect 2503 1705 2507 1706
rect 2711 1710 2715 1711
rect 2711 1705 2715 1706
rect 1822 1678 1828 1679
rect 2030 1679 2036 1680
rect 1824 1676 1826 1678
rect 1670 1674 1676 1675
rect 1734 1675 1740 1676
rect 1672 1671 1674 1674
rect 1734 1671 1735 1675
rect 1739 1671 1740 1675
rect 1630 1670 1636 1671
rect 1671 1670 1675 1671
rect 1632 1655 1634 1670
rect 1695 1670 1699 1671
rect 1734 1670 1740 1671
rect 1822 1675 1828 1676
rect 1822 1671 1823 1675
rect 1827 1671 1828 1675
rect 1822 1670 1828 1671
rect 1878 1675 1884 1676
rect 1878 1671 1879 1675
rect 1883 1671 1884 1675
rect 2022 1675 2028 1676
rect 2022 1671 2023 1675
rect 2027 1671 2028 1675
rect 2030 1675 2031 1679
rect 2035 1675 2036 1679
rect 2030 1674 2036 1675
rect 2106 1679 2112 1680
rect 2106 1675 2107 1679
rect 2111 1675 2112 1679
rect 2322 1679 2328 1680
rect 2106 1674 2112 1675
rect 2166 1675 2172 1676
rect 1878 1670 1884 1671
rect 1895 1670 1899 1671
rect 2022 1670 2028 1671
rect 1671 1665 1675 1666
rect 1694 1665 1700 1666
rect 1735 1665 1739 1666
rect 1879 1665 1883 1666
rect 1894 1665 1900 1666
rect 2023 1665 2027 1666
rect 1672 1662 1674 1665
rect 1670 1661 1676 1662
rect 1670 1657 1671 1661
rect 1675 1657 1676 1661
rect 1694 1661 1695 1665
rect 1699 1661 1700 1665
rect 1694 1660 1700 1661
rect 1894 1661 1895 1665
rect 1899 1661 1900 1665
rect 1894 1660 1900 1661
rect 2108 1660 2110 1674
rect 2166 1671 2167 1675
rect 2171 1671 2172 1675
rect 2127 1670 2131 1671
rect 2166 1670 2172 1671
rect 2310 1675 2316 1676
rect 2310 1671 2311 1675
rect 2315 1671 2316 1675
rect 2322 1675 2323 1679
rect 2327 1675 2328 1679
rect 2474 1679 2480 1680
rect 2322 1674 2328 1675
rect 2462 1675 2468 1676
rect 2310 1670 2316 1671
rect 2126 1665 2132 1666
rect 2167 1665 2171 1666
rect 2311 1665 2315 1666
rect 2126 1661 2127 1665
rect 2131 1661 2132 1665
rect 2126 1660 2132 1661
rect 2324 1660 2326 1674
rect 2462 1671 2463 1675
rect 2467 1671 2468 1675
rect 2474 1675 2475 1679
rect 2479 1675 2480 1679
rect 2474 1674 2480 1675
rect 2367 1670 2371 1671
rect 2462 1670 2468 1671
rect 2615 1670 2619 1671
rect 2366 1665 2372 1666
rect 2463 1665 2467 1666
rect 2614 1665 2620 1666
rect 2366 1661 2367 1665
rect 2371 1661 2372 1665
rect 2366 1660 2372 1661
rect 2614 1661 2615 1665
rect 2619 1661 2620 1665
rect 2614 1660 2620 1661
rect 2720 1660 2722 1734
rect 2934 1716 2940 1717
rect 2934 1712 2935 1716
rect 2939 1712 2940 1716
rect 2934 1711 2940 1712
rect 3158 1716 3164 1717
rect 3158 1712 3159 1716
rect 3163 1712 3164 1716
rect 3158 1711 3164 1712
rect 2935 1710 2939 1711
rect 2935 1705 2939 1706
rect 3159 1710 3163 1711
rect 3159 1705 3163 1706
rect 2871 1670 2875 1671
rect 3135 1670 3139 1671
rect 2870 1665 2876 1666
rect 2870 1661 2871 1665
rect 2875 1661 2876 1665
rect 2870 1660 2876 1661
rect 3134 1665 3140 1666
rect 3134 1661 3135 1665
rect 3139 1661 3140 1665
rect 3168 1664 3170 1738
rect 3190 1737 3191 1741
rect 3195 1737 3196 1741
rect 3190 1736 3196 1737
rect 3190 1723 3196 1724
rect 3190 1719 3191 1723
rect 3195 1719 3196 1723
rect 3190 1718 3196 1719
rect 3192 1711 3194 1718
rect 3191 1710 3195 1711
rect 3191 1705 3195 1706
rect 3192 1698 3194 1705
rect 3190 1697 3196 1698
rect 3190 1693 3191 1697
rect 3195 1693 3196 1697
rect 3190 1692 3196 1693
rect 3190 1679 3196 1680
rect 3190 1675 3191 1679
rect 3195 1675 3196 1679
rect 3190 1674 3196 1675
rect 3192 1671 3194 1674
rect 3191 1670 3195 1671
rect 3191 1665 3195 1666
rect 3134 1660 3140 1661
rect 3142 1663 3148 1664
rect 1670 1656 1676 1657
rect 2106 1659 2112 1660
rect 2106 1655 2107 1659
rect 2111 1655 2112 1659
rect 1383 1654 1387 1655
rect 1599 1654 1603 1655
rect 1631 1654 1635 1655
rect 2106 1654 2112 1655
rect 2322 1659 2328 1660
rect 2322 1655 2323 1659
rect 2327 1655 2328 1659
rect 2322 1654 2328 1655
rect 2398 1659 2404 1660
rect 2398 1655 2399 1659
rect 2403 1655 2404 1659
rect 2398 1654 2404 1655
rect 2718 1659 2724 1660
rect 2718 1655 2719 1659
rect 2723 1655 2724 1659
rect 2718 1654 2724 1655
rect 2918 1659 2924 1660
rect 2918 1655 2919 1659
rect 2923 1655 2924 1659
rect 3142 1659 3143 1663
rect 3147 1659 3148 1663
rect 3142 1658 3148 1659
rect 3166 1663 3172 1664
rect 3166 1659 3167 1663
rect 3171 1659 3172 1663
rect 3192 1662 3194 1665
rect 3166 1658 3172 1659
rect 3190 1661 3196 1662
rect 2918 1654 2924 1655
rect 1382 1649 1388 1650
rect 1142 1644 1148 1645
rect 1166 1647 1172 1648
rect 1166 1643 1167 1647
rect 1171 1643 1172 1647
rect 1382 1645 1383 1649
rect 1387 1645 1388 1649
rect 1382 1644 1388 1645
rect 1598 1649 1604 1650
rect 1631 1649 1635 1650
rect 1598 1645 1599 1649
rect 1603 1645 1604 1649
rect 1598 1644 1604 1645
rect 1606 1647 1612 1648
rect 1166 1642 1172 1643
rect 1422 1643 1428 1644
rect 1142 1620 1148 1621
rect 1142 1616 1143 1620
rect 1147 1616 1148 1620
rect 1142 1615 1148 1616
rect 1144 1607 1146 1615
rect 1143 1606 1147 1607
rect 1143 1601 1147 1602
rect 1168 1580 1170 1642
rect 1422 1639 1423 1643
rect 1427 1639 1428 1643
rect 1606 1643 1607 1647
rect 1611 1643 1612 1647
rect 1632 1646 1634 1649
rect 1606 1642 1612 1643
rect 1630 1645 1636 1646
rect 1422 1638 1428 1639
rect 1382 1620 1388 1621
rect 1382 1616 1383 1620
rect 1387 1616 1388 1620
rect 1382 1615 1388 1616
rect 1384 1607 1386 1615
rect 1239 1606 1243 1607
rect 1239 1601 1243 1602
rect 1383 1606 1387 1607
rect 1383 1601 1387 1602
rect 1415 1606 1419 1607
rect 1415 1601 1419 1602
rect 1238 1600 1244 1601
rect 1238 1596 1239 1600
rect 1243 1596 1244 1600
rect 1238 1595 1244 1596
rect 1414 1600 1420 1601
rect 1414 1596 1415 1600
rect 1419 1596 1420 1600
rect 1414 1595 1420 1596
rect 1166 1579 1172 1580
rect 1070 1575 1076 1576
rect 718 1570 724 1571
rect 886 1571 892 1572
rect 694 1566 700 1567
rect 136 1555 138 1566
rect 304 1555 306 1566
rect 504 1555 506 1566
rect 696 1555 698 1566
rect 111 1554 115 1555
rect 111 1549 115 1550
rect 135 1554 139 1555
rect 135 1549 139 1550
rect 303 1554 307 1555
rect 303 1549 307 1550
rect 503 1554 507 1555
rect 679 1554 683 1555
rect 695 1554 699 1555
rect 503 1549 507 1550
rect 678 1549 684 1550
rect 695 1549 699 1550
rect 112 1546 114 1549
rect 110 1545 116 1546
rect 110 1541 111 1545
rect 115 1541 116 1545
rect 678 1545 679 1549
rect 683 1545 684 1549
rect 720 1548 722 1570
rect 886 1567 887 1571
rect 891 1567 892 1571
rect 886 1566 892 1567
rect 894 1571 900 1572
rect 894 1567 895 1571
rect 899 1567 900 1571
rect 894 1566 900 1567
rect 926 1571 932 1572
rect 926 1567 927 1571
rect 931 1567 932 1571
rect 926 1566 932 1567
rect 1062 1571 1068 1572
rect 1062 1567 1063 1571
rect 1067 1567 1068 1571
rect 1070 1571 1071 1575
rect 1075 1571 1076 1575
rect 1166 1575 1167 1579
rect 1171 1575 1172 1579
rect 1166 1574 1172 1575
rect 1286 1575 1292 1576
rect 1070 1570 1076 1571
rect 1062 1566 1068 1567
rect 888 1555 890 1566
rect 807 1554 811 1555
rect 887 1554 891 1555
rect 806 1549 812 1550
rect 887 1549 891 1550
rect 678 1544 684 1545
rect 718 1547 724 1548
rect 718 1543 719 1547
rect 723 1543 724 1547
rect 806 1545 807 1549
rect 811 1545 812 1549
rect 806 1544 812 1545
rect 896 1544 898 1566
rect 1064 1555 1066 1566
rect 927 1554 931 1555
rect 1047 1554 1051 1555
rect 1063 1554 1067 1555
rect 926 1549 932 1550
rect 926 1545 927 1549
rect 931 1545 932 1549
rect 926 1544 932 1545
rect 1046 1549 1052 1550
rect 1063 1549 1067 1550
rect 1046 1545 1047 1549
rect 1051 1545 1052 1549
rect 1072 1548 1074 1570
rect 1168 1563 1170 1574
rect 1238 1571 1244 1572
rect 1238 1567 1239 1571
rect 1243 1567 1244 1571
rect 1286 1571 1287 1575
rect 1291 1571 1292 1575
rect 1424 1572 1426 1638
rect 1598 1620 1604 1621
rect 1598 1616 1599 1620
rect 1603 1616 1604 1620
rect 1598 1615 1604 1616
rect 1600 1607 1602 1615
rect 1591 1606 1595 1607
rect 1591 1601 1595 1602
rect 1599 1606 1603 1607
rect 1599 1601 1603 1602
rect 1590 1600 1596 1601
rect 1590 1596 1591 1600
rect 1595 1596 1596 1600
rect 1590 1595 1596 1596
rect 1286 1570 1292 1571
rect 1414 1571 1420 1572
rect 1238 1566 1244 1567
rect 1168 1561 1178 1563
rect 1167 1554 1171 1555
rect 1166 1549 1172 1550
rect 1046 1544 1052 1545
rect 1070 1547 1076 1548
rect 718 1542 724 1543
rect 838 1543 844 1544
rect 110 1540 116 1541
rect 838 1539 839 1543
rect 843 1539 844 1543
rect 838 1538 844 1539
rect 894 1543 900 1544
rect 894 1539 895 1543
rect 899 1539 900 1543
rect 1070 1543 1071 1547
rect 1075 1543 1076 1547
rect 1166 1545 1167 1549
rect 1171 1545 1172 1549
rect 1176 1548 1178 1561
rect 1240 1555 1242 1566
rect 1239 1554 1243 1555
rect 1279 1554 1283 1555
rect 1239 1549 1243 1550
rect 1278 1549 1284 1550
rect 1166 1544 1172 1545
rect 1174 1547 1180 1548
rect 1070 1542 1076 1543
rect 1174 1543 1175 1547
rect 1179 1543 1180 1547
rect 1174 1542 1180 1543
rect 1190 1547 1196 1548
rect 1190 1543 1191 1547
rect 1195 1543 1196 1547
rect 1278 1545 1279 1549
rect 1283 1545 1284 1549
rect 1288 1548 1290 1570
rect 1414 1567 1415 1571
rect 1419 1567 1420 1571
rect 1414 1566 1420 1567
rect 1422 1571 1428 1572
rect 1422 1567 1423 1571
rect 1427 1567 1428 1571
rect 1422 1566 1428 1567
rect 1590 1571 1596 1572
rect 1590 1567 1591 1571
rect 1595 1567 1596 1571
rect 1590 1566 1596 1567
rect 1599 1571 1605 1572
rect 1599 1567 1600 1571
rect 1604 1570 1605 1571
rect 1608 1570 1610 1642
rect 1630 1641 1631 1645
rect 1635 1641 1636 1645
rect 1630 1640 1636 1641
rect 1670 1643 1676 1644
rect 1670 1639 1671 1643
rect 1675 1639 1676 1643
rect 1670 1638 1676 1639
rect 1630 1627 1636 1628
rect 1672 1627 1674 1638
rect 1694 1636 1700 1637
rect 1694 1632 1695 1636
rect 1699 1632 1700 1636
rect 1694 1631 1700 1632
rect 1894 1636 1900 1637
rect 1894 1632 1895 1636
rect 1899 1632 1900 1636
rect 1894 1631 1900 1632
rect 1696 1627 1698 1631
rect 1896 1627 1898 1631
rect 1630 1623 1631 1627
rect 1635 1623 1636 1627
rect 1630 1622 1636 1623
rect 1671 1626 1675 1627
rect 1632 1607 1634 1622
rect 1671 1621 1675 1622
rect 1695 1626 1699 1627
rect 1695 1621 1699 1622
rect 1895 1626 1899 1627
rect 1895 1621 1899 1622
rect 1672 1614 1674 1621
rect 1670 1613 1676 1614
rect 1670 1609 1671 1613
rect 1675 1609 1676 1613
rect 1670 1608 1676 1609
rect 1631 1606 1635 1607
rect 1631 1601 1635 1602
rect 1632 1594 1634 1601
rect 1670 1595 1676 1596
rect 1630 1593 1636 1594
rect 1630 1589 1631 1593
rect 1635 1589 1636 1593
rect 1670 1591 1671 1595
rect 1675 1591 1676 1595
rect 1670 1590 1676 1591
rect 1630 1588 1636 1589
rect 1672 1587 1674 1590
rect 1671 1586 1675 1587
rect 1671 1581 1675 1582
rect 1672 1578 1674 1581
rect 1670 1577 1676 1578
rect 1630 1575 1636 1576
rect 1630 1571 1631 1575
rect 1635 1571 1636 1575
rect 1670 1573 1671 1577
rect 1675 1573 1676 1577
rect 1670 1572 1676 1573
rect 1630 1570 1636 1571
rect 1604 1568 1610 1570
rect 1604 1567 1605 1568
rect 1599 1566 1605 1567
rect 1416 1555 1418 1566
rect 1399 1554 1403 1555
rect 1415 1554 1419 1555
rect 1398 1549 1404 1550
rect 1415 1549 1419 1550
rect 1278 1544 1284 1545
rect 1286 1547 1292 1548
rect 1190 1542 1196 1543
rect 1286 1543 1287 1547
rect 1291 1543 1292 1547
rect 1398 1545 1399 1549
rect 1403 1545 1404 1549
rect 1398 1544 1404 1545
rect 1424 1544 1426 1566
rect 1592 1555 1594 1566
rect 1519 1554 1523 1555
rect 1591 1554 1595 1555
rect 1518 1549 1524 1550
rect 1591 1549 1595 1550
rect 1518 1545 1519 1549
rect 1523 1545 1524 1549
rect 1518 1544 1524 1545
rect 1600 1544 1602 1566
rect 1632 1555 1634 1570
rect 1670 1559 1676 1560
rect 1670 1555 1671 1559
rect 1675 1555 1676 1559
rect 1631 1554 1635 1555
rect 1670 1554 1676 1555
rect 1631 1549 1635 1550
rect 1632 1546 1634 1549
rect 1630 1545 1636 1546
rect 1286 1542 1292 1543
rect 1406 1543 1412 1544
rect 894 1538 900 1539
rect 110 1527 116 1528
rect 110 1523 111 1527
rect 115 1523 116 1527
rect 110 1522 116 1523
rect 112 1507 114 1522
rect 678 1520 684 1521
rect 678 1516 679 1520
rect 683 1516 684 1520
rect 678 1515 684 1516
rect 806 1520 812 1521
rect 806 1516 807 1520
rect 811 1516 812 1520
rect 806 1515 812 1516
rect 680 1507 682 1515
rect 808 1507 810 1515
rect 111 1506 115 1507
rect 111 1501 115 1502
rect 575 1506 579 1507
rect 575 1501 579 1502
rect 679 1506 683 1507
rect 679 1501 683 1502
rect 703 1506 707 1507
rect 703 1501 707 1502
rect 807 1506 811 1507
rect 807 1501 811 1502
rect 831 1506 835 1507
rect 831 1501 835 1502
rect 112 1494 114 1501
rect 574 1500 580 1501
rect 574 1496 575 1500
rect 579 1496 580 1500
rect 574 1495 580 1496
rect 702 1500 708 1501
rect 702 1496 703 1500
rect 707 1496 708 1500
rect 702 1495 708 1496
rect 830 1500 836 1501
rect 830 1496 831 1500
rect 835 1496 836 1500
rect 830 1495 836 1496
rect 110 1493 116 1494
rect 110 1489 111 1493
rect 115 1489 116 1493
rect 110 1488 116 1489
rect 110 1475 116 1476
rect 110 1471 111 1475
rect 115 1471 116 1475
rect 840 1472 842 1538
rect 926 1520 932 1521
rect 926 1516 927 1520
rect 931 1516 932 1520
rect 926 1515 932 1516
rect 1046 1520 1052 1521
rect 1046 1516 1047 1520
rect 1051 1516 1052 1520
rect 1046 1515 1052 1516
rect 1166 1520 1172 1521
rect 1166 1516 1167 1520
rect 1171 1516 1172 1520
rect 1166 1515 1172 1516
rect 928 1507 930 1515
rect 1048 1507 1050 1515
rect 1168 1507 1170 1515
rect 927 1506 931 1507
rect 927 1501 931 1502
rect 951 1506 955 1507
rect 951 1501 955 1502
rect 1047 1506 1051 1507
rect 1047 1501 1051 1502
rect 1071 1506 1075 1507
rect 1071 1501 1075 1502
rect 1167 1506 1171 1507
rect 1167 1501 1171 1502
rect 1183 1506 1187 1507
rect 1183 1501 1187 1502
rect 950 1500 956 1501
rect 950 1496 951 1500
rect 955 1496 956 1500
rect 950 1495 956 1496
rect 1070 1500 1076 1501
rect 1070 1496 1071 1500
rect 1075 1496 1076 1500
rect 1070 1495 1076 1496
rect 1182 1500 1188 1501
rect 1182 1496 1183 1500
rect 1187 1496 1188 1500
rect 1182 1495 1188 1496
rect 1192 1472 1194 1542
rect 1278 1520 1284 1521
rect 1278 1516 1279 1520
rect 1283 1516 1284 1520
rect 1278 1515 1284 1516
rect 1280 1507 1282 1515
rect 1279 1506 1283 1507
rect 1279 1501 1283 1502
rect 1288 1480 1290 1542
rect 1406 1539 1407 1543
rect 1411 1539 1412 1543
rect 1406 1538 1412 1539
rect 1422 1543 1428 1544
rect 1422 1539 1423 1543
rect 1427 1539 1428 1543
rect 1422 1538 1428 1539
rect 1598 1543 1604 1544
rect 1598 1539 1599 1543
rect 1603 1539 1604 1543
rect 1630 1541 1631 1545
rect 1635 1541 1636 1545
rect 1630 1540 1636 1541
rect 1672 1539 1674 1554
rect 1598 1538 1604 1539
rect 1671 1538 1675 1539
rect 1398 1520 1404 1521
rect 1398 1516 1399 1520
rect 1403 1516 1404 1520
rect 1398 1515 1404 1516
rect 1400 1507 1402 1515
rect 1295 1506 1299 1507
rect 1295 1501 1299 1502
rect 1399 1506 1403 1507
rect 1399 1501 1403 1502
rect 1294 1500 1300 1501
rect 1294 1496 1295 1500
rect 1299 1496 1300 1500
rect 1294 1495 1300 1496
rect 1408 1480 1410 1538
rect 1671 1533 1675 1534
rect 1630 1527 1636 1528
rect 1630 1523 1631 1527
rect 1635 1523 1636 1527
rect 1672 1526 1674 1533
rect 1630 1522 1636 1523
rect 1670 1525 1676 1526
rect 1518 1520 1524 1521
rect 1518 1516 1519 1520
rect 1523 1516 1524 1520
rect 1518 1515 1524 1516
rect 1520 1507 1522 1515
rect 1632 1507 1634 1522
rect 1670 1521 1671 1525
rect 1675 1521 1676 1525
rect 1670 1520 1676 1521
rect 1670 1507 1676 1508
rect 1415 1506 1419 1507
rect 1415 1501 1419 1502
rect 1519 1506 1523 1507
rect 1519 1501 1523 1502
rect 1631 1506 1635 1507
rect 1670 1503 1671 1507
rect 1675 1503 1676 1507
rect 1670 1502 1676 1503
rect 1631 1501 1635 1502
rect 1414 1500 1420 1501
rect 1414 1496 1415 1500
rect 1419 1496 1420 1500
rect 1414 1495 1420 1496
rect 1632 1494 1634 1501
rect 1672 1495 1674 1502
rect 2108 1496 2110 1654
rect 2126 1636 2132 1637
rect 2126 1632 2127 1636
rect 2131 1632 2132 1636
rect 2126 1631 2132 1632
rect 2366 1636 2372 1637
rect 2366 1632 2367 1636
rect 2371 1632 2372 1636
rect 2366 1631 2372 1632
rect 2128 1627 2130 1631
rect 2368 1627 2370 1631
rect 2127 1626 2131 1627
rect 2127 1621 2131 1622
rect 2319 1626 2323 1627
rect 2319 1621 2323 1622
rect 2367 1626 2371 1627
rect 2367 1621 2371 1622
rect 2318 1620 2324 1621
rect 2318 1616 2319 1620
rect 2323 1616 2324 1620
rect 2318 1615 2324 1616
rect 2318 1591 2324 1592
rect 2318 1587 2319 1591
rect 2323 1587 2324 1591
rect 2271 1586 2275 1587
rect 2318 1586 2324 1587
rect 2290 1583 2296 1584
rect 2270 1581 2276 1582
rect 2270 1577 2271 1581
rect 2275 1577 2276 1581
rect 2290 1579 2291 1583
rect 2295 1579 2296 1583
rect 2319 1581 2323 1582
rect 2290 1578 2296 1579
rect 2270 1576 2276 1577
rect 2270 1552 2276 1553
rect 2270 1548 2271 1552
rect 2275 1548 2276 1552
rect 2270 1547 2276 1548
rect 2272 1539 2274 1547
rect 2167 1538 2171 1539
rect 2167 1533 2171 1534
rect 2271 1538 2275 1539
rect 2271 1533 2275 1534
rect 2279 1538 2283 1539
rect 2279 1533 2283 1534
rect 2166 1532 2172 1533
rect 2166 1528 2167 1532
rect 2171 1528 2172 1532
rect 2166 1527 2172 1528
rect 2278 1532 2284 1533
rect 2278 1528 2279 1532
rect 2283 1528 2284 1532
rect 2278 1527 2284 1528
rect 2292 1508 2294 1578
rect 2400 1576 2402 1654
rect 2614 1636 2620 1637
rect 2614 1632 2615 1636
rect 2619 1632 2620 1636
rect 2614 1631 2620 1632
rect 2616 1627 2618 1631
rect 2519 1626 2523 1627
rect 2519 1621 2523 1622
rect 2615 1626 2619 1627
rect 2615 1621 2619 1622
rect 2711 1626 2715 1627
rect 2711 1621 2715 1622
rect 2518 1620 2524 1621
rect 2518 1616 2519 1620
rect 2523 1616 2524 1620
rect 2518 1615 2524 1616
rect 2710 1620 2716 1621
rect 2710 1616 2711 1620
rect 2715 1616 2716 1620
rect 2710 1615 2716 1616
rect 2720 1592 2722 1654
rect 2870 1636 2876 1637
rect 2870 1632 2871 1636
rect 2875 1632 2876 1636
rect 2870 1631 2876 1632
rect 2872 1627 2874 1631
rect 2871 1626 2875 1627
rect 2871 1621 2875 1622
rect 2911 1626 2915 1627
rect 2911 1621 2915 1622
rect 2910 1620 2916 1621
rect 2910 1616 2911 1620
rect 2915 1616 2916 1620
rect 2910 1615 2916 1616
rect 2920 1592 2922 1654
rect 3134 1636 3140 1637
rect 3134 1632 3135 1636
rect 3139 1632 3140 1636
rect 3134 1631 3140 1632
rect 3136 1627 3138 1631
rect 3111 1626 3115 1627
rect 3111 1621 3115 1622
rect 3135 1626 3139 1627
rect 3135 1621 3139 1622
rect 3110 1620 3116 1621
rect 3110 1616 3111 1620
rect 3115 1616 3116 1620
rect 3110 1615 3116 1616
rect 3144 1596 3146 1658
rect 3190 1657 3191 1661
rect 3195 1657 3196 1661
rect 3190 1656 3196 1657
rect 3190 1643 3196 1644
rect 3190 1639 3191 1643
rect 3195 1639 3196 1643
rect 3190 1638 3196 1639
rect 3192 1627 3194 1638
rect 3191 1626 3195 1627
rect 3191 1621 3195 1622
rect 3192 1614 3194 1621
rect 3190 1613 3196 1614
rect 3190 1609 3191 1613
rect 3195 1609 3196 1613
rect 3190 1608 3196 1609
rect 3118 1595 3124 1596
rect 2518 1591 2524 1592
rect 2518 1587 2519 1591
rect 2523 1587 2524 1591
rect 2415 1586 2419 1587
rect 2518 1586 2524 1587
rect 2526 1591 2532 1592
rect 2526 1587 2527 1591
rect 2531 1587 2532 1591
rect 2710 1591 2716 1592
rect 2710 1587 2711 1591
rect 2715 1587 2716 1591
rect 2526 1586 2532 1587
rect 2559 1586 2563 1587
rect 2414 1581 2420 1582
rect 2519 1581 2523 1582
rect 2414 1577 2415 1581
rect 2419 1577 2420 1581
rect 2414 1576 2420 1577
rect 2528 1576 2530 1586
rect 2695 1586 2699 1587
rect 2710 1586 2716 1587
rect 2718 1591 2724 1592
rect 2718 1587 2719 1591
rect 2723 1587 2724 1591
rect 2910 1591 2916 1592
rect 2910 1587 2911 1591
rect 2915 1587 2916 1591
rect 2718 1586 2724 1587
rect 2839 1586 2843 1587
rect 2910 1586 2916 1587
rect 2918 1591 2924 1592
rect 2918 1587 2919 1591
rect 2923 1587 2924 1591
rect 3006 1591 3012 1592
rect 3006 1587 3007 1591
rect 3011 1587 3012 1591
rect 2918 1586 2924 1587
rect 2983 1586 2987 1587
rect 3006 1586 3012 1587
rect 3110 1591 3116 1592
rect 3110 1587 3111 1591
rect 3115 1587 3116 1591
rect 3118 1591 3119 1595
rect 3123 1591 3124 1595
rect 3118 1590 3124 1591
rect 3142 1595 3148 1596
rect 3142 1591 3143 1595
rect 3147 1591 3148 1595
rect 3142 1590 3148 1591
rect 3190 1595 3196 1596
rect 3190 1591 3191 1595
rect 3195 1591 3196 1595
rect 3190 1590 3196 1591
rect 3110 1586 3116 1587
rect 2558 1581 2564 1582
rect 2558 1577 2559 1581
rect 2563 1577 2564 1581
rect 2558 1576 2564 1577
rect 2694 1581 2700 1582
rect 2711 1581 2715 1582
rect 2694 1577 2695 1581
rect 2699 1577 2700 1581
rect 2694 1576 2700 1577
rect 2720 1576 2722 1586
rect 2838 1581 2844 1582
rect 2911 1581 2915 1582
rect 2838 1577 2839 1581
rect 2843 1577 2844 1581
rect 2838 1576 2844 1577
rect 2920 1576 2922 1586
rect 2982 1581 2988 1582
rect 2982 1577 2983 1581
rect 2987 1577 2988 1581
rect 2982 1576 2988 1577
rect 3008 1576 3010 1586
rect 3111 1581 3115 1582
rect 2398 1575 2404 1576
rect 2398 1571 2399 1575
rect 2403 1571 2404 1575
rect 2398 1570 2404 1571
rect 2526 1575 2532 1576
rect 2526 1571 2527 1575
rect 2531 1571 2532 1575
rect 2526 1570 2532 1571
rect 2662 1575 2668 1576
rect 2662 1571 2663 1575
rect 2667 1571 2668 1575
rect 2662 1570 2668 1571
rect 2718 1575 2724 1576
rect 2718 1571 2719 1575
rect 2723 1571 2724 1575
rect 2718 1570 2724 1571
rect 2918 1575 2924 1576
rect 2918 1571 2919 1575
rect 2923 1571 2924 1575
rect 2918 1570 2924 1571
rect 3006 1575 3012 1576
rect 3006 1571 3007 1575
rect 3011 1571 3012 1575
rect 3006 1570 3012 1571
rect 2391 1538 2395 1539
rect 2391 1533 2395 1534
rect 2390 1532 2396 1533
rect 2390 1528 2391 1532
rect 2395 1528 2396 1532
rect 2390 1527 2396 1528
rect 2400 1508 2402 1570
rect 2414 1552 2420 1553
rect 2414 1548 2415 1552
rect 2419 1548 2420 1552
rect 2414 1547 2420 1548
rect 2416 1539 2418 1547
rect 2415 1538 2419 1539
rect 2415 1533 2419 1534
rect 2503 1538 2507 1539
rect 2503 1533 2507 1534
rect 2502 1532 2508 1533
rect 2502 1528 2503 1532
rect 2507 1528 2508 1532
rect 2502 1527 2508 1528
rect 2528 1512 2530 1570
rect 2558 1552 2564 1553
rect 2558 1548 2559 1552
rect 2563 1548 2564 1552
rect 2558 1547 2564 1548
rect 2560 1539 2562 1547
rect 2559 1538 2563 1539
rect 2559 1533 2563 1534
rect 2615 1538 2619 1539
rect 2615 1533 2619 1534
rect 2614 1532 2620 1533
rect 2614 1528 2615 1532
rect 2619 1528 2620 1532
rect 2614 1527 2620 1528
rect 2526 1511 2532 1512
rect 2290 1507 2296 1508
rect 2166 1503 2172 1504
rect 2166 1499 2167 1503
rect 2171 1499 2172 1503
rect 2166 1498 2172 1499
rect 2278 1503 2284 1504
rect 2278 1499 2279 1503
rect 2283 1499 2284 1503
rect 2290 1503 2291 1507
rect 2295 1503 2296 1507
rect 2398 1507 2404 1508
rect 2290 1502 2296 1503
rect 2390 1503 2396 1504
rect 2278 1498 2284 1499
rect 2106 1495 2112 1496
rect 2168 1495 2170 1498
rect 2280 1495 2282 1498
rect 1671 1494 1675 1495
rect 1630 1493 1636 1494
rect 1630 1489 1631 1493
rect 1635 1489 1636 1493
rect 2087 1494 2091 1495
rect 2106 1491 2107 1495
rect 2111 1491 2112 1495
rect 2106 1490 2112 1491
rect 2167 1494 2171 1495
rect 2231 1494 2235 1495
rect 2279 1494 2283 1495
rect 1671 1489 1675 1490
rect 2086 1489 2092 1490
rect 1630 1488 1636 1489
rect 1672 1486 1674 1489
rect 1670 1485 1676 1486
rect 1670 1481 1671 1485
rect 1675 1481 1676 1485
rect 2086 1485 2087 1489
rect 2091 1485 2092 1489
rect 2086 1484 2092 1485
rect 2108 1484 2110 1490
rect 2167 1489 2171 1490
rect 2230 1489 2236 1490
rect 2279 1489 2283 1490
rect 2230 1485 2231 1489
rect 2235 1485 2236 1489
rect 2292 1488 2294 1502
rect 2390 1499 2391 1503
rect 2395 1499 2396 1503
rect 2398 1503 2399 1507
rect 2403 1503 2404 1507
rect 2526 1507 2527 1511
rect 2531 1507 2532 1511
rect 2664 1508 2666 1570
rect 2694 1552 2700 1553
rect 2694 1548 2695 1552
rect 2699 1548 2700 1552
rect 2694 1547 2700 1548
rect 2838 1552 2844 1553
rect 2838 1548 2839 1552
rect 2843 1548 2844 1552
rect 2838 1547 2844 1548
rect 2696 1539 2698 1547
rect 2840 1539 2842 1547
rect 2695 1538 2699 1539
rect 2695 1533 2699 1534
rect 2735 1538 2739 1539
rect 2735 1533 2739 1534
rect 2839 1538 2843 1539
rect 2839 1533 2843 1534
rect 2855 1538 2859 1539
rect 2855 1533 2859 1534
rect 2734 1532 2740 1533
rect 2734 1528 2735 1532
rect 2739 1528 2740 1532
rect 2734 1527 2740 1528
rect 2854 1532 2860 1533
rect 2854 1528 2855 1532
rect 2859 1528 2860 1532
rect 2854 1527 2860 1528
rect 2920 1508 2922 1570
rect 2982 1552 2988 1553
rect 2982 1548 2983 1552
rect 2987 1548 2988 1552
rect 2982 1547 2988 1548
rect 2984 1539 2986 1547
rect 2983 1538 2987 1539
rect 2983 1533 2987 1534
rect 2982 1532 2988 1533
rect 2982 1528 2983 1532
rect 2987 1528 2988 1532
rect 2982 1527 2988 1528
rect 2526 1506 2532 1507
rect 2662 1507 2668 1508
rect 2528 1504 2530 1506
rect 2398 1502 2404 1503
rect 2502 1503 2508 1504
rect 2390 1498 2396 1499
rect 2392 1495 2394 1498
rect 2400 1496 2402 1502
rect 2502 1499 2503 1503
rect 2507 1499 2508 1503
rect 2502 1498 2508 1499
rect 2526 1503 2532 1504
rect 2526 1499 2527 1503
rect 2531 1499 2532 1503
rect 2526 1498 2532 1499
rect 2614 1503 2620 1504
rect 2614 1499 2615 1503
rect 2619 1499 2620 1503
rect 2662 1503 2663 1507
rect 2667 1503 2668 1507
rect 2806 1507 2812 1508
rect 2662 1502 2668 1503
rect 2734 1503 2740 1504
rect 2614 1498 2620 1499
rect 2398 1495 2404 1496
rect 2375 1494 2379 1495
rect 2391 1494 2395 1495
rect 2398 1491 2399 1495
rect 2403 1491 2404 1495
rect 2398 1490 2404 1491
rect 2486 1495 2492 1496
rect 2504 1495 2506 1498
rect 2616 1495 2618 1498
rect 2486 1491 2487 1495
rect 2491 1491 2492 1495
rect 2486 1490 2492 1491
rect 2503 1494 2507 1495
rect 2511 1494 2515 1495
rect 2615 1494 2619 1495
rect 2655 1494 2659 1495
rect 2374 1489 2380 1490
rect 2391 1489 2395 1490
rect 2230 1484 2236 1485
rect 2238 1487 2244 1488
rect 1670 1480 1676 1481
rect 2106 1483 2112 1484
rect 1286 1479 1292 1480
rect 1286 1475 1287 1479
rect 1291 1475 1292 1479
rect 1406 1479 1412 1480
rect 1286 1474 1292 1475
rect 1318 1475 1324 1476
rect 110 1470 116 1471
rect 574 1471 580 1472
rect 112 1455 114 1470
rect 574 1467 575 1471
rect 579 1467 580 1471
rect 574 1466 580 1467
rect 586 1471 592 1472
rect 586 1467 587 1471
rect 591 1467 592 1471
rect 586 1466 592 1467
rect 702 1471 708 1472
rect 702 1467 703 1471
rect 707 1467 708 1471
rect 702 1466 708 1467
rect 734 1471 740 1472
rect 734 1467 735 1471
rect 739 1467 740 1471
rect 734 1466 740 1467
rect 830 1471 836 1472
rect 830 1467 831 1471
rect 835 1467 836 1471
rect 830 1466 836 1467
rect 838 1471 844 1472
rect 838 1467 839 1471
rect 843 1467 844 1471
rect 838 1466 844 1467
rect 950 1471 956 1472
rect 950 1467 951 1471
rect 955 1467 956 1471
rect 950 1466 956 1467
rect 958 1471 964 1472
rect 958 1467 959 1471
rect 963 1467 964 1471
rect 958 1466 964 1467
rect 1070 1471 1076 1472
rect 1070 1467 1071 1471
rect 1075 1467 1076 1471
rect 1070 1466 1076 1467
rect 1078 1471 1084 1472
rect 1078 1467 1079 1471
rect 1083 1467 1084 1471
rect 1182 1471 1188 1472
rect 1182 1467 1183 1471
rect 1187 1467 1188 1471
rect 1078 1466 1090 1467
rect 1182 1466 1188 1467
rect 1190 1471 1196 1472
rect 1190 1467 1191 1471
rect 1195 1467 1196 1471
rect 1294 1471 1300 1472
rect 1294 1467 1295 1471
rect 1299 1467 1300 1471
rect 1318 1471 1319 1475
rect 1323 1471 1324 1475
rect 1406 1475 1407 1479
rect 1411 1475 1412 1479
rect 2106 1479 2107 1483
rect 2111 1479 2112 1483
rect 2238 1483 2239 1487
rect 2243 1483 2244 1487
rect 2238 1482 2244 1483
rect 2290 1487 2296 1488
rect 2290 1483 2291 1487
rect 2295 1483 2296 1487
rect 2374 1485 2375 1489
rect 2379 1485 2380 1489
rect 2400 1488 2402 1490
rect 2374 1484 2380 1485
rect 2398 1487 2404 1488
rect 2290 1482 2296 1483
rect 2398 1483 2399 1487
rect 2403 1483 2404 1487
rect 2398 1482 2404 1483
rect 2106 1478 2112 1479
rect 1406 1474 1412 1475
rect 1630 1475 1636 1476
rect 1318 1470 1324 1471
rect 1414 1471 1420 1472
rect 1190 1466 1202 1467
rect 1294 1466 1300 1467
rect 576 1455 578 1466
rect 111 1454 115 1455
rect 479 1454 483 1455
rect 575 1454 579 1455
rect 111 1449 115 1450
rect 478 1449 484 1450
rect 575 1449 579 1450
rect 112 1446 114 1449
rect 110 1445 116 1446
rect 110 1441 111 1445
rect 115 1441 116 1445
rect 478 1445 479 1449
rect 483 1445 484 1449
rect 478 1444 484 1445
rect 588 1444 590 1466
rect 704 1455 706 1466
rect 607 1454 611 1455
rect 703 1454 707 1455
rect 727 1454 731 1455
rect 606 1449 612 1450
rect 703 1449 707 1450
rect 726 1449 732 1450
rect 606 1445 607 1449
rect 611 1445 612 1449
rect 606 1444 612 1445
rect 726 1445 727 1449
rect 731 1445 732 1449
rect 726 1444 732 1445
rect 736 1444 738 1466
rect 832 1455 834 1466
rect 831 1454 835 1455
rect 831 1449 835 1450
rect 840 1444 842 1466
rect 952 1455 954 1466
rect 847 1454 851 1455
rect 951 1454 955 1455
rect 846 1449 852 1450
rect 951 1449 955 1450
rect 846 1445 847 1449
rect 851 1445 852 1449
rect 846 1444 852 1445
rect 960 1444 962 1466
rect 1072 1455 1074 1466
rect 1080 1465 1090 1466
rect 967 1454 971 1455
rect 1071 1454 1075 1455
rect 1079 1454 1083 1455
rect 966 1449 972 1450
rect 1071 1449 1075 1450
rect 1078 1449 1084 1450
rect 966 1445 967 1449
rect 971 1445 972 1449
rect 966 1444 972 1445
rect 1078 1445 1079 1449
rect 1083 1445 1084 1449
rect 1078 1444 1084 1445
rect 1088 1444 1090 1465
rect 1184 1455 1186 1466
rect 1192 1465 1202 1466
rect 1183 1454 1187 1455
rect 1191 1454 1195 1455
rect 1183 1449 1187 1450
rect 1190 1449 1196 1450
rect 1190 1445 1191 1449
rect 1195 1445 1196 1449
rect 1200 1448 1202 1465
rect 1296 1455 1298 1466
rect 1295 1454 1299 1455
rect 1311 1454 1315 1455
rect 1295 1449 1299 1450
rect 1310 1449 1316 1450
rect 1190 1444 1196 1445
rect 1198 1447 1204 1448
rect 110 1440 116 1441
rect 586 1443 592 1444
rect 586 1439 587 1443
rect 591 1439 592 1443
rect 586 1438 592 1439
rect 634 1443 640 1444
rect 634 1439 635 1443
rect 639 1439 640 1443
rect 634 1438 640 1439
rect 734 1443 740 1444
rect 734 1439 735 1443
rect 739 1439 740 1443
rect 734 1438 740 1439
rect 838 1443 844 1444
rect 838 1439 839 1443
rect 843 1439 844 1443
rect 838 1438 844 1439
rect 886 1443 892 1444
rect 886 1439 887 1443
rect 891 1439 892 1443
rect 886 1438 892 1439
rect 958 1443 964 1444
rect 958 1439 959 1443
rect 963 1439 964 1443
rect 958 1438 964 1439
rect 1086 1443 1092 1444
rect 1086 1439 1087 1443
rect 1091 1439 1092 1443
rect 1086 1438 1092 1439
rect 1102 1443 1108 1444
rect 1102 1439 1103 1443
rect 1107 1439 1108 1443
rect 1198 1443 1199 1447
rect 1203 1443 1204 1447
rect 1310 1445 1311 1449
rect 1315 1445 1316 1449
rect 1320 1448 1322 1470
rect 1414 1467 1415 1471
rect 1419 1467 1420 1471
rect 1630 1471 1631 1475
rect 1635 1471 1636 1475
rect 1630 1470 1636 1471
rect 1414 1466 1420 1467
rect 1416 1455 1418 1466
rect 1632 1455 1634 1470
rect 1670 1467 1676 1468
rect 1670 1463 1671 1467
rect 1675 1463 1676 1467
rect 1670 1462 1676 1463
rect 1415 1454 1419 1455
rect 1415 1449 1419 1450
rect 1631 1454 1635 1455
rect 1672 1451 1674 1462
rect 2086 1460 2092 1461
rect 2086 1456 2087 1460
rect 2091 1456 2092 1460
rect 2086 1455 2092 1456
rect 2088 1451 2090 1455
rect 1631 1449 1635 1450
rect 1671 1450 1675 1451
rect 1310 1444 1316 1445
rect 1318 1447 1324 1448
rect 1198 1442 1204 1443
rect 1318 1443 1319 1447
rect 1323 1443 1324 1447
rect 1632 1446 1634 1449
rect 1318 1442 1324 1443
rect 1630 1445 1636 1446
rect 1671 1445 1675 1446
rect 1983 1450 1987 1451
rect 1983 1445 1987 1446
rect 2087 1450 2091 1451
rect 2087 1445 2091 1446
rect 2095 1450 2099 1451
rect 2095 1445 2099 1446
rect 1630 1441 1631 1445
rect 1635 1441 1636 1445
rect 1630 1440 1636 1441
rect 1102 1438 1108 1439
rect 1672 1438 1674 1445
rect 1982 1444 1988 1445
rect 1982 1440 1983 1444
rect 1987 1440 1988 1444
rect 1982 1439 1988 1440
rect 2094 1444 2100 1445
rect 2094 1440 2095 1444
rect 2099 1440 2100 1444
rect 2094 1439 2100 1440
rect 110 1427 116 1428
rect 110 1423 111 1427
rect 115 1423 116 1427
rect 110 1422 116 1423
rect 112 1403 114 1422
rect 478 1420 484 1421
rect 478 1416 479 1420
rect 483 1416 484 1420
rect 478 1415 484 1416
rect 606 1420 612 1421
rect 606 1416 607 1420
rect 611 1416 612 1420
rect 606 1415 612 1416
rect 480 1403 482 1415
rect 608 1403 610 1415
rect 111 1402 115 1403
rect 111 1397 115 1398
rect 375 1402 379 1403
rect 375 1397 379 1398
rect 479 1402 483 1403
rect 479 1397 483 1398
rect 503 1402 507 1403
rect 503 1397 507 1398
rect 607 1402 611 1403
rect 607 1397 611 1398
rect 623 1402 627 1403
rect 623 1397 627 1398
rect 112 1390 114 1397
rect 374 1396 380 1397
rect 374 1392 375 1396
rect 379 1392 380 1396
rect 374 1391 380 1392
rect 502 1396 508 1397
rect 502 1392 503 1396
rect 507 1392 508 1396
rect 502 1391 508 1392
rect 622 1396 628 1397
rect 622 1392 623 1396
rect 627 1392 628 1396
rect 622 1391 628 1392
rect 110 1389 116 1390
rect 110 1385 111 1389
rect 115 1385 116 1389
rect 110 1384 116 1385
rect 110 1371 116 1372
rect 110 1367 111 1371
rect 115 1367 116 1371
rect 636 1368 638 1438
rect 726 1420 732 1421
rect 726 1416 727 1420
rect 731 1416 732 1420
rect 726 1415 732 1416
rect 846 1420 852 1421
rect 846 1416 847 1420
rect 851 1416 852 1420
rect 846 1415 852 1416
rect 728 1403 730 1415
rect 848 1403 850 1415
rect 727 1402 731 1403
rect 727 1397 731 1398
rect 743 1402 747 1403
rect 743 1397 747 1398
rect 847 1402 851 1403
rect 847 1397 851 1398
rect 863 1402 867 1403
rect 863 1397 867 1398
rect 742 1396 748 1397
rect 742 1392 743 1396
rect 747 1392 748 1396
rect 742 1391 748 1392
rect 862 1396 868 1397
rect 862 1392 863 1396
rect 867 1392 868 1396
rect 862 1391 868 1392
rect 888 1368 890 1438
rect 966 1420 972 1421
rect 966 1416 967 1420
rect 971 1416 972 1420
rect 966 1415 972 1416
rect 1078 1420 1084 1421
rect 1078 1416 1079 1420
rect 1083 1416 1084 1420
rect 1078 1415 1084 1416
rect 968 1403 970 1415
rect 1080 1403 1082 1415
rect 967 1402 971 1403
rect 967 1397 971 1398
rect 975 1402 979 1403
rect 975 1397 979 1398
rect 1079 1402 1083 1403
rect 1079 1397 1083 1398
rect 1095 1402 1099 1403
rect 1095 1397 1099 1398
rect 974 1396 980 1397
rect 974 1392 975 1396
rect 979 1392 980 1396
rect 974 1391 980 1392
rect 1094 1396 1100 1397
rect 1094 1392 1095 1396
rect 1099 1392 1100 1396
rect 1094 1391 1100 1392
rect 1104 1368 1106 1438
rect 1670 1437 1676 1438
rect 1670 1433 1671 1437
rect 1675 1433 1676 1437
rect 1670 1432 1676 1433
rect 1630 1427 1636 1428
rect 1630 1423 1631 1427
rect 1635 1423 1636 1427
rect 1630 1422 1636 1423
rect 1190 1420 1196 1421
rect 1190 1416 1191 1420
rect 1195 1416 1196 1420
rect 1190 1415 1196 1416
rect 1310 1420 1316 1421
rect 1310 1416 1311 1420
rect 1315 1416 1316 1420
rect 1310 1415 1316 1416
rect 1192 1403 1194 1415
rect 1312 1403 1314 1415
rect 1632 1403 1634 1422
rect 2108 1420 2110 1478
rect 2230 1460 2236 1461
rect 2230 1456 2231 1460
rect 2235 1456 2236 1460
rect 2230 1455 2236 1456
rect 2232 1451 2234 1455
rect 2207 1450 2211 1451
rect 2207 1445 2211 1446
rect 2231 1450 2235 1451
rect 2231 1445 2235 1446
rect 2206 1444 2212 1445
rect 2206 1440 2207 1444
rect 2211 1440 2212 1444
rect 2206 1439 2212 1440
rect 2240 1424 2242 1482
rect 2374 1460 2380 1461
rect 2374 1456 2375 1460
rect 2379 1456 2380 1460
rect 2374 1455 2380 1456
rect 2376 1451 2378 1455
rect 2335 1450 2339 1451
rect 2335 1445 2339 1446
rect 2375 1450 2379 1451
rect 2375 1445 2379 1446
rect 2334 1444 2340 1445
rect 2334 1440 2335 1444
rect 2339 1440 2340 1444
rect 2334 1439 2340 1440
rect 2238 1423 2244 1424
rect 1670 1419 1676 1420
rect 1670 1415 1671 1419
rect 1675 1415 1676 1419
rect 2106 1419 2112 1420
rect 1670 1414 1676 1415
rect 1982 1415 1988 1416
rect 1191 1402 1195 1403
rect 1191 1397 1195 1398
rect 1215 1402 1219 1403
rect 1215 1397 1219 1398
rect 1311 1402 1315 1403
rect 1311 1397 1315 1398
rect 1631 1402 1635 1403
rect 1631 1397 1635 1398
rect 1214 1396 1220 1397
rect 1214 1392 1215 1396
rect 1219 1392 1220 1396
rect 1214 1391 1220 1392
rect 1632 1390 1634 1397
rect 1672 1395 1674 1414
rect 1982 1411 1983 1415
rect 1987 1411 1988 1415
rect 1982 1410 1988 1411
rect 1990 1415 1996 1416
rect 1990 1411 1991 1415
rect 1995 1411 1996 1415
rect 2094 1415 2100 1416
rect 2094 1411 2095 1415
rect 2099 1411 2100 1415
rect 2106 1415 2107 1419
rect 2111 1415 2112 1419
rect 2238 1419 2239 1423
rect 2243 1419 2244 1423
rect 2400 1420 2402 1482
rect 2479 1450 2483 1451
rect 2479 1445 2483 1446
rect 2478 1444 2484 1445
rect 2478 1440 2479 1444
rect 2483 1440 2484 1444
rect 2478 1439 2484 1440
rect 2488 1420 2490 1490
rect 2503 1489 2507 1490
rect 2510 1489 2516 1490
rect 2615 1489 2619 1490
rect 2654 1489 2660 1490
rect 2510 1485 2511 1489
rect 2515 1485 2516 1489
rect 2510 1484 2516 1485
rect 2654 1485 2655 1489
rect 2659 1485 2660 1489
rect 2664 1488 2666 1502
rect 2734 1499 2735 1503
rect 2739 1499 2740 1503
rect 2806 1503 2807 1507
rect 2811 1503 2812 1507
rect 2862 1507 2868 1508
rect 2806 1502 2812 1503
rect 2854 1503 2860 1504
rect 2734 1498 2740 1499
rect 2736 1495 2738 1498
rect 2735 1494 2739 1495
rect 2799 1494 2803 1495
rect 2735 1489 2739 1490
rect 2798 1489 2804 1490
rect 2654 1484 2660 1485
rect 2662 1487 2668 1488
rect 2662 1483 2663 1487
rect 2667 1483 2668 1487
rect 2798 1485 2799 1489
rect 2803 1485 2804 1489
rect 2808 1488 2810 1502
rect 2854 1499 2855 1503
rect 2859 1499 2860 1503
rect 2862 1503 2863 1507
rect 2867 1503 2868 1507
rect 2862 1502 2868 1503
rect 2918 1507 2924 1508
rect 2918 1503 2919 1507
rect 2923 1503 2924 1507
rect 3008 1504 3010 1570
rect 3111 1538 3115 1539
rect 3111 1533 3115 1534
rect 3110 1532 3116 1533
rect 3110 1528 3111 1532
rect 3115 1528 3116 1532
rect 3110 1527 3116 1528
rect 3120 1508 3122 1590
rect 3192 1587 3194 1590
rect 3191 1586 3195 1587
rect 3191 1581 3195 1582
rect 3192 1578 3194 1581
rect 3190 1577 3196 1578
rect 3190 1573 3191 1577
rect 3195 1573 3196 1577
rect 3190 1572 3196 1573
rect 3190 1559 3196 1560
rect 3190 1555 3191 1559
rect 3195 1555 3196 1559
rect 3190 1554 3196 1555
rect 3192 1539 3194 1554
rect 3191 1538 3195 1539
rect 3191 1533 3195 1534
rect 3192 1526 3194 1533
rect 3190 1525 3196 1526
rect 3190 1521 3191 1525
rect 3195 1521 3196 1525
rect 3190 1520 3196 1521
rect 3118 1507 3124 1508
rect 2918 1502 2924 1503
rect 2982 1503 2988 1504
rect 2854 1498 2860 1499
rect 2856 1495 2858 1498
rect 2855 1494 2859 1495
rect 2855 1489 2859 1490
rect 2798 1484 2804 1485
rect 2806 1487 2812 1488
rect 2662 1482 2668 1483
rect 2806 1483 2807 1487
rect 2811 1483 2812 1487
rect 2864 1484 2866 1502
rect 2982 1499 2983 1503
rect 2987 1499 2988 1503
rect 2982 1498 2988 1499
rect 3006 1503 3012 1504
rect 3006 1499 3007 1503
rect 3011 1499 3012 1503
rect 3006 1498 3012 1499
rect 3110 1503 3116 1504
rect 3110 1499 3111 1503
rect 3115 1499 3116 1503
rect 3118 1503 3119 1507
rect 3123 1503 3124 1507
rect 3118 1502 3124 1503
rect 3190 1507 3196 1508
rect 3190 1503 3191 1507
rect 3195 1503 3196 1507
rect 3190 1502 3196 1503
rect 3110 1498 3116 1499
rect 2984 1495 2986 1498
rect 2983 1494 2987 1495
rect 2983 1489 2987 1490
rect 2806 1482 2812 1483
rect 2862 1483 2868 1484
rect 2510 1460 2516 1461
rect 2510 1456 2511 1460
rect 2515 1456 2516 1460
rect 2510 1455 2516 1456
rect 2654 1460 2660 1461
rect 2654 1456 2655 1460
rect 2659 1456 2660 1460
rect 2654 1455 2660 1456
rect 2512 1451 2514 1455
rect 2656 1451 2658 1455
rect 2511 1450 2515 1451
rect 2511 1445 2515 1446
rect 2639 1450 2643 1451
rect 2639 1445 2643 1446
rect 2655 1450 2659 1451
rect 2655 1445 2659 1446
rect 2638 1444 2644 1445
rect 2638 1440 2639 1444
rect 2643 1440 2644 1444
rect 2638 1439 2644 1440
rect 2664 1420 2666 1482
rect 2862 1479 2863 1483
rect 2867 1479 2868 1483
rect 2862 1478 2868 1479
rect 2798 1460 2804 1461
rect 2798 1456 2799 1460
rect 2803 1456 2804 1460
rect 2798 1455 2804 1456
rect 2800 1451 2802 1455
rect 2799 1450 2803 1451
rect 2799 1445 2803 1446
rect 2815 1450 2819 1451
rect 2815 1445 2819 1446
rect 2814 1444 2820 1445
rect 2814 1440 2815 1444
rect 2819 1440 2820 1444
rect 2814 1439 2820 1440
rect 2864 1420 2866 1478
rect 2999 1450 3003 1451
rect 2999 1445 3003 1446
rect 2998 1444 3004 1445
rect 2998 1440 2999 1444
rect 3003 1440 3004 1444
rect 2998 1439 3004 1440
rect 3008 1424 3010 1498
rect 3112 1495 3114 1498
rect 3111 1494 3115 1495
rect 3111 1489 3115 1490
rect 3120 1424 3122 1502
rect 3192 1495 3194 1502
rect 3191 1494 3195 1495
rect 3191 1489 3195 1490
rect 3192 1486 3194 1489
rect 3190 1485 3196 1486
rect 3190 1481 3191 1485
rect 3195 1481 3196 1485
rect 3190 1480 3196 1481
rect 3190 1467 3196 1468
rect 3190 1463 3191 1467
rect 3195 1463 3196 1467
rect 3190 1462 3196 1463
rect 3192 1451 3194 1462
rect 3159 1450 3163 1451
rect 3159 1445 3163 1446
rect 3191 1450 3195 1451
rect 3191 1445 3195 1446
rect 3158 1444 3164 1445
rect 3158 1440 3159 1444
rect 3163 1440 3164 1444
rect 3158 1439 3164 1440
rect 3192 1438 3194 1445
rect 3190 1437 3196 1438
rect 3190 1433 3191 1437
rect 3195 1433 3196 1437
rect 3190 1432 3196 1433
rect 3006 1423 3012 1424
rect 2238 1418 2244 1419
rect 2398 1419 2404 1420
rect 2106 1414 2112 1415
rect 2206 1415 2212 1416
rect 1990 1410 2002 1411
rect 2094 1410 2100 1411
rect 2108 1411 2110 1414
rect 2206 1411 2207 1415
rect 2211 1411 2212 1415
rect 1984 1395 1986 1410
rect 1992 1409 2002 1410
rect 1671 1394 1675 1395
rect 1879 1394 1883 1395
rect 1983 1394 1987 1395
rect 1991 1394 1995 1395
rect 1630 1389 1636 1390
rect 1671 1389 1675 1390
rect 1878 1389 1884 1390
rect 1983 1389 1987 1390
rect 1990 1389 1996 1390
rect 1630 1385 1631 1389
rect 1635 1385 1636 1389
rect 1672 1386 1674 1389
rect 1630 1384 1636 1385
rect 1670 1385 1676 1386
rect 1670 1381 1671 1385
rect 1675 1381 1676 1385
rect 1878 1385 1879 1389
rect 1883 1385 1884 1389
rect 1878 1384 1884 1385
rect 1990 1385 1991 1389
rect 1995 1385 1996 1389
rect 1990 1384 1996 1385
rect 2000 1384 2002 1409
rect 2096 1395 2098 1410
rect 2108 1409 2114 1411
rect 2206 1410 2212 1411
rect 2095 1394 2099 1395
rect 2103 1394 2107 1395
rect 2095 1389 2099 1390
rect 2102 1389 2108 1390
rect 2102 1385 2103 1389
rect 2107 1385 2108 1389
rect 2102 1384 2108 1385
rect 2112 1384 2114 1409
rect 2208 1395 2210 1410
rect 2240 1403 2242 1418
rect 2334 1415 2340 1416
rect 2334 1411 2335 1415
rect 2339 1411 2340 1415
rect 2398 1415 2399 1419
rect 2403 1415 2404 1419
rect 2486 1419 2492 1420
rect 2398 1414 2404 1415
rect 2478 1415 2484 1416
rect 2334 1410 2340 1411
rect 2240 1401 2250 1403
rect 2207 1394 2211 1395
rect 2239 1394 2243 1395
rect 2207 1389 2211 1390
rect 2238 1389 2244 1390
rect 2238 1385 2239 1389
rect 2243 1385 2244 1389
rect 2248 1388 2250 1401
rect 2336 1395 2338 1410
rect 2335 1394 2339 1395
rect 2391 1394 2395 1395
rect 2335 1389 2339 1390
rect 2390 1389 2396 1390
rect 2238 1384 2244 1385
rect 2246 1387 2252 1388
rect 1670 1380 1676 1381
rect 1886 1383 1892 1384
rect 1886 1379 1887 1383
rect 1891 1379 1892 1383
rect 1998 1383 2004 1384
rect 1998 1379 1999 1383
rect 2003 1379 2004 1383
rect 1886 1378 1898 1379
rect 1998 1378 2004 1379
rect 2110 1383 2116 1384
rect 2110 1379 2111 1383
rect 2115 1379 2116 1383
rect 2246 1383 2247 1387
rect 2251 1383 2252 1387
rect 2390 1385 2391 1389
rect 2395 1385 2396 1389
rect 2400 1388 2402 1414
rect 2478 1411 2479 1415
rect 2483 1411 2484 1415
rect 2486 1415 2487 1419
rect 2491 1415 2492 1419
rect 2662 1419 2668 1420
rect 2486 1414 2492 1415
rect 2638 1415 2644 1416
rect 2478 1410 2484 1411
rect 2638 1411 2639 1415
rect 2643 1411 2644 1415
rect 2662 1415 2663 1419
rect 2667 1415 2668 1419
rect 2862 1419 2868 1420
rect 2662 1414 2668 1415
rect 2814 1415 2820 1416
rect 2638 1410 2644 1411
rect 2480 1395 2482 1410
rect 2640 1395 2642 1410
rect 2479 1394 2483 1395
rect 2567 1394 2571 1395
rect 2639 1394 2643 1395
rect 2479 1389 2483 1390
rect 2566 1389 2572 1390
rect 2639 1389 2643 1390
rect 2390 1384 2396 1385
rect 2398 1387 2404 1388
rect 2246 1382 2252 1383
rect 2398 1383 2399 1387
rect 2403 1383 2404 1387
rect 2566 1385 2567 1389
rect 2571 1385 2572 1389
rect 2664 1388 2666 1414
rect 2814 1411 2815 1415
rect 2819 1411 2820 1415
rect 2814 1410 2820 1411
rect 2822 1415 2828 1416
rect 2822 1411 2823 1415
rect 2827 1411 2828 1415
rect 2862 1415 2863 1419
rect 2867 1415 2868 1419
rect 3006 1419 3007 1423
rect 3011 1419 3012 1423
rect 3006 1418 3012 1419
rect 3118 1423 3124 1424
rect 3118 1419 3119 1423
rect 3123 1419 3124 1423
rect 3118 1418 3124 1419
rect 3166 1419 3172 1420
rect 2862 1414 2868 1415
rect 2998 1415 3004 1416
rect 2822 1410 2828 1411
rect 2998 1411 2999 1415
rect 3003 1411 3004 1415
rect 2998 1410 3004 1411
rect 2816 1395 2818 1410
rect 2767 1394 2771 1395
rect 2815 1394 2819 1395
rect 2766 1389 2772 1390
rect 2815 1389 2819 1390
rect 2566 1384 2572 1385
rect 2662 1387 2668 1388
rect 2398 1382 2404 1383
rect 2662 1383 2663 1387
rect 2667 1383 2668 1387
rect 2766 1385 2767 1389
rect 2771 1385 2772 1389
rect 2824 1388 2826 1410
rect 3000 1395 3002 1410
rect 2975 1394 2979 1395
rect 2999 1394 3003 1395
rect 2974 1389 2980 1390
rect 2999 1389 3003 1390
rect 2766 1384 2772 1385
rect 2822 1387 2828 1388
rect 2662 1382 2668 1383
rect 2822 1383 2823 1387
rect 2827 1383 2828 1387
rect 2974 1385 2975 1389
rect 2979 1385 2980 1389
rect 3008 1388 3010 1418
rect 3158 1415 3164 1416
rect 3158 1411 3159 1415
rect 3163 1411 3164 1415
rect 3166 1415 3167 1419
rect 3171 1415 3172 1419
rect 3166 1414 3172 1415
rect 3190 1419 3196 1420
rect 3190 1415 3191 1419
rect 3195 1415 3196 1419
rect 3190 1414 3196 1415
rect 3158 1410 3164 1411
rect 3160 1395 3162 1410
rect 3159 1394 3163 1395
rect 3158 1389 3164 1390
rect 2974 1384 2980 1385
rect 2982 1387 2988 1388
rect 2822 1382 2828 1383
rect 2982 1383 2983 1387
rect 2987 1383 2988 1387
rect 2982 1382 2988 1383
rect 3006 1387 3012 1388
rect 3006 1383 3007 1387
rect 3011 1383 3012 1387
rect 3158 1385 3159 1389
rect 3163 1385 3164 1389
rect 3168 1388 3170 1414
rect 3192 1395 3194 1414
rect 3191 1394 3195 1395
rect 3191 1389 3195 1390
rect 3158 1384 3164 1385
rect 3166 1387 3172 1388
rect 3006 1382 3012 1383
rect 3166 1383 3167 1387
rect 3171 1383 3172 1387
rect 3192 1386 3194 1389
rect 3166 1382 3172 1383
rect 3190 1385 3196 1386
rect 2110 1378 2116 1379
rect 1888 1377 1898 1378
rect 1630 1371 1636 1372
rect 110 1366 116 1367
rect 374 1367 380 1368
rect 112 1355 114 1366
rect 374 1363 375 1367
rect 379 1363 380 1367
rect 374 1362 380 1363
rect 382 1367 388 1368
rect 382 1363 383 1367
rect 387 1363 388 1367
rect 382 1362 388 1363
rect 502 1367 508 1368
rect 502 1363 503 1367
rect 507 1363 508 1367
rect 502 1362 508 1363
rect 534 1367 540 1368
rect 534 1363 535 1367
rect 539 1363 540 1367
rect 534 1362 540 1363
rect 622 1367 628 1368
rect 622 1363 623 1367
rect 627 1363 628 1367
rect 622 1362 628 1363
rect 634 1367 640 1368
rect 634 1363 635 1367
rect 639 1363 640 1367
rect 634 1362 640 1363
rect 742 1367 748 1368
rect 742 1363 743 1367
rect 747 1363 748 1367
rect 742 1362 748 1363
rect 786 1367 792 1368
rect 786 1363 787 1367
rect 791 1363 792 1367
rect 786 1362 792 1363
rect 862 1367 868 1368
rect 862 1363 863 1367
rect 867 1363 868 1367
rect 862 1362 868 1363
rect 886 1367 892 1368
rect 886 1363 887 1367
rect 891 1363 892 1367
rect 886 1362 892 1363
rect 974 1367 980 1368
rect 974 1363 975 1367
rect 979 1363 980 1367
rect 974 1362 980 1363
rect 1014 1367 1020 1368
rect 1014 1363 1015 1367
rect 1019 1363 1020 1367
rect 1014 1362 1020 1363
rect 1094 1367 1100 1368
rect 1094 1363 1095 1367
rect 1099 1363 1100 1367
rect 1094 1362 1100 1363
rect 1102 1367 1108 1368
rect 1102 1363 1103 1367
rect 1107 1363 1108 1367
rect 1102 1362 1108 1363
rect 1214 1367 1220 1368
rect 1214 1363 1215 1367
rect 1219 1363 1220 1367
rect 1630 1367 1631 1371
rect 1635 1367 1636 1371
rect 1630 1366 1636 1367
rect 1670 1367 1676 1368
rect 1214 1362 1220 1363
rect 376 1355 378 1362
rect 111 1354 115 1355
rect 271 1354 275 1355
rect 375 1354 379 1355
rect 111 1349 115 1350
rect 270 1349 276 1350
rect 375 1349 379 1350
rect 112 1346 114 1349
rect 110 1345 116 1346
rect 110 1341 111 1345
rect 115 1341 116 1345
rect 270 1345 271 1349
rect 275 1345 276 1349
rect 270 1344 276 1345
rect 384 1344 386 1362
rect 504 1355 506 1362
rect 399 1354 403 1355
rect 503 1354 507 1355
rect 527 1354 531 1355
rect 398 1349 404 1350
rect 503 1349 507 1350
rect 526 1349 532 1350
rect 398 1345 399 1349
rect 403 1345 404 1349
rect 398 1344 404 1345
rect 526 1345 527 1349
rect 531 1345 532 1349
rect 526 1344 532 1345
rect 536 1344 538 1362
rect 624 1355 626 1362
rect 623 1354 627 1355
rect 623 1349 627 1350
rect 636 1344 638 1362
rect 744 1355 746 1362
rect 647 1354 651 1355
rect 743 1354 747 1355
rect 767 1354 771 1355
rect 646 1349 652 1350
rect 743 1349 747 1350
rect 766 1349 772 1350
rect 646 1345 647 1349
rect 651 1345 652 1349
rect 646 1344 652 1345
rect 766 1345 767 1349
rect 771 1345 772 1349
rect 766 1344 772 1345
rect 788 1344 790 1362
rect 864 1355 866 1362
rect 863 1354 867 1355
rect 879 1354 883 1355
rect 863 1349 867 1350
rect 878 1349 884 1350
rect 878 1345 879 1349
rect 883 1345 884 1349
rect 878 1344 884 1345
rect 888 1344 890 1362
rect 976 1355 978 1362
rect 975 1354 979 1355
rect 991 1354 995 1355
rect 975 1349 979 1350
rect 990 1349 996 1350
rect 990 1345 991 1349
rect 995 1345 996 1349
rect 990 1344 996 1345
rect 1016 1344 1018 1362
rect 1096 1355 1098 1362
rect 1095 1354 1099 1355
rect 1095 1349 1099 1350
rect 1104 1344 1106 1362
rect 1216 1355 1218 1362
rect 1632 1355 1634 1366
rect 1670 1363 1671 1367
rect 1675 1363 1676 1367
rect 1670 1362 1676 1363
rect 1111 1354 1115 1355
rect 1215 1354 1219 1355
rect 1110 1349 1116 1350
rect 1215 1349 1219 1350
rect 1631 1354 1635 1355
rect 1631 1349 1635 1350
rect 1110 1345 1111 1349
rect 1115 1345 1116 1349
rect 1632 1346 1634 1349
rect 1110 1344 1116 1345
rect 1630 1345 1636 1346
rect 110 1340 116 1341
rect 310 1343 316 1344
rect 310 1339 311 1343
rect 315 1339 316 1343
rect 310 1338 316 1339
rect 382 1343 388 1344
rect 382 1339 383 1343
rect 387 1339 388 1343
rect 382 1338 388 1339
rect 534 1343 540 1344
rect 534 1339 535 1343
rect 539 1339 540 1343
rect 534 1338 540 1339
rect 634 1343 640 1344
rect 634 1339 635 1343
rect 639 1339 640 1343
rect 634 1338 640 1339
rect 786 1343 792 1344
rect 786 1339 787 1343
rect 791 1339 792 1343
rect 786 1338 792 1339
rect 887 1343 893 1344
rect 887 1339 888 1343
rect 892 1342 893 1343
rect 1014 1343 1020 1344
rect 892 1340 898 1342
rect 892 1339 893 1340
rect 887 1338 893 1339
rect 110 1327 116 1328
rect 110 1323 111 1327
rect 115 1323 116 1327
rect 110 1322 116 1323
rect 112 1303 114 1322
rect 270 1320 276 1321
rect 270 1316 271 1320
rect 275 1316 276 1320
rect 270 1315 276 1316
rect 272 1303 274 1315
rect 111 1302 115 1303
rect 111 1297 115 1298
rect 175 1302 179 1303
rect 175 1297 179 1298
rect 271 1302 275 1303
rect 271 1297 275 1298
rect 303 1302 307 1303
rect 303 1297 307 1298
rect 112 1290 114 1297
rect 174 1296 180 1297
rect 174 1292 175 1296
rect 179 1292 180 1296
rect 174 1291 180 1292
rect 302 1296 308 1297
rect 302 1292 303 1296
rect 307 1292 308 1296
rect 302 1291 308 1292
rect 110 1289 116 1290
rect 110 1285 111 1289
rect 115 1285 116 1289
rect 110 1284 116 1285
rect 312 1272 314 1338
rect 398 1320 404 1321
rect 398 1316 399 1320
rect 403 1316 404 1320
rect 398 1315 404 1316
rect 526 1320 532 1321
rect 526 1316 527 1320
rect 531 1316 532 1320
rect 526 1315 532 1316
rect 400 1303 402 1315
rect 528 1303 530 1315
rect 399 1302 403 1303
rect 399 1297 403 1298
rect 423 1302 427 1303
rect 423 1297 427 1298
rect 527 1302 531 1303
rect 527 1297 531 1298
rect 543 1302 547 1303
rect 543 1297 547 1298
rect 422 1296 428 1297
rect 422 1292 423 1296
rect 427 1292 428 1296
rect 422 1291 428 1292
rect 542 1296 548 1297
rect 542 1292 543 1296
rect 547 1292 548 1296
rect 542 1291 548 1292
rect 636 1272 638 1338
rect 646 1320 652 1321
rect 646 1316 647 1320
rect 651 1316 652 1320
rect 646 1315 652 1316
rect 766 1320 772 1321
rect 766 1316 767 1320
rect 771 1316 772 1320
rect 766 1315 772 1316
rect 648 1303 650 1315
rect 768 1303 770 1315
rect 647 1302 651 1303
rect 647 1297 651 1298
rect 663 1302 667 1303
rect 663 1297 667 1298
rect 767 1302 771 1303
rect 767 1297 771 1298
rect 775 1302 779 1303
rect 775 1297 779 1298
rect 662 1296 668 1297
rect 662 1292 663 1296
rect 667 1292 668 1296
rect 662 1291 668 1292
rect 774 1296 780 1297
rect 774 1292 775 1296
rect 779 1292 780 1296
rect 774 1291 780 1292
rect 110 1271 116 1272
rect 110 1267 111 1271
rect 115 1267 116 1271
rect 310 1271 316 1272
rect 110 1266 116 1267
rect 174 1267 180 1268
rect 112 1251 114 1266
rect 174 1263 175 1267
rect 179 1263 180 1267
rect 174 1262 180 1263
rect 186 1267 192 1268
rect 186 1263 187 1267
rect 191 1263 192 1267
rect 186 1262 192 1263
rect 302 1267 308 1268
rect 302 1263 303 1267
rect 307 1263 308 1267
rect 310 1267 311 1271
rect 315 1267 316 1271
rect 550 1271 556 1272
rect 310 1266 316 1267
rect 422 1267 428 1268
rect 302 1262 308 1263
rect 176 1251 178 1262
rect 111 1250 115 1251
rect 135 1250 139 1251
rect 175 1250 179 1251
rect 111 1245 115 1246
rect 134 1245 140 1246
rect 175 1245 179 1246
rect 112 1242 114 1245
rect 110 1241 116 1242
rect 110 1237 111 1241
rect 115 1237 116 1241
rect 134 1241 135 1245
rect 139 1241 140 1245
rect 134 1240 140 1241
rect 188 1240 190 1262
rect 304 1251 306 1262
rect 231 1250 235 1251
rect 303 1250 307 1251
rect 230 1245 236 1246
rect 303 1245 307 1246
rect 230 1241 231 1245
rect 235 1241 236 1245
rect 230 1240 236 1241
rect 312 1240 314 1266
rect 422 1263 423 1267
rect 427 1263 428 1267
rect 422 1262 428 1263
rect 430 1267 436 1268
rect 430 1263 431 1267
rect 435 1263 436 1267
rect 430 1262 436 1263
rect 542 1267 548 1268
rect 542 1263 543 1267
rect 547 1263 548 1267
rect 550 1267 551 1271
rect 555 1267 556 1271
rect 550 1266 556 1267
rect 634 1271 640 1272
rect 634 1267 635 1271
rect 639 1267 640 1271
rect 788 1268 790 1338
rect 878 1320 884 1321
rect 878 1316 879 1320
rect 883 1316 884 1320
rect 878 1315 884 1316
rect 880 1303 882 1315
rect 879 1302 883 1303
rect 879 1297 883 1298
rect 887 1302 891 1303
rect 887 1297 891 1298
rect 886 1296 892 1297
rect 886 1292 887 1296
rect 891 1292 892 1296
rect 886 1291 892 1292
rect 896 1268 898 1340
rect 1014 1339 1015 1343
rect 1019 1339 1020 1343
rect 1014 1338 1020 1339
rect 1102 1343 1108 1344
rect 1102 1339 1103 1343
rect 1107 1339 1108 1343
rect 1630 1341 1631 1345
rect 1635 1341 1636 1345
rect 1672 1343 1674 1362
rect 1878 1360 1884 1361
rect 1878 1356 1879 1360
rect 1883 1356 1884 1360
rect 1878 1355 1884 1356
rect 1880 1343 1882 1355
rect 1630 1340 1636 1341
rect 1671 1342 1675 1343
rect 1102 1338 1108 1339
rect 990 1320 996 1321
rect 990 1316 991 1320
rect 995 1316 996 1320
rect 990 1315 996 1316
rect 992 1303 994 1315
rect 991 1302 995 1303
rect 991 1297 995 1298
rect 1007 1302 1011 1303
rect 1007 1297 1011 1298
rect 1006 1296 1012 1297
rect 1006 1292 1007 1296
rect 1011 1292 1012 1296
rect 1006 1291 1012 1292
rect 1016 1268 1018 1338
rect 1671 1337 1675 1338
rect 1775 1342 1779 1343
rect 1775 1337 1779 1338
rect 1879 1342 1883 1343
rect 1879 1337 1883 1338
rect 1887 1342 1891 1343
rect 1887 1337 1891 1338
rect 1672 1330 1674 1337
rect 1774 1336 1780 1337
rect 1774 1332 1775 1336
rect 1779 1332 1780 1336
rect 1774 1331 1780 1332
rect 1886 1336 1892 1337
rect 1886 1332 1887 1336
rect 1891 1332 1892 1336
rect 1886 1331 1892 1332
rect 1670 1329 1676 1330
rect 1630 1327 1636 1328
rect 1630 1323 1631 1327
rect 1635 1323 1636 1327
rect 1670 1325 1671 1329
rect 1675 1325 1676 1329
rect 1670 1324 1676 1325
rect 1630 1322 1636 1323
rect 1110 1320 1116 1321
rect 1110 1316 1111 1320
rect 1115 1316 1116 1320
rect 1110 1315 1116 1316
rect 1112 1303 1114 1315
rect 1632 1303 1634 1322
rect 1896 1316 1898 1377
rect 1990 1360 1996 1361
rect 1990 1356 1991 1360
rect 1995 1356 1996 1360
rect 1990 1355 1996 1356
rect 1992 1343 1994 1355
rect 1991 1342 1995 1343
rect 1991 1337 1995 1338
rect 1990 1336 1996 1337
rect 1990 1332 1991 1336
rect 1995 1332 1996 1336
rect 1990 1331 1996 1332
rect 2000 1316 2002 1378
rect 2102 1360 2108 1361
rect 2102 1356 2103 1360
rect 2107 1356 2108 1360
rect 2102 1355 2108 1356
rect 2238 1360 2244 1361
rect 2238 1356 2239 1360
rect 2243 1356 2244 1360
rect 2238 1355 2244 1356
rect 2390 1360 2396 1361
rect 2390 1356 2391 1360
rect 2395 1356 2396 1360
rect 2390 1355 2396 1356
rect 2104 1343 2106 1355
rect 2240 1343 2242 1355
rect 2392 1343 2394 1355
rect 2095 1342 2099 1343
rect 2095 1337 2099 1338
rect 2103 1342 2107 1343
rect 2103 1337 2107 1338
rect 2199 1342 2203 1343
rect 2199 1337 2203 1338
rect 2239 1342 2243 1343
rect 2239 1337 2243 1338
rect 2303 1342 2307 1343
rect 2303 1337 2307 1338
rect 2391 1342 2395 1343
rect 2391 1337 2395 1338
rect 2094 1336 2100 1337
rect 2094 1332 2095 1336
rect 2099 1332 2100 1336
rect 2094 1331 2100 1332
rect 2198 1336 2204 1337
rect 2198 1332 2199 1336
rect 2203 1332 2204 1336
rect 2198 1331 2204 1332
rect 2302 1336 2308 1337
rect 2302 1332 2303 1336
rect 2307 1332 2308 1336
rect 2302 1331 2308 1332
rect 2400 1316 2402 1382
rect 2566 1360 2572 1361
rect 2566 1356 2567 1360
rect 2571 1356 2572 1360
rect 2566 1355 2572 1356
rect 2766 1360 2772 1361
rect 2766 1356 2767 1360
rect 2771 1356 2772 1360
rect 2766 1355 2772 1356
rect 2974 1360 2980 1361
rect 2974 1356 2975 1360
rect 2979 1356 2980 1360
rect 2974 1355 2980 1356
rect 2568 1343 2570 1355
rect 2768 1343 2770 1355
rect 2976 1343 2978 1355
rect 2407 1342 2411 1343
rect 2407 1337 2411 1338
rect 2511 1342 2515 1343
rect 2511 1337 2515 1338
rect 2567 1342 2571 1343
rect 2567 1337 2571 1338
rect 2767 1342 2771 1343
rect 2767 1337 2771 1338
rect 2975 1342 2979 1343
rect 2975 1337 2979 1338
rect 2406 1336 2412 1337
rect 2406 1332 2407 1336
rect 2411 1332 2412 1336
rect 2406 1331 2412 1332
rect 2510 1336 2516 1337
rect 2510 1332 2511 1336
rect 2515 1332 2516 1336
rect 2510 1331 2516 1332
rect 1894 1315 1900 1316
rect 1670 1311 1676 1312
rect 1670 1307 1671 1311
rect 1675 1307 1676 1311
rect 1894 1311 1895 1315
rect 1899 1311 1900 1315
rect 1998 1315 2004 1316
rect 1894 1310 1900 1311
rect 1942 1311 1948 1312
rect 1670 1306 1676 1307
rect 1774 1307 1780 1308
rect 1111 1302 1115 1303
rect 1111 1297 1115 1298
rect 1631 1302 1635 1303
rect 1631 1297 1635 1298
rect 1632 1290 1634 1297
rect 1672 1295 1674 1306
rect 1774 1303 1775 1307
rect 1779 1303 1780 1307
rect 1774 1302 1780 1303
rect 1782 1307 1788 1308
rect 1782 1303 1783 1307
rect 1787 1303 1788 1307
rect 1782 1302 1788 1303
rect 1886 1307 1892 1308
rect 1886 1303 1887 1307
rect 1891 1303 1892 1307
rect 1942 1307 1943 1311
rect 1947 1307 1948 1311
rect 1998 1311 1999 1315
rect 2003 1311 2004 1315
rect 1998 1310 2004 1311
rect 2102 1315 2108 1316
rect 2102 1311 2103 1315
rect 2107 1311 2108 1315
rect 2102 1310 2108 1311
rect 2398 1315 2404 1316
rect 2398 1311 2399 1315
rect 2403 1311 2404 1315
rect 2398 1310 2404 1311
rect 2502 1315 2508 1316
rect 2502 1311 2503 1315
rect 2507 1311 2508 1315
rect 2502 1310 2508 1311
rect 1942 1306 1948 1307
rect 1990 1307 1996 1308
rect 1886 1302 1892 1303
rect 1776 1295 1778 1302
rect 1671 1294 1675 1295
rect 1695 1294 1699 1295
rect 1775 1294 1779 1295
rect 1630 1289 1636 1290
rect 1671 1289 1675 1290
rect 1694 1289 1700 1290
rect 1775 1289 1779 1290
rect 1630 1285 1631 1289
rect 1635 1285 1636 1289
rect 1672 1286 1674 1289
rect 1630 1284 1636 1285
rect 1670 1285 1676 1286
rect 1670 1281 1671 1285
rect 1675 1281 1676 1285
rect 1694 1285 1695 1289
rect 1699 1285 1700 1289
rect 1694 1284 1700 1285
rect 1784 1284 1786 1302
rect 1888 1295 1890 1302
rect 1791 1294 1795 1295
rect 1887 1294 1891 1295
rect 1935 1294 1939 1295
rect 1790 1289 1796 1290
rect 1887 1289 1891 1290
rect 1934 1289 1940 1290
rect 1790 1285 1791 1289
rect 1795 1285 1796 1289
rect 1790 1284 1796 1285
rect 1934 1285 1935 1289
rect 1939 1285 1940 1289
rect 1944 1288 1946 1306
rect 1990 1303 1991 1307
rect 1995 1303 1996 1307
rect 1990 1302 1996 1303
rect 2094 1307 2100 1308
rect 2094 1303 2095 1307
rect 2099 1303 2100 1307
rect 2094 1302 2100 1303
rect 1992 1295 1994 1302
rect 2096 1295 2098 1302
rect 2104 1299 2106 1310
rect 2198 1307 2204 1308
rect 2198 1303 2199 1307
rect 2203 1303 2204 1307
rect 2198 1302 2204 1303
rect 2302 1307 2308 1308
rect 2302 1303 2303 1307
rect 2307 1303 2308 1307
rect 2302 1302 2308 1303
rect 2406 1307 2412 1308
rect 2406 1303 2407 1307
rect 2411 1303 2412 1307
rect 2406 1302 2412 1303
rect 2110 1299 2116 1300
rect 2104 1297 2111 1299
rect 2110 1295 2111 1297
rect 2115 1295 2116 1299
rect 2200 1295 2202 1302
rect 2304 1295 2306 1302
rect 2408 1295 2410 1302
rect 1991 1294 1995 1295
rect 1991 1289 1995 1290
rect 2095 1294 2099 1295
rect 2103 1294 2107 1295
rect 2110 1294 2116 1295
rect 2199 1294 2203 1295
rect 2095 1289 2099 1290
rect 2102 1289 2108 1290
rect 1934 1284 1940 1285
rect 1942 1287 1948 1288
rect 1670 1280 1676 1281
rect 1702 1283 1708 1284
rect 1702 1279 1703 1283
rect 1707 1279 1708 1283
rect 1702 1278 1708 1279
rect 1782 1283 1788 1284
rect 1782 1279 1783 1283
rect 1787 1279 1788 1283
rect 1942 1283 1943 1287
rect 1947 1283 1948 1287
rect 2102 1285 2103 1289
rect 2107 1285 2108 1289
rect 2112 1288 2114 1294
rect 2295 1294 2299 1295
rect 2303 1294 2307 1295
rect 2199 1289 2203 1290
rect 2294 1289 2300 1290
rect 2303 1289 2307 1290
rect 2407 1294 2411 1295
rect 2495 1294 2499 1295
rect 2407 1289 2411 1290
rect 2494 1289 2500 1290
rect 2102 1284 2108 1285
rect 2110 1287 2116 1288
rect 1942 1282 1948 1283
rect 2110 1283 2111 1287
rect 2115 1283 2116 1287
rect 2294 1285 2295 1289
rect 2299 1285 2300 1289
rect 2294 1284 2300 1285
rect 2494 1285 2495 1289
rect 2499 1285 2500 1289
rect 2504 1288 2506 1310
rect 2510 1307 2516 1308
rect 2510 1303 2511 1307
rect 2515 1303 2516 1307
rect 2510 1302 2516 1303
rect 2512 1295 2514 1302
rect 2511 1294 2515 1295
rect 2711 1294 2715 1295
rect 2935 1294 2939 1295
rect 2511 1289 2515 1290
rect 2710 1289 2716 1290
rect 2494 1284 2500 1285
rect 2502 1287 2508 1288
rect 2110 1282 2116 1283
rect 2502 1283 2503 1287
rect 2507 1283 2508 1287
rect 2710 1285 2711 1289
rect 2715 1285 2716 1289
rect 2710 1284 2716 1285
rect 2934 1289 2940 1290
rect 2934 1285 2935 1289
rect 2939 1285 2940 1289
rect 2984 1288 2986 1382
rect 3158 1360 3164 1361
rect 3158 1356 3159 1360
rect 3163 1356 3164 1360
rect 3158 1355 3164 1356
rect 3160 1343 3162 1355
rect 3159 1342 3163 1343
rect 3159 1337 3163 1338
rect 3159 1294 3163 1295
rect 3158 1289 3164 1290
rect 2934 1284 2940 1285
rect 2982 1287 2988 1288
rect 2502 1282 2508 1283
rect 2718 1283 2724 1284
rect 1782 1278 1788 1279
rect 1630 1271 1636 1272
rect 634 1266 640 1267
rect 662 1267 668 1268
rect 542 1262 548 1263
rect 424 1251 426 1262
rect 359 1250 363 1251
rect 423 1250 427 1251
rect 358 1245 364 1246
rect 423 1245 427 1246
rect 358 1241 359 1245
rect 363 1241 364 1245
rect 358 1240 364 1241
rect 432 1240 434 1262
rect 544 1251 546 1262
rect 503 1250 507 1251
rect 543 1250 547 1251
rect 502 1245 508 1246
rect 543 1245 547 1246
rect 502 1241 503 1245
rect 507 1241 508 1245
rect 552 1244 554 1266
rect 662 1263 663 1267
rect 667 1263 668 1267
rect 662 1262 668 1263
rect 670 1267 676 1268
rect 670 1263 671 1267
rect 675 1263 676 1267
rect 670 1262 676 1263
rect 774 1267 780 1268
rect 774 1263 775 1267
rect 779 1263 780 1267
rect 774 1262 780 1263
rect 786 1267 792 1268
rect 786 1263 787 1267
rect 791 1263 792 1267
rect 786 1262 792 1263
rect 886 1267 892 1268
rect 886 1263 887 1267
rect 891 1263 892 1267
rect 886 1262 892 1263
rect 894 1267 900 1268
rect 894 1263 895 1267
rect 899 1263 900 1267
rect 894 1262 900 1263
rect 1006 1267 1012 1268
rect 1006 1263 1007 1267
rect 1011 1263 1012 1267
rect 1006 1262 1012 1263
rect 1015 1267 1021 1268
rect 1015 1263 1016 1267
rect 1020 1266 1021 1267
rect 1630 1267 1631 1271
rect 1635 1267 1636 1271
rect 1630 1266 1636 1267
rect 1670 1267 1676 1268
rect 1020 1264 1026 1266
rect 1020 1263 1021 1264
rect 1015 1262 1021 1263
rect 664 1251 666 1262
rect 663 1250 667 1251
rect 662 1245 668 1246
rect 502 1240 508 1241
rect 550 1243 556 1244
rect 110 1236 116 1237
rect 186 1239 192 1240
rect 186 1235 187 1239
rect 191 1235 192 1239
rect 186 1234 192 1235
rect 258 1239 264 1240
rect 258 1235 259 1239
rect 263 1235 264 1239
rect 258 1234 264 1235
rect 310 1239 316 1240
rect 310 1235 311 1239
rect 315 1235 316 1239
rect 310 1234 316 1235
rect 430 1239 436 1240
rect 430 1235 431 1239
rect 435 1235 436 1239
rect 550 1239 551 1243
rect 555 1239 556 1243
rect 662 1241 663 1245
rect 667 1241 668 1245
rect 662 1240 668 1241
rect 672 1240 674 1262
rect 776 1251 778 1262
rect 775 1250 779 1251
rect 775 1245 779 1246
rect 788 1240 790 1262
rect 866 1259 872 1260
rect 866 1255 867 1259
rect 871 1255 872 1259
rect 866 1254 872 1255
rect 831 1250 835 1251
rect 830 1245 836 1246
rect 830 1241 831 1245
rect 835 1241 836 1245
rect 830 1240 836 1241
rect 868 1240 870 1254
rect 888 1251 890 1262
rect 1008 1251 1010 1262
rect 887 1250 891 1251
rect 887 1245 891 1246
rect 1007 1250 1011 1251
rect 1015 1250 1019 1251
rect 1007 1245 1011 1246
rect 1014 1245 1020 1246
rect 1014 1241 1015 1245
rect 1019 1241 1020 1245
rect 1014 1240 1020 1241
rect 1024 1240 1026 1264
rect 1632 1251 1634 1266
rect 1670 1263 1671 1267
rect 1675 1263 1676 1267
rect 1670 1262 1676 1263
rect 1207 1250 1211 1251
rect 1407 1250 1411 1251
rect 1599 1250 1603 1251
rect 1631 1250 1635 1251
rect 1206 1245 1212 1246
rect 1206 1241 1207 1245
rect 1211 1241 1212 1245
rect 1206 1240 1212 1241
rect 1406 1245 1412 1246
rect 1406 1241 1407 1245
rect 1411 1241 1412 1245
rect 1406 1240 1412 1241
rect 1598 1245 1604 1246
rect 1631 1245 1635 1246
rect 1598 1241 1599 1245
rect 1603 1241 1604 1245
rect 1632 1242 1634 1245
rect 1598 1240 1604 1241
rect 1630 1241 1636 1242
rect 550 1238 556 1239
rect 670 1239 676 1240
rect 430 1234 436 1235
rect 670 1235 671 1239
rect 675 1235 676 1239
rect 670 1234 676 1235
rect 786 1239 792 1240
rect 786 1235 787 1239
rect 791 1235 792 1239
rect 786 1234 792 1235
rect 866 1239 872 1240
rect 866 1235 867 1239
rect 871 1235 872 1239
rect 866 1234 872 1235
rect 1006 1239 1012 1240
rect 1006 1235 1007 1239
rect 1011 1235 1012 1239
rect 1006 1234 1012 1235
rect 1022 1239 1028 1240
rect 1022 1235 1023 1239
rect 1027 1235 1028 1239
rect 1022 1234 1028 1235
rect 1230 1239 1236 1240
rect 1230 1235 1231 1239
rect 1235 1235 1236 1239
rect 1230 1234 1236 1235
rect 1454 1239 1460 1240
rect 1454 1235 1455 1239
rect 1459 1235 1460 1239
rect 1454 1234 1460 1235
rect 1606 1239 1612 1240
rect 1606 1235 1607 1239
rect 1611 1235 1612 1239
rect 1630 1237 1631 1241
rect 1635 1237 1636 1241
rect 1672 1239 1674 1262
rect 1694 1260 1700 1261
rect 1694 1256 1695 1260
rect 1699 1256 1700 1260
rect 1694 1255 1700 1256
rect 1696 1239 1698 1255
rect 1630 1236 1636 1237
rect 1671 1238 1675 1239
rect 1606 1234 1612 1235
rect 110 1223 116 1224
rect 110 1219 111 1223
rect 115 1219 116 1223
rect 110 1218 116 1219
rect 112 1203 114 1218
rect 134 1216 140 1217
rect 134 1212 135 1216
rect 139 1212 140 1216
rect 134 1211 140 1212
rect 230 1216 236 1217
rect 230 1212 231 1216
rect 235 1212 236 1216
rect 230 1211 236 1212
rect 136 1203 138 1211
rect 232 1203 234 1211
rect 111 1202 115 1203
rect 111 1197 115 1198
rect 135 1202 139 1203
rect 135 1197 139 1198
rect 231 1202 235 1203
rect 231 1197 235 1198
rect 112 1190 114 1197
rect 110 1189 116 1190
rect 110 1185 111 1189
rect 115 1185 116 1189
rect 110 1184 116 1185
rect 110 1171 116 1172
rect 110 1167 111 1171
rect 115 1167 116 1171
rect 110 1166 116 1167
rect 112 1151 114 1166
rect 111 1150 115 1151
rect 111 1145 115 1146
rect 112 1142 114 1145
rect 110 1141 116 1142
rect 110 1137 111 1141
rect 115 1137 116 1141
rect 110 1136 116 1137
rect 110 1123 116 1124
rect 110 1119 111 1123
rect 115 1119 116 1123
rect 110 1118 116 1119
rect 112 1099 114 1118
rect 111 1098 115 1099
rect 111 1093 115 1094
rect 112 1086 114 1093
rect 110 1085 116 1086
rect 110 1081 111 1085
rect 115 1081 116 1085
rect 110 1080 116 1081
rect 110 1067 116 1068
rect 110 1063 111 1067
rect 115 1063 116 1067
rect 110 1062 116 1063
rect 112 1051 114 1062
rect 111 1050 115 1051
rect 111 1045 115 1046
rect 112 1042 114 1045
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 110 1036 116 1037
rect 110 1023 116 1024
rect 110 1019 111 1023
rect 115 1019 116 1023
rect 110 1018 116 1019
rect 112 999 114 1018
rect 111 998 115 999
rect 111 993 115 994
rect 112 986 114 993
rect 110 985 116 986
rect 110 981 111 985
rect 115 981 116 985
rect 110 980 116 981
rect 110 967 116 968
rect 110 963 111 967
rect 115 963 116 967
rect 110 962 116 963
rect 112 947 114 962
rect 111 946 115 947
rect 223 946 227 947
rect 111 941 115 942
rect 222 941 228 942
rect 112 938 114 941
rect 110 937 116 938
rect 110 933 111 937
rect 115 933 116 937
rect 222 937 223 941
rect 227 937 228 941
rect 260 940 262 1234
rect 358 1216 364 1217
rect 358 1212 359 1216
rect 363 1212 364 1216
rect 358 1211 364 1212
rect 502 1216 508 1217
rect 502 1212 503 1216
rect 507 1212 508 1216
rect 502 1211 508 1212
rect 662 1216 668 1217
rect 662 1212 663 1216
rect 667 1212 668 1216
rect 662 1211 668 1212
rect 360 1203 362 1211
rect 504 1203 506 1211
rect 664 1203 666 1211
rect 359 1202 363 1203
rect 359 1197 363 1198
rect 503 1202 507 1203
rect 503 1197 507 1198
rect 663 1202 667 1203
rect 663 1197 667 1198
rect 631 1150 635 1151
rect 630 1145 636 1146
rect 630 1141 631 1145
rect 635 1141 636 1145
rect 630 1140 636 1141
rect 672 1140 674 1234
rect 830 1216 836 1217
rect 830 1212 831 1216
rect 835 1212 836 1216
rect 830 1211 836 1212
rect 832 1203 834 1211
rect 727 1202 731 1203
rect 727 1197 731 1198
rect 831 1202 835 1203
rect 831 1197 835 1198
rect 855 1202 859 1203
rect 855 1197 859 1198
rect 726 1196 732 1197
rect 726 1192 727 1196
rect 731 1192 732 1196
rect 726 1191 732 1192
rect 854 1196 860 1197
rect 854 1192 855 1196
rect 859 1192 860 1196
rect 854 1191 860 1192
rect 868 1168 870 1234
rect 983 1202 987 1203
rect 983 1197 987 1198
rect 982 1196 988 1197
rect 982 1192 983 1196
rect 987 1192 988 1196
rect 982 1191 988 1192
rect 1008 1168 1010 1234
rect 1014 1216 1020 1217
rect 1014 1212 1015 1216
rect 1019 1212 1020 1216
rect 1014 1211 1020 1212
rect 1206 1216 1212 1217
rect 1206 1212 1207 1216
rect 1211 1212 1212 1216
rect 1206 1211 1212 1212
rect 1016 1203 1018 1211
rect 1208 1203 1210 1211
rect 1015 1202 1019 1203
rect 1015 1197 1019 1198
rect 1103 1202 1107 1203
rect 1103 1197 1107 1198
rect 1207 1202 1211 1203
rect 1207 1197 1211 1198
rect 1223 1202 1227 1203
rect 1223 1197 1227 1198
rect 1102 1196 1108 1197
rect 1102 1192 1103 1196
rect 1107 1192 1108 1196
rect 1102 1191 1108 1192
rect 1222 1196 1228 1197
rect 1222 1192 1223 1196
rect 1227 1192 1228 1196
rect 1222 1191 1228 1192
rect 1232 1172 1234 1234
rect 1406 1216 1412 1217
rect 1406 1212 1407 1216
rect 1411 1212 1412 1216
rect 1406 1211 1412 1212
rect 1408 1203 1410 1211
rect 1335 1202 1339 1203
rect 1335 1197 1339 1198
rect 1407 1202 1411 1203
rect 1407 1197 1411 1198
rect 1447 1202 1451 1203
rect 1447 1197 1451 1198
rect 1334 1196 1340 1197
rect 1334 1192 1335 1196
rect 1339 1192 1340 1196
rect 1334 1191 1340 1192
rect 1446 1196 1452 1197
rect 1446 1192 1447 1196
rect 1451 1192 1452 1196
rect 1446 1191 1452 1192
rect 1230 1171 1236 1172
rect 726 1167 732 1168
rect 726 1163 727 1167
rect 731 1163 732 1167
rect 726 1162 732 1163
rect 734 1167 740 1168
rect 734 1163 735 1167
rect 739 1163 740 1167
rect 734 1162 740 1163
rect 854 1167 860 1168
rect 854 1163 855 1167
rect 859 1163 860 1167
rect 854 1162 860 1163
rect 866 1167 872 1168
rect 866 1163 867 1167
rect 871 1163 872 1167
rect 866 1162 872 1163
rect 982 1167 988 1168
rect 982 1163 983 1167
rect 987 1163 988 1167
rect 982 1162 988 1163
rect 1006 1167 1012 1168
rect 1006 1163 1007 1167
rect 1011 1163 1012 1167
rect 1006 1162 1012 1163
rect 1102 1167 1108 1168
rect 1102 1163 1103 1167
rect 1107 1163 1108 1167
rect 1102 1162 1108 1163
rect 1110 1167 1116 1168
rect 1110 1163 1111 1167
rect 1115 1163 1116 1167
rect 1110 1162 1116 1163
rect 1222 1167 1228 1168
rect 1222 1163 1223 1167
rect 1227 1163 1228 1167
rect 1230 1167 1231 1171
rect 1235 1167 1236 1171
rect 1230 1166 1236 1167
rect 1254 1171 1260 1172
rect 1254 1167 1255 1171
rect 1259 1167 1260 1171
rect 1456 1168 1458 1234
rect 1598 1216 1604 1217
rect 1608 1216 1610 1234
rect 1671 1233 1675 1234
rect 1695 1238 1699 1239
rect 1695 1233 1699 1234
rect 1672 1226 1674 1233
rect 1694 1232 1700 1233
rect 1694 1228 1695 1232
rect 1699 1228 1700 1232
rect 1694 1227 1700 1228
rect 1670 1225 1676 1226
rect 1630 1223 1636 1224
rect 1630 1219 1631 1223
rect 1635 1219 1636 1223
rect 1670 1221 1671 1225
rect 1675 1221 1676 1225
rect 1670 1220 1676 1221
rect 1630 1218 1636 1219
rect 1598 1212 1599 1216
rect 1603 1212 1604 1216
rect 1598 1211 1604 1212
rect 1606 1215 1612 1216
rect 1606 1211 1607 1215
rect 1611 1211 1612 1215
rect 1600 1203 1602 1211
rect 1606 1210 1612 1211
rect 1567 1202 1571 1203
rect 1567 1197 1571 1198
rect 1599 1202 1603 1203
rect 1599 1197 1603 1198
rect 1566 1196 1572 1197
rect 1566 1192 1567 1196
rect 1571 1192 1572 1196
rect 1566 1191 1572 1192
rect 1608 1172 1610 1210
rect 1632 1203 1634 1218
rect 1704 1216 1706 1278
rect 1790 1260 1796 1261
rect 1790 1256 1791 1260
rect 1795 1256 1796 1260
rect 1790 1255 1796 1256
rect 1934 1260 1940 1261
rect 1934 1256 1935 1260
rect 1939 1256 1940 1260
rect 1934 1255 1940 1256
rect 1792 1239 1794 1255
rect 1936 1239 1938 1255
rect 1791 1238 1795 1239
rect 1791 1233 1795 1234
rect 1935 1238 1939 1239
rect 1935 1233 1939 1234
rect 1702 1215 1708 1216
rect 1702 1211 1703 1215
rect 1707 1211 1708 1215
rect 1944 1212 1946 1282
rect 2718 1279 2719 1283
rect 2723 1279 2724 1283
rect 2982 1283 2983 1287
rect 2987 1283 2988 1287
rect 3158 1285 3159 1289
rect 3163 1285 3164 1289
rect 3168 1288 3170 1382
rect 3190 1381 3191 1385
rect 3195 1381 3196 1385
rect 3190 1380 3196 1381
rect 3190 1367 3196 1368
rect 3190 1363 3191 1367
rect 3195 1363 3196 1367
rect 3190 1362 3196 1363
rect 3192 1343 3194 1362
rect 3191 1342 3195 1343
rect 3191 1337 3195 1338
rect 3192 1330 3194 1337
rect 3190 1329 3196 1330
rect 3190 1325 3191 1329
rect 3195 1325 3196 1329
rect 3190 1324 3196 1325
rect 3190 1311 3196 1312
rect 3190 1307 3191 1311
rect 3195 1307 3196 1311
rect 3190 1306 3196 1307
rect 3192 1295 3194 1306
rect 3191 1294 3195 1295
rect 3191 1289 3195 1290
rect 3158 1284 3164 1285
rect 3166 1287 3172 1288
rect 2982 1282 2988 1283
rect 3166 1283 3167 1287
rect 3171 1283 3172 1287
rect 3192 1286 3194 1289
rect 3166 1282 3172 1283
rect 3190 1285 3196 1286
rect 2718 1278 2724 1279
rect 2102 1260 2108 1261
rect 2102 1256 2103 1260
rect 2107 1256 2108 1260
rect 2102 1255 2108 1256
rect 2294 1260 2300 1261
rect 2294 1256 2295 1260
rect 2299 1256 2300 1260
rect 2294 1255 2300 1256
rect 2494 1260 2500 1261
rect 2494 1256 2495 1260
rect 2499 1256 2500 1260
rect 2494 1255 2500 1256
rect 2710 1260 2716 1261
rect 2710 1256 2711 1260
rect 2715 1256 2716 1260
rect 2710 1255 2716 1256
rect 2104 1239 2106 1255
rect 2296 1239 2298 1255
rect 2496 1239 2498 1255
rect 2712 1239 2714 1255
rect 1983 1238 1987 1239
rect 1983 1233 1987 1234
rect 2103 1238 2107 1239
rect 2103 1233 2107 1234
rect 2255 1238 2259 1239
rect 2255 1233 2259 1234
rect 2295 1238 2299 1239
rect 2295 1233 2299 1234
rect 2495 1238 2499 1239
rect 2495 1233 2499 1234
rect 2711 1238 2715 1239
rect 2711 1233 2715 1234
rect 1982 1232 1988 1233
rect 1982 1228 1983 1232
rect 1987 1228 1988 1232
rect 1982 1227 1988 1228
rect 2254 1232 2260 1233
rect 2254 1228 2255 1232
rect 2259 1228 2260 1232
rect 2254 1227 2260 1228
rect 2494 1232 2500 1233
rect 2494 1228 2495 1232
rect 2499 1228 2500 1232
rect 2494 1227 2500 1228
rect 2710 1232 2716 1233
rect 2710 1228 2711 1232
rect 2715 1228 2716 1232
rect 2710 1227 2716 1228
rect 1702 1210 1708 1211
rect 1942 1211 1948 1212
rect 1670 1207 1676 1208
rect 1670 1203 1671 1207
rect 1675 1203 1676 1207
rect 1942 1207 1943 1211
rect 1947 1207 1948 1211
rect 1942 1206 1948 1207
rect 2720 1204 2722 1278
rect 2934 1260 2940 1261
rect 2934 1256 2935 1260
rect 2939 1256 2940 1260
rect 2934 1255 2940 1256
rect 3158 1260 3164 1261
rect 3158 1256 3159 1260
rect 3163 1256 3164 1260
rect 3158 1255 3164 1256
rect 2936 1239 2938 1255
rect 3160 1239 3162 1255
rect 2919 1238 2923 1239
rect 2919 1233 2923 1234
rect 2935 1238 2939 1239
rect 2935 1233 2939 1234
rect 3135 1238 3139 1239
rect 3135 1233 3139 1234
rect 3159 1238 3163 1239
rect 3159 1233 3163 1234
rect 2918 1232 2924 1233
rect 2918 1228 2919 1232
rect 2923 1228 2924 1232
rect 2918 1227 2924 1228
rect 3134 1232 3140 1233
rect 3134 1228 3135 1232
rect 3139 1228 3140 1232
rect 3134 1227 3140 1228
rect 3168 1208 3170 1282
rect 3190 1281 3191 1285
rect 3195 1281 3196 1285
rect 3190 1280 3196 1281
rect 3190 1267 3196 1268
rect 3190 1263 3191 1267
rect 3195 1263 3196 1267
rect 3190 1262 3196 1263
rect 3192 1239 3194 1262
rect 3191 1238 3195 1239
rect 3191 1233 3195 1234
rect 3192 1226 3194 1233
rect 3190 1225 3196 1226
rect 3190 1221 3191 1225
rect 3195 1221 3196 1225
rect 3190 1220 3196 1221
rect 3142 1207 3148 1208
rect 1631 1202 1635 1203
rect 1670 1202 1676 1203
rect 1694 1203 1700 1204
rect 1631 1197 1635 1198
rect 1632 1190 1634 1197
rect 1672 1195 1674 1202
rect 1694 1199 1695 1203
rect 1699 1199 1700 1203
rect 1694 1198 1700 1199
rect 1982 1203 1988 1204
rect 1982 1199 1983 1203
rect 1987 1199 1988 1203
rect 1982 1198 1988 1199
rect 2254 1203 2260 1204
rect 2254 1199 2255 1203
rect 2259 1199 2260 1203
rect 2254 1198 2260 1199
rect 2494 1203 2500 1204
rect 2494 1199 2495 1203
rect 2499 1199 2500 1203
rect 2494 1198 2500 1199
rect 2506 1203 2512 1204
rect 2506 1199 2507 1203
rect 2511 1199 2512 1203
rect 2506 1198 2512 1199
rect 2710 1203 2716 1204
rect 2710 1199 2711 1203
rect 2715 1199 2716 1203
rect 2710 1198 2716 1199
rect 2718 1203 2724 1204
rect 2718 1199 2719 1203
rect 2723 1199 2724 1203
rect 2718 1198 2724 1199
rect 2854 1203 2860 1204
rect 2854 1199 2855 1203
rect 2859 1199 2860 1203
rect 2854 1198 2860 1199
rect 2918 1203 2924 1204
rect 2918 1199 2919 1203
rect 2923 1199 2924 1203
rect 2918 1198 2924 1199
rect 3006 1203 3012 1204
rect 3006 1199 3007 1203
rect 3011 1199 3012 1203
rect 3006 1198 3012 1199
rect 3134 1203 3140 1204
rect 3134 1199 3135 1203
rect 3139 1199 3140 1203
rect 3142 1203 3143 1207
rect 3147 1203 3148 1207
rect 3142 1202 3148 1203
rect 3166 1207 3172 1208
rect 3166 1203 3167 1207
rect 3171 1203 3172 1207
rect 3166 1202 3172 1203
rect 3190 1207 3196 1208
rect 3190 1203 3191 1207
rect 3195 1203 3196 1207
rect 3190 1202 3196 1203
rect 3134 1198 3140 1199
rect 1696 1195 1698 1198
rect 1984 1195 1986 1198
rect 2182 1195 2188 1196
rect 2256 1195 2258 1198
rect 2496 1195 2498 1198
rect 1671 1194 1675 1195
rect 1630 1189 1636 1190
rect 1671 1189 1675 1190
rect 1695 1194 1699 1195
rect 1695 1189 1699 1190
rect 1983 1194 1987 1195
rect 2182 1191 2183 1195
rect 2187 1191 2188 1195
rect 2182 1190 2188 1191
rect 2247 1194 2251 1195
rect 2255 1194 2259 1195
rect 2399 1194 2403 1195
rect 2495 1194 2499 1195
rect 1983 1189 1987 1190
rect 1630 1185 1631 1189
rect 1635 1185 1636 1189
rect 1672 1186 1674 1189
rect 1630 1184 1636 1185
rect 1670 1185 1676 1186
rect 1670 1181 1671 1185
rect 1675 1181 1676 1185
rect 1670 1180 1676 1181
rect 1606 1171 1612 1172
rect 1254 1166 1260 1167
rect 1334 1167 1340 1168
rect 1222 1162 1228 1163
rect 728 1151 730 1162
rect 727 1150 731 1151
rect 727 1145 731 1146
rect 736 1140 738 1162
rect 856 1151 858 1162
rect 759 1150 763 1151
rect 855 1150 859 1151
rect 758 1145 764 1146
rect 855 1145 859 1146
rect 758 1141 759 1145
rect 763 1141 764 1145
rect 758 1140 764 1141
rect 868 1140 870 1162
rect 984 1151 986 1162
rect 879 1150 883 1151
rect 983 1150 987 1151
rect 999 1150 1003 1151
rect 878 1145 884 1146
rect 983 1145 987 1146
rect 998 1145 1004 1146
rect 878 1141 879 1145
rect 883 1141 884 1145
rect 878 1140 884 1141
rect 998 1141 999 1145
rect 1003 1141 1004 1145
rect 998 1140 1004 1141
rect 1008 1140 1010 1162
rect 1104 1151 1106 1162
rect 1103 1150 1107 1151
rect 1103 1145 1107 1146
rect 1112 1140 1114 1162
rect 1224 1151 1226 1162
rect 1119 1150 1123 1151
rect 1223 1150 1227 1151
rect 1231 1150 1235 1151
rect 1118 1145 1124 1146
rect 1223 1145 1227 1146
rect 1230 1145 1236 1146
rect 1118 1141 1119 1145
rect 1123 1141 1124 1145
rect 1118 1140 1124 1141
rect 1230 1141 1231 1145
rect 1235 1141 1236 1145
rect 1230 1140 1236 1141
rect 1256 1140 1258 1166
rect 1334 1163 1335 1167
rect 1339 1163 1340 1167
rect 1334 1162 1340 1163
rect 1343 1167 1349 1168
rect 1343 1163 1344 1167
rect 1348 1166 1349 1167
rect 1446 1167 1452 1168
rect 1348 1164 1354 1166
rect 1348 1163 1349 1164
rect 1343 1162 1349 1163
rect 1336 1151 1338 1162
rect 1335 1150 1339 1151
rect 1343 1150 1347 1151
rect 1335 1145 1339 1146
rect 1342 1145 1348 1146
rect 1342 1141 1343 1145
rect 1347 1141 1348 1145
rect 1342 1140 1348 1141
rect 1352 1140 1354 1164
rect 1446 1163 1447 1167
rect 1451 1163 1452 1167
rect 1446 1162 1452 1163
rect 1454 1167 1460 1168
rect 1454 1163 1455 1167
rect 1459 1163 1460 1167
rect 1454 1162 1460 1163
rect 1566 1167 1572 1168
rect 1566 1163 1567 1167
rect 1571 1163 1572 1167
rect 1606 1167 1607 1171
rect 1611 1167 1612 1171
rect 1606 1166 1612 1167
rect 1630 1171 1636 1172
rect 1630 1167 1631 1171
rect 1635 1167 1636 1171
rect 1630 1166 1636 1167
rect 1670 1167 1676 1168
rect 1566 1162 1572 1163
rect 1448 1151 1450 1162
rect 1447 1150 1451 1151
rect 1447 1145 1451 1146
rect 1456 1140 1458 1162
rect 1568 1151 1570 1162
rect 1632 1151 1634 1166
rect 1670 1163 1671 1167
rect 1675 1163 1676 1167
rect 1670 1162 1676 1163
rect 1672 1155 1674 1162
rect 1671 1154 1675 1155
rect 1463 1150 1467 1151
rect 1567 1150 1571 1151
rect 1462 1145 1468 1146
rect 1567 1145 1571 1146
rect 1631 1150 1635 1151
rect 1671 1149 1675 1150
rect 2175 1154 2179 1155
rect 2175 1149 2179 1150
rect 1631 1145 1635 1146
rect 1462 1141 1463 1145
rect 1467 1141 1468 1145
rect 1632 1142 1634 1145
rect 1672 1142 1674 1149
rect 2174 1148 2180 1149
rect 2174 1144 2175 1148
rect 2179 1144 2180 1148
rect 2174 1143 2180 1144
rect 1462 1140 1468 1141
rect 1630 1141 1636 1142
rect 638 1139 644 1140
rect 638 1135 639 1139
rect 643 1135 644 1139
rect 638 1134 644 1135
rect 670 1139 676 1140
rect 670 1135 671 1139
rect 675 1135 676 1139
rect 670 1134 676 1135
rect 734 1139 740 1140
rect 734 1135 735 1139
rect 739 1135 740 1139
rect 734 1134 740 1135
rect 782 1139 788 1140
rect 782 1135 783 1139
rect 787 1135 788 1139
rect 782 1134 788 1135
rect 866 1139 872 1140
rect 866 1135 867 1139
rect 871 1135 872 1139
rect 866 1134 872 1135
rect 906 1139 912 1140
rect 906 1135 907 1139
rect 911 1135 912 1139
rect 906 1134 912 1135
rect 1006 1139 1012 1140
rect 1006 1135 1007 1139
rect 1011 1135 1012 1139
rect 1006 1134 1012 1135
rect 1110 1139 1116 1140
rect 1110 1135 1111 1139
rect 1115 1135 1116 1139
rect 1110 1134 1116 1135
rect 1127 1139 1133 1140
rect 1127 1135 1128 1139
rect 1132 1138 1133 1139
rect 1254 1139 1260 1140
rect 1132 1136 1138 1138
rect 1132 1135 1133 1136
rect 1127 1134 1133 1135
rect 630 1116 636 1117
rect 630 1112 631 1116
rect 635 1112 636 1116
rect 630 1111 636 1112
rect 632 1099 634 1111
rect 527 1098 531 1099
rect 527 1093 531 1094
rect 631 1098 635 1099
rect 631 1093 635 1094
rect 526 1092 532 1093
rect 526 1088 527 1092
rect 531 1088 532 1092
rect 526 1087 532 1088
rect 526 1063 532 1064
rect 526 1059 527 1063
rect 531 1059 532 1063
rect 526 1058 532 1059
rect 534 1063 540 1064
rect 534 1059 535 1063
rect 539 1059 540 1063
rect 534 1058 540 1059
rect 528 1051 530 1058
rect 423 1050 427 1051
rect 527 1050 531 1051
rect 422 1045 428 1046
rect 527 1045 531 1046
rect 422 1041 423 1045
rect 427 1041 428 1045
rect 422 1040 428 1041
rect 536 1040 538 1058
rect 640 1056 642 1134
rect 758 1116 764 1117
rect 758 1112 759 1116
rect 763 1112 764 1116
rect 758 1111 764 1112
rect 760 1099 762 1111
rect 655 1098 659 1099
rect 655 1093 659 1094
rect 759 1098 763 1099
rect 759 1093 763 1094
rect 775 1098 779 1099
rect 775 1093 779 1094
rect 654 1092 660 1093
rect 654 1088 655 1092
rect 659 1088 660 1092
rect 654 1087 660 1088
rect 774 1092 780 1093
rect 774 1088 775 1092
rect 779 1088 780 1092
rect 774 1087 780 1088
rect 784 1068 786 1134
rect 878 1116 884 1117
rect 878 1112 879 1116
rect 883 1112 884 1116
rect 878 1111 884 1112
rect 880 1099 882 1111
rect 879 1098 883 1099
rect 879 1093 883 1094
rect 895 1098 899 1099
rect 895 1093 899 1094
rect 894 1092 900 1093
rect 894 1088 895 1092
rect 899 1088 900 1092
rect 894 1087 900 1088
rect 782 1067 788 1068
rect 654 1063 660 1064
rect 654 1059 655 1063
rect 659 1059 660 1063
rect 654 1058 660 1059
rect 774 1063 780 1064
rect 774 1059 775 1063
rect 779 1059 780 1063
rect 782 1063 783 1067
rect 787 1063 788 1067
rect 908 1064 910 1134
rect 998 1116 1004 1117
rect 998 1112 999 1116
rect 1003 1112 1004 1116
rect 998 1111 1004 1112
rect 1118 1116 1124 1117
rect 1118 1112 1119 1116
rect 1123 1112 1124 1116
rect 1118 1111 1124 1112
rect 1000 1099 1002 1111
rect 1120 1099 1122 1111
rect 999 1098 1003 1099
rect 999 1093 1003 1094
rect 1015 1098 1019 1099
rect 1015 1093 1019 1094
rect 1119 1098 1123 1099
rect 1119 1093 1123 1094
rect 1127 1098 1131 1099
rect 1127 1093 1131 1094
rect 1014 1092 1020 1093
rect 1014 1088 1015 1092
rect 1019 1088 1020 1092
rect 1014 1087 1020 1088
rect 1126 1092 1132 1093
rect 1126 1088 1127 1092
rect 1131 1088 1132 1092
rect 1126 1087 1132 1088
rect 1136 1064 1138 1136
rect 1254 1135 1255 1139
rect 1259 1135 1260 1139
rect 1254 1134 1260 1135
rect 1350 1139 1356 1140
rect 1350 1135 1351 1139
rect 1355 1135 1356 1139
rect 1350 1134 1356 1135
rect 1454 1139 1460 1140
rect 1454 1135 1455 1139
rect 1459 1135 1460 1139
rect 1630 1137 1631 1141
rect 1635 1137 1636 1141
rect 1630 1136 1636 1137
rect 1670 1141 1676 1142
rect 1670 1137 1671 1141
rect 1675 1137 1676 1141
rect 1670 1136 1676 1137
rect 1454 1134 1460 1135
rect 1230 1116 1236 1117
rect 1230 1112 1231 1116
rect 1235 1112 1236 1116
rect 1230 1111 1236 1112
rect 1232 1099 1234 1111
rect 1231 1098 1235 1099
rect 1231 1093 1235 1094
rect 1247 1098 1251 1099
rect 1247 1093 1251 1094
rect 1246 1092 1252 1093
rect 1246 1088 1247 1092
rect 1251 1088 1252 1092
rect 1246 1087 1252 1088
rect 1256 1064 1258 1134
rect 1630 1123 1636 1124
rect 1630 1119 1631 1123
rect 1635 1119 1636 1123
rect 1630 1118 1636 1119
rect 1670 1123 1676 1124
rect 1670 1119 1671 1123
rect 1675 1119 1676 1123
rect 2184 1120 2186 1190
rect 2246 1189 2252 1190
rect 2255 1189 2259 1190
rect 2398 1189 2404 1190
rect 2495 1189 2499 1190
rect 2246 1185 2247 1189
rect 2251 1185 2252 1189
rect 2246 1184 2252 1185
rect 2398 1185 2399 1189
rect 2403 1185 2404 1189
rect 2398 1184 2404 1185
rect 2508 1184 2510 1198
rect 2712 1195 2714 1198
rect 2551 1194 2555 1195
rect 2695 1194 2699 1195
rect 2711 1194 2715 1195
rect 2847 1194 2851 1195
rect 2550 1189 2556 1190
rect 2550 1185 2551 1189
rect 2555 1185 2556 1189
rect 2550 1184 2556 1185
rect 2694 1189 2700 1190
rect 2711 1189 2715 1190
rect 2846 1189 2852 1190
rect 2694 1185 2695 1189
rect 2699 1185 2700 1189
rect 2694 1184 2700 1185
rect 2702 1187 2708 1188
rect 2506 1183 2512 1184
rect 2506 1179 2507 1183
rect 2511 1179 2512 1183
rect 2702 1183 2703 1187
rect 2707 1183 2708 1187
rect 2846 1185 2847 1189
rect 2851 1185 2852 1189
rect 2856 1188 2858 1198
rect 2920 1195 2922 1198
rect 2919 1194 2923 1195
rect 2999 1194 3003 1195
rect 2919 1189 2923 1190
rect 2998 1189 3004 1190
rect 2846 1184 2852 1185
rect 2854 1187 2860 1188
rect 2702 1182 2708 1183
rect 2854 1183 2855 1187
rect 2859 1183 2860 1187
rect 2998 1185 2999 1189
rect 3003 1185 3004 1189
rect 2998 1184 3004 1185
rect 3008 1184 3010 1198
rect 3136 1195 3138 1198
rect 3135 1194 3139 1195
rect 3135 1189 3139 1190
rect 2854 1182 2860 1183
rect 3006 1183 3012 1184
rect 2506 1178 2512 1179
rect 2246 1160 2252 1161
rect 2246 1156 2247 1160
rect 2251 1156 2252 1160
rect 2246 1155 2252 1156
rect 2398 1160 2404 1161
rect 2398 1156 2399 1160
rect 2403 1156 2404 1160
rect 2398 1155 2404 1156
rect 2247 1154 2251 1155
rect 2247 1149 2251 1150
rect 2335 1154 2339 1155
rect 2335 1149 2339 1150
rect 2399 1154 2403 1155
rect 2399 1149 2403 1150
rect 2495 1154 2499 1155
rect 2495 1149 2499 1150
rect 2334 1148 2340 1149
rect 2334 1144 2335 1148
rect 2339 1144 2340 1148
rect 2334 1143 2340 1144
rect 2494 1148 2500 1149
rect 2494 1144 2495 1148
rect 2499 1144 2500 1148
rect 2494 1143 2500 1144
rect 2508 1124 2510 1178
rect 2550 1160 2556 1161
rect 2550 1156 2551 1160
rect 2555 1156 2556 1160
rect 2550 1155 2556 1156
rect 2694 1160 2700 1161
rect 2694 1156 2695 1160
rect 2699 1156 2700 1160
rect 2694 1155 2700 1156
rect 2551 1154 2555 1155
rect 2551 1149 2555 1150
rect 2655 1154 2659 1155
rect 2655 1149 2659 1150
rect 2695 1154 2699 1155
rect 2695 1149 2699 1150
rect 2654 1148 2660 1149
rect 2654 1144 2655 1148
rect 2659 1144 2660 1148
rect 2654 1143 2660 1144
rect 2704 1124 2706 1182
rect 2846 1160 2852 1161
rect 2846 1156 2847 1160
rect 2851 1156 2852 1160
rect 2846 1155 2852 1156
rect 2815 1154 2819 1155
rect 2815 1149 2819 1150
rect 2847 1154 2851 1155
rect 2847 1149 2851 1150
rect 2814 1148 2820 1149
rect 2814 1144 2815 1148
rect 2819 1144 2820 1148
rect 2814 1143 2820 1144
rect 2856 1124 2858 1182
rect 3006 1179 3007 1183
rect 3011 1179 3012 1183
rect 3006 1178 3012 1179
rect 2998 1160 3004 1161
rect 2998 1156 2999 1160
rect 3003 1156 3004 1160
rect 2998 1155 3004 1156
rect 2975 1154 2979 1155
rect 2975 1149 2979 1150
rect 2999 1154 3003 1155
rect 2999 1149 3003 1150
rect 2974 1148 2980 1149
rect 2974 1144 2975 1148
rect 2979 1144 2980 1148
rect 2974 1143 2980 1144
rect 3008 1124 3010 1178
rect 3135 1154 3139 1155
rect 3135 1149 3139 1150
rect 3134 1148 3140 1149
rect 3134 1144 3135 1148
rect 3139 1144 3140 1148
rect 3134 1143 3140 1144
rect 3144 1124 3146 1202
rect 3192 1195 3194 1202
rect 3191 1194 3195 1195
rect 3191 1189 3195 1190
rect 3192 1186 3194 1189
rect 3190 1185 3196 1186
rect 3190 1181 3191 1185
rect 3195 1181 3196 1185
rect 3190 1180 3196 1181
rect 3190 1167 3196 1168
rect 3190 1163 3191 1167
rect 3195 1163 3196 1167
rect 3190 1162 3196 1163
rect 3192 1155 3194 1162
rect 3191 1154 3195 1155
rect 3191 1149 3195 1150
rect 3192 1142 3194 1149
rect 3190 1141 3196 1142
rect 3190 1137 3191 1141
rect 3195 1137 3196 1141
rect 3190 1136 3196 1137
rect 2506 1123 2512 1124
rect 1670 1118 1676 1119
rect 2174 1119 2180 1120
rect 1342 1116 1348 1117
rect 1342 1112 1343 1116
rect 1347 1112 1348 1116
rect 1342 1111 1348 1112
rect 1462 1116 1468 1117
rect 1462 1112 1463 1116
rect 1467 1112 1468 1116
rect 1462 1111 1468 1112
rect 1344 1099 1346 1111
rect 1464 1099 1466 1111
rect 1632 1099 1634 1118
rect 1672 1111 1674 1118
rect 2174 1115 2175 1119
rect 2179 1115 2180 1119
rect 2174 1114 2180 1115
rect 2182 1119 2188 1120
rect 2182 1115 2183 1119
rect 2187 1115 2188 1119
rect 2182 1114 2188 1115
rect 2334 1119 2340 1120
rect 2334 1115 2335 1119
rect 2339 1115 2340 1119
rect 2334 1114 2340 1115
rect 2494 1119 2500 1120
rect 2494 1115 2495 1119
rect 2499 1115 2500 1119
rect 2506 1119 2507 1123
rect 2511 1119 2512 1123
rect 2662 1123 2668 1124
rect 2506 1118 2512 1119
rect 2654 1119 2660 1120
rect 2494 1114 2500 1115
rect 2176 1111 2178 1114
rect 1671 1110 1675 1111
rect 2071 1110 2075 1111
rect 2175 1110 2179 1111
rect 1671 1105 1675 1106
rect 2070 1105 2076 1106
rect 2175 1105 2179 1106
rect 1672 1102 1674 1105
rect 1670 1101 1676 1102
rect 1343 1098 1347 1099
rect 1343 1093 1347 1094
rect 1367 1098 1371 1099
rect 1367 1093 1371 1094
rect 1463 1098 1467 1099
rect 1463 1093 1467 1094
rect 1631 1098 1635 1099
rect 1670 1097 1671 1101
rect 1675 1097 1676 1101
rect 2070 1101 2071 1105
rect 2075 1101 2076 1105
rect 2070 1100 2076 1101
rect 2184 1100 2186 1114
rect 2336 1111 2338 1114
rect 2496 1111 2498 1114
rect 2191 1110 2195 1111
rect 2327 1110 2331 1111
rect 2335 1110 2339 1111
rect 2479 1110 2483 1111
rect 2495 1110 2499 1111
rect 2190 1105 2196 1106
rect 2190 1101 2191 1105
rect 2195 1101 2196 1105
rect 2190 1100 2196 1101
rect 2326 1105 2332 1106
rect 2335 1105 2339 1106
rect 2478 1105 2484 1106
rect 2495 1105 2499 1106
rect 2326 1101 2327 1105
rect 2331 1101 2332 1105
rect 2326 1100 2332 1101
rect 2350 1103 2356 1104
rect 1670 1096 1676 1097
rect 2078 1099 2084 1100
rect 2078 1095 2079 1099
rect 2083 1095 2084 1099
rect 2078 1094 2084 1095
rect 2182 1099 2188 1100
rect 2182 1095 2183 1099
rect 2187 1095 2188 1099
rect 2350 1099 2351 1103
rect 2355 1099 2356 1103
rect 2478 1101 2479 1105
rect 2483 1101 2484 1105
rect 2508 1104 2510 1118
rect 2654 1115 2655 1119
rect 2659 1115 2660 1119
rect 2662 1119 2663 1123
rect 2667 1119 2668 1123
rect 2662 1118 2668 1119
rect 2702 1123 2708 1124
rect 2702 1119 2703 1123
rect 2707 1119 2708 1123
rect 2822 1123 2828 1124
rect 2702 1118 2708 1119
rect 2814 1119 2820 1120
rect 2654 1114 2660 1115
rect 2656 1111 2658 1114
rect 2639 1110 2643 1111
rect 2655 1110 2659 1111
rect 2638 1105 2644 1106
rect 2655 1105 2659 1106
rect 2478 1100 2484 1101
rect 2506 1103 2512 1104
rect 2350 1098 2356 1099
rect 2506 1099 2507 1103
rect 2511 1099 2512 1103
rect 2638 1101 2639 1105
rect 2643 1101 2644 1105
rect 2664 1104 2666 1118
rect 2814 1115 2815 1119
rect 2819 1115 2820 1119
rect 2822 1119 2823 1123
rect 2827 1119 2828 1123
rect 2822 1118 2828 1119
rect 2854 1123 2860 1124
rect 2854 1119 2855 1123
rect 2859 1119 2860 1123
rect 3006 1123 3012 1124
rect 2854 1118 2860 1119
rect 2974 1119 2980 1120
rect 2814 1114 2820 1115
rect 2816 1111 2818 1114
rect 2815 1110 2819 1111
rect 2814 1105 2820 1106
rect 2638 1100 2644 1101
rect 2662 1103 2668 1104
rect 2506 1098 2512 1099
rect 2662 1099 2663 1103
rect 2667 1099 2668 1103
rect 2814 1101 2815 1105
rect 2819 1101 2820 1105
rect 2824 1104 2826 1118
rect 2974 1115 2975 1119
rect 2979 1115 2980 1119
rect 3006 1119 3007 1123
rect 3011 1119 3012 1123
rect 3142 1123 3148 1124
rect 3006 1118 3012 1119
rect 3134 1119 3140 1120
rect 2974 1114 2980 1115
rect 2976 1111 2978 1114
rect 2975 1110 2979 1111
rect 2999 1110 3003 1111
rect 2975 1105 2979 1106
rect 2998 1105 3004 1106
rect 2814 1100 2820 1101
rect 2822 1103 2828 1104
rect 2662 1098 2668 1099
rect 2822 1099 2823 1103
rect 2827 1099 2828 1103
rect 2998 1101 2999 1105
rect 3003 1101 3004 1105
rect 2998 1100 3004 1101
rect 3008 1100 3010 1118
rect 3134 1115 3135 1119
rect 3139 1115 3140 1119
rect 3142 1119 3143 1123
rect 3147 1119 3148 1123
rect 3142 1118 3148 1119
rect 3190 1123 3196 1124
rect 3190 1119 3191 1123
rect 3195 1119 3196 1123
rect 3190 1118 3196 1119
rect 3134 1114 3140 1115
rect 3136 1111 3138 1114
rect 3135 1110 3139 1111
rect 3135 1105 3139 1106
rect 3144 1100 3146 1118
rect 3192 1111 3194 1118
rect 3159 1110 3163 1111
rect 3191 1110 3195 1111
rect 3158 1105 3164 1106
rect 3191 1105 3195 1106
rect 3158 1101 3159 1105
rect 3163 1101 3164 1105
rect 3192 1102 3194 1105
rect 3158 1100 3164 1101
rect 3190 1101 3196 1102
rect 2822 1098 2828 1099
rect 3006 1099 3012 1100
rect 2182 1094 2188 1095
rect 1631 1093 1635 1094
rect 1366 1092 1372 1093
rect 1366 1088 1367 1092
rect 1371 1088 1372 1092
rect 1366 1087 1372 1088
rect 1632 1086 1634 1093
rect 1630 1085 1636 1086
rect 1630 1081 1631 1085
rect 1635 1081 1636 1085
rect 1630 1080 1636 1081
rect 1670 1083 1676 1084
rect 1670 1079 1671 1083
rect 1675 1079 1676 1083
rect 1670 1078 1676 1079
rect 1630 1067 1636 1068
rect 782 1062 788 1063
rect 894 1063 900 1064
rect 774 1058 780 1059
rect 582 1055 588 1056
rect 582 1051 583 1055
rect 587 1051 588 1055
rect 551 1050 555 1051
rect 582 1050 588 1051
rect 638 1055 644 1056
rect 638 1051 639 1055
rect 643 1051 644 1055
rect 656 1051 658 1058
rect 776 1051 778 1058
rect 638 1050 644 1051
rect 655 1050 659 1051
rect 550 1045 556 1046
rect 550 1041 551 1045
rect 555 1041 556 1045
rect 550 1040 556 1041
rect 584 1040 586 1050
rect 679 1050 683 1051
rect 775 1050 779 1051
rect 655 1045 659 1046
rect 678 1045 684 1046
rect 775 1045 779 1046
rect 678 1041 679 1045
rect 683 1041 684 1045
rect 678 1040 684 1041
rect 702 1043 708 1044
rect 462 1039 468 1040
rect 462 1035 463 1039
rect 467 1035 468 1039
rect 462 1034 468 1035
rect 534 1039 540 1040
rect 534 1035 535 1039
rect 539 1035 540 1039
rect 534 1034 540 1035
rect 582 1039 588 1040
rect 582 1035 583 1039
rect 587 1035 588 1039
rect 702 1039 703 1043
rect 707 1039 708 1043
rect 784 1040 786 1062
rect 894 1059 895 1063
rect 899 1059 900 1063
rect 894 1058 900 1059
rect 906 1063 912 1064
rect 906 1059 907 1063
rect 911 1059 912 1063
rect 906 1058 912 1059
rect 1014 1063 1020 1064
rect 1014 1059 1015 1063
rect 1019 1059 1020 1063
rect 1014 1058 1020 1059
rect 1038 1063 1044 1064
rect 1038 1059 1039 1063
rect 1043 1059 1044 1063
rect 1038 1058 1044 1059
rect 1126 1063 1132 1064
rect 1126 1059 1127 1063
rect 1131 1059 1132 1063
rect 1126 1058 1132 1059
rect 1134 1063 1140 1064
rect 1134 1059 1135 1063
rect 1139 1059 1140 1063
rect 1134 1058 1140 1059
rect 1246 1063 1252 1064
rect 1246 1059 1247 1063
rect 1251 1059 1252 1063
rect 1246 1058 1252 1059
rect 1254 1063 1260 1064
rect 1254 1059 1255 1063
rect 1259 1059 1260 1063
rect 1254 1058 1260 1059
rect 1366 1063 1372 1064
rect 1366 1059 1367 1063
rect 1371 1059 1372 1063
rect 1630 1063 1631 1067
rect 1635 1063 1636 1067
rect 1630 1062 1636 1063
rect 1366 1058 1372 1059
rect 896 1051 898 1058
rect 799 1050 803 1051
rect 895 1050 899 1051
rect 798 1045 804 1046
rect 895 1045 899 1046
rect 798 1041 799 1045
rect 803 1041 804 1045
rect 798 1040 804 1041
rect 908 1040 910 1058
rect 1016 1051 1018 1058
rect 919 1050 923 1051
rect 1015 1050 1019 1051
rect 1031 1050 1035 1051
rect 918 1045 924 1046
rect 1015 1045 1019 1046
rect 1030 1045 1036 1046
rect 918 1041 919 1045
rect 923 1041 924 1045
rect 918 1040 924 1041
rect 1030 1041 1031 1045
rect 1035 1041 1036 1045
rect 1030 1040 1036 1041
rect 1040 1040 1042 1058
rect 1128 1051 1130 1058
rect 1127 1050 1131 1051
rect 1127 1045 1131 1046
rect 1136 1040 1138 1058
rect 1248 1051 1250 1058
rect 1143 1050 1147 1051
rect 1247 1050 1251 1051
rect 1142 1045 1148 1046
rect 1247 1045 1251 1046
rect 1142 1041 1143 1045
rect 1147 1041 1148 1045
rect 1142 1040 1148 1041
rect 1256 1040 1258 1058
rect 1368 1051 1370 1058
rect 1632 1051 1634 1062
rect 1672 1059 1674 1078
rect 2070 1076 2076 1077
rect 2070 1072 2071 1076
rect 2075 1072 2076 1076
rect 2070 1071 2076 1072
rect 2072 1059 2074 1071
rect 1671 1058 1675 1059
rect 1671 1053 1675 1054
rect 1975 1058 1979 1059
rect 1975 1053 1979 1054
rect 2071 1058 2075 1059
rect 2071 1053 2075 1054
rect 1263 1050 1267 1051
rect 1367 1050 1371 1051
rect 1262 1045 1268 1046
rect 1367 1045 1371 1046
rect 1631 1050 1635 1051
rect 1672 1046 1674 1053
rect 1974 1052 1980 1053
rect 1974 1048 1975 1052
rect 1979 1048 1980 1052
rect 1974 1047 1980 1048
rect 1631 1045 1635 1046
rect 1670 1045 1676 1046
rect 1262 1041 1263 1045
rect 1267 1041 1268 1045
rect 1632 1042 1634 1045
rect 1262 1040 1268 1041
rect 1630 1041 1636 1042
rect 702 1038 708 1039
rect 782 1039 788 1040
rect 582 1034 588 1035
rect 422 1016 428 1017
rect 422 1012 423 1016
rect 427 1012 428 1016
rect 422 1011 428 1012
rect 424 999 426 1011
rect 327 998 331 999
rect 327 993 331 994
rect 423 998 427 999
rect 423 993 427 994
rect 455 998 459 999
rect 455 993 459 994
rect 326 992 332 993
rect 326 988 327 992
rect 331 988 332 992
rect 326 987 332 988
rect 454 992 460 993
rect 454 988 455 992
rect 459 988 460 992
rect 454 987 460 988
rect 464 964 466 1034
rect 550 1016 556 1017
rect 550 1012 551 1016
rect 555 1012 556 1016
rect 550 1011 556 1012
rect 552 999 554 1011
rect 551 998 555 999
rect 551 993 555 994
rect 575 998 579 999
rect 575 993 579 994
rect 574 992 580 993
rect 574 988 575 992
rect 579 988 580 992
rect 574 987 580 988
rect 584 968 586 1034
rect 678 1016 684 1017
rect 678 1012 679 1016
rect 683 1012 684 1016
rect 678 1011 684 1012
rect 680 999 682 1011
rect 679 998 683 999
rect 679 993 683 994
rect 695 998 699 999
rect 695 993 699 994
rect 694 992 700 993
rect 694 988 695 992
rect 699 988 700 992
rect 694 987 700 988
rect 704 968 706 1038
rect 782 1035 783 1039
rect 787 1035 788 1039
rect 782 1034 788 1035
rect 906 1039 912 1040
rect 906 1035 907 1039
rect 911 1035 912 1039
rect 906 1034 912 1035
rect 1038 1039 1044 1040
rect 1038 1035 1039 1039
rect 1043 1035 1044 1039
rect 1038 1034 1044 1035
rect 1134 1039 1140 1040
rect 1134 1035 1135 1039
rect 1139 1035 1140 1039
rect 1134 1034 1140 1035
rect 1166 1039 1172 1040
rect 1166 1035 1167 1039
rect 1171 1035 1172 1039
rect 1166 1034 1172 1035
rect 1254 1039 1260 1040
rect 1254 1035 1255 1039
rect 1259 1035 1260 1039
rect 1630 1037 1631 1041
rect 1635 1037 1636 1041
rect 1670 1041 1671 1045
rect 1675 1041 1676 1045
rect 1670 1040 1676 1041
rect 1630 1036 1636 1037
rect 1254 1034 1260 1035
rect 798 1016 804 1017
rect 798 1012 799 1016
rect 803 1012 804 1016
rect 798 1011 804 1012
rect 918 1016 924 1017
rect 918 1012 919 1016
rect 923 1012 924 1016
rect 918 1011 924 1012
rect 1030 1016 1036 1017
rect 1030 1012 1031 1016
rect 1035 1012 1036 1016
rect 1030 1011 1036 1012
rect 1142 1016 1148 1017
rect 1142 1012 1143 1016
rect 1147 1012 1148 1016
rect 1142 1011 1148 1012
rect 800 999 802 1011
rect 920 999 922 1011
rect 1032 999 1034 1011
rect 1144 999 1146 1011
rect 799 998 803 999
rect 799 993 803 994
rect 815 998 819 999
rect 815 993 819 994
rect 919 998 923 999
rect 919 993 923 994
rect 927 998 931 999
rect 927 993 931 994
rect 1031 998 1035 999
rect 1031 993 1035 994
rect 1039 998 1043 999
rect 1039 993 1043 994
rect 1143 998 1147 999
rect 1143 993 1147 994
rect 1159 998 1163 999
rect 1159 993 1163 994
rect 814 992 820 993
rect 814 988 815 992
rect 819 988 820 992
rect 814 987 820 988
rect 926 992 932 993
rect 926 988 927 992
rect 931 988 932 992
rect 926 987 932 988
rect 1038 992 1044 993
rect 1038 988 1039 992
rect 1043 988 1044 992
rect 1038 987 1044 988
rect 1158 992 1164 993
rect 1158 988 1159 992
rect 1163 988 1164 992
rect 1158 987 1164 988
rect 582 967 588 968
rect 326 963 332 964
rect 326 959 327 963
rect 331 959 332 963
rect 326 958 332 959
rect 334 963 340 964
rect 334 959 335 963
rect 339 959 340 963
rect 334 958 340 959
rect 454 963 460 964
rect 454 959 455 963
rect 459 959 460 963
rect 454 958 460 959
rect 462 963 468 964
rect 462 959 463 963
rect 467 959 468 963
rect 462 958 468 959
rect 574 963 580 964
rect 574 959 575 963
rect 579 959 580 963
rect 582 963 583 967
rect 587 963 588 967
rect 702 967 708 968
rect 582 962 588 963
rect 694 963 700 964
rect 574 958 580 959
rect 328 947 330 958
rect 327 946 331 947
rect 327 941 331 942
rect 336 940 338 958
rect 456 947 458 958
rect 351 946 355 947
rect 455 946 459 947
rect 350 941 356 942
rect 455 941 459 942
rect 222 936 228 937
rect 258 939 264 940
rect 258 935 259 939
rect 263 935 264 939
rect 258 934 264 935
rect 334 939 340 940
rect 334 935 335 939
rect 339 935 340 939
rect 350 937 351 941
rect 355 937 356 941
rect 350 936 356 937
rect 464 936 466 958
rect 576 947 578 958
rect 471 946 475 947
rect 575 946 579 947
rect 470 941 476 942
rect 575 941 579 942
rect 470 937 471 941
rect 475 937 476 941
rect 470 936 476 937
rect 584 936 586 962
rect 694 959 695 963
rect 699 959 700 963
rect 702 963 703 967
rect 707 963 708 967
rect 1168 964 1170 1034
rect 1670 1027 1676 1028
rect 1630 1023 1636 1024
rect 1630 1019 1631 1023
rect 1635 1019 1636 1023
rect 1670 1023 1671 1027
rect 1675 1023 1676 1027
rect 1670 1022 1676 1023
rect 1974 1023 1980 1024
rect 1630 1018 1636 1019
rect 1262 1016 1268 1017
rect 1262 1012 1263 1016
rect 1267 1012 1268 1016
rect 1262 1011 1268 1012
rect 1264 999 1266 1011
rect 1632 999 1634 1018
rect 1672 1015 1674 1022
rect 1974 1019 1975 1023
rect 1979 1019 1980 1023
rect 1974 1018 1980 1019
rect 1926 1015 1932 1016
rect 1976 1015 1978 1018
rect 2080 1016 2082 1094
rect 2190 1076 2196 1077
rect 2190 1072 2191 1076
rect 2195 1072 2196 1076
rect 2190 1071 2196 1072
rect 2326 1076 2332 1077
rect 2326 1072 2327 1076
rect 2331 1072 2332 1076
rect 2326 1071 2332 1072
rect 2192 1059 2194 1071
rect 2328 1059 2330 1071
rect 2095 1058 2099 1059
rect 2095 1053 2099 1054
rect 2191 1058 2195 1059
rect 2191 1053 2195 1054
rect 2215 1058 2219 1059
rect 2215 1053 2219 1054
rect 2327 1058 2331 1059
rect 2327 1053 2331 1054
rect 2343 1058 2347 1059
rect 2343 1053 2347 1054
rect 2094 1052 2100 1053
rect 2094 1048 2095 1052
rect 2099 1048 2100 1052
rect 2094 1047 2100 1048
rect 2214 1052 2220 1053
rect 2214 1048 2215 1052
rect 2219 1048 2220 1052
rect 2214 1047 2220 1048
rect 2342 1052 2348 1053
rect 2342 1048 2343 1052
rect 2347 1048 2348 1052
rect 2342 1047 2348 1048
rect 2352 1028 2354 1098
rect 3006 1095 3007 1099
rect 3011 1095 3012 1099
rect 3006 1094 3012 1095
rect 3142 1099 3148 1100
rect 3142 1095 3143 1099
rect 3147 1095 3148 1099
rect 3142 1094 3148 1095
rect 3166 1099 3172 1100
rect 3166 1095 3167 1099
rect 3171 1095 3172 1099
rect 3190 1097 3191 1101
rect 3195 1097 3196 1101
rect 3190 1096 3196 1097
rect 3166 1094 3172 1095
rect 2478 1076 2484 1077
rect 2478 1072 2479 1076
rect 2483 1072 2484 1076
rect 2478 1071 2484 1072
rect 2638 1076 2644 1077
rect 2638 1072 2639 1076
rect 2643 1072 2644 1076
rect 2638 1071 2644 1072
rect 2814 1076 2820 1077
rect 2814 1072 2815 1076
rect 2819 1072 2820 1076
rect 2814 1071 2820 1072
rect 2998 1076 3004 1077
rect 2998 1072 2999 1076
rect 3003 1072 3004 1076
rect 2998 1071 3004 1072
rect 2480 1059 2482 1071
rect 2640 1059 2642 1071
rect 2816 1059 2818 1071
rect 3000 1059 3002 1071
rect 2479 1058 2483 1059
rect 2479 1053 2483 1054
rect 2487 1058 2491 1059
rect 2487 1053 2491 1054
rect 2639 1058 2643 1059
rect 2639 1053 2643 1054
rect 2647 1058 2651 1059
rect 2647 1053 2651 1054
rect 2815 1058 2819 1059
rect 2815 1053 2819 1054
rect 2823 1058 2827 1059
rect 2823 1053 2827 1054
rect 2999 1058 3003 1059
rect 2999 1053 3003 1054
rect 2486 1052 2492 1053
rect 2486 1048 2487 1052
rect 2491 1048 2492 1052
rect 2486 1047 2492 1048
rect 2646 1052 2652 1053
rect 2646 1048 2647 1052
rect 2651 1048 2652 1052
rect 2646 1047 2652 1048
rect 2822 1052 2828 1053
rect 2822 1048 2823 1052
rect 2827 1048 2828 1052
rect 2822 1047 2828 1048
rect 2998 1052 3004 1053
rect 2998 1048 2999 1052
rect 3003 1048 3004 1052
rect 2998 1047 3004 1048
rect 3008 1032 3010 1094
rect 3158 1076 3164 1077
rect 3158 1072 3159 1076
rect 3163 1072 3164 1076
rect 3158 1071 3164 1072
rect 3160 1059 3162 1071
rect 3159 1058 3163 1059
rect 3159 1053 3163 1054
rect 3158 1052 3164 1053
rect 3158 1048 3159 1052
rect 3163 1048 3164 1052
rect 3158 1047 3164 1048
rect 3006 1031 3012 1032
rect 2350 1027 2356 1028
rect 2094 1023 2100 1024
rect 2094 1019 2095 1023
rect 2099 1019 2100 1023
rect 2094 1018 2100 1019
rect 2214 1023 2220 1024
rect 2214 1019 2215 1023
rect 2219 1019 2220 1023
rect 2214 1018 2220 1019
rect 2342 1023 2348 1024
rect 2342 1019 2343 1023
rect 2347 1019 2348 1023
rect 2350 1023 2351 1027
rect 2355 1023 2356 1027
rect 2830 1027 2836 1028
rect 2350 1022 2356 1023
rect 2486 1023 2492 1024
rect 2342 1018 2348 1019
rect 2078 1015 2084 1016
rect 2096 1015 2098 1018
rect 2216 1015 2218 1018
rect 2230 1015 2236 1016
rect 2344 1015 2346 1018
rect 1671 1014 1675 1015
rect 1895 1014 1899 1015
rect 1926 1011 1927 1015
rect 1931 1011 1932 1015
rect 1926 1010 1932 1011
rect 1975 1014 1979 1015
rect 2047 1014 2051 1015
rect 2078 1011 2079 1015
rect 2083 1011 2084 1015
rect 2078 1010 2084 1011
rect 2095 1014 2099 1015
rect 2199 1014 2203 1015
rect 2215 1014 2219 1015
rect 2230 1011 2231 1015
rect 2235 1011 2236 1015
rect 2230 1010 2236 1011
rect 2343 1014 2347 1015
rect 1671 1009 1675 1010
rect 1894 1009 1900 1010
rect 1672 1006 1674 1009
rect 1670 1005 1676 1006
rect 1670 1001 1671 1005
rect 1675 1001 1676 1005
rect 1894 1005 1895 1009
rect 1899 1005 1900 1009
rect 1894 1004 1900 1005
rect 1928 1004 1930 1010
rect 1975 1009 1979 1010
rect 2046 1009 2052 1010
rect 2095 1009 2099 1010
rect 2198 1009 2204 1010
rect 2215 1009 2219 1010
rect 2046 1005 2047 1009
rect 2051 1005 2052 1009
rect 2046 1004 2052 1005
rect 2198 1005 2199 1009
rect 2203 1005 2204 1009
rect 2198 1004 2204 1005
rect 1670 1000 1676 1001
rect 1926 1003 1932 1004
rect 1926 999 1927 1003
rect 1931 999 1932 1003
rect 1263 998 1267 999
rect 1263 993 1267 994
rect 1631 998 1635 999
rect 1926 998 1932 999
rect 1631 993 1635 994
rect 1632 986 1634 993
rect 1670 987 1676 988
rect 1630 985 1636 986
rect 1630 981 1631 985
rect 1635 981 1636 985
rect 1670 983 1671 987
rect 1675 983 1676 987
rect 1670 982 1676 983
rect 1630 980 1636 981
rect 1672 975 1674 982
rect 1894 980 1900 981
rect 1894 976 1895 980
rect 1899 976 1900 980
rect 1894 975 1900 976
rect 1671 974 1675 975
rect 1671 969 1675 970
rect 1791 974 1795 975
rect 1791 969 1795 970
rect 1895 974 1899 975
rect 1895 969 1899 970
rect 1919 974 1923 975
rect 1919 969 1923 970
rect 1630 967 1636 968
rect 702 962 708 963
rect 814 963 820 964
rect 694 958 700 959
rect 696 947 698 958
rect 591 946 595 947
rect 695 946 699 947
rect 590 941 596 942
rect 695 941 699 942
rect 590 937 591 941
rect 595 937 596 941
rect 590 936 596 937
rect 704 936 706 962
rect 814 959 815 963
rect 819 959 820 963
rect 814 958 820 959
rect 823 963 829 964
rect 823 959 824 963
rect 828 962 829 963
rect 926 963 932 964
rect 828 960 834 962
rect 828 959 829 960
rect 823 958 829 959
rect 816 947 818 958
rect 711 946 715 947
rect 815 946 819 947
rect 823 946 827 947
rect 710 941 716 942
rect 815 941 819 942
rect 822 941 828 942
rect 710 937 711 941
rect 715 937 716 941
rect 710 936 716 937
rect 822 937 823 941
rect 827 937 828 941
rect 822 936 828 937
rect 832 936 834 960
rect 926 959 927 963
rect 931 959 932 963
rect 926 958 932 959
rect 950 963 956 964
rect 950 959 951 963
rect 955 959 956 963
rect 950 958 956 959
rect 1038 963 1044 964
rect 1038 959 1039 963
rect 1043 959 1044 963
rect 1038 958 1044 959
rect 1070 963 1076 964
rect 1070 959 1071 963
rect 1075 959 1076 963
rect 1070 958 1076 959
rect 1158 963 1164 964
rect 1158 959 1159 963
rect 1163 959 1164 963
rect 1158 958 1164 959
rect 1166 963 1172 964
rect 1166 959 1167 963
rect 1171 959 1172 963
rect 1630 963 1631 967
rect 1635 963 1636 967
rect 1630 962 1636 963
rect 1672 962 1674 969
rect 1790 968 1796 969
rect 1790 964 1791 968
rect 1795 964 1796 968
rect 1790 963 1796 964
rect 1918 968 1924 969
rect 1918 964 1919 968
rect 1923 964 1924 968
rect 1918 963 1924 964
rect 1166 958 1172 959
rect 928 947 930 958
rect 927 946 931 947
rect 943 946 947 947
rect 927 941 931 942
rect 942 941 948 942
rect 942 937 943 941
rect 947 937 948 941
rect 942 936 948 937
rect 952 936 954 958
rect 1040 947 1042 958
rect 1039 946 1043 947
rect 1063 946 1067 947
rect 1039 941 1043 942
rect 1062 941 1068 942
rect 1062 937 1063 941
rect 1067 937 1068 941
rect 1062 936 1068 937
rect 1072 936 1074 958
rect 1160 947 1162 958
rect 1159 946 1163 947
rect 1159 941 1163 942
rect 334 934 340 935
rect 462 935 468 936
rect 110 932 116 933
rect 110 919 116 920
rect 110 915 111 919
rect 115 915 116 919
rect 110 914 116 915
rect 112 895 114 914
rect 222 912 228 913
rect 222 908 223 912
rect 227 908 228 912
rect 222 907 228 908
rect 224 895 226 907
rect 111 894 115 895
rect 111 889 115 890
rect 135 894 139 895
rect 135 889 139 890
rect 223 894 227 895
rect 223 889 227 890
rect 247 894 251 895
rect 247 889 251 890
rect 112 882 114 889
rect 134 888 140 889
rect 134 884 135 888
rect 139 884 140 888
rect 134 883 140 884
rect 246 888 252 889
rect 246 884 247 888
rect 251 884 252 888
rect 246 883 252 884
rect 110 881 116 882
rect 110 877 111 881
rect 115 877 116 881
rect 110 876 116 877
rect 260 864 262 934
rect 462 931 463 935
rect 467 931 468 935
rect 462 930 468 931
rect 582 935 588 936
rect 582 931 583 935
rect 587 931 588 935
rect 582 930 588 931
rect 702 935 708 936
rect 702 931 703 935
rect 707 931 708 935
rect 702 930 708 931
rect 830 935 836 936
rect 830 931 831 935
rect 835 931 836 935
rect 830 930 836 931
rect 950 935 956 936
rect 950 931 951 935
rect 955 931 956 935
rect 950 930 956 931
rect 1070 935 1076 936
rect 1070 931 1071 935
rect 1075 931 1076 935
rect 1070 930 1076 931
rect 350 912 356 913
rect 350 908 351 912
rect 355 908 356 912
rect 350 907 356 908
rect 470 912 476 913
rect 470 908 471 912
rect 475 908 476 912
rect 470 907 476 908
rect 590 912 596 913
rect 590 908 591 912
rect 595 908 596 912
rect 590 907 596 908
rect 710 912 716 913
rect 710 908 711 912
rect 715 908 716 912
rect 710 907 716 908
rect 822 912 828 913
rect 822 908 823 912
rect 827 908 828 912
rect 822 907 828 908
rect 942 912 948 913
rect 942 908 943 912
rect 947 908 948 912
rect 942 907 948 908
rect 1062 912 1068 913
rect 1062 908 1063 912
rect 1067 908 1068 912
rect 1062 907 1068 908
rect 352 895 354 907
rect 472 895 474 907
rect 592 895 594 907
rect 712 895 714 907
rect 824 895 826 907
rect 944 895 946 907
rect 1064 895 1066 907
rect 351 894 355 895
rect 351 889 355 890
rect 383 894 387 895
rect 383 889 387 890
rect 471 894 475 895
rect 471 889 475 890
rect 535 894 539 895
rect 535 889 539 890
rect 591 894 595 895
rect 591 889 595 890
rect 711 894 715 895
rect 711 889 715 890
rect 823 894 827 895
rect 823 889 827 890
rect 919 894 923 895
rect 919 889 923 890
rect 943 894 947 895
rect 943 889 947 890
rect 1063 894 1067 895
rect 1063 889 1067 890
rect 382 888 388 889
rect 382 884 383 888
rect 387 884 388 888
rect 382 883 388 884
rect 534 888 540 889
rect 534 884 535 888
rect 539 884 540 888
rect 534 883 540 884
rect 710 888 716 889
rect 710 884 711 888
rect 715 884 716 888
rect 710 883 716 884
rect 918 888 924 889
rect 918 884 919 888
rect 923 884 924 888
rect 918 883 924 884
rect 110 863 116 864
rect 110 859 111 863
rect 115 859 116 863
rect 258 863 264 864
rect 110 858 116 859
rect 134 859 140 860
rect 112 851 114 858
rect 134 855 135 859
rect 139 855 140 859
rect 134 854 140 855
rect 246 859 252 860
rect 246 855 247 859
rect 251 855 252 859
rect 258 859 259 863
rect 263 859 264 863
rect 258 858 264 859
rect 382 859 388 860
rect 246 854 252 855
rect 136 851 138 854
rect 248 851 250 854
rect 260 852 262 858
rect 382 855 383 859
rect 387 855 388 859
rect 382 854 388 855
rect 534 859 540 860
rect 534 855 535 859
rect 539 855 540 859
rect 534 854 540 855
rect 710 859 716 860
rect 710 855 711 859
rect 715 855 716 859
rect 710 854 716 855
rect 718 859 724 860
rect 718 855 719 859
rect 723 855 724 859
rect 718 854 724 855
rect 918 859 924 860
rect 918 855 919 859
rect 923 855 924 859
rect 918 854 924 855
rect 926 859 932 860
rect 926 855 927 859
rect 931 855 932 859
rect 926 854 932 855
rect 258 851 264 852
rect 384 851 386 854
rect 536 851 538 854
rect 582 851 588 852
rect 712 851 714 854
rect 111 850 115 851
rect 135 850 139 851
rect 247 850 251 851
rect 258 847 259 851
rect 263 847 264 851
rect 258 846 264 847
rect 303 850 307 851
rect 383 850 387 851
rect 503 850 507 851
rect 535 850 539 851
rect 582 847 583 851
rect 587 847 588 851
rect 582 846 588 847
rect 695 850 699 851
rect 711 850 715 851
rect 111 845 115 846
rect 134 845 140 846
rect 247 845 251 846
rect 302 845 308 846
rect 383 845 387 846
rect 502 845 508 846
rect 535 845 539 846
rect 112 842 114 845
rect 110 841 116 842
rect 110 837 111 841
rect 115 837 116 841
rect 134 841 135 845
rect 139 841 140 845
rect 134 840 140 841
rect 302 841 303 845
rect 307 841 308 845
rect 302 840 308 841
rect 502 841 503 845
rect 507 841 508 845
rect 502 840 508 841
rect 110 836 116 837
rect 110 823 116 824
rect 110 819 111 823
rect 115 819 116 823
rect 110 818 116 819
rect 112 795 114 818
rect 134 816 140 817
rect 134 812 135 816
rect 139 812 140 816
rect 134 811 140 812
rect 302 816 308 817
rect 302 812 303 816
rect 307 812 308 816
rect 302 811 308 812
rect 502 816 508 817
rect 502 812 503 816
rect 507 812 508 816
rect 502 811 508 812
rect 136 795 138 811
rect 304 795 306 811
rect 504 795 506 811
rect 111 794 115 795
rect 111 789 115 790
rect 135 794 139 795
rect 135 789 139 790
rect 303 794 307 795
rect 303 789 307 790
rect 503 794 507 795
rect 503 789 507 790
rect 112 782 114 789
rect 110 781 116 782
rect 110 777 111 781
rect 115 777 116 781
rect 110 776 116 777
rect 110 763 116 764
rect 110 759 111 763
rect 115 759 116 763
rect 110 758 116 759
rect 112 747 114 758
rect 111 746 115 747
rect 575 746 579 747
rect 111 741 115 742
rect 574 741 580 742
rect 112 738 114 741
rect 110 737 116 738
rect 110 733 111 737
rect 115 733 116 737
rect 574 737 575 741
rect 579 737 580 741
rect 574 736 580 737
rect 584 736 586 846
rect 694 845 700 846
rect 711 845 715 846
rect 694 841 695 845
rect 699 841 700 845
rect 694 840 700 841
rect 720 840 722 854
rect 920 851 922 854
rect 879 850 883 851
rect 919 850 923 851
rect 878 845 884 846
rect 919 845 923 846
rect 878 841 879 845
rect 883 841 884 845
rect 878 840 884 841
rect 928 840 930 854
rect 1047 850 1051 851
rect 1046 845 1052 846
rect 1046 841 1047 845
rect 1051 841 1052 845
rect 1046 840 1052 841
rect 1072 840 1074 930
rect 1143 894 1147 895
rect 1143 889 1147 890
rect 1142 888 1148 889
rect 1142 884 1143 888
rect 1147 884 1148 888
rect 1142 883 1148 884
rect 1168 860 1170 958
rect 1632 947 1634 962
rect 1670 961 1676 962
rect 1670 957 1671 961
rect 1675 957 1676 961
rect 1670 956 1676 957
rect 1631 946 1635 947
rect 1631 941 1635 942
rect 1670 943 1676 944
rect 1632 938 1634 941
rect 1670 939 1671 943
rect 1675 939 1676 943
rect 1928 940 1930 998
rect 2046 980 2052 981
rect 2046 976 2047 980
rect 2051 976 2052 980
rect 2046 975 2052 976
rect 2198 980 2204 981
rect 2198 976 2199 980
rect 2203 976 2204 980
rect 2198 975 2204 976
rect 2047 974 2051 975
rect 2047 969 2051 970
rect 2071 974 2075 975
rect 2071 969 2075 970
rect 2199 974 2203 975
rect 2199 969 2203 970
rect 2070 968 2076 969
rect 2070 964 2071 968
rect 2075 964 2076 968
rect 2070 963 2076 964
rect 2232 948 2234 1010
rect 2342 1009 2348 1010
rect 2342 1005 2343 1009
rect 2347 1005 2348 1009
rect 2352 1008 2354 1022
rect 2486 1019 2487 1023
rect 2491 1019 2492 1023
rect 2486 1018 2492 1019
rect 2646 1023 2652 1024
rect 2646 1019 2647 1023
rect 2651 1019 2652 1023
rect 2646 1018 2652 1019
rect 2654 1023 2660 1024
rect 2654 1019 2655 1023
rect 2659 1019 2660 1023
rect 2654 1018 2660 1019
rect 2822 1023 2828 1024
rect 2822 1019 2823 1023
rect 2827 1019 2828 1023
rect 2830 1023 2831 1027
rect 2835 1023 2836 1027
rect 3006 1027 3007 1031
rect 3011 1027 3012 1031
rect 3168 1028 3170 1094
rect 3190 1083 3196 1084
rect 3190 1079 3191 1083
rect 3195 1079 3196 1083
rect 3190 1078 3196 1079
rect 3192 1059 3194 1078
rect 3191 1058 3195 1059
rect 3191 1053 3195 1054
rect 3192 1046 3194 1053
rect 3190 1045 3196 1046
rect 3190 1041 3191 1045
rect 3195 1041 3196 1045
rect 3190 1040 3196 1041
rect 3006 1026 3012 1027
rect 3166 1027 3172 1028
rect 2830 1022 2836 1023
rect 2998 1023 3004 1024
rect 2822 1018 2828 1019
rect 2488 1015 2490 1018
rect 2648 1015 2650 1018
rect 2487 1014 2491 1015
rect 2495 1014 2499 1015
rect 2647 1014 2651 1015
rect 2487 1009 2491 1010
rect 2494 1009 2500 1010
rect 2342 1004 2348 1005
rect 2350 1007 2356 1008
rect 2350 1003 2351 1007
rect 2355 1003 2356 1007
rect 2494 1005 2495 1009
rect 2499 1005 2500 1009
rect 2494 1004 2500 1005
rect 2646 1009 2652 1010
rect 2646 1005 2647 1009
rect 2651 1005 2652 1009
rect 2646 1004 2652 1005
rect 2656 1004 2658 1018
rect 2824 1015 2826 1018
rect 2823 1014 2827 1015
rect 2823 1009 2827 1010
rect 2350 1002 2356 1003
rect 2654 1003 2660 1004
rect 2654 999 2655 1003
rect 2659 999 2660 1003
rect 2654 998 2660 999
rect 2702 1003 2708 1004
rect 2702 999 2703 1003
rect 2707 999 2708 1003
rect 2702 998 2708 999
rect 2342 980 2348 981
rect 2342 976 2343 980
rect 2347 976 2348 980
rect 2342 975 2348 976
rect 2494 980 2500 981
rect 2494 976 2495 980
rect 2499 976 2500 980
rect 2494 975 2500 976
rect 2646 980 2652 981
rect 2646 976 2647 980
rect 2651 976 2652 980
rect 2646 975 2652 976
rect 2255 974 2259 975
rect 2255 969 2259 970
rect 2343 974 2347 975
rect 2343 969 2347 970
rect 2463 974 2467 975
rect 2463 969 2467 970
rect 2495 974 2499 975
rect 2495 969 2499 970
rect 2647 974 2651 975
rect 2647 969 2651 970
rect 2695 974 2699 975
rect 2695 969 2699 970
rect 2254 968 2260 969
rect 2254 964 2255 968
rect 2259 964 2260 968
rect 2254 963 2260 964
rect 2462 968 2468 969
rect 2462 964 2463 968
rect 2467 964 2468 968
rect 2462 963 2468 964
rect 2694 968 2700 969
rect 2694 964 2695 968
rect 2699 964 2700 968
rect 2694 963 2700 964
rect 2230 947 2236 948
rect 2230 943 2231 947
rect 2235 943 2236 947
rect 2704 944 2706 998
rect 2832 944 2834 1022
rect 2998 1019 2999 1023
rect 3003 1019 3004 1023
rect 2998 1018 3004 1019
rect 3000 1015 3002 1018
rect 2999 1014 3003 1015
rect 2999 1009 3003 1010
rect 2935 974 2939 975
rect 2935 969 2939 970
rect 2934 968 2940 969
rect 2934 964 2935 968
rect 2939 964 2940 968
rect 2934 963 2940 964
rect 3008 944 3010 1026
rect 3158 1023 3164 1024
rect 3158 1019 3159 1023
rect 3163 1019 3164 1023
rect 3166 1023 3167 1027
rect 3171 1023 3172 1027
rect 3166 1022 3172 1023
rect 3190 1027 3196 1028
rect 3190 1023 3191 1027
rect 3195 1023 3196 1027
rect 3190 1022 3196 1023
rect 3158 1018 3164 1019
rect 3160 1015 3162 1018
rect 3159 1014 3163 1015
rect 3159 1009 3163 1010
rect 3159 974 3163 975
rect 3159 969 3163 970
rect 3158 968 3164 969
rect 3158 964 3159 968
rect 3163 964 3164 968
rect 3158 963 3164 964
rect 3168 944 3170 1022
rect 3192 1015 3194 1022
rect 3191 1014 3195 1015
rect 3191 1009 3195 1010
rect 3192 1006 3194 1009
rect 3190 1005 3196 1006
rect 3190 1001 3191 1005
rect 3195 1001 3196 1005
rect 3190 1000 3196 1001
rect 3190 987 3196 988
rect 3190 983 3191 987
rect 3195 983 3196 987
rect 3190 982 3196 983
rect 3192 975 3194 982
rect 3191 974 3195 975
rect 3191 969 3195 970
rect 3192 962 3194 969
rect 3190 961 3196 962
rect 3190 957 3191 961
rect 3195 957 3196 961
rect 3190 956 3196 957
rect 2230 942 2236 943
rect 2702 943 2708 944
rect 1670 938 1676 939
rect 1790 939 1796 940
rect 1630 937 1636 938
rect 1630 933 1631 937
rect 1635 933 1636 937
rect 1630 932 1636 933
rect 1672 927 1674 938
rect 1790 935 1791 939
rect 1795 935 1796 939
rect 1790 934 1796 935
rect 1802 939 1808 940
rect 1802 935 1803 939
rect 1807 935 1808 939
rect 1802 934 1808 935
rect 1918 939 1924 940
rect 1918 935 1919 939
rect 1923 935 1924 939
rect 1918 934 1924 935
rect 1926 939 1932 940
rect 1926 935 1927 939
rect 1931 935 1932 939
rect 1926 934 1932 935
rect 2070 939 2076 940
rect 2070 935 2071 939
rect 2075 935 2076 939
rect 2070 934 2076 935
rect 2078 939 2084 940
rect 2078 935 2079 939
rect 2083 935 2084 939
rect 2078 934 2084 935
rect 1792 927 1794 934
rect 1671 926 1675 927
rect 1719 926 1723 927
rect 1791 926 1795 927
rect 1671 921 1675 922
rect 1718 921 1724 922
rect 1791 921 1795 922
rect 1630 919 1636 920
rect 1630 915 1631 919
rect 1635 915 1636 919
rect 1672 918 1674 921
rect 1630 914 1636 915
rect 1670 917 1676 918
rect 1632 895 1634 914
rect 1670 913 1671 917
rect 1675 913 1676 917
rect 1718 917 1719 921
rect 1723 917 1724 921
rect 1718 916 1724 917
rect 1804 916 1806 934
rect 1920 927 1922 934
rect 1871 926 1875 927
rect 1919 926 1923 927
rect 1870 921 1876 922
rect 1919 921 1923 922
rect 1870 917 1871 921
rect 1875 917 1876 921
rect 1870 916 1876 917
rect 1928 916 1930 934
rect 2072 927 2074 934
rect 2039 926 2043 927
rect 2071 926 2075 927
rect 2038 921 2044 922
rect 2071 921 2075 922
rect 2038 917 2039 921
rect 2043 917 2044 921
rect 2038 916 2044 917
rect 2080 916 2082 934
rect 2223 926 2227 927
rect 2222 921 2228 922
rect 2222 917 2223 921
rect 2227 917 2228 921
rect 2232 920 2234 942
rect 2254 939 2260 940
rect 2254 935 2255 939
rect 2259 935 2260 939
rect 2254 934 2260 935
rect 2462 939 2468 940
rect 2462 935 2463 939
rect 2467 935 2468 939
rect 2462 934 2468 935
rect 2470 939 2476 940
rect 2470 935 2471 939
rect 2475 935 2476 939
rect 2470 934 2476 935
rect 2694 939 2700 940
rect 2694 935 2695 939
rect 2699 935 2700 939
rect 2702 939 2703 943
rect 2707 939 2708 943
rect 2702 938 2708 939
rect 2830 943 2836 944
rect 2830 939 2831 943
rect 2835 939 2836 943
rect 2942 943 2948 944
rect 2830 938 2836 939
rect 2934 939 2940 940
rect 2694 934 2700 935
rect 2256 927 2258 934
rect 2464 927 2466 934
rect 2255 926 2259 927
rect 2439 926 2443 927
rect 2463 926 2467 927
rect 2255 921 2259 922
rect 2438 921 2444 922
rect 2463 921 2467 922
rect 2222 916 2228 917
rect 2230 919 2236 920
rect 1670 912 1676 913
rect 1802 915 1808 916
rect 1802 911 1803 915
rect 1807 911 1808 915
rect 1802 910 1808 911
rect 1926 915 1932 916
rect 1926 911 1927 915
rect 1931 911 1932 915
rect 1926 910 1932 911
rect 2022 915 2028 916
rect 2022 911 2023 915
rect 2027 911 2028 915
rect 2022 910 2028 911
rect 2078 915 2084 916
rect 2078 911 2079 915
rect 2083 911 2084 915
rect 2230 915 2231 919
rect 2235 915 2236 919
rect 2438 917 2439 921
rect 2443 917 2444 921
rect 2472 920 2474 934
rect 2696 927 2698 934
rect 2671 926 2675 927
rect 2695 926 2699 927
rect 2670 921 2676 922
rect 2695 921 2699 922
rect 2438 916 2444 917
rect 2446 919 2452 920
rect 2230 914 2236 915
rect 2446 915 2447 919
rect 2451 915 2452 919
rect 2446 914 2452 915
rect 2470 919 2476 920
rect 2470 915 2471 919
rect 2475 915 2476 919
rect 2670 917 2671 921
rect 2675 917 2676 921
rect 2704 920 2706 938
rect 2934 935 2935 939
rect 2939 935 2940 939
rect 2942 939 2943 943
rect 2947 939 2948 943
rect 2942 938 2948 939
rect 3006 943 3012 944
rect 3006 939 3007 943
rect 3011 939 3012 943
rect 3166 943 3172 944
rect 3006 938 3012 939
rect 3158 939 3164 940
rect 2934 934 2940 935
rect 2936 927 2938 934
rect 2911 926 2915 927
rect 2935 926 2939 927
rect 2910 921 2916 922
rect 2935 921 2939 922
rect 2670 916 2676 917
rect 2702 919 2708 920
rect 2470 914 2476 915
rect 2702 915 2703 919
rect 2707 915 2708 919
rect 2910 917 2911 921
rect 2915 917 2916 921
rect 2944 920 2946 938
rect 3158 935 3159 939
rect 3163 935 3164 939
rect 3166 939 3167 943
rect 3171 939 3172 943
rect 3166 938 3172 939
rect 3190 943 3196 944
rect 3190 939 3191 943
rect 3195 939 3196 943
rect 3190 938 3196 939
rect 3158 934 3164 935
rect 3160 927 3162 934
rect 3159 926 3163 927
rect 3158 921 3164 922
rect 2910 916 2916 917
rect 2942 919 2948 920
rect 2702 914 2708 915
rect 2942 915 2943 919
rect 2947 915 2948 919
rect 3158 917 3159 921
rect 3163 917 3164 921
rect 3168 920 3170 938
rect 3192 927 3194 938
rect 3191 926 3195 927
rect 3191 921 3195 922
rect 3158 916 3164 917
rect 3166 919 3172 920
rect 2942 914 2948 915
rect 3166 915 3167 919
rect 3171 915 3172 919
rect 3192 918 3194 921
rect 3166 914 3172 915
rect 3190 917 3196 918
rect 2078 910 2084 911
rect 1670 899 1676 900
rect 1670 895 1671 899
rect 1675 895 1676 899
rect 1383 894 1387 895
rect 1383 889 1387 890
rect 1599 894 1603 895
rect 1599 889 1603 890
rect 1631 894 1635 895
rect 1670 894 1676 895
rect 1631 889 1635 890
rect 1382 888 1388 889
rect 1382 884 1383 888
rect 1387 884 1388 888
rect 1382 883 1388 884
rect 1598 888 1604 889
rect 1598 884 1599 888
rect 1603 884 1604 888
rect 1598 883 1604 884
rect 1632 882 1634 889
rect 1672 887 1674 894
rect 1718 892 1724 893
rect 1718 888 1719 892
rect 1723 888 1724 892
rect 1718 887 1724 888
rect 1870 892 1876 893
rect 1870 888 1871 892
rect 1875 888 1876 892
rect 1870 887 1876 888
rect 1671 886 1675 887
rect 1630 881 1636 882
rect 1671 881 1675 882
rect 1695 886 1699 887
rect 1695 881 1699 882
rect 1719 886 1723 887
rect 1719 881 1723 882
rect 1871 886 1875 887
rect 1871 881 1875 882
rect 2015 886 2019 887
rect 2015 881 2019 882
rect 1630 877 1631 881
rect 1635 877 1636 881
rect 1630 876 1636 877
rect 1672 874 1674 881
rect 1694 880 1700 881
rect 1694 876 1695 880
rect 1699 876 1700 880
rect 1694 875 1700 876
rect 2014 880 2020 881
rect 2014 876 2015 880
rect 2019 876 2020 880
rect 2014 875 2020 876
rect 1670 873 1676 874
rect 1670 869 1671 873
rect 1675 869 1676 873
rect 1670 868 1676 869
rect 1630 863 1636 864
rect 1142 859 1148 860
rect 1142 855 1143 859
rect 1147 855 1148 859
rect 1142 854 1148 855
rect 1154 859 1160 860
rect 1154 855 1155 859
rect 1159 855 1160 859
rect 1154 854 1160 855
rect 1166 859 1172 860
rect 1166 855 1167 859
rect 1171 855 1172 859
rect 1166 854 1172 855
rect 1382 859 1388 860
rect 1382 855 1383 859
rect 1387 855 1388 859
rect 1382 854 1388 855
rect 1394 859 1400 860
rect 1394 855 1395 859
rect 1399 855 1400 859
rect 1394 854 1400 855
rect 1598 859 1604 860
rect 1598 855 1599 859
rect 1603 855 1604 859
rect 1630 859 1631 863
rect 1635 859 1636 863
rect 1630 858 1636 859
rect 1598 854 1604 855
rect 1144 851 1146 854
rect 1143 850 1147 851
rect 1143 845 1147 846
rect 1156 840 1158 854
rect 1384 851 1386 854
rect 1199 850 1203 851
rect 1335 850 1339 851
rect 1383 850 1387 851
rect 1198 845 1204 846
rect 1198 841 1199 845
rect 1203 841 1204 845
rect 1198 840 1204 841
rect 1334 845 1340 846
rect 1383 845 1387 846
rect 1334 841 1335 845
rect 1339 841 1340 845
rect 1334 840 1340 841
rect 1396 840 1398 854
rect 1600 851 1602 854
rect 1632 851 1634 858
rect 2024 856 2026 910
rect 2038 892 2044 893
rect 2038 888 2039 892
rect 2043 888 2044 892
rect 2038 887 2044 888
rect 2222 892 2228 893
rect 2222 888 2223 892
rect 2227 888 2228 892
rect 2222 887 2228 888
rect 2039 886 2043 887
rect 2039 881 2043 882
rect 2223 886 2227 887
rect 2223 881 2227 882
rect 1670 855 1676 856
rect 1670 851 1671 855
rect 1675 851 1676 855
rect 2022 855 2028 856
rect 1471 850 1475 851
rect 1599 850 1603 851
rect 1631 850 1635 851
rect 1670 850 1676 851
rect 1694 851 1700 852
rect 1470 845 1476 846
rect 1470 841 1471 845
rect 1475 841 1476 845
rect 1470 840 1476 841
rect 1598 845 1604 846
rect 1631 845 1635 846
rect 1598 841 1599 845
rect 1603 841 1604 845
rect 1632 842 1634 845
rect 1598 840 1604 841
rect 1630 841 1636 842
rect 686 839 692 840
rect 686 835 687 839
rect 691 835 692 839
rect 686 834 692 835
rect 718 839 724 840
rect 718 835 719 839
rect 723 835 724 839
rect 718 834 724 835
rect 886 839 892 840
rect 886 835 887 839
rect 891 835 892 839
rect 886 834 892 835
rect 926 839 932 840
rect 926 835 927 839
rect 931 835 932 839
rect 926 834 932 835
rect 1070 839 1076 840
rect 1070 835 1071 839
rect 1075 835 1076 839
rect 1070 834 1076 835
rect 1154 839 1160 840
rect 1154 835 1155 839
rect 1159 835 1160 839
rect 1154 834 1160 835
rect 1394 839 1400 840
rect 1394 835 1395 839
rect 1399 835 1400 839
rect 1394 834 1400 835
rect 1526 839 1532 840
rect 1526 835 1527 839
rect 1531 835 1532 839
rect 1630 837 1631 841
rect 1635 837 1636 841
rect 1630 836 1636 837
rect 1672 835 1674 850
rect 1694 847 1695 851
rect 1699 847 1700 851
rect 1694 846 1700 847
rect 2014 851 2020 852
rect 2014 847 2015 851
rect 2019 847 2020 851
rect 2022 851 2023 855
rect 2027 851 2028 855
rect 2022 850 2028 851
rect 2014 846 2020 847
rect 1696 835 1698 846
rect 2016 835 2018 846
rect 1526 834 1532 835
rect 1671 834 1675 835
rect 679 794 683 795
rect 679 789 683 790
rect 678 788 684 789
rect 678 784 679 788
rect 683 784 684 788
rect 678 783 684 784
rect 688 760 690 834
rect 694 816 700 817
rect 694 812 695 816
rect 699 812 700 816
rect 694 811 700 812
rect 878 816 884 817
rect 878 812 879 816
rect 883 812 884 816
rect 878 811 884 812
rect 696 795 698 811
rect 880 795 882 811
rect 695 794 699 795
rect 695 789 699 790
rect 807 794 811 795
rect 807 789 811 790
rect 879 794 883 795
rect 879 789 883 790
rect 806 788 812 789
rect 806 784 807 788
rect 811 784 812 788
rect 806 783 812 784
rect 678 759 684 760
rect 678 755 679 759
rect 683 755 684 759
rect 678 754 684 755
rect 686 759 692 760
rect 686 755 687 759
rect 691 755 692 759
rect 686 754 692 755
rect 806 759 812 760
rect 806 755 807 759
rect 811 755 812 759
rect 806 754 812 755
rect 814 759 820 760
rect 814 755 815 759
rect 819 755 820 759
rect 814 754 820 755
rect 614 751 620 752
rect 614 747 615 751
rect 619 747 620 751
rect 680 747 682 754
rect 808 747 810 754
rect 614 746 620 747
rect 679 746 683 747
rect 616 736 618 746
rect 703 746 707 747
rect 807 746 811 747
rect 679 741 683 742
rect 702 741 708 742
rect 807 741 811 742
rect 702 737 703 741
rect 707 737 708 741
rect 702 736 708 737
rect 816 736 818 754
rect 831 746 835 747
rect 830 741 836 742
rect 830 737 831 741
rect 835 737 836 741
rect 830 736 836 737
rect 888 736 890 834
rect 1046 816 1052 817
rect 1046 812 1047 816
rect 1051 812 1052 816
rect 1046 811 1052 812
rect 1198 816 1204 817
rect 1198 812 1199 816
rect 1203 812 1204 816
rect 1198 811 1204 812
rect 1334 816 1340 817
rect 1334 812 1335 816
rect 1339 812 1340 816
rect 1334 811 1340 812
rect 1470 816 1476 817
rect 1470 812 1471 816
rect 1475 812 1476 816
rect 1470 811 1476 812
rect 1048 795 1050 811
rect 1200 795 1202 811
rect 1336 795 1338 811
rect 1472 795 1474 811
rect 927 794 931 795
rect 927 789 931 790
rect 1047 794 1051 795
rect 1047 789 1051 790
rect 1167 794 1171 795
rect 1167 789 1171 790
rect 1199 794 1203 795
rect 1199 789 1203 790
rect 1279 794 1283 795
rect 1279 789 1283 790
rect 1335 794 1339 795
rect 1335 789 1339 790
rect 1399 794 1403 795
rect 1399 789 1403 790
rect 1471 794 1475 795
rect 1471 789 1475 790
rect 1519 794 1523 795
rect 1519 789 1523 790
rect 926 788 932 789
rect 926 784 927 788
rect 931 784 932 788
rect 926 783 932 784
rect 1046 788 1052 789
rect 1046 784 1047 788
rect 1051 784 1052 788
rect 1046 783 1052 784
rect 1166 788 1172 789
rect 1166 784 1167 788
rect 1171 784 1172 788
rect 1166 783 1172 784
rect 1278 788 1284 789
rect 1278 784 1279 788
rect 1283 784 1284 788
rect 1278 783 1284 784
rect 1398 788 1404 789
rect 1398 784 1399 788
rect 1403 784 1404 788
rect 1398 783 1404 784
rect 1518 788 1524 789
rect 1518 784 1519 788
rect 1523 784 1524 788
rect 1518 783 1524 784
rect 1422 767 1428 768
rect 1422 763 1423 767
rect 1427 763 1428 767
rect 1528 764 1530 834
rect 1671 829 1675 830
rect 1695 834 1699 835
rect 1695 829 1699 830
rect 2015 834 2019 835
rect 2015 829 2019 830
rect 1672 826 1674 829
rect 1670 825 1676 826
rect 1630 823 1636 824
rect 1630 819 1631 823
rect 1635 819 1636 823
rect 1670 821 1671 825
rect 1675 821 1676 825
rect 2232 824 2234 914
rect 2438 892 2444 893
rect 2438 888 2439 892
rect 2443 888 2444 892
rect 2438 887 2444 888
rect 2367 886 2371 887
rect 2367 881 2371 882
rect 2439 886 2443 887
rect 2439 881 2443 882
rect 2366 880 2372 881
rect 2366 876 2367 880
rect 2371 876 2372 880
rect 2366 875 2372 876
rect 2448 856 2450 914
rect 2670 892 2676 893
rect 2670 888 2671 892
rect 2675 888 2676 892
rect 2670 887 2676 888
rect 2910 892 2916 893
rect 2910 888 2911 892
rect 2915 888 2916 892
rect 2910 887 2916 888
rect 3158 892 3164 893
rect 3158 888 3159 892
rect 3163 888 3164 892
rect 3158 887 3164 888
rect 2671 886 2675 887
rect 2671 881 2675 882
rect 2727 886 2731 887
rect 2727 881 2731 882
rect 2911 886 2915 887
rect 2911 881 2915 882
rect 3087 886 3091 887
rect 3087 881 3091 882
rect 3159 886 3163 887
rect 3159 881 3163 882
rect 2726 880 2732 881
rect 2726 876 2727 880
rect 2731 876 2732 880
rect 2726 875 2732 876
rect 3086 880 3092 881
rect 3086 876 3087 880
rect 3091 876 3092 880
rect 3086 875 3092 876
rect 3168 856 3170 914
rect 3190 913 3191 917
rect 3195 913 3196 917
rect 3190 912 3196 913
rect 3190 899 3196 900
rect 3190 895 3191 899
rect 3195 895 3196 899
rect 3190 894 3196 895
rect 3192 887 3194 894
rect 3191 886 3195 887
rect 3191 881 3195 882
rect 3192 874 3194 881
rect 3190 873 3196 874
rect 3190 869 3191 873
rect 3195 869 3196 873
rect 3190 868 3196 869
rect 2446 855 2452 856
rect 2366 851 2372 852
rect 2366 847 2367 851
rect 2371 847 2372 851
rect 2446 851 2447 855
rect 2451 851 2452 855
rect 3118 855 3124 856
rect 2446 850 2452 851
rect 2726 851 2732 852
rect 2366 846 2372 847
rect 2368 835 2370 846
rect 2279 834 2283 835
rect 2367 834 2371 835
rect 2439 834 2443 835
rect 2278 829 2284 830
rect 2367 829 2371 830
rect 2438 829 2444 830
rect 2278 825 2279 829
rect 2283 825 2284 829
rect 2278 824 2284 825
rect 2438 825 2439 829
rect 2443 825 2444 829
rect 2448 828 2450 850
rect 2726 847 2727 851
rect 2731 847 2732 851
rect 2726 846 2732 847
rect 2738 851 2744 852
rect 2738 847 2739 851
rect 2743 847 2744 851
rect 2738 846 2744 847
rect 3086 851 3092 852
rect 3086 847 3087 851
rect 3091 847 3092 851
rect 3118 851 3119 855
rect 3123 851 3124 855
rect 3118 850 3124 851
rect 3166 855 3172 856
rect 3166 851 3167 855
rect 3171 851 3172 855
rect 3166 850 3172 851
rect 3190 855 3196 856
rect 3190 851 3191 855
rect 3195 851 3196 855
rect 3190 850 3196 851
rect 3086 846 3092 847
rect 2728 835 2730 846
rect 2583 834 2587 835
rect 2719 834 2723 835
rect 2727 834 2731 835
rect 2582 829 2588 830
rect 2438 824 2444 825
rect 2446 827 2452 828
rect 1670 820 1676 821
rect 2230 823 2236 824
rect 1630 818 1636 819
rect 2230 819 2231 823
rect 2235 819 2236 823
rect 2230 818 2236 819
rect 2306 823 2312 824
rect 2306 819 2307 823
rect 2311 819 2312 823
rect 2446 823 2447 827
rect 2451 823 2452 827
rect 2446 822 2452 823
rect 2458 827 2464 828
rect 2458 823 2459 827
rect 2463 823 2464 827
rect 2582 825 2583 829
rect 2587 825 2588 829
rect 2582 824 2588 825
rect 2718 829 2724 830
rect 2727 829 2731 830
rect 2718 825 2719 829
rect 2723 825 2724 829
rect 2718 824 2724 825
rect 2740 824 2742 846
rect 3088 835 3090 846
rect 2847 834 2851 835
rect 2975 834 2979 835
rect 3087 834 3091 835
rect 3111 834 3115 835
rect 2846 829 2852 830
rect 2846 825 2847 829
rect 2851 825 2852 829
rect 2846 824 2852 825
rect 2974 829 2980 830
rect 3087 829 3091 830
rect 3110 829 3116 830
rect 2974 825 2975 829
rect 2979 825 2980 829
rect 2974 824 2980 825
rect 3110 825 3111 829
rect 3115 825 3116 829
rect 3120 828 3122 850
rect 3192 835 3194 850
rect 3191 834 3195 835
rect 3191 829 3195 830
rect 3110 824 3116 825
rect 3118 827 3124 828
rect 2458 822 2464 823
rect 2622 823 2628 824
rect 2306 818 2312 819
rect 1598 816 1604 817
rect 1598 812 1599 816
rect 1603 812 1604 816
rect 1598 811 1604 812
rect 1600 795 1602 811
rect 1632 795 1634 818
rect 1670 807 1676 808
rect 1670 803 1671 807
rect 1675 803 1676 807
rect 1670 802 1676 803
rect 1599 794 1603 795
rect 1599 789 1603 790
rect 1631 794 1635 795
rect 1672 791 1674 802
rect 2278 800 2284 801
rect 2278 796 2279 800
rect 2283 796 2284 800
rect 2278 795 2284 796
rect 2280 791 2282 795
rect 1631 789 1635 790
rect 1671 790 1675 791
rect 1632 782 1634 789
rect 1671 785 1675 786
rect 2199 790 2203 791
rect 2199 785 2203 786
rect 2279 790 2283 791
rect 2279 785 2283 786
rect 1630 781 1636 782
rect 1630 777 1631 781
rect 1635 777 1636 781
rect 1672 778 1674 785
rect 2198 784 2204 785
rect 2198 780 2199 784
rect 2203 780 2204 784
rect 2198 779 2204 780
rect 1630 776 1636 777
rect 1670 777 1676 778
rect 1670 773 1671 777
rect 1675 773 1676 777
rect 1670 772 1676 773
rect 1422 762 1428 763
rect 1526 763 1532 764
rect 926 759 932 760
rect 926 755 927 759
rect 931 755 932 759
rect 926 754 932 755
rect 934 759 940 760
rect 934 755 935 759
rect 939 755 940 759
rect 934 754 940 755
rect 1046 759 1052 760
rect 1046 755 1047 759
rect 1051 755 1052 759
rect 1046 754 1052 755
rect 1058 759 1064 760
rect 1058 755 1059 759
rect 1063 755 1064 759
rect 1058 754 1064 755
rect 1166 759 1172 760
rect 1166 755 1167 759
rect 1171 755 1172 759
rect 1166 754 1172 755
rect 1190 759 1196 760
rect 1190 755 1191 759
rect 1195 755 1196 759
rect 1190 754 1196 755
rect 1278 759 1284 760
rect 1278 755 1279 759
rect 1283 755 1284 759
rect 1278 754 1284 755
rect 1302 759 1308 760
rect 1302 755 1303 759
rect 1307 755 1308 759
rect 1302 754 1308 755
rect 1398 759 1404 760
rect 1398 755 1399 759
rect 1403 755 1404 759
rect 1398 754 1404 755
rect 928 747 930 754
rect 927 746 931 747
rect 927 741 931 742
rect 936 736 938 754
rect 1048 747 1050 754
rect 951 746 955 747
rect 1047 746 1051 747
rect 950 741 956 742
rect 1047 741 1051 742
rect 950 737 951 741
rect 955 737 956 741
rect 950 736 956 737
rect 1060 736 1062 754
rect 1168 747 1170 754
rect 1071 746 1075 747
rect 1167 746 1171 747
rect 1183 746 1187 747
rect 1070 741 1076 742
rect 1167 741 1171 742
rect 1182 741 1188 742
rect 1070 737 1071 741
rect 1075 737 1076 741
rect 1070 736 1076 737
rect 1182 737 1183 741
rect 1187 737 1188 741
rect 1182 736 1188 737
rect 1192 736 1194 754
rect 1280 747 1282 754
rect 1279 746 1283 747
rect 1295 746 1299 747
rect 1279 741 1283 742
rect 1294 741 1300 742
rect 1294 737 1295 741
rect 1299 737 1300 741
rect 1294 736 1300 737
rect 1304 736 1306 754
rect 1400 747 1402 754
rect 1399 746 1403 747
rect 1415 746 1419 747
rect 1399 741 1403 742
rect 1414 741 1420 742
rect 1414 737 1415 741
rect 1419 737 1420 741
rect 1424 740 1426 762
rect 1518 759 1524 760
rect 1518 755 1519 759
rect 1523 755 1524 759
rect 1526 759 1527 763
rect 1531 759 1532 763
rect 1526 758 1532 759
rect 1630 763 1636 764
rect 1630 759 1631 763
rect 1635 759 1636 763
rect 1630 758 1636 759
rect 1670 759 1676 760
rect 1518 754 1524 755
rect 1520 747 1522 754
rect 1632 747 1634 758
rect 1670 755 1671 759
rect 1675 755 1676 759
rect 1670 754 1676 755
rect 2198 755 2204 756
rect 1672 747 1674 754
rect 2198 751 2199 755
rect 2203 751 2204 755
rect 2198 750 2204 751
rect 2158 747 2164 748
rect 2200 747 2202 750
rect 1519 746 1523 747
rect 1519 741 1523 742
rect 1631 746 1635 747
rect 1631 741 1635 742
rect 1671 746 1675 747
rect 2127 746 2131 747
rect 2158 743 2159 747
rect 2163 743 2164 747
rect 2158 742 2164 743
rect 2199 746 2203 747
rect 2287 746 2291 747
rect 1671 741 1675 742
rect 2126 741 2132 742
rect 1414 736 1420 737
rect 1422 739 1428 740
rect 110 732 116 733
rect 582 735 588 736
rect 582 731 583 735
rect 587 731 588 735
rect 582 730 588 731
rect 614 735 620 736
rect 614 731 615 735
rect 619 731 620 735
rect 614 730 620 731
rect 814 735 820 736
rect 814 731 815 735
rect 819 731 820 735
rect 814 730 820 731
rect 854 735 860 736
rect 854 731 855 735
rect 859 731 860 735
rect 854 730 860 731
rect 886 735 892 736
rect 886 731 887 735
rect 891 731 892 735
rect 886 730 892 731
rect 934 735 940 736
rect 934 731 935 735
rect 939 731 940 735
rect 934 730 940 731
rect 1058 735 1064 736
rect 1058 731 1059 735
rect 1063 731 1064 735
rect 1058 730 1064 731
rect 1190 735 1196 736
rect 1190 731 1191 735
rect 1195 731 1196 735
rect 1190 730 1196 731
rect 1302 735 1308 736
rect 1302 731 1303 735
rect 1307 731 1308 735
rect 1302 730 1308 731
rect 1318 735 1324 736
rect 1318 731 1319 735
rect 1323 731 1324 735
rect 1422 735 1423 739
rect 1427 735 1428 739
rect 1632 738 1634 741
rect 1672 738 1674 741
rect 1422 734 1428 735
rect 1630 737 1636 738
rect 1630 733 1631 737
rect 1635 733 1636 737
rect 1630 732 1636 733
rect 1670 737 1676 738
rect 1670 733 1671 737
rect 1675 733 1676 737
rect 2126 737 2127 741
rect 2131 737 2132 741
rect 2126 736 2132 737
rect 2160 736 2162 742
rect 2199 741 2203 742
rect 2286 741 2292 742
rect 2286 737 2287 741
rect 2291 737 2292 741
rect 2286 736 2292 737
rect 2308 736 2310 818
rect 2438 800 2444 801
rect 2438 796 2439 800
rect 2443 796 2444 800
rect 2438 795 2444 796
rect 2440 791 2442 795
rect 2359 790 2363 791
rect 2359 785 2363 786
rect 2439 790 2443 791
rect 2439 785 2443 786
rect 2358 784 2364 785
rect 2358 780 2359 784
rect 2363 780 2364 784
rect 2358 779 2364 780
rect 2460 760 2462 822
rect 2622 819 2623 823
rect 2627 819 2628 823
rect 2622 818 2628 819
rect 2738 823 2744 824
rect 2738 819 2739 823
rect 2743 819 2744 823
rect 2738 818 2744 819
rect 2798 823 2804 824
rect 2798 819 2799 823
rect 2803 819 2804 823
rect 2798 818 2804 819
rect 2930 823 2936 824
rect 2930 819 2931 823
rect 2935 819 2936 823
rect 2930 818 2936 819
rect 3054 823 3060 824
rect 3054 819 3055 823
rect 3059 819 3060 823
rect 3118 823 3119 827
rect 3123 823 3124 827
rect 3192 826 3194 829
rect 3118 822 3124 823
rect 3190 825 3196 826
rect 3190 821 3191 825
rect 3195 821 3196 825
rect 3190 820 3196 821
rect 3054 818 3060 819
rect 2582 800 2588 801
rect 2582 796 2583 800
rect 2587 796 2588 800
rect 2582 795 2588 796
rect 2584 791 2586 795
rect 2511 790 2515 791
rect 2511 785 2515 786
rect 2583 790 2587 791
rect 2583 785 2587 786
rect 2510 784 2516 785
rect 2510 780 2511 784
rect 2515 780 2516 784
rect 2510 779 2516 780
rect 2624 760 2626 818
rect 2718 800 2724 801
rect 2718 796 2719 800
rect 2723 796 2724 800
rect 2718 795 2724 796
rect 2720 791 2722 795
rect 2655 790 2659 791
rect 2655 785 2659 786
rect 2719 790 2723 791
rect 2719 785 2723 786
rect 2791 790 2795 791
rect 2791 785 2795 786
rect 2654 784 2660 785
rect 2654 780 2655 784
rect 2659 780 2660 784
rect 2654 779 2660 780
rect 2790 784 2796 785
rect 2790 780 2791 784
rect 2795 780 2796 784
rect 2790 779 2796 780
rect 2458 759 2464 760
rect 2358 755 2364 756
rect 2358 751 2359 755
rect 2363 751 2364 755
rect 2458 755 2459 759
rect 2463 755 2464 759
rect 2622 759 2628 760
rect 2458 754 2464 755
rect 2510 755 2516 756
rect 2358 750 2364 751
rect 2360 747 2362 750
rect 2359 746 2363 747
rect 2447 746 2451 747
rect 2359 741 2363 742
rect 2446 741 2452 742
rect 2446 737 2447 741
rect 2451 737 2452 741
rect 2446 736 2452 737
rect 2460 736 2462 754
rect 2510 751 2511 755
rect 2515 751 2516 755
rect 2622 755 2623 759
rect 2627 755 2628 759
rect 2800 756 2802 818
rect 2846 800 2852 801
rect 2846 796 2847 800
rect 2851 796 2852 800
rect 2846 795 2852 796
rect 2848 791 2850 795
rect 2847 790 2851 791
rect 2847 785 2851 786
rect 2919 790 2923 791
rect 2919 785 2923 786
rect 2918 784 2924 785
rect 2918 780 2919 784
rect 2923 780 2924 784
rect 2918 779 2924 780
rect 2932 760 2934 818
rect 2974 800 2980 801
rect 2974 796 2975 800
rect 2979 796 2980 800
rect 2974 795 2980 796
rect 2976 791 2978 795
rect 2975 790 2979 791
rect 2975 785 2979 786
rect 3047 790 3051 791
rect 3047 785 3051 786
rect 3046 784 3052 785
rect 3046 780 3047 784
rect 3051 780 3052 784
rect 3046 779 3052 780
rect 3056 760 3058 818
rect 3190 807 3196 808
rect 3190 803 3191 807
rect 3195 803 3196 807
rect 3190 802 3196 803
rect 3110 800 3116 801
rect 3110 796 3111 800
rect 3115 796 3116 800
rect 3110 795 3116 796
rect 3112 791 3114 795
rect 3192 791 3194 802
rect 3111 790 3115 791
rect 3111 785 3115 786
rect 3159 790 3163 791
rect 3159 785 3163 786
rect 3191 790 3195 791
rect 3191 785 3195 786
rect 3158 784 3164 785
rect 3158 780 3159 784
rect 3163 780 3164 784
rect 3158 779 3164 780
rect 3192 778 3194 785
rect 3190 777 3196 778
rect 3190 773 3191 777
rect 3195 773 3196 777
rect 3190 772 3196 773
rect 2930 759 2936 760
rect 2622 754 2628 755
rect 2654 755 2660 756
rect 2510 750 2516 751
rect 2512 747 2514 750
rect 2511 746 2515 747
rect 2599 746 2603 747
rect 2511 741 2515 742
rect 2598 741 2604 742
rect 2598 737 2599 741
rect 2603 737 2604 741
rect 2598 736 2604 737
rect 2624 736 2626 754
rect 2654 751 2655 755
rect 2659 751 2660 755
rect 2654 750 2660 751
rect 2766 755 2772 756
rect 2766 751 2767 755
rect 2771 751 2772 755
rect 2766 750 2772 751
rect 2790 755 2796 756
rect 2790 751 2791 755
rect 2795 751 2796 755
rect 2790 750 2796 751
rect 2798 755 2804 756
rect 2798 751 2799 755
rect 2803 751 2804 755
rect 2798 750 2804 751
rect 2918 755 2924 756
rect 2918 751 2919 755
rect 2923 751 2924 755
rect 2930 755 2931 759
rect 2935 755 2936 759
rect 3054 759 3060 760
rect 2930 754 2936 755
rect 3046 755 3052 756
rect 2918 750 2924 751
rect 2656 747 2658 750
rect 2655 746 2659 747
rect 2759 746 2763 747
rect 2655 741 2659 742
rect 2758 741 2764 742
rect 2758 737 2759 741
rect 2763 737 2764 741
rect 2758 736 2764 737
rect 2768 736 2770 750
rect 2792 747 2794 750
rect 2791 746 2795 747
rect 2791 741 2795 742
rect 2800 736 2802 750
rect 2920 747 2922 750
rect 2919 746 2923 747
rect 2918 741 2924 742
rect 2918 737 2919 741
rect 2923 737 2924 741
rect 2932 740 2934 754
rect 3046 751 3047 755
rect 3051 751 3052 755
rect 3054 755 3055 759
rect 3059 755 3060 759
rect 3190 759 3196 760
rect 3054 754 3060 755
rect 3158 755 3164 756
rect 3046 750 3052 751
rect 3158 751 3159 755
rect 3163 751 3164 755
rect 3158 750 3164 751
rect 3166 755 3172 756
rect 3166 751 3167 755
rect 3171 751 3172 755
rect 3190 755 3191 759
rect 3195 755 3196 759
rect 3190 754 3196 755
rect 3166 750 3172 751
rect 3048 747 3050 750
rect 3160 747 3162 750
rect 3047 746 3051 747
rect 3047 741 3051 742
rect 3159 746 3163 747
rect 3159 741 3163 742
rect 2918 736 2924 737
rect 2930 739 2936 740
rect 1670 732 1676 733
rect 2158 735 2164 736
rect 1318 730 1324 731
rect 2158 731 2159 735
rect 2163 731 2164 735
rect 2158 730 2164 731
rect 2306 735 2312 736
rect 2306 731 2307 735
rect 2311 731 2312 735
rect 2306 730 2312 731
rect 2458 735 2464 736
rect 2458 731 2459 735
rect 2463 731 2464 735
rect 2458 730 2464 731
rect 2622 735 2628 736
rect 2622 731 2623 735
rect 2627 731 2628 735
rect 2622 730 2628 731
rect 2766 735 2772 736
rect 2766 731 2767 735
rect 2771 731 2772 735
rect 2766 730 2772 731
rect 2798 735 2804 736
rect 2798 731 2799 735
rect 2803 731 2804 735
rect 2930 735 2931 739
rect 2935 735 2936 739
rect 2930 734 2936 735
rect 2798 730 2804 731
rect 110 719 116 720
rect 110 715 111 719
rect 115 715 116 719
rect 110 714 116 715
rect 112 695 114 714
rect 574 712 580 713
rect 574 708 575 712
rect 579 708 580 712
rect 574 707 580 708
rect 576 695 578 707
rect 111 694 115 695
rect 111 689 115 690
rect 479 694 483 695
rect 479 689 483 690
rect 575 694 579 695
rect 575 689 579 690
rect 607 694 611 695
rect 607 689 611 690
rect 112 682 114 689
rect 478 688 484 689
rect 478 684 479 688
rect 483 684 484 688
rect 478 683 484 684
rect 606 688 612 689
rect 606 684 607 688
rect 611 684 612 688
rect 606 683 612 684
rect 110 681 116 682
rect 110 677 111 681
rect 115 677 116 681
rect 110 676 116 677
rect 110 663 116 664
rect 110 659 111 663
rect 115 659 116 663
rect 616 660 618 730
rect 702 712 708 713
rect 702 708 703 712
rect 707 708 708 712
rect 702 707 708 708
rect 830 712 836 713
rect 830 708 831 712
rect 835 708 836 712
rect 830 707 836 708
rect 704 695 706 707
rect 832 695 834 707
rect 703 694 707 695
rect 703 689 707 690
rect 727 694 731 695
rect 727 689 731 690
rect 831 694 835 695
rect 831 689 835 690
rect 847 694 851 695
rect 847 689 851 690
rect 726 688 732 689
rect 726 684 727 688
rect 731 684 732 688
rect 726 683 732 684
rect 846 688 852 689
rect 846 684 847 688
rect 851 684 852 688
rect 846 683 852 684
rect 856 660 858 730
rect 950 712 956 713
rect 950 708 951 712
rect 955 708 956 712
rect 950 707 956 708
rect 1070 712 1076 713
rect 1070 708 1071 712
rect 1075 708 1076 712
rect 1070 707 1076 708
rect 1182 712 1188 713
rect 1182 708 1183 712
rect 1187 708 1188 712
rect 1182 707 1188 708
rect 1294 712 1300 713
rect 1294 708 1295 712
rect 1299 708 1300 712
rect 1294 707 1300 708
rect 952 695 954 707
rect 1072 695 1074 707
rect 1184 695 1186 707
rect 1296 695 1298 707
rect 951 694 955 695
rect 951 689 955 690
rect 967 694 971 695
rect 967 689 971 690
rect 1071 694 1075 695
rect 1071 689 1075 690
rect 1079 694 1083 695
rect 1079 689 1083 690
rect 1183 694 1187 695
rect 1183 689 1187 690
rect 1191 694 1195 695
rect 1191 689 1195 690
rect 1295 694 1299 695
rect 1295 689 1299 690
rect 1311 694 1315 695
rect 1311 689 1315 690
rect 966 688 972 689
rect 966 684 967 688
rect 971 684 972 688
rect 966 683 972 684
rect 1078 688 1084 689
rect 1078 684 1079 688
rect 1083 684 1084 688
rect 1078 683 1084 684
rect 1190 688 1196 689
rect 1190 684 1191 688
rect 1195 684 1196 688
rect 1190 683 1196 684
rect 1310 688 1316 689
rect 1310 684 1311 688
rect 1315 684 1316 688
rect 1310 683 1316 684
rect 1320 664 1322 730
rect 1630 719 1636 720
rect 1630 715 1631 719
rect 1635 715 1636 719
rect 1630 714 1636 715
rect 1670 719 1676 720
rect 1670 715 1671 719
rect 1675 715 1676 719
rect 1670 714 1676 715
rect 1414 712 1420 713
rect 1414 708 1415 712
rect 1419 708 1420 712
rect 1414 707 1420 708
rect 1416 695 1418 707
rect 1632 695 1634 714
rect 1672 707 1674 714
rect 2126 712 2132 713
rect 2126 708 2127 712
rect 2131 708 2132 712
rect 2126 707 2132 708
rect 1671 706 1675 707
rect 1671 701 1675 702
rect 2023 706 2027 707
rect 2023 701 2027 702
rect 2127 706 2131 707
rect 2127 701 2131 702
rect 2151 706 2155 707
rect 2151 701 2155 702
rect 1415 694 1419 695
rect 1415 689 1419 690
rect 1631 694 1635 695
rect 1672 694 1674 701
rect 2022 700 2028 701
rect 2022 696 2023 700
rect 2027 696 2028 700
rect 2022 695 2028 696
rect 2150 700 2156 701
rect 2150 696 2151 700
rect 2155 696 2156 700
rect 2150 695 2156 696
rect 1631 689 1635 690
rect 1670 693 1676 694
rect 1670 689 1671 693
rect 1675 689 1676 693
rect 1632 682 1634 689
rect 1670 688 1676 689
rect 1630 681 1636 682
rect 1630 677 1631 681
rect 1635 677 1636 681
rect 1630 676 1636 677
rect 1670 675 1676 676
rect 1670 671 1671 675
rect 1675 671 1676 675
rect 2160 672 2162 730
rect 2286 712 2292 713
rect 2286 708 2287 712
rect 2291 708 2292 712
rect 2286 707 2292 708
rect 2287 706 2291 707
rect 2287 701 2291 702
rect 2295 706 2299 707
rect 2295 701 2299 702
rect 2294 700 2300 701
rect 2294 696 2295 700
rect 2299 696 2300 700
rect 2294 695 2300 696
rect 2308 672 2310 730
rect 2446 712 2452 713
rect 2446 708 2447 712
rect 2451 708 2452 712
rect 2446 707 2452 708
rect 2447 706 2451 707
rect 2447 701 2451 702
rect 2446 700 2452 701
rect 2446 696 2447 700
rect 2451 696 2452 700
rect 2446 695 2452 696
rect 2460 672 2462 730
rect 2598 712 2604 713
rect 2598 708 2599 712
rect 2603 708 2604 712
rect 2598 707 2604 708
rect 2599 706 2603 707
rect 2599 701 2603 702
rect 2615 706 2619 707
rect 2615 701 2619 702
rect 2614 700 2620 701
rect 2614 696 2615 700
rect 2619 696 2620 700
rect 2614 695 2620 696
rect 2624 672 2626 730
rect 2758 712 2764 713
rect 2758 708 2759 712
rect 2763 708 2764 712
rect 2758 707 2764 708
rect 2759 706 2763 707
rect 2759 701 2763 702
rect 1670 670 1676 671
rect 2022 671 2028 672
rect 1222 663 1228 664
rect 110 658 116 659
rect 478 659 484 660
rect 112 643 114 658
rect 478 655 479 659
rect 483 655 484 659
rect 478 654 484 655
rect 486 659 492 660
rect 486 655 487 659
rect 491 655 492 659
rect 486 654 492 655
rect 606 659 612 660
rect 606 655 607 659
rect 611 655 612 659
rect 606 654 612 655
rect 614 659 620 660
rect 614 655 615 659
rect 619 655 620 659
rect 614 654 620 655
rect 630 659 636 660
rect 630 655 631 659
rect 635 655 636 659
rect 630 654 636 655
rect 726 659 732 660
rect 726 655 727 659
rect 731 655 732 659
rect 726 654 732 655
rect 750 659 756 660
rect 750 655 751 659
rect 755 655 756 659
rect 750 654 756 655
rect 846 659 852 660
rect 846 655 847 659
rect 851 655 852 659
rect 846 654 852 655
rect 854 659 860 660
rect 854 655 855 659
rect 859 655 860 659
rect 854 654 860 655
rect 966 659 972 660
rect 966 655 967 659
rect 971 655 972 659
rect 966 654 972 655
rect 998 659 1004 660
rect 998 655 999 659
rect 1003 655 1004 659
rect 998 654 1004 655
rect 1078 659 1084 660
rect 1078 655 1079 659
rect 1083 655 1084 659
rect 1078 654 1084 655
rect 1102 659 1108 660
rect 1102 655 1103 659
rect 1107 655 1108 659
rect 1102 654 1108 655
rect 1190 659 1196 660
rect 1190 655 1191 659
rect 1195 655 1196 659
rect 1222 659 1223 663
rect 1227 659 1228 663
rect 1318 663 1324 664
rect 1222 658 1228 659
rect 1310 659 1316 660
rect 1190 654 1196 655
rect 480 643 482 654
rect 111 642 115 643
rect 375 642 379 643
rect 479 642 483 643
rect 111 637 115 638
rect 374 637 380 638
rect 479 637 483 638
rect 112 634 114 637
rect 110 633 116 634
rect 110 629 111 633
rect 115 629 116 633
rect 374 633 375 637
rect 379 633 380 637
rect 374 632 380 633
rect 488 632 490 654
rect 608 643 610 654
rect 503 642 507 643
rect 607 642 611 643
rect 623 642 627 643
rect 502 637 508 638
rect 607 637 611 638
rect 622 637 628 638
rect 502 633 503 637
rect 507 633 508 637
rect 502 632 508 633
rect 622 633 623 637
rect 627 633 628 637
rect 622 632 628 633
rect 632 632 634 654
rect 728 643 730 654
rect 727 642 731 643
rect 743 642 747 643
rect 727 637 731 638
rect 742 637 748 638
rect 742 633 743 637
rect 747 633 748 637
rect 752 636 754 654
rect 848 643 850 654
rect 847 642 851 643
rect 847 637 851 638
rect 742 632 748 633
rect 750 635 756 636
rect 110 628 116 629
rect 406 631 412 632
rect 406 627 407 631
rect 411 627 412 631
rect 406 626 412 627
rect 486 631 492 632
rect 486 627 487 631
rect 491 627 492 631
rect 486 626 492 627
rect 630 631 636 632
rect 630 627 631 631
rect 635 627 636 631
rect 630 626 636 627
rect 670 631 676 632
rect 670 627 671 631
rect 675 627 676 631
rect 750 631 751 635
rect 755 631 756 635
rect 750 630 756 631
rect 774 635 780 636
rect 774 631 775 635
rect 779 631 780 635
rect 856 632 858 654
rect 968 643 970 654
rect 863 642 867 643
rect 967 642 971 643
rect 975 642 979 643
rect 862 637 868 638
rect 967 637 971 638
rect 974 637 980 638
rect 862 633 863 637
rect 867 633 868 637
rect 862 632 868 633
rect 974 633 975 637
rect 979 633 980 637
rect 974 632 980 633
rect 1000 632 1002 654
rect 1080 643 1082 654
rect 1079 642 1083 643
rect 1095 642 1099 643
rect 1079 637 1083 638
rect 1094 637 1100 638
rect 1094 633 1095 637
rect 1099 633 1100 637
rect 1094 632 1100 633
rect 1104 632 1106 654
rect 1192 643 1194 654
rect 1191 642 1195 643
rect 1215 642 1219 643
rect 1191 637 1195 638
rect 1214 637 1220 638
rect 1214 633 1215 637
rect 1219 633 1220 637
rect 1224 636 1226 658
rect 1310 655 1311 659
rect 1315 655 1316 659
rect 1318 659 1319 663
rect 1323 659 1324 663
rect 1318 658 1324 659
rect 1630 663 1636 664
rect 1630 659 1631 663
rect 1635 659 1636 663
rect 1672 659 1674 670
rect 2022 667 2023 671
rect 2027 667 2028 671
rect 2022 666 2028 667
rect 2030 671 2036 672
rect 2030 667 2031 671
rect 2035 667 2036 671
rect 2030 666 2036 667
rect 2150 671 2156 672
rect 2150 667 2151 671
rect 2155 667 2156 671
rect 2150 666 2156 667
rect 2158 671 2164 672
rect 2158 667 2159 671
rect 2163 667 2164 671
rect 2158 666 2164 667
rect 2294 671 2300 672
rect 2294 667 2295 671
rect 2299 667 2300 671
rect 2294 666 2300 667
rect 2306 671 2312 672
rect 2306 667 2307 671
rect 2311 667 2312 671
rect 2306 666 2312 667
rect 2446 671 2452 672
rect 2446 667 2447 671
rect 2451 667 2452 671
rect 2446 666 2452 667
rect 2458 671 2464 672
rect 2458 667 2459 671
rect 2463 667 2464 671
rect 2458 666 2464 667
rect 2614 671 2620 672
rect 2614 667 2615 671
rect 2619 667 2620 671
rect 2614 666 2620 667
rect 2622 671 2628 672
rect 2622 667 2623 671
rect 2627 667 2628 671
rect 2622 666 2628 667
rect 2024 659 2026 666
rect 1630 658 1636 659
rect 1671 658 1675 659
rect 1310 654 1316 655
rect 1312 643 1314 654
rect 1632 643 1634 658
rect 1919 658 1923 659
rect 2023 658 2027 659
rect 1671 653 1675 654
rect 1918 653 1924 654
rect 2023 653 2027 654
rect 1672 650 1674 653
rect 1670 649 1676 650
rect 1670 645 1671 649
rect 1675 645 1676 649
rect 1918 649 1919 653
rect 1923 649 1924 653
rect 1918 648 1924 649
rect 2032 648 2034 666
rect 2152 659 2154 666
rect 2047 658 2051 659
rect 2151 658 2155 659
rect 2046 653 2052 654
rect 2151 653 2155 654
rect 2046 649 2047 653
rect 2051 649 2052 653
rect 2046 648 2052 649
rect 2160 648 2162 666
rect 2296 659 2298 666
rect 2183 658 2187 659
rect 2295 658 2299 659
rect 2182 653 2188 654
rect 2295 653 2299 654
rect 2182 649 2183 653
rect 2187 649 2188 653
rect 2182 648 2188 649
rect 2308 648 2310 666
rect 2448 659 2450 666
rect 2327 658 2331 659
rect 2447 658 2451 659
rect 2326 653 2332 654
rect 2447 653 2451 654
rect 2326 649 2327 653
rect 2331 649 2332 653
rect 2326 648 2332 649
rect 2460 648 2462 666
rect 2616 659 2618 666
rect 2471 658 2475 659
rect 2615 658 2619 659
rect 2470 653 2476 654
rect 2470 649 2471 653
rect 2475 649 2476 653
rect 2470 648 2476 649
rect 2614 653 2620 654
rect 2614 649 2615 653
rect 2619 649 2620 653
rect 2614 648 2620 649
rect 2624 648 2626 666
rect 2759 658 2763 659
rect 2758 653 2764 654
rect 2758 649 2759 653
rect 2763 649 2764 653
rect 2768 652 2770 730
rect 2918 712 2924 713
rect 2918 708 2919 712
rect 2923 708 2924 712
rect 2918 707 2924 708
rect 2799 706 2803 707
rect 2799 701 2803 702
rect 2919 706 2923 707
rect 2919 701 2923 702
rect 2798 700 2804 701
rect 2798 696 2799 700
rect 2803 696 2804 700
rect 2798 695 2804 696
rect 2932 680 2934 734
rect 2991 706 2995 707
rect 2991 701 2995 702
rect 3159 706 3163 707
rect 3159 701 3163 702
rect 2990 700 2996 701
rect 2990 696 2991 700
rect 2995 696 2996 700
rect 2990 695 2996 696
rect 3158 700 3164 701
rect 3158 696 3159 700
rect 3163 696 3164 700
rect 3158 695 3164 696
rect 2930 679 2936 680
rect 2930 675 2931 679
rect 2935 675 2936 679
rect 3168 676 3170 750
rect 3192 747 3194 754
rect 3191 746 3195 747
rect 3191 741 3195 742
rect 3192 738 3194 741
rect 3190 737 3196 738
rect 3190 733 3191 737
rect 3195 733 3196 737
rect 3190 732 3196 733
rect 3190 719 3196 720
rect 3190 715 3191 719
rect 3195 715 3196 719
rect 3190 714 3196 715
rect 3192 707 3194 714
rect 3191 706 3195 707
rect 3191 701 3195 702
rect 3192 694 3194 701
rect 3190 693 3196 694
rect 3190 689 3191 693
rect 3195 689 3196 693
rect 3190 688 3196 689
rect 2930 674 2936 675
rect 3166 675 3172 676
rect 2798 671 2804 672
rect 2798 667 2799 671
rect 2803 667 2804 671
rect 2798 666 2804 667
rect 2806 671 2812 672
rect 2806 667 2807 671
rect 2811 667 2812 671
rect 2806 666 2812 667
rect 2870 671 2876 672
rect 2870 667 2871 671
rect 2875 667 2876 671
rect 2870 666 2876 667
rect 2990 671 2996 672
rect 2990 667 2991 671
rect 2995 667 2996 671
rect 2990 666 2996 667
rect 3158 671 3164 672
rect 3158 667 3159 671
rect 3163 667 3164 671
rect 3166 671 3167 675
rect 3171 671 3172 675
rect 3166 670 3172 671
rect 3190 675 3196 676
rect 3190 671 3191 675
rect 3195 671 3196 675
rect 3190 670 3196 671
rect 3158 666 3164 667
rect 2800 659 2802 666
rect 2799 658 2803 659
rect 2799 653 2803 654
rect 2808 652 2810 666
rect 2758 648 2764 649
rect 2766 651 2772 652
rect 1670 644 1676 645
rect 1894 647 1900 648
rect 1894 643 1895 647
rect 1899 643 1900 647
rect 1311 642 1315 643
rect 1311 637 1315 638
rect 1631 642 1635 643
rect 1894 642 1900 643
rect 2030 647 2036 648
rect 2030 643 2031 647
rect 2035 643 2036 647
rect 2030 642 2036 643
rect 2158 647 2164 648
rect 2158 643 2159 647
rect 2163 643 2164 647
rect 2158 642 2164 643
rect 2190 647 2196 648
rect 2190 643 2191 647
rect 2195 643 2196 647
rect 2190 642 2196 643
rect 2306 647 2312 648
rect 2306 643 2307 647
rect 2311 643 2312 647
rect 2306 642 2312 643
rect 2458 647 2464 648
rect 2458 643 2459 647
rect 2463 643 2464 647
rect 2458 642 2464 643
rect 2622 647 2628 648
rect 2622 643 2623 647
rect 2627 643 2628 647
rect 2766 647 2767 651
rect 2771 647 2772 651
rect 2766 646 2772 647
rect 2806 651 2812 652
rect 2806 647 2807 651
rect 2811 647 2812 651
rect 2806 646 2812 647
rect 2622 642 2628 643
rect 1631 637 1635 638
rect 1214 632 1220 633
rect 1222 635 1228 636
rect 774 630 780 631
rect 854 631 860 632
rect 670 626 676 627
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 110 610 116 611
rect 112 595 114 610
rect 374 608 380 609
rect 374 604 375 608
rect 379 604 380 608
rect 374 603 380 604
rect 376 595 378 603
rect 111 594 115 595
rect 111 589 115 590
rect 271 594 275 595
rect 271 589 275 590
rect 375 594 379 595
rect 375 589 379 590
rect 399 594 403 595
rect 399 589 403 590
rect 112 582 114 589
rect 270 588 276 589
rect 270 584 271 588
rect 275 584 276 588
rect 270 583 276 584
rect 398 588 404 589
rect 398 584 399 588
rect 403 584 404 588
rect 398 583 404 584
rect 110 581 116 582
rect 110 577 111 581
rect 115 577 116 581
rect 110 576 116 577
rect 110 563 116 564
rect 110 559 111 563
rect 115 559 116 563
rect 408 560 410 626
rect 502 608 508 609
rect 502 604 503 608
rect 507 604 508 608
rect 502 603 508 604
rect 622 608 628 609
rect 622 604 623 608
rect 627 604 628 608
rect 622 603 628 604
rect 504 595 506 603
rect 624 595 626 603
rect 503 594 507 595
rect 503 589 507 590
rect 527 594 531 595
rect 527 589 531 590
rect 623 594 627 595
rect 623 589 627 590
rect 647 594 651 595
rect 647 589 651 590
rect 526 588 532 589
rect 526 584 527 588
rect 531 584 532 588
rect 526 583 532 584
rect 646 588 652 589
rect 646 584 647 588
rect 651 584 652 588
rect 646 583 652 584
rect 672 560 674 626
rect 742 608 748 609
rect 742 604 743 608
rect 747 604 748 608
rect 742 603 748 604
rect 744 595 746 603
rect 743 594 747 595
rect 743 589 747 590
rect 767 594 771 595
rect 767 589 771 590
rect 766 588 772 589
rect 766 584 767 588
rect 771 584 772 588
rect 766 583 772 584
rect 776 564 778 630
rect 854 627 855 631
rect 859 627 860 631
rect 854 626 860 627
rect 998 631 1004 632
rect 998 627 999 631
rect 1003 627 1004 631
rect 998 626 1004 627
rect 1102 631 1108 632
rect 1102 627 1103 631
rect 1107 627 1108 631
rect 1222 631 1223 635
rect 1227 631 1228 635
rect 1632 634 1634 637
rect 1222 630 1228 631
rect 1630 633 1636 634
rect 1630 629 1631 633
rect 1635 629 1636 633
rect 1630 628 1636 629
rect 1670 631 1676 632
rect 1102 626 1108 627
rect 1670 627 1671 631
rect 1675 627 1676 631
rect 1670 626 1676 627
rect 862 608 868 609
rect 862 604 863 608
rect 867 604 868 608
rect 862 603 868 604
rect 974 608 980 609
rect 974 604 975 608
rect 979 604 980 608
rect 974 603 980 604
rect 864 595 866 603
rect 976 595 978 603
rect 863 594 867 595
rect 863 589 867 590
rect 879 594 883 595
rect 879 589 883 590
rect 975 594 979 595
rect 975 589 979 590
rect 991 594 995 595
rect 991 589 995 590
rect 878 588 884 589
rect 878 584 879 588
rect 883 584 884 588
rect 878 583 884 584
rect 990 588 996 589
rect 990 584 991 588
rect 995 584 996 588
rect 990 583 996 584
rect 775 563 781 564
rect 110 558 116 559
rect 270 559 276 560
rect 112 543 114 558
rect 270 555 271 559
rect 275 555 276 559
rect 270 554 276 555
rect 310 559 316 560
rect 310 555 311 559
rect 315 555 316 559
rect 310 554 316 555
rect 398 559 404 560
rect 398 555 399 559
rect 403 555 404 559
rect 398 554 404 555
rect 406 559 412 560
rect 406 555 407 559
rect 411 555 412 559
rect 406 554 412 555
rect 430 559 436 560
rect 430 555 431 559
rect 435 555 436 559
rect 430 554 436 555
rect 526 559 532 560
rect 526 555 527 559
rect 531 555 532 559
rect 526 554 532 555
rect 550 559 556 560
rect 550 555 551 559
rect 555 555 556 559
rect 550 554 556 555
rect 646 559 652 560
rect 646 555 647 559
rect 651 555 652 559
rect 646 554 652 555
rect 670 559 676 560
rect 670 555 671 559
rect 675 555 676 559
rect 670 554 676 555
rect 766 559 772 560
rect 766 555 767 559
rect 771 555 772 559
rect 775 559 776 563
rect 780 561 786 563
rect 780 559 781 561
rect 775 558 781 559
rect 766 554 772 555
rect 272 543 274 554
rect 312 552 314 554
rect 310 551 316 552
rect 310 547 311 551
rect 315 547 316 551
rect 310 546 316 547
rect 111 542 115 543
rect 175 542 179 543
rect 271 542 275 543
rect 303 542 307 543
rect 111 537 115 538
rect 174 537 180 538
rect 271 537 275 538
rect 302 537 308 538
rect 112 534 114 537
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 174 533 175 537
rect 179 533 180 537
rect 174 532 180 533
rect 302 533 303 537
rect 307 533 308 537
rect 302 532 308 533
rect 312 532 314 546
rect 400 543 402 554
rect 432 552 434 554
rect 430 551 436 552
rect 430 547 431 551
rect 435 547 436 551
rect 430 546 436 547
rect 399 542 403 543
rect 423 542 427 543
rect 399 537 403 538
rect 422 537 428 538
rect 422 533 423 537
rect 427 533 428 537
rect 432 536 434 546
rect 528 543 530 554
rect 527 542 531 543
rect 543 542 547 543
rect 527 537 531 538
rect 542 537 548 538
rect 422 532 428 533
rect 430 535 436 536
rect 110 528 116 529
rect 146 531 152 532
rect 146 527 147 531
rect 151 527 152 531
rect 146 526 152 527
rect 310 531 316 532
rect 310 527 311 531
rect 315 527 316 531
rect 430 531 431 535
rect 435 531 436 535
rect 542 533 543 537
rect 547 533 548 537
rect 542 532 548 533
rect 552 532 554 554
rect 648 543 650 554
rect 647 542 651 543
rect 663 542 667 543
rect 647 537 651 538
rect 662 537 668 538
rect 662 533 663 537
rect 667 533 668 537
rect 662 532 668 533
rect 672 532 674 554
rect 768 543 770 554
rect 767 542 771 543
rect 775 542 779 543
rect 767 537 771 538
rect 774 537 780 538
rect 774 533 775 537
rect 779 533 780 537
rect 784 536 786 561
rect 1000 560 1002 626
rect 1630 615 1636 616
rect 1672 615 1674 626
rect 1630 611 1631 615
rect 1635 611 1636 615
rect 1630 610 1636 611
rect 1671 614 1675 615
rect 1094 608 1100 609
rect 1094 604 1095 608
rect 1099 604 1100 608
rect 1094 603 1100 604
rect 1214 608 1220 609
rect 1214 604 1215 608
rect 1219 604 1220 608
rect 1214 603 1220 604
rect 1096 595 1098 603
rect 1216 595 1218 603
rect 1632 595 1634 610
rect 1671 609 1675 610
rect 1847 614 1851 615
rect 1847 609 1851 610
rect 1672 602 1674 609
rect 1846 608 1852 609
rect 1846 604 1847 608
rect 1851 604 1852 608
rect 1846 603 1852 604
rect 1670 601 1676 602
rect 1670 597 1671 601
rect 1675 597 1676 601
rect 1670 596 1676 597
rect 1095 594 1099 595
rect 1095 589 1099 590
rect 1111 594 1115 595
rect 1111 589 1115 590
rect 1215 594 1219 595
rect 1215 589 1219 590
rect 1631 594 1635 595
rect 1631 589 1635 590
rect 1110 588 1116 589
rect 1110 584 1111 588
rect 1115 584 1116 588
rect 1110 583 1116 584
rect 1632 582 1634 589
rect 1670 583 1676 584
rect 1630 581 1636 582
rect 1630 577 1631 581
rect 1635 577 1636 581
rect 1670 579 1671 583
rect 1675 579 1676 583
rect 1670 578 1676 579
rect 1846 579 1852 580
rect 1630 576 1636 577
rect 1672 575 1674 578
rect 1846 575 1847 579
rect 1851 575 1852 579
rect 1671 574 1675 575
rect 1767 574 1771 575
rect 1846 574 1852 575
rect 1671 569 1675 570
rect 1766 569 1772 570
rect 1847 569 1851 570
rect 1672 566 1674 569
rect 1670 565 1676 566
rect 1630 563 1636 564
rect 878 559 884 560
rect 878 555 879 559
rect 883 555 884 559
rect 878 554 884 555
rect 886 559 892 560
rect 886 555 887 559
rect 891 555 892 559
rect 990 559 996 560
rect 990 555 991 559
rect 995 555 996 559
rect 886 554 898 555
rect 990 554 996 555
rect 998 559 1004 560
rect 998 555 999 559
rect 1003 555 1004 559
rect 998 554 1004 555
rect 1110 559 1116 560
rect 1110 555 1111 559
rect 1115 555 1116 559
rect 1110 554 1116 555
rect 1142 559 1148 560
rect 1142 555 1143 559
rect 1147 555 1148 559
rect 1630 559 1631 563
rect 1635 559 1636 563
rect 1670 561 1671 565
rect 1675 561 1676 565
rect 1766 565 1767 569
rect 1771 565 1772 569
rect 1896 568 1898 642
rect 1918 624 1924 625
rect 1918 620 1919 624
rect 1923 620 1924 624
rect 1918 619 1924 620
rect 1920 615 1922 619
rect 1919 614 1923 615
rect 1919 609 1923 610
rect 2015 614 2019 615
rect 2015 609 2019 610
rect 2014 608 2020 609
rect 2014 604 2015 608
rect 2019 604 2020 608
rect 2014 603 2020 604
rect 2014 579 2020 580
rect 2014 575 2015 579
rect 2019 575 2020 579
rect 1927 574 1931 575
rect 2014 574 2020 575
rect 1926 569 1932 570
rect 2015 569 2019 570
rect 1766 564 1772 565
rect 1894 567 1900 568
rect 1894 563 1895 567
rect 1899 563 1900 567
rect 1926 565 1927 569
rect 1931 565 1932 569
rect 1926 564 1932 565
rect 2032 564 2034 642
rect 2046 624 2052 625
rect 2046 620 2047 624
rect 2051 620 2052 624
rect 2046 619 2052 620
rect 2182 624 2188 625
rect 2182 620 2183 624
rect 2187 620 2188 624
rect 2182 619 2188 620
rect 2048 615 2050 619
rect 2184 615 2186 619
rect 2047 614 2051 615
rect 2047 609 2051 610
rect 2183 614 2187 615
rect 2183 609 2187 610
rect 2182 608 2188 609
rect 2182 604 2183 608
rect 2187 604 2188 608
rect 2182 603 2188 604
rect 2192 584 2194 642
rect 2326 624 2332 625
rect 2326 620 2327 624
rect 2331 620 2332 624
rect 2326 619 2332 620
rect 2328 615 2330 619
rect 2327 614 2331 615
rect 2327 609 2331 610
rect 2359 614 2363 615
rect 2359 609 2363 610
rect 2358 608 2364 609
rect 2358 604 2359 608
rect 2363 604 2364 608
rect 2358 603 2364 604
rect 2190 583 2196 584
rect 2182 579 2188 580
rect 2182 575 2183 579
rect 2187 575 2188 579
rect 2190 579 2191 583
rect 2195 579 2196 583
rect 2190 578 2196 579
rect 2358 579 2364 580
rect 2358 575 2359 579
rect 2363 575 2364 579
rect 2414 579 2420 580
rect 2414 575 2415 579
rect 2419 575 2420 579
rect 2087 574 2091 575
rect 2182 574 2188 575
rect 2247 574 2251 575
rect 2358 574 2364 575
rect 2407 574 2411 575
rect 2414 574 2420 575
rect 2086 569 2092 570
rect 2183 569 2187 570
rect 2246 569 2252 570
rect 2359 569 2363 570
rect 2406 569 2412 570
rect 2086 565 2087 569
rect 2091 565 2092 569
rect 2086 564 2092 565
rect 2246 565 2247 569
rect 2251 565 2252 569
rect 2246 564 2252 565
rect 2406 565 2407 569
rect 2411 565 2412 569
rect 2416 568 2418 574
rect 2460 568 2462 642
rect 2470 624 2476 625
rect 2470 620 2471 624
rect 2475 620 2476 624
rect 2470 619 2476 620
rect 2614 624 2620 625
rect 2614 620 2615 624
rect 2619 620 2620 624
rect 2614 619 2620 620
rect 2758 624 2764 625
rect 2758 620 2759 624
rect 2763 620 2764 624
rect 2758 619 2764 620
rect 2472 615 2474 619
rect 2616 615 2618 619
rect 2760 615 2762 619
rect 2471 614 2475 615
rect 2471 609 2475 610
rect 2551 614 2555 615
rect 2551 609 2555 610
rect 2615 614 2619 615
rect 2615 609 2619 610
rect 2751 614 2755 615
rect 2751 609 2755 610
rect 2759 614 2763 615
rect 2759 609 2763 610
rect 2550 608 2556 609
rect 2550 604 2551 608
rect 2555 604 2556 608
rect 2550 603 2556 604
rect 2750 608 2756 609
rect 2750 604 2751 608
rect 2755 604 2756 608
rect 2750 603 2756 604
rect 2759 583 2765 584
rect 2550 579 2556 580
rect 2550 575 2551 579
rect 2555 575 2556 579
rect 2750 579 2756 580
rect 2750 575 2751 579
rect 2755 575 2756 579
rect 2759 579 2760 583
rect 2764 582 2765 583
rect 2768 582 2770 646
rect 2764 580 2770 582
rect 2764 579 2765 580
rect 2759 578 2765 579
rect 2550 574 2556 575
rect 2567 574 2571 575
rect 2750 574 2756 575
rect 2551 569 2555 570
rect 2566 569 2572 570
rect 2751 569 2755 570
rect 2406 564 2412 565
rect 2414 567 2420 568
rect 1894 562 1900 563
rect 2030 563 2036 564
rect 1670 560 1676 561
rect 1630 558 1636 559
rect 1142 554 1148 555
rect 880 543 882 554
rect 888 553 898 554
rect 879 542 883 543
rect 887 542 891 543
rect 879 537 883 538
rect 886 537 892 538
rect 774 532 780 533
rect 782 535 788 536
rect 430 530 436 531
rect 550 531 556 532
rect 310 526 316 527
rect 550 527 551 531
rect 555 527 556 531
rect 550 526 556 527
rect 670 531 676 532
rect 670 527 671 531
rect 675 527 676 531
rect 782 531 783 535
rect 787 531 788 535
rect 886 533 887 537
rect 891 533 892 537
rect 886 532 892 533
rect 896 532 898 553
rect 992 543 994 554
rect 991 542 995 543
rect 991 537 995 538
rect 1000 532 1002 554
rect 1112 543 1114 554
rect 1007 542 1011 543
rect 1111 542 1115 543
rect 1006 537 1012 538
rect 1111 537 1115 538
rect 1006 533 1007 537
rect 1011 533 1012 537
rect 1006 532 1012 533
rect 782 530 788 531
rect 826 531 832 532
rect 670 526 676 527
rect 826 527 827 531
rect 831 527 832 531
rect 826 526 832 527
rect 894 531 900 532
rect 894 527 895 531
rect 899 527 900 531
rect 894 526 900 527
rect 998 531 1004 532
rect 998 527 999 531
rect 1003 527 1004 531
rect 998 526 1004 527
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 110 510 116 511
rect 112 491 114 510
rect 111 490 115 491
rect 111 485 115 486
rect 135 490 139 491
rect 135 485 139 486
rect 112 478 114 485
rect 134 484 140 485
rect 134 480 135 484
rect 139 480 140 484
rect 134 479 140 480
rect 110 477 116 478
rect 110 473 111 477
rect 115 473 116 477
rect 110 472 116 473
rect 148 460 150 526
rect 174 508 180 509
rect 174 504 175 508
rect 179 504 180 508
rect 174 503 180 504
rect 302 508 308 509
rect 302 504 303 508
rect 307 504 308 508
rect 302 503 308 504
rect 422 508 428 509
rect 422 504 423 508
rect 427 504 428 508
rect 422 503 428 504
rect 542 508 548 509
rect 542 504 543 508
rect 547 504 548 508
rect 542 503 548 504
rect 662 508 668 509
rect 662 504 663 508
rect 667 504 668 508
rect 662 503 668 504
rect 176 491 178 503
rect 304 491 306 503
rect 424 491 426 503
rect 544 491 546 503
rect 664 491 666 503
rect 175 490 179 491
rect 175 485 179 486
rect 231 490 235 491
rect 231 485 235 486
rect 303 490 307 491
rect 303 485 307 486
rect 359 490 363 491
rect 359 485 363 486
rect 423 490 427 491
rect 423 485 427 486
rect 503 490 507 491
rect 503 485 507 486
rect 543 490 547 491
rect 543 485 547 486
rect 655 490 659 491
rect 655 485 659 486
rect 663 490 667 491
rect 663 485 667 486
rect 230 484 236 485
rect 230 480 231 484
rect 235 480 236 484
rect 230 479 236 480
rect 358 484 364 485
rect 358 480 359 484
rect 363 480 364 484
rect 358 479 364 480
rect 502 484 508 485
rect 502 480 503 484
rect 507 480 508 484
rect 502 479 508 480
rect 654 484 660 485
rect 654 480 655 484
rect 659 480 660 484
rect 672 483 674 526
rect 774 508 780 509
rect 774 504 775 508
rect 779 504 780 508
rect 774 503 780 504
rect 776 491 778 503
rect 775 490 779 491
rect 775 485 779 486
rect 815 490 819 491
rect 815 485 819 486
rect 654 479 660 480
rect 664 481 674 483
rect 814 484 820 485
rect 470 463 476 464
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 146 459 152 460
rect 110 454 116 455
rect 134 455 140 456
rect 112 439 114 454
rect 134 451 135 455
rect 139 451 140 455
rect 146 455 147 459
rect 151 455 152 459
rect 470 459 471 463
rect 475 459 476 463
rect 470 458 476 459
rect 146 454 152 455
rect 230 455 236 456
rect 134 450 140 451
rect 230 451 231 455
rect 235 451 236 455
rect 230 450 236 451
rect 358 455 364 456
rect 358 451 359 455
rect 363 451 364 455
rect 358 450 364 451
rect 136 439 138 450
rect 232 439 234 450
rect 360 439 362 450
rect 111 438 115 439
rect 111 433 115 434
rect 135 438 139 439
rect 135 433 139 434
rect 231 438 235 439
rect 231 433 235 434
rect 359 438 363 439
rect 359 433 363 434
rect 112 430 114 433
rect 110 429 116 430
rect 110 425 111 429
rect 115 425 116 429
rect 110 424 116 425
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 110 406 116 407
rect 112 391 114 406
rect 111 390 115 391
rect 111 385 115 386
rect 112 378 114 385
rect 110 377 116 378
rect 110 373 111 377
rect 115 373 116 377
rect 110 372 116 373
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 110 354 116 355
rect 112 347 114 354
rect 111 346 115 347
rect 111 341 115 342
rect 112 338 114 341
rect 110 337 116 338
rect 110 333 111 337
rect 115 333 116 337
rect 110 332 116 333
rect 110 319 116 320
rect 110 315 111 319
rect 115 315 116 319
rect 110 314 116 315
rect 112 303 114 314
rect 111 302 115 303
rect 111 297 115 298
rect 463 302 467 303
rect 463 297 467 298
rect 112 290 114 297
rect 462 296 468 297
rect 462 292 463 296
rect 467 292 468 296
rect 462 291 468 292
rect 110 289 116 290
rect 110 285 111 289
rect 115 285 116 289
rect 110 284 116 285
rect 472 272 474 458
rect 664 456 666 481
rect 814 480 815 484
rect 819 480 820 484
rect 814 479 820 480
rect 828 456 830 526
rect 886 508 892 509
rect 886 504 887 508
rect 891 504 892 508
rect 886 503 892 504
rect 1006 508 1012 509
rect 1006 504 1007 508
rect 1011 504 1012 508
rect 1006 503 1012 504
rect 888 491 890 503
rect 1008 491 1010 503
rect 887 490 891 491
rect 887 485 891 486
rect 975 490 979 491
rect 975 485 979 486
rect 1007 490 1011 491
rect 1007 485 1011 486
rect 1135 490 1139 491
rect 1135 485 1139 486
rect 974 484 980 485
rect 974 480 975 484
rect 979 480 980 484
rect 974 479 980 480
rect 1134 484 1140 485
rect 1134 480 1135 484
rect 1139 480 1140 484
rect 1134 479 1140 480
rect 1144 460 1146 554
rect 1632 543 1634 558
rect 1670 547 1676 548
rect 1670 543 1671 547
rect 1675 543 1676 547
rect 1631 542 1635 543
rect 1670 542 1676 543
rect 1631 537 1635 538
rect 1632 534 1634 537
rect 1672 535 1674 542
rect 1766 540 1772 541
rect 1766 536 1767 540
rect 1771 536 1772 540
rect 1766 535 1772 536
rect 1671 534 1675 535
rect 1630 533 1636 534
rect 1630 529 1631 533
rect 1635 529 1636 533
rect 1671 529 1675 530
rect 1695 534 1699 535
rect 1695 529 1699 530
rect 1767 534 1771 535
rect 1767 529 1771 530
rect 1887 534 1891 535
rect 1887 529 1891 530
rect 1630 528 1636 529
rect 1672 522 1674 529
rect 1694 528 1700 529
rect 1694 524 1695 528
rect 1699 524 1700 528
rect 1694 523 1700 524
rect 1886 528 1892 529
rect 1886 524 1887 528
rect 1891 524 1892 528
rect 1886 523 1892 524
rect 1670 521 1676 522
rect 1670 517 1671 521
rect 1675 517 1676 521
rect 1670 516 1676 517
rect 1630 515 1636 516
rect 1630 511 1631 515
rect 1635 511 1636 515
rect 1630 510 1636 511
rect 1632 491 1634 510
rect 1896 504 1898 562
rect 2030 559 2031 563
rect 2035 559 2036 563
rect 2030 558 2036 559
rect 2110 563 2116 564
rect 2110 559 2111 563
rect 2115 559 2116 563
rect 2414 563 2415 567
rect 2419 563 2420 567
rect 2414 562 2420 563
rect 2458 567 2464 568
rect 2458 563 2459 567
rect 2463 563 2464 567
rect 2566 565 2567 569
rect 2571 565 2572 569
rect 2566 564 2572 565
rect 2458 562 2464 563
rect 2606 563 2612 564
rect 2110 558 2116 559
rect 1926 540 1932 541
rect 1926 536 1927 540
rect 1931 536 1932 540
rect 1926 535 1932 536
rect 1927 534 1931 535
rect 1927 529 1931 530
rect 1670 503 1676 504
rect 1670 499 1671 503
rect 1675 499 1676 503
rect 1894 503 1900 504
rect 1670 498 1676 499
rect 1694 499 1700 500
rect 1295 490 1299 491
rect 1295 485 1299 486
rect 1455 490 1459 491
rect 1455 485 1459 486
rect 1599 490 1603 491
rect 1599 485 1603 486
rect 1631 490 1635 491
rect 1672 487 1674 498
rect 1694 495 1695 499
rect 1699 495 1700 499
rect 1694 494 1700 495
rect 1702 499 1708 500
rect 1702 495 1703 499
rect 1707 495 1708 499
rect 1702 494 1708 495
rect 1886 499 1892 500
rect 1886 495 1887 499
rect 1891 495 1892 499
rect 1894 499 1895 503
rect 1899 499 1900 503
rect 1894 498 1900 499
rect 1886 494 1892 495
rect 1696 487 1698 494
rect 1631 485 1635 486
rect 1671 486 1675 487
rect 1294 484 1300 485
rect 1294 480 1295 484
rect 1299 480 1300 484
rect 1294 479 1300 480
rect 1454 484 1460 485
rect 1454 480 1455 484
rect 1459 480 1460 484
rect 1454 479 1460 480
rect 1598 484 1604 485
rect 1598 480 1599 484
rect 1603 480 1604 484
rect 1598 479 1604 480
rect 1632 478 1634 485
rect 1695 486 1699 487
rect 1671 481 1675 482
rect 1694 481 1700 482
rect 1672 478 1674 481
rect 1630 477 1636 478
rect 1630 473 1631 477
rect 1635 473 1636 477
rect 1630 472 1636 473
rect 1670 477 1676 478
rect 1670 473 1671 477
rect 1675 473 1676 477
rect 1694 477 1695 481
rect 1699 477 1700 481
rect 1704 480 1706 494
rect 1888 487 1890 494
rect 1887 486 1891 487
rect 2023 486 2027 487
rect 1887 481 1891 482
rect 2022 481 2028 482
rect 1694 476 1700 477
rect 1702 479 1708 480
rect 1702 475 1703 479
rect 1707 475 1708 479
rect 2022 477 2023 481
rect 2027 477 2028 481
rect 2032 480 2034 558
rect 2086 540 2092 541
rect 2086 536 2087 540
rect 2091 536 2092 540
rect 2086 535 2092 536
rect 2087 534 2091 535
rect 2087 529 2091 530
rect 2103 534 2107 535
rect 2103 529 2107 530
rect 2102 528 2108 529
rect 2102 524 2103 528
rect 2107 524 2108 528
rect 2102 523 2108 524
rect 2112 504 2114 558
rect 2246 540 2252 541
rect 2246 536 2247 540
rect 2251 536 2252 540
rect 2246 535 2252 536
rect 2406 540 2412 541
rect 2406 536 2407 540
rect 2411 536 2412 540
rect 2406 535 2412 536
rect 2247 534 2251 535
rect 2247 529 2251 530
rect 2343 534 2347 535
rect 2343 529 2347 530
rect 2407 534 2411 535
rect 2407 529 2411 530
rect 2342 528 2348 529
rect 2342 524 2343 528
rect 2347 524 2348 528
rect 2342 523 2348 524
rect 2416 504 2418 562
rect 2606 559 2607 563
rect 2611 559 2612 563
rect 2606 558 2612 559
rect 2566 540 2572 541
rect 2566 536 2567 540
rect 2571 536 2572 540
rect 2566 535 2572 536
rect 2567 534 2571 535
rect 2567 529 2571 530
rect 2599 534 2603 535
rect 2599 529 2603 530
rect 2598 528 2604 529
rect 2598 524 2599 528
rect 2603 524 2604 528
rect 2598 523 2604 524
rect 2110 503 2116 504
rect 2102 499 2108 500
rect 2102 495 2103 499
rect 2107 495 2108 499
rect 2110 499 2111 503
rect 2115 499 2116 503
rect 2414 503 2420 504
rect 2110 498 2116 499
rect 2342 499 2348 500
rect 2102 494 2108 495
rect 2342 495 2343 499
rect 2347 495 2348 499
rect 2414 499 2415 503
rect 2419 499 2420 503
rect 2608 500 2610 558
rect 2863 534 2867 535
rect 2863 529 2867 530
rect 2862 528 2868 529
rect 2862 524 2863 528
rect 2867 524 2868 528
rect 2862 523 2868 524
rect 2872 500 2874 666
rect 2992 659 2994 666
rect 3160 659 3162 666
rect 2991 658 2995 659
rect 2991 653 2995 654
rect 3159 658 3163 659
rect 3159 653 3163 654
rect 2959 614 2963 615
rect 2959 609 2963 610
rect 3159 614 3163 615
rect 3159 609 3163 610
rect 2958 608 2964 609
rect 2958 604 2959 608
rect 2963 604 2964 608
rect 2958 603 2964 604
rect 3158 608 3164 609
rect 3158 604 3159 608
rect 3163 604 3164 608
rect 3158 603 3164 604
rect 3168 584 3170 670
rect 3192 659 3194 670
rect 3191 658 3195 659
rect 3191 653 3195 654
rect 3192 650 3194 653
rect 3190 649 3196 650
rect 3190 645 3191 649
rect 3195 645 3196 649
rect 3190 644 3196 645
rect 3190 631 3196 632
rect 3190 627 3191 631
rect 3195 627 3196 631
rect 3190 626 3196 627
rect 3192 615 3194 626
rect 3191 614 3195 615
rect 3191 609 3195 610
rect 3192 602 3194 609
rect 3190 601 3196 602
rect 3190 597 3191 601
rect 3195 597 3196 601
rect 3190 596 3196 597
rect 3166 583 3172 584
rect 2958 579 2964 580
rect 2958 575 2959 579
rect 2963 575 2964 579
rect 2958 574 2964 575
rect 3158 579 3164 580
rect 3158 575 3159 579
rect 3163 575 3164 579
rect 3166 579 3167 583
rect 3171 579 3172 583
rect 3166 578 3172 579
rect 3190 583 3196 584
rect 3190 579 3191 583
rect 3195 579 3196 583
rect 3190 578 3196 579
rect 3158 574 3164 575
rect 2959 569 2963 570
rect 3159 569 3163 570
rect 3135 534 3139 535
rect 3135 529 3139 530
rect 3134 528 3140 529
rect 3134 524 3135 528
rect 3139 524 3140 528
rect 3134 523 3140 524
rect 3168 504 3170 578
rect 3192 575 3194 578
rect 3191 574 3195 575
rect 3191 569 3195 570
rect 3192 566 3194 569
rect 3190 565 3196 566
rect 3190 561 3191 565
rect 3195 561 3196 565
rect 3190 560 3196 561
rect 3190 547 3196 548
rect 3190 543 3191 547
rect 3195 543 3196 547
rect 3190 542 3196 543
rect 3192 535 3194 542
rect 3191 534 3195 535
rect 3191 529 3195 530
rect 3192 522 3194 529
rect 3190 521 3196 522
rect 3190 517 3191 521
rect 3195 517 3196 521
rect 3190 516 3196 517
rect 3142 503 3148 504
rect 2414 498 2420 499
rect 2598 499 2604 500
rect 2342 494 2348 495
rect 2104 487 2106 494
rect 2344 487 2346 494
rect 2103 486 2107 487
rect 2103 481 2107 482
rect 2343 486 2347 487
rect 2383 486 2387 487
rect 2343 481 2347 482
rect 2382 481 2388 482
rect 2022 476 2028 477
rect 2030 479 2036 480
rect 1702 474 1708 475
rect 2030 475 2031 479
rect 2035 475 2036 479
rect 2030 474 2036 475
rect 2058 479 2064 480
rect 2058 475 2059 479
rect 2063 475 2064 479
rect 2382 477 2383 481
rect 2387 477 2388 481
rect 2416 480 2418 498
rect 2598 495 2599 499
rect 2603 495 2604 499
rect 2598 494 2604 495
rect 2606 499 2612 500
rect 2606 495 2607 499
rect 2611 495 2612 499
rect 2606 494 2612 495
rect 2630 499 2636 500
rect 2630 495 2631 499
rect 2635 495 2636 499
rect 2630 494 2636 495
rect 2862 499 2868 500
rect 2862 495 2863 499
rect 2867 495 2868 499
rect 2862 494 2868 495
rect 2870 499 2876 500
rect 2870 495 2871 499
rect 2875 495 2876 499
rect 2870 494 2876 495
rect 2926 499 2932 500
rect 2926 495 2927 499
rect 2931 495 2932 499
rect 2926 494 2932 495
rect 3134 499 3140 500
rect 3134 495 3135 499
rect 3139 495 3140 499
rect 3142 499 3143 503
rect 3147 499 3148 503
rect 3142 498 3148 499
rect 3166 503 3172 504
rect 3166 499 3167 503
rect 3171 499 3172 503
rect 3166 498 3172 499
rect 3190 503 3196 504
rect 3190 499 3191 503
rect 3195 499 3196 503
rect 3190 498 3196 499
rect 3134 494 3140 495
rect 2600 487 2602 494
rect 2599 486 2603 487
rect 2599 481 2603 482
rect 2382 476 2388 477
rect 2414 479 2420 480
rect 2058 474 2064 475
rect 2414 475 2415 479
rect 2419 475 2420 479
rect 2414 474 2420 475
rect 1670 472 1676 473
rect 1704 468 1706 474
rect 1606 467 1612 468
rect 1606 463 1607 467
rect 1611 463 1612 467
rect 1606 462 1612 463
rect 1702 467 1708 468
rect 1702 463 1703 467
rect 1707 463 1708 467
rect 1702 462 1708 463
rect 1142 459 1148 460
rect 502 455 508 456
rect 502 451 503 455
rect 507 451 508 455
rect 502 450 508 451
rect 654 455 660 456
rect 654 451 655 455
rect 659 451 660 455
rect 654 450 660 451
rect 662 455 668 456
rect 662 451 663 455
rect 667 451 668 455
rect 662 450 668 451
rect 814 455 820 456
rect 814 451 815 455
rect 819 451 820 455
rect 814 450 820 451
rect 826 455 832 456
rect 826 451 827 455
rect 831 451 832 455
rect 826 450 832 451
rect 974 455 980 456
rect 974 451 975 455
rect 979 451 980 455
rect 974 450 980 451
rect 982 455 988 456
rect 982 451 983 455
rect 987 451 988 455
rect 1134 455 1140 456
rect 1134 451 1135 455
rect 1139 451 1140 455
rect 1142 455 1143 459
rect 1147 455 1148 459
rect 1608 456 1610 462
rect 1630 459 1636 460
rect 1142 454 1148 455
rect 1294 455 1300 456
rect 982 450 994 451
rect 1134 450 1140 451
rect 504 439 506 450
rect 656 439 658 450
rect 503 438 507 439
rect 503 433 507 434
rect 655 438 659 439
rect 655 433 659 434
rect 664 427 666 450
rect 816 439 818 450
rect 727 438 731 439
rect 815 438 819 439
rect 726 433 732 434
rect 815 433 819 434
rect 726 429 727 433
rect 731 429 732 433
rect 726 428 732 429
rect 828 428 830 450
rect 976 439 978 450
rect 984 449 994 450
rect 855 438 859 439
rect 975 438 979 439
rect 983 438 987 439
rect 854 433 860 434
rect 975 433 979 434
rect 982 433 988 434
rect 854 429 855 433
rect 859 429 860 433
rect 854 428 860 429
rect 982 429 983 433
rect 987 429 988 433
rect 982 428 988 429
rect 992 428 994 449
rect 1136 439 1138 450
rect 1144 440 1146 454
rect 1294 451 1295 455
rect 1299 451 1300 455
rect 1294 450 1300 451
rect 1342 455 1348 456
rect 1342 451 1343 455
rect 1347 451 1348 455
rect 1342 450 1348 451
rect 1454 455 1460 456
rect 1454 451 1455 455
rect 1459 451 1460 455
rect 1454 450 1460 451
rect 1466 455 1472 456
rect 1466 451 1467 455
rect 1471 451 1472 455
rect 1466 450 1472 451
rect 1598 455 1604 456
rect 1598 451 1599 455
rect 1603 451 1604 455
rect 1598 450 1604 451
rect 1606 455 1612 456
rect 1606 451 1607 455
rect 1611 451 1612 455
rect 1630 455 1631 459
rect 1635 455 1636 459
rect 1630 454 1636 455
rect 1670 459 1676 460
rect 1670 455 1671 459
rect 1675 455 1676 459
rect 1670 454 1676 455
rect 1606 450 1612 451
rect 1142 439 1148 440
rect 1230 439 1236 440
rect 1296 439 1298 450
rect 1103 438 1107 439
rect 1135 438 1139 439
rect 1142 435 1143 439
rect 1147 435 1148 439
rect 1142 434 1148 435
rect 1223 438 1227 439
rect 1230 435 1231 439
rect 1235 435 1236 439
rect 1230 434 1236 435
rect 1295 438 1299 439
rect 1335 438 1339 439
rect 1102 433 1108 434
rect 1135 433 1139 434
rect 1102 429 1103 433
rect 1107 429 1108 433
rect 1144 432 1146 434
rect 1222 433 1228 434
rect 1102 428 1108 429
rect 1142 431 1148 432
rect 660 425 666 427
rect 814 427 820 428
rect 647 390 651 391
rect 647 385 651 386
rect 646 384 652 385
rect 646 380 647 384
rect 651 380 652 384
rect 646 379 652 380
rect 660 360 662 425
rect 814 423 815 427
rect 819 423 820 427
rect 814 422 820 423
rect 826 427 832 428
rect 826 423 827 427
rect 831 423 832 427
rect 826 422 832 423
rect 990 427 996 428
rect 990 423 991 427
rect 995 423 996 427
rect 1142 427 1143 431
rect 1147 427 1148 431
rect 1222 429 1223 433
rect 1227 429 1228 433
rect 1232 432 1234 434
rect 1295 433 1299 434
rect 1334 433 1340 434
rect 1222 428 1228 429
rect 1230 431 1236 432
rect 1142 426 1148 427
rect 1230 427 1231 431
rect 1235 427 1236 431
rect 1334 429 1335 433
rect 1339 429 1340 433
rect 1334 428 1340 429
rect 1344 428 1346 450
rect 1456 439 1458 450
rect 1468 440 1470 450
rect 1466 439 1472 440
rect 1600 439 1602 450
rect 1608 440 1610 450
rect 1606 439 1612 440
rect 1632 439 1634 454
rect 1672 443 1674 454
rect 1694 452 1700 453
rect 1694 448 1695 452
rect 1699 448 1700 452
rect 1694 447 1700 448
rect 2022 452 2028 453
rect 2022 448 2023 452
rect 2027 448 2028 452
rect 2022 447 2028 448
rect 1696 443 1698 447
rect 2024 443 2026 447
rect 1671 442 1675 443
rect 1447 438 1451 439
rect 1455 438 1459 439
rect 1466 435 1467 439
rect 1471 435 1472 439
rect 1466 434 1472 435
rect 1567 438 1571 439
rect 1599 438 1603 439
rect 1606 435 1607 439
rect 1611 435 1612 439
rect 1606 434 1612 435
rect 1631 438 1635 439
rect 1671 437 1675 438
rect 1695 442 1699 443
rect 1695 437 1699 438
rect 2023 442 2027 443
rect 2023 437 2027 438
rect 1446 433 1452 434
rect 1455 433 1459 434
rect 1446 429 1447 433
rect 1451 429 1452 433
rect 1468 432 1470 434
rect 1566 433 1572 434
rect 1599 433 1603 434
rect 1446 428 1452 429
rect 1466 431 1472 432
rect 1230 426 1236 427
rect 1342 427 1348 428
rect 990 422 996 423
rect 1342 423 1343 427
rect 1347 423 1348 427
rect 1466 427 1467 431
rect 1471 427 1472 431
rect 1566 429 1567 433
rect 1571 429 1572 433
rect 1608 432 1610 434
rect 1631 433 1635 434
rect 1566 428 1572 429
rect 1606 431 1612 432
rect 1466 426 1472 427
rect 1606 427 1607 431
rect 1611 427 1612 431
rect 1632 430 1634 433
rect 1672 430 1674 437
rect 1606 426 1612 427
rect 1630 429 1636 430
rect 1342 422 1348 423
rect 726 404 732 405
rect 726 400 727 404
rect 731 400 732 404
rect 726 399 732 400
rect 728 391 730 399
rect 727 390 731 391
rect 727 385 731 386
rect 807 390 811 391
rect 807 385 811 386
rect 806 384 812 385
rect 806 380 807 384
rect 811 380 812 384
rect 806 379 812 380
rect 654 359 662 360
rect 646 355 652 356
rect 646 351 647 355
rect 651 351 652 355
rect 654 355 655 359
rect 659 356 662 359
rect 816 356 818 422
rect 854 404 860 405
rect 854 400 855 404
rect 859 400 860 404
rect 854 399 860 400
rect 982 404 988 405
rect 982 400 983 404
rect 987 400 988 404
rect 982 399 988 400
rect 856 391 858 399
rect 984 391 986 399
rect 855 390 859 391
rect 855 385 859 386
rect 951 390 955 391
rect 951 385 955 386
rect 983 390 987 391
rect 983 385 987 386
rect 950 384 956 385
rect 950 380 951 384
rect 955 380 956 384
rect 950 379 956 380
rect 992 356 994 422
rect 1102 404 1108 405
rect 1102 400 1103 404
rect 1107 400 1108 404
rect 1102 399 1108 400
rect 1222 404 1228 405
rect 1222 400 1223 404
rect 1227 400 1228 404
rect 1222 399 1228 400
rect 1334 404 1340 405
rect 1334 400 1335 404
rect 1339 400 1340 404
rect 1334 399 1340 400
rect 1104 391 1106 399
rect 1224 391 1226 399
rect 1336 391 1338 399
rect 1087 390 1091 391
rect 1087 385 1091 386
rect 1103 390 1107 391
rect 1103 385 1107 386
rect 1215 390 1219 391
rect 1215 385 1219 386
rect 1223 390 1227 391
rect 1223 385 1227 386
rect 1335 390 1339 391
rect 1335 385 1339 386
rect 1086 384 1092 385
rect 1086 380 1087 384
rect 1091 380 1092 384
rect 1086 379 1092 380
rect 1214 384 1220 385
rect 1214 380 1215 384
rect 1219 380 1220 384
rect 1214 379 1220 380
rect 1334 384 1340 385
rect 1334 380 1335 384
rect 1339 380 1340 384
rect 1334 379 1340 380
rect 1344 356 1346 422
rect 1446 404 1452 405
rect 1446 400 1447 404
rect 1451 400 1452 404
rect 1446 399 1452 400
rect 1448 391 1450 399
rect 1468 395 1470 426
rect 1630 425 1631 429
rect 1635 425 1636 429
rect 1630 424 1636 425
rect 1670 429 1676 430
rect 1670 425 1671 429
rect 1675 425 1676 429
rect 1670 424 1676 425
rect 1630 411 1636 412
rect 1630 407 1631 411
rect 1635 407 1636 411
rect 1630 406 1636 407
rect 1670 411 1676 412
rect 1670 407 1671 411
rect 1675 407 1676 411
rect 1670 406 1676 407
rect 1566 404 1572 405
rect 1566 400 1567 404
rect 1571 400 1572 404
rect 1566 399 1572 400
rect 1468 393 1474 395
rect 1447 390 1451 391
rect 1447 385 1451 386
rect 1463 390 1467 391
rect 1463 385 1467 386
rect 1462 384 1468 385
rect 1462 380 1463 384
rect 1467 380 1468 384
rect 1462 379 1468 380
rect 1472 360 1474 393
rect 1568 391 1570 399
rect 1632 391 1634 406
rect 1672 391 1674 406
rect 1567 390 1571 391
rect 1567 385 1571 386
rect 1631 390 1635 391
rect 1631 385 1635 386
rect 1671 390 1675 391
rect 1671 385 1675 386
rect 1632 378 1634 385
rect 1672 382 1674 385
rect 1670 381 1676 382
rect 1630 377 1636 378
rect 1630 373 1631 377
rect 1635 373 1636 377
rect 1670 377 1671 381
rect 1675 377 1676 381
rect 1670 376 1676 377
rect 1630 372 1636 373
rect 1670 363 1676 364
rect 1470 359 1476 360
rect 659 355 660 356
rect 654 354 660 355
rect 806 355 812 356
rect 646 350 652 351
rect 648 347 650 350
rect 543 346 547 347
rect 647 346 651 347
rect 542 341 548 342
rect 647 341 651 342
rect 542 337 543 341
rect 547 337 548 341
rect 542 336 548 337
rect 656 336 658 354
rect 806 351 807 355
rect 811 351 812 355
rect 806 350 812 351
rect 814 355 820 356
rect 814 351 815 355
rect 819 351 820 355
rect 814 350 820 351
rect 950 355 956 356
rect 950 351 951 355
rect 955 351 956 355
rect 950 350 956 351
rect 990 355 996 356
rect 990 351 991 355
rect 995 351 996 355
rect 990 350 996 351
rect 1086 355 1092 356
rect 1086 351 1087 355
rect 1091 351 1092 355
rect 1086 350 1092 351
rect 1214 355 1220 356
rect 1214 351 1215 355
rect 1219 351 1220 355
rect 1214 350 1220 351
rect 1334 355 1340 356
rect 1334 351 1335 355
rect 1339 351 1340 355
rect 1334 350 1340 351
rect 1342 355 1348 356
rect 1342 351 1343 355
rect 1347 351 1348 355
rect 1342 350 1348 351
rect 1462 355 1468 356
rect 1462 351 1463 355
rect 1467 351 1468 355
rect 1470 355 1471 359
rect 1475 355 1476 359
rect 1470 354 1476 355
rect 1630 359 1636 360
rect 1630 355 1631 359
rect 1635 355 1636 359
rect 1670 359 1671 363
rect 1675 359 1676 363
rect 1670 358 1676 359
rect 1630 354 1636 355
rect 1462 350 1468 351
rect 808 347 810 350
rect 671 346 675 347
rect 807 346 811 347
rect 670 341 676 342
rect 670 337 671 341
rect 675 337 676 341
rect 670 336 676 337
rect 806 341 812 342
rect 806 337 807 341
rect 811 337 812 341
rect 806 336 812 337
rect 816 336 818 350
rect 952 347 954 350
rect 1088 347 1090 350
rect 1216 347 1218 350
rect 1336 347 1338 350
rect 943 346 947 347
rect 951 346 955 347
rect 1079 346 1083 347
rect 1087 346 1091 347
rect 942 341 948 342
rect 951 341 955 342
rect 1078 341 1084 342
rect 1087 341 1091 342
rect 1215 346 1219 347
rect 1223 346 1227 347
rect 1335 346 1339 347
rect 1215 341 1219 342
rect 1222 341 1228 342
rect 1335 341 1339 342
rect 942 337 943 341
rect 947 337 948 341
rect 942 336 948 337
rect 1078 337 1079 341
rect 1083 337 1084 341
rect 1078 336 1084 337
rect 1222 337 1223 341
rect 1227 337 1228 341
rect 1344 340 1346 350
rect 1464 347 1466 350
rect 1367 346 1371 347
rect 1463 346 1467 347
rect 1366 341 1372 342
rect 1463 341 1467 342
rect 1222 336 1228 337
rect 1294 339 1300 340
rect 630 335 636 336
rect 630 331 631 335
rect 635 331 636 335
rect 630 330 636 331
rect 654 335 660 336
rect 654 331 655 335
rect 659 331 660 335
rect 654 330 660 331
rect 814 335 820 336
rect 814 331 815 335
rect 819 331 820 335
rect 1294 335 1295 339
rect 1299 335 1300 339
rect 1294 334 1300 335
rect 1342 339 1348 340
rect 1342 335 1343 339
rect 1347 335 1348 339
rect 1366 337 1367 341
rect 1371 337 1372 341
rect 1472 340 1474 354
rect 1632 347 1634 354
rect 1631 346 1635 347
rect 1631 341 1635 342
rect 1366 336 1372 337
rect 1470 339 1476 340
rect 1342 334 1348 335
rect 1470 335 1471 339
rect 1475 335 1476 339
rect 1632 338 1634 341
rect 1672 339 1674 358
rect 1671 338 1675 339
rect 1470 334 1476 335
rect 1630 337 1636 338
rect 814 330 820 331
rect 542 312 548 313
rect 542 308 543 312
rect 547 308 548 312
rect 542 307 548 308
rect 544 303 546 307
rect 543 302 547 303
rect 543 297 547 298
rect 623 302 627 303
rect 623 297 627 298
rect 622 296 628 297
rect 622 292 623 296
rect 627 292 628 296
rect 622 291 628 292
rect 110 271 116 272
rect 110 267 111 271
rect 115 267 116 271
rect 470 271 476 272
rect 110 266 116 267
rect 462 267 468 268
rect 112 259 114 266
rect 462 263 463 267
rect 467 263 468 267
rect 470 267 471 271
rect 475 267 476 271
rect 632 268 634 330
rect 670 312 676 313
rect 670 308 671 312
rect 675 308 676 312
rect 670 307 676 308
rect 806 312 812 313
rect 806 308 807 312
rect 811 308 812 312
rect 806 307 812 308
rect 672 303 674 307
rect 808 303 810 307
rect 671 302 675 303
rect 671 297 675 298
rect 767 302 771 303
rect 767 297 771 298
rect 807 302 811 303
rect 807 297 811 298
rect 766 296 772 297
rect 766 292 767 296
rect 771 292 772 296
rect 766 291 772 292
rect 816 272 818 330
rect 942 312 948 313
rect 942 308 943 312
rect 947 308 948 312
rect 942 307 948 308
rect 1078 312 1084 313
rect 1078 308 1079 312
rect 1083 308 1084 312
rect 1078 307 1084 308
rect 1222 312 1228 313
rect 1222 308 1223 312
rect 1227 308 1228 312
rect 1222 307 1228 308
rect 944 303 946 307
rect 1080 303 1082 307
rect 1224 303 1226 307
rect 903 302 907 303
rect 903 297 907 298
rect 943 302 947 303
rect 943 297 947 298
rect 1031 302 1035 303
rect 1031 297 1035 298
rect 1079 302 1083 303
rect 1079 297 1083 298
rect 1159 302 1163 303
rect 1159 297 1163 298
rect 1223 302 1227 303
rect 1223 297 1227 298
rect 1287 302 1291 303
rect 1287 297 1291 298
rect 902 296 908 297
rect 902 292 903 296
rect 907 292 908 296
rect 902 291 908 292
rect 1030 296 1036 297
rect 1030 292 1031 296
rect 1035 292 1036 296
rect 1030 291 1036 292
rect 1158 296 1164 297
rect 1158 292 1159 296
rect 1163 292 1164 296
rect 1158 291 1164 292
rect 1286 296 1292 297
rect 1286 292 1287 296
rect 1291 292 1292 296
rect 1286 291 1292 292
rect 1296 272 1298 334
rect 1630 333 1631 337
rect 1635 333 1636 337
rect 1671 333 1675 334
rect 2047 338 2051 339
rect 2047 333 2051 334
rect 1630 332 1636 333
rect 1672 326 1674 333
rect 2046 332 2052 333
rect 2046 328 2047 332
rect 2051 328 2052 332
rect 2046 327 2052 328
rect 1670 325 1676 326
rect 1670 321 1671 325
rect 1675 321 1676 325
rect 1670 320 1676 321
rect 1630 319 1636 320
rect 1630 315 1631 319
rect 1635 315 1636 319
rect 1630 314 1636 315
rect 1366 312 1372 313
rect 1366 308 1367 312
rect 1371 308 1372 312
rect 1366 307 1372 308
rect 1368 303 1370 307
rect 1632 303 1634 314
rect 1670 307 1676 308
rect 1670 303 1671 307
rect 1675 303 1676 307
rect 2060 304 2062 474
rect 2382 452 2388 453
rect 2382 448 2383 452
rect 2387 448 2388 452
rect 2382 447 2388 448
rect 2384 443 2386 447
rect 2247 442 2251 443
rect 2247 437 2251 438
rect 2375 442 2379 443
rect 2375 437 2379 438
rect 2383 442 2387 443
rect 2383 437 2387 438
rect 2503 442 2507 443
rect 2503 437 2507 438
rect 2623 442 2627 443
rect 2623 437 2627 438
rect 2246 436 2252 437
rect 2246 432 2247 436
rect 2251 432 2252 436
rect 2246 431 2252 432
rect 2374 436 2380 437
rect 2374 432 2375 436
rect 2379 432 2380 436
rect 2374 431 2380 432
rect 2502 436 2508 437
rect 2502 432 2503 436
rect 2507 432 2508 436
rect 2502 431 2508 432
rect 2622 436 2628 437
rect 2622 432 2623 436
rect 2627 432 2628 436
rect 2622 431 2628 432
rect 2632 408 2634 494
rect 2864 487 2866 494
rect 2743 486 2747 487
rect 2863 486 2867 487
rect 2742 481 2748 482
rect 2863 481 2867 482
rect 2742 477 2743 481
rect 2747 477 2748 481
rect 2742 476 2748 477
rect 2750 475 2756 476
rect 2750 471 2751 475
rect 2755 471 2756 475
rect 2750 470 2756 471
rect 2742 452 2748 453
rect 2742 448 2743 452
rect 2747 448 2748 452
rect 2742 447 2748 448
rect 2744 443 2746 447
rect 2743 442 2747 443
rect 2743 437 2747 438
rect 2742 436 2748 437
rect 2742 432 2743 436
rect 2747 432 2748 436
rect 2742 431 2748 432
rect 2752 408 2754 470
rect 2855 442 2859 443
rect 2855 437 2859 438
rect 2854 436 2860 437
rect 2854 432 2855 436
rect 2859 432 2860 436
rect 2854 431 2860 432
rect 2928 412 2930 494
rect 3136 487 3138 494
rect 3111 486 3115 487
rect 3135 486 3139 487
rect 3110 481 3116 482
rect 3135 481 3139 482
rect 3110 477 3111 481
rect 3115 477 3116 481
rect 3144 480 3146 498
rect 3192 487 3194 498
rect 3191 486 3195 487
rect 3191 481 3195 482
rect 3110 476 3116 477
rect 3118 479 3124 480
rect 3118 475 3119 479
rect 3123 475 3124 479
rect 3118 474 3124 475
rect 3142 479 3148 480
rect 3142 475 3143 479
rect 3147 475 3148 479
rect 3192 478 3194 481
rect 3142 474 3148 475
rect 3190 477 3196 478
rect 3110 452 3116 453
rect 3110 448 3111 452
rect 3115 448 3116 452
rect 3110 447 3116 448
rect 3112 443 3114 447
rect 2967 442 2971 443
rect 2967 437 2971 438
rect 3087 442 3091 443
rect 3087 437 3091 438
rect 3111 442 3115 443
rect 3111 437 3115 438
rect 2966 436 2972 437
rect 2966 432 2967 436
rect 2971 432 2972 436
rect 2966 431 2972 432
rect 3086 436 3092 437
rect 3086 432 3087 436
rect 3091 432 3092 436
rect 3086 431 3092 432
rect 3120 412 3122 474
rect 3190 473 3191 477
rect 3195 473 3196 477
rect 3190 472 3196 473
rect 3190 459 3196 460
rect 3190 455 3191 459
rect 3195 455 3196 459
rect 3190 454 3196 455
rect 3192 443 3194 454
rect 3191 442 3195 443
rect 3191 437 3195 438
rect 3192 430 3194 437
rect 3190 429 3196 430
rect 3190 425 3191 429
rect 3195 425 3196 429
rect 3190 424 3196 425
rect 2862 411 2868 412
rect 2246 407 2252 408
rect 2246 403 2247 407
rect 2251 403 2252 407
rect 2246 402 2252 403
rect 2258 407 2264 408
rect 2258 403 2259 407
rect 2263 403 2264 407
rect 2258 402 2264 403
rect 2374 407 2380 408
rect 2374 403 2375 407
rect 2379 403 2380 407
rect 2374 402 2380 403
rect 2386 407 2392 408
rect 2386 403 2387 407
rect 2391 403 2392 407
rect 2386 402 2392 403
rect 2502 407 2508 408
rect 2502 403 2503 407
rect 2507 403 2508 407
rect 2502 402 2508 403
rect 2514 407 2520 408
rect 2514 403 2515 407
rect 2519 403 2520 407
rect 2514 402 2520 403
rect 2622 407 2628 408
rect 2622 403 2623 407
rect 2627 403 2628 407
rect 2622 402 2628 403
rect 2630 407 2636 408
rect 2630 403 2631 407
rect 2635 403 2636 407
rect 2630 402 2636 403
rect 2670 407 2676 408
rect 2670 403 2671 407
rect 2675 403 2676 407
rect 2670 402 2676 403
rect 2742 407 2748 408
rect 2742 403 2743 407
rect 2747 403 2748 407
rect 2742 402 2748 403
rect 2750 407 2756 408
rect 2750 403 2751 407
rect 2755 403 2756 407
rect 2750 402 2756 403
rect 2798 407 2804 408
rect 2798 403 2799 407
rect 2803 403 2804 407
rect 2798 402 2804 403
rect 2854 407 2860 408
rect 2854 403 2855 407
rect 2859 403 2860 407
rect 2862 407 2863 411
rect 2867 407 2868 411
rect 2862 406 2868 407
rect 2926 411 2932 412
rect 2926 407 2927 411
rect 2931 407 2932 411
rect 3118 411 3124 412
rect 2926 406 2932 407
rect 2966 407 2972 408
rect 2854 402 2860 403
rect 2248 391 2250 402
rect 2151 390 2155 391
rect 2247 390 2251 391
rect 2150 385 2156 386
rect 2247 385 2251 386
rect 2150 381 2151 385
rect 2155 381 2156 385
rect 2150 380 2156 381
rect 2260 380 2262 402
rect 2376 391 2378 402
rect 2279 390 2283 391
rect 2375 390 2379 391
rect 2278 385 2284 386
rect 2375 385 2379 386
rect 2278 381 2279 385
rect 2283 381 2284 385
rect 2278 380 2284 381
rect 2388 380 2390 402
rect 2504 391 2506 402
rect 2407 390 2411 391
rect 2503 390 2507 391
rect 2406 385 2412 386
rect 2503 385 2507 386
rect 2406 381 2407 385
rect 2411 381 2412 385
rect 2406 380 2412 381
rect 2516 380 2518 402
rect 2624 391 2626 402
rect 2535 390 2539 391
rect 2623 390 2627 391
rect 2663 390 2667 391
rect 2534 385 2540 386
rect 2623 385 2627 386
rect 2662 385 2668 386
rect 2534 381 2535 385
rect 2539 381 2540 385
rect 2534 380 2540 381
rect 2662 381 2663 385
rect 2667 381 2668 385
rect 2672 384 2674 402
rect 2744 391 2746 402
rect 2743 390 2747 391
rect 2743 385 2747 386
rect 2752 384 2754 402
rect 2791 390 2795 391
rect 2790 385 2796 386
rect 2662 380 2668 381
rect 2670 383 2676 384
rect 2258 379 2264 380
rect 2258 375 2259 379
rect 2263 375 2264 379
rect 2258 374 2264 375
rect 2386 379 2392 380
rect 2386 375 2387 379
rect 2391 375 2392 379
rect 2386 374 2392 375
rect 2514 379 2520 380
rect 2514 375 2515 379
rect 2519 375 2520 379
rect 2514 374 2520 375
rect 2574 379 2580 380
rect 2574 375 2575 379
rect 2579 375 2580 379
rect 2670 379 2671 383
rect 2675 379 2676 383
rect 2670 378 2676 379
rect 2750 383 2756 384
rect 2750 379 2751 383
rect 2755 379 2756 383
rect 2790 381 2791 385
rect 2795 381 2796 385
rect 2800 384 2802 402
rect 2856 391 2858 402
rect 2855 390 2859 391
rect 2855 385 2859 386
rect 2864 384 2866 406
rect 2919 390 2923 391
rect 2918 385 2924 386
rect 2790 380 2796 381
rect 2798 383 2804 384
rect 2750 378 2756 379
rect 2798 379 2799 383
rect 2803 379 2804 383
rect 2798 378 2804 379
rect 2862 383 2868 384
rect 2862 379 2863 383
rect 2867 379 2868 383
rect 2918 381 2919 385
rect 2923 381 2924 385
rect 2928 384 2930 406
rect 2966 403 2967 407
rect 2971 403 2972 407
rect 2966 402 2972 403
rect 2974 407 2980 408
rect 2974 403 2975 407
rect 2979 403 2980 407
rect 2974 402 2980 403
rect 3034 407 3040 408
rect 3034 403 3035 407
rect 3039 403 3040 407
rect 3034 402 3040 403
rect 3086 407 3092 408
rect 3086 403 3087 407
rect 3091 403 3092 407
rect 3118 407 3119 411
rect 3123 407 3124 411
rect 3118 406 3124 407
rect 3190 411 3196 412
rect 3190 407 3191 411
rect 3195 407 3196 411
rect 3190 406 3196 407
rect 3086 402 3092 403
rect 2968 391 2970 402
rect 2967 390 2971 391
rect 2967 385 2971 386
rect 2976 384 2978 402
rect 2918 380 2924 381
rect 2926 383 2932 384
rect 2862 378 2868 379
rect 2926 379 2927 383
rect 2931 379 2932 383
rect 2926 378 2932 379
rect 2974 383 2980 384
rect 2974 379 2975 383
rect 2979 379 2980 383
rect 3036 380 3038 402
rect 3088 391 3090 402
rect 3047 390 3051 391
rect 3087 390 3091 391
rect 3046 385 3052 386
rect 3087 385 3091 386
rect 3046 381 3047 385
rect 3051 381 3052 385
rect 3046 380 3052 381
rect 3120 380 3122 406
rect 3192 391 3194 406
rect 3159 390 3163 391
rect 3191 390 3195 391
rect 3158 385 3164 386
rect 3191 385 3195 386
rect 3158 381 3159 385
rect 3163 381 3164 385
rect 3192 382 3194 385
rect 3158 380 3164 381
rect 3190 381 3196 382
rect 2974 378 2980 379
rect 3034 379 3040 380
rect 2574 374 2580 375
rect 2150 356 2156 357
rect 2150 352 2151 356
rect 2155 352 2156 356
rect 2150 351 2156 352
rect 2278 356 2284 357
rect 2278 352 2279 356
rect 2283 352 2284 356
rect 2278 351 2284 352
rect 2406 356 2412 357
rect 2406 352 2407 356
rect 2411 352 2412 356
rect 2406 351 2412 352
rect 2534 356 2540 357
rect 2534 352 2535 356
rect 2539 352 2540 356
rect 2534 351 2540 352
rect 2152 339 2154 351
rect 2280 339 2282 351
rect 2408 339 2410 351
rect 2536 339 2538 351
rect 2151 338 2155 339
rect 2151 333 2155 334
rect 2175 338 2179 339
rect 2175 333 2179 334
rect 2279 338 2283 339
rect 2279 333 2283 334
rect 2303 338 2307 339
rect 2303 333 2307 334
rect 2407 338 2411 339
rect 2407 333 2411 334
rect 2431 338 2435 339
rect 2431 333 2435 334
rect 2535 338 2539 339
rect 2535 333 2539 334
rect 2567 338 2571 339
rect 2567 333 2571 334
rect 2174 332 2180 333
rect 2174 328 2175 332
rect 2179 328 2180 332
rect 2174 327 2180 328
rect 2302 332 2308 333
rect 2302 328 2303 332
rect 2307 328 2308 332
rect 2302 327 2308 328
rect 2430 332 2436 333
rect 2430 328 2431 332
rect 2435 328 2436 332
rect 2430 327 2436 328
rect 2566 332 2572 333
rect 2566 328 2567 332
rect 2571 328 2572 332
rect 2566 327 2572 328
rect 2439 307 2445 308
rect 1367 302 1371 303
rect 1367 297 1371 298
rect 1631 302 1635 303
rect 1670 302 1676 303
rect 2046 303 2052 304
rect 1631 297 1635 298
rect 1632 290 1634 297
rect 1672 291 1674 302
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 2046 298 2052 299
rect 2058 303 2064 304
rect 2058 299 2059 303
rect 2063 299 2064 303
rect 2058 298 2064 299
rect 2174 303 2180 304
rect 2174 299 2175 303
rect 2179 299 2180 303
rect 2174 298 2180 299
rect 2186 303 2192 304
rect 2186 299 2187 303
rect 2191 299 2192 303
rect 2186 298 2192 299
rect 2302 303 2308 304
rect 2302 299 2303 303
rect 2307 299 2308 303
rect 2302 298 2308 299
rect 2326 303 2332 304
rect 2326 299 2327 303
rect 2331 299 2332 303
rect 2326 298 2332 299
rect 2430 303 2436 304
rect 2430 299 2431 303
rect 2435 299 2436 303
rect 2439 303 2440 307
rect 2444 306 2445 307
rect 2444 304 2450 306
rect 2576 304 2578 374
rect 2662 356 2668 357
rect 2662 352 2663 356
rect 2667 352 2668 356
rect 2662 351 2668 352
rect 2790 356 2796 357
rect 2790 352 2791 356
rect 2795 352 2796 356
rect 2790 351 2796 352
rect 2918 356 2924 357
rect 2918 352 2919 356
rect 2923 352 2924 356
rect 2918 351 2924 352
rect 2664 339 2666 351
rect 2792 339 2794 351
rect 2920 339 2922 351
rect 2663 338 2667 339
rect 2663 333 2667 334
rect 2711 338 2715 339
rect 2711 333 2715 334
rect 2791 338 2795 339
rect 2791 333 2795 334
rect 2863 338 2867 339
rect 2863 333 2867 334
rect 2919 338 2923 339
rect 2919 333 2923 334
rect 2710 332 2716 333
rect 2710 328 2711 332
rect 2715 328 2716 332
rect 2710 327 2716 328
rect 2862 332 2868 333
rect 2862 328 2863 332
rect 2867 328 2868 332
rect 2862 327 2868 328
rect 2928 308 2930 378
rect 3034 375 3035 379
rect 3039 375 3040 379
rect 3034 374 3040 375
rect 3118 379 3124 380
rect 3118 375 3119 379
rect 3123 375 3124 379
rect 3118 374 3124 375
rect 3166 379 3172 380
rect 3166 375 3167 379
rect 3171 375 3172 379
rect 3190 377 3191 381
rect 3195 377 3196 381
rect 3190 376 3196 377
rect 3166 374 3172 375
rect 3023 338 3027 339
rect 3023 333 3027 334
rect 3022 332 3028 333
rect 3022 328 3023 332
rect 3027 328 3028 332
rect 3022 327 3028 328
rect 3036 308 3038 374
rect 3046 356 3052 357
rect 3046 352 3047 356
rect 3051 352 3052 356
rect 3046 351 3052 352
rect 3158 356 3164 357
rect 3158 352 3159 356
rect 3163 352 3164 356
rect 3158 351 3164 352
rect 3048 339 3050 351
rect 3160 339 3162 351
rect 3047 338 3051 339
rect 3047 333 3051 334
rect 3159 338 3163 339
rect 3159 333 3163 334
rect 3158 332 3164 333
rect 3158 328 3159 332
rect 3163 328 3164 332
rect 3158 327 3164 328
rect 3168 308 3170 374
rect 3190 363 3196 364
rect 3190 359 3191 363
rect 3195 359 3196 363
rect 3190 358 3196 359
rect 3192 339 3194 358
rect 3191 338 3195 339
rect 3191 333 3195 334
rect 3192 326 3194 333
rect 3190 325 3196 326
rect 3190 321 3191 325
rect 3195 321 3196 325
rect 3190 320 3196 321
rect 2870 307 2876 308
rect 2444 303 2445 304
rect 2439 302 2445 303
rect 2430 298 2436 299
rect 2048 291 2050 298
rect 1671 290 1675 291
rect 1630 289 1636 290
rect 1630 285 1631 289
rect 1635 285 1636 289
rect 1943 290 1947 291
rect 2047 290 2051 291
rect 1671 285 1675 286
rect 1942 285 1948 286
rect 2047 285 2051 286
rect 1630 284 1636 285
rect 1672 282 1674 285
rect 1670 281 1676 282
rect 1670 277 1671 281
rect 1675 277 1676 281
rect 1942 281 1943 285
rect 1947 281 1948 285
rect 1942 280 1948 281
rect 2060 280 2062 298
rect 2176 291 2178 298
rect 2071 290 2075 291
rect 2175 290 2179 291
rect 2070 285 2076 286
rect 2175 285 2179 286
rect 2070 281 2071 285
rect 2075 281 2076 285
rect 2070 280 2076 281
rect 2188 280 2190 298
rect 2304 291 2306 298
rect 2199 290 2203 291
rect 2303 290 2307 291
rect 2319 290 2323 291
rect 2198 285 2204 286
rect 2303 285 2307 286
rect 2318 285 2324 286
rect 2198 281 2199 285
rect 2203 281 2204 285
rect 2198 280 2204 281
rect 2318 281 2319 285
rect 2323 281 2324 285
rect 2318 280 2324 281
rect 2328 280 2330 298
rect 2432 291 2434 298
rect 2431 290 2435 291
rect 2439 290 2443 291
rect 2431 285 2435 286
rect 2438 285 2444 286
rect 2438 281 2439 285
rect 2443 281 2444 285
rect 2438 280 2444 281
rect 2448 280 2450 304
rect 2566 303 2572 304
rect 2566 299 2567 303
rect 2571 299 2572 303
rect 2566 298 2572 299
rect 2574 303 2580 304
rect 2574 299 2575 303
rect 2579 299 2580 303
rect 2574 298 2580 299
rect 2670 303 2676 304
rect 2670 299 2671 303
rect 2675 299 2676 303
rect 2670 298 2676 299
rect 2710 303 2716 304
rect 2710 299 2711 303
rect 2715 299 2716 303
rect 2710 298 2716 299
rect 2718 303 2724 304
rect 2718 299 2719 303
rect 2723 299 2724 303
rect 2718 298 2724 299
rect 2790 303 2796 304
rect 2790 299 2791 303
rect 2795 299 2796 303
rect 2790 298 2796 299
rect 2862 303 2868 304
rect 2862 299 2863 303
rect 2867 299 2868 303
rect 2870 303 2871 307
rect 2875 303 2876 307
rect 2870 302 2876 303
rect 2926 307 2932 308
rect 2926 303 2927 307
rect 2931 303 2932 307
rect 3034 307 3040 308
rect 2926 302 2932 303
rect 3022 303 3028 304
rect 2862 298 2868 299
rect 2568 291 2570 298
rect 2551 290 2555 291
rect 2567 290 2571 291
rect 2550 285 2556 286
rect 2567 285 2571 286
rect 2550 281 2551 285
rect 2555 281 2556 285
rect 2576 284 2578 298
rect 2663 290 2667 291
rect 2662 285 2668 286
rect 2550 280 2556 281
rect 2574 283 2580 284
rect 1670 276 1676 277
rect 2058 279 2064 280
rect 2058 275 2059 279
rect 2063 275 2064 279
rect 2058 274 2064 275
rect 2186 279 2192 280
rect 2186 275 2187 279
rect 2191 275 2192 279
rect 2186 274 2192 275
rect 2326 279 2332 280
rect 2326 275 2327 279
rect 2331 275 2332 279
rect 2326 274 2332 275
rect 2446 279 2452 280
rect 2446 275 2447 279
rect 2451 275 2452 279
rect 2446 274 2452 275
rect 2526 279 2532 280
rect 2526 275 2527 279
rect 2531 275 2532 279
rect 2574 279 2575 283
rect 2579 279 2580 283
rect 2662 281 2663 285
rect 2667 281 2668 285
rect 2672 284 2674 298
rect 2712 291 2714 298
rect 2711 290 2715 291
rect 2711 285 2715 286
rect 2720 284 2722 298
rect 2783 290 2787 291
rect 2782 285 2788 286
rect 2662 280 2668 281
rect 2670 283 2676 284
rect 2574 278 2580 279
rect 2670 279 2671 283
rect 2675 279 2676 283
rect 2670 278 2676 279
rect 2718 283 2724 284
rect 2718 279 2719 283
rect 2723 279 2724 283
rect 2782 281 2783 285
rect 2787 281 2788 285
rect 2792 284 2794 298
rect 2864 291 2866 298
rect 2863 290 2867 291
rect 2863 285 2867 286
rect 2872 284 2874 302
rect 2782 280 2788 281
rect 2790 283 2796 284
rect 2718 278 2724 279
rect 2790 279 2791 283
rect 2795 279 2796 283
rect 2790 278 2796 279
rect 2870 283 2876 284
rect 2870 279 2871 283
rect 2875 279 2876 283
rect 2870 278 2876 279
rect 2526 274 2532 275
rect 774 271 780 272
rect 470 266 476 267
rect 622 267 628 268
rect 462 262 468 263
rect 464 259 466 262
rect 111 258 115 259
rect 359 258 363 259
rect 463 258 467 259
rect 111 253 115 254
rect 358 253 364 254
rect 463 253 467 254
rect 112 250 114 253
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 358 249 359 253
rect 363 249 364 253
rect 472 252 474 266
rect 622 263 623 267
rect 627 263 628 267
rect 622 262 628 263
rect 630 267 636 268
rect 630 263 631 267
rect 635 263 636 267
rect 630 262 636 263
rect 766 267 772 268
rect 766 263 767 267
rect 771 263 772 267
rect 774 267 775 271
rect 779 267 780 271
rect 774 266 780 267
rect 814 271 820 272
rect 814 267 815 271
rect 819 267 820 271
rect 1294 271 1300 272
rect 814 266 820 267
rect 902 267 908 268
rect 766 262 772 263
rect 624 259 626 262
rect 487 258 491 259
rect 623 258 627 259
rect 486 253 492 254
rect 358 248 364 249
rect 366 251 372 252
rect 366 247 367 251
rect 371 247 372 251
rect 366 246 372 247
rect 470 251 476 252
rect 470 247 471 251
rect 475 247 476 251
rect 486 249 487 253
rect 491 249 492 253
rect 486 248 492 249
rect 622 253 628 254
rect 622 249 623 253
rect 627 249 628 253
rect 622 248 628 249
rect 632 248 634 262
rect 768 259 770 262
rect 759 258 763 259
rect 767 258 771 259
rect 758 253 764 254
rect 767 253 771 254
rect 758 249 759 253
rect 763 249 764 253
rect 758 248 764 249
rect 470 246 476 247
rect 630 247 636 248
rect 110 244 116 245
rect 110 231 116 232
rect 110 227 111 231
rect 115 227 116 231
rect 110 226 116 227
rect 112 215 114 226
rect 358 224 364 225
rect 358 220 359 224
rect 363 220 364 224
rect 358 219 364 220
rect 360 215 362 219
rect 111 214 115 215
rect 111 209 115 210
rect 279 214 283 215
rect 279 209 283 210
rect 359 214 363 215
rect 359 209 363 210
rect 112 202 114 209
rect 278 208 284 209
rect 278 204 279 208
rect 283 204 284 208
rect 278 203 284 204
rect 110 201 116 202
rect 110 197 111 201
rect 115 197 116 201
rect 110 196 116 197
rect 368 184 370 246
rect 447 214 451 215
rect 447 209 451 210
rect 446 208 452 209
rect 446 204 447 208
rect 451 204 452 208
rect 446 203 452 204
rect 472 184 474 246
rect 630 243 631 247
rect 635 243 636 247
rect 630 242 636 243
rect 766 243 772 244
rect 776 243 778 266
rect 902 263 903 267
rect 907 263 908 267
rect 902 262 908 263
rect 1030 267 1036 268
rect 1030 263 1031 267
rect 1035 263 1036 267
rect 1030 262 1036 263
rect 1158 267 1164 268
rect 1158 263 1159 267
rect 1163 263 1164 267
rect 1158 262 1164 263
rect 1286 267 1292 268
rect 1286 263 1287 267
rect 1291 263 1292 267
rect 1294 267 1295 271
rect 1299 267 1300 271
rect 1294 266 1300 267
rect 1630 271 1636 272
rect 1630 267 1631 271
rect 1635 267 1636 271
rect 1630 266 1636 267
rect 1286 262 1292 263
rect 904 259 906 262
rect 1032 259 1034 262
rect 1160 259 1162 262
rect 1288 259 1290 262
rect 895 258 899 259
rect 903 258 907 259
rect 894 253 900 254
rect 903 253 907 254
rect 1031 258 1035 259
rect 1039 258 1043 259
rect 1159 258 1163 259
rect 1183 258 1187 259
rect 1287 258 1291 259
rect 1031 253 1035 254
rect 1038 253 1044 254
rect 1159 253 1163 254
rect 1182 253 1188 254
rect 1287 253 1291 254
rect 894 249 895 253
rect 899 249 900 253
rect 894 248 900 249
rect 1038 249 1039 253
rect 1043 249 1044 253
rect 1038 248 1044 249
rect 1182 249 1183 253
rect 1187 249 1188 253
rect 1296 252 1298 266
rect 1632 259 1634 266
rect 1670 263 1676 264
rect 1670 259 1671 263
rect 1675 259 1676 263
rect 1631 258 1635 259
rect 1670 258 1676 259
rect 1631 253 1635 254
rect 1182 248 1188 249
rect 1294 251 1300 252
rect 486 224 492 225
rect 486 220 487 224
rect 491 220 492 224
rect 486 219 492 220
rect 622 224 628 225
rect 622 220 623 224
rect 627 220 628 224
rect 622 219 628 220
rect 488 215 490 219
rect 624 215 626 219
rect 487 214 491 215
rect 487 209 491 210
rect 615 214 619 215
rect 615 209 619 210
rect 623 214 627 215
rect 623 209 627 210
rect 614 208 620 209
rect 614 204 615 208
rect 619 204 620 208
rect 614 203 620 204
rect 110 183 116 184
rect 110 179 111 183
rect 115 179 116 183
rect 366 183 372 184
rect 110 178 116 179
rect 278 179 284 180
rect 112 175 114 178
rect 278 175 279 179
rect 283 175 284 179
rect 366 179 367 183
rect 371 179 372 183
rect 470 183 476 184
rect 366 178 372 179
rect 446 179 452 180
rect 446 175 447 179
rect 451 175 452 179
rect 470 179 471 183
rect 475 179 476 183
rect 470 178 476 179
rect 614 179 620 180
rect 111 174 115 175
rect 199 174 203 175
rect 278 174 284 175
rect 367 174 371 175
rect 446 174 452 175
rect 111 169 115 170
rect 198 169 204 170
rect 279 169 283 170
rect 366 169 372 170
rect 447 169 451 170
rect 112 166 114 169
rect 110 165 116 166
rect 110 161 111 165
rect 115 161 116 165
rect 198 165 199 169
rect 203 165 204 169
rect 198 164 204 165
rect 366 165 367 169
rect 371 165 372 169
rect 366 164 372 165
rect 472 164 474 178
rect 614 175 615 179
rect 619 175 620 179
rect 535 174 539 175
rect 614 174 620 175
rect 623 179 629 180
rect 623 175 624 179
rect 628 178 629 179
rect 632 178 634 242
rect 766 239 767 243
rect 771 241 778 243
rect 902 247 908 248
rect 902 243 903 247
rect 907 243 908 247
rect 1294 247 1295 251
rect 1299 247 1300 251
rect 1632 250 1634 253
rect 1294 246 1300 247
rect 1630 249 1636 250
rect 1630 245 1631 249
rect 1635 245 1636 249
rect 1630 244 1636 245
rect 902 242 908 243
rect 771 239 772 241
rect 766 238 772 239
rect 758 224 764 225
rect 758 220 759 224
rect 763 220 764 224
rect 758 219 764 220
rect 760 215 762 219
rect 759 214 763 215
rect 759 209 763 210
rect 628 176 634 178
rect 628 175 629 176
rect 623 174 629 175
rect 695 174 699 175
rect 534 169 540 170
rect 615 169 619 170
rect 694 169 700 170
rect 534 165 535 169
rect 539 165 540 169
rect 534 164 540 165
rect 694 165 695 169
rect 699 165 700 169
rect 694 164 700 165
rect 768 164 770 238
rect 894 224 900 225
rect 894 220 895 224
rect 899 220 900 224
rect 894 219 900 220
rect 896 215 898 219
rect 775 214 779 215
rect 775 209 779 210
rect 895 214 899 215
rect 895 209 899 210
rect 774 208 780 209
rect 774 204 775 208
rect 779 204 780 208
rect 774 203 780 204
rect 904 188 906 242
rect 1672 239 1674 258
rect 1942 256 1948 257
rect 1942 252 1943 256
rect 1947 252 1948 256
rect 1942 251 1948 252
rect 2070 256 2076 257
rect 2070 252 2071 256
rect 2075 252 2076 256
rect 2070 251 2076 252
rect 2198 256 2204 257
rect 2198 252 2199 256
rect 2203 252 2204 256
rect 2198 251 2204 252
rect 2318 256 2324 257
rect 2318 252 2319 256
rect 2323 252 2324 256
rect 2318 251 2324 252
rect 2438 256 2444 257
rect 2438 252 2439 256
rect 2443 252 2444 256
rect 2438 251 2444 252
rect 1944 239 1946 251
rect 2072 239 2074 251
rect 2200 239 2202 251
rect 2320 239 2322 251
rect 2440 239 2442 251
rect 1671 238 1675 239
rect 1671 233 1675 234
rect 1847 238 1851 239
rect 1847 233 1851 234
rect 1943 238 1947 239
rect 1943 233 1947 234
rect 1975 238 1979 239
rect 1975 233 1979 234
rect 2071 238 2075 239
rect 2071 233 2075 234
rect 2103 238 2107 239
rect 2103 233 2107 234
rect 2199 238 2203 239
rect 2199 233 2203 234
rect 2247 238 2251 239
rect 2247 233 2251 234
rect 2319 238 2323 239
rect 2319 233 2323 234
rect 2407 238 2411 239
rect 2407 233 2411 234
rect 2439 238 2443 239
rect 2439 233 2443 234
rect 1630 231 1636 232
rect 1630 227 1631 231
rect 1635 227 1636 231
rect 1630 226 1636 227
rect 1672 226 1674 233
rect 1846 232 1852 233
rect 1846 228 1847 232
rect 1851 228 1852 232
rect 1846 227 1852 228
rect 1974 232 1980 233
rect 1974 228 1975 232
rect 1979 228 1980 232
rect 1974 227 1980 228
rect 2102 232 2108 233
rect 2102 228 2103 232
rect 2107 228 2108 232
rect 2102 227 2108 228
rect 2246 232 2252 233
rect 2246 228 2247 232
rect 2251 228 2252 232
rect 2246 227 2252 228
rect 2406 232 2412 233
rect 2406 228 2407 232
rect 2411 228 2412 232
rect 2406 227 2412 228
rect 1038 224 1044 225
rect 1038 220 1039 224
rect 1043 220 1044 224
rect 1038 219 1044 220
rect 1182 224 1188 225
rect 1182 220 1183 224
rect 1187 220 1188 224
rect 1182 219 1188 220
rect 1040 215 1042 219
rect 1184 215 1186 219
rect 1632 215 1634 226
rect 1670 225 1676 226
rect 1670 221 1671 225
rect 1675 221 1676 225
rect 1670 220 1676 221
rect 943 214 947 215
rect 943 209 947 210
rect 1039 214 1043 215
rect 1039 209 1043 210
rect 1111 214 1115 215
rect 1111 209 1115 210
rect 1183 214 1187 215
rect 1183 209 1187 210
rect 1631 214 1635 215
rect 1631 209 1635 210
rect 942 208 948 209
rect 942 204 943 208
rect 947 204 948 208
rect 942 203 948 204
rect 1110 208 1116 209
rect 1110 204 1111 208
rect 1115 204 1116 208
rect 1110 203 1116 204
rect 1632 202 1634 209
rect 1670 207 1676 208
rect 1670 203 1671 207
rect 1675 203 1676 207
rect 1670 202 1676 203
rect 1846 203 1852 204
rect 1630 201 1636 202
rect 1630 197 1631 201
rect 1635 197 1636 201
rect 1630 196 1636 197
rect 902 187 908 188
rect 1672 187 1674 202
rect 1846 199 1847 203
rect 1851 199 1852 203
rect 1846 198 1852 199
rect 1854 203 1860 204
rect 1854 199 1855 203
rect 1859 199 1860 203
rect 1854 198 1860 199
rect 1974 203 1980 204
rect 1974 199 1975 203
rect 1979 199 1980 203
rect 1974 198 1980 199
rect 1982 203 1988 204
rect 1982 199 1983 203
rect 1987 199 1988 203
rect 1982 198 1988 199
rect 2102 203 2108 204
rect 2102 199 2103 203
rect 2107 199 2108 203
rect 2102 198 2108 199
rect 2110 203 2116 204
rect 2110 199 2111 203
rect 2115 199 2116 203
rect 2110 198 2116 199
rect 2246 203 2252 204
rect 2246 199 2247 203
rect 2251 199 2252 203
rect 2246 198 2252 199
rect 2254 203 2260 204
rect 2254 199 2255 203
rect 2259 199 2260 203
rect 2254 198 2260 199
rect 2318 203 2324 204
rect 2318 199 2319 203
rect 2323 199 2324 203
rect 2318 198 2324 199
rect 2406 203 2412 204
rect 2406 199 2407 203
rect 2411 199 2412 203
rect 2406 198 2412 199
rect 2414 203 2420 204
rect 2414 199 2415 203
rect 2419 199 2420 203
rect 2414 198 2420 199
rect 2502 203 2508 204
rect 2502 199 2503 203
rect 2507 199 2508 203
rect 2502 198 2508 199
rect 1848 187 1850 198
rect 902 183 903 187
rect 907 183 908 187
rect 1671 186 1675 187
rect 902 182 908 183
rect 1630 183 1636 184
rect 774 179 780 180
rect 774 175 775 179
rect 779 175 780 179
rect 774 174 780 175
rect 863 174 867 175
rect 775 169 779 170
rect 862 169 868 170
rect 862 165 863 169
rect 867 165 868 169
rect 862 164 868 165
rect 904 164 906 182
rect 942 179 948 180
rect 942 175 943 179
rect 947 175 948 179
rect 1110 179 1116 180
rect 1110 175 1111 179
rect 1115 175 1116 179
rect 1630 179 1631 183
rect 1635 179 1636 183
rect 1743 186 1747 187
rect 1847 186 1851 187
rect 1671 181 1675 182
rect 1742 181 1748 182
rect 1847 181 1851 182
rect 1630 178 1636 179
rect 1672 178 1674 181
rect 1632 175 1634 178
rect 1670 177 1676 178
rect 942 174 948 175
rect 1031 174 1035 175
rect 1110 174 1116 175
rect 1631 174 1635 175
rect 943 169 947 170
rect 1030 169 1036 170
rect 1111 169 1115 170
rect 1670 173 1671 177
rect 1675 173 1676 177
rect 1742 177 1743 181
rect 1747 177 1748 181
rect 1742 176 1748 177
rect 1856 176 1858 198
rect 1976 187 1978 198
rect 1871 186 1875 187
rect 1975 186 1979 187
rect 1870 181 1876 182
rect 1975 181 1979 182
rect 1870 177 1871 181
rect 1875 177 1876 181
rect 1870 176 1876 177
rect 1984 176 1986 198
rect 2104 187 2106 198
rect 1999 186 2003 187
rect 2103 186 2107 187
rect 1998 181 2004 182
rect 2103 181 2107 182
rect 1998 177 1999 181
rect 2003 177 2004 181
rect 1998 176 2004 177
rect 2112 176 2114 198
rect 2248 187 2250 198
rect 2143 186 2147 187
rect 2247 186 2251 187
rect 2142 181 2148 182
rect 2247 181 2251 182
rect 2142 177 2143 181
rect 2147 177 2148 181
rect 2256 180 2258 198
rect 2311 186 2315 187
rect 2310 181 2316 182
rect 2142 176 2148 177
rect 2254 179 2260 180
rect 1670 172 1676 173
rect 1750 175 1756 176
rect 1750 171 1751 175
rect 1755 171 1756 175
rect 1750 170 1756 171
rect 1854 175 1860 176
rect 1854 171 1855 175
rect 1859 171 1860 175
rect 1854 170 1860 171
rect 1982 175 1988 176
rect 1982 171 1983 175
rect 1987 171 1988 175
rect 1982 170 1988 171
rect 2110 175 2116 176
rect 2110 171 2111 175
rect 2115 171 2116 175
rect 2254 175 2255 179
rect 2259 175 2260 179
rect 2310 177 2311 181
rect 2315 177 2316 181
rect 2320 180 2322 198
rect 2408 187 2410 198
rect 2407 186 2411 187
rect 2407 181 2411 182
rect 2416 180 2418 198
rect 2495 186 2499 187
rect 2494 181 2500 182
rect 2310 176 2316 177
rect 2318 179 2324 180
rect 2254 174 2260 175
rect 2318 175 2319 179
rect 2323 175 2324 179
rect 2318 174 2324 175
rect 2358 179 2364 180
rect 2358 175 2359 179
rect 2363 175 2364 179
rect 2358 174 2364 175
rect 2414 179 2420 180
rect 2414 175 2415 179
rect 2419 175 2420 179
rect 2494 177 2495 181
rect 2499 177 2500 181
rect 2504 180 2506 198
rect 2494 176 2500 177
rect 2502 179 2508 180
rect 2414 174 2420 175
rect 2502 175 2503 179
rect 2507 175 2508 179
rect 2502 174 2508 175
rect 2110 170 2116 171
rect 1631 169 1635 170
rect 1030 165 1031 169
rect 1035 165 1036 169
rect 1632 166 1634 169
rect 1030 164 1036 165
rect 1630 165 1636 166
rect 110 160 116 161
rect 146 163 152 164
rect 146 159 147 163
rect 151 159 152 163
rect 146 158 152 159
rect 470 163 476 164
rect 470 159 471 163
rect 475 159 476 163
rect 470 158 476 159
rect 546 163 552 164
rect 546 159 547 163
rect 551 159 552 163
rect 546 158 552 159
rect 702 163 708 164
rect 702 159 703 163
rect 707 159 708 163
rect 702 158 708 159
rect 766 163 772 164
rect 766 159 767 163
rect 771 159 772 163
rect 766 158 772 159
rect 902 163 908 164
rect 902 159 903 163
rect 907 159 908 163
rect 902 158 908 159
rect 1022 163 1028 164
rect 1022 159 1023 163
rect 1027 159 1028 163
rect 1630 161 1631 165
rect 1635 161 1636 165
rect 1630 160 1636 161
rect 1022 158 1028 159
rect 1670 159 1676 160
rect 110 147 116 148
rect 110 143 111 147
rect 115 143 116 147
rect 110 142 116 143
rect 112 123 114 142
rect 111 122 115 123
rect 111 117 115 118
rect 135 122 139 123
rect 135 117 139 118
rect 112 110 114 117
rect 134 116 140 117
rect 134 112 135 116
rect 139 112 140 116
rect 134 111 140 112
rect 110 109 116 110
rect 110 105 111 109
rect 115 105 116 109
rect 110 104 116 105
rect 148 92 150 158
rect 198 140 204 141
rect 198 136 199 140
rect 203 136 204 140
rect 198 135 204 136
rect 366 140 372 141
rect 366 136 367 140
rect 371 136 372 140
rect 366 135 372 136
rect 534 140 540 141
rect 534 136 535 140
rect 539 136 540 140
rect 534 135 540 136
rect 200 123 202 135
rect 368 123 370 135
rect 536 123 538 135
rect 191 122 195 123
rect 191 117 195 118
rect 199 122 203 123
rect 199 117 203 118
rect 287 122 291 123
rect 287 117 291 118
rect 367 122 371 123
rect 367 117 371 118
rect 383 122 387 123
rect 383 117 387 118
rect 479 122 483 123
rect 479 117 483 118
rect 535 122 539 123
rect 535 117 539 118
rect 190 116 196 117
rect 190 112 191 116
rect 195 112 196 116
rect 190 111 196 112
rect 286 116 292 117
rect 286 112 287 116
rect 291 112 292 116
rect 286 111 292 112
rect 382 116 388 117
rect 382 112 383 116
rect 387 112 388 116
rect 382 111 388 112
rect 478 116 484 117
rect 478 112 479 116
rect 483 112 484 116
rect 478 111 484 112
rect 548 96 550 158
rect 694 140 700 141
rect 694 136 695 140
rect 699 136 700 140
rect 694 135 700 136
rect 696 123 698 135
rect 583 122 587 123
rect 583 117 587 118
rect 695 122 699 123
rect 695 117 699 118
rect 582 116 588 117
rect 582 112 583 116
rect 587 112 588 116
rect 582 111 588 112
rect 694 116 700 117
rect 694 112 695 116
rect 699 112 700 116
rect 694 111 700 112
rect 546 95 552 96
rect 110 91 116 92
rect 110 87 111 91
rect 115 87 116 91
rect 146 91 152 92
rect 110 86 116 87
rect 134 87 140 88
rect 112 83 114 86
rect 134 83 135 87
rect 139 83 140 87
rect 146 87 147 91
rect 151 87 152 91
rect 546 91 547 95
rect 551 91 552 95
rect 704 92 706 158
rect 862 140 868 141
rect 862 136 863 140
rect 867 136 868 140
rect 862 135 868 136
rect 864 123 866 135
rect 815 122 819 123
rect 815 117 819 118
rect 863 122 867 123
rect 863 117 867 118
rect 943 122 947 123
rect 943 117 947 118
rect 814 116 820 117
rect 814 112 815 116
rect 819 112 820 116
rect 814 111 820 112
rect 942 116 948 117
rect 942 112 943 116
rect 947 112 948 116
rect 942 111 948 112
rect 1024 96 1026 158
rect 1670 155 1671 159
rect 1675 155 1676 159
rect 1670 154 1676 155
rect 1630 147 1636 148
rect 1630 143 1631 147
rect 1635 143 1636 147
rect 1630 142 1636 143
rect 1030 140 1036 141
rect 1030 136 1031 140
rect 1035 136 1036 140
rect 1030 135 1036 136
rect 1032 123 1034 135
rect 1632 123 1634 142
rect 1672 131 1674 154
rect 1742 152 1748 153
rect 1742 148 1743 152
rect 1747 148 1748 152
rect 1742 147 1748 148
rect 1744 131 1746 147
rect 1671 130 1675 131
rect 1671 125 1675 126
rect 1695 130 1699 131
rect 1695 125 1699 126
rect 1743 130 1747 131
rect 1743 125 1747 126
rect 1031 122 1035 123
rect 1031 117 1035 118
rect 1079 122 1083 123
rect 1079 117 1083 118
rect 1215 122 1219 123
rect 1215 117 1219 118
rect 1351 122 1355 123
rect 1351 117 1355 118
rect 1487 122 1491 123
rect 1487 117 1491 118
rect 1599 122 1603 123
rect 1599 117 1603 118
rect 1631 122 1635 123
rect 1672 118 1674 125
rect 1694 124 1700 125
rect 1694 120 1695 124
rect 1699 120 1700 124
rect 1694 119 1700 120
rect 1631 117 1635 118
rect 1670 117 1676 118
rect 1078 116 1084 117
rect 1078 112 1079 116
rect 1083 112 1084 116
rect 1078 111 1084 112
rect 1214 116 1220 117
rect 1214 112 1215 116
rect 1219 112 1220 116
rect 1214 111 1220 112
rect 1350 116 1356 117
rect 1350 112 1351 116
rect 1355 112 1356 116
rect 1350 111 1356 112
rect 1486 116 1492 117
rect 1486 112 1487 116
rect 1491 112 1492 116
rect 1486 111 1492 112
rect 1598 116 1604 117
rect 1598 112 1599 116
rect 1603 112 1604 116
rect 1598 111 1604 112
rect 1632 110 1634 117
rect 1670 113 1671 117
rect 1675 113 1676 117
rect 1670 112 1676 113
rect 1630 109 1636 110
rect 1630 105 1631 109
rect 1635 105 1636 109
rect 1630 104 1636 105
rect 1670 99 1676 100
rect 1022 95 1028 96
rect 546 90 552 91
rect 702 91 708 92
rect 146 86 152 87
rect 190 87 196 88
rect 111 82 115 83
rect 134 82 140 83
rect 190 83 191 87
rect 195 83 196 87
rect 190 82 196 83
rect 286 87 292 88
rect 286 83 287 87
rect 291 83 292 87
rect 286 82 292 83
rect 382 87 388 88
rect 382 83 383 87
rect 387 83 388 87
rect 382 82 388 83
rect 478 87 484 88
rect 478 83 479 87
rect 483 83 484 87
rect 478 82 484 83
rect 582 87 588 88
rect 582 83 583 87
rect 587 83 588 87
rect 582 82 588 83
rect 694 87 700 88
rect 694 83 695 87
rect 699 83 700 87
rect 702 87 703 91
rect 707 87 708 91
rect 1022 91 1023 95
rect 1027 91 1028 95
rect 1670 95 1671 99
rect 1675 95 1676 99
rect 1670 94 1676 95
rect 1694 95 1700 96
rect 1022 90 1028 91
rect 1630 91 1636 92
rect 1672 91 1674 94
rect 1694 91 1695 95
rect 1699 91 1700 95
rect 702 86 708 87
rect 814 87 820 88
rect 694 82 700 83
rect 814 83 815 87
rect 819 83 820 87
rect 814 82 820 83
rect 942 87 948 88
rect 942 83 943 87
rect 947 83 948 87
rect 942 82 948 83
rect 1078 87 1084 88
rect 1078 83 1079 87
rect 1083 83 1084 87
rect 1078 82 1084 83
rect 1214 87 1220 88
rect 1214 83 1215 87
rect 1219 83 1220 87
rect 1214 82 1220 83
rect 1350 87 1356 88
rect 1350 83 1351 87
rect 1355 83 1356 87
rect 1350 82 1356 83
rect 1486 87 1492 88
rect 1486 83 1487 87
rect 1491 83 1492 87
rect 1486 82 1492 83
rect 1598 87 1604 88
rect 1598 83 1599 87
rect 1603 83 1604 87
rect 1630 87 1631 91
rect 1635 87 1636 91
rect 1630 86 1636 87
rect 1671 90 1675 91
rect 1694 90 1700 91
rect 1632 83 1634 86
rect 1671 85 1675 86
rect 1752 88 1754 170
rect 1870 152 1876 153
rect 1870 148 1871 152
rect 1875 148 1876 152
rect 1870 147 1876 148
rect 1998 152 2004 153
rect 1998 148 1999 152
rect 2003 148 2004 152
rect 1998 147 2004 148
rect 2142 152 2148 153
rect 2142 148 2143 152
rect 2147 148 2148 152
rect 2142 147 2148 148
rect 2310 152 2316 153
rect 2310 148 2311 152
rect 2315 148 2316 152
rect 2310 147 2316 148
rect 1872 131 1874 147
rect 2000 131 2002 147
rect 2144 131 2146 147
rect 2312 131 2314 147
rect 1815 130 1819 131
rect 1815 125 1819 126
rect 1871 130 1875 131
rect 1871 125 1875 126
rect 1943 130 1947 131
rect 1943 125 1947 126
rect 1999 130 2003 131
rect 1999 125 2003 126
rect 2071 130 2075 131
rect 2071 125 2075 126
rect 2143 130 2147 131
rect 2143 125 2147 126
rect 2199 130 2203 131
rect 2199 125 2203 126
rect 2311 130 2315 131
rect 2311 125 2315 126
rect 2351 130 2355 131
rect 2351 125 2355 126
rect 1814 124 1820 125
rect 1814 120 1815 124
rect 1819 120 1820 124
rect 1814 119 1820 120
rect 1942 124 1948 125
rect 1942 120 1943 124
rect 1947 120 1948 124
rect 1942 119 1948 120
rect 2070 124 2076 125
rect 2070 120 2071 124
rect 2075 120 2076 124
rect 2070 119 2076 120
rect 2198 124 2204 125
rect 2198 120 2199 124
rect 2203 120 2204 124
rect 2198 119 2204 120
rect 2350 124 2356 125
rect 2350 120 2351 124
rect 2355 120 2356 124
rect 2350 119 2356 120
rect 2360 100 2362 174
rect 2494 152 2500 153
rect 2494 148 2495 152
rect 2499 148 2500 152
rect 2494 147 2500 148
rect 2496 131 2498 147
rect 2495 130 2499 131
rect 2495 125 2499 126
rect 2519 130 2523 131
rect 2519 125 2523 126
rect 2518 124 2524 125
rect 2518 120 2519 124
rect 2523 120 2524 124
rect 2518 119 2524 120
rect 2528 100 2530 274
rect 2550 256 2556 257
rect 2550 252 2551 256
rect 2555 252 2556 256
rect 2550 251 2556 252
rect 2662 256 2668 257
rect 2662 252 2663 256
rect 2667 252 2668 256
rect 2662 251 2668 252
rect 2552 239 2554 251
rect 2664 239 2666 251
rect 2551 238 2555 239
rect 2551 233 2555 234
rect 2583 238 2587 239
rect 2583 233 2587 234
rect 2663 238 2667 239
rect 2663 233 2667 234
rect 2582 232 2588 233
rect 2582 228 2583 232
rect 2587 228 2588 232
rect 2582 227 2588 228
rect 2582 203 2588 204
rect 2582 199 2583 203
rect 2587 199 2588 203
rect 2582 198 2588 199
rect 2590 203 2596 204
rect 2590 199 2591 203
rect 2595 199 2596 203
rect 2590 198 2596 199
rect 2584 187 2586 198
rect 2583 186 2587 187
rect 2583 181 2587 182
rect 2592 180 2594 198
rect 2703 186 2707 187
rect 2702 181 2708 182
rect 2590 179 2596 180
rect 2590 175 2591 179
rect 2595 175 2596 179
rect 2702 177 2703 181
rect 2707 177 2708 181
rect 2720 180 2722 278
rect 2782 256 2788 257
rect 2782 252 2783 256
rect 2787 252 2788 256
rect 2782 251 2788 252
rect 2784 239 2786 251
rect 2767 238 2771 239
rect 2767 233 2771 234
rect 2783 238 2787 239
rect 2783 233 2787 234
rect 2766 232 2772 233
rect 2766 228 2767 232
rect 2771 228 2772 232
rect 2766 227 2772 228
rect 2792 208 2794 278
rect 2928 212 2930 302
rect 3022 299 3023 303
rect 3027 299 3028 303
rect 3034 303 3035 307
rect 3039 303 3040 307
rect 3166 307 3172 308
rect 3034 302 3040 303
rect 3158 303 3164 304
rect 3022 298 3028 299
rect 3158 299 3159 303
rect 3163 299 3164 303
rect 3166 303 3167 307
rect 3171 303 3172 307
rect 3166 302 3172 303
rect 3190 307 3196 308
rect 3190 303 3191 307
rect 3195 303 3196 307
rect 3190 302 3196 303
rect 3158 298 3164 299
rect 3024 291 3026 298
rect 3160 291 3162 298
rect 3023 290 3027 291
rect 3023 285 3027 286
rect 3159 290 3163 291
rect 3159 285 3163 286
rect 2967 238 2971 239
rect 2967 233 2971 234
rect 3159 238 3163 239
rect 3159 233 3163 234
rect 2966 232 2972 233
rect 2966 228 2967 232
rect 2971 228 2972 232
rect 2966 227 2972 228
rect 3158 232 3164 233
rect 3158 228 3159 232
rect 3163 228 3164 232
rect 3158 227 3164 228
rect 2926 211 2932 212
rect 2790 207 2796 208
rect 2766 203 2772 204
rect 2766 199 2767 203
rect 2771 199 2772 203
rect 2790 203 2791 207
rect 2795 203 2796 207
rect 2926 207 2927 211
rect 2931 207 2932 211
rect 3168 208 3170 302
rect 3192 291 3194 302
rect 3191 290 3195 291
rect 3191 285 3195 286
rect 3192 282 3194 285
rect 3190 281 3196 282
rect 3190 277 3191 281
rect 3195 277 3196 281
rect 3190 276 3196 277
rect 3190 263 3196 264
rect 3190 259 3191 263
rect 3195 259 3196 263
rect 3190 258 3196 259
rect 3192 239 3194 258
rect 3191 238 3195 239
rect 3191 233 3195 234
rect 3192 226 3194 233
rect 3190 225 3196 226
rect 3190 221 3191 225
rect 3195 221 3196 225
rect 3190 220 3196 221
rect 2926 206 2932 207
rect 3166 207 3172 208
rect 2790 202 2796 203
rect 2766 198 2772 199
rect 2768 187 2770 198
rect 2767 186 2771 187
rect 2919 186 2923 187
rect 2767 181 2771 182
rect 2918 181 2924 182
rect 2702 176 2708 177
rect 2714 179 2722 180
rect 2590 174 2596 175
rect 2714 175 2715 179
rect 2719 175 2722 179
rect 2918 177 2919 181
rect 2923 177 2924 181
rect 2928 180 2930 206
rect 2966 203 2972 204
rect 2966 199 2967 203
rect 2971 199 2972 203
rect 2966 198 2972 199
rect 3158 203 3164 204
rect 3158 199 3159 203
rect 3163 199 3164 203
rect 3166 203 3167 207
rect 3171 203 3172 207
rect 3166 202 3172 203
rect 3190 207 3196 208
rect 3190 203 3191 207
rect 3195 203 3196 207
rect 3190 202 3196 203
rect 3158 198 3164 199
rect 2968 187 2970 198
rect 3160 187 3162 198
rect 2967 186 2971 187
rect 3135 186 3139 187
rect 3159 186 3163 187
rect 2967 181 2971 182
rect 3134 181 3140 182
rect 3159 181 3163 182
rect 2918 176 2924 177
rect 2926 179 2932 180
rect 2714 174 2722 175
rect 2926 175 2927 179
rect 2931 175 2932 179
rect 3134 177 3135 181
rect 3139 177 3140 181
rect 3168 180 3170 202
rect 3192 187 3194 202
rect 3191 186 3195 187
rect 3191 181 3195 182
rect 3134 176 3140 177
rect 3142 179 3148 180
rect 2926 174 2932 175
rect 3142 175 3143 179
rect 3147 175 3148 179
rect 3142 174 3148 175
rect 3166 179 3172 180
rect 3166 175 3167 179
rect 3171 175 3172 179
rect 3192 178 3194 181
rect 3166 174 3172 175
rect 3190 177 3196 178
rect 2702 152 2708 153
rect 2702 148 2703 152
rect 2707 148 2708 152
rect 2702 147 2708 148
rect 2704 131 2706 147
rect 2703 130 2707 131
rect 2703 125 2707 126
rect 2711 130 2715 131
rect 2711 125 2715 126
rect 2710 124 2716 125
rect 2710 120 2711 124
rect 2715 120 2716 124
rect 2710 119 2716 120
rect 2720 100 2722 174
rect 2918 152 2924 153
rect 2918 148 2919 152
rect 2923 148 2924 152
rect 2918 147 2924 148
rect 2920 131 2922 147
rect 2911 130 2915 131
rect 2911 125 2915 126
rect 2919 130 2923 131
rect 2919 125 2923 126
rect 2910 124 2916 125
rect 2910 120 2911 124
rect 2915 120 2916 124
rect 2910 119 2916 120
rect 2358 99 2364 100
rect 1814 95 1820 96
rect 1814 91 1815 95
rect 1819 91 1820 95
rect 1814 90 1820 91
rect 1942 95 1948 96
rect 1942 91 1943 95
rect 1947 91 1948 95
rect 1942 90 1948 91
rect 2070 95 2076 96
rect 2070 91 2071 95
rect 2075 91 2076 95
rect 2070 90 2076 91
rect 2198 95 2204 96
rect 2198 91 2199 95
rect 2203 91 2204 95
rect 2198 90 2204 91
rect 2350 95 2356 96
rect 2350 91 2351 95
rect 2355 91 2356 95
rect 2358 95 2359 99
rect 2363 95 2364 99
rect 2526 99 2532 100
rect 2358 94 2364 95
rect 2518 95 2524 96
rect 2350 90 2356 91
rect 2518 91 2519 95
rect 2523 91 2524 95
rect 2526 95 2527 99
rect 2531 95 2532 99
rect 2718 99 2724 100
rect 2526 94 2532 95
rect 2710 95 2716 96
rect 2518 90 2524 91
rect 2710 91 2711 95
rect 2715 91 2716 95
rect 2718 95 2719 99
rect 2723 95 2724 99
rect 2919 99 2925 100
rect 2718 94 2724 95
rect 2910 95 2916 96
rect 2710 90 2716 91
rect 2910 91 2911 95
rect 2915 91 2916 95
rect 2919 95 2920 99
rect 2924 98 2925 99
rect 2928 98 2930 174
rect 3134 152 3140 153
rect 3134 148 3135 152
rect 3139 148 3140 152
rect 3134 147 3140 148
rect 3136 131 3138 147
rect 3111 130 3115 131
rect 3111 125 3115 126
rect 3135 130 3139 131
rect 3135 125 3139 126
rect 3110 124 3116 125
rect 3110 120 3111 124
rect 3115 120 3116 124
rect 3110 119 3116 120
rect 3144 100 3146 174
rect 3190 173 3191 177
rect 3195 173 3196 177
rect 3190 172 3196 173
rect 3190 159 3196 160
rect 3190 155 3191 159
rect 3195 155 3196 159
rect 3190 154 3196 155
rect 3192 131 3194 154
rect 3191 130 3195 131
rect 3191 125 3195 126
rect 3192 118 3194 125
rect 3190 117 3196 118
rect 3190 113 3191 117
rect 3195 113 3196 117
rect 3190 112 3196 113
rect 2924 96 2930 98
rect 3142 99 3148 100
rect 2924 95 2925 96
rect 2919 94 2925 95
rect 3110 95 3116 96
rect 2910 90 2916 91
rect 3110 91 3111 95
rect 3115 91 3116 95
rect 3142 95 3143 99
rect 3147 95 3148 99
rect 3142 94 3148 95
rect 3190 99 3196 100
rect 3190 95 3191 99
rect 3195 95 3196 99
rect 3190 94 3196 95
rect 3192 91 3194 94
rect 3110 90 3116 91
rect 3191 90 3195 91
rect 1695 85 1699 86
rect 1750 87 1756 88
rect 1750 83 1751 87
rect 1755 83 1756 87
rect 1815 85 1819 86
rect 1943 85 1947 86
rect 2071 85 2075 86
rect 2199 85 2203 86
rect 2351 85 2355 86
rect 2519 85 2523 86
rect 2711 85 2715 86
rect 2911 85 2915 86
rect 3111 85 3115 86
rect 3191 85 3195 86
rect 1598 82 1604 83
rect 1631 82 1635 83
rect 1750 82 1756 83
rect 111 77 115 78
rect 135 77 139 78
rect 191 77 195 78
rect 287 77 291 78
rect 383 77 387 78
rect 479 77 483 78
rect 583 77 587 78
rect 695 77 699 78
rect 815 77 819 78
rect 943 77 947 78
rect 1079 77 1083 78
rect 1215 77 1219 78
rect 1351 77 1355 78
rect 1487 77 1491 78
rect 1599 77 1603 78
rect 1631 77 1635 78
<< m4c >>
rect 1671 3306 1675 3310
rect 3055 3306 3059 3310
rect 3191 3306 3195 3310
rect 1671 3266 1675 3270
rect 2151 3266 2155 3270
rect 2287 3266 2291 3270
rect 2423 3266 2427 3270
rect 2567 3266 2571 3270
rect 2711 3266 2715 3270
rect 2855 3266 2859 3270
rect 2999 3266 3003 3270
rect 3055 3266 3059 3270
rect 1671 3226 1675 3230
rect 1999 3226 2003 3230
rect 2151 3226 2155 3230
rect 2175 3226 2179 3230
rect 2287 3226 2291 3230
rect 2359 3226 2363 3230
rect 2423 3226 2427 3230
rect 2543 3226 2547 3230
rect 2567 3226 2571 3230
rect 2711 3226 2715 3230
rect 2727 3226 2731 3230
rect 2855 3226 2859 3230
rect 2919 3226 2923 3230
rect 2999 3226 3003 3230
rect 3111 3226 3115 3230
rect 1671 3186 1675 3190
rect 1847 3186 1851 3190
rect 1999 3186 2003 3190
rect 2039 3186 2043 3190
rect 2175 3186 2179 3190
rect 2247 3186 2251 3190
rect 2359 3186 2363 3190
rect 2463 3186 2467 3190
rect 2543 3186 2547 3190
rect 3191 3266 3195 3270
rect 3191 3226 3195 3230
rect 2695 3186 2699 3190
rect 2727 3186 2731 3190
rect 2919 3186 2923 3190
rect 1671 3146 1675 3150
rect 1695 3146 1699 3150
rect 1847 3146 1851 3150
rect 111 3126 115 3130
rect 807 3126 811 3130
rect 1079 3126 1083 3130
rect 1351 3126 1355 3130
rect 1599 3126 1603 3130
rect 1631 3126 1635 3130
rect 1863 3146 1867 3150
rect 2023 3146 2027 3150
rect 2039 3146 2043 3150
rect 2935 3186 2939 3190
rect 3111 3186 3115 3190
rect 3159 3186 3163 3190
rect 3191 3186 3195 3190
rect 2183 3146 2187 3150
rect 111 3082 115 3086
rect 703 3082 707 3086
rect 807 3082 811 3086
rect 831 3082 835 3086
rect 959 3082 963 3086
rect 1079 3082 1083 3086
rect 1199 3082 1203 3086
rect 1311 3082 1315 3086
rect 111 3034 115 3038
rect 623 3034 627 3038
rect 703 3034 707 3038
rect 783 3034 787 3038
rect 831 3034 835 3038
rect 927 3034 931 3038
rect 959 3034 963 3038
rect 1063 3034 1067 3038
rect 1079 3034 1083 3038
rect 1191 3034 1195 3038
rect 1199 3034 1203 3038
rect 111 2990 115 2994
rect 519 2990 523 2994
rect 623 2990 627 2994
rect 647 2990 651 2994
rect 783 2990 787 2994
rect 919 2990 923 2994
rect 927 2990 931 2994
rect 111 2942 115 2946
rect 439 2942 443 2946
rect 519 2942 523 2946
rect 599 2942 603 2946
rect 647 2942 651 2946
rect 759 2942 763 2946
rect 783 2942 787 2946
rect 1055 2990 1059 2994
rect 1063 2990 1067 2994
rect 1311 3034 1315 3038
rect 1671 3106 1675 3110
rect 1695 3106 1699 3110
rect 1351 3082 1355 3086
rect 1423 3082 1427 3086
rect 1543 3082 1547 3086
rect 1599 3082 1603 3086
rect 1631 3082 1635 3086
rect 2247 3146 2251 3150
rect 2343 3146 2347 3150
rect 2463 3146 2467 3150
rect 2511 3146 2515 3150
rect 2695 3146 2699 3150
rect 1863 3106 1867 3110
rect 1959 3106 1963 3110
rect 2023 3106 2027 3110
rect 2183 3106 2187 3110
rect 2343 3106 2347 3110
rect 2415 3106 2419 3110
rect 2511 3106 2515 3110
rect 2655 3106 2659 3110
rect 2903 3106 2907 3110
rect 2935 3146 2939 3150
rect 3159 3146 3163 3150
rect 3191 3146 3195 3150
rect 3159 3106 3163 3110
rect 3191 3106 3195 3110
rect 1671 3066 1675 3070
rect 1423 3034 1427 3038
rect 1439 3034 1443 3038
rect 1543 3034 1547 3038
rect 1631 3034 1635 3038
rect 1191 2990 1195 2994
rect 1311 2990 1315 2994
rect 1335 2990 1339 2994
rect 919 2942 923 2946
rect 927 2942 931 2946
rect 1439 2990 1443 2994
rect 1055 2942 1059 2946
rect 1095 2942 1099 2946
rect 1191 2942 1195 2946
rect 1263 2942 1267 2946
rect 1335 2942 1339 2946
rect 1439 2942 1443 2946
rect 1671 3026 1675 3030
rect 1871 3066 1875 3070
rect 1959 3066 1963 3070
rect 2111 3066 2115 3070
rect 2183 3066 2187 3070
rect 2367 3066 2371 3070
rect 2415 3066 2419 3070
rect 2631 3066 2635 3070
rect 2655 3066 2659 3070
rect 2903 3066 2907 3070
rect 1791 3026 1795 3030
rect 1871 3026 1875 3030
rect 3159 3066 3163 3070
rect 3191 3066 3195 3070
rect 1959 3026 1963 3030
rect 2111 3026 2115 3030
rect 2127 3026 2131 3030
rect 2287 3026 2291 3030
rect 2367 3026 2371 3030
rect 2455 3026 2459 3030
rect 2623 3026 2627 3030
rect 2631 3026 2635 3030
rect 2903 3026 2907 3030
rect 1631 2990 1635 2994
rect 1671 2986 1675 2990
rect 1703 2986 1707 2990
rect 1791 2986 1795 2990
rect 1903 2986 1907 2990
rect 1959 2986 1963 2990
rect 2127 2986 2131 2990
rect 1599 2942 1603 2946
rect 1631 2942 1635 2946
rect 1671 2946 1675 2950
rect 1695 2946 1699 2950
rect 1703 2946 1707 2950
rect 2287 2986 2291 2990
rect 1903 2946 1907 2950
rect 1935 2946 1939 2950
rect 2127 2946 2131 2950
rect 2223 2946 2227 2950
rect 2367 2986 2371 2990
rect 2455 2986 2459 2990
rect 2367 2946 2371 2950
rect 2519 2946 2523 2950
rect 2623 2986 2627 2990
rect 2887 2986 2891 2990
rect 3159 3026 3163 3030
rect 3159 2986 3163 2990
rect 3191 3026 3195 3030
rect 3191 2986 3195 2990
rect 2623 2946 2627 2950
rect 2823 2946 2827 2950
rect 2887 2946 2891 2950
rect 3135 2946 3139 2950
rect 3159 2946 3163 2950
rect 3191 2946 3195 2950
rect 111 2902 115 2906
rect 335 2902 339 2906
rect 439 2902 443 2906
rect 471 2902 475 2906
rect 599 2902 603 2906
rect 623 2902 627 2906
rect 759 2902 763 2906
rect 791 2902 795 2906
rect 927 2902 931 2906
rect 111 2854 115 2858
rect 255 2854 259 2858
rect 335 2854 339 2858
rect 415 2854 419 2858
rect 471 2854 475 2858
rect 559 2854 563 2858
rect 623 2854 627 2858
rect 695 2854 699 2858
rect 791 2854 795 2858
rect 823 2854 827 2858
rect 975 2902 979 2906
rect 1095 2902 1099 2906
rect 951 2854 955 2858
rect 975 2854 979 2858
rect 1175 2902 1179 2906
rect 1263 2902 1267 2906
rect 1383 2902 1387 2906
rect 1439 2902 1443 2906
rect 1591 2902 1595 2906
rect 1599 2902 1603 2906
rect 1631 2902 1635 2906
rect 1671 2906 1675 2910
rect 1695 2906 1699 2910
rect 1935 2906 1939 2910
rect 2223 2906 2227 2910
rect 1087 2854 1091 2858
rect 1175 2854 1179 2858
rect 111 2806 115 2810
rect 151 2806 155 2810
rect 255 2806 259 2810
rect 279 2806 283 2810
rect 399 2806 403 2810
rect 415 2806 419 2810
rect 519 2806 523 2810
rect 559 2806 563 2810
rect 639 2806 643 2810
rect 695 2806 699 2810
rect 751 2806 755 2810
rect 823 2806 827 2810
rect 863 2806 867 2810
rect 951 2806 955 2810
rect 983 2806 987 2810
rect 1087 2806 1091 2810
rect 111 2754 115 2758
rect 135 2754 139 2758
rect 151 2754 155 2758
rect 263 2754 267 2758
rect 279 2754 283 2758
rect 399 2754 403 2758
rect 431 2754 435 2758
rect 519 2754 523 2758
rect 623 2754 627 2758
rect 639 2754 643 2758
rect 751 2754 755 2758
rect 839 2754 843 2758
rect 863 2754 867 2758
rect 111 2702 115 2706
rect 135 2702 139 2706
rect 263 2702 267 2706
rect 431 2702 435 2706
rect 623 2702 627 2706
rect 703 2702 707 2706
rect 831 2702 835 2706
rect 839 2702 843 2706
rect 959 2702 963 2706
rect 983 2754 987 2758
rect 1071 2754 1075 2758
rect 1319 2754 1323 2758
rect 1383 2854 1387 2858
rect 1591 2854 1595 2858
rect 1567 2754 1571 2758
rect 1671 2866 1675 2870
rect 2207 2866 2211 2870
rect 1631 2854 1635 2858
rect 1671 2818 1675 2822
rect 2127 2818 2131 2822
rect 2207 2818 2211 2822
rect 1631 2806 1635 2810
rect 1671 2778 1675 2782
rect 2039 2778 2043 2782
rect 2127 2778 2131 2782
rect 2207 2778 2211 2782
rect 2295 2906 2299 2910
rect 2519 2906 2523 2910
rect 2551 2906 2555 2910
rect 2815 2906 2819 2910
rect 2823 2906 2827 2910
rect 2295 2866 2299 2870
rect 2375 2866 2379 2870
rect 2535 2866 2539 2870
rect 3079 2906 3083 2910
rect 3135 2906 3139 2910
rect 2551 2866 2555 2870
rect 2679 2866 2683 2870
rect 2815 2866 2819 2870
rect 2823 2866 2827 2870
rect 2967 2866 2971 2870
rect 3079 2866 3083 2870
rect 3111 2866 3115 2870
rect 3191 2906 3195 2910
rect 3191 2866 3195 2870
rect 2303 2818 2307 2822
rect 2375 2818 2379 2822
rect 2479 2818 2483 2822
rect 2535 2818 2539 2822
rect 2655 2818 2659 2822
rect 2679 2818 2683 2822
rect 2823 2818 2827 2822
rect 2831 2818 2835 2822
rect 2967 2818 2971 2822
rect 3007 2818 3011 2822
rect 3111 2818 3115 2822
rect 3159 2818 3163 2822
rect 3191 2818 3195 2822
rect 2303 2778 2307 2782
rect 1631 2754 1635 2758
rect 1071 2702 1075 2706
rect 1079 2702 1083 2706
rect 111 2654 115 2658
rect 607 2654 611 2658
rect 703 2654 707 2658
rect 735 2654 739 2658
rect 1199 2702 1203 2706
rect 1311 2702 1315 2706
rect 1319 2702 1323 2706
rect 1423 2702 1427 2706
rect 1543 2702 1547 2706
rect 1567 2702 1571 2706
rect 1671 2734 1675 2738
rect 2015 2734 2019 2738
rect 1631 2702 1635 2706
rect 2039 2734 2043 2738
rect 2199 2734 2203 2738
rect 2207 2734 2211 2738
rect 1671 2686 1675 2690
rect 1999 2686 2003 2690
rect 2015 2686 2019 2690
rect 2175 2686 2179 2690
rect 2199 2686 2203 2690
rect 2375 2778 2379 2782
rect 2479 2778 2483 2782
rect 2535 2778 2539 2782
rect 2655 2778 2659 2782
rect 2703 2778 2707 2782
rect 2831 2778 2835 2782
rect 2871 2778 2875 2782
rect 3007 2778 3011 2782
rect 2375 2734 2379 2738
rect 2383 2734 2387 2738
rect 2535 2734 2539 2738
rect 2575 2734 2579 2738
rect 2703 2734 2707 2738
rect 2775 2734 2779 2738
rect 2871 2734 2875 2738
rect 2975 2734 2979 2738
rect 2359 2686 2363 2690
rect 2383 2686 2387 2690
rect 831 2654 835 2658
rect 855 2654 859 2658
rect 959 2654 963 2658
rect 975 2654 979 2658
rect 1079 2654 1083 2658
rect 1095 2654 1099 2658
rect 1199 2654 1203 2658
rect 1207 2654 1211 2658
rect 1311 2654 1315 2658
rect 1319 2654 1323 2658
rect 1423 2654 1427 2658
rect 1439 2654 1443 2658
rect 1543 2654 1547 2658
rect 1631 2654 1635 2658
rect 111 2602 115 2606
rect 503 2602 507 2606
rect 607 2602 611 2606
rect 631 2602 635 2606
rect 735 2602 739 2606
rect 751 2602 755 2606
rect 855 2602 859 2606
rect 871 2602 875 2606
rect 975 2602 979 2606
rect 991 2602 995 2606
rect 1095 2602 1099 2606
rect 1103 2602 1107 2606
rect 1207 2602 1211 2606
rect 1215 2602 1219 2606
rect 1319 2602 1323 2606
rect 1335 2602 1339 2606
rect 1671 2646 1675 2650
rect 1911 2646 1915 2650
rect 1999 2646 2003 2650
rect 1439 2602 1443 2606
rect 1631 2602 1635 2606
rect 1671 2606 1675 2610
rect 1823 2606 1827 2610
rect 1911 2606 1915 2610
rect 2103 2646 2107 2650
rect 2175 2646 2179 2650
rect 2015 2606 2019 2610
rect 2103 2606 2107 2610
rect 2295 2646 2299 2650
rect 2359 2646 2363 2650
rect 2215 2606 2219 2610
rect 2295 2606 2299 2610
rect 111 2550 115 2554
rect 399 2550 403 2554
rect 503 2550 507 2554
rect 527 2550 531 2554
rect 631 2550 635 2554
rect 655 2550 659 2554
rect 751 2550 755 2554
rect 775 2550 779 2554
rect 871 2550 875 2554
rect 895 2550 899 2554
rect 991 2550 995 2554
rect 1007 2550 1011 2554
rect 1103 2550 1107 2554
rect 1119 2550 1123 2554
rect 1215 2550 1219 2554
rect 1239 2550 1243 2554
rect 1671 2562 1675 2566
rect 1735 2562 1739 2566
rect 1823 2562 1827 2566
rect 1335 2550 1339 2554
rect 1631 2550 1635 2554
rect 111 2498 115 2502
rect 303 2498 307 2502
rect 399 2498 403 2502
rect 431 2498 435 2502
rect 527 2498 531 2502
rect 559 2498 563 2502
rect 655 2498 659 2502
rect 703 2498 707 2502
rect 775 2498 779 2502
rect 863 2498 867 2502
rect 895 2498 899 2502
rect 1007 2498 1011 2502
rect 1039 2498 1043 2502
rect 1119 2498 1123 2502
rect 1223 2498 1227 2502
rect 1239 2498 1243 2502
rect 1671 2518 1675 2522
rect 1695 2518 1699 2522
rect 1735 2518 1739 2522
rect 1895 2562 1899 2566
rect 2015 2562 2019 2566
rect 2055 2562 2059 2566
rect 2215 2562 2219 2566
rect 1863 2518 1867 2522
rect 1895 2518 1899 2522
rect 2055 2518 2059 2522
rect 2079 2518 2083 2522
rect 2215 2518 2219 2522
rect 2319 2518 2323 2522
rect 2439 2606 2443 2610
rect 2551 2686 2555 2690
rect 3159 2778 3163 2782
rect 3159 2734 3163 2738
rect 3191 2778 3195 2782
rect 3191 2734 3195 2738
rect 2575 2686 2579 2690
rect 2759 2686 2763 2690
rect 2775 2686 2779 2690
rect 2967 2686 2971 2690
rect 2975 2686 2979 2690
rect 3159 2686 3163 2690
rect 3191 2686 3195 2690
rect 2487 2646 2491 2650
rect 2551 2646 2555 2650
rect 2687 2646 2691 2650
rect 2759 2646 2763 2650
rect 2487 2606 2491 2610
rect 2671 2606 2675 2610
rect 2687 2606 2691 2610
rect 2919 2606 2923 2610
rect 2967 2646 2971 2650
rect 3159 2646 3163 2650
rect 3159 2606 3163 2610
rect 3191 2646 3195 2650
rect 3191 2606 3195 2610
rect 2375 2562 2379 2566
rect 2439 2562 2443 2566
rect 2535 2562 2539 2566
rect 2671 2562 2675 2566
rect 2919 2562 2923 2566
rect 2375 2518 2379 2522
rect 2535 2518 2539 2522
rect 2583 2518 2587 2522
rect 2855 2518 2859 2522
rect 1423 2498 1427 2502
rect 1599 2498 1603 2502
rect 1631 2498 1635 2502
rect 111 2454 115 2458
rect 199 2454 203 2458
rect 303 2454 307 2458
rect 327 2454 331 2458
rect 431 2454 435 2458
rect 455 2454 459 2458
rect 559 2454 563 2458
rect 599 2454 603 2458
rect 703 2454 707 2458
rect 767 2454 771 2458
rect 863 2454 867 2458
rect 951 2454 955 2458
rect 1039 2454 1043 2458
rect 1159 2454 1163 2458
rect 1223 2454 1227 2458
rect 1375 2454 1379 2458
rect 1423 2454 1427 2458
rect 111 2398 115 2402
rect 135 2398 139 2402
rect 199 2398 203 2402
rect 239 2398 243 2402
rect 327 2398 331 2402
rect 359 2398 363 2402
rect 455 2398 459 2402
rect 479 2398 483 2402
rect 591 2398 595 2402
rect 599 2398 603 2402
rect 703 2398 707 2402
rect 767 2398 771 2402
rect 815 2398 819 2402
rect 935 2398 939 2402
rect 951 2398 955 2402
rect 1159 2398 1163 2402
rect 111 2350 115 2354
rect 135 2350 139 2354
rect 239 2350 243 2354
rect 343 2350 347 2354
rect 359 2350 363 2354
rect 479 2350 483 2354
rect 567 2350 571 2354
rect 591 2350 595 2354
rect 703 2350 707 2354
rect 775 2350 779 2354
rect 815 2350 819 2354
rect 935 2350 939 2354
rect 111 2298 115 2302
rect 135 2298 139 2302
rect 111 2246 115 2250
rect 111 2198 115 2202
rect 111 2146 115 2150
rect 111 2094 115 2098
rect 111 2046 115 2050
rect 175 2046 179 2050
rect 343 2298 347 2302
rect 567 2298 571 2302
rect 551 2246 555 2250
rect 655 2298 659 2302
rect 775 2298 779 2302
rect 783 2298 787 2302
rect 903 2298 907 2302
rect 975 2350 979 2354
rect 1175 2350 1179 2354
rect 1375 2398 1379 2402
rect 1367 2350 1371 2354
rect 1567 2350 1571 2354
rect 1671 2470 1675 2474
rect 1695 2470 1699 2474
rect 1863 2470 1867 2474
rect 2079 2470 2083 2474
rect 2319 2470 2323 2474
rect 1591 2454 1595 2458
rect 1599 2454 1603 2458
rect 1631 2454 1635 2458
rect 2567 2470 2571 2474
rect 3135 2518 3139 2522
rect 3159 2562 3163 2566
rect 3191 2562 3195 2566
rect 3191 2518 3195 2522
rect 2583 2470 2587 2474
rect 2823 2470 2827 2474
rect 2855 2470 2859 2474
rect 1671 2430 1675 2434
rect 2231 2430 2235 2434
rect 2319 2430 2323 2434
rect 2391 2430 2395 2434
rect 2543 2430 2547 2434
rect 2567 2430 2571 2434
rect 2687 2430 2691 2434
rect 2823 2430 2827 2434
rect 2967 2430 2971 2434
rect 3079 2470 3083 2474
rect 3135 2470 3139 2474
rect 3079 2430 3083 2434
rect 3111 2430 3115 2434
rect 3191 2470 3195 2474
rect 3191 2430 3195 2434
rect 1591 2398 1595 2402
rect 1631 2398 1635 2402
rect 1671 2382 1675 2386
rect 2143 2382 2147 2386
rect 2231 2382 2235 2386
rect 2311 2382 2315 2386
rect 2391 2382 2395 2386
rect 2479 2382 2483 2386
rect 2543 2382 2547 2386
rect 2655 2382 2659 2386
rect 2687 2382 2691 2386
rect 2823 2382 2827 2386
rect 2831 2382 2835 2386
rect 2967 2382 2971 2386
rect 3007 2382 3011 2386
rect 3111 2382 3115 2386
rect 3159 2382 3163 2386
rect 3191 2382 3195 2386
rect 1631 2350 1635 2354
rect 975 2298 979 2302
rect 1023 2298 1027 2302
rect 1143 2298 1147 2302
rect 1175 2298 1179 2302
rect 1255 2298 1259 2302
rect 1367 2298 1371 2302
rect 655 2246 659 2250
rect 679 2246 683 2250
rect 783 2246 787 2250
rect 807 2246 811 2250
rect 903 2246 907 2250
rect 927 2246 931 2250
rect 1023 2246 1027 2250
rect 1047 2246 1051 2250
rect 1143 2246 1147 2250
rect 1159 2246 1163 2250
rect 1671 2342 1675 2346
rect 2143 2342 2147 2346
rect 2183 2342 2187 2346
rect 2311 2342 2315 2346
rect 2335 2342 2339 2346
rect 2479 2342 2483 2346
rect 2623 2342 2627 2346
rect 2655 2342 2659 2346
rect 2767 2342 2771 2346
rect 2831 2342 2835 2346
rect 2919 2342 2923 2346
rect 3007 2342 3011 2346
rect 3159 2342 3163 2346
rect 1487 2298 1491 2302
rect 1567 2298 1571 2302
rect 1631 2298 1635 2302
rect 1671 2298 1675 2302
rect 2095 2298 2099 2302
rect 1255 2246 1259 2250
rect 1271 2246 1275 2250
rect 455 2198 459 2202
rect 551 2198 555 2202
rect 583 2198 587 2202
rect 679 2198 683 2202
rect 703 2198 707 2202
rect 807 2198 811 2202
rect 823 2198 827 2202
rect 927 2198 931 2202
rect 943 2198 947 2202
rect 1367 2246 1371 2250
rect 1391 2246 1395 2250
rect 1671 2258 1675 2262
rect 2015 2258 2019 2262
rect 1487 2246 1491 2250
rect 1631 2246 1635 2250
rect 2095 2258 2099 2262
rect 2167 2258 2171 2262
rect 2183 2298 2187 2302
rect 2263 2298 2267 2302
rect 2335 2298 2339 2302
rect 2431 2298 2435 2302
rect 2479 2298 2483 2302
rect 2607 2298 2611 2302
rect 2623 2298 2627 2302
rect 2767 2298 2771 2302
rect 2791 2298 2795 2302
rect 2919 2298 2923 2302
rect 2983 2298 2987 2302
rect 3159 2298 3163 2302
rect 2263 2258 2267 2262
rect 2319 2258 2323 2262
rect 2431 2258 2435 2262
rect 2463 2258 2467 2262
rect 2607 2258 2611 2262
rect 2759 2258 2763 2262
rect 2791 2258 2795 2262
rect 3191 2342 3195 2346
rect 3191 2298 3195 2302
rect 2983 2258 2987 2262
rect 1047 2198 1051 2202
rect 1055 2198 1059 2202
rect 1159 2198 1163 2202
rect 1167 2198 1171 2202
rect 1271 2198 1275 2202
rect 1671 2214 1675 2218
rect 1927 2214 1931 2218
rect 2015 2214 2019 2218
rect 1287 2198 1291 2202
rect 1391 2198 1395 2202
rect 1631 2198 1635 2202
rect 2103 2214 2107 2218
rect 2167 2214 2171 2218
rect 2295 2214 2299 2218
rect 1671 2174 1675 2178
rect 1847 2174 1851 2178
rect 1927 2174 1931 2178
rect 1999 2174 2003 2178
rect 351 2146 355 2150
rect 455 2146 459 2150
rect 479 2146 483 2150
rect 583 2146 587 2150
rect 599 2146 603 2150
rect 703 2146 707 2150
rect 719 2146 723 2150
rect 823 2146 827 2150
rect 839 2146 843 2150
rect 943 2146 947 2150
rect 951 2146 955 2150
rect 1055 2146 1059 2150
rect 1063 2146 1067 2150
rect 1167 2146 1171 2150
rect 2103 2174 2107 2178
rect 1183 2146 1187 2150
rect 1287 2146 1291 2150
rect 1631 2146 1635 2150
rect 247 2094 251 2098
rect 351 2094 355 2098
rect 375 2094 379 2098
rect 479 2094 483 2098
rect 503 2094 507 2098
rect 599 2094 603 2098
rect 623 2094 627 2098
rect 719 2094 723 2098
rect 743 2094 747 2098
rect 839 2094 843 2098
rect 855 2094 859 2098
rect 951 2094 955 2098
rect 967 2094 971 2098
rect 1063 2094 1067 2098
rect 1671 2130 1675 2134
rect 1759 2130 1763 2134
rect 1847 2130 1851 2134
rect 1911 2130 1915 2134
rect 1999 2130 2003 2134
rect 1087 2094 1091 2098
rect 1183 2094 1187 2098
rect 1631 2094 1635 2098
rect 1671 2090 1675 2094
rect 1695 2090 1699 2094
rect 1759 2090 1763 2094
rect 1823 2090 1827 2094
rect 1911 2090 1915 2094
rect 1967 2090 1971 2094
rect 2071 2130 2075 2134
rect 2151 2174 2155 2178
rect 2319 2214 2323 2218
rect 2463 2214 2467 2218
rect 2503 2214 2507 2218
rect 2607 2214 2611 2218
rect 2719 2214 2723 2218
rect 2759 2214 2763 2218
rect 2951 2214 2955 2218
rect 3159 2258 3163 2262
rect 3159 2214 3163 2218
rect 2295 2174 2299 2178
rect 2447 2174 2451 2178
rect 2503 2174 2507 2178
rect 2599 2174 2603 2178
rect 2719 2174 2723 2178
rect 2151 2130 2155 2134
rect 2255 2130 2259 2134
rect 2295 2130 2299 2134
rect 2447 2130 2451 2134
rect 2463 2130 2467 2134
rect 2599 2130 2603 2134
rect 2687 2130 2691 2134
rect 3191 2258 3195 2262
rect 3191 2214 3195 2218
rect 2951 2174 2955 2178
rect 2927 2130 2931 2134
rect 3159 2174 3163 2178
rect 3159 2130 3163 2134
rect 2071 2090 2075 2094
rect 2111 2090 2115 2094
rect 2255 2090 2259 2094
rect 2407 2090 2411 2094
rect 2463 2090 2467 2094
rect 2687 2090 2691 2094
rect 247 2046 251 2050
rect 111 2006 115 2010
rect 135 2006 139 2010
rect 175 2006 179 2010
rect 231 2006 235 2010
rect 367 2046 371 2050
rect 375 2046 379 2050
rect 503 2046 507 2050
rect 559 2046 563 2050
rect 623 2046 627 2050
rect 743 2046 747 2050
rect 759 2046 763 2050
rect 855 2046 859 2050
rect 351 2006 355 2010
rect 367 2006 371 2010
rect 463 2006 467 2010
rect 559 2006 563 2010
rect 575 2006 579 2010
rect 687 2006 691 2010
rect 759 2006 763 2010
rect 111 1958 115 1962
rect 135 1958 139 1962
rect 111 1906 115 1910
rect 111 1854 115 1858
rect 111 1806 115 1810
rect 111 1754 115 1758
rect 111 1702 115 1706
rect 111 1650 115 1654
rect 135 1650 139 1654
rect 799 2006 803 2010
rect 967 2046 971 2050
rect 1087 2046 1091 2050
rect 1183 2046 1187 2050
rect 1399 2046 1403 2050
rect 1599 2046 1603 2050
rect 1631 2046 1635 2050
rect 1671 2050 1675 2054
rect 1695 2050 1699 2054
rect 1823 2050 1827 2054
rect 1967 2050 1971 2054
rect 911 2006 915 2010
rect 967 2006 971 2010
rect 1183 2006 1187 2010
rect 1399 2006 1403 2010
rect 231 1958 235 1962
rect 351 1958 355 1962
rect 463 1958 467 1962
rect 575 1958 579 1962
rect 687 1958 691 1962
rect 727 1958 731 1962
rect 799 1958 803 1962
rect 855 1958 859 1962
rect 911 1958 915 1962
rect 983 1958 987 1962
rect 1103 1958 1107 1962
rect 1223 1958 1227 1962
rect 1335 1958 1339 1962
rect 1599 2006 1603 2010
rect 1447 1958 1451 1962
rect 1567 1958 1571 1962
rect 2039 2050 2043 2054
rect 2111 2050 2115 2054
rect 1631 2006 1635 2010
rect 1671 2002 1675 2006
rect 1695 2002 1699 2006
rect 2039 2002 2043 2006
rect 2255 2050 2259 2054
rect 2407 2050 2411 2054
rect 3191 2174 3195 2178
rect 3191 2130 3195 2134
rect 2927 2090 2931 2094
rect 3159 2090 3163 2094
rect 2767 2050 2771 2054
rect 3135 2050 3139 2054
rect 2263 2002 2267 2006
rect 2407 2002 2411 2006
rect 2415 2002 2419 2006
rect 2559 2002 2563 2006
rect 2703 2002 2707 2006
rect 2767 2002 2771 2006
rect 2839 2002 2843 2006
rect 1631 1958 1635 1962
rect 1671 1962 1675 1966
rect 2239 1962 2243 1966
rect 631 1906 635 1910
rect 727 1906 731 1910
rect 759 1906 763 1910
rect 855 1906 859 1910
rect 879 1906 883 1910
rect 983 1906 987 1910
rect 999 1906 1003 1910
rect 1103 1906 1107 1910
rect 1119 1906 1123 1910
rect 1223 1906 1227 1910
rect 1231 1906 1235 1910
rect 1335 1906 1339 1910
rect 1343 1906 1347 1910
rect 1447 1906 1451 1910
rect 1463 1906 1467 1910
rect 2263 1962 2267 1966
rect 2391 1962 2395 1966
rect 2415 1962 2419 1966
rect 2975 2002 2979 2006
rect 3111 2002 3115 2006
rect 3135 2002 3139 2006
rect 3191 2090 3195 2094
rect 3191 2050 3195 2054
rect 3191 2002 3195 2006
rect 2543 1962 2547 1966
rect 2559 1962 2563 1966
rect 2695 1962 2699 1966
rect 2703 1962 2707 1966
rect 2839 1962 2843 1966
rect 2847 1962 2851 1966
rect 2975 1962 2979 1966
rect 2999 1962 3003 1966
rect 3111 1962 3115 1966
rect 1671 1918 1675 1922
rect 2151 1918 2155 1922
rect 2239 1918 2243 1922
rect 1567 1906 1571 1910
rect 1631 1906 1635 1910
rect 2311 1918 2315 1922
rect 2391 1918 2395 1922
rect 2471 1918 2475 1922
rect 2543 1918 2547 1922
rect 527 1854 531 1858
rect 631 1854 635 1858
rect 655 1854 659 1858
rect 759 1854 763 1858
rect 775 1854 779 1858
rect 879 1854 883 1858
rect 895 1854 899 1858
rect 999 1854 1003 1858
rect 1015 1854 1019 1858
rect 1119 1854 1123 1858
rect 1127 1854 1131 1858
rect 1231 1854 1235 1858
rect 1247 1854 1251 1858
rect 1343 1854 1347 1858
rect 1671 1874 1675 1878
rect 2071 1874 2075 1878
rect 2151 1874 2155 1878
rect 1367 1854 1371 1858
rect 1463 1854 1467 1858
rect 1631 1854 1635 1858
rect 2239 1874 2243 1878
rect 2311 1874 2315 1878
rect 2415 1874 2419 1878
rect 423 1806 427 1810
rect 527 1806 531 1810
rect 551 1806 555 1810
rect 655 1806 659 1810
rect 679 1806 683 1810
rect 775 1806 779 1810
rect 799 1806 803 1810
rect 895 1806 899 1810
rect 919 1806 923 1810
rect 1015 1806 1019 1810
rect 1031 1806 1035 1810
rect 1127 1806 1131 1810
rect 1143 1806 1147 1810
rect 1247 1806 1251 1810
rect 2471 1874 2475 1878
rect 2639 1918 2643 1922
rect 2695 1918 2699 1922
rect 2815 1918 2819 1922
rect 2847 1918 2851 1922
rect 2999 1918 3003 1922
rect 3159 1918 3163 1922
rect 3191 1962 3195 1966
rect 3191 1918 3195 1922
rect 2599 1874 2603 1878
rect 2639 1874 2643 1878
rect 2791 1874 2795 1878
rect 2815 1874 2819 1878
rect 1671 1834 1675 1838
rect 1983 1834 1987 1838
rect 2071 1834 2075 1838
rect 2135 1834 2139 1838
rect 2239 1834 2243 1838
rect 2983 1874 2987 1878
rect 2999 1874 3003 1878
rect 3159 1874 3163 1878
rect 3191 1874 3195 1878
rect 2287 1834 2291 1838
rect 2415 1834 2419 1838
rect 2431 1834 2435 1838
rect 2583 1834 2587 1838
rect 2599 1834 2603 1838
rect 2735 1834 2739 1838
rect 2791 1834 2795 1838
rect 2983 1834 2987 1838
rect 1263 1806 1267 1810
rect 1367 1806 1371 1810
rect 1631 1806 1635 1810
rect 1671 1794 1675 1798
rect 1903 1794 1907 1798
rect 1983 1794 1987 1798
rect 327 1754 331 1758
rect 423 1754 427 1758
rect 455 1754 459 1758
rect 551 1754 555 1758
rect 2079 1794 2083 1798
rect 2135 1794 2139 1798
rect 2271 1794 2275 1798
rect 2287 1794 2291 1798
rect 2431 1794 2435 1798
rect 2487 1794 2491 1798
rect 575 1754 579 1758
rect 679 1754 683 1758
rect 695 1754 699 1758
rect 799 1754 803 1758
rect 815 1754 819 1758
rect 919 1754 923 1758
rect 927 1754 931 1758
rect 1031 1754 1035 1758
rect 1039 1754 1043 1758
rect 1143 1754 1147 1758
rect 1159 1754 1163 1758
rect 1263 1754 1267 1758
rect 1631 1754 1635 1758
rect 2583 1794 2587 1798
rect 2711 1794 2715 1798
rect 2735 1794 2739 1798
rect 2943 1794 2947 1798
rect 3159 1834 3163 1838
rect 3159 1794 3163 1798
rect 3191 1834 3195 1838
rect 3191 1794 3195 1798
rect 223 1702 227 1706
rect 327 1702 331 1706
rect 223 1650 227 1654
rect 351 1702 355 1706
rect 455 1702 459 1706
rect 471 1702 475 1706
rect 575 1702 579 1706
rect 591 1702 595 1706
rect 695 1702 699 1706
rect 711 1702 715 1706
rect 815 1702 819 1706
rect 823 1702 827 1706
rect 1671 1746 1675 1750
rect 1815 1746 1819 1750
rect 1903 1746 1907 1750
rect 1967 1746 1971 1750
rect 2079 1746 2083 1750
rect 2127 1746 2131 1750
rect 2271 1746 2275 1750
rect 2303 1746 2307 1750
rect 2487 1746 2491 1750
rect 2503 1746 2507 1750
rect 2711 1746 2715 1750
rect 2935 1746 2939 1750
rect 2943 1746 2947 1750
rect 927 1702 931 1706
rect 943 1702 947 1706
rect 247 1650 251 1654
rect 351 1650 355 1654
rect 383 1650 387 1654
rect 471 1650 475 1654
rect 535 1650 539 1654
rect 591 1650 595 1654
rect 711 1650 715 1654
rect 1039 1702 1043 1706
rect 1063 1702 1067 1706
rect 1159 1702 1163 1706
rect 823 1650 827 1654
rect 919 1650 923 1654
rect 111 1602 115 1606
rect 135 1602 139 1606
rect 247 1602 251 1606
rect 303 1602 307 1606
rect 383 1602 387 1606
rect 943 1650 947 1654
rect 1063 1650 1067 1654
rect 503 1602 507 1606
rect 535 1602 539 1606
rect 695 1602 699 1606
rect 711 1602 715 1606
rect 887 1602 891 1606
rect 919 1602 923 1606
rect 1063 1602 1067 1606
rect 1143 1650 1147 1654
rect 3159 1746 3163 1750
rect 3191 1746 3195 1750
rect 1631 1702 1635 1706
rect 1671 1706 1675 1710
rect 1735 1706 1739 1710
rect 1815 1706 1819 1710
rect 1879 1706 1883 1710
rect 1967 1706 1971 1710
rect 2023 1706 2027 1710
rect 2127 1706 2131 1710
rect 2167 1706 2171 1710
rect 2303 1706 2307 1710
rect 2311 1706 2315 1710
rect 2463 1706 2467 1710
rect 2503 1706 2507 1710
rect 2711 1706 2715 1710
rect 1671 1666 1675 1670
rect 1695 1666 1699 1670
rect 1735 1666 1739 1670
rect 1879 1666 1883 1670
rect 1895 1666 1899 1670
rect 2023 1666 2027 1670
rect 2127 1666 2131 1670
rect 2167 1666 2171 1670
rect 2311 1666 2315 1670
rect 2367 1666 2371 1670
rect 2463 1666 2467 1670
rect 2615 1666 2619 1670
rect 2935 1706 2939 1710
rect 3159 1706 3163 1710
rect 2871 1666 2875 1670
rect 3135 1666 3139 1670
rect 3191 1706 3195 1710
rect 3191 1666 3195 1670
rect 1383 1650 1387 1654
rect 1599 1650 1603 1654
rect 1631 1650 1635 1654
rect 1143 1602 1147 1606
rect 1239 1602 1243 1606
rect 1383 1602 1387 1606
rect 1415 1602 1419 1606
rect 111 1550 115 1554
rect 135 1550 139 1554
rect 303 1550 307 1554
rect 503 1550 507 1554
rect 679 1550 683 1554
rect 695 1550 699 1554
rect 807 1550 811 1554
rect 887 1550 891 1554
rect 927 1550 931 1554
rect 1047 1550 1051 1554
rect 1063 1550 1067 1554
rect 1591 1602 1595 1606
rect 1599 1602 1603 1606
rect 1167 1550 1171 1554
rect 1239 1550 1243 1554
rect 1279 1550 1283 1554
rect 1671 1622 1675 1626
rect 1695 1622 1699 1626
rect 1895 1622 1899 1626
rect 1631 1602 1635 1606
rect 1671 1582 1675 1586
rect 1399 1550 1403 1554
rect 1415 1550 1419 1554
rect 1519 1550 1523 1554
rect 1591 1550 1595 1554
rect 1631 1550 1635 1554
rect 111 1502 115 1506
rect 575 1502 579 1506
rect 679 1502 683 1506
rect 703 1502 707 1506
rect 807 1502 811 1506
rect 831 1502 835 1506
rect 927 1502 931 1506
rect 951 1502 955 1506
rect 1047 1502 1051 1506
rect 1071 1502 1075 1506
rect 1167 1502 1171 1506
rect 1183 1502 1187 1506
rect 1279 1502 1283 1506
rect 1295 1502 1299 1506
rect 1399 1502 1403 1506
rect 1671 1534 1675 1538
rect 1415 1502 1419 1506
rect 1519 1502 1523 1506
rect 1631 1502 1635 1506
rect 2127 1622 2131 1626
rect 2319 1622 2323 1626
rect 2367 1622 2371 1626
rect 2271 1582 2275 1586
rect 2319 1582 2323 1586
rect 2167 1534 2171 1538
rect 2271 1534 2275 1538
rect 2279 1534 2283 1538
rect 2519 1622 2523 1626
rect 2615 1622 2619 1626
rect 2711 1622 2715 1626
rect 2871 1622 2875 1626
rect 2911 1622 2915 1626
rect 3111 1622 3115 1626
rect 3135 1622 3139 1626
rect 3191 1622 3195 1626
rect 2415 1582 2419 1586
rect 2519 1582 2523 1586
rect 2559 1582 2563 1586
rect 2695 1582 2699 1586
rect 2711 1582 2715 1586
rect 2839 1582 2843 1586
rect 2911 1582 2915 1586
rect 2983 1582 2987 1586
rect 3111 1582 3115 1586
rect 2391 1534 2395 1538
rect 2415 1534 2419 1538
rect 2503 1534 2507 1538
rect 2559 1534 2563 1538
rect 2615 1534 2619 1538
rect 1671 1490 1675 1494
rect 2087 1490 2091 1494
rect 2167 1490 2171 1494
rect 2231 1490 2235 1494
rect 2279 1490 2283 1494
rect 2695 1534 2699 1538
rect 2735 1534 2739 1538
rect 2839 1534 2843 1538
rect 2855 1534 2859 1538
rect 2983 1534 2987 1538
rect 2375 1490 2379 1494
rect 2391 1490 2395 1494
rect 2503 1490 2507 1494
rect 2511 1490 2515 1494
rect 2615 1490 2619 1494
rect 2655 1490 2659 1494
rect 111 1450 115 1454
rect 479 1450 483 1454
rect 575 1450 579 1454
rect 607 1450 611 1454
rect 703 1450 707 1454
rect 727 1450 731 1454
rect 831 1450 835 1454
rect 847 1450 851 1454
rect 951 1450 955 1454
rect 967 1450 971 1454
rect 1071 1450 1075 1454
rect 1079 1450 1083 1454
rect 1183 1450 1187 1454
rect 1191 1450 1195 1454
rect 1295 1450 1299 1454
rect 1311 1450 1315 1454
rect 1415 1450 1419 1454
rect 1631 1450 1635 1454
rect 1671 1446 1675 1450
rect 1983 1446 1987 1450
rect 2087 1446 2091 1450
rect 2095 1446 2099 1450
rect 111 1398 115 1402
rect 375 1398 379 1402
rect 479 1398 483 1402
rect 503 1398 507 1402
rect 607 1398 611 1402
rect 623 1398 627 1402
rect 727 1398 731 1402
rect 743 1398 747 1402
rect 847 1398 851 1402
rect 863 1398 867 1402
rect 967 1398 971 1402
rect 975 1398 979 1402
rect 1079 1398 1083 1402
rect 1095 1398 1099 1402
rect 2207 1446 2211 1450
rect 2231 1446 2235 1450
rect 2335 1446 2339 1450
rect 2375 1446 2379 1450
rect 1191 1398 1195 1402
rect 1215 1398 1219 1402
rect 1311 1398 1315 1402
rect 1631 1398 1635 1402
rect 2479 1446 2483 1450
rect 2735 1490 2739 1494
rect 2799 1490 2803 1494
rect 3111 1534 3115 1538
rect 3191 1582 3195 1586
rect 3191 1534 3195 1538
rect 2855 1490 2859 1494
rect 2983 1490 2987 1494
rect 2511 1446 2515 1450
rect 2639 1446 2643 1450
rect 2655 1446 2659 1450
rect 2799 1446 2803 1450
rect 2815 1446 2819 1450
rect 2999 1446 3003 1450
rect 3111 1490 3115 1494
rect 3191 1490 3195 1494
rect 3159 1446 3163 1450
rect 3191 1446 3195 1450
rect 1671 1390 1675 1394
rect 1879 1390 1883 1394
rect 1983 1390 1987 1394
rect 1991 1390 1995 1394
rect 2095 1390 2099 1394
rect 2103 1390 2107 1394
rect 2207 1390 2211 1394
rect 2239 1390 2243 1394
rect 2335 1390 2339 1394
rect 2391 1390 2395 1394
rect 2479 1390 2483 1394
rect 2567 1390 2571 1394
rect 2639 1390 2643 1394
rect 2767 1390 2771 1394
rect 2815 1390 2819 1394
rect 2975 1390 2979 1394
rect 2999 1390 3003 1394
rect 3159 1390 3163 1394
rect 3191 1390 3195 1394
rect 111 1350 115 1354
rect 271 1350 275 1354
rect 375 1350 379 1354
rect 399 1350 403 1354
rect 503 1350 507 1354
rect 527 1350 531 1354
rect 623 1350 627 1354
rect 647 1350 651 1354
rect 743 1350 747 1354
rect 767 1350 771 1354
rect 863 1350 867 1354
rect 879 1350 883 1354
rect 975 1350 979 1354
rect 991 1350 995 1354
rect 1095 1350 1099 1354
rect 1111 1350 1115 1354
rect 1215 1350 1219 1354
rect 1631 1350 1635 1354
rect 111 1298 115 1302
rect 175 1298 179 1302
rect 271 1298 275 1302
rect 303 1298 307 1302
rect 399 1298 403 1302
rect 423 1298 427 1302
rect 527 1298 531 1302
rect 543 1298 547 1302
rect 647 1298 651 1302
rect 663 1298 667 1302
rect 767 1298 771 1302
rect 775 1298 779 1302
rect 111 1246 115 1250
rect 135 1246 139 1250
rect 175 1246 179 1250
rect 231 1246 235 1250
rect 303 1246 307 1250
rect 879 1298 883 1302
rect 887 1298 891 1302
rect 1671 1338 1675 1342
rect 991 1298 995 1302
rect 1007 1298 1011 1302
rect 1775 1338 1779 1342
rect 1879 1338 1883 1342
rect 1887 1338 1891 1342
rect 1991 1338 1995 1342
rect 2095 1338 2099 1342
rect 2103 1338 2107 1342
rect 2199 1338 2203 1342
rect 2239 1338 2243 1342
rect 2303 1338 2307 1342
rect 2391 1338 2395 1342
rect 2407 1338 2411 1342
rect 2511 1338 2515 1342
rect 2567 1338 2571 1342
rect 2767 1338 2771 1342
rect 2975 1338 2979 1342
rect 1111 1298 1115 1302
rect 1631 1298 1635 1302
rect 1671 1290 1675 1294
rect 1695 1290 1699 1294
rect 1775 1290 1779 1294
rect 1791 1290 1795 1294
rect 1887 1290 1891 1294
rect 1935 1290 1939 1294
rect 1991 1290 1995 1294
rect 2095 1290 2099 1294
rect 2103 1290 2107 1294
rect 2199 1290 2203 1294
rect 2295 1290 2299 1294
rect 2303 1290 2307 1294
rect 2407 1290 2411 1294
rect 2495 1290 2499 1294
rect 2511 1290 2515 1294
rect 2711 1290 2715 1294
rect 2935 1290 2939 1294
rect 3159 1338 3163 1342
rect 3159 1290 3163 1294
rect 359 1246 363 1250
rect 423 1246 427 1250
rect 503 1246 507 1250
rect 543 1246 547 1250
rect 663 1246 667 1250
rect 775 1246 779 1250
rect 831 1246 835 1250
rect 887 1246 891 1250
rect 1007 1246 1011 1250
rect 1015 1246 1019 1250
rect 1207 1246 1211 1250
rect 1407 1246 1411 1250
rect 1599 1246 1603 1250
rect 1631 1246 1635 1250
rect 1671 1234 1675 1238
rect 111 1198 115 1202
rect 135 1198 139 1202
rect 231 1198 235 1202
rect 111 1146 115 1150
rect 111 1094 115 1098
rect 111 1046 115 1050
rect 111 994 115 998
rect 111 942 115 946
rect 223 942 227 946
rect 359 1198 363 1202
rect 503 1198 507 1202
rect 663 1198 667 1202
rect 631 1146 635 1150
rect 727 1198 731 1202
rect 831 1198 835 1202
rect 855 1198 859 1202
rect 983 1198 987 1202
rect 1015 1198 1019 1202
rect 1103 1198 1107 1202
rect 1207 1198 1211 1202
rect 1223 1198 1227 1202
rect 1335 1198 1339 1202
rect 1407 1198 1411 1202
rect 1447 1198 1451 1202
rect 1695 1234 1699 1238
rect 1567 1198 1571 1202
rect 1599 1198 1603 1202
rect 1791 1234 1795 1238
rect 1935 1234 1939 1238
rect 3191 1338 3195 1342
rect 3191 1290 3195 1294
rect 1983 1234 1987 1238
rect 2103 1234 2107 1238
rect 2255 1234 2259 1238
rect 2295 1234 2299 1238
rect 2495 1234 2499 1238
rect 2711 1234 2715 1238
rect 2919 1234 2923 1238
rect 2935 1234 2939 1238
rect 3135 1234 3139 1238
rect 3159 1234 3163 1238
rect 3191 1234 3195 1238
rect 1631 1198 1635 1202
rect 1671 1190 1675 1194
rect 1695 1190 1699 1194
rect 1983 1190 1987 1194
rect 2247 1190 2251 1194
rect 2255 1190 2259 1194
rect 2399 1190 2403 1194
rect 2495 1190 2499 1194
rect 727 1146 731 1150
rect 759 1146 763 1150
rect 855 1146 859 1150
rect 879 1146 883 1150
rect 983 1146 987 1150
rect 999 1146 1003 1150
rect 1103 1146 1107 1150
rect 1119 1146 1123 1150
rect 1223 1146 1227 1150
rect 1231 1146 1235 1150
rect 1335 1146 1339 1150
rect 1343 1146 1347 1150
rect 1447 1146 1451 1150
rect 1463 1146 1467 1150
rect 1567 1146 1571 1150
rect 1631 1146 1635 1150
rect 1671 1150 1675 1154
rect 2175 1150 2179 1154
rect 527 1094 531 1098
rect 631 1094 635 1098
rect 423 1046 427 1050
rect 527 1046 531 1050
rect 655 1094 659 1098
rect 759 1094 763 1098
rect 775 1094 779 1098
rect 879 1094 883 1098
rect 895 1094 899 1098
rect 999 1094 1003 1098
rect 1015 1094 1019 1098
rect 1119 1094 1123 1098
rect 1127 1094 1131 1098
rect 1231 1094 1235 1098
rect 1247 1094 1251 1098
rect 2551 1190 2555 1194
rect 2695 1190 2699 1194
rect 2711 1190 2715 1194
rect 2847 1190 2851 1194
rect 2919 1190 2923 1194
rect 2999 1190 3003 1194
rect 3135 1190 3139 1194
rect 2247 1150 2251 1154
rect 2335 1150 2339 1154
rect 2399 1150 2403 1154
rect 2495 1150 2499 1154
rect 2551 1150 2555 1154
rect 2655 1150 2659 1154
rect 2695 1150 2699 1154
rect 2815 1150 2819 1154
rect 2847 1150 2851 1154
rect 2975 1150 2979 1154
rect 2999 1150 3003 1154
rect 3135 1150 3139 1154
rect 3191 1190 3195 1194
rect 3191 1150 3195 1154
rect 1671 1106 1675 1110
rect 2071 1106 2075 1110
rect 2175 1106 2179 1110
rect 1343 1094 1347 1098
rect 1367 1094 1371 1098
rect 1463 1094 1467 1098
rect 1631 1094 1635 1098
rect 2191 1106 2195 1110
rect 2327 1106 2331 1110
rect 2335 1106 2339 1110
rect 2479 1106 2483 1110
rect 2495 1106 2499 1110
rect 2639 1106 2643 1110
rect 2655 1106 2659 1110
rect 2815 1106 2819 1110
rect 2975 1106 2979 1110
rect 2999 1106 3003 1110
rect 3135 1106 3139 1110
rect 3159 1106 3163 1110
rect 3191 1106 3195 1110
rect 551 1046 555 1050
rect 655 1046 659 1050
rect 679 1046 683 1050
rect 775 1046 779 1050
rect 799 1046 803 1050
rect 895 1046 899 1050
rect 919 1046 923 1050
rect 1015 1046 1019 1050
rect 1031 1046 1035 1050
rect 1127 1046 1131 1050
rect 1143 1046 1147 1050
rect 1247 1046 1251 1050
rect 1671 1054 1675 1058
rect 1975 1054 1979 1058
rect 2071 1054 2075 1058
rect 1263 1046 1267 1050
rect 1367 1046 1371 1050
rect 1631 1046 1635 1050
rect 327 994 331 998
rect 423 994 427 998
rect 455 994 459 998
rect 551 994 555 998
rect 575 994 579 998
rect 679 994 683 998
rect 695 994 699 998
rect 799 994 803 998
rect 815 994 819 998
rect 919 994 923 998
rect 927 994 931 998
rect 1031 994 1035 998
rect 1039 994 1043 998
rect 1143 994 1147 998
rect 1159 994 1163 998
rect 327 942 331 946
rect 351 942 355 946
rect 455 942 459 946
rect 471 942 475 946
rect 575 942 579 946
rect 2095 1054 2099 1058
rect 2191 1054 2195 1058
rect 2215 1054 2219 1058
rect 2327 1054 2331 1058
rect 2343 1054 2347 1058
rect 2479 1054 2483 1058
rect 2487 1054 2491 1058
rect 2639 1054 2643 1058
rect 2647 1054 2651 1058
rect 2815 1054 2819 1058
rect 2823 1054 2827 1058
rect 2999 1054 3003 1058
rect 3159 1054 3163 1058
rect 1671 1010 1675 1014
rect 1895 1010 1899 1014
rect 1975 1010 1979 1014
rect 2047 1010 2051 1014
rect 2095 1010 2099 1014
rect 2199 1010 2203 1014
rect 2215 1010 2219 1014
rect 2343 1010 2347 1014
rect 1263 994 1267 998
rect 1631 994 1635 998
rect 1671 970 1675 974
rect 1791 970 1795 974
rect 1895 970 1899 974
rect 1919 970 1923 974
rect 591 942 595 946
rect 695 942 699 946
rect 711 942 715 946
rect 815 942 819 946
rect 823 942 827 946
rect 927 942 931 946
rect 943 942 947 946
rect 1039 942 1043 946
rect 1063 942 1067 946
rect 1159 942 1163 946
rect 111 890 115 894
rect 135 890 139 894
rect 223 890 227 894
rect 247 890 251 894
rect 351 890 355 894
rect 383 890 387 894
rect 471 890 475 894
rect 535 890 539 894
rect 591 890 595 894
rect 711 890 715 894
rect 823 890 827 894
rect 919 890 923 894
rect 943 890 947 894
rect 1063 890 1067 894
rect 111 846 115 850
rect 135 846 139 850
rect 247 846 251 850
rect 303 846 307 850
rect 383 846 387 850
rect 503 846 507 850
rect 535 846 539 850
rect 695 846 699 850
rect 711 846 715 850
rect 111 790 115 794
rect 135 790 139 794
rect 303 790 307 794
rect 503 790 507 794
rect 111 742 115 746
rect 575 742 579 746
rect 879 846 883 850
rect 919 846 923 850
rect 1047 846 1051 850
rect 1143 890 1147 894
rect 1631 942 1635 946
rect 2047 970 2051 974
rect 2071 970 2075 974
rect 2199 970 2203 974
rect 3191 1054 3195 1058
rect 2487 1010 2491 1014
rect 2495 1010 2499 1014
rect 2647 1010 2651 1014
rect 2823 1010 2827 1014
rect 2255 970 2259 974
rect 2343 970 2347 974
rect 2463 970 2467 974
rect 2495 970 2499 974
rect 2647 970 2651 974
rect 2695 970 2699 974
rect 2999 1010 3003 1014
rect 2935 970 2939 974
rect 3159 1010 3163 1014
rect 3159 970 3163 974
rect 3191 1010 3195 1014
rect 3191 970 3195 974
rect 1671 922 1675 926
rect 1719 922 1723 926
rect 1791 922 1795 926
rect 1871 922 1875 926
rect 1919 922 1923 926
rect 2039 922 2043 926
rect 2071 922 2075 926
rect 2223 922 2227 926
rect 2255 922 2259 926
rect 2439 922 2443 926
rect 2463 922 2467 926
rect 2671 922 2675 926
rect 2695 922 2699 926
rect 2911 922 2915 926
rect 2935 922 2939 926
rect 3159 922 3163 926
rect 3191 922 3195 926
rect 1383 890 1387 894
rect 1599 890 1603 894
rect 1631 890 1635 894
rect 1671 882 1675 886
rect 1695 882 1699 886
rect 1719 882 1723 886
rect 1871 882 1875 886
rect 2015 882 2019 886
rect 1143 846 1147 850
rect 1199 846 1203 850
rect 1335 846 1339 850
rect 1383 846 1387 850
rect 2039 882 2043 886
rect 2223 882 2227 886
rect 1471 846 1475 850
rect 1599 846 1603 850
rect 1631 846 1635 850
rect 679 790 683 794
rect 695 790 699 794
rect 807 790 811 794
rect 879 790 883 794
rect 679 742 683 746
rect 703 742 707 746
rect 807 742 811 746
rect 831 742 835 746
rect 927 790 931 794
rect 1047 790 1051 794
rect 1167 790 1171 794
rect 1199 790 1203 794
rect 1279 790 1283 794
rect 1335 790 1339 794
rect 1399 790 1403 794
rect 1471 790 1475 794
rect 1519 790 1523 794
rect 1671 830 1675 834
rect 1695 830 1699 834
rect 2015 830 2019 834
rect 2367 882 2371 886
rect 2439 882 2443 886
rect 2671 882 2675 886
rect 2727 882 2731 886
rect 2911 882 2915 886
rect 3087 882 3091 886
rect 3159 882 3163 886
rect 3191 882 3195 886
rect 2279 830 2283 834
rect 2367 830 2371 834
rect 2439 830 2443 834
rect 2583 830 2587 834
rect 2719 830 2723 834
rect 2727 830 2731 834
rect 2847 830 2851 834
rect 2975 830 2979 834
rect 3087 830 3091 834
rect 3111 830 3115 834
rect 3191 830 3195 834
rect 1599 790 1603 794
rect 1631 790 1635 794
rect 1671 786 1675 790
rect 2199 786 2203 790
rect 2279 786 2283 790
rect 927 742 931 746
rect 951 742 955 746
rect 1047 742 1051 746
rect 1071 742 1075 746
rect 1167 742 1171 746
rect 1183 742 1187 746
rect 1279 742 1283 746
rect 1295 742 1299 746
rect 1399 742 1403 746
rect 1415 742 1419 746
rect 1519 742 1523 746
rect 1631 742 1635 746
rect 1671 742 1675 746
rect 2127 742 2131 746
rect 2199 742 2203 746
rect 2287 742 2291 746
rect 2359 786 2363 790
rect 2439 786 2443 790
rect 2511 786 2515 790
rect 2583 786 2587 790
rect 2655 786 2659 790
rect 2719 786 2723 790
rect 2791 786 2795 790
rect 2359 742 2363 746
rect 2447 742 2451 746
rect 2847 786 2851 790
rect 2919 786 2923 790
rect 2975 786 2979 790
rect 3047 786 3051 790
rect 3111 786 3115 790
rect 3159 786 3163 790
rect 3191 786 3195 790
rect 2511 742 2515 746
rect 2599 742 2603 746
rect 2655 742 2659 746
rect 2759 742 2763 746
rect 2791 742 2795 746
rect 2919 742 2923 746
rect 3047 742 3051 746
rect 3159 742 3163 746
rect 111 690 115 694
rect 479 690 483 694
rect 575 690 579 694
rect 607 690 611 694
rect 703 690 707 694
rect 727 690 731 694
rect 831 690 835 694
rect 847 690 851 694
rect 951 690 955 694
rect 967 690 971 694
rect 1071 690 1075 694
rect 1079 690 1083 694
rect 1183 690 1187 694
rect 1191 690 1195 694
rect 1295 690 1299 694
rect 1311 690 1315 694
rect 1671 702 1675 706
rect 2023 702 2027 706
rect 2127 702 2131 706
rect 2151 702 2155 706
rect 1415 690 1419 694
rect 1631 690 1635 694
rect 2287 702 2291 706
rect 2295 702 2299 706
rect 2447 702 2451 706
rect 2599 702 2603 706
rect 2615 702 2619 706
rect 2759 702 2763 706
rect 111 638 115 642
rect 375 638 379 642
rect 479 638 483 642
rect 503 638 507 642
rect 607 638 611 642
rect 623 638 627 642
rect 727 638 731 642
rect 743 638 747 642
rect 847 638 851 642
rect 863 638 867 642
rect 967 638 971 642
rect 975 638 979 642
rect 1079 638 1083 642
rect 1095 638 1099 642
rect 1191 638 1195 642
rect 1215 638 1219 642
rect 1671 654 1675 658
rect 1919 654 1923 658
rect 2023 654 2027 658
rect 2047 654 2051 658
rect 2151 654 2155 658
rect 2183 654 2187 658
rect 2295 654 2299 658
rect 2327 654 2331 658
rect 2447 654 2451 658
rect 2471 654 2475 658
rect 2615 654 2619 658
rect 2759 654 2763 658
rect 2799 702 2803 706
rect 2919 702 2923 706
rect 2991 702 2995 706
rect 3159 702 3163 706
rect 3191 742 3195 746
rect 3191 702 3195 706
rect 2799 654 2803 658
rect 1311 638 1315 642
rect 1631 638 1635 642
rect 111 590 115 594
rect 271 590 275 594
rect 375 590 379 594
rect 399 590 403 594
rect 503 590 507 594
rect 527 590 531 594
rect 623 590 627 594
rect 647 590 651 594
rect 743 590 747 594
rect 767 590 771 594
rect 863 590 867 594
rect 879 590 883 594
rect 975 590 979 594
rect 991 590 995 594
rect 111 538 115 542
rect 175 538 179 542
rect 271 538 275 542
rect 303 538 307 542
rect 399 538 403 542
rect 423 538 427 542
rect 527 538 531 542
rect 543 538 547 542
rect 647 538 651 542
rect 663 538 667 542
rect 767 538 771 542
rect 775 538 779 542
rect 1671 610 1675 614
rect 1847 610 1851 614
rect 1095 590 1099 594
rect 1111 590 1115 594
rect 1215 590 1219 594
rect 1631 590 1635 594
rect 1671 570 1675 574
rect 1767 570 1771 574
rect 1847 570 1851 574
rect 1919 610 1923 614
rect 2015 610 2019 614
rect 1927 570 1931 574
rect 2015 570 2019 574
rect 2047 610 2051 614
rect 2183 610 2187 614
rect 2327 610 2331 614
rect 2359 610 2363 614
rect 2087 570 2091 574
rect 2183 570 2187 574
rect 2247 570 2251 574
rect 2359 570 2363 574
rect 2407 570 2411 574
rect 2471 610 2475 614
rect 2551 610 2555 614
rect 2615 610 2619 614
rect 2751 610 2755 614
rect 2759 610 2763 614
rect 2551 570 2555 574
rect 2567 570 2571 574
rect 2751 570 2755 574
rect 879 538 883 542
rect 887 538 891 542
rect 991 538 995 542
rect 1007 538 1011 542
rect 1111 538 1115 542
rect 111 486 115 490
rect 135 486 139 490
rect 175 486 179 490
rect 231 486 235 490
rect 303 486 307 490
rect 359 486 363 490
rect 423 486 427 490
rect 503 486 507 490
rect 543 486 547 490
rect 655 486 659 490
rect 663 486 667 490
rect 775 486 779 490
rect 815 486 819 490
rect 111 434 115 438
rect 135 434 139 438
rect 231 434 235 438
rect 359 434 363 438
rect 111 386 115 390
rect 111 342 115 346
rect 111 298 115 302
rect 463 298 467 302
rect 887 486 891 490
rect 975 486 979 490
rect 1007 486 1011 490
rect 1135 486 1139 490
rect 1631 538 1635 542
rect 1671 530 1675 534
rect 1695 530 1699 534
rect 1767 530 1771 534
rect 1887 530 1891 534
rect 1927 530 1931 534
rect 1295 486 1299 490
rect 1455 486 1459 490
rect 1599 486 1603 490
rect 1631 486 1635 490
rect 1671 482 1675 486
rect 1695 482 1699 486
rect 1887 482 1891 486
rect 2023 482 2027 486
rect 2087 530 2091 534
rect 2103 530 2107 534
rect 2247 530 2251 534
rect 2343 530 2347 534
rect 2407 530 2411 534
rect 2567 530 2571 534
rect 2599 530 2603 534
rect 2863 530 2867 534
rect 2991 654 2995 658
rect 3159 654 3163 658
rect 2959 610 2963 614
rect 3159 610 3163 614
rect 3191 654 3195 658
rect 3191 610 3195 614
rect 2959 570 2963 574
rect 3159 570 3163 574
rect 3135 530 3139 534
rect 3191 570 3195 574
rect 3191 530 3195 534
rect 2103 482 2107 486
rect 2343 482 2347 486
rect 2383 482 2387 486
rect 2599 482 2603 486
rect 503 434 507 438
rect 655 434 659 438
rect 727 434 731 438
rect 815 434 819 438
rect 855 434 859 438
rect 975 434 979 438
rect 983 434 987 438
rect 1103 434 1107 438
rect 1135 434 1139 438
rect 1223 434 1227 438
rect 1295 434 1299 438
rect 1335 434 1339 438
rect 647 386 651 390
rect 1447 434 1451 438
rect 1455 434 1459 438
rect 1567 434 1571 438
rect 1599 434 1603 438
rect 1631 434 1635 438
rect 1671 438 1675 442
rect 1695 438 1699 442
rect 2023 438 2027 442
rect 727 386 731 390
rect 807 386 811 390
rect 855 386 859 390
rect 951 386 955 390
rect 983 386 987 390
rect 1087 386 1091 390
rect 1103 386 1107 390
rect 1215 386 1219 390
rect 1223 386 1227 390
rect 1335 386 1339 390
rect 1447 386 1451 390
rect 1463 386 1467 390
rect 1567 386 1571 390
rect 1631 386 1635 390
rect 1671 386 1675 390
rect 543 342 547 346
rect 647 342 651 346
rect 671 342 675 346
rect 807 342 811 346
rect 943 342 947 346
rect 951 342 955 346
rect 1079 342 1083 346
rect 1087 342 1091 346
rect 1215 342 1219 346
rect 1223 342 1227 346
rect 1335 342 1339 346
rect 1367 342 1371 346
rect 1463 342 1467 346
rect 1631 342 1635 346
rect 543 298 547 302
rect 623 298 627 302
rect 671 298 675 302
rect 767 298 771 302
rect 807 298 811 302
rect 903 298 907 302
rect 943 298 947 302
rect 1031 298 1035 302
rect 1079 298 1083 302
rect 1159 298 1163 302
rect 1223 298 1227 302
rect 1287 298 1291 302
rect 1671 334 1675 338
rect 2047 334 2051 338
rect 2247 438 2251 442
rect 2375 438 2379 442
rect 2383 438 2387 442
rect 2503 438 2507 442
rect 2623 438 2627 442
rect 2743 482 2747 486
rect 2863 482 2867 486
rect 2743 438 2747 442
rect 2855 438 2859 442
rect 3111 482 3115 486
rect 3135 482 3139 486
rect 3191 482 3195 486
rect 2967 438 2971 442
rect 3087 438 3091 442
rect 3111 438 3115 442
rect 3191 438 3195 442
rect 2151 386 2155 390
rect 2247 386 2251 390
rect 2279 386 2283 390
rect 2375 386 2379 390
rect 2407 386 2411 390
rect 2503 386 2507 390
rect 2535 386 2539 390
rect 2623 386 2627 390
rect 2663 386 2667 390
rect 2743 386 2747 390
rect 2791 386 2795 390
rect 2855 386 2859 390
rect 2919 386 2923 390
rect 2967 386 2971 390
rect 3047 386 3051 390
rect 3087 386 3091 390
rect 3159 386 3163 390
rect 3191 386 3195 390
rect 2151 334 2155 338
rect 2175 334 2179 338
rect 2279 334 2283 338
rect 2303 334 2307 338
rect 2407 334 2411 338
rect 2431 334 2435 338
rect 2535 334 2539 338
rect 2567 334 2571 338
rect 1367 298 1371 302
rect 1631 298 1635 302
rect 2663 334 2667 338
rect 2711 334 2715 338
rect 2791 334 2795 338
rect 2863 334 2867 338
rect 2919 334 2923 338
rect 3023 334 3027 338
rect 3047 334 3051 338
rect 3159 334 3163 338
rect 3191 334 3195 338
rect 1671 286 1675 290
rect 1943 286 1947 290
rect 2047 286 2051 290
rect 2071 286 2075 290
rect 2175 286 2179 290
rect 2199 286 2203 290
rect 2303 286 2307 290
rect 2319 286 2323 290
rect 2431 286 2435 290
rect 2439 286 2443 290
rect 2551 286 2555 290
rect 2567 286 2571 290
rect 2663 286 2667 290
rect 2711 286 2715 290
rect 2783 286 2787 290
rect 2863 286 2867 290
rect 111 254 115 258
rect 359 254 363 258
rect 463 254 467 258
rect 487 254 491 258
rect 623 254 627 258
rect 759 254 763 258
rect 767 254 771 258
rect 111 210 115 214
rect 279 210 283 214
rect 359 210 363 214
rect 447 210 451 214
rect 895 254 899 258
rect 903 254 907 258
rect 1031 254 1035 258
rect 1039 254 1043 258
rect 1159 254 1163 258
rect 1183 254 1187 258
rect 1287 254 1291 258
rect 1631 254 1635 258
rect 487 210 491 214
rect 615 210 619 214
rect 623 210 627 214
rect 111 170 115 174
rect 199 170 203 174
rect 279 170 283 174
rect 367 170 371 174
rect 447 170 451 174
rect 759 210 763 214
rect 535 170 539 174
rect 615 170 619 174
rect 695 170 699 174
rect 775 210 779 214
rect 895 210 899 214
rect 1671 234 1675 238
rect 1847 234 1851 238
rect 1943 234 1947 238
rect 1975 234 1979 238
rect 2071 234 2075 238
rect 2103 234 2107 238
rect 2199 234 2203 238
rect 2247 234 2251 238
rect 2319 234 2323 238
rect 2407 234 2411 238
rect 2439 234 2443 238
rect 943 210 947 214
rect 1039 210 1043 214
rect 1111 210 1115 214
rect 1183 210 1187 214
rect 1631 210 1635 214
rect 775 170 779 174
rect 863 170 867 174
rect 1671 182 1675 186
rect 1743 182 1747 186
rect 1847 182 1851 186
rect 943 170 947 174
rect 1031 170 1035 174
rect 1111 170 1115 174
rect 1631 170 1635 174
rect 1871 182 1875 186
rect 1975 182 1979 186
rect 1999 182 2003 186
rect 2103 182 2107 186
rect 2143 182 2147 186
rect 2247 182 2251 186
rect 2311 182 2315 186
rect 2407 182 2411 186
rect 2495 182 2499 186
rect 111 118 115 122
rect 135 118 139 122
rect 191 118 195 122
rect 199 118 203 122
rect 287 118 291 122
rect 367 118 371 122
rect 383 118 387 122
rect 479 118 483 122
rect 535 118 539 122
rect 583 118 587 122
rect 695 118 699 122
rect 815 118 819 122
rect 863 118 867 122
rect 943 118 947 122
rect 1671 126 1675 130
rect 1695 126 1699 130
rect 1743 126 1747 130
rect 1031 118 1035 122
rect 1079 118 1083 122
rect 1215 118 1219 122
rect 1351 118 1355 122
rect 1487 118 1491 122
rect 1599 118 1603 122
rect 1631 118 1635 122
rect 1671 86 1675 90
rect 1695 86 1699 90
rect 1815 126 1819 130
rect 1871 126 1875 130
rect 1943 126 1947 130
rect 1999 126 2003 130
rect 2071 126 2075 130
rect 2143 126 2147 130
rect 2199 126 2203 130
rect 2311 126 2315 130
rect 2351 126 2355 130
rect 2495 126 2499 130
rect 2519 126 2523 130
rect 2551 234 2555 238
rect 2583 234 2587 238
rect 2663 234 2667 238
rect 2583 182 2587 186
rect 2703 182 2707 186
rect 2767 234 2771 238
rect 2783 234 2787 238
rect 3023 286 3027 290
rect 3159 286 3163 290
rect 2967 234 2971 238
rect 3159 234 3163 238
rect 3191 286 3195 290
rect 3191 234 3195 238
rect 2767 182 2771 186
rect 2919 182 2923 186
rect 2967 182 2971 186
rect 3135 182 3139 186
rect 3159 182 3163 186
rect 3191 182 3195 186
rect 2703 126 2707 130
rect 2711 126 2715 130
rect 2911 126 2915 130
rect 2919 126 2923 130
rect 3111 126 3115 130
rect 3135 126 3139 130
rect 3191 126 3195 130
rect 1815 86 1819 90
rect 1943 86 1947 90
rect 2071 86 2075 90
rect 2199 86 2203 90
rect 2351 86 2355 90
rect 2519 86 2523 90
rect 2711 86 2715 90
rect 2911 86 2915 90
rect 3111 86 3115 90
rect 3191 86 3195 90
rect 111 78 115 82
rect 135 78 139 82
rect 191 78 195 82
rect 287 78 291 82
rect 383 78 387 82
rect 479 78 483 82
rect 583 78 587 82
rect 695 78 699 82
rect 815 78 819 82
rect 943 78 947 82
rect 1079 78 1083 82
rect 1215 78 1219 82
rect 1351 78 1355 82
rect 1487 78 1491 82
rect 1599 78 1603 82
rect 1631 78 1635 82
<< m4 >>
rect 1654 3305 1655 3311
rect 1661 3310 3231 3311
rect 1661 3306 1671 3310
rect 1675 3306 3055 3310
rect 3059 3306 3191 3310
rect 3195 3306 3231 3310
rect 1661 3305 3231 3306
rect 3237 3305 3238 3311
rect 1642 3265 1643 3271
rect 1649 3270 3219 3271
rect 1649 3266 1671 3270
rect 1675 3266 2151 3270
rect 2155 3266 2287 3270
rect 2291 3266 2423 3270
rect 2427 3266 2567 3270
rect 2571 3266 2711 3270
rect 2715 3266 2855 3270
rect 2859 3266 2999 3270
rect 3003 3266 3055 3270
rect 3059 3266 3191 3270
rect 3195 3266 3219 3270
rect 1649 3265 3219 3266
rect 3225 3265 3226 3271
rect 1654 3225 1655 3231
rect 1661 3230 3231 3231
rect 1661 3226 1671 3230
rect 1675 3226 1999 3230
rect 2003 3226 2151 3230
rect 2155 3226 2175 3230
rect 2179 3226 2287 3230
rect 2291 3226 2359 3230
rect 2363 3226 2423 3230
rect 2427 3226 2543 3230
rect 2547 3226 2567 3230
rect 2571 3226 2711 3230
rect 2715 3226 2727 3230
rect 2731 3226 2855 3230
rect 2859 3226 2919 3230
rect 2923 3226 2999 3230
rect 3003 3226 3111 3230
rect 3115 3226 3191 3230
rect 3195 3226 3231 3230
rect 1661 3225 3231 3226
rect 3237 3225 3238 3231
rect 1642 3185 1643 3191
rect 1649 3190 3219 3191
rect 1649 3186 1671 3190
rect 1675 3186 1847 3190
rect 1851 3186 1999 3190
rect 2003 3186 2039 3190
rect 2043 3186 2175 3190
rect 2179 3186 2247 3190
rect 2251 3186 2359 3190
rect 2363 3186 2463 3190
rect 2467 3186 2543 3190
rect 2547 3186 2695 3190
rect 2699 3186 2727 3190
rect 2731 3186 2919 3190
rect 2923 3186 2935 3190
rect 2939 3186 3111 3190
rect 3115 3186 3159 3190
rect 3163 3186 3191 3190
rect 3195 3186 3219 3190
rect 1649 3185 3219 3186
rect 3225 3185 3226 3191
rect 1654 3145 1655 3151
rect 1661 3150 3231 3151
rect 1661 3146 1671 3150
rect 1675 3146 1695 3150
rect 1699 3146 1847 3150
rect 1851 3146 1863 3150
rect 1867 3146 2023 3150
rect 2027 3146 2039 3150
rect 2043 3146 2183 3150
rect 2187 3146 2247 3150
rect 2251 3146 2343 3150
rect 2347 3146 2463 3150
rect 2467 3146 2511 3150
rect 2515 3146 2695 3150
rect 2699 3146 2935 3150
rect 2939 3146 3159 3150
rect 3163 3146 3191 3150
rect 3195 3146 3231 3150
rect 1661 3145 3231 3146
rect 3237 3145 3238 3151
rect 84 3125 85 3131
rect 91 3130 1643 3131
rect 91 3126 111 3130
rect 115 3126 807 3130
rect 811 3126 1079 3130
rect 1083 3126 1351 3130
rect 1355 3126 1599 3130
rect 1603 3126 1631 3130
rect 1635 3126 1643 3130
rect 91 3125 1643 3126
rect 1649 3125 1650 3131
rect 1642 3105 1643 3111
rect 1649 3110 3219 3111
rect 1649 3106 1671 3110
rect 1675 3106 1695 3110
rect 1699 3106 1863 3110
rect 1867 3106 1959 3110
rect 1963 3106 2023 3110
rect 2027 3106 2183 3110
rect 2187 3106 2343 3110
rect 2347 3106 2415 3110
rect 2419 3106 2511 3110
rect 2515 3106 2655 3110
rect 2659 3106 2903 3110
rect 2907 3106 3159 3110
rect 3163 3106 3191 3110
rect 3195 3106 3219 3110
rect 1649 3105 3219 3106
rect 3225 3105 3226 3111
rect 96 3081 97 3087
rect 103 3086 1655 3087
rect 103 3082 111 3086
rect 115 3082 703 3086
rect 707 3082 807 3086
rect 811 3082 831 3086
rect 835 3082 959 3086
rect 963 3082 1079 3086
rect 1083 3082 1199 3086
rect 1203 3082 1311 3086
rect 1315 3082 1351 3086
rect 1355 3082 1423 3086
rect 1427 3082 1543 3086
rect 1547 3082 1599 3086
rect 1603 3082 1631 3086
rect 1635 3082 1655 3086
rect 103 3081 1655 3082
rect 1661 3081 1662 3087
rect 1654 3065 1655 3071
rect 1661 3070 3231 3071
rect 1661 3066 1671 3070
rect 1675 3066 1871 3070
rect 1875 3066 1959 3070
rect 1963 3066 2111 3070
rect 2115 3066 2183 3070
rect 2187 3066 2367 3070
rect 2371 3066 2415 3070
rect 2419 3066 2631 3070
rect 2635 3066 2655 3070
rect 2659 3066 2903 3070
rect 2907 3066 3159 3070
rect 3163 3066 3191 3070
rect 3195 3066 3231 3070
rect 1661 3065 3231 3066
rect 3237 3065 3238 3071
rect 84 3033 85 3039
rect 91 3038 1643 3039
rect 91 3034 111 3038
rect 115 3034 623 3038
rect 627 3034 703 3038
rect 707 3034 783 3038
rect 787 3034 831 3038
rect 835 3034 927 3038
rect 931 3034 959 3038
rect 963 3034 1063 3038
rect 1067 3034 1079 3038
rect 1083 3034 1191 3038
rect 1195 3034 1199 3038
rect 1203 3034 1311 3038
rect 1315 3034 1423 3038
rect 1427 3034 1439 3038
rect 1443 3034 1543 3038
rect 1547 3034 1631 3038
rect 1635 3034 1643 3038
rect 91 3033 1643 3034
rect 1649 3033 1650 3039
rect 1642 3031 1650 3033
rect 1642 3025 1643 3031
rect 1649 3030 3219 3031
rect 1649 3026 1671 3030
rect 1675 3026 1791 3030
rect 1795 3026 1871 3030
rect 1875 3026 1959 3030
rect 1963 3026 2111 3030
rect 2115 3026 2127 3030
rect 2131 3026 2287 3030
rect 2291 3026 2367 3030
rect 2371 3026 2455 3030
rect 2459 3026 2623 3030
rect 2627 3026 2631 3030
rect 2635 3026 2903 3030
rect 2907 3026 3159 3030
rect 3163 3026 3191 3030
rect 3195 3026 3219 3030
rect 1649 3025 3219 3026
rect 3225 3025 3226 3031
rect 96 2989 97 2995
rect 103 2994 1655 2995
rect 103 2990 111 2994
rect 115 2990 519 2994
rect 523 2990 623 2994
rect 627 2990 647 2994
rect 651 2990 783 2994
rect 787 2990 919 2994
rect 923 2990 927 2994
rect 931 2990 1055 2994
rect 1059 2990 1063 2994
rect 1067 2990 1191 2994
rect 1195 2990 1311 2994
rect 1315 2990 1335 2994
rect 1339 2990 1439 2994
rect 1443 2990 1631 2994
rect 1635 2990 1655 2994
rect 103 2989 1655 2990
rect 1661 2991 1662 2995
rect 1661 2990 3238 2991
rect 1661 2989 1671 2990
rect 1654 2986 1671 2989
rect 1675 2986 1703 2990
rect 1707 2986 1791 2990
rect 1795 2986 1903 2990
rect 1907 2986 1959 2990
rect 1963 2986 2127 2990
rect 2131 2986 2287 2990
rect 2291 2986 2367 2990
rect 2371 2986 2455 2990
rect 2459 2986 2623 2990
rect 2627 2986 2887 2990
rect 2891 2986 3159 2990
rect 3163 2986 3191 2990
rect 3195 2986 3238 2990
rect 1654 2985 3238 2986
rect 1642 2950 3226 2951
rect 1642 2947 1671 2950
rect 84 2941 85 2947
rect 91 2946 1643 2947
rect 91 2942 111 2946
rect 115 2942 439 2946
rect 443 2942 519 2946
rect 523 2942 599 2946
rect 603 2942 647 2946
rect 651 2942 759 2946
rect 763 2942 783 2946
rect 787 2942 919 2946
rect 923 2942 927 2946
rect 931 2942 1055 2946
rect 1059 2942 1095 2946
rect 1099 2942 1191 2946
rect 1195 2942 1263 2946
rect 1267 2942 1335 2946
rect 1339 2942 1439 2946
rect 1443 2942 1599 2946
rect 1603 2942 1631 2946
rect 1635 2942 1643 2946
rect 91 2941 1643 2942
rect 1649 2946 1671 2947
rect 1675 2946 1695 2950
rect 1699 2946 1703 2950
rect 1707 2946 1903 2950
rect 1907 2946 1935 2950
rect 1939 2946 2127 2950
rect 2131 2946 2223 2950
rect 2227 2946 2367 2950
rect 2371 2946 2519 2950
rect 2523 2946 2623 2950
rect 2627 2946 2823 2950
rect 2827 2946 2887 2950
rect 2891 2946 3135 2950
rect 3139 2946 3159 2950
rect 3163 2946 3191 2950
rect 3195 2946 3226 2950
rect 1649 2945 3226 2946
rect 1649 2941 1650 2945
rect 1654 2910 3238 2911
rect 1654 2907 1671 2910
rect 96 2901 97 2907
rect 103 2906 1655 2907
rect 103 2902 111 2906
rect 115 2902 335 2906
rect 339 2902 439 2906
rect 443 2902 471 2906
rect 475 2902 599 2906
rect 603 2902 623 2906
rect 627 2902 759 2906
rect 763 2902 791 2906
rect 795 2902 927 2906
rect 931 2902 975 2906
rect 979 2902 1095 2906
rect 1099 2902 1175 2906
rect 1179 2902 1263 2906
rect 1267 2902 1383 2906
rect 1387 2902 1439 2906
rect 1443 2902 1591 2906
rect 1595 2902 1599 2906
rect 1603 2902 1631 2906
rect 1635 2902 1655 2906
rect 103 2901 1655 2902
rect 1661 2906 1671 2907
rect 1675 2906 1695 2910
rect 1699 2906 1935 2910
rect 1939 2906 2223 2910
rect 2227 2906 2295 2910
rect 2299 2906 2519 2910
rect 2523 2906 2551 2910
rect 2555 2906 2815 2910
rect 2819 2906 2823 2910
rect 2827 2906 3079 2910
rect 3083 2906 3135 2910
rect 3139 2906 3191 2910
rect 3195 2906 3238 2910
rect 1661 2905 3238 2906
rect 1661 2901 1662 2905
rect 1642 2865 1643 2871
rect 1649 2870 3219 2871
rect 1649 2866 1671 2870
rect 1675 2866 2207 2870
rect 2211 2866 2295 2870
rect 2299 2866 2375 2870
rect 2379 2866 2535 2870
rect 2539 2866 2551 2870
rect 2555 2866 2679 2870
rect 2683 2866 2815 2870
rect 2819 2866 2823 2870
rect 2827 2866 2967 2870
rect 2971 2866 3079 2870
rect 3083 2866 3111 2870
rect 3115 2866 3191 2870
rect 3195 2866 3219 2870
rect 1649 2865 3219 2866
rect 3225 2865 3226 2871
rect 84 2853 85 2859
rect 91 2858 1643 2859
rect 91 2854 111 2858
rect 115 2854 255 2858
rect 259 2854 335 2858
rect 339 2854 415 2858
rect 419 2854 471 2858
rect 475 2854 559 2858
rect 563 2854 623 2858
rect 627 2854 695 2858
rect 699 2854 791 2858
rect 795 2854 823 2858
rect 827 2854 951 2858
rect 955 2854 975 2858
rect 979 2854 1087 2858
rect 1091 2854 1175 2858
rect 1179 2854 1383 2858
rect 1387 2854 1591 2858
rect 1595 2854 1631 2858
rect 1635 2854 1643 2858
rect 91 2853 1643 2854
rect 1649 2853 1650 2859
rect 1654 2817 1655 2823
rect 1661 2822 3231 2823
rect 1661 2818 1671 2822
rect 1675 2818 2127 2822
rect 2131 2818 2207 2822
rect 2211 2818 2303 2822
rect 2307 2818 2375 2822
rect 2379 2818 2479 2822
rect 2483 2818 2535 2822
rect 2539 2818 2655 2822
rect 2659 2818 2679 2822
rect 2683 2818 2823 2822
rect 2827 2818 2831 2822
rect 2835 2818 2967 2822
rect 2971 2818 3007 2822
rect 3011 2818 3111 2822
rect 3115 2818 3159 2822
rect 3163 2818 3191 2822
rect 3195 2818 3231 2822
rect 1661 2817 3231 2818
rect 3237 2817 3238 2823
rect 96 2805 97 2811
rect 103 2810 1655 2811
rect 103 2806 111 2810
rect 115 2806 151 2810
rect 155 2806 255 2810
rect 259 2806 279 2810
rect 283 2806 399 2810
rect 403 2806 415 2810
rect 419 2806 519 2810
rect 523 2806 559 2810
rect 563 2806 639 2810
rect 643 2806 695 2810
rect 699 2806 751 2810
rect 755 2806 823 2810
rect 827 2806 863 2810
rect 867 2806 951 2810
rect 955 2806 983 2810
rect 987 2806 1087 2810
rect 1091 2806 1631 2810
rect 1635 2806 1655 2810
rect 103 2805 1655 2806
rect 1661 2805 1662 2811
rect 1642 2777 1643 2783
rect 1649 2782 3219 2783
rect 1649 2778 1671 2782
rect 1675 2778 2039 2782
rect 2043 2778 2127 2782
rect 2131 2778 2207 2782
rect 2211 2778 2303 2782
rect 2307 2778 2375 2782
rect 2379 2778 2479 2782
rect 2483 2778 2535 2782
rect 2539 2778 2655 2782
rect 2659 2778 2703 2782
rect 2707 2778 2831 2782
rect 2835 2778 2871 2782
rect 2875 2778 3007 2782
rect 3011 2778 3159 2782
rect 3163 2778 3191 2782
rect 3195 2778 3219 2782
rect 1649 2777 3219 2778
rect 3225 2777 3226 2783
rect 84 2753 85 2759
rect 91 2758 1643 2759
rect 91 2754 111 2758
rect 115 2754 135 2758
rect 139 2754 151 2758
rect 155 2754 263 2758
rect 267 2754 279 2758
rect 283 2754 399 2758
rect 403 2754 431 2758
rect 435 2754 519 2758
rect 523 2754 623 2758
rect 627 2754 639 2758
rect 643 2754 751 2758
rect 755 2754 839 2758
rect 843 2754 863 2758
rect 867 2754 983 2758
rect 987 2754 1071 2758
rect 1075 2754 1319 2758
rect 1323 2754 1567 2758
rect 1571 2754 1631 2758
rect 1635 2754 1643 2758
rect 91 2753 1643 2754
rect 1649 2753 1650 2759
rect 1654 2733 1655 2739
rect 1661 2738 3231 2739
rect 1661 2734 1671 2738
rect 1675 2734 2015 2738
rect 2019 2734 2039 2738
rect 2043 2734 2199 2738
rect 2203 2734 2207 2738
rect 2211 2734 2375 2738
rect 2379 2734 2383 2738
rect 2387 2734 2535 2738
rect 2539 2734 2575 2738
rect 2579 2734 2703 2738
rect 2707 2734 2775 2738
rect 2779 2734 2871 2738
rect 2875 2734 2975 2738
rect 2979 2734 3159 2738
rect 3163 2734 3191 2738
rect 3195 2734 3231 2738
rect 1661 2733 3231 2734
rect 3237 2733 3238 2739
rect 96 2701 97 2707
rect 103 2706 1655 2707
rect 103 2702 111 2706
rect 115 2702 135 2706
rect 139 2702 263 2706
rect 267 2702 431 2706
rect 435 2702 623 2706
rect 627 2702 703 2706
rect 707 2702 831 2706
rect 835 2702 839 2706
rect 843 2702 959 2706
rect 963 2702 1071 2706
rect 1075 2702 1079 2706
rect 1083 2702 1199 2706
rect 1203 2702 1311 2706
rect 1315 2702 1319 2706
rect 1323 2702 1423 2706
rect 1427 2702 1543 2706
rect 1547 2702 1567 2706
rect 1571 2702 1631 2706
rect 1635 2702 1655 2706
rect 103 2701 1655 2702
rect 1661 2701 1662 2707
rect 1642 2685 1643 2691
rect 1649 2690 3219 2691
rect 1649 2686 1671 2690
rect 1675 2686 1999 2690
rect 2003 2686 2015 2690
rect 2019 2686 2175 2690
rect 2179 2686 2199 2690
rect 2203 2686 2359 2690
rect 2363 2686 2383 2690
rect 2387 2686 2551 2690
rect 2555 2686 2575 2690
rect 2579 2686 2759 2690
rect 2763 2686 2775 2690
rect 2779 2686 2967 2690
rect 2971 2686 2975 2690
rect 2979 2686 3159 2690
rect 3163 2686 3191 2690
rect 3195 2686 3219 2690
rect 1649 2685 3219 2686
rect 3225 2685 3226 2691
rect 84 2653 85 2659
rect 91 2658 1643 2659
rect 91 2654 111 2658
rect 115 2654 607 2658
rect 611 2654 703 2658
rect 707 2654 735 2658
rect 739 2654 831 2658
rect 835 2654 855 2658
rect 859 2654 959 2658
rect 963 2654 975 2658
rect 979 2654 1079 2658
rect 1083 2654 1095 2658
rect 1099 2654 1199 2658
rect 1203 2654 1207 2658
rect 1211 2654 1311 2658
rect 1315 2654 1319 2658
rect 1323 2654 1423 2658
rect 1427 2654 1439 2658
rect 1443 2654 1543 2658
rect 1547 2654 1631 2658
rect 1635 2654 1643 2658
rect 91 2653 1643 2654
rect 1649 2653 1650 2659
rect 1654 2645 1655 2651
rect 1661 2650 3231 2651
rect 1661 2646 1671 2650
rect 1675 2646 1911 2650
rect 1915 2646 1999 2650
rect 2003 2646 2103 2650
rect 2107 2646 2175 2650
rect 2179 2646 2295 2650
rect 2299 2646 2359 2650
rect 2363 2646 2487 2650
rect 2491 2646 2551 2650
rect 2555 2646 2687 2650
rect 2691 2646 2759 2650
rect 2763 2646 2967 2650
rect 2971 2646 3159 2650
rect 3163 2646 3191 2650
rect 3195 2646 3231 2650
rect 1661 2645 3231 2646
rect 3237 2645 3238 2651
rect 1642 2611 1643 2617
rect 1649 2611 1674 2617
rect 1668 2610 3219 2611
rect 96 2601 97 2607
rect 103 2606 1655 2607
rect 103 2602 111 2606
rect 115 2602 503 2606
rect 507 2602 607 2606
rect 611 2602 631 2606
rect 635 2602 735 2606
rect 739 2602 751 2606
rect 755 2602 855 2606
rect 859 2602 871 2606
rect 875 2602 975 2606
rect 979 2602 991 2606
rect 995 2602 1095 2606
rect 1099 2602 1103 2606
rect 1107 2602 1207 2606
rect 1211 2602 1215 2606
rect 1219 2602 1319 2606
rect 1323 2602 1335 2606
rect 1339 2602 1439 2606
rect 1443 2602 1631 2606
rect 1635 2602 1655 2606
rect 103 2601 1655 2602
rect 1661 2601 1662 2607
rect 1668 2606 1671 2610
rect 1675 2606 1823 2610
rect 1827 2606 1911 2610
rect 1915 2606 2015 2610
rect 2019 2606 2103 2610
rect 2107 2606 2215 2610
rect 2219 2606 2295 2610
rect 2299 2606 2439 2610
rect 2443 2606 2487 2610
rect 2491 2606 2671 2610
rect 2675 2606 2687 2610
rect 2691 2606 2919 2610
rect 2923 2606 3159 2610
rect 3163 2606 3191 2610
rect 3195 2606 3219 2610
rect 1668 2605 3219 2606
rect 3225 2605 3226 2611
rect 1654 2561 1655 2567
rect 1661 2566 3231 2567
rect 1661 2562 1671 2566
rect 1675 2562 1735 2566
rect 1739 2562 1823 2566
rect 1827 2562 1895 2566
rect 1899 2562 2015 2566
rect 2019 2562 2055 2566
rect 2059 2562 2215 2566
rect 2219 2562 2375 2566
rect 2379 2562 2439 2566
rect 2443 2562 2535 2566
rect 2539 2562 2671 2566
rect 2675 2562 2919 2566
rect 2923 2562 3159 2566
rect 3163 2562 3191 2566
rect 3195 2562 3231 2566
rect 1661 2561 3231 2562
rect 3237 2561 3238 2567
rect 84 2549 85 2555
rect 91 2554 1643 2555
rect 91 2550 111 2554
rect 115 2550 399 2554
rect 403 2550 503 2554
rect 507 2550 527 2554
rect 531 2550 631 2554
rect 635 2550 655 2554
rect 659 2550 751 2554
rect 755 2550 775 2554
rect 779 2550 871 2554
rect 875 2550 895 2554
rect 899 2550 991 2554
rect 995 2550 1007 2554
rect 1011 2550 1103 2554
rect 1107 2550 1119 2554
rect 1123 2550 1215 2554
rect 1219 2550 1239 2554
rect 1243 2550 1335 2554
rect 1339 2550 1631 2554
rect 1635 2550 1643 2554
rect 91 2549 1643 2550
rect 1649 2549 1650 2555
rect 1642 2517 1643 2523
rect 1649 2522 3219 2523
rect 1649 2518 1671 2522
rect 1675 2518 1695 2522
rect 1699 2518 1735 2522
rect 1739 2518 1863 2522
rect 1867 2518 1895 2522
rect 1899 2518 2055 2522
rect 2059 2518 2079 2522
rect 2083 2518 2215 2522
rect 2219 2518 2319 2522
rect 2323 2518 2375 2522
rect 2379 2518 2535 2522
rect 2539 2518 2583 2522
rect 2587 2518 2855 2522
rect 2859 2518 3135 2522
rect 3139 2518 3191 2522
rect 3195 2518 3219 2522
rect 1649 2517 3219 2518
rect 3225 2517 3226 2523
rect 96 2497 97 2503
rect 103 2502 1655 2503
rect 103 2498 111 2502
rect 115 2498 303 2502
rect 307 2498 399 2502
rect 403 2498 431 2502
rect 435 2498 527 2502
rect 531 2498 559 2502
rect 563 2498 655 2502
rect 659 2498 703 2502
rect 707 2498 775 2502
rect 779 2498 863 2502
rect 867 2498 895 2502
rect 899 2498 1007 2502
rect 1011 2498 1039 2502
rect 1043 2498 1119 2502
rect 1123 2498 1223 2502
rect 1227 2498 1239 2502
rect 1243 2498 1423 2502
rect 1427 2498 1599 2502
rect 1603 2498 1631 2502
rect 1635 2498 1655 2502
rect 103 2497 1655 2498
rect 1661 2497 1662 2503
rect 1654 2469 1655 2475
rect 1661 2474 3231 2475
rect 1661 2470 1671 2474
rect 1675 2470 1695 2474
rect 1699 2470 1863 2474
rect 1867 2470 2079 2474
rect 2083 2470 2319 2474
rect 2323 2470 2567 2474
rect 2571 2470 2583 2474
rect 2587 2470 2823 2474
rect 2827 2470 2855 2474
rect 2859 2470 3079 2474
rect 3083 2470 3135 2474
rect 3139 2470 3191 2474
rect 3195 2470 3231 2474
rect 1661 2469 3231 2470
rect 3237 2469 3238 2475
rect 84 2453 85 2459
rect 91 2458 1643 2459
rect 91 2454 111 2458
rect 115 2454 199 2458
rect 203 2454 303 2458
rect 307 2454 327 2458
rect 331 2454 431 2458
rect 435 2454 455 2458
rect 459 2454 559 2458
rect 563 2454 599 2458
rect 603 2454 703 2458
rect 707 2454 767 2458
rect 771 2454 863 2458
rect 867 2454 951 2458
rect 955 2454 1039 2458
rect 1043 2454 1159 2458
rect 1163 2454 1223 2458
rect 1227 2454 1375 2458
rect 1379 2454 1423 2458
rect 1427 2454 1591 2458
rect 1595 2454 1599 2458
rect 1603 2454 1631 2458
rect 1635 2454 1643 2458
rect 91 2453 1643 2454
rect 1649 2453 1650 2459
rect 1642 2429 1643 2435
rect 1649 2434 3219 2435
rect 1649 2430 1671 2434
rect 1675 2430 2231 2434
rect 2235 2430 2319 2434
rect 2323 2430 2391 2434
rect 2395 2430 2543 2434
rect 2547 2430 2567 2434
rect 2571 2430 2687 2434
rect 2691 2430 2823 2434
rect 2827 2430 2967 2434
rect 2971 2430 3079 2434
rect 3083 2430 3111 2434
rect 3115 2430 3191 2434
rect 3195 2430 3219 2434
rect 1649 2429 3219 2430
rect 3225 2429 3226 2435
rect 96 2397 97 2403
rect 103 2402 1655 2403
rect 103 2398 111 2402
rect 115 2398 135 2402
rect 139 2398 199 2402
rect 203 2398 239 2402
rect 243 2398 327 2402
rect 331 2398 359 2402
rect 363 2398 455 2402
rect 459 2398 479 2402
rect 483 2398 591 2402
rect 595 2398 599 2402
rect 603 2398 703 2402
rect 707 2398 767 2402
rect 771 2398 815 2402
rect 819 2398 935 2402
rect 939 2398 951 2402
rect 955 2398 1159 2402
rect 1163 2398 1375 2402
rect 1379 2398 1591 2402
rect 1595 2398 1631 2402
rect 1635 2398 1655 2402
rect 103 2397 1655 2398
rect 1661 2397 1662 2403
rect 1654 2381 1655 2387
rect 1661 2386 3231 2387
rect 1661 2382 1671 2386
rect 1675 2382 2143 2386
rect 2147 2382 2231 2386
rect 2235 2382 2311 2386
rect 2315 2382 2391 2386
rect 2395 2382 2479 2386
rect 2483 2382 2543 2386
rect 2547 2382 2655 2386
rect 2659 2382 2687 2386
rect 2691 2382 2823 2386
rect 2827 2382 2831 2386
rect 2835 2382 2967 2386
rect 2971 2382 3007 2386
rect 3011 2382 3111 2386
rect 3115 2382 3159 2386
rect 3163 2382 3191 2386
rect 3195 2382 3231 2386
rect 1661 2381 3231 2382
rect 3237 2381 3238 2387
rect 84 2349 85 2355
rect 91 2354 1643 2355
rect 91 2350 111 2354
rect 115 2350 135 2354
rect 139 2350 239 2354
rect 243 2350 343 2354
rect 347 2350 359 2354
rect 363 2350 479 2354
rect 483 2350 567 2354
rect 571 2350 591 2354
rect 595 2350 703 2354
rect 707 2350 775 2354
rect 779 2350 815 2354
rect 819 2350 935 2354
rect 939 2350 975 2354
rect 979 2350 1175 2354
rect 1179 2350 1367 2354
rect 1371 2350 1567 2354
rect 1571 2350 1631 2354
rect 1635 2350 1643 2354
rect 91 2349 1643 2350
rect 1649 2349 1650 2355
rect 1642 2347 1650 2349
rect 1642 2341 1643 2347
rect 1649 2346 3219 2347
rect 1649 2342 1671 2346
rect 1675 2342 2143 2346
rect 2147 2342 2183 2346
rect 2187 2342 2311 2346
rect 2315 2342 2335 2346
rect 2339 2342 2479 2346
rect 2483 2342 2623 2346
rect 2627 2342 2655 2346
rect 2659 2342 2767 2346
rect 2771 2342 2831 2346
rect 2835 2342 2919 2346
rect 2923 2342 3007 2346
rect 3011 2342 3159 2346
rect 3163 2342 3191 2346
rect 3195 2342 3219 2346
rect 1649 2341 3219 2342
rect 3225 2341 3226 2347
rect 96 2297 97 2303
rect 103 2302 1655 2303
rect 103 2298 111 2302
rect 115 2298 135 2302
rect 139 2298 343 2302
rect 347 2298 567 2302
rect 571 2298 655 2302
rect 659 2298 775 2302
rect 779 2298 783 2302
rect 787 2298 903 2302
rect 907 2298 975 2302
rect 979 2298 1023 2302
rect 1027 2298 1143 2302
rect 1147 2298 1175 2302
rect 1179 2298 1255 2302
rect 1259 2298 1367 2302
rect 1371 2298 1487 2302
rect 1491 2298 1567 2302
rect 1571 2298 1631 2302
rect 1635 2298 1655 2302
rect 103 2297 1655 2298
rect 1661 2302 3238 2303
rect 1661 2298 1671 2302
rect 1675 2298 2095 2302
rect 2099 2298 2183 2302
rect 2187 2298 2263 2302
rect 2267 2298 2335 2302
rect 2339 2298 2431 2302
rect 2435 2298 2479 2302
rect 2483 2298 2607 2302
rect 2611 2298 2623 2302
rect 2627 2298 2767 2302
rect 2771 2298 2791 2302
rect 2795 2298 2919 2302
rect 2923 2298 2983 2302
rect 2987 2298 3159 2302
rect 3163 2298 3191 2302
rect 3195 2298 3238 2302
rect 1661 2297 3238 2298
rect 1642 2257 1643 2263
rect 1649 2262 3219 2263
rect 1649 2258 1671 2262
rect 1675 2258 2015 2262
rect 2019 2258 2095 2262
rect 2099 2258 2167 2262
rect 2171 2258 2263 2262
rect 2267 2258 2319 2262
rect 2323 2258 2431 2262
rect 2435 2258 2463 2262
rect 2467 2258 2607 2262
rect 2611 2258 2759 2262
rect 2763 2258 2791 2262
rect 2795 2258 2983 2262
rect 2987 2258 3159 2262
rect 3163 2258 3191 2262
rect 3195 2258 3219 2262
rect 1649 2257 3219 2258
rect 3225 2257 3226 2263
rect 84 2245 85 2251
rect 91 2250 1643 2251
rect 91 2246 111 2250
rect 115 2246 551 2250
rect 555 2246 655 2250
rect 659 2246 679 2250
rect 683 2246 783 2250
rect 787 2246 807 2250
rect 811 2246 903 2250
rect 907 2246 927 2250
rect 931 2246 1023 2250
rect 1027 2246 1047 2250
rect 1051 2246 1143 2250
rect 1147 2246 1159 2250
rect 1163 2246 1255 2250
rect 1259 2246 1271 2250
rect 1275 2246 1367 2250
rect 1371 2246 1391 2250
rect 1395 2246 1487 2250
rect 1491 2246 1631 2250
rect 1635 2246 1643 2250
rect 91 2245 1643 2246
rect 1649 2245 1650 2251
rect 1654 2213 1655 2219
rect 1661 2218 3231 2219
rect 1661 2214 1671 2218
rect 1675 2214 1927 2218
rect 1931 2214 2015 2218
rect 2019 2214 2103 2218
rect 2107 2214 2167 2218
rect 2171 2214 2295 2218
rect 2299 2214 2319 2218
rect 2323 2214 2463 2218
rect 2467 2214 2503 2218
rect 2507 2214 2607 2218
rect 2611 2214 2719 2218
rect 2723 2214 2759 2218
rect 2763 2214 2951 2218
rect 2955 2214 3159 2218
rect 3163 2214 3191 2218
rect 3195 2214 3231 2218
rect 1661 2213 3231 2214
rect 3237 2213 3238 2219
rect 96 2197 97 2203
rect 103 2202 1655 2203
rect 103 2198 111 2202
rect 115 2198 455 2202
rect 459 2198 551 2202
rect 555 2198 583 2202
rect 587 2198 679 2202
rect 683 2198 703 2202
rect 707 2198 807 2202
rect 811 2198 823 2202
rect 827 2198 927 2202
rect 931 2198 943 2202
rect 947 2198 1047 2202
rect 1051 2198 1055 2202
rect 1059 2198 1159 2202
rect 1163 2198 1167 2202
rect 1171 2198 1271 2202
rect 1275 2198 1287 2202
rect 1291 2198 1391 2202
rect 1395 2198 1631 2202
rect 1635 2198 1655 2202
rect 103 2197 1655 2198
rect 1661 2197 1662 2203
rect 1642 2173 1643 2179
rect 1649 2178 3219 2179
rect 1649 2174 1671 2178
rect 1675 2174 1847 2178
rect 1851 2174 1927 2178
rect 1931 2174 1999 2178
rect 2003 2174 2103 2178
rect 2107 2174 2151 2178
rect 2155 2174 2295 2178
rect 2299 2174 2447 2178
rect 2451 2174 2503 2178
rect 2507 2174 2599 2178
rect 2603 2174 2719 2178
rect 2723 2174 2951 2178
rect 2955 2174 3159 2178
rect 3163 2174 3191 2178
rect 3195 2174 3219 2178
rect 1649 2173 3219 2174
rect 3225 2173 3226 2179
rect 84 2145 85 2151
rect 91 2150 1643 2151
rect 91 2146 111 2150
rect 115 2146 351 2150
rect 355 2146 455 2150
rect 459 2146 479 2150
rect 483 2146 583 2150
rect 587 2146 599 2150
rect 603 2146 703 2150
rect 707 2146 719 2150
rect 723 2146 823 2150
rect 827 2146 839 2150
rect 843 2146 943 2150
rect 947 2146 951 2150
rect 955 2146 1055 2150
rect 1059 2146 1063 2150
rect 1067 2146 1167 2150
rect 1171 2146 1183 2150
rect 1187 2146 1287 2150
rect 1291 2146 1631 2150
rect 1635 2146 1643 2150
rect 91 2145 1643 2146
rect 1649 2145 1650 2151
rect 1654 2129 1655 2135
rect 1661 2134 3231 2135
rect 1661 2130 1671 2134
rect 1675 2130 1759 2134
rect 1763 2130 1847 2134
rect 1851 2130 1911 2134
rect 1915 2130 1999 2134
rect 2003 2130 2071 2134
rect 2075 2130 2151 2134
rect 2155 2130 2255 2134
rect 2259 2130 2295 2134
rect 2299 2130 2447 2134
rect 2451 2130 2463 2134
rect 2467 2130 2599 2134
rect 2603 2130 2687 2134
rect 2691 2130 2927 2134
rect 2931 2130 3159 2134
rect 3163 2130 3191 2134
rect 3195 2130 3231 2134
rect 1661 2129 3231 2130
rect 3237 2129 3238 2135
rect 1642 2103 1643 2109
rect 1649 2103 1674 2109
rect 96 2093 97 2099
rect 103 2098 1655 2099
rect 103 2094 111 2098
rect 115 2094 247 2098
rect 251 2094 351 2098
rect 355 2094 375 2098
rect 379 2094 479 2098
rect 483 2094 503 2098
rect 507 2094 599 2098
rect 603 2094 623 2098
rect 627 2094 719 2098
rect 723 2094 743 2098
rect 747 2094 839 2098
rect 843 2094 855 2098
rect 859 2094 951 2098
rect 955 2094 967 2098
rect 971 2094 1063 2098
rect 1067 2094 1087 2098
rect 1091 2094 1183 2098
rect 1187 2094 1631 2098
rect 1635 2094 1655 2098
rect 103 2093 1655 2094
rect 1661 2093 1662 2099
rect 1668 2095 1674 2103
rect 1668 2094 3219 2095
rect 1668 2090 1671 2094
rect 1675 2090 1695 2094
rect 1699 2090 1759 2094
rect 1763 2090 1823 2094
rect 1827 2090 1911 2094
rect 1915 2090 1967 2094
rect 1971 2090 2071 2094
rect 2075 2090 2111 2094
rect 2115 2090 2255 2094
rect 2259 2090 2407 2094
rect 2411 2090 2463 2094
rect 2467 2090 2687 2094
rect 2691 2090 2927 2094
rect 2931 2090 3159 2094
rect 3163 2090 3191 2094
rect 3195 2090 3219 2094
rect 1668 2089 3219 2090
rect 3225 2089 3226 2095
rect 84 2045 85 2051
rect 91 2050 1643 2051
rect 91 2046 111 2050
rect 115 2046 175 2050
rect 179 2046 247 2050
rect 251 2046 367 2050
rect 371 2046 375 2050
rect 379 2046 503 2050
rect 507 2046 559 2050
rect 563 2046 623 2050
rect 627 2046 743 2050
rect 747 2046 759 2050
rect 763 2046 855 2050
rect 859 2046 967 2050
rect 971 2046 1087 2050
rect 1091 2046 1183 2050
rect 1187 2046 1399 2050
rect 1403 2046 1599 2050
rect 1603 2046 1631 2050
rect 1635 2046 1643 2050
rect 91 2045 1643 2046
rect 1649 2045 1650 2051
rect 1654 2049 1655 2055
rect 1661 2054 3231 2055
rect 1661 2050 1671 2054
rect 1675 2050 1695 2054
rect 1699 2050 1823 2054
rect 1827 2050 1967 2054
rect 1971 2050 2039 2054
rect 2043 2050 2111 2054
rect 2115 2050 2255 2054
rect 2259 2050 2407 2054
rect 2411 2050 2767 2054
rect 2771 2050 3135 2054
rect 3139 2050 3191 2054
rect 3195 2050 3231 2054
rect 1661 2049 3231 2050
rect 3237 2049 3238 2055
rect 1642 2015 1643 2021
rect 1649 2015 1674 2021
rect 96 2005 97 2011
rect 103 2010 1655 2011
rect 103 2006 111 2010
rect 115 2006 135 2010
rect 139 2006 175 2010
rect 179 2006 231 2010
rect 235 2006 351 2010
rect 355 2006 367 2010
rect 371 2006 463 2010
rect 467 2006 559 2010
rect 563 2006 575 2010
rect 579 2006 687 2010
rect 691 2006 759 2010
rect 763 2006 799 2010
rect 803 2006 911 2010
rect 915 2006 967 2010
rect 971 2006 1183 2010
rect 1187 2006 1399 2010
rect 1403 2006 1599 2010
rect 1603 2006 1631 2010
rect 1635 2006 1655 2010
rect 103 2005 1655 2006
rect 1661 2005 1662 2011
rect 1668 2007 1674 2015
rect 1668 2006 3219 2007
rect 1668 2002 1671 2006
rect 1675 2002 1695 2006
rect 1699 2002 2039 2006
rect 2043 2002 2263 2006
rect 2267 2002 2407 2006
rect 2411 2002 2415 2006
rect 2419 2002 2559 2006
rect 2563 2002 2703 2006
rect 2707 2002 2767 2006
rect 2771 2002 2839 2006
rect 2843 2002 2975 2006
rect 2979 2002 3111 2006
rect 3115 2002 3135 2006
rect 3139 2002 3191 2006
rect 3195 2002 3219 2006
rect 1668 2001 3219 2002
rect 3225 2001 3226 2007
rect 84 1957 85 1963
rect 91 1962 1643 1963
rect 91 1958 111 1962
rect 115 1958 135 1962
rect 139 1958 231 1962
rect 235 1958 351 1962
rect 355 1958 463 1962
rect 467 1958 575 1962
rect 579 1958 687 1962
rect 691 1958 727 1962
rect 731 1958 799 1962
rect 803 1958 855 1962
rect 859 1958 911 1962
rect 915 1958 983 1962
rect 987 1958 1103 1962
rect 1107 1958 1223 1962
rect 1227 1958 1335 1962
rect 1339 1958 1447 1962
rect 1451 1958 1567 1962
rect 1571 1958 1631 1962
rect 1635 1958 1643 1962
rect 91 1957 1643 1958
rect 1649 1957 1650 1963
rect 1654 1961 1655 1967
rect 1661 1966 3231 1967
rect 1661 1962 1671 1966
rect 1675 1962 2239 1966
rect 2243 1962 2263 1966
rect 2267 1962 2391 1966
rect 2395 1962 2415 1966
rect 2419 1962 2543 1966
rect 2547 1962 2559 1966
rect 2563 1962 2695 1966
rect 2699 1962 2703 1966
rect 2707 1962 2839 1966
rect 2843 1962 2847 1966
rect 2851 1962 2975 1966
rect 2979 1962 2999 1966
rect 3003 1962 3111 1966
rect 3115 1962 3191 1966
rect 3195 1962 3231 1966
rect 1661 1961 3231 1962
rect 3237 1961 3238 1967
rect 1642 1917 1643 1923
rect 1649 1922 3219 1923
rect 1649 1918 1671 1922
rect 1675 1918 2151 1922
rect 2155 1918 2239 1922
rect 2243 1918 2311 1922
rect 2315 1918 2391 1922
rect 2395 1918 2471 1922
rect 2475 1918 2543 1922
rect 2547 1918 2639 1922
rect 2643 1918 2695 1922
rect 2699 1918 2815 1922
rect 2819 1918 2847 1922
rect 2851 1918 2999 1922
rect 3003 1918 3159 1922
rect 3163 1918 3191 1922
rect 3195 1918 3219 1922
rect 1649 1917 3219 1918
rect 3225 1917 3226 1923
rect 96 1905 97 1911
rect 103 1910 1655 1911
rect 103 1906 111 1910
rect 115 1906 631 1910
rect 635 1906 727 1910
rect 731 1906 759 1910
rect 763 1906 855 1910
rect 859 1906 879 1910
rect 883 1906 983 1910
rect 987 1906 999 1910
rect 1003 1906 1103 1910
rect 1107 1906 1119 1910
rect 1123 1906 1223 1910
rect 1227 1906 1231 1910
rect 1235 1906 1335 1910
rect 1339 1906 1343 1910
rect 1347 1906 1447 1910
rect 1451 1906 1463 1910
rect 1467 1906 1567 1910
rect 1571 1906 1631 1910
rect 1635 1906 1655 1910
rect 103 1905 1655 1906
rect 1661 1905 1662 1911
rect 1654 1873 1655 1879
rect 1661 1878 3231 1879
rect 1661 1874 1671 1878
rect 1675 1874 2071 1878
rect 2075 1874 2151 1878
rect 2155 1874 2239 1878
rect 2243 1874 2311 1878
rect 2315 1874 2415 1878
rect 2419 1874 2471 1878
rect 2475 1874 2599 1878
rect 2603 1874 2639 1878
rect 2643 1874 2791 1878
rect 2795 1874 2815 1878
rect 2819 1874 2983 1878
rect 2987 1874 2999 1878
rect 3003 1874 3159 1878
rect 3163 1874 3191 1878
rect 3195 1874 3231 1878
rect 1661 1873 3231 1874
rect 3237 1873 3238 1879
rect 84 1853 85 1859
rect 91 1858 1643 1859
rect 91 1854 111 1858
rect 115 1854 527 1858
rect 531 1854 631 1858
rect 635 1854 655 1858
rect 659 1854 759 1858
rect 763 1854 775 1858
rect 779 1854 879 1858
rect 883 1854 895 1858
rect 899 1854 999 1858
rect 1003 1854 1015 1858
rect 1019 1854 1119 1858
rect 1123 1854 1127 1858
rect 1131 1854 1231 1858
rect 1235 1854 1247 1858
rect 1251 1854 1343 1858
rect 1347 1854 1367 1858
rect 1371 1854 1463 1858
rect 1467 1854 1631 1858
rect 1635 1854 1643 1858
rect 91 1853 1643 1854
rect 1649 1853 1650 1859
rect 1642 1833 1643 1839
rect 1649 1838 3219 1839
rect 1649 1834 1671 1838
rect 1675 1834 1983 1838
rect 1987 1834 2071 1838
rect 2075 1834 2135 1838
rect 2139 1834 2239 1838
rect 2243 1834 2287 1838
rect 2291 1834 2415 1838
rect 2419 1834 2431 1838
rect 2435 1834 2583 1838
rect 2587 1834 2599 1838
rect 2603 1834 2735 1838
rect 2739 1834 2791 1838
rect 2795 1834 2983 1838
rect 2987 1834 3159 1838
rect 3163 1834 3191 1838
rect 3195 1834 3219 1838
rect 1649 1833 3219 1834
rect 3225 1833 3226 1839
rect 96 1805 97 1811
rect 103 1810 1655 1811
rect 103 1806 111 1810
rect 115 1806 423 1810
rect 427 1806 527 1810
rect 531 1806 551 1810
rect 555 1806 655 1810
rect 659 1806 679 1810
rect 683 1806 775 1810
rect 779 1806 799 1810
rect 803 1806 895 1810
rect 899 1806 919 1810
rect 923 1806 1015 1810
rect 1019 1806 1031 1810
rect 1035 1806 1127 1810
rect 1131 1806 1143 1810
rect 1147 1806 1247 1810
rect 1251 1806 1263 1810
rect 1267 1806 1367 1810
rect 1371 1806 1631 1810
rect 1635 1806 1655 1810
rect 103 1805 1655 1806
rect 1661 1805 1662 1811
rect 1654 1793 1655 1799
rect 1661 1798 3231 1799
rect 1661 1794 1671 1798
rect 1675 1794 1903 1798
rect 1907 1794 1983 1798
rect 1987 1794 2079 1798
rect 2083 1794 2135 1798
rect 2139 1794 2271 1798
rect 2275 1794 2287 1798
rect 2291 1794 2431 1798
rect 2435 1794 2487 1798
rect 2491 1794 2583 1798
rect 2587 1794 2711 1798
rect 2715 1794 2735 1798
rect 2739 1794 2943 1798
rect 2947 1794 3159 1798
rect 3163 1794 3191 1798
rect 3195 1794 3231 1798
rect 1661 1793 3231 1794
rect 3237 1793 3238 1799
rect 84 1753 85 1759
rect 91 1758 1643 1759
rect 91 1754 111 1758
rect 115 1754 327 1758
rect 331 1754 423 1758
rect 427 1754 455 1758
rect 459 1754 551 1758
rect 555 1754 575 1758
rect 579 1754 679 1758
rect 683 1754 695 1758
rect 699 1754 799 1758
rect 803 1754 815 1758
rect 819 1754 919 1758
rect 923 1754 927 1758
rect 931 1754 1031 1758
rect 1035 1754 1039 1758
rect 1043 1754 1143 1758
rect 1147 1754 1159 1758
rect 1163 1754 1263 1758
rect 1267 1754 1631 1758
rect 1635 1754 1643 1758
rect 91 1753 1643 1754
rect 1649 1753 1650 1759
rect 1642 1751 1650 1753
rect 1642 1745 1643 1751
rect 1649 1750 3219 1751
rect 1649 1746 1671 1750
rect 1675 1746 1815 1750
rect 1819 1746 1903 1750
rect 1907 1746 1967 1750
rect 1971 1746 2079 1750
rect 2083 1746 2127 1750
rect 2131 1746 2271 1750
rect 2275 1746 2303 1750
rect 2307 1746 2487 1750
rect 2491 1746 2503 1750
rect 2507 1746 2711 1750
rect 2715 1746 2935 1750
rect 2939 1746 2943 1750
rect 2947 1746 3159 1750
rect 3163 1746 3191 1750
rect 3195 1746 3219 1750
rect 1649 1745 3219 1746
rect 3225 1745 3226 1751
rect 1654 1710 3238 1711
rect 1654 1707 1671 1710
rect 96 1701 97 1707
rect 103 1706 1655 1707
rect 103 1702 111 1706
rect 115 1702 223 1706
rect 227 1702 327 1706
rect 331 1702 351 1706
rect 355 1702 455 1706
rect 459 1702 471 1706
rect 475 1702 575 1706
rect 579 1702 591 1706
rect 595 1702 695 1706
rect 699 1702 711 1706
rect 715 1702 815 1706
rect 819 1702 823 1706
rect 827 1702 927 1706
rect 931 1702 943 1706
rect 947 1702 1039 1706
rect 1043 1702 1063 1706
rect 1067 1702 1159 1706
rect 1163 1702 1631 1706
rect 1635 1702 1655 1706
rect 103 1701 1655 1702
rect 1661 1706 1671 1707
rect 1675 1706 1735 1710
rect 1739 1706 1815 1710
rect 1819 1706 1879 1710
rect 1883 1706 1967 1710
rect 1971 1706 2023 1710
rect 2027 1706 2127 1710
rect 2131 1706 2167 1710
rect 2171 1706 2303 1710
rect 2307 1706 2311 1710
rect 2315 1706 2463 1710
rect 2467 1706 2503 1710
rect 2507 1706 2711 1710
rect 2715 1706 2935 1710
rect 2939 1706 3159 1710
rect 3163 1706 3191 1710
rect 3195 1706 3238 1710
rect 1661 1705 3238 1706
rect 1661 1701 1662 1705
rect 1642 1665 1643 1671
rect 1649 1670 3219 1671
rect 1649 1666 1671 1670
rect 1675 1666 1695 1670
rect 1699 1666 1735 1670
rect 1739 1666 1879 1670
rect 1883 1666 1895 1670
rect 1899 1666 2023 1670
rect 2027 1666 2127 1670
rect 2131 1666 2167 1670
rect 2171 1666 2311 1670
rect 2315 1666 2367 1670
rect 2371 1666 2463 1670
rect 2467 1666 2615 1670
rect 2619 1666 2871 1670
rect 2875 1666 3135 1670
rect 3139 1666 3191 1670
rect 3195 1666 3219 1670
rect 1649 1665 3219 1666
rect 3225 1665 3226 1671
rect 84 1649 85 1655
rect 91 1654 1643 1655
rect 91 1650 111 1654
rect 115 1650 135 1654
rect 139 1650 223 1654
rect 227 1650 247 1654
rect 251 1650 351 1654
rect 355 1650 383 1654
rect 387 1650 471 1654
rect 475 1650 535 1654
rect 539 1650 591 1654
rect 595 1650 711 1654
rect 715 1650 823 1654
rect 827 1650 919 1654
rect 923 1650 943 1654
rect 947 1650 1063 1654
rect 1067 1650 1143 1654
rect 1147 1650 1383 1654
rect 1387 1650 1599 1654
rect 1603 1650 1631 1654
rect 1635 1650 1643 1654
rect 91 1649 1643 1650
rect 1649 1649 1650 1655
rect 1654 1621 1655 1627
rect 1661 1626 3231 1627
rect 1661 1622 1671 1626
rect 1675 1622 1695 1626
rect 1699 1622 1895 1626
rect 1899 1622 2127 1626
rect 2131 1622 2319 1626
rect 2323 1622 2367 1626
rect 2371 1622 2519 1626
rect 2523 1622 2615 1626
rect 2619 1622 2711 1626
rect 2715 1622 2871 1626
rect 2875 1622 2911 1626
rect 2915 1622 3111 1626
rect 3115 1622 3135 1626
rect 3139 1622 3191 1626
rect 3195 1622 3231 1626
rect 1661 1621 3231 1622
rect 3237 1621 3238 1627
rect 96 1601 97 1607
rect 103 1606 1655 1607
rect 103 1602 111 1606
rect 115 1602 135 1606
rect 139 1602 247 1606
rect 251 1602 303 1606
rect 307 1602 383 1606
rect 387 1602 503 1606
rect 507 1602 535 1606
rect 539 1602 695 1606
rect 699 1602 711 1606
rect 715 1602 887 1606
rect 891 1602 919 1606
rect 923 1602 1063 1606
rect 1067 1602 1143 1606
rect 1147 1602 1239 1606
rect 1243 1602 1383 1606
rect 1387 1602 1415 1606
rect 1419 1602 1591 1606
rect 1595 1602 1599 1606
rect 1603 1602 1631 1606
rect 1635 1602 1655 1606
rect 103 1601 1655 1602
rect 1661 1601 1662 1607
rect 1642 1581 1643 1587
rect 1649 1586 3219 1587
rect 1649 1582 1671 1586
rect 1675 1582 2271 1586
rect 2275 1582 2319 1586
rect 2323 1582 2415 1586
rect 2419 1582 2519 1586
rect 2523 1582 2559 1586
rect 2563 1582 2695 1586
rect 2699 1582 2711 1586
rect 2715 1582 2839 1586
rect 2843 1582 2911 1586
rect 2915 1582 2983 1586
rect 2987 1582 3111 1586
rect 3115 1582 3191 1586
rect 3195 1582 3219 1586
rect 1649 1581 3219 1582
rect 3225 1581 3226 1587
rect 84 1549 85 1555
rect 91 1554 1643 1555
rect 91 1550 111 1554
rect 115 1550 135 1554
rect 139 1550 303 1554
rect 307 1550 503 1554
rect 507 1550 679 1554
rect 683 1550 695 1554
rect 699 1550 807 1554
rect 811 1550 887 1554
rect 891 1550 927 1554
rect 931 1550 1047 1554
rect 1051 1550 1063 1554
rect 1067 1550 1167 1554
rect 1171 1550 1239 1554
rect 1243 1550 1279 1554
rect 1283 1550 1399 1554
rect 1403 1550 1415 1554
rect 1419 1550 1519 1554
rect 1523 1550 1591 1554
rect 1595 1550 1631 1554
rect 1635 1550 1643 1554
rect 91 1549 1643 1550
rect 1649 1549 1650 1555
rect 1654 1533 1655 1539
rect 1661 1538 3231 1539
rect 1661 1534 1671 1538
rect 1675 1534 2167 1538
rect 2171 1534 2271 1538
rect 2275 1534 2279 1538
rect 2283 1534 2391 1538
rect 2395 1534 2415 1538
rect 2419 1534 2503 1538
rect 2507 1534 2559 1538
rect 2563 1534 2615 1538
rect 2619 1534 2695 1538
rect 2699 1534 2735 1538
rect 2739 1534 2839 1538
rect 2843 1534 2855 1538
rect 2859 1534 2983 1538
rect 2987 1534 3111 1538
rect 3115 1534 3191 1538
rect 3195 1534 3231 1538
rect 1661 1533 3231 1534
rect 3237 1533 3238 1539
rect 96 1501 97 1507
rect 103 1506 1655 1507
rect 103 1502 111 1506
rect 115 1502 575 1506
rect 579 1502 679 1506
rect 683 1502 703 1506
rect 707 1502 807 1506
rect 811 1502 831 1506
rect 835 1502 927 1506
rect 931 1502 951 1506
rect 955 1502 1047 1506
rect 1051 1502 1071 1506
rect 1075 1502 1167 1506
rect 1171 1502 1183 1506
rect 1187 1502 1279 1506
rect 1283 1502 1295 1506
rect 1299 1502 1399 1506
rect 1403 1502 1415 1506
rect 1419 1502 1519 1506
rect 1523 1502 1631 1506
rect 1635 1502 1655 1506
rect 103 1501 1655 1502
rect 1661 1501 1662 1507
rect 1642 1489 1643 1495
rect 1649 1494 3219 1495
rect 1649 1490 1671 1494
rect 1675 1490 2087 1494
rect 2091 1490 2167 1494
rect 2171 1490 2231 1494
rect 2235 1490 2279 1494
rect 2283 1490 2375 1494
rect 2379 1490 2391 1494
rect 2395 1490 2503 1494
rect 2507 1490 2511 1494
rect 2515 1490 2615 1494
rect 2619 1490 2655 1494
rect 2659 1490 2735 1494
rect 2739 1490 2799 1494
rect 2803 1490 2855 1494
rect 2859 1490 2983 1494
rect 2987 1490 3111 1494
rect 3115 1490 3191 1494
rect 3195 1490 3219 1494
rect 1649 1489 3219 1490
rect 3225 1489 3226 1495
rect 84 1449 85 1455
rect 91 1454 1643 1455
rect 91 1450 111 1454
rect 115 1450 479 1454
rect 483 1450 575 1454
rect 579 1450 607 1454
rect 611 1450 703 1454
rect 707 1450 727 1454
rect 731 1450 831 1454
rect 835 1450 847 1454
rect 851 1450 951 1454
rect 955 1450 967 1454
rect 971 1450 1071 1454
rect 1075 1450 1079 1454
rect 1083 1450 1183 1454
rect 1187 1450 1191 1454
rect 1195 1450 1295 1454
rect 1299 1450 1311 1454
rect 1315 1450 1415 1454
rect 1419 1450 1631 1454
rect 1635 1450 1643 1454
rect 91 1449 1643 1450
rect 1649 1449 1650 1455
rect 1654 1445 1655 1451
rect 1661 1450 3231 1451
rect 1661 1446 1671 1450
rect 1675 1446 1983 1450
rect 1987 1446 2087 1450
rect 2091 1446 2095 1450
rect 2099 1446 2207 1450
rect 2211 1446 2231 1450
rect 2235 1446 2335 1450
rect 2339 1446 2375 1450
rect 2379 1446 2479 1450
rect 2483 1446 2511 1450
rect 2515 1446 2639 1450
rect 2643 1446 2655 1450
rect 2659 1446 2799 1450
rect 2803 1446 2815 1450
rect 2819 1446 2999 1450
rect 3003 1446 3159 1450
rect 3163 1446 3191 1450
rect 3195 1446 3231 1450
rect 1661 1445 3231 1446
rect 3237 1445 3238 1451
rect 1642 1407 1643 1413
rect 1649 1407 1674 1413
rect 96 1397 97 1403
rect 103 1402 1655 1403
rect 103 1398 111 1402
rect 115 1398 375 1402
rect 379 1398 479 1402
rect 483 1398 503 1402
rect 507 1398 607 1402
rect 611 1398 623 1402
rect 627 1398 727 1402
rect 731 1398 743 1402
rect 747 1398 847 1402
rect 851 1398 863 1402
rect 867 1398 967 1402
rect 971 1398 975 1402
rect 979 1398 1079 1402
rect 1083 1398 1095 1402
rect 1099 1398 1191 1402
rect 1195 1398 1215 1402
rect 1219 1398 1311 1402
rect 1315 1398 1631 1402
rect 1635 1398 1655 1402
rect 103 1397 1655 1398
rect 1661 1397 1662 1403
rect 1668 1395 1674 1407
rect 1668 1394 3219 1395
rect 1668 1390 1671 1394
rect 1675 1390 1879 1394
rect 1883 1390 1983 1394
rect 1987 1390 1991 1394
rect 1995 1390 2095 1394
rect 2099 1390 2103 1394
rect 2107 1390 2207 1394
rect 2211 1390 2239 1394
rect 2243 1390 2335 1394
rect 2339 1390 2391 1394
rect 2395 1390 2479 1394
rect 2483 1390 2567 1394
rect 2571 1390 2639 1394
rect 2643 1390 2767 1394
rect 2771 1390 2815 1394
rect 2819 1390 2975 1394
rect 2979 1390 2999 1394
rect 3003 1390 3159 1394
rect 3163 1390 3191 1394
rect 3195 1390 3219 1394
rect 1668 1389 3219 1390
rect 3225 1389 3226 1395
rect 84 1349 85 1355
rect 91 1354 1643 1355
rect 91 1350 111 1354
rect 115 1350 271 1354
rect 275 1350 375 1354
rect 379 1350 399 1354
rect 403 1350 503 1354
rect 507 1350 527 1354
rect 531 1350 623 1354
rect 627 1350 647 1354
rect 651 1350 743 1354
rect 747 1350 767 1354
rect 771 1350 863 1354
rect 867 1350 879 1354
rect 883 1350 975 1354
rect 979 1350 991 1354
rect 995 1350 1095 1354
rect 1099 1350 1111 1354
rect 1115 1350 1215 1354
rect 1219 1350 1631 1354
rect 1635 1350 1643 1354
rect 91 1349 1643 1350
rect 1649 1349 1650 1355
rect 1654 1337 1655 1343
rect 1661 1342 3231 1343
rect 1661 1338 1671 1342
rect 1675 1338 1775 1342
rect 1779 1338 1879 1342
rect 1883 1338 1887 1342
rect 1891 1338 1991 1342
rect 1995 1338 2095 1342
rect 2099 1338 2103 1342
rect 2107 1338 2199 1342
rect 2203 1338 2239 1342
rect 2243 1338 2303 1342
rect 2307 1338 2391 1342
rect 2395 1338 2407 1342
rect 2411 1338 2511 1342
rect 2515 1338 2567 1342
rect 2571 1338 2767 1342
rect 2771 1338 2975 1342
rect 2979 1338 3159 1342
rect 3163 1338 3191 1342
rect 3195 1338 3231 1342
rect 1661 1337 3231 1338
rect 3237 1337 3238 1343
rect 1642 1307 1643 1313
rect 1649 1307 1674 1313
rect 96 1297 97 1303
rect 103 1302 1655 1303
rect 103 1298 111 1302
rect 115 1298 175 1302
rect 179 1298 271 1302
rect 275 1298 303 1302
rect 307 1298 399 1302
rect 403 1298 423 1302
rect 427 1298 527 1302
rect 531 1298 543 1302
rect 547 1298 647 1302
rect 651 1298 663 1302
rect 667 1298 767 1302
rect 771 1298 775 1302
rect 779 1298 879 1302
rect 883 1298 887 1302
rect 891 1298 991 1302
rect 995 1298 1007 1302
rect 1011 1298 1111 1302
rect 1115 1298 1631 1302
rect 1635 1298 1655 1302
rect 103 1297 1655 1298
rect 1661 1297 1662 1303
rect 1668 1295 1674 1307
rect 1668 1294 3219 1295
rect 1668 1290 1671 1294
rect 1675 1290 1695 1294
rect 1699 1290 1775 1294
rect 1779 1290 1791 1294
rect 1795 1290 1887 1294
rect 1891 1290 1935 1294
rect 1939 1290 1991 1294
rect 1995 1290 2095 1294
rect 2099 1290 2103 1294
rect 2107 1290 2199 1294
rect 2203 1290 2295 1294
rect 2299 1290 2303 1294
rect 2307 1290 2407 1294
rect 2411 1290 2495 1294
rect 2499 1290 2511 1294
rect 2515 1290 2711 1294
rect 2715 1290 2935 1294
rect 2939 1290 3159 1294
rect 3163 1290 3191 1294
rect 3195 1290 3219 1294
rect 1668 1289 3219 1290
rect 3225 1289 3226 1295
rect 84 1245 85 1251
rect 91 1250 1643 1251
rect 91 1246 111 1250
rect 115 1246 135 1250
rect 139 1246 175 1250
rect 179 1246 231 1250
rect 235 1246 303 1250
rect 307 1246 359 1250
rect 363 1246 423 1250
rect 427 1246 503 1250
rect 507 1246 543 1250
rect 547 1246 663 1250
rect 667 1246 775 1250
rect 779 1246 831 1250
rect 835 1246 887 1250
rect 891 1246 1007 1250
rect 1011 1246 1015 1250
rect 1019 1246 1207 1250
rect 1211 1246 1407 1250
rect 1411 1246 1599 1250
rect 1603 1246 1631 1250
rect 1635 1246 1643 1250
rect 91 1245 1643 1246
rect 1649 1245 1650 1251
rect 1654 1233 1655 1239
rect 1661 1238 3231 1239
rect 1661 1234 1671 1238
rect 1675 1234 1695 1238
rect 1699 1234 1791 1238
rect 1795 1234 1935 1238
rect 1939 1234 1983 1238
rect 1987 1234 2103 1238
rect 2107 1234 2255 1238
rect 2259 1234 2295 1238
rect 2299 1234 2495 1238
rect 2499 1234 2711 1238
rect 2715 1234 2919 1238
rect 2923 1234 2935 1238
rect 2939 1234 3135 1238
rect 3139 1234 3159 1238
rect 3163 1234 3191 1238
rect 3195 1234 3231 1238
rect 1661 1233 3231 1234
rect 3237 1233 3238 1239
rect 1642 1207 1643 1213
rect 1649 1207 1674 1213
rect 96 1197 97 1203
rect 103 1202 1655 1203
rect 103 1198 111 1202
rect 115 1198 135 1202
rect 139 1198 231 1202
rect 235 1198 359 1202
rect 363 1198 503 1202
rect 507 1198 663 1202
rect 667 1198 727 1202
rect 731 1198 831 1202
rect 835 1198 855 1202
rect 859 1198 983 1202
rect 987 1198 1015 1202
rect 1019 1198 1103 1202
rect 1107 1198 1207 1202
rect 1211 1198 1223 1202
rect 1227 1198 1335 1202
rect 1339 1198 1407 1202
rect 1411 1198 1447 1202
rect 1451 1198 1567 1202
rect 1571 1198 1599 1202
rect 1603 1198 1631 1202
rect 1635 1198 1655 1202
rect 103 1197 1655 1198
rect 1661 1197 1662 1203
rect 1668 1195 1674 1207
rect 1668 1194 3219 1195
rect 1668 1190 1671 1194
rect 1675 1190 1695 1194
rect 1699 1190 1983 1194
rect 1987 1190 2247 1194
rect 2251 1190 2255 1194
rect 2259 1190 2399 1194
rect 2403 1190 2495 1194
rect 2499 1190 2551 1194
rect 2555 1190 2695 1194
rect 2699 1190 2711 1194
rect 2715 1190 2847 1194
rect 2851 1190 2919 1194
rect 2923 1190 2999 1194
rect 3003 1190 3135 1194
rect 3139 1190 3191 1194
rect 3195 1190 3219 1194
rect 1668 1189 3219 1190
rect 3225 1189 3226 1195
rect 84 1145 85 1151
rect 91 1150 1643 1151
rect 91 1146 111 1150
rect 115 1146 631 1150
rect 635 1146 727 1150
rect 731 1146 759 1150
rect 763 1146 855 1150
rect 859 1146 879 1150
rect 883 1146 983 1150
rect 987 1146 999 1150
rect 1003 1146 1103 1150
rect 1107 1146 1119 1150
rect 1123 1146 1223 1150
rect 1227 1146 1231 1150
rect 1235 1146 1335 1150
rect 1339 1146 1343 1150
rect 1347 1146 1447 1150
rect 1451 1146 1463 1150
rect 1467 1146 1567 1150
rect 1571 1146 1631 1150
rect 1635 1146 1643 1150
rect 91 1145 1643 1146
rect 1649 1145 1650 1151
rect 1654 1149 1655 1155
rect 1661 1154 3231 1155
rect 1661 1150 1671 1154
rect 1675 1150 2175 1154
rect 2179 1150 2247 1154
rect 2251 1150 2335 1154
rect 2339 1150 2399 1154
rect 2403 1150 2495 1154
rect 2499 1150 2551 1154
rect 2555 1150 2655 1154
rect 2659 1150 2695 1154
rect 2699 1150 2815 1154
rect 2819 1150 2847 1154
rect 2851 1150 2975 1154
rect 2979 1150 2999 1154
rect 3003 1150 3135 1154
rect 3139 1150 3191 1154
rect 3195 1150 3231 1154
rect 1661 1149 3231 1150
rect 3237 1149 3238 1155
rect 1642 1105 1643 1111
rect 1649 1110 3219 1111
rect 1649 1106 1671 1110
rect 1675 1106 2071 1110
rect 2075 1106 2175 1110
rect 2179 1106 2191 1110
rect 2195 1106 2327 1110
rect 2331 1106 2335 1110
rect 2339 1106 2479 1110
rect 2483 1106 2495 1110
rect 2499 1106 2639 1110
rect 2643 1106 2655 1110
rect 2659 1106 2815 1110
rect 2819 1106 2975 1110
rect 2979 1106 2999 1110
rect 3003 1106 3135 1110
rect 3139 1106 3159 1110
rect 3163 1106 3191 1110
rect 3195 1106 3219 1110
rect 1649 1105 3219 1106
rect 3225 1105 3226 1111
rect 96 1093 97 1099
rect 103 1098 1655 1099
rect 103 1094 111 1098
rect 115 1094 527 1098
rect 531 1094 631 1098
rect 635 1094 655 1098
rect 659 1094 759 1098
rect 763 1094 775 1098
rect 779 1094 879 1098
rect 883 1094 895 1098
rect 899 1094 999 1098
rect 1003 1094 1015 1098
rect 1019 1094 1119 1098
rect 1123 1094 1127 1098
rect 1131 1094 1231 1098
rect 1235 1094 1247 1098
rect 1251 1094 1343 1098
rect 1347 1094 1367 1098
rect 1371 1094 1463 1098
rect 1467 1094 1631 1098
rect 1635 1094 1655 1098
rect 103 1093 1655 1094
rect 1661 1093 1662 1099
rect 1654 1053 1655 1059
rect 1661 1058 3231 1059
rect 1661 1054 1671 1058
rect 1675 1054 1975 1058
rect 1979 1054 2071 1058
rect 2075 1054 2095 1058
rect 2099 1054 2191 1058
rect 2195 1054 2215 1058
rect 2219 1054 2327 1058
rect 2331 1054 2343 1058
rect 2347 1054 2479 1058
rect 2483 1054 2487 1058
rect 2491 1054 2639 1058
rect 2643 1054 2647 1058
rect 2651 1054 2815 1058
rect 2819 1054 2823 1058
rect 2827 1054 2999 1058
rect 3003 1054 3159 1058
rect 3163 1054 3191 1058
rect 3195 1054 3231 1058
rect 1661 1053 3231 1054
rect 3237 1053 3238 1059
rect 84 1045 85 1051
rect 91 1050 1643 1051
rect 91 1046 111 1050
rect 115 1046 423 1050
rect 427 1046 527 1050
rect 531 1046 551 1050
rect 555 1046 655 1050
rect 659 1046 679 1050
rect 683 1046 775 1050
rect 779 1046 799 1050
rect 803 1046 895 1050
rect 899 1046 919 1050
rect 923 1046 1015 1050
rect 1019 1046 1031 1050
rect 1035 1046 1127 1050
rect 1131 1046 1143 1050
rect 1147 1046 1247 1050
rect 1251 1046 1263 1050
rect 1267 1046 1367 1050
rect 1371 1046 1631 1050
rect 1635 1046 1643 1050
rect 91 1045 1643 1046
rect 1649 1045 1650 1051
rect 1642 1009 1643 1015
rect 1649 1014 3219 1015
rect 1649 1010 1671 1014
rect 1675 1010 1895 1014
rect 1899 1010 1975 1014
rect 1979 1010 2047 1014
rect 2051 1010 2095 1014
rect 2099 1010 2199 1014
rect 2203 1010 2215 1014
rect 2219 1010 2343 1014
rect 2347 1010 2487 1014
rect 2491 1010 2495 1014
rect 2499 1010 2647 1014
rect 2651 1010 2823 1014
rect 2827 1010 2999 1014
rect 3003 1010 3159 1014
rect 3163 1010 3191 1014
rect 3195 1010 3219 1014
rect 1649 1009 3219 1010
rect 3225 1009 3226 1015
rect 96 993 97 999
rect 103 998 1655 999
rect 103 994 111 998
rect 115 994 327 998
rect 331 994 423 998
rect 427 994 455 998
rect 459 994 551 998
rect 555 994 575 998
rect 579 994 679 998
rect 683 994 695 998
rect 699 994 799 998
rect 803 994 815 998
rect 819 994 919 998
rect 923 994 927 998
rect 931 994 1031 998
rect 1035 994 1039 998
rect 1043 994 1143 998
rect 1147 994 1159 998
rect 1163 994 1263 998
rect 1267 994 1631 998
rect 1635 994 1655 998
rect 103 993 1655 994
rect 1661 993 1662 999
rect 1654 969 1655 975
rect 1661 974 3231 975
rect 1661 970 1671 974
rect 1675 970 1791 974
rect 1795 970 1895 974
rect 1899 970 1919 974
rect 1923 970 2047 974
rect 2051 970 2071 974
rect 2075 970 2199 974
rect 2203 970 2255 974
rect 2259 970 2343 974
rect 2347 970 2463 974
rect 2467 970 2495 974
rect 2499 970 2647 974
rect 2651 970 2695 974
rect 2699 970 2935 974
rect 2939 970 3159 974
rect 3163 970 3191 974
rect 3195 970 3231 974
rect 1661 969 3231 970
rect 3237 969 3238 975
rect 84 941 85 947
rect 91 946 1643 947
rect 91 942 111 946
rect 115 942 223 946
rect 227 942 327 946
rect 331 942 351 946
rect 355 942 455 946
rect 459 942 471 946
rect 475 942 575 946
rect 579 942 591 946
rect 595 942 695 946
rect 699 942 711 946
rect 715 942 815 946
rect 819 942 823 946
rect 827 942 927 946
rect 931 942 943 946
rect 947 942 1039 946
rect 1043 942 1063 946
rect 1067 942 1159 946
rect 1163 942 1631 946
rect 1635 942 1643 946
rect 91 941 1643 942
rect 1649 941 1650 947
rect 1642 921 1643 927
rect 1649 926 3219 927
rect 1649 922 1671 926
rect 1675 922 1719 926
rect 1723 922 1791 926
rect 1795 922 1871 926
rect 1875 922 1919 926
rect 1923 922 2039 926
rect 2043 922 2071 926
rect 2075 922 2223 926
rect 2227 922 2255 926
rect 2259 922 2439 926
rect 2443 922 2463 926
rect 2467 922 2671 926
rect 2675 922 2695 926
rect 2699 922 2911 926
rect 2915 922 2935 926
rect 2939 922 3159 926
rect 3163 922 3191 926
rect 3195 922 3219 926
rect 1649 921 3219 922
rect 3225 921 3226 927
rect 96 889 97 895
rect 103 894 1655 895
rect 103 890 111 894
rect 115 890 135 894
rect 139 890 223 894
rect 227 890 247 894
rect 251 890 351 894
rect 355 890 383 894
rect 387 890 471 894
rect 475 890 535 894
rect 539 890 591 894
rect 595 890 711 894
rect 715 890 823 894
rect 827 890 919 894
rect 923 890 943 894
rect 947 890 1063 894
rect 1067 890 1143 894
rect 1147 890 1383 894
rect 1387 890 1599 894
rect 1603 890 1631 894
rect 1635 890 1655 894
rect 103 889 1655 890
rect 1661 889 1662 895
rect 1654 887 1662 889
rect 1654 881 1655 887
rect 1661 886 3231 887
rect 1661 882 1671 886
rect 1675 882 1695 886
rect 1699 882 1719 886
rect 1723 882 1871 886
rect 1875 882 2015 886
rect 2019 882 2039 886
rect 2043 882 2223 886
rect 2227 882 2367 886
rect 2371 882 2439 886
rect 2443 882 2671 886
rect 2675 882 2727 886
rect 2731 882 2911 886
rect 2915 882 3087 886
rect 3091 882 3159 886
rect 3163 882 3191 886
rect 3195 882 3231 886
rect 1661 881 3231 882
rect 3237 881 3238 887
rect 84 845 85 851
rect 91 850 1643 851
rect 91 846 111 850
rect 115 846 135 850
rect 139 846 247 850
rect 251 846 303 850
rect 307 846 383 850
rect 387 846 503 850
rect 507 846 535 850
rect 539 846 695 850
rect 699 846 711 850
rect 715 846 879 850
rect 883 846 919 850
rect 923 846 1047 850
rect 1051 846 1143 850
rect 1147 846 1199 850
rect 1203 846 1335 850
rect 1339 846 1383 850
rect 1387 846 1471 850
rect 1475 846 1599 850
rect 1603 846 1631 850
rect 1635 846 1643 850
rect 91 845 1643 846
rect 1649 845 1650 851
rect 1642 829 1643 835
rect 1649 834 3219 835
rect 1649 830 1671 834
rect 1675 830 1695 834
rect 1699 830 2015 834
rect 2019 830 2279 834
rect 2283 830 2367 834
rect 2371 830 2439 834
rect 2443 830 2583 834
rect 2587 830 2719 834
rect 2723 830 2727 834
rect 2731 830 2847 834
rect 2851 830 2975 834
rect 2979 830 3087 834
rect 3091 830 3111 834
rect 3115 830 3191 834
rect 3195 830 3219 834
rect 1649 829 3219 830
rect 3225 829 3226 835
rect 96 789 97 795
rect 103 794 1655 795
rect 103 790 111 794
rect 115 790 135 794
rect 139 790 303 794
rect 307 790 503 794
rect 507 790 679 794
rect 683 790 695 794
rect 699 790 807 794
rect 811 790 879 794
rect 883 790 927 794
rect 931 790 1047 794
rect 1051 790 1167 794
rect 1171 790 1199 794
rect 1203 790 1279 794
rect 1283 790 1335 794
rect 1339 790 1399 794
rect 1403 790 1471 794
rect 1475 790 1519 794
rect 1523 790 1599 794
rect 1603 790 1631 794
rect 1635 790 1655 794
rect 103 789 1655 790
rect 1661 791 1662 795
rect 1661 790 3238 791
rect 1661 789 1671 790
rect 1654 786 1671 789
rect 1675 786 2199 790
rect 2203 786 2279 790
rect 2283 786 2359 790
rect 2363 786 2439 790
rect 2443 786 2511 790
rect 2515 786 2583 790
rect 2587 786 2655 790
rect 2659 786 2719 790
rect 2723 786 2791 790
rect 2795 786 2847 790
rect 2851 786 2919 790
rect 2923 786 2975 790
rect 2979 786 3047 790
rect 3051 786 3111 790
rect 3115 786 3159 790
rect 3163 786 3191 790
rect 3195 786 3238 790
rect 1654 785 3238 786
rect 84 741 85 747
rect 91 746 1643 747
rect 91 742 111 746
rect 115 742 575 746
rect 579 742 679 746
rect 683 742 703 746
rect 707 742 807 746
rect 811 742 831 746
rect 835 742 927 746
rect 931 742 951 746
rect 955 742 1047 746
rect 1051 742 1071 746
rect 1075 742 1167 746
rect 1171 742 1183 746
rect 1187 742 1279 746
rect 1283 742 1295 746
rect 1299 742 1399 746
rect 1403 742 1415 746
rect 1419 742 1519 746
rect 1523 742 1631 746
rect 1635 742 1643 746
rect 91 741 1643 742
rect 1649 746 3226 747
rect 1649 742 1671 746
rect 1675 742 2127 746
rect 2131 742 2199 746
rect 2203 742 2287 746
rect 2291 742 2359 746
rect 2363 742 2447 746
rect 2451 742 2511 746
rect 2515 742 2599 746
rect 2603 742 2655 746
rect 2659 742 2759 746
rect 2763 742 2791 746
rect 2795 742 2919 746
rect 2923 742 3047 746
rect 3051 742 3159 746
rect 3163 742 3191 746
rect 3195 742 3226 746
rect 1649 741 3226 742
rect 1654 701 1655 707
rect 1661 706 3231 707
rect 1661 702 1671 706
rect 1675 702 2023 706
rect 2027 702 2127 706
rect 2131 702 2151 706
rect 2155 702 2287 706
rect 2291 702 2295 706
rect 2299 702 2447 706
rect 2451 702 2599 706
rect 2603 702 2615 706
rect 2619 702 2759 706
rect 2763 702 2799 706
rect 2803 702 2919 706
rect 2923 702 2991 706
rect 2995 702 3159 706
rect 3163 702 3191 706
rect 3195 702 3231 706
rect 1661 701 3231 702
rect 3237 701 3238 707
rect 96 689 97 695
rect 103 694 1655 695
rect 103 690 111 694
rect 115 690 479 694
rect 483 690 575 694
rect 579 690 607 694
rect 611 690 703 694
rect 707 690 727 694
rect 731 690 831 694
rect 835 690 847 694
rect 851 690 951 694
rect 955 690 967 694
rect 971 690 1071 694
rect 1075 690 1079 694
rect 1083 690 1183 694
rect 1187 690 1191 694
rect 1195 690 1295 694
rect 1299 690 1311 694
rect 1315 690 1415 694
rect 1419 690 1631 694
rect 1635 690 1655 694
rect 103 689 1655 690
rect 1661 689 1662 695
rect 1642 653 1643 659
rect 1649 658 3219 659
rect 1649 654 1671 658
rect 1675 654 1919 658
rect 1923 654 2023 658
rect 2027 654 2047 658
rect 2051 654 2151 658
rect 2155 654 2183 658
rect 2187 654 2295 658
rect 2299 654 2327 658
rect 2331 654 2447 658
rect 2451 654 2471 658
rect 2475 654 2615 658
rect 2619 654 2759 658
rect 2763 654 2799 658
rect 2803 654 2991 658
rect 2995 654 3159 658
rect 3163 654 3191 658
rect 3195 654 3219 658
rect 1649 653 3219 654
rect 3225 653 3226 659
rect 84 637 85 643
rect 91 642 1643 643
rect 91 638 111 642
rect 115 638 375 642
rect 379 638 479 642
rect 483 638 503 642
rect 507 638 607 642
rect 611 638 623 642
rect 627 638 727 642
rect 731 638 743 642
rect 747 638 847 642
rect 851 638 863 642
rect 867 638 967 642
rect 971 638 975 642
rect 979 638 1079 642
rect 1083 638 1095 642
rect 1099 638 1191 642
rect 1195 638 1215 642
rect 1219 638 1311 642
rect 1315 638 1631 642
rect 1635 638 1643 642
rect 91 637 1643 638
rect 1649 637 1650 643
rect 1654 609 1655 615
rect 1661 614 3231 615
rect 1661 610 1671 614
rect 1675 610 1847 614
rect 1851 610 1919 614
rect 1923 610 2015 614
rect 2019 610 2047 614
rect 2051 610 2183 614
rect 2187 610 2327 614
rect 2331 610 2359 614
rect 2363 610 2471 614
rect 2475 610 2551 614
rect 2555 610 2615 614
rect 2619 610 2751 614
rect 2755 610 2759 614
rect 2763 610 2959 614
rect 2963 610 3159 614
rect 3163 610 3191 614
rect 3195 610 3231 614
rect 1661 609 3231 610
rect 3237 609 3238 615
rect 96 589 97 595
rect 103 594 1655 595
rect 103 590 111 594
rect 115 590 271 594
rect 275 590 375 594
rect 379 590 399 594
rect 403 590 503 594
rect 507 590 527 594
rect 531 590 623 594
rect 627 590 647 594
rect 651 590 743 594
rect 747 590 767 594
rect 771 590 863 594
rect 867 590 879 594
rect 883 590 975 594
rect 979 590 991 594
rect 995 590 1095 594
rect 1099 590 1111 594
rect 1115 590 1215 594
rect 1219 590 1631 594
rect 1635 590 1655 594
rect 103 589 1655 590
rect 1661 589 1662 595
rect 1642 569 1643 575
rect 1649 574 3219 575
rect 1649 570 1671 574
rect 1675 570 1767 574
rect 1771 570 1847 574
rect 1851 570 1927 574
rect 1931 570 2015 574
rect 2019 570 2087 574
rect 2091 570 2183 574
rect 2187 570 2247 574
rect 2251 570 2359 574
rect 2363 570 2407 574
rect 2411 570 2551 574
rect 2555 570 2567 574
rect 2571 570 2751 574
rect 2755 570 2959 574
rect 2963 570 3159 574
rect 3163 570 3191 574
rect 3195 570 3219 574
rect 1649 569 3219 570
rect 3225 569 3226 575
rect 84 537 85 543
rect 91 542 1643 543
rect 91 538 111 542
rect 115 538 175 542
rect 179 538 271 542
rect 275 538 303 542
rect 307 538 399 542
rect 403 538 423 542
rect 427 538 527 542
rect 531 538 543 542
rect 547 538 647 542
rect 651 538 663 542
rect 667 538 767 542
rect 771 538 775 542
rect 779 538 879 542
rect 883 538 887 542
rect 891 538 991 542
rect 995 538 1007 542
rect 1011 538 1111 542
rect 1115 538 1631 542
rect 1635 538 1643 542
rect 91 537 1643 538
rect 1649 537 1650 543
rect 1654 529 1655 535
rect 1661 534 3231 535
rect 1661 530 1671 534
rect 1675 530 1695 534
rect 1699 530 1767 534
rect 1771 530 1887 534
rect 1891 530 1927 534
rect 1931 530 2087 534
rect 2091 530 2103 534
rect 2107 530 2247 534
rect 2251 530 2343 534
rect 2347 530 2407 534
rect 2411 530 2567 534
rect 2571 530 2599 534
rect 2603 530 2863 534
rect 2867 530 3135 534
rect 3139 530 3191 534
rect 3195 530 3231 534
rect 1661 529 3231 530
rect 3237 529 3238 535
rect 1642 495 1643 501
rect 1649 495 1674 501
rect 96 485 97 491
rect 103 490 1655 491
rect 103 486 111 490
rect 115 486 135 490
rect 139 486 175 490
rect 179 486 231 490
rect 235 486 303 490
rect 307 486 359 490
rect 363 486 423 490
rect 427 486 503 490
rect 507 486 543 490
rect 547 486 655 490
rect 659 486 663 490
rect 667 486 775 490
rect 779 486 815 490
rect 819 486 887 490
rect 891 486 975 490
rect 979 486 1007 490
rect 1011 486 1135 490
rect 1139 486 1295 490
rect 1299 486 1455 490
rect 1459 486 1599 490
rect 1603 486 1631 490
rect 1635 486 1655 490
rect 103 485 1655 486
rect 1661 485 1662 491
rect 1668 487 1674 495
rect 1668 486 3219 487
rect 1668 482 1671 486
rect 1675 482 1695 486
rect 1699 482 1887 486
rect 1891 482 2023 486
rect 2027 482 2103 486
rect 2107 482 2343 486
rect 2347 482 2383 486
rect 2387 482 2599 486
rect 2603 482 2743 486
rect 2747 482 2863 486
rect 2867 482 3111 486
rect 3115 482 3135 486
rect 3139 482 3191 486
rect 3195 482 3219 486
rect 1668 481 3219 482
rect 3225 481 3226 487
rect 84 433 85 439
rect 91 438 1643 439
rect 91 434 111 438
rect 115 434 135 438
rect 139 434 231 438
rect 235 434 359 438
rect 363 434 503 438
rect 507 434 655 438
rect 659 434 727 438
rect 731 434 815 438
rect 819 434 855 438
rect 859 434 975 438
rect 979 434 983 438
rect 987 434 1103 438
rect 1107 434 1135 438
rect 1139 434 1223 438
rect 1227 434 1295 438
rect 1299 434 1335 438
rect 1339 434 1447 438
rect 1451 434 1455 438
rect 1459 434 1567 438
rect 1571 434 1599 438
rect 1603 434 1631 438
rect 1635 434 1643 438
rect 91 433 1643 434
rect 1649 433 1650 439
rect 1654 437 1655 443
rect 1661 442 3231 443
rect 1661 438 1671 442
rect 1675 438 1695 442
rect 1699 438 2023 442
rect 2027 438 2247 442
rect 2251 438 2375 442
rect 2379 438 2383 442
rect 2387 438 2503 442
rect 2507 438 2623 442
rect 2627 438 2743 442
rect 2747 438 2855 442
rect 2859 438 2967 442
rect 2971 438 3087 442
rect 3091 438 3111 442
rect 3115 438 3191 442
rect 3195 438 3231 442
rect 1661 437 3231 438
rect 3237 437 3238 443
rect 1642 395 1643 401
rect 1649 395 1674 401
rect 1668 391 1674 395
rect 96 385 97 391
rect 103 390 1655 391
rect 103 386 111 390
rect 115 386 647 390
rect 651 386 727 390
rect 731 386 807 390
rect 811 386 855 390
rect 859 386 951 390
rect 955 386 983 390
rect 987 386 1087 390
rect 1091 386 1103 390
rect 1107 386 1215 390
rect 1219 386 1223 390
rect 1227 386 1335 390
rect 1339 386 1447 390
rect 1451 386 1463 390
rect 1467 386 1567 390
rect 1571 386 1631 390
rect 1635 386 1655 390
rect 103 385 1655 386
rect 1661 385 1662 391
rect 1668 390 3219 391
rect 1668 386 1671 390
rect 1675 386 2151 390
rect 2155 386 2247 390
rect 2251 386 2279 390
rect 2283 386 2375 390
rect 2379 386 2407 390
rect 2411 386 2503 390
rect 2507 386 2535 390
rect 2539 386 2623 390
rect 2627 386 2663 390
rect 2667 386 2743 390
rect 2747 386 2791 390
rect 2795 386 2855 390
rect 2859 386 2919 390
rect 2923 386 2967 390
rect 2971 386 3047 390
rect 3051 386 3087 390
rect 3091 386 3159 390
rect 3163 386 3191 390
rect 3195 386 3219 390
rect 1668 385 3219 386
rect 3225 385 3226 391
rect 84 341 85 347
rect 91 346 1643 347
rect 91 342 111 346
rect 115 342 543 346
rect 547 342 647 346
rect 651 342 671 346
rect 675 342 807 346
rect 811 342 943 346
rect 947 342 951 346
rect 955 342 1079 346
rect 1083 342 1087 346
rect 1091 342 1215 346
rect 1219 342 1223 346
rect 1227 342 1335 346
rect 1339 342 1367 346
rect 1371 342 1463 346
rect 1467 342 1631 346
rect 1635 342 1643 346
rect 91 341 1643 342
rect 1649 341 1650 347
rect 1654 333 1655 339
rect 1661 338 3231 339
rect 1661 334 1671 338
rect 1675 334 2047 338
rect 2051 334 2151 338
rect 2155 334 2175 338
rect 2179 334 2279 338
rect 2283 334 2303 338
rect 2307 334 2407 338
rect 2411 334 2431 338
rect 2435 334 2535 338
rect 2539 334 2567 338
rect 2571 334 2663 338
rect 2667 334 2711 338
rect 2715 334 2791 338
rect 2795 334 2863 338
rect 2867 334 2919 338
rect 2923 334 3023 338
rect 3027 334 3047 338
rect 3051 334 3159 338
rect 3163 334 3191 338
rect 3195 334 3231 338
rect 1661 333 3231 334
rect 3237 333 3238 339
rect 96 297 97 303
rect 103 302 1655 303
rect 103 298 111 302
rect 115 298 463 302
rect 467 298 543 302
rect 547 298 623 302
rect 627 298 671 302
rect 675 298 767 302
rect 771 298 807 302
rect 811 298 903 302
rect 907 298 943 302
rect 947 298 1031 302
rect 1035 298 1079 302
rect 1083 298 1159 302
rect 1163 298 1223 302
rect 1227 298 1287 302
rect 1291 298 1367 302
rect 1371 298 1631 302
rect 1635 298 1655 302
rect 103 297 1655 298
rect 1661 297 1662 303
rect 1642 285 1643 291
rect 1649 290 3219 291
rect 1649 286 1671 290
rect 1675 286 1943 290
rect 1947 286 2047 290
rect 2051 286 2071 290
rect 2075 286 2175 290
rect 2179 286 2199 290
rect 2203 286 2303 290
rect 2307 286 2319 290
rect 2323 286 2431 290
rect 2435 286 2439 290
rect 2443 286 2551 290
rect 2555 286 2567 290
rect 2571 286 2663 290
rect 2667 286 2711 290
rect 2715 286 2783 290
rect 2787 286 2863 290
rect 2867 286 3023 290
rect 3027 286 3159 290
rect 3163 286 3191 290
rect 3195 286 3219 290
rect 1649 285 3219 286
rect 3225 285 3226 291
rect 84 253 85 259
rect 91 258 1643 259
rect 91 254 111 258
rect 115 254 359 258
rect 363 254 463 258
rect 467 254 487 258
rect 491 254 623 258
rect 627 254 759 258
rect 763 254 767 258
rect 771 254 895 258
rect 899 254 903 258
rect 907 254 1031 258
rect 1035 254 1039 258
rect 1043 254 1159 258
rect 1163 254 1183 258
rect 1187 254 1287 258
rect 1291 254 1631 258
rect 1635 254 1643 258
rect 91 253 1643 254
rect 1649 253 1650 259
rect 1654 233 1655 239
rect 1661 238 3231 239
rect 1661 234 1671 238
rect 1675 234 1847 238
rect 1851 234 1943 238
rect 1947 234 1975 238
rect 1979 234 2071 238
rect 2075 234 2103 238
rect 2107 234 2199 238
rect 2203 234 2247 238
rect 2251 234 2319 238
rect 2323 234 2407 238
rect 2411 234 2439 238
rect 2443 234 2551 238
rect 2555 234 2583 238
rect 2587 234 2663 238
rect 2667 234 2767 238
rect 2771 234 2783 238
rect 2787 234 2967 238
rect 2971 234 3159 238
rect 3163 234 3191 238
rect 3195 234 3231 238
rect 1661 233 3231 234
rect 3237 233 3238 239
rect 96 209 97 215
rect 103 214 1655 215
rect 103 210 111 214
rect 115 210 279 214
rect 283 210 359 214
rect 363 210 447 214
rect 451 210 487 214
rect 491 210 615 214
rect 619 210 623 214
rect 627 210 759 214
rect 763 210 775 214
rect 779 210 895 214
rect 899 210 943 214
rect 947 210 1039 214
rect 1043 210 1111 214
rect 1115 210 1183 214
rect 1187 210 1631 214
rect 1635 210 1655 214
rect 103 209 1655 210
rect 1661 209 1662 215
rect 1642 181 1643 187
rect 1649 186 3219 187
rect 1649 182 1671 186
rect 1675 182 1743 186
rect 1747 182 1847 186
rect 1851 182 1871 186
rect 1875 182 1975 186
rect 1979 182 1999 186
rect 2003 182 2103 186
rect 2107 182 2143 186
rect 2147 182 2247 186
rect 2251 182 2311 186
rect 2315 182 2407 186
rect 2411 182 2495 186
rect 2499 182 2583 186
rect 2587 182 2703 186
rect 2707 182 2767 186
rect 2771 182 2919 186
rect 2923 182 2967 186
rect 2971 182 3135 186
rect 3139 182 3159 186
rect 3163 182 3191 186
rect 3195 182 3219 186
rect 1649 181 3219 182
rect 3225 181 3226 187
rect 84 169 85 175
rect 91 174 1643 175
rect 91 170 111 174
rect 115 170 199 174
rect 203 170 279 174
rect 283 170 367 174
rect 371 170 447 174
rect 451 170 535 174
rect 539 170 615 174
rect 619 170 695 174
rect 699 170 775 174
rect 779 170 863 174
rect 867 170 943 174
rect 947 170 1031 174
rect 1035 170 1111 174
rect 1115 170 1631 174
rect 1635 170 1643 174
rect 91 169 1643 170
rect 1649 169 1650 175
rect 1654 125 1655 131
rect 1661 130 3231 131
rect 1661 126 1671 130
rect 1675 126 1695 130
rect 1699 126 1743 130
rect 1747 126 1815 130
rect 1819 126 1871 130
rect 1875 126 1943 130
rect 1947 126 1999 130
rect 2003 126 2071 130
rect 2075 126 2143 130
rect 2147 126 2199 130
rect 2203 126 2311 130
rect 2315 126 2351 130
rect 2355 126 2495 130
rect 2499 126 2519 130
rect 2523 126 2703 130
rect 2707 126 2711 130
rect 2715 126 2911 130
rect 2915 126 2919 130
rect 2923 126 3111 130
rect 3115 126 3135 130
rect 3139 126 3191 130
rect 3195 126 3231 130
rect 1661 125 3231 126
rect 3237 125 3238 131
rect 1654 123 1662 125
rect 96 117 97 123
rect 103 122 1655 123
rect 103 118 111 122
rect 115 118 135 122
rect 139 118 191 122
rect 195 118 199 122
rect 203 118 287 122
rect 291 118 367 122
rect 371 118 383 122
rect 387 118 479 122
rect 483 118 535 122
rect 539 118 583 122
rect 587 118 695 122
rect 699 118 815 122
rect 819 118 863 122
rect 867 118 943 122
rect 947 118 1031 122
rect 1035 118 1079 122
rect 1083 118 1215 122
rect 1219 118 1351 122
rect 1355 118 1487 122
rect 1491 118 1599 122
rect 1603 118 1631 122
rect 1635 118 1655 122
rect 103 117 1655 118
rect 1661 117 1662 123
rect 1642 85 1643 91
rect 1649 90 3219 91
rect 1649 86 1671 90
rect 1675 86 1695 90
rect 1699 86 1815 90
rect 1819 86 1943 90
rect 1947 86 2071 90
rect 2075 86 2199 90
rect 2203 86 2351 90
rect 2355 86 2519 90
rect 2523 86 2711 90
rect 2715 86 2911 90
rect 2915 86 3111 90
rect 3115 86 3191 90
rect 3195 86 3219 90
rect 1649 85 3219 86
rect 3225 85 3226 91
rect 1642 83 1650 85
rect 84 77 85 83
rect 91 82 1643 83
rect 91 78 111 82
rect 115 78 135 82
rect 139 78 191 82
rect 195 78 287 82
rect 291 78 383 82
rect 387 78 479 82
rect 483 78 583 82
rect 587 78 695 82
rect 699 78 815 82
rect 819 78 943 82
rect 947 78 1079 82
rect 1083 78 1215 82
rect 1219 78 1351 82
rect 1355 78 1487 82
rect 1491 78 1599 82
rect 1603 78 1631 82
rect 1635 78 1643 82
rect 91 77 1643 78
rect 1649 77 1650 83
<< m5c >>
rect 1655 3305 1661 3311
rect 3231 3305 3237 3311
rect 1643 3265 1649 3271
rect 3219 3265 3225 3271
rect 1655 3225 1661 3231
rect 3231 3225 3237 3231
rect 1643 3185 1649 3191
rect 3219 3185 3225 3191
rect 1655 3145 1661 3151
rect 3231 3145 3237 3151
rect 85 3125 91 3131
rect 1643 3125 1649 3131
rect 1643 3105 1649 3111
rect 3219 3105 3225 3111
rect 97 3081 103 3087
rect 1655 3081 1661 3087
rect 1655 3065 1661 3071
rect 3231 3065 3237 3071
rect 85 3033 91 3039
rect 1643 3033 1649 3039
rect 1643 3025 1649 3031
rect 3219 3025 3225 3031
rect 97 2989 103 2995
rect 1655 2989 1661 2995
rect 85 2941 91 2947
rect 1643 2941 1649 2947
rect 97 2901 103 2907
rect 1655 2901 1661 2907
rect 1643 2865 1649 2871
rect 3219 2865 3225 2871
rect 85 2853 91 2859
rect 1643 2853 1649 2859
rect 1655 2817 1661 2823
rect 3231 2817 3237 2823
rect 97 2805 103 2811
rect 1655 2805 1661 2811
rect 1643 2777 1649 2783
rect 3219 2777 3225 2783
rect 85 2753 91 2759
rect 1643 2753 1649 2759
rect 1655 2733 1661 2739
rect 3231 2733 3237 2739
rect 97 2701 103 2707
rect 1655 2701 1661 2707
rect 1643 2685 1649 2691
rect 3219 2685 3225 2691
rect 85 2653 91 2659
rect 1643 2653 1649 2659
rect 1655 2645 1661 2651
rect 3231 2645 3237 2651
rect 1643 2611 1649 2617
rect 97 2601 103 2607
rect 1655 2601 1661 2607
rect 3219 2605 3225 2611
rect 1655 2561 1661 2567
rect 3231 2561 3237 2567
rect 85 2549 91 2555
rect 1643 2549 1649 2555
rect 1643 2517 1649 2523
rect 3219 2517 3225 2523
rect 97 2497 103 2503
rect 1655 2497 1661 2503
rect 1655 2469 1661 2475
rect 3231 2469 3237 2475
rect 85 2453 91 2459
rect 1643 2453 1649 2459
rect 1643 2429 1649 2435
rect 3219 2429 3225 2435
rect 97 2397 103 2403
rect 1655 2397 1661 2403
rect 1655 2381 1661 2387
rect 3231 2381 3237 2387
rect 85 2349 91 2355
rect 1643 2349 1649 2355
rect 1643 2341 1649 2347
rect 3219 2341 3225 2347
rect 97 2297 103 2303
rect 1655 2297 1661 2303
rect 1643 2257 1649 2263
rect 3219 2257 3225 2263
rect 85 2245 91 2251
rect 1643 2245 1649 2251
rect 1655 2213 1661 2219
rect 3231 2213 3237 2219
rect 97 2197 103 2203
rect 1655 2197 1661 2203
rect 1643 2173 1649 2179
rect 3219 2173 3225 2179
rect 85 2145 91 2151
rect 1643 2145 1649 2151
rect 1655 2129 1661 2135
rect 3231 2129 3237 2135
rect 1643 2103 1649 2109
rect 97 2093 103 2099
rect 1655 2093 1661 2099
rect 3219 2089 3225 2095
rect 85 2045 91 2051
rect 1643 2045 1649 2051
rect 1655 2049 1661 2055
rect 3231 2049 3237 2055
rect 1643 2015 1649 2021
rect 97 2005 103 2011
rect 1655 2005 1661 2011
rect 3219 2001 3225 2007
rect 85 1957 91 1963
rect 1643 1957 1649 1963
rect 1655 1961 1661 1967
rect 3231 1961 3237 1967
rect 1643 1917 1649 1923
rect 3219 1917 3225 1923
rect 97 1905 103 1911
rect 1655 1905 1661 1911
rect 1655 1873 1661 1879
rect 3231 1873 3237 1879
rect 85 1853 91 1859
rect 1643 1853 1649 1859
rect 1643 1833 1649 1839
rect 3219 1833 3225 1839
rect 97 1805 103 1811
rect 1655 1805 1661 1811
rect 1655 1793 1661 1799
rect 3231 1793 3237 1799
rect 85 1753 91 1759
rect 1643 1753 1649 1759
rect 1643 1745 1649 1751
rect 3219 1745 3225 1751
rect 97 1701 103 1707
rect 1655 1701 1661 1707
rect 1643 1665 1649 1671
rect 3219 1665 3225 1671
rect 85 1649 91 1655
rect 1643 1649 1649 1655
rect 1655 1621 1661 1627
rect 3231 1621 3237 1627
rect 97 1601 103 1607
rect 1655 1601 1661 1607
rect 1643 1581 1649 1587
rect 3219 1581 3225 1587
rect 85 1549 91 1555
rect 1643 1549 1649 1555
rect 1655 1533 1661 1539
rect 3231 1533 3237 1539
rect 97 1501 103 1507
rect 1655 1501 1661 1507
rect 1643 1489 1649 1495
rect 3219 1489 3225 1495
rect 85 1449 91 1455
rect 1643 1449 1649 1455
rect 1655 1445 1661 1451
rect 3231 1445 3237 1451
rect 1643 1407 1649 1413
rect 97 1397 103 1403
rect 1655 1397 1661 1403
rect 3219 1389 3225 1395
rect 85 1349 91 1355
rect 1643 1349 1649 1355
rect 1655 1337 1661 1343
rect 3231 1337 3237 1343
rect 1643 1307 1649 1313
rect 97 1297 103 1303
rect 1655 1297 1661 1303
rect 3219 1289 3225 1295
rect 85 1245 91 1251
rect 1643 1245 1649 1251
rect 1655 1233 1661 1239
rect 3231 1233 3237 1239
rect 1643 1207 1649 1213
rect 97 1197 103 1203
rect 1655 1197 1661 1203
rect 3219 1189 3225 1195
rect 85 1145 91 1151
rect 1643 1145 1649 1151
rect 1655 1149 1661 1155
rect 3231 1149 3237 1155
rect 1643 1105 1649 1111
rect 3219 1105 3225 1111
rect 97 1093 103 1099
rect 1655 1093 1661 1099
rect 1655 1053 1661 1059
rect 3231 1053 3237 1059
rect 85 1045 91 1051
rect 1643 1045 1649 1051
rect 1643 1009 1649 1015
rect 3219 1009 3225 1015
rect 97 993 103 999
rect 1655 993 1661 999
rect 1655 969 1661 975
rect 3231 969 3237 975
rect 85 941 91 947
rect 1643 941 1649 947
rect 1643 921 1649 927
rect 3219 921 3225 927
rect 97 889 103 895
rect 1655 889 1661 895
rect 1655 881 1661 887
rect 3231 881 3237 887
rect 85 845 91 851
rect 1643 845 1649 851
rect 1643 829 1649 835
rect 3219 829 3225 835
rect 97 789 103 795
rect 1655 789 1661 795
rect 85 741 91 747
rect 1643 741 1649 747
rect 1655 701 1661 707
rect 3231 701 3237 707
rect 97 689 103 695
rect 1655 689 1661 695
rect 1643 653 1649 659
rect 3219 653 3225 659
rect 85 637 91 643
rect 1643 637 1649 643
rect 1655 609 1661 615
rect 3231 609 3237 615
rect 97 589 103 595
rect 1655 589 1661 595
rect 1643 569 1649 575
rect 3219 569 3225 575
rect 85 537 91 543
rect 1643 537 1649 543
rect 1655 529 1661 535
rect 3231 529 3237 535
rect 1643 495 1649 501
rect 97 485 103 491
rect 1655 485 1661 491
rect 3219 481 3225 487
rect 85 433 91 439
rect 1643 433 1649 439
rect 1655 437 1661 443
rect 3231 437 3237 443
rect 1643 395 1649 401
rect 97 385 103 391
rect 1655 385 1661 391
rect 3219 385 3225 391
rect 85 341 91 347
rect 1643 341 1649 347
rect 1655 333 1661 339
rect 3231 333 3237 339
rect 97 297 103 303
rect 1655 297 1661 303
rect 1643 285 1649 291
rect 3219 285 3225 291
rect 85 253 91 259
rect 1643 253 1649 259
rect 1655 233 1661 239
rect 3231 233 3237 239
rect 97 209 103 215
rect 1655 209 1661 215
rect 1643 181 1649 187
rect 3219 181 3225 187
rect 85 169 91 175
rect 1643 169 1649 175
rect 1655 125 1661 131
rect 3231 125 3237 131
rect 97 117 103 123
rect 1655 117 1661 123
rect 1643 85 1649 91
rect 3219 85 3225 91
rect 85 77 91 83
rect 1643 77 1649 83
<< m5 >>
rect 84 3131 92 3312
rect 84 3125 85 3131
rect 91 3125 92 3131
rect 84 3039 92 3125
rect 84 3033 85 3039
rect 91 3033 92 3039
rect 84 2947 92 3033
rect 84 2941 85 2947
rect 91 2941 92 2947
rect 84 2859 92 2941
rect 84 2853 85 2859
rect 91 2853 92 2859
rect 84 2759 92 2853
rect 84 2753 85 2759
rect 91 2753 92 2759
rect 84 2659 92 2753
rect 84 2653 85 2659
rect 91 2653 92 2659
rect 84 2555 92 2653
rect 84 2549 85 2555
rect 91 2549 92 2555
rect 84 2459 92 2549
rect 84 2453 85 2459
rect 91 2453 92 2459
rect 84 2355 92 2453
rect 84 2349 85 2355
rect 91 2349 92 2355
rect 84 2251 92 2349
rect 84 2245 85 2251
rect 91 2245 92 2251
rect 84 2151 92 2245
rect 84 2145 85 2151
rect 91 2145 92 2151
rect 84 2051 92 2145
rect 84 2045 85 2051
rect 91 2045 92 2051
rect 84 1963 92 2045
rect 84 1957 85 1963
rect 91 1957 92 1963
rect 84 1859 92 1957
rect 84 1853 85 1859
rect 91 1853 92 1859
rect 84 1759 92 1853
rect 84 1753 85 1759
rect 91 1753 92 1759
rect 84 1655 92 1753
rect 84 1649 85 1655
rect 91 1649 92 1655
rect 84 1555 92 1649
rect 84 1549 85 1555
rect 91 1549 92 1555
rect 84 1455 92 1549
rect 84 1449 85 1455
rect 91 1449 92 1455
rect 84 1355 92 1449
rect 84 1349 85 1355
rect 91 1349 92 1355
rect 84 1251 92 1349
rect 84 1245 85 1251
rect 91 1245 92 1251
rect 84 1151 92 1245
rect 84 1145 85 1151
rect 91 1145 92 1151
rect 84 1051 92 1145
rect 84 1045 85 1051
rect 91 1045 92 1051
rect 84 947 92 1045
rect 84 941 85 947
rect 91 941 92 947
rect 84 851 92 941
rect 84 845 85 851
rect 91 845 92 851
rect 84 747 92 845
rect 84 741 85 747
rect 91 741 92 747
rect 84 643 92 741
rect 84 637 85 643
rect 91 637 92 643
rect 84 543 92 637
rect 84 537 85 543
rect 91 537 92 543
rect 84 439 92 537
rect 84 433 85 439
rect 91 433 92 439
rect 84 347 92 433
rect 84 341 85 347
rect 91 341 92 347
rect 84 259 92 341
rect 84 253 85 259
rect 91 253 92 259
rect 84 175 92 253
rect 84 169 85 175
rect 91 169 92 175
rect 84 83 92 169
rect 84 77 85 83
rect 91 77 92 83
rect 84 72 92 77
rect 96 3087 104 3312
rect 96 3081 97 3087
rect 103 3081 104 3087
rect 96 2995 104 3081
rect 96 2989 97 2995
rect 103 2989 104 2995
rect 96 2907 104 2989
rect 96 2901 97 2907
rect 103 2901 104 2907
rect 96 2811 104 2901
rect 96 2805 97 2811
rect 103 2805 104 2811
rect 96 2707 104 2805
rect 96 2701 97 2707
rect 103 2701 104 2707
rect 96 2607 104 2701
rect 96 2601 97 2607
rect 103 2601 104 2607
rect 96 2503 104 2601
rect 96 2497 97 2503
rect 103 2497 104 2503
rect 96 2403 104 2497
rect 96 2397 97 2403
rect 103 2397 104 2403
rect 96 2303 104 2397
rect 96 2297 97 2303
rect 103 2297 104 2303
rect 96 2203 104 2297
rect 96 2197 97 2203
rect 103 2197 104 2203
rect 96 2099 104 2197
rect 96 2093 97 2099
rect 103 2093 104 2099
rect 96 2011 104 2093
rect 96 2005 97 2011
rect 103 2005 104 2011
rect 96 1911 104 2005
rect 96 1905 97 1911
rect 103 1905 104 1911
rect 96 1811 104 1905
rect 96 1805 97 1811
rect 103 1805 104 1811
rect 96 1707 104 1805
rect 96 1701 97 1707
rect 103 1701 104 1707
rect 96 1607 104 1701
rect 96 1601 97 1607
rect 103 1601 104 1607
rect 96 1507 104 1601
rect 96 1501 97 1507
rect 103 1501 104 1507
rect 96 1403 104 1501
rect 96 1397 97 1403
rect 103 1397 104 1403
rect 96 1303 104 1397
rect 96 1297 97 1303
rect 103 1297 104 1303
rect 96 1203 104 1297
rect 96 1197 97 1203
rect 103 1197 104 1203
rect 96 1099 104 1197
rect 96 1093 97 1099
rect 103 1093 104 1099
rect 96 999 104 1093
rect 96 993 97 999
rect 103 993 104 999
rect 96 895 104 993
rect 96 889 97 895
rect 103 889 104 895
rect 96 795 104 889
rect 96 789 97 795
rect 103 789 104 795
rect 96 695 104 789
rect 96 689 97 695
rect 103 689 104 695
rect 96 595 104 689
rect 96 589 97 595
rect 103 589 104 595
rect 96 491 104 589
rect 96 485 97 491
rect 103 485 104 491
rect 96 391 104 485
rect 96 385 97 391
rect 103 385 104 391
rect 96 303 104 385
rect 96 297 97 303
rect 103 297 104 303
rect 96 215 104 297
rect 96 209 97 215
rect 103 209 104 215
rect 96 123 104 209
rect 96 117 97 123
rect 103 117 104 123
rect 96 72 104 117
rect 1642 3271 1650 3312
rect 1642 3265 1643 3271
rect 1649 3265 1650 3271
rect 1642 3191 1650 3265
rect 1642 3185 1643 3191
rect 1649 3185 1650 3191
rect 1642 3131 1650 3185
rect 1642 3125 1643 3131
rect 1649 3125 1650 3131
rect 1642 3111 1650 3125
rect 1642 3105 1643 3111
rect 1649 3105 1650 3111
rect 1642 3039 1650 3105
rect 1642 3033 1643 3039
rect 1649 3033 1650 3039
rect 1642 3031 1650 3033
rect 1642 3025 1643 3031
rect 1649 3025 1650 3031
rect 1642 2947 1650 3025
rect 1642 2941 1643 2947
rect 1649 2941 1650 2947
rect 1642 2871 1650 2941
rect 1642 2865 1643 2871
rect 1649 2865 1650 2871
rect 1642 2859 1650 2865
rect 1642 2853 1643 2859
rect 1649 2853 1650 2859
rect 1642 2783 1650 2853
rect 1642 2777 1643 2783
rect 1649 2777 1650 2783
rect 1642 2759 1650 2777
rect 1642 2753 1643 2759
rect 1649 2753 1650 2759
rect 1642 2691 1650 2753
rect 1642 2685 1643 2691
rect 1649 2685 1650 2691
rect 1642 2659 1650 2685
rect 1642 2653 1643 2659
rect 1649 2653 1650 2659
rect 1642 2617 1650 2653
rect 1642 2611 1643 2617
rect 1649 2611 1650 2617
rect 1642 2555 1650 2611
rect 1642 2549 1643 2555
rect 1649 2549 1650 2555
rect 1642 2523 1650 2549
rect 1642 2517 1643 2523
rect 1649 2517 1650 2523
rect 1642 2459 1650 2517
rect 1642 2453 1643 2459
rect 1649 2453 1650 2459
rect 1642 2435 1650 2453
rect 1642 2429 1643 2435
rect 1649 2429 1650 2435
rect 1642 2355 1650 2429
rect 1642 2349 1643 2355
rect 1649 2349 1650 2355
rect 1642 2347 1650 2349
rect 1642 2341 1643 2347
rect 1649 2341 1650 2347
rect 1642 2263 1650 2341
rect 1642 2257 1643 2263
rect 1649 2257 1650 2263
rect 1642 2251 1650 2257
rect 1642 2245 1643 2251
rect 1649 2245 1650 2251
rect 1642 2179 1650 2245
rect 1642 2173 1643 2179
rect 1649 2173 1650 2179
rect 1642 2151 1650 2173
rect 1642 2145 1643 2151
rect 1649 2145 1650 2151
rect 1642 2109 1650 2145
rect 1642 2103 1643 2109
rect 1649 2103 1650 2109
rect 1642 2051 1650 2103
rect 1642 2045 1643 2051
rect 1649 2045 1650 2051
rect 1642 2021 1650 2045
rect 1642 2015 1643 2021
rect 1649 2015 1650 2021
rect 1642 1963 1650 2015
rect 1642 1957 1643 1963
rect 1649 1957 1650 1963
rect 1642 1923 1650 1957
rect 1642 1917 1643 1923
rect 1649 1917 1650 1923
rect 1642 1859 1650 1917
rect 1642 1853 1643 1859
rect 1649 1853 1650 1859
rect 1642 1839 1650 1853
rect 1642 1833 1643 1839
rect 1649 1833 1650 1839
rect 1642 1759 1650 1833
rect 1642 1753 1643 1759
rect 1649 1753 1650 1759
rect 1642 1751 1650 1753
rect 1642 1745 1643 1751
rect 1649 1745 1650 1751
rect 1642 1671 1650 1745
rect 1642 1665 1643 1671
rect 1649 1665 1650 1671
rect 1642 1655 1650 1665
rect 1642 1649 1643 1655
rect 1649 1649 1650 1655
rect 1642 1587 1650 1649
rect 1642 1581 1643 1587
rect 1649 1581 1650 1587
rect 1642 1555 1650 1581
rect 1642 1549 1643 1555
rect 1649 1549 1650 1555
rect 1642 1495 1650 1549
rect 1642 1489 1643 1495
rect 1649 1489 1650 1495
rect 1642 1455 1650 1489
rect 1642 1449 1643 1455
rect 1649 1449 1650 1455
rect 1642 1413 1650 1449
rect 1642 1407 1643 1413
rect 1649 1407 1650 1413
rect 1642 1355 1650 1407
rect 1642 1349 1643 1355
rect 1649 1349 1650 1355
rect 1642 1313 1650 1349
rect 1642 1307 1643 1313
rect 1649 1307 1650 1313
rect 1642 1251 1650 1307
rect 1642 1245 1643 1251
rect 1649 1245 1650 1251
rect 1642 1213 1650 1245
rect 1642 1207 1643 1213
rect 1649 1207 1650 1213
rect 1642 1151 1650 1207
rect 1642 1145 1643 1151
rect 1649 1145 1650 1151
rect 1642 1111 1650 1145
rect 1642 1105 1643 1111
rect 1649 1105 1650 1111
rect 1642 1051 1650 1105
rect 1642 1045 1643 1051
rect 1649 1045 1650 1051
rect 1642 1015 1650 1045
rect 1642 1009 1643 1015
rect 1649 1009 1650 1015
rect 1642 947 1650 1009
rect 1642 941 1643 947
rect 1649 941 1650 947
rect 1642 927 1650 941
rect 1642 921 1643 927
rect 1649 921 1650 927
rect 1642 851 1650 921
rect 1642 845 1643 851
rect 1649 845 1650 851
rect 1642 835 1650 845
rect 1642 829 1643 835
rect 1649 829 1650 835
rect 1642 747 1650 829
rect 1642 741 1643 747
rect 1649 741 1650 747
rect 1642 659 1650 741
rect 1642 653 1643 659
rect 1649 653 1650 659
rect 1642 643 1650 653
rect 1642 637 1643 643
rect 1649 637 1650 643
rect 1642 575 1650 637
rect 1642 569 1643 575
rect 1649 569 1650 575
rect 1642 543 1650 569
rect 1642 537 1643 543
rect 1649 537 1650 543
rect 1642 501 1650 537
rect 1642 495 1643 501
rect 1649 495 1650 501
rect 1642 439 1650 495
rect 1642 433 1643 439
rect 1649 433 1650 439
rect 1642 401 1650 433
rect 1642 395 1643 401
rect 1649 395 1650 401
rect 1642 347 1650 395
rect 1642 341 1643 347
rect 1649 341 1650 347
rect 1642 291 1650 341
rect 1642 285 1643 291
rect 1649 285 1650 291
rect 1642 259 1650 285
rect 1642 253 1643 259
rect 1649 253 1650 259
rect 1642 187 1650 253
rect 1642 181 1643 187
rect 1649 181 1650 187
rect 1642 175 1650 181
rect 1642 169 1643 175
rect 1649 169 1650 175
rect 1642 91 1650 169
rect 1642 85 1643 91
rect 1649 85 1650 91
rect 1642 83 1650 85
rect 1642 77 1643 83
rect 1649 77 1650 83
rect 1642 72 1650 77
rect 1654 3311 1662 3312
rect 1654 3305 1655 3311
rect 1661 3305 1662 3311
rect 1654 3231 1662 3305
rect 1654 3225 1655 3231
rect 1661 3225 1662 3231
rect 1654 3151 1662 3225
rect 1654 3145 1655 3151
rect 1661 3145 1662 3151
rect 1654 3087 1662 3145
rect 1654 3081 1655 3087
rect 1661 3081 1662 3087
rect 1654 3071 1662 3081
rect 1654 3065 1655 3071
rect 1661 3065 1662 3071
rect 1654 2995 1662 3065
rect 1654 2989 1655 2995
rect 1661 2989 1662 2995
rect 1654 2907 1662 2989
rect 1654 2901 1655 2907
rect 1661 2901 1662 2907
rect 1654 2823 1662 2901
rect 1654 2817 1655 2823
rect 1661 2817 1662 2823
rect 1654 2811 1662 2817
rect 1654 2805 1655 2811
rect 1661 2805 1662 2811
rect 1654 2739 1662 2805
rect 1654 2733 1655 2739
rect 1661 2733 1662 2739
rect 1654 2707 1662 2733
rect 1654 2701 1655 2707
rect 1661 2701 1662 2707
rect 1654 2651 1662 2701
rect 1654 2645 1655 2651
rect 1661 2645 1662 2651
rect 1654 2607 1662 2645
rect 1654 2601 1655 2607
rect 1661 2601 1662 2607
rect 1654 2567 1662 2601
rect 1654 2561 1655 2567
rect 1661 2561 1662 2567
rect 1654 2503 1662 2561
rect 1654 2497 1655 2503
rect 1661 2497 1662 2503
rect 1654 2475 1662 2497
rect 1654 2469 1655 2475
rect 1661 2469 1662 2475
rect 1654 2403 1662 2469
rect 1654 2397 1655 2403
rect 1661 2397 1662 2403
rect 1654 2387 1662 2397
rect 1654 2381 1655 2387
rect 1661 2381 1662 2387
rect 1654 2303 1662 2381
rect 1654 2297 1655 2303
rect 1661 2297 1662 2303
rect 1654 2219 1662 2297
rect 1654 2213 1655 2219
rect 1661 2213 1662 2219
rect 1654 2203 1662 2213
rect 1654 2197 1655 2203
rect 1661 2197 1662 2203
rect 1654 2135 1662 2197
rect 1654 2129 1655 2135
rect 1661 2129 1662 2135
rect 1654 2099 1662 2129
rect 1654 2093 1655 2099
rect 1661 2093 1662 2099
rect 1654 2055 1662 2093
rect 1654 2049 1655 2055
rect 1661 2049 1662 2055
rect 1654 2011 1662 2049
rect 1654 2005 1655 2011
rect 1661 2005 1662 2011
rect 1654 1967 1662 2005
rect 1654 1961 1655 1967
rect 1661 1961 1662 1967
rect 1654 1911 1662 1961
rect 1654 1905 1655 1911
rect 1661 1905 1662 1911
rect 1654 1879 1662 1905
rect 1654 1873 1655 1879
rect 1661 1873 1662 1879
rect 1654 1811 1662 1873
rect 1654 1805 1655 1811
rect 1661 1805 1662 1811
rect 1654 1799 1662 1805
rect 1654 1793 1655 1799
rect 1661 1793 1662 1799
rect 1654 1707 1662 1793
rect 1654 1701 1655 1707
rect 1661 1701 1662 1707
rect 1654 1627 1662 1701
rect 1654 1621 1655 1627
rect 1661 1621 1662 1627
rect 1654 1607 1662 1621
rect 1654 1601 1655 1607
rect 1661 1601 1662 1607
rect 1654 1539 1662 1601
rect 1654 1533 1655 1539
rect 1661 1533 1662 1539
rect 1654 1507 1662 1533
rect 1654 1501 1655 1507
rect 1661 1501 1662 1507
rect 1654 1451 1662 1501
rect 1654 1445 1655 1451
rect 1661 1445 1662 1451
rect 1654 1403 1662 1445
rect 1654 1397 1655 1403
rect 1661 1397 1662 1403
rect 1654 1343 1662 1397
rect 1654 1337 1655 1343
rect 1661 1337 1662 1343
rect 1654 1303 1662 1337
rect 1654 1297 1655 1303
rect 1661 1297 1662 1303
rect 1654 1239 1662 1297
rect 1654 1233 1655 1239
rect 1661 1233 1662 1239
rect 1654 1203 1662 1233
rect 1654 1197 1655 1203
rect 1661 1197 1662 1203
rect 1654 1155 1662 1197
rect 1654 1149 1655 1155
rect 1661 1149 1662 1155
rect 1654 1099 1662 1149
rect 1654 1093 1655 1099
rect 1661 1093 1662 1099
rect 1654 1059 1662 1093
rect 1654 1053 1655 1059
rect 1661 1053 1662 1059
rect 1654 999 1662 1053
rect 1654 993 1655 999
rect 1661 993 1662 999
rect 1654 975 1662 993
rect 1654 969 1655 975
rect 1661 969 1662 975
rect 1654 895 1662 969
rect 1654 889 1655 895
rect 1661 889 1662 895
rect 1654 887 1662 889
rect 1654 881 1655 887
rect 1661 881 1662 887
rect 1654 795 1662 881
rect 1654 789 1655 795
rect 1661 789 1662 795
rect 1654 707 1662 789
rect 1654 701 1655 707
rect 1661 701 1662 707
rect 1654 695 1662 701
rect 1654 689 1655 695
rect 1661 689 1662 695
rect 1654 615 1662 689
rect 1654 609 1655 615
rect 1661 609 1662 615
rect 1654 595 1662 609
rect 1654 589 1655 595
rect 1661 589 1662 595
rect 1654 535 1662 589
rect 1654 529 1655 535
rect 1661 529 1662 535
rect 1654 491 1662 529
rect 1654 485 1655 491
rect 1661 485 1662 491
rect 1654 443 1662 485
rect 1654 437 1655 443
rect 1661 437 1662 443
rect 1654 391 1662 437
rect 1654 385 1655 391
rect 1661 385 1662 391
rect 1654 339 1662 385
rect 1654 333 1655 339
rect 1661 333 1662 339
rect 1654 303 1662 333
rect 1654 297 1655 303
rect 1661 297 1662 303
rect 1654 239 1662 297
rect 1654 233 1655 239
rect 1661 233 1662 239
rect 1654 215 1662 233
rect 1654 209 1655 215
rect 1661 209 1662 215
rect 1654 131 1662 209
rect 1654 125 1655 131
rect 1661 125 1662 131
rect 1654 123 1662 125
rect 1654 117 1655 123
rect 1661 117 1662 123
rect 1654 72 1662 117
rect 3218 3271 3226 3312
rect 3218 3265 3219 3271
rect 3225 3265 3226 3271
rect 3218 3191 3226 3265
rect 3218 3185 3219 3191
rect 3225 3185 3226 3191
rect 3218 3111 3226 3185
rect 3218 3105 3219 3111
rect 3225 3105 3226 3111
rect 3218 3031 3226 3105
rect 3218 3025 3219 3031
rect 3225 3025 3226 3031
rect 3218 2871 3226 3025
rect 3218 2865 3219 2871
rect 3225 2865 3226 2871
rect 3218 2783 3226 2865
rect 3218 2777 3219 2783
rect 3225 2777 3226 2783
rect 3218 2691 3226 2777
rect 3218 2685 3219 2691
rect 3225 2685 3226 2691
rect 3218 2611 3226 2685
rect 3218 2605 3219 2611
rect 3225 2605 3226 2611
rect 3218 2523 3226 2605
rect 3218 2517 3219 2523
rect 3225 2517 3226 2523
rect 3218 2435 3226 2517
rect 3218 2429 3219 2435
rect 3225 2429 3226 2435
rect 3218 2347 3226 2429
rect 3218 2341 3219 2347
rect 3225 2341 3226 2347
rect 3218 2263 3226 2341
rect 3218 2257 3219 2263
rect 3225 2257 3226 2263
rect 3218 2179 3226 2257
rect 3218 2173 3219 2179
rect 3225 2173 3226 2179
rect 3218 2095 3226 2173
rect 3218 2089 3219 2095
rect 3225 2089 3226 2095
rect 3218 2007 3226 2089
rect 3218 2001 3219 2007
rect 3225 2001 3226 2007
rect 3218 1923 3226 2001
rect 3218 1917 3219 1923
rect 3225 1917 3226 1923
rect 3218 1839 3226 1917
rect 3218 1833 3219 1839
rect 3225 1833 3226 1839
rect 3218 1751 3226 1833
rect 3218 1745 3219 1751
rect 3225 1745 3226 1751
rect 3218 1671 3226 1745
rect 3218 1665 3219 1671
rect 3225 1665 3226 1671
rect 3218 1587 3226 1665
rect 3218 1581 3219 1587
rect 3225 1581 3226 1587
rect 3218 1495 3226 1581
rect 3218 1489 3219 1495
rect 3225 1489 3226 1495
rect 3218 1395 3226 1489
rect 3218 1389 3219 1395
rect 3225 1389 3226 1395
rect 3218 1295 3226 1389
rect 3218 1289 3219 1295
rect 3225 1289 3226 1295
rect 3218 1195 3226 1289
rect 3218 1189 3219 1195
rect 3225 1189 3226 1195
rect 3218 1111 3226 1189
rect 3218 1105 3219 1111
rect 3225 1105 3226 1111
rect 3218 1015 3226 1105
rect 3218 1009 3219 1015
rect 3225 1009 3226 1015
rect 3218 927 3226 1009
rect 3218 921 3219 927
rect 3225 921 3226 927
rect 3218 835 3226 921
rect 3218 829 3219 835
rect 3225 829 3226 835
rect 3218 659 3226 829
rect 3218 653 3219 659
rect 3225 653 3226 659
rect 3218 575 3226 653
rect 3218 569 3219 575
rect 3225 569 3226 575
rect 3218 487 3226 569
rect 3218 481 3219 487
rect 3225 481 3226 487
rect 3218 391 3226 481
rect 3218 385 3219 391
rect 3225 385 3226 391
rect 3218 291 3226 385
rect 3218 285 3219 291
rect 3225 285 3226 291
rect 3218 187 3226 285
rect 3218 181 3219 187
rect 3225 181 3226 187
rect 3218 91 3226 181
rect 3218 85 3219 91
rect 3225 85 3226 91
rect 3218 72 3226 85
rect 3230 3311 3238 3312
rect 3230 3305 3231 3311
rect 3237 3305 3238 3311
rect 3230 3231 3238 3305
rect 3230 3225 3231 3231
rect 3237 3225 3238 3231
rect 3230 3151 3238 3225
rect 3230 3145 3231 3151
rect 3237 3145 3238 3151
rect 3230 3071 3238 3145
rect 3230 3065 3231 3071
rect 3237 3065 3238 3071
rect 3230 2823 3238 3065
rect 3230 2817 3231 2823
rect 3237 2817 3238 2823
rect 3230 2739 3238 2817
rect 3230 2733 3231 2739
rect 3237 2733 3238 2739
rect 3230 2651 3238 2733
rect 3230 2645 3231 2651
rect 3237 2645 3238 2651
rect 3230 2567 3238 2645
rect 3230 2561 3231 2567
rect 3237 2561 3238 2567
rect 3230 2475 3238 2561
rect 3230 2469 3231 2475
rect 3237 2469 3238 2475
rect 3230 2387 3238 2469
rect 3230 2381 3231 2387
rect 3237 2381 3238 2387
rect 3230 2219 3238 2381
rect 3230 2213 3231 2219
rect 3237 2213 3238 2219
rect 3230 2135 3238 2213
rect 3230 2129 3231 2135
rect 3237 2129 3238 2135
rect 3230 2055 3238 2129
rect 3230 2049 3231 2055
rect 3237 2049 3238 2055
rect 3230 1967 3238 2049
rect 3230 1961 3231 1967
rect 3237 1961 3238 1967
rect 3230 1879 3238 1961
rect 3230 1873 3231 1879
rect 3237 1873 3238 1879
rect 3230 1799 3238 1873
rect 3230 1793 3231 1799
rect 3237 1793 3238 1799
rect 3230 1627 3238 1793
rect 3230 1621 3231 1627
rect 3237 1621 3238 1627
rect 3230 1539 3238 1621
rect 3230 1533 3231 1539
rect 3237 1533 3238 1539
rect 3230 1451 3238 1533
rect 3230 1445 3231 1451
rect 3237 1445 3238 1451
rect 3230 1343 3238 1445
rect 3230 1337 3231 1343
rect 3237 1337 3238 1343
rect 3230 1239 3238 1337
rect 3230 1233 3231 1239
rect 3237 1233 3238 1239
rect 3230 1155 3238 1233
rect 3230 1149 3231 1155
rect 3237 1149 3238 1155
rect 3230 1059 3238 1149
rect 3230 1053 3231 1059
rect 3237 1053 3238 1059
rect 3230 975 3238 1053
rect 3230 969 3231 975
rect 3237 969 3238 975
rect 3230 887 3238 969
rect 3230 881 3231 887
rect 3237 881 3238 887
rect 3230 707 3238 881
rect 3230 701 3231 707
rect 3237 701 3238 707
rect 3230 615 3238 701
rect 3230 609 3231 615
rect 3237 609 3238 615
rect 3230 535 3238 609
rect 3230 529 3231 535
rect 3237 529 3238 535
rect 3230 443 3238 529
rect 3230 437 3231 443
rect 3237 437 3238 443
rect 3230 339 3238 437
rect 3230 333 3231 339
rect 3237 333 3238 339
rect 3230 239 3238 333
rect 3230 233 3231 239
rect 3237 233 3238 239
rect 3230 131 3238 233
rect 3230 125 3231 131
rect 3237 125 3238 131
rect 3230 72 3238 125
use _0_0std_0_0cells_0_0TIELOX1  tielo_5672_6
timestamp 1730814361
transform 1 0 128 0 1 80
box 7 3 20 38
use welltap_svt  __well_tap__0
timestamp 1730814361
transform 1 0 104 0 1 84
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0TIELOX1  tielo_5672_6
timestamp 1730814361
transform 1 0 128 0 1 80
box 7 3 20 38
use welltap_svt  __well_tap__0
timestamp 1730814361
transform 1 0 104 0 1 84
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0TIELOX1  tielo_5657_6
timestamp 1730814361
transform 1 0 184 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5657_6
timestamp 1730814361
transform 1 0 184 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5658_6
timestamp 1730814361
transform 1 0 280 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5658_6
timestamp 1730814361
transform 1 0 280 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5659_6
timestamp 1730814361
transform 1 0 376 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5659_6
timestamp 1730814361
transform 1 0 376 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5660_6
timestamp 1730814361
transform 1 0 472 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5660_6
timestamp 1730814361
transform 1 0 472 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5555_6
timestamp 1730814361
transform 1 0 576 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5555_6
timestamp 1730814361
transform 1 0 576 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5556_6
timestamp 1730814361
transform 1 0 688 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5556_6
timestamp 1730814361
transform 1 0 688 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5557_6
timestamp 1730814361
transform 1 0 808 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5557_6
timestamp 1730814361
transform 1 0 808 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5558_6
timestamp 1730814361
transform 1 0 936 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5558_6
timestamp 1730814361
transform 1 0 936 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5559_6
timestamp 1730814361
transform 1 0 1072 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5559_6
timestamp 1730814361
transform 1 0 1072 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5560_6
timestamp 1730814361
transform 1 0 1208 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5560_6
timestamp 1730814361
transform 1 0 1208 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5583_6
timestamp 1730814361
transform 1 0 1344 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5583_6
timestamp 1730814361
transform 1 0 1344 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5584_6
timestamp 1730814361
transform 1 0 1480 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5584_6
timestamp 1730814361
transform 1 0 1480 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5585_6
timestamp 1730814361
transform 1 0 1592 0 1 80
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5585_6
timestamp 1730814361
transform 1 0 1592 0 1 80
box 7 3 20 38
use welltap_svt  __well_tap__1
timestamp 1730814361
transform 1 0 1624 0 1 84
box 8 4 12 24
use welltap_svt  __well_tap__124
timestamp 1730814361
transform 1 0 1664 0 1 92
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730814361
transform 1 0 1624 0 1 84
box 8 4 12 24
use welltap_svt  __well_tap__124
timestamp 1730814361
transform 1 0 1664 0 1 92
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5586_6
timestamp 1730814361
transform 1 0 1688 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5586_6
timestamp 1730814361
transform 1 0 1688 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5587_6
timestamp 1730814361
transform 1 0 1808 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5587_6
timestamp 1730814361
transform 1 0 1808 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5588_6
timestamp 1730814361
transform 1 0 1936 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5588_6
timestamp 1730814361
transform 1 0 1936 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5124_6
timestamp 1730814361
transform 1 0 2064 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5124_6
timestamp 1730814361
transform 1 0 2064 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_579_6
timestamp 1730814361
transform 1 0 2192 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_579_6
timestamp 1730814361
transform 1 0 2192 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_564_6
timestamp 1730814361
transform 1 0 2344 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_564_6
timestamp 1730814361
transform 1 0 2344 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_565_6
timestamp 1730814361
transform 1 0 2512 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_565_6
timestamp 1730814361
transform 1 0 2512 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_566_6
timestamp 1730814361
transform 1 0 2704 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_566_6
timestamp 1730814361
transform 1 0 2704 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_567_6
timestamp 1730814361
transform 1 0 2904 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_567_6
timestamp 1730814361
transform 1 0 2904 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5463_6
timestamp 1730814361
transform 1 0 3104 0 1 88
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5463_6
timestamp 1730814361
transform 1 0 3104 0 1 88
box 7 3 20 38
use welltap_svt  __well_tap__125
timestamp 1730814361
transform 1 0 3184 0 1 92
box 8 4 12 24
use welltap_svt  __well_tap__125
timestamp 1730814361
transform 1 0 3184 0 1 92
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730814361
transform 1 0 104 0 -1 168
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730814361
transform 1 0 104 0 1 176
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730814361
transform 1 0 104 0 -1 168
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730814361
transform 1 0 104 0 1 176
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5661_6
timestamp 1730814361
transform 1 0 192 0 -1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5661_6
timestamp 1730814361
transform 1 0 192 0 -1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5664_6
timestamp 1730814361
transform 1 0 272 0 1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5664_6
timestamp 1730814361
transform 1 0 272 0 1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5662_6
timestamp 1730814361
transform 1 0 360 0 -1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5662_6
timestamp 1730814361
transform 1 0 360 0 -1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5665_6
timestamp 1730814361
transform 1 0 440 0 1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5665_6
timestamp 1730814361
transform 1 0 440 0 1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5663_6
timestamp 1730814361
transform 1 0 528 0 -1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5663_6
timestamp 1730814361
transform 1 0 528 0 -1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5666_6
timestamp 1730814361
transform 1 0 608 0 1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5666_6
timestamp 1730814361
transform 1 0 608 0 1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5561_6
timestamp 1730814361
transform 1 0 688 0 -1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5561_6
timestamp 1730814361
transform 1 0 688 0 -1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5501_6
timestamp 1730814361
transform 1 0 768 0 1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5501_6
timestamp 1730814361
transform 1 0 768 0 1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5562_6
timestamp 1730814361
transform 1 0 856 0 -1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5562_6
timestamp 1730814361
transform 1 0 856 0 -1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5502_6
timestamp 1730814361
transform 1 0 936 0 1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5502_6
timestamp 1730814361
transform 1 0 936 0 1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5516_6
timestamp 1730814361
transform 1 0 1024 0 -1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5516_6
timestamp 1730814361
transform 1 0 1024 0 -1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5503_6
timestamp 1730814361
transform 1 0 1104 0 1 172
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5503_6
timestamp 1730814361
transform 1 0 1104 0 1 172
box 7 3 20 38
use welltap_svt  __well_tap__3
timestamp 1730814361
transform 1 0 1624 0 -1 168
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730814361
transform 1 0 1624 0 1 176
box 8 4 12 24
use welltap_svt  __well_tap__126
timestamp 1730814361
transform 1 0 1664 0 -1 180
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730814361
transform 1 0 1624 0 -1 168
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730814361
transform 1 0 1624 0 1 176
box 8 4 12 24
use welltap_svt  __well_tap__126
timestamp 1730814361
transform 1 0 1664 0 -1 180
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5589_6
timestamp 1730814361
transform 1 0 1736 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5589_6
timestamp 1730814361
transform 1 0 1736 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5590_6
timestamp 1730814361
transform 1 0 1864 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5590_6
timestamp 1730814361
transform 1 0 1864 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5591_6
timestamp 1730814361
transform 1 0 1992 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5591_6
timestamp 1730814361
transform 1 0 1992 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5592_6
timestamp 1730814361
transform 1 0 2136 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5592_6
timestamp 1730814361
transform 1 0 2136 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_568_6
timestamp 1730814361
transform 1 0 2304 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_568_6
timestamp 1730814361
transform 1 0 2304 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_569_6
timestamp 1730814361
transform 1 0 2488 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_569_6
timestamp 1730814361
transform 1 0 2488 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_570_6
timestamp 1730814361
transform 1 0 2696 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_570_6
timestamp 1730814361
transform 1 0 2696 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_571_6
timestamp 1730814361
transform 1 0 2912 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_571_6
timestamp 1730814361
transform 1 0 2912 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5464_6
timestamp 1730814361
transform 1 0 3128 0 -1 184
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5464_6
timestamp 1730814361
transform 1 0 3128 0 -1 184
box 7 3 20 38
use welltap_svt  __well_tap__127
timestamp 1730814361
transform 1 0 3184 0 -1 180
box 8 4 12 24
use welltap_svt  __well_tap__127
timestamp 1730814361
transform 1 0 3184 0 -1 180
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730814361
transform 1 0 104 0 -1 252
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730814361
transform 1 0 104 0 -1 252
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5667_6
timestamp 1730814361
transform 1 0 352 0 -1 256
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5667_6
timestamp 1730814361
transform 1 0 352 0 -1 256
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5668_6
timestamp 1730814361
transform 1 0 480 0 -1 256
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5668_6
timestamp 1730814361
transform 1 0 480 0 -1 256
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5669_6
timestamp 1730814361
transform 1 0 616 0 -1 256
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5669_6
timestamp 1730814361
transform 1 0 616 0 -1 256
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5670_6
timestamp 1730814361
transform 1 0 752 0 -1 256
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5670_6
timestamp 1730814361
transform 1 0 752 0 -1 256
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5504_6
timestamp 1730814361
transform 1 0 888 0 -1 256
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5504_6
timestamp 1730814361
transform 1 0 888 0 -1 256
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5505_6
timestamp 1730814361
transform 1 0 1032 0 -1 256
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5505_6
timestamp 1730814361
transform 1 0 1032 0 -1 256
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5506_6
timestamp 1730814361
transform 1 0 1176 0 -1 256
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5506_6
timestamp 1730814361
transform 1 0 1176 0 -1 256
box 7 3 20 38
use welltap_svt  __well_tap__7
timestamp 1730814361
transform 1 0 1624 0 -1 252
box 8 4 12 24
use welltap_svt  __well_tap__128
timestamp 1730814361
transform 1 0 1664 0 1 200
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730814361
transform 1 0 1624 0 -1 252
box 8 4 12 24
use welltap_svt  __well_tap__128
timestamp 1730814361
transform 1 0 1664 0 1 200
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5593_6
timestamp 1730814361
transform 1 0 1840 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5593_6
timestamp 1730814361
transform 1 0 1840 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5909_6
timestamp 1730814361
transform 1 0 1936 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5922_6
timestamp 1730814361
transform 1 0 1968 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5909_6
timestamp 1730814361
transform 1 0 1936 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5922_6
timestamp 1730814361
transform 1 0 1968 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5907_6
timestamp 1730814361
transform 1 0 2096 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5910_6
timestamp 1730814361
transform 1 0 2064 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5907_6
timestamp 1730814361
transform 1 0 2096 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5910_6
timestamp 1730814361
transform 1 0 2064 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5908_6
timestamp 1730814361
transform 1 0 2240 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5911_6
timestamp 1730814361
transform 1 0 2192 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5908_6
timestamp 1730814361
transform 1 0 2240 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5911_6
timestamp 1730814361
transform 1 0 2192 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5912_6
timestamp 1730814361
transform 1 0 2312 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5912_6
timestamp 1730814361
transform 1 0 2312 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_572_6
timestamp 1730814361
transform 1 0 2400 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_572_6
timestamp 1730814361
transform 1 0 2400 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_576_6
timestamp 1730814361
transform 1 0 2432 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_576_6
timestamp 1730814361
transform 1 0 2432 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_577_6
timestamp 1730814361
transform 1 0 2544 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_577_6
timestamp 1730814361
transform 1 0 2544 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_573_6
timestamp 1730814361
transform 1 0 2576 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_573_6
timestamp 1730814361
transform 1 0 2576 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_578_6
timestamp 1730814361
transform 1 0 2656 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_578_6
timestamp 1730814361
transform 1 0 2656 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_574_6
timestamp 1730814361
transform 1 0 2760 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5250_6
timestamp 1730814361
transform 1 0 2776 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_574_6
timestamp 1730814361
transform 1 0 2760 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5250_6
timestamp 1730814361
transform 1 0 2776 0 -1 288
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_575_6
timestamp 1730814361
transform 1 0 2960 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_575_6
timestamp 1730814361
transform 1 0 2960 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5465_6
timestamp 1730814361
transform 1 0 3152 0 1 196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5465_6
timestamp 1730814361
transform 1 0 3152 0 1 196
box 7 3 20 38
use welltap_svt  __well_tap__129
timestamp 1730814361
transform 1 0 3184 0 1 200
box 8 4 12 24
use welltap_svt  __well_tap__129
timestamp 1730814361
transform 1 0 3184 0 1 200
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730814361
transform 1 0 104 0 1 264
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730814361
transform 1 0 104 0 -1 340
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730814361
transform 1 0 104 0 1 264
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730814361
transform 1 0 104 0 -1 340
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5671_6
timestamp 1730814361
transform 1 0 456 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5671_6
timestamp 1730814361
transform 1 0 456 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5674_6
timestamp 1730814361
transform 1 0 536 0 -1 344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5674_6
timestamp 1730814361
transform 1 0 536 0 -1 344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5656_6
timestamp 1730814361
transform 1 0 616 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5656_6
timestamp 1730814361
transform 1 0 616 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5675_6
timestamp 1730814361
transform 1 0 664 0 -1 344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5675_6
timestamp 1730814361
transform 1 0 664 0 -1 344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5673_6
timestamp 1730814361
transform 1 0 760 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5676_6
timestamp 1730814361
transform 1 0 800 0 -1 344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5673_6
timestamp 1730814361
transform 1 0 760 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5676_6
timestamp 1730814361
transform 1 0 800 0 -1 344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5507_6
timestamp 1730814361
transform 1 0 896 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5677_6
timestamp 1730814361
transform 1 0 936 0 -1 344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5507_6
timestamp 1730814361
transform 1 0 896 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5677_6
timestamp 1730814361
transform 1 0 936 0 -1 344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5508_6
timestamp 1730814361
transform 1 0 1024 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5508_6
timestamp 1730814361
transform 1 0 1024 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5511_6
timestamp 1730814361
transform 1 0 1072 0 -1 344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5511_6
timestamp 1730814361
transform 1 0 1072 0 -1 344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5509_6
timestamp 1730814361
transform 1 0 1152 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5509_6
timestamp 1730814361
transform 1 0 1152 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5512_6
timestamp 1730814361
transform 1 0 1216 0 -1 344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5512_6
timestamp 1730814361
transform 1 0 1216 0 -1 344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5510_6
timestamp 1730814361
transform 1 0 1280 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5510_6
timestamp 1730814361
transform 1 0 1280 0 1 260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5513_6
timestamp 1730814361
transform 1 0 1360 0 -1 344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5513_6
timestamp 1730814361
transform 1 0 1360 0 -1 344
box 7 3 20 38
use welltap_svt  __well_tap__9
timestamp 1730814361
transform 1 0 1624 0 1 264
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730814361
transform 1 0 1624 0 -1 340
box 8 4 12 24
use welltap_svt  __well_tap__130
timestamp 1730814361
transform 1 0 1664 0 -1 284
box 8 4 12 24
use welltap_svt  __well_tap__132
timestamp 1730814361
transform 1 0 1664 0 1 300
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730814361
transform 1 0 1624 0 1 264
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730814361
transform 1 0 1624 0 -1 340
box 8 4 12 24
use welltap_svt  __well_tap__130
timestamp 1730814361
transform 1 0 1664 0 -1 284
box 8 4 12 24
use welltap_svt  __well_tap__132
timestamp 1730814361
transform 1 0 1664 0 1 300
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5913_6
timestamp 1730814361
transform 1 0 2040 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5913_6
timestamp 1730814361
transform 1 0 2040 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5914_6
timestamp 1730814361
transform 1 0 2168 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5914_6
timestamp 1730814361
transform 1 0 2168 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5915_6
timestamp 1730814361
transform 1 0 2296 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5915_6
timestamp 1730814361
transform 1 0 2296 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5916_6
timestamp 1730814361
transform 1 0 2424 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5916_6
timestamp 1730814361
transform 1 0 2424 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_580_6
timestamp 1730814361
transform 1 0 2560 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_580_6
timestamp 1730814361
transform 1 0 2560 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_581_6
timestamp 1730814361
transform 1 0 2704 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_581_6
timestamp 1730814361
transform 1 0 2704 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_582_6
timestamp 1730814361
transform 1 0 2856 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_582_6
timestamp 1730814361
transform 1 0 2856 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_583_6
timestamp 1730814361
transform 1 0 3016 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_583_6
timestamp 1730814361
transform 1 0 3016 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5466_6
timestamp 1730814361
transform 1 0 3152 0 1 296
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5466_6
timestamp 1730814361
transform 1 0 3152 0 1 296
box 7 3 20 38
use welltap_svt  __well_tap__131
timestamp 1730814361
transform 1 0 3184 0 -1 284
box 8 4 12 24
use welltap_svt  __well_tap__133
timestamp 1730814361
transform 1 0 3184 0 1 300
box 8 4 12 24
use welltap_svt  __well_tap__131
timestamp 1730814361
transform 1 0 3184 0 -1 284
box 8 4 12 24
use welltap_svt  __well_tap__133
timestamp 1730814361
transform 1 0 3184 0 1 300
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730814361
transform 1 0 104 0 1 352
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730814361
transform 1 0 104 0 1 352
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5678_6
timestamp 1730814361
transform 1 0 640 0 1 348
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5678_6
timestamp 1730814361
transform 1 0 640 0 1 348
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5679_6
timestamp 1730814361
transform 1 0 800 0 1 348
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5679_6
timestamp 1730814361
transform 1 0 800 0 1 348
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5680_6
timestamp 1730814361
transform 1 0 944 0 1 348
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5680_6
timestamp 1730814361
transform 1 0 944 0 1 348
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5514_6
timestamp 1730814361
transform 1 0 1080 0 1 348
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5514_6
timestamp 1730814361
transform 1 0 1080 0 1 348
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5515_6
timestamp 1730814361
transform 1 0 1208 0 1 348
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5515_6
timestamp 1730814361
transform 1 0 1208 0 1 348
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5563_6
timestamp 1730814361
transform 1 0 1328 0 1 348
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5563_6
timestamp 1730814361
transform 1 0 1328 0 1 348
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5517_6
timestamp 1730814361
transform 1 0 1456 0 1 348
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5517_6
timestamp 1730814361
transform 1 0 1456 0 1 348
box 7 3 20 38
use welltap_svt  __well_tap__13
timestamp 1730814361
transform 1 0 1624 0 1 352
box 8 4 12 24
use welltap_svt  __well_tap__134
timestamp 1730814361
transform 1 0 1664 0 -1 384
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730814361
transform 1 0 1624 0 1 352
box 8 4 12 24
use welltap_svt  __well_tap__134
timestamp 1730814361
transform 1 0 1664 0 -1 384
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5917_6
timestamp 1730814361
transform 1 0 2144 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5917_6
timestamp 1730814361
transform 1 0 2144 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5918_6
timestamp 1730814361
transform 1 0 2272 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5918_6
timestamp 1730814361
transform 1 0 2272 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5919_6
timestamp 1730814361
transform 1 0 2400 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5919_6
timestamp 1730814361
transform 1 0 2400 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5920_6
timestamp 1730814361
transform 1 0 2528 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5920_6
timestamp 1730814361
transform 1 0 2528 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_584_6
timestamp 1730814361
transform 1 0 2656 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_584_6
timestamp 1730814361
transform 1 0 2656 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_585_6
timestamp 1730814361
transform 1 0 2784 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_585_6
timestamp 1730814361
transform 1 0 2784 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_586_6
timestamp 1730814361
transform 1 0 2912 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_586_6
timestamp 1730814361
transform 1 0 2912 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_587_6
timestamp 1730814361
transform 1 0 3040 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_587_6
timestamp 1730814361
transform 1 0 3040 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5467_6
timestamp 1730814361
transform 1 0 3152 0 -1 388
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5467_6
timestamp 1730814361
transform 1 0 3152 0 -1 388
box 7 3 20 38
use welltap_svt  __well_tap__135
timestamp 1730814361
transform 1 0 3184 0 -1 384
box 8 4 12 24
use welltap_svt  __well_tap__135
timestamp 1730814361
transform 1 0 3184 0 -1 384
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730814361
transform 1 0 104 0 -1 432
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730814361
transform 1 0 104 0 -1 432
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5681_6
timestamp 1730814361
transform 1 0 720 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5681_6
timestamp 1730814361
transform 1 0 720 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5682_6
timestamp 1730814361
transform 1 0 848 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5682_6
timestamp 1730814361
transform 1 0 848 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5683_6
timestamp 1730814361
transform 1 0 976 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5683_6
timestamp 1730814361
transform 1 0 976 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5684_6
timestamp 1730814361
transform 1 0 1096 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5684_6
timestamp 1730814361
transform 1 0 1096 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5518_6
timestamp 1730814361
transform 1 0 1216 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5518_6
timestamp 1730814361
transform 1 0 1216 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5519_6
timestamp 1730814361
transform 1 0 1328 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5519_6
timestamp 1730814361
transform 1 0 1328 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5520_6
timestamp 1730814361
transform 1 0 1440 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5520_6
timestamp 1730814361
transform 1 0 1440 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5521_6
timestamp 1730814361
transform 1 0 1560 0 -1 436
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5521_6
timestamp 1730814361
transform 1 0 1560 0 -1 436
box 7 3 20 38
use welltap_svt  __well_tap__15
timestamp 1730814361
transform 1 0 1624 0 -1 432
box 8 4 12 24
use welltap_svt  __well_tap__136
timestamp 1730814361
transform 1 0 1664 0 1 404
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730814361
transform 1 0 1624 0 -1 432
box 8 4 12 24
use welltap_svt  __well_tap__136
timestamp 1730814361
transform 1 0 1664 0 1 404
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5921_6
timestamp 1730814361
transform 1 0 2240 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5921_6
timestamp 1730814361
transform 1 0 2240 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5906_6
timestamp 1730814361
transform 1 0 2368 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5906_6
timestamp 1730814361
transform 1 0 2368 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5923_6
timestamp 1730814361
transform 1 0 2496 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5923_6
timestamp 1730814361
transform 1 0 2496 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5924_6
timestamp 1730814361
transform 1 0 2616 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5924_6
timestamp 1730814361
transform 1 0 2616 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_588_6
timestamp 1730814361
transform 1 0 2736 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_588_6
timestamp 1730814361
transform 1 0 2736 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_589_6
timestamp 1730814361
transform 1 0 2848 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_589_6
timestamp 1730814361
transform 1 0 2848 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_590_6
timestamp 1730814361
transform 1 0 2960 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_590_6
timestamp 1730814361
transform 1 0 2960 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_591_6
timestamp 1730814361
transform 1 0 3080 0 1 400
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_591_6
timestamp 1730814361
transform 1 0 3080 0 1 400
box 7 3 20 38
use welltap_svt  __well_tap__137
timestamp 1730814361
transform 1 0 3184 0 1 404
box 8 4 12 24
use welltap_svt  __well_tap__137
timestamp 1730814361
transform 1 0 3184 0 1 404
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5685_6
timestamp 1730814361
transform 1 0 128 0 1 448
box 7 3 20 38
use welltap_svt  __well_tap__16
timestamp 1730814361
transform 1 0 104 0 1 452
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5685_6
timestamp 1730814361
transform 1 0 128 0 1 448
box 7 3 20 38
use welltap_svt  __well_tap__16
timestamp 1730814361
transform 1 0 104 0 1 452
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5626_6
timestamp 1730814361
transform 1 0 168 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5626_6
timestamp 1730814361
transform 1 0 168 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5686_6
timestamp 1730814361
transform 1 0 224 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5686_6
timestamp 1730814361
transform 1 0 224 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5627_6
timestamp 1730814361
transform 1 0 296 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5627_6
timestamp 1730814361
transform 1 0 296 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5687_6
timestamp 1730814361
transform 1 0 352 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5687_6
timestamp 1730814361
transform 1 0 352 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5628_6
timestamp 1730814361
transform 1 0 416 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5628_6
timestamp 1730814361
transform 1 0 416 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5641_6
timestamp 1730814361
transform 1 0 496 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5641_6
timestamp 1730814361
transform 1 0 496 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5629_6
timestamp 1730814361
transform 1 0 536 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5629_6
timestamp 1730814361
transform 1 0 536 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5522_6
timestamp 1730814361
transform 1 0 648 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5526_6
timestamp 1730814361
transform 1 0 656 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5522_6
timestamp 1730814361
transform 1 0 648 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5526_6
timestamp 1730814361
transform 1 0 656 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5523_6
timestamp 1730814361
transform 1 0 808 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5527_6
timestamp 1730814361
transform 1 0 768 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5523_6
timestamp 1730814361
transform 1 0 808 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5527_6
timestamp 1730814361
transform 1 0 768 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5528_6
timestamp 1730814361
transform 1 0 880 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5528_6
timestamp 1730814361
transform 1 0 880 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5524_6
timestamp 1730814361
transform 1 0 968 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5529_6
timestamp 1730814361
transform 1 0 1000 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5524_6
timestamp 1730814361
transform 1 0 968 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5529_6
timestamp 1730814361
transform 1 0 1000 0 -1 540
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5525_6
timestamp 1730814361
transform 1 0 1128 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5525_6
timestamp 1730814361
transform 1 0 1128 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5925_6
timestamp 1730814361
transform 1 0 1288 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5925_6
timestamp 1730814361
transform 1 0 1288 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5926_6
timestamp 1730814361
transform 1 0 1448 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5926_6
timestamp 1730814361
transform 1 0 1448 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5927_6
timestamp 1730814361
transform 1 0 1592 0 1 448
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5927_6
timestamp 1730814361
transform 1 0 1592 0 1 448
box 7 3 20 38
use welltap_svt  __well_tap__17
timestamp 1730814361
transform 1 0 1624 0 1 452
box 8 4 12 24
use welltap_svt  __well_tap__138
timestamp 1730814361
transform 1 0 1664 0 -1 480
box 8 4 12 24
use welltap_svt  __well_tap__140
timestamp 1730814361
transform 1 0 1664 0 1 496
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730814361
transform 1 0 1624 0 1 452
box 8 4 12 24
use welltap_svt  __well_tap__138
timestamp 1730814361
transform 1 0 1664 0 -1 480
box 8 4 12 24
use welltap_svt  __well_tap__140
timestamp 1730814361
transform 1 0 1664 0 1 496
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5928_6
timestamp 1730814361
transform 1 0 1688 0 -1 484
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5929_6
timestamp 1730814361
transform 1 0 1688 0 1 492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5928_6
timestamp 1730814361
transform 1 0 1688 0 -1 484
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5929_6
timestamp 1730814361
transform 1 0 1688 0 1 492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5930_6
timestamp 1730814361
transform 1 0 1880 0 1 492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5930_6
timestamp 1730814361
transform 1 0 1880 0 1 492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_592_6
timestamp 1730814361
transform 1 0 2016 0 -1 484
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_592_6
timestamp 1730814361
transform 1 0 2016 0 -1 484
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5931_6
timestamp 1730814361
transform 1 0 2096 0 1 492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5931_6
timestamp 1730814361
transform 1 0 2096 0 1 492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5407_6
timestamp 1730814361
transform 1 0 2336 0 1 492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5407_6
timestamp 1730814361
transform 1 0 2336 0 1 492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_593_6
timestamp 1730814361
transform 1 0 2376 0 -1 484
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_593_6
timestamp 1730814361
transform 1 0 2376 0 -1 484
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5408_6
timestamp 1730814361
transform 1 0 2592 0 1 492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5408_6
timestamp 1730814361
transform 1 0 2592 0 1 492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5422_6
timestamp 1730814361
transform 1 0 2736 0 -1 484
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5422_6
timestamp 1730814361
transform 1 0 2736 0 -1 484
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5409_6
timestamp 1730814361
transform 1 0 2856 0 1 492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5409_6
timestamp 1730814361
transform 1 0 2856 0 1 492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5468_6
timestamp 1730814361
transform 1 0 3104 0 -1 484
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5468_6
timestamp 1730814361
transform 1 0 3104 0 -1 484
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5297_6
timestamp 1730814361
transform 1 0 3128 0 1 492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5297_6
timestamp 1730814361
transform 1 0 3128 0 1 492
box 7 3 20 38
use welltap_svt  __well_tap__139
timestamp 1730814361
transform 1 0 3184 0 -1 480
box 8 4 12 24
use welltap_svt  __well_tap__141
timestamp 1730814361
transform 1 0 3184 0 1 496
box 8 4 12 24
use welltap_svt  __well_tap__139
timestamp 1730814361
transform 1 0 3184 0 -1 480
box 8 4 12 24
use welltap_svt  __well_tap__141
timestamp 1730814361
transform 1 0 3184 0 1 496
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730814361
transform 1 0 104 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730814361
transform 1 0 104 0 1 556
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730814361
transform 1 0 104 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730814361
transform 1 0 104 0 1 556
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5630_6
timestamp 1730814361
transform 1 0 264 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5630_6
timestamp 1730814361
transform 1 0 264 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5631_6
timestamp 1730814361
transform 1 0 392 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5631_6
timestamp 1730814361
transform 1 0 392 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5632_6
timestamp 1730814361
transform 1 0 520 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5632_6
timestamp 1730814361
transform 1 0 520 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5633_6
timestamp 1730814361
transform 1 0 640 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5633_6
timestamp 1730814361
transform 1 0 640 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5530_6
timestamp 1730814361
transform 1 0 760 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5530_6
timestamp 1730814361
transform 1 0 760 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5610_6
timestamp 1730814361
transform 1 0 872 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5610_6
timestamp 1730814361
transform 1 0 872 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5595_6
timestamp 1730814361
transform 1 0 984 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5595_6
timestamp 1730814361
transform 1 0 984 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5596_6
timestamp 1730814361
transform 1 0 1104 0 1 552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5596_6
timestamp 1730814361
transform 1 0 1104 0 1 552
box 7 3 20 38
use welltap_svt  __well_tap__19
timestamp 1730814361
transform 1 0 1624 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730814361
transform 1 0 1624 0 1 556
box 8 4 12 24
use welltap_svt  __well_tap__142
timestamp 1730814361
transform 1 0 1664 0 -1 568
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730814361
transform 1 0 1624 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730814361
transform 1 0 1624 0 1 556
box 8 4 12 24
use welltap_svt  __well_tap__142
timestamp 1730814361
transform 1 0 1664 0 -1 568
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5932_6
timestamp 1730814361
transform 1 0 1760 0 -1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5932_6
timestamp 1730814361
transform 1 0 1760 0 -1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5933_6
timestamp 1730814361
transform 1 0 1920 0 -1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5933_6
timestamp 1730814361
transform 1 0 1920 0 -1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5934_6
timestamp 1730814361
transform 1 0 2080 0 -1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5934_6
timestamp 1730814361
transform 1 0 2080 0 -1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5410_6
timestamp 1730814361
transform 1 0 2240 0 -1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5410_6
timestamp 1730814361
transform 1 0 2240 0 -1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5411_6
timestamp 1730814361
transform 1 0 2400 0 -1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5411_6
timestamp 1730814361
transform 1 0 2400 0 -1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5412_6
timestamp 1730814361
transform 1 0 2560 0 -1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5412_6
timestamp 1730814361
transform 1 0 2560 0 -1 572
box 7 3 20 38
use welltap_svt  __well_tap__143
timestamp 1730814361
transform 1 0 3184 0 -1 568
box 8 4 12 24
use welltap_svt  __well_tap__143
timestamp 1730814361
transform 1 0 3184 0 -1 568
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730814361
transform 1 0 104 0 -1 636
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730814361
transform 1 0 104 0 -1 636
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5634_6
timestamp 1730814361
transform 1 0 368 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5634_6
timestamp 1730814361
transform 1 0 368 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5635_6
timestamp 1730814361
transform 1 0 496 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5635_6
timestamp 1730814361
transform 1 0 496 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5636_6
timestamp 1730814361
transform 1 0 616 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5636_6
timestamp 1730814361
transform 1 0 616 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5637_6
timestamp 1730814361
transform 1 0 736 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5637_6
timestamp 1730814361
transform 1 0 736 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5597_6
timestamp 1730814361
transform 1 0 856 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5597_6
timestamp 1730814361
transform 1 0 856 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5598_6
timestamp 1730814361
transform 1 0 968 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5598_6
timestamp 1730814361
transform 1 0 968 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5599_6
timestamp 1730814361
transform 1 0 1088 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5599_6
timestamp 1730814361
transform 1 0 1088 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5600_6
timestamp 1730814361
transform 1 0 1208 0 -1 640
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5600_6
timestamp 1730814361
transform 1 0 1208 0 -1 640
box 7 3 20 38
use welltap_svt  __well_tap__23
timestamp 1730814361
transform 1 0 1624 0 -1 636
box 8 4 12 24
use welltap_svt  __well_tap__144
timestamp 1730814361
transform 1 0 1664 0 1 576
box 8 4 12 24
use welltap_svt  __well_tap__146
timestamp 1730814361
transform 1 0 1664 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730814361
transform 1 0 1624 0 -1 636
box 8 4 12 24
use welltap_svt  __well_tap__144
timestamp 1730814361
transform 1 0 1664 0 1 576
box 8 4 12 24
use welltap_svt  __well_tap__146
timestamp 1730814361
transform 1 0 1664 0 -1 652
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5935_6
timestamp 1730814361
transform 1 0 1840 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5935_6
timestamp 1730814361
transform 1 0 1840 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5891_6
timestamp 1730814361
transform 1 0 1912 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5891_6
timestamp 1730814361
transform 1 0 1912 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5876_6
timestamp 1730814361
transform 1 0 2040 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5936_6
timestamp 1730814361
transform 1 0 2008 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5876_6
timestamp 1730814361
transform 1 0 2040 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5936_6
timestamp 1730814361
transform 1 0 2008 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5877_6
timestamp 1730814361
transform 1 0 2176 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5937_6
timestamp 1730814361
transform 1 0 2176 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5877_6
timestamp 1730814361
transform 1 0 2176 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5937_6
timestamp 1730814361
transform 1 0 2176 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5413_6
timestamp 1730814361
transform 1 0 2352 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5878_6
timestamp 1730814361
transform 1 0 2320 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5413_6
timestamp 1730814361
transform 1 0 2352 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5878_6
timestamp 1730814361
transform 1 0 2320 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5417_6
timestamp 1730814361
transform 1 0 2464 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5417_6
timestamp 1730814361
transform 1 0 2464 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5414_6
timestamp 1730814361
transform 1 0 2544 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5414_6
timestamp 1730814361
transform 1 0 2544 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5418_6
timestamp 1730814361
transform 1 0 2608 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5418_6
timestamp 1730814361
transform 1 0 2608 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5415_6
timestamp 1730814361
transform 1 0 2744 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5419_6
timestamp 1730814361
transform 1 0 2752 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5415_6
timestamp 1730814361
transform 1 0 2744 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5419_6
timestamp 1730814361
transform 1 0 2752 0 -1 656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5416_6
timestamp 1730814361
transform 1 0 2952 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5416_6
timestamp 1730814361
transform 1 0 2952 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5282_6
timestamp 1730814361
transform 1 0 3152 0 1 572
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5282_6
timestamp 1730814361
transform 1 0 3152 0 1 572
box 7 3 20 38
use welltap_svt  __well_tap__145
timestamp 1730814361
transform 1 0 3184 0 1 576
box 8 4 12 24
use welltap_svt  __well_tap__147
timestamp 1730814361
transform 1 0 3184 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__145
timestamp 1730814361
transform 1 0 3184 0 1 576
box 8 4 12 24
use welltap_svt  __well_tap__147
timestamp 1730814361
transform 1 0 3184 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730814361
transform 1 0 104 0 1 656
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730814361
transform 1 0 104 0 1 656
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5638_6
timestamp 1730814361
transform 1 0 472 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5638_6
timestamp 1730814361
transform 1 0 472 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5639_6
timestamp 1730814361
transform 1 0 600 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5639_6
timestamp 1730814361
transform 1 0 600 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5640_6
timestamp 1730814361
transform 1 0 720 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5640_6
timestamp 1730814361
transform 1 0 720 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5688_6
timestamp 1730814361
transform 1 0 840 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5688_6
timestamp 1730814361
transform 1 0 840 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5601_6
timestamp 1730814361
transform 1 0 960 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5601_6
timestamp 1730814361
transform 1 0 960 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5602_6
timestamp 1730814361
transform 1 0 1072 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5602_6
timestamp 1730814361
transform 1 0 1072 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5603_6
timestamp 1730814361
transform 1 0 1184 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5603_6
timestamp 1730814361
transform 1 0 1184 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5604_6
timestamp 1730814361
transform 1 0 1304 0 1 652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5604_6
timestamp 1730814361
transform 1 0 1304 0 1 652
box 7 3 20 38
use welltap_svt  __well_tap__25
timestamp 1730814361
transform 1 0 1624 0 1 656
box 8 4 12 24
use welltap_svt  __well_tap__148
timestamp 1730814361
transform 1 0 1664 0 1 668
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730814361
transform 1 0 1624 0 1 656
box 8 4 12 24
use welltap_svt  __well_tap__148
timestamp 1730814361
transform 1 0 1664 0 1 668
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5879_6
timestamp 1730814361
transform 1 0 2016 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5879_6
timestamp 1730814361
transform 1 0 2016 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5880_6
timestamp 1730814361
transform 1 0 2144 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5880_6
timestamp 1730814361
transform 1 0 2144 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5881_6
timestamp 1730814361
transform 1 0 2288 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5881_6
timestamp 1730814361
transform 1 0 2288 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5882_6
timestamp 1730814361
transform 1 0 2440 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5882_6
timestamp 1730814361
transform 1 0 2440 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5420_6
timestamp 1730814361
transform 1 0 2608 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5420_6
timestamp 1730814361
transform 1 0 2608 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5421_6
timestamp 1730814361
transform 1 0 2792 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5421_6
timestamp 1730814361
transform 1 0 2792 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5406_6
timestamp 1730814361
transform 1 0 2984 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5406_6
timestamp 1730814361
transform 1 0 2984 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5283_6
timestamp 1730814361
transform 1 0 3152 0 1 664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5283_6
timestamp 1730814361
transform 1 0 3152 0 1 664
box 7 3 20 38
use welltap_svt  __well_tap__149
timestamp 1730814361
transform 1 0 3184 0 1 668
box 8 4 12 24
use welltap_svt  __well_tap__149
timestamp 1730814361
transform 1 0 3184 0 1 668
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730814361
transform 1 0 104 0 -1 740
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730814361
transform 1 0 104 0 -1 740
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5642_6
timestamp 1730814361
transform 1 0 568 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5642_6
timestamp 1730814361
transform 1 0 568 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5643_6
timestamp 1730814361
transform 1 0 696 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5643_6
timestamp 1730814361
transform 1 0 696 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5644_6
timestamp 1730814361
transform 1 0 824 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5644_6
timestamp 1730814361
transform 1 0 824 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5645_6
timestamp 1730814361
transform 1 0 944 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5645_6
timestamp 1730814361
transform 1 0 944 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5605_6
timestamp 1730814361
transform 1 0 1064 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5605_6
timestamp 1730814361
transform 1 0 1064 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5606_6
timestamp 1730814361
transform 1 0 1176 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5606_6
timestamp 1730814361
transform 1 0 1176 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5607_6
timestamp 1730814361
transform 1 0 1288 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5607_6
timestamp 1730814361
transform 1 0 1288 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5608_6
timestamp 1730814361
transform 1 0 1408 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5608_6
timestamp 1730814361
transform 1 0 1408 0 -1 744
box 7 3 20 38
use welltap_svt  __well_tap__27
timestamp 1730814361
transform 1 0 1624 0 -1 740
box 8 4 12 24
use welltap_svt  __well_tap__150
timestamp 1730814361
transform 1 0 1664 0 -1 740
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730814361
transform 1 0 1624 0 -1 740
box 8 4 12 24
use welltap_svt  __well_tap__150
timestamp 1730814361
transform 1 0 1664 0 -1 740
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5883_6
timestamp 1730814361
transform 1 0 2120 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5883_6
timestamp 1730814361
transform 1 0 2120 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5886_6
timestamp 1730814361
transform 1 0 2192 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5886_6
timestamp 1730814361
transform 1 0 2192 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5884_6
timestamp 1730814361
transform 1 0 2280 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5884_6
timestamp 1730814361
transform 1 0 2280 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5887_6
timestamp 1730814361
transform 1 0 2352 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5887_6
timestamp 1730814361
transform 1 0 2352 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5885_6
timestamp 1730814361
transform 1 0 2440 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5885_6
timestamp 1730814361
transform 1 0 2440 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5888_6
timestamp 1730814361
transform 1 0 2504 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5888_6
timestamp 1730814361
transform 1 0 2504 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5423_6
timestamp 1730814361
transform 1 0 2592 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5423_6
timestamp 1730814361
transform 1 0 2592 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5426_6
timestamp 1730814361
transform 1 0 2648 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5426_6
timestamp 1730814361
transform 1 0 2648 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5424_6
timestamp 1730814361
transform 1 0 2752 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5427_6
timestamp 1730814361
transform 1 0 2784 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5424_6
timestamp 1730814361
transform 1 0 2752 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5427_6
timestamp 1730814361
transform 1 0 2784 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5425_6
timestamp 1730814361
transform 1 0 2912 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5428_6
timestamp 1730814361
transform 1 0 2912 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5425_6
timestamp 1730814361
transform 1 0 2912 0 -1 744
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5428_6
timestamp 1730814361
transform 1 0 2912 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5429_6
timestamp 1730814361
transform 1 0 3040 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5429_6
timestamp 1730814361
transform 1 0 3040 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5284_6
timestamp 1730814361
transform 1 0 3152 0 1 748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5284_6
timestamp 1730814361
transform 1 0 3152 0 1 748
box 7 3 20 38
use welltap_svt  __well_tap__151
timestamp 1730814361
transform 1 0 3184 0 -1 740
box 8 4 12 24
use welltap_svt  __well_tap__151
timestamp 1730814361
transform 1 0 3184 0 -1 740
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5652_6
timestamp 1730814361
transform 1 0 128 0 -1 848
box 7 3 20 38
use welltap_svt  __well_tap__28
timestamp 1730814361
transform 1 0 104 0 1 756
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5652_6
timestamp 1730814361
transform 1 0 128 0 -1 848
box 7 3 20 38
use welltap_svt  __well_tap__28
timestamp 1730814361
transform 1 0 104 0 1 756
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5653_6
timestamp 1730814361
transform 1 0 296 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5653_6
timestamp 1730814361
transform 1 0 296 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5650_6
timestamp 1730814361
transform 1 0 496 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5650_6
timestamp 1730814361
transform 1 0 496 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5646_6
timestamp 1730814361
transform 1 0 672 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5651_6
timestamp 1730814361
transform 1 0 688 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5646_6
timestamp 1730814361
transform 1 0 672 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5651_6
timestamp 1730814361
transform 1 0 688 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5647_6
timestamp 1730814361
transform 1 0 800 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5647_6
timestamp 1730814361
transform 1 0 800 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5615_6
timestamp 1730814361
transform 1 0 872 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5615_6
timestamp 1730814361
transform 1 0 872 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5648_6
timestamp 1730814361
transform 1 0 920 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5648_6
timestamp 1730814361
transform 1 0 920 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5616_6
timestamp 1730814361
transform 1 0 1040 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5649_6
timestamp 1730814361
transform 1 0 1040 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5616_6
timestamp 1730814361
transform 1 0 1040 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5649_6
timestamp 1730814361
transform 1 0 1040 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5609_6
timestamp 1730814361
transform 1 0 1160 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5609_6
timestamp 1730814361
transform 1 0 1160 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5613_6
timestamp 1730814361
transform 1 0 1192 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5613_6
timestamp 1730814361
transform 1 0 1192 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5594_6
timestamp 1730814361
transform 1 0 1272 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5594_6
timestamp 1730814361
transform 1 0 1272 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5614_6
timestamp 1730814361
transform 1 0 1328 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5614_6
timestamp 1730814361
transform 1 0 1328 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5611_6
timestamp 1730814361
transform 1 0 1392 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5611_6
timestamp 1730814361
transform 1 0 1392 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5892_6
timestamp 1730814361
transform 1 0 1464 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5892_6
timestamp 1730814361
transform 1 0 1464 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5612_6
timestamp 1730814361
transform 1 0 1512 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5612_6
timestamp 1730814361
transform 1 0 1512 0 1 752
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5893_6
timestamp 1730814361
transform 1 0 1592 0 -1 848
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5893_6
timestamp 1730814361
transform 1 0 1592 0 -1 848
box 7 3 20 38
use welltap_svt  __well_tap__29
timestamp 1730814361
transform 1 0 1624 0 1 756
box 8 4 12 24
use welltap_svt  __well_tap__152
timestamp 1730814361
transform 1 0 1664 0 1 752
box 8 4 12 24
use welltap_svt  __well_tap__154
timestamp 1730814361
transform 1 0 1664 0 -1 828
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1730814361
transform 1 0 1624 0 1 756
box 8 4 12 24
use welltap_svt  __well_tap__152
timestamp 1730814361
transform 1 0 1664 0 1 752
box 8 4 12 24
use welltap_svt  __well_tap__154
timestamp 1730814361
transform 1 0 1664 0 -1 828
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5889_6
timestamp 1730814361
transform 1 0 2272 0 -1 832
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5889_6
timestamp 1730814361
transform 1 0 2272 0 -1 832
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5890_6
timestamp 1730814361
transform 1 0 2432 0 -1 832
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5890_6
timestamp 1730814361
transform 1 0 2432 0 -1 832
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5938_6
timestamp 1730814361
transform 1 0 2576 0 -1 832
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5938_6
timestamp 1730814361
transform 1 0 2576 0 -1 832
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5430_6
timestamp 1730814361
transform 1 0 2712 0 -1 832
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5430_6
timestamp 1730814361
transform 1 0 2712 0 -1 832
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5432_6
timestamp 1730814361
transform 1 0 2840 0 -1 832
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5432_6
timestamp 1730814361
transform 1 0 2840 0 -1 832
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5431_6
timestamp 1730814361
transform 1 0 2968 0 -1 832
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5431_6
timestamp 1730814361
transform 1 0 2968 0 -1 832
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5285_6
timestamp 1730814361
transform 1 0 3104 0 -1 832
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5285_6
timestamp 1730814361
transform 1 0 3104 0 -1 832
box 7 3 20 38
use welltap_svt  __well_tap__153
timestamp 1730814361
transform 1 0 3184 0 1 752
box 8 4 12 24
use welltap_svt  __well_tap__155
timestamp 1730814361
transform 1 0 3184 0 -1 828
box 8 4 12 24
use welltap_svt  __well_tap__153
timestamp 1730814361
transform 1 0 3184 0 1 752
box 8 4 12 24
use welltap_svt  __well_tap__155
timestamp 1730814361
transform 1 0 3184 0 -1 828
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5654_6
timestamp 1730814361
transform 1 0 128 0 1 852
box 7 3 20 38
use welltap_svt  __well_tap__30
timestamp 1730814361
transform 1 0 104 0 -1 844
box 8 4 12 24
use welltap_svt  __well_tap__32
timestamp 1730814361
transform 1 0 104 0 1 856
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5654_6
timestamp 1730814361
transform 1 0 128 0 1 852
box 7 3 20 38
use welltap_svt  __well_tap__30
timestamp 1730814361
transform 1 0 104 0 -1 844
box 8 4 12 24
use welltap_svt  __well_tap__32
timestamp 1730814361
transform 1 0 104 0 1 856
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5655_6
timestamp 1730814361
transform 1 0 240 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5655_6
timestamp 1730814361
transform 1 0 240 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5735_6
timestamp 1730814361
transform 1 0 376 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5735_6
timestamp 1730814361
transform 1 0 376 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5720_6
timestamp 1730814361
transform 1 0 528 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5720_6
timestamp 1730814361
transform 1 0 528 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5617_6
timestamp 1730814361
transform 1 0 704 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5617_6
timestamp 1730814361
transform 1 0 704 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5618_6
timestamp 1730814361
transform 1 0 912 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5618_6
timestamp 1730814361
transform 1 0 912 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5619_6
timestamp 1730814361
transform 1 0 1136 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5619_6
timestamp 1730814361
transform 1 0 1136 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5620_6
timestamp 1730814361
transform 1 0 1376 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5620_6
timestamp 1730814361
transform 1 0 1376 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5894_6
timestamp 1730814361
transform 1 0 1592 0 1 852
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5894_6
timestamp 1730814361
transform 1 0 1592 0 1 852
box 7 3 20 38
use welltap_svt  __well_tap__31
timestamp 1730814361
transform 1 0 1624 0 -1 844
box 8 4 12 24
use welltap_svt  __well_tap__33
timestamp 1730814361
transform 1 0 1624 0 1 856
box 8 4 12 24
use welltap_svt  __well_tap__156
timestamp 1730814361
transform 1 0 1664 0 1 848
box 8 4 12 24
use welltap_svt  __well_tap__31
timestamp 1730814361
transform 1 0 1624 0 -1 844
box 8 4 12 24
use welltap_svt  __well_tap__33
timestamp 1730814361
transform 1 0 1624 0 1 856
box 8 4 12 24
use welltap_svt  __well_tap__156
timestamp 1730814361
transform 1 0 1664 0 1 848
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5895_6
timestamp 1730814361
transform 1 0 1688 0 1 844
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5895_6
timestamp 1730814361
transform 1 0 1688 0 1 844
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5896_6
timestamp 1730814361
transform 1 0 2008 0 1 844
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5896_6
timestamp 1730814361
transform 1 0 2008 0 1 844
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5434_6
timestamp 1730814361
transform 1 0 2360 0 1 844
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5434_6
timestamp 1730814361
transform 1 0 2360 0 1 844
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5435_6
timestamp 1730814361
transform 1 0 2720 0 1 844
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5435_6
timestamp 1730814361
transform 1 0 2720 0 1 844
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5433_6
timestamp 1730814361
transform 1 0 3080 0 1 844
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5433_6
timestamp 1730814361
transform 1 0 3080 0 1 844
box 7 3 20 38
use welltap_svt  __well_tap__157
timestamp 1730814361
transform 1 0 3184 0 1 848
box 8 4 12 24
use welltap_svt  __well_tap__157
timestamp 1730814361
transform 1 0 3184 0 1 848
box 8 4 12 24
use welltap_svt  __well_tap__34
timestamp 1730814361
transform 1 0 104 0 -1 940
box 8 4 12 24
use welltap_svt  __well_tap__34
timestamp 1730814361
transform 1 0 104 0 -1 940
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5721_6
timestamp 1730814361
transform 1 0 216 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5721_6
timestamp 1730814361
transform 1 0 216 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5722_6
timestamp 1730814361
transform 1 0 344 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5722_6
timestamp 1730814361
transform 1 0 344 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5723_6
timestamp 1730814361
transform 1 0 464 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5723_6
timestamp 1730814361
transform 1 0 464 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5724_6
timestamp 1730814361
transform 1 0 584 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5724_6
timestamp 1730814361
transform 1 0 584 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5621_6
timestamp 1730814361
transform 1 0 704 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5621_6
timestamp 1730814361
transform 1 0 704 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5622_6
timestamp 1730814361
transform 1 0 816 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5622_6
timestamp 1730814361
transform 1 0 816 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5623_6
timestamp 1730814361
transform 1 0 936 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5623_6
timestamp 1730814361
transform 1 0 936 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5624_6
timestamp 1730814361
transform 1 0 1056 0 -1 944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5624_6
timestamp 1730814361
transform 1 0 1056 0 -1 944
box 7 3 20 38
use welltap_svt  __well_tap__35
timestamp 1730814361
transform 1 0 1624 0 -1 940
box 8 4 12 24
use welltap_svt  __well_tap__158
timestamp 1730814361
transform 1 0 1664 0 -1 920
box 8 4 12 24
use welltap_svt  __well_tap__35
timestamp 1730814361
transform 1 0 1624 0 -1 940
box 8 4 12 24
use welltap_svt  __well_tap__158
timestamp 1730814361
transform 1 0 1664 0 -1 920
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5897_6
timestamp 1730814361
transform 1 0 1712 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5897_6
timestamp 1730814361
transform 1 0 1712 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5900_6
timestamp 1730814361
transform 1 0 1784 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5900_6
timestamp 1730814361
transform 1 0 1784 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5898_6
timestamp 1730814361
transform 1 0 1864 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5898_6
timestamp 1730814361
transform 1 0 1864 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5901_6
timestamp 1730814361
transform 1 0 1912 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5901_6
timestamp 1730814361
transform 1 0 1912 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5899_6
timestamp 1730814361
transform 1 0 2032 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5899_6
timestamp 1730814361
transform 1 0 2032 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5902_6
timestamp 1730814361
transform 1 0 2064 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5902_6
timestamp 1730814361
transform 1 0 2064 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5436_6
timestamp 1730814361
transform 1 0 2216 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5436_6
timestamp 1730814361
transform 1 0 2216 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5903_6
timestamp 1730814361
transform 1 0 2248 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5903_6
timestamp 1730814361
transform 1 0 2248 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5377_6
timestamp 1730814361
transform 1 0 2456 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5437_6
timestamp 1730814361
transform 1 0 2432 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5377_6
timestamp 1730814361
transform 1 0 2456 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5437_6
timestamp 1730814361
transform 1 0 2432 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5391_6
timestamp 1730814361
transform 1 0 2664 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5391_6
timestamp 1730814361
transform 1 0 2664 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5378_6
timestamp 1730814361
transform 1 0 2688 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5378_6
timestamp 1730814361
transform 1 0 2688 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5376_6
timestamp 1730814361
transform 1 0 2904 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5376_6
timestamp 1730814361
transform 1 0 2904 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5379_6
timestamp 1730814361
transform 1 0 2928 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5379_6
timestamp 1730814361
transform 1 0 2928 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5286_6
timestamp 1730814361
transform 1 0 3152 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5287_6
timestamp 1730814361
transform 1 0 3152 0 1 932
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5286_6
timestamp 1730814361
transform 1 0 3152 0 -1 924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5287_6
timestamp 1730814361
transform 1 0 3152 0 1 932
box 7 3 20 38
use welltap_svt  __well_tap__159
timestamp 1730814361
transform 1 0 3184 0 -1 920
box 8 4 12 24
use welltap_svt  __well_tap__159
timestamp 1730814361
transform 1 0 3184 0 -1 920
box 8 4 12 24
use welltap_svt  __well_tap__36
timestamp 1730814361
transform 1 0 104 0 1 960
box 8 4 12 24
use welltap_svt  __well_tap__36
timestamp 1730814361
transform 1 0 104 0 1 960
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5725_6
timestamp 1730814361
transform 1 0 320 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5725_6
timestamp 1730814361
transform 1 0 320 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5726_6
timestamp 1730814361
transform 1 0 448 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5726_6
timestamp 1730814361
transform 1 0 448 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5727_6
timestamp 1730814361
transform 1 0 568 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5727_6
timestamp 1730814361
transform 1 0 568 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5728_6
timestamp 1730814361
transform 1 0 688 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5728_6
timestamp 1730814361
transform 1 0 688 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5579_6
timestamp 1730814361
transform 1 0 808 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5579_6
timestamp 1730814361
transform 1 0 808 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5564_6
timestamp 1730814361
transform 1 0 920 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5564_6
timestamp 1730814361
transform 1 0 920 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5565_6
timestamp 1730814361
transform 1 0 1032 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5565_6
timestamp 1730814361
transform 1 0 1032 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5566_6
timestamp 1730814361
transform 1 0 1152 0 1 956
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5566_6
timestamp 1730814361
transform 1 0 1152 0 1 956
box 7 3 20 38
use welltap_svt  __well_tap__37
timestamp 1730814361
transform 1 0 1624 0 1 960
box 8 4 12 24
use welltap_svt  __well_tap__160
timestamp 1730814361
transform 1 0 1664 0 1 936
box 8 4 12 24
use welltap_svt  __well_tap__162
timestamp 1730814361
transform 1 0 1664 0 -1 1008
box 8 4 12 24
use welltap_svt  __well_tap__37
timestamp 1730814361
transform 1 0 1624 0 1 960
box 8 4 12 24
use welltap_svt  __well_tap__160
timestamp 1730814361
transform 1 0 1664 0 1 936
box 8 4 12 24
use welltap_svt  __well_tap__162
timestamp 1730814361
transform 1 0 1664 0 -1 1008
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5904_6
timestamp 1730814361
transform 1 0 1888 0 -1 1012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5904_6
timestamp 1730814361
transform 1 0 1888 0 -1 1012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5905_6
timestamp 1730814361
transform 1 0 2040 0 -1 1012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5905_6
timestamp 1730814361
transform 1 0 2040 0 -1 1012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5985_6
timestamp 1730814361
transform 1 0 2192 0 -1 1012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5985_6
timestamp 1730814361
transform 1 0 2192 0 -1 1012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5380_6
timestamp 1730814361
transform 1 0 2336 0 -1 1012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5380_6
timestamp 1730814361
transform 1 0 2336 0 -1 1012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5381_6
timestamp 1730814361
transform 1 0 2488 0 -1 1012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5381_6
timestamp 1730814361
transform 1 0 2488 0 -1 1012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5382_6
timestamp 1730814361
transform 1 0 2640 0 -1 1012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5382_6
timestamp 1730814361
transform 1 0 2640 0 -1 1012
box 7 3 20 38
use welltap_svt  __well_tap__161
timestamp 1730814361
transform 1 0 3184 0 1 936
box 8 4 12 24
use welltap_svt  __well_tap__163
timestamp 1730814361
transform 1 0 3184 0 -1 1008
box 8 4 12 24
use welltap_svt  __well_tap__161
timestamp 1730814361
transform 1 0 3184 0 1 936
box 8 4 12 24
use welltap_svt  __well_tap__163
timestamp 1730814361
transform 1 0 3184 0 -1 1008
box 8 4 12 24
use welltap_svt  __well_tap__38
timestamp 1730814361
transform 1 0 104 0 -1 1044
box 8 4 12 24
use welltap_svt  __well_tap__38
timestamp 1730814361
transform 1 0 104 0 -1 1044
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5729_6
timestamp 1730814361
transform 1 0 416 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5729_6
timestamp 1730814361
transform 1 0 416 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5730_6
timestamp 1730814361
transform 1 0 544 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5733_6
timestamp 1730814361
transform 1 0 520 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5730_6
timestamp 1730814361
transform 1 0 544 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5733_6
timestamp 1730814361
transform 1 0 520 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5731_6
timestamp 1730814361
transform 1 0 672 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5734_6
timestamp 1730814361
transform 1 0 648 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5731_6
timestamp 1730814361
transform 1 0 672 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5734_6
timestamp 1730814361
transform 1 0 648 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5719_6
timestamp 1730814361
transform 1 0 768 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5732_6
timestamp 1730814361
transform 1 0 792 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5719_6
timestamp 1730814361
transform 1 0 768 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5732_6
timestamp 1730814361
transform 1 0 792 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5567_6
timestamp 1730814361
transform 1 0 912 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5736_6
timestamp 1730814361
transform 1 0 888 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5567_6
timestamp 1730814361
transform 1 0 912 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5736_6
timestamp 1730814361
transform 1 0 888 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5568_6
timestamp 1730814361
transform 1 0 1024 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5571_6
timestamp 1730814361
transform 1 0 1008 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5568_6
timestamp 1730814361
transform 1 0 1024 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5571_6
timestamp 1730814361
transform 1 0 1008 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5572_6
timestamp 1730814361
transform 1 0 1120 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5572_6
timestamp 1730814361
transform 1 0 1120 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5569_6
timestamp 1730814361
transform 1 0 1136 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5569_6
timestamp 1730814361
transform 1 0 1136 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5573_6
timestamp 1730814361
transform 1 0 1240 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5573_6
timestamp 1730814361
transform 1 0 1240 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5570_6
timestamp 1730814361
transform 1 0 1256 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5570_6
timestamp 1730814361
transform 1 0 1256 0 -1 1048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5574_6
timestamp 1730814361
transform 1 0 1360 0 1 1056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5574_6
timestamp 1730814361
transform 1 0 1360 0 1 1056
box 7 3 20 38
use welltap_svt  __well_tap__39
timestamp 1730814361
transform 1 0 1624 0 -1 1044
box 8 4 12 24
use welltap_svt  __well_tap__164
timestamp 1730814361
transform 1 0 1664 0 1 1020
box 8 4 12 24
use welltap_svt  __well_tap__39
timestamp 1730814361
transform 1 0 1624 0 -1 1044
box 8 4 12 24
use welltap_svt  __well_tap__164
timestamp 1730814361
transform 1 0 1664 0 1 1020
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5970_6
timestamp 1730814361
transform 1 0 1968 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5970_6
timestamp 1730814361
transform 1 0 1968 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5971_6
timestamp 1730814361
transform 1 0 2088 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5971_6
timestamp 1730814361
transform 1 0 2088 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5972_6
timestamp 1730814361
transform 1 0 2208 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5972_6
timestamp 1730814361
transform 1 0 2208 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5973_6
timestamp 1730814361
transform 1 0 2336 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5973_6
timestamp 1730814361
transform 1 0 2336 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5383_6
timestamp 1730814361
transform 1 0 2480 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5383_6
timestamp 1730814361
transform 1 0 2480 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5384_6
timestamp 1730814361
transform 1 0 2640 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5384_6
timestamp 1730814361
transform 1 0 2640 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5385_6
timestamp 1730814361
transform 1 0 2816 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5385_6
timestamp 1730814361
transform 1 0 2816 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5386_6
timestamp 1730814361
transform 1 0 2992 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5386_6
timestamp 1730814361
transform 1 0 2992 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5288_6
timestamp 1730814361
transform 1 0 3152 0 1 1016
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5288_6
timestamp 1730814361
transform 1 0 3152 0 1 1016
box 7 3 20 38
use welltap_svt  __well_tap__165
timestamp 1730814361
transform 1 0 3184 0 1 1020
box 8 4 12 24
use welltap_svt  __well_tap__165
timestamp 1730814361
transform 1 0 3184 0 1 1020
box 8 4 12 24
use welltap_svt  __well_tap__40
timestamp 1730814361
transform 1 0 104 0 1 1060
box 8 4 12 24
use welltap_svt  __well_tap__42
timestamp 1730814361
transform 1 0 104 0 -1 1144
box 8 4 12 24
use welltap_svt  __well_tap__40
timestamp 1730814361
transform 1 0 104 0 1 1060
box 8 4 12 24
use welltap_svt  __well_tap__42
timestamp 1730814361
transform 1 0 104 0 -1 1144
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5737_6
timestamp 1730814361
transform 1 0 624 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5737_6
timestamp 1730814361
transform 1 0 624 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5738_6
timestamp 1730814361
transform 1 0 752 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5738_6
timestamp 1730814361
transform 1 0 752 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5739_6
timestamp 1730814361
transform 1 0 872 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5739_6
timestamp 1730814361
transform 1 0 872 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5740_6
timestamp 1730814361
transform 1 0 992 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5740_6
timestamp 1730814361
transform 1 0 992 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5575_6
timestamp 1730814361
transform 1 0 1112 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5575_6
timestamp 1730814361
transform 1 0 1112 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5576_6
timestamp 1730814361
transform 1 0 1224 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5576_6
timestamp 1730814361
transform 1 0 1224 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5577_6
timestamp 1730814361
transform 1 0 1336 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5577_6
timestamp 1730814361
transform 1 0 1336 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5578_6
timestamp 1730814361
transform 1 0 1456 0 -1 1148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5578_6
timestamp 1730814361
transform 1 0 1456 0 -1 1148
box 7 3 20 38
use welltap_svt  __well_tap__41
timestamp 1730814361
transform 1 0 1624 0 1 1060
box 8 4 12 24
use welltap_svt  __well_tap__43
timestamp 1730814361
transform 1 0 1624 0 -1 1144
box 8 4 12 24
use welltap_svt  __well_tap__166
timestamp 1730814361
transform 1 0 1664 0 -1 1104
box 8 4 12 24
use welltap_svt  __well_tap__168
timestamp 1730814361
transform 1 0 1664 0 1 1116
box 8 4 12 24
use welltap_svt  __well_tap__41
timestamp 1730814361
transform 1 0 1624 0 1 1060
box 8 4 12 24
use welltap_svt  __well_tap__43
timestamp 1730814361
transform 1 0 1624 0 -1 1144
box 8 4 12 24
use welltap_svt  __well_tap__166
timestamp 1730814361
transform 1 0 1664 0 -1 1104
box 8 4 12 24
use welltap_svt  __well_tap__168
timestamp 1730814361
transform 1 0 1664 0 1 1116
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5974_6
timestamp 1730814361
transform 1 0 2064 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5974_6
timestamp 1730814361
transform 1 0 2064 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5978_6
timestamp 1730814361
transform 1 0 2168 0 1 1112
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5978_6
timestamp 1730814361
transform 1 0 2168 0 1 1112
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5975_6
timestamp 1730814361
transform 1 0 2184 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5975_6
timestamp 1730814361
transform 1 0 2184 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5976_6
timestamp 1730814361
transform 1 0 2320 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5979_6
timestamp 1730814361
transform 1 0 2328 0 1 1112
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5976_6
timestamp 1730814361
transform 1 0 2320 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5979_6
timestamp 1730814361
transform 1 0 2328 0 1 1112
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5977_6
timestamp 1730814361
transform 1 0 2472 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5980_6
timestamp 1730814361
transform 1 0 2488 0 1 1112
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5977_6
timestamp 1730814361
transform 1 0 2472 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5980_6
timestamp 1730814361
transform 1 0 2488 0 1 1112
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5387_6
timestamp 1730814361
transform 1 0 2632 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5390_6
timestamp 1730814361
transform 1 0 2648 0 1 1112
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5387_6
timestamp 1730814361
transform 1 0 2632 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5390_6
timestamp 1730814361
transform 1 0 2648 0 1 1112
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5388_6
timestamp 1730814361
transform 1 0 2808 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5438_6
timestamp 1730814361
transform 1 0 2808 0 1 1112
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5388_6
timestamp 1730814361
transform 1 0 2808 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5438_6
timestamp 1730814361
transform 1 0 2808 0 1 1112
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5392_6
timestamp 1730814361
transform 1 0 2968 0 1 1112
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5392_6
timestamp 1730814361
transform 1 0 2968 0 1 1112
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5389_6
timestamp 1730814361
transform 1 0 2992 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5389_6
timestamp 1730814361
transform 1 0 2992 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5289_6
timestamp 1730814361
transform 1 0 3152 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5290_6
timestamp 1730814361
transform 1 0 3128 0 1 1112
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5289_6
timestamp 1730814361
transform 1 0 3152 0 -1 1108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5290_6
timestamp 1730814361
transform 1 0 3128 0 1 1112
box 7 3 20 38
use welltap_svt  __well_tap__167
timestamp 1730814361
transform 1 0 3184 0 -1 1104
box 8 4 12 24
use welltap_svt  __well_tap__169
timestamp 1730814361
transform 1 0 3184 0 1 1116
box 8 4 12 24
use welltap_svt  __well_tap__167
timestamp 1730814361
transform 1 0 3184 0 -1 1104
box 8 4 12 24
use welltap_svt  __well_tap__169
timestamp 1730814361
transform 1 0 3184 0 1 1116
box 8 4 12 24
use welltap_svt  __well_tap__44
timestamp 1730814361
transform 1 0 104 0 1 1164
box 8 4 12 24
use welltap_svt  __well_tap__44
timestamp 1730814361
transform 1 0 104 0 1 1164
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5741_6
timestamp 1730814361
transform 1 0 720 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5741_6
timestamp 1730814361
transform 1 0 720 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5742_6
timestamp 1730814361
transform 1 0 848 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5742_6
timestamp 1730814361
transform 1 0 848 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5743_6
timestamp 1730814361
transform 1 0 976 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5743_6
timestamp 1730814361
transform 1 0 976 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5744_6
timestamp 1730814361
transform 1 0 1096 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5744_6
timestamp 1730814361
transform 1 0 1096 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5750_6
timestamp 1730814361
transform 1 0 1216 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5750_6
timestamp 1730814361
transform 1 0 1216 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5580_6
timestamp 1730814361
transform 1 0 1328 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5580_6
timestamp 1730814361
transform 1 0 1328 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5581_6
timestamp 1730814361
transform 1 0 1440 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5581_6
timestamp 1730814361
transform 1 0 1440 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5582_6
timestamp 1730814361
transform 1 0 1560 0 1 1160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5582_6
timestamp 1730814361
transform 1 0 1560 0 1 1160
box 7 3 20 38
use welltap_svt  __well_tap__45
timestamp 1730814361
transform 1 0 1624 0 1 1164
box 8 4 12 24
use welltap_svt  __well_tap__170
timestamp 1730814361
transform 1 0 1664 0 -1 1188
box 8 4 12 24
use welltap_svt  __well_tap__45
timestamp 1730814361
transform 1 0 1624 0 1 1164
box 8 4 12 24
use welltap_svt  __well_tap__170
timestamp 1730814361
transform 1 0 1664 0 -1 1188
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5981_6
timestamp 1730814361
transform 1 0 2240 0 -1 1192
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5981_6
timestamp 1730814361
transform 1 0 2240 0 -1 1192
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5982_6
timestamp 1730814361
transform 1 0 2392 0 -1 1192
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5982_6
timestamp 1730814361
transform 1 0 2392 0 -1 1192
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5983_6
timestamp 1730814361
transform 1 0 2544 0 -1 1192
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5983_6
timestamp 1730814361
transform 1 0 2544 0 -1 1192
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5393_6
timestamp 1730814361
transform 1 0 2688 0 -1 1192
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5393_6
timestamp 1730814361
transform 1 0 2688 0 -1 1192
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5394_6
timestamp 1730814361
transform 1 0 2840 0 -1 1192
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5394_6
timestamp 1730814361
transform 1 0 2840 0 -1 1192
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5395_6
timestamp 1730814361
transform 1 0 2992 0 -1 1192
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5395_6
timestamp 1730814361
transform 1 0 2992 0 -1 1192
box 7 3 20 38
use welltap_svt  __well_tap__171
timestamp 1730814361
transform 1 0 3184 0 -1 1188
box 8 4 12 24
use welltap_svt  __well_tap__171
timestamp 1730814361
transform 1 0 3184 0 -1 1188
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5745_6
timestamp 1730814361
transform 1 0 128 0 -1 1248
box 7 3 20 38
use welltap_svt  __well_tap__46
timestamp 1730814361
transform 1 0 104 0 -1 1244
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5745_6
timestamp 1730814361
transform 1 0 128 0 -1 1248
box 7 3 20 38
use welltap_svt  __well_tap__46
timestamp 1730814361
transform 1 0 104 0 -1 1244
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5746_6
timestamp 1730814361
transform 1 0 224 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5746_6
timestamp 1730814361
transform 1 0 224 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5747_6
timestamp 1730814361
transform 1 0 352 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5747_6
timestamp 1730814361
transform 1 0 352 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5748_6
timestamp 1730814361
transform 1 0 496 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5748_6
timestamp 1730814361
transform 1 0 496 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5969_6
timestamp 1730814361
transform 1 0 656 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5969_6
timestamp 1730814361
transform 1 0 656 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5986_6
timestamp 1730814361
transform 1 0 824 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5986_6
timestamp 1730814361
transform 1 0 824 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5987_6
timestamp 1730814361
transform 1 0 1008 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5987_6
timestamp 1730814361
transform 1 0 1008 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5988_6
timestamp 1730814361
transform 1 0 1200 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5988_6
timestamp 1730814361
transform 1 0 1200 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5795_6
timestamp 1730814361
transform 1 0 1400 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5795_6
timestamp 1730814361
transform 1 0 1400 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5796_6
timestamp 1730814361
transform 1 0 1592 0 -1 1248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5796_6
timestamp 1730814361
transform 1 0 1592 0 -1 1248
box 7 3 20 38
use welltap_svt  __well_tap__47
timestamp 1730814361
transform 1 0 1624 0 -1 1244
box 8 4 12 24
use welltap_svt  __well_tap__172
timestamp 1730814361
transform 1 0 1664 0 1 1200
box 8 4 12 24
use welltap_svt  __well_tap__47
timestamp 1730814361
transform 1 0 1624 0 -1 1244
box 8 4 12 24
use welltap_svt  __well_tap__172
timestamp 1730814361
transform 1 0 1664 0 1 1200
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5781_6
timestamp 1730814361
transform 1 0 1688 0 1 1196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5781_6
timestamp 1730814361
transform 1 0 1688 0 1 1196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5984_6
timestamp 1730814361
transform 1 0 1976 0 1 1196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5984_6
timestamp 1730814361
transform 1 0 1976 0 1 1196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5398_6
timestamp 1730814361
transform 1 0 2248 0 1 1196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5398_6
timestamp 1730814361
transform 1 0 2248 0 1 1196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5396_6
timestamp 1730814361
transform 1 0 2488 0 1 1196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5396_6
timestamp 1730814361
transform 1 0 2488 0 1 1196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5399_6
timestamp 1730814361
transform 1 0 2704 0 1 1196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5399_6
timestamp 1730814361
transform 1 0 2704 0 1 1196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5397_6
timestamp 1730814361
transform 1 0 2912 0 1 1196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5397_6
timestamp 1730814361
transform 1 0 2912 0 1 1196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5291_6
timestamp 1730814361
transform 1 0 3128 0 1 1196
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5291_6
timestamp 1730814361
transform 1 0 3128 0 1 1196
box 7 3 20 38
use welltap_svt  __well_tap__173
timestamp 1730814361
transform 1 0 3184 0 1 1200
box 8 4 12 24
use welltap_svt  __well_tap__173
timestamp 1730814361
transform 1 0 3184 0 1 1200
box 8 4 12 24
use welltap_svt  __well_tap__48
timestamp 1730814361
transform 1 0 104 0 1 1264
box 8 4 12 24
use welltap_svt  __well_tap__48
timestamp 1730814361
transform 1 0 104 0 1 1264
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5749_6
timestamp 1730814361
transform 1 0 168 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5749_6
timestamp 1730814361
transform 1 0 168 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5704_6
timestamp 1730814361
transform 1 0 296 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5704_6
timestamp 1730814361
transform 1 0 296 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5689_6
timestamp 1730814361
transform 1 0 416 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5689_6
timestamp 1730814361
transform 1 0 416 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5690_6
timestamp 1730814361
transform 1 0 536 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5690_6
timestamp 1730814361
transform 1 0 536 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5989_6
timestamp 1730814361
transform 1 0 656 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5989_6
timestamp 1730814361
transform 1 0 656 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5990_6
timestamp 1730814361
transform 1 0 768 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5990_6
timestamp 1730814361
transform 1 0 768 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5991_6
timestamp 1730814361
transform 1 0 880 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5991_6
timestamp 1730814361
transform 1 0 880 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5992_6
timestamp 1730814361
transform 1 0 1000 0 1 1260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5992_6
timestamp 1730814361
transform 1 0 1000 0 1 1260
box 7 3 20 38
use welltap_svt  __well_tap__49
timestamp 1730814361
transform 1 0 1624 0 1 1264
box 8 4 12 24
use welltap_svt  __well_tap__174
timestamp 1730814361
transform 1 0 1664 0 -1 1288
box 8 4 12 24
use welltap_svt  __well_tap__176
timestamp 1730814361
transform 1 0 1664 0 1 1304
box 8 4 12 24
use welltap_svt  __well_tap__49
timestamp 1730814361
transform 1 0 1624 0 1 1264
box 8 4 12 24
use welltap_svt  __well_tap__174
timestamp 1730814361
transform 1 0 1664 0 -1 1288
box 8 4 12 24
use welltap_svt  __well_tap__176
timestamp 1730814361
transform 1 0 1664 0 1 1304
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5798_6
timestamp 1730814361
transform 1 0 1688 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5798_6
timestamp 1730814361
transform 1 0 1688 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5799_6
timestamp 1730814361
transform 1 0 1784 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5802_6
timestamp 1730814361
transform 1 0 1768 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5799_6
timestamp 1730814361
transform 1 0 1784 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5802_6
timestamp 1730814361
transform 1 0 1768 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5800_6
timestamp 1730814361
transform 1 0 1928 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5803_6
timestamp 1730814361
transform 1 0 1880 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5800_6
timestamp 1730814361
transform 1 0 1928 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5803_6
timestamp 1730814361
transform 1 0 1880 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5804_6
timestamp 1730814361
transform 1 0 1984 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5804_6
timestamp 1730814361
transform 1 0 1984 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5801_6
timestamp 1730814361
transform 1 0 2096 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5805_6
timestamp 1730814361
transform 1 0 2088 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5801_6
timestamp 1730814361
transform 1 0 2096 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5805_6
timestamp 1730814361
transform 1 0 2088 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5404_6
timestamp 1730814361
transform 1 0 2192 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5404_6
timestamp 1730814361
transform 1 0 2192 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5401_6
timestamp 1730814361
transform 1 0 2288 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5405_6
timestamp 1730814361
transform 1 0 2296 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5401_6
timestamp 1730814361
transform 1 0 2288 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5405_6
timestamp 1730814361
transform 1 0 2296 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5485_6
timestamp 1730814361
transform 1 0 2400 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5485_6
timestamp 1730814361
transform 1 0 2400 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5402_6
timestamp 1730814361
transform 1 0 2488 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5402_6
timestamp 1730814361
transform 1 0 2488 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5470_6
timestamp 1730814361
transform 1 0 2504 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5470_6
timestamp 1730814361
transform 1 0 2504 0 1 1300
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5403_6
timestamp 1730814361
transform 1 0 2704 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5403_6
timestamp 1730814361
transform 1 0 2704 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5400_6
timestamp 1730814361
transform 1 0 2928 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5400_6
timestamp 1730814361
transform 1 0 2928 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5292_6
timestamp 1730814361
transform 1 0 3152 0 -1 1292
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5292_6
timestamp 1730814361
transform 1 0 3152 0 -1 1292
box 7 3 20 38
use welltap_svt  __well_tap__175
timestamp 1730814361
transform 1 0 3184 0 -1 1288
box 8 4 12 24
use welltap_svt  __well_tap__177
timestamp 1730814361
transform 1 0 3184 0 1 1304
box 8 4 12 24
use welltap_svt  __well_tap__175
timestamp 1730814361
transform 1 0 3184 0 -1 1288
box 8 4 12 24
use welltap_svt  __well_tap__177
timestamp 1730814361
transform 1 0 3184 0 1 1304
box 8 4 12 24
use welltap_svt  __well_tap__50
timestamp 1730814361
transform 1 0 104 0 -1 1348
box 8 4 12 24
use welltap_svt  __well_tap__52
timestamp 1730814361
transform 1 0 104 0 1 1364
box 8 4 12 24
use welltap_svt  __well_tap__50
timestamp 1730814361
transform 1 0 104 0 -1 1348
box 8 4 12 24
use welltap_svt  __well_tap__52
timestamp 1730814361
transform 1 0 104 0 1 1364
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5691_6
timestamp 1730814361
transform 1 0 264 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5691_6
timestamp 1730814361
transform 1 0 264 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5695_6
timestamp 1730814361
transform 1 0 368 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5695_6
timestamp 1730814361
transform 1 0 368 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5692_6
timestamp 1730814361
transform 1 0 392 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5692_6
timestamp 1730814361
transform 1 0 392 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5696_6
timestamp 1730814361
transform 1 0 496 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5696_6
timestamp 1730814361
transform 1 0 496 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5693_6
timestamp 1730814361
transform 1 0 520 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5693_6
timestamp 1730814361
transform 1 0 520 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5697_6
timestamp 1730814361
transform 1 0 616 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5697_6
timestamp 1730814361
transform 1 0 616 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5694_6
timestamp 1730814361
transform 1 0 640 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5694_6
timestamp 1730814361
transform 1 0 640 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5698_6
timestamp 1730814361
transform 1 0 736 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5698_6
timestamp 1730814361
transform 1 0 736 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5993_6
timestamp 1730814361
transform 1 0 760 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5993_6
timestamp 1730814361
transform 1 0 760 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5994_6
timestamp 1730814361
transform 1 0 872 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5997_6
timestamp 1730814361
transform 1 0 856 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5994_6
timestamp 1730814361
transform 1 0 872 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5997_6
timestamp 1730814361
transform 1 0 856 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5995_6
timestamp 1730814361
transform 1 0 984 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5998_6
timestamp 1730814361
transform 1 0 968 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5995_6
timestamp 1730814361
transform 1 0 984 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5998_6
timestamp 1730814361
transform 1 0 968 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5996_6
timestamp 1730814361
transform 1 0 1104 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5999_6
timestamp 1730814361
transform 1 0 1088 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5996_6
timestamp 1730814361
transform 1 0 1104 0 -1 1352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5999_6
timestamp 1730814361
transform 1 0 1088 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5954_6
timestamp 1730814361
transform 1 0 1208 0 1 1360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5954_6
timestamp 1730814361
transform 1 0 1208 0 1 1360
box 7 3 20 38
use welltap_svt  __well_tap__51
timestamp 1730814361
transform 1 0 1624 0 -1 1348
box 8 4 12 24
use welltap_svt  __well_tap__53
timestamp 1730814361
transform 1 0 1624 0 1 1364
box 8 4 12 24
use welltap_svt  __well_tap__178
timestamp 1730814361
transform 1 0 1664 0 -1 1388
box 8 4 12 24
use welltap_svt  __well_tap__51
timestamp 1730814361
transform 1 0 1624 0 -1 1348
box 8 4 12 24
use welltap_svt  __well_tap__53
timestamp 1730814361
transform 1 0 1624 0 1 1364
box 8 4 12 24
use welltap_svt  __well_tap__178
timestamp 1730814361
transform 1 0 1664 0 -1 1388
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5806_6
timestamp 1730814361
transform 1 0 1872 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5806_6
timestamp 1730814361
transform 1 0 1872 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5807_6
timestamp 1730814361
transform 1 0 1984 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5807_6
timestamp 1730814361
transform 1 0 1984 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5808_6
timestamp 1730814361
transform 1 0 2096 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5808_6
timestamp 1730814361
transform 1 0 2096 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5809_6
timestamp 1730814361
transform 1 0 2232 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5809_6
timestamp 1730814361
transform 1 0 2232 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5471_6
timestamp 1730814361
transform 1 0 2384 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5471_6
timestamp 1730814361
transform 1 0 2384 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5472_6
timestamp 1730814361
transform 1 0 2560 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5472_6
timestamp 1730814361
transform 1 0 2560 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5473_6
timestamp 1730814361
transform 1 0 2760 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5473_6
timestamp 1730814361
transform 1 0 2760 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5474_6
timestamp 1730814361
transform 1 0 2968 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5474_6
timestamp 1730814361
transform 1 0 2968 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5293_6
timestamp 1730814361
transform 1 0 3152 0 -1 1392
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5293_6
timestamp 1730814361
transform 1 0 3152 0 -1 1392
box 7 3 20 38
use welltap_svt  __well_tap__179
timestamp 1730814361
transform 1 0 3184 0 -1 1388
box 8 4 12 24
use welltap_svt  __well_tap__179
timestamp 1730814361
transform 1 0 3184 0 -1 1388
box 8 4 12 24
use welltap_svt  __well_tap__54
timestamp 1730814361
transform 1 0 104 0 -1 1448
box 8 4 12 24
use welltap_svt  __well_tap__54
timestamp 1730814361
transform 1 0 104 0 -1 1448
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5699_6
timestamp 1730814361
transform 1 0 472 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5699_6
timestamp 1730814361
transform 1 0 472 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5700_6
timestamp 1730814361
transform 1 0 600 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5700_6
timestamp 1730814361
transform 1 0 600 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5701_6
timestamp 1730814361
transform 1 0 720 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5701_6
timestamp 1730814361
transform 1 0 720 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5702_6
timestamp 1730814361
transform 1 0 840 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5702_6
timestamp 1730814361
transform 1 0 840 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5939_6
timestamp 1730814361
transform 1 0 960 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5939_6
timestamp 1730814361
transform 1 0 960 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5940_6
timestamp 1730814361
transform 1 0 1072 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5940_6
timestamp 1730814361
transform 1 0 1072 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5941_6
timestamp 1730814361
transform 1 0 1184 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5941_6
timestamp 1730814361
transform 1 0 1184 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5942_6
timestamp 1730814361
transform 1 0 1304 0 -1 1452
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5942_6
timestamp 1730814361
transform 1 0 1304 0 -1 1452
box 7 3 20 38
use welltap_svt  __well_tap__55
timestamp 1730814361
transform 1 0 1624 0 -1 1448
box 8 4 12 24
use welltap_svt  __well_tap__180
timestamp 1730814361
transform 1 0 1664 0 1 1412
box 8 4 12 24
use welltap_svt  __well_tap__55
timestamp 1730814361
transform 1 0 1624 0 -1 1448
box 8 4 12 24
use welltap_svt  __well_tap__180
timestamp 1730814361
transform 1 0 1664 0 1 1412
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5810_6
timestamp 1730814361
transform 1 0 1976 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5810_6
timestamp 1730814361
transform 1 0 1976 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5811_6
timestamp 1730814361
transform 1 0 2088 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5811_6
timestamp 1730814361
transform 1 0 2088 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5812_6
timestamp 1730814361
transform 1 0 2200 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5812_6
timestamp 1730814361
transform 1 0 2200 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5766_6
timestamp 1730814361
transform 1 0 2328 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5766_6
timestamp 1730814361
transform 1 0 2328 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5475_6
timestamp 1730814361
transform 1 0 2472 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5475_6
timestamp 1730814361
transform 1 0 2472 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5476_6
timestamp 1730814361
transform 1 0 2632 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5476_6
timestamp 1730814361
transform 1 0 2632 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5477_6
timestamp 1730814361
transform 1 0 2808 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5477_6
timestamp 1730814361
transform 1 0 2808 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5478_6
timestamp 1730814361
transform 1 0 2992 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5478_6
timestamp 1730814361
transform 1 0 2992 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5294_6
timestamp 1730814361
transform 1 0 3152 0 1 1408
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5294_6
timestamp 1730814361
transform 1 0 3152 0 1 1408
box 7 3 20 38
use welltap_svt  __well_tap__181
timestamp 1730814361
transform 1 0 3184 0 1 1412
box 8 4 12 24
use welltap_svt  __well_tap__181
timestamp 1730814361
transform 1 0 3184 0 1 1412
box 8 4 12 24
use welltap_svt  __well_tap__56
timestamp 1730814361
transform 1 0 104 0 1 1468
box 8 4 12 24
use welltap_svt  __well_tap__56
timestamp 1730814361
transform 1 0 104 0 1 1468
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5703_6
timestamp 1730814361
transform 1 0 568 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5703_6
timestamp 1730814361
transform 1 0 568 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5625_6
timestamp 1730814361
transform 1 0 696 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5625_6
timestamp 1730814361
transform 1 0 696 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5705_6
timestamp 1730814361
transform 1 0 824 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5705_6
timestamp 1730814361
transform 1 0 824 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5706_6
timestamp 1730814361
transform 1 0 944 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5706_6
timestamp 1730814361
transform 1 0 944 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5943_6
timestamp 1730814361
transform 1 0 1064 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5943_6
timestamp 1730814361
transform 1 0 1064 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5944_6
timestamp 1730814361
transform 1 0 1176 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5944_6
timestamp 1730814361
transform 1 0 1176 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5945_6
timestamp 1730814361
transform 1 0 1288 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5945_6
timestamp 1730814361
transform 1 0 1288 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5946_6
timestamp 1730814361
transform 1 0 1408 0 1 1464
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5946_6
timestamp 1730814361
transform 1 0 1408 0 1 1464
box 7 3 20 38
use welltap_svt  __well_tap__57
timestamp 1730814361
transform 1 0 1624 0 1 1468
box 8 4 12 24
use welltap_svt  __well_tap__182
timestamp 1730814361
transform 1 0 1664 0 -1 1488
box 8 4 12 24
use welltap_svt  __well_tap__57
timestamp 1730814361
transform 1 0 1624 0 1 1468
box 8 4 12 24
use welltap_svt  __well_tap__182
timestamp 1730814361
transform 1 0 1664 0 -1 1488
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5751_6
timestamp 1730814361
transform 1 0 2080 0 -1 1492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5751_6
timestamp 1730814361
transform 1 0 2080 0 -1 1492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5752_6
timestamp 1730814361
transform 1 0 2224 0 -1 1492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5752_6
timestamp 1730814361
transform 1 0 2224 0 -1 1492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5753_6
timestamp 1730814361
transform 1 0 2368 0 -1 1492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5753_6
timestamp 1730814361
transform 1 0 2368 0 -1 1492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5479_6
timestamp 1730814361
transform 1 0 2504 0 -1 1492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5479_6
timestamp 1730814361
transform 1 0 2504 0 -1 1492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5480_6
timestamp 1730814361
transform 1 0 2648 0 -1 1492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5480_6
timestamp 1730814361
transform 1 0 2648 0 -1 1492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5481_6
timestamp 1730814361
transform 1 0 2792 0 -1 1492
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5481_6
timestamp 1730814361
transform 1 0 2792 0 -1 1492
box 7 3 20 38
use welltap_svt  __well_tap__183
timestamp 1730814361
transform 1 0 3184 0 -1 1488
box 8 4 12 24
use welltap_svt  __well_tap__183
timestamp 1730814361
transform 1 0 3184 0 -1 1488
box 8 4 12 24
use welltap_svt  __well_tap__58
timestamp 1730814361
transform 1 0 104 0 -1 1548
box 8 4 12 24
use welltap_svt  __well_tap__58
timestamp 1730814361
transform 1 0 104 0 -1 1548
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5707_6
timestamp 1730814361
transform 1 0 672 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5707_6
timestamp 1730814361
transform 1 0 672 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5708_6
timestamp 1730814361
transform 1 0 800 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5708_6
timestamp 1730814361
transform 1 0 800 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5709_6
timestamp 1730814361
transform 1 0 920 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5709_6
timestamp 1730814361
transform 1 0 920 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5710_6
timestamp 1730814361
transform 1 0 1040 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5710_6
timestamp 1730814361
transform 1 0 1040 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5947_6
timestamp 1730814361
transform 1 0 1160 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5947_6
timestamp 1730814361
transform 1 0 1160 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5948_6
timestamp 1730814361
transform 1 0 1272 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5948_6
timestamp 1730814361
transform 1 0 1272 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5949_6
timestamp 1730814361
transform 1 0 1392 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5949_6
timestamp 1730814361
transform 1 0 1392 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5950_6
timestamp 1730814361
transform 1 0 1512 0 -1 1552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5950_6
timestamp 1730814361
transform 1 0 1512 0 -1 1552
box 7 3 20 38
use welltap_svt  __well_tap__59
timestamp 1730814361
transform 1 0 1624 0 -1 1548
box 8 4 12 24
use welltap_svt  __well_tap__184
timestamp 1730814361
transform 1 0 1664 0 1 1500
box 8 4 12 24
use welltap_svt  __well_tap__186
timestamp 1730814361
transform 1 0 1664 0 -1 1580
box 8 4 12 24
use welltap_svt  __well_tap__59
timestamp 1730814361
transform 1 0 1624 0 -1 1548
box 8 4 12 24
use welltap_svt  __well_tap__184
timestamp 1730814361
transform 1 0 1664 0 1 1500
box 8 4 12 24
use welltap_svt  __well_tap__186
timestamp 1730814361
transform 1 0 1664 0 -1 1580
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5754_6
timestamp 1730814361
transform 1 0 2160 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5754_6
timestamp 1730814361
transform 1 0 2160 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5755_6
timestamp 1730814361
transform 1 0 2272 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5758_6
timestamp 1730814361
transform 1 0 2264 0 -1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5755_6
timestamp 1730814361
transform 1 0 2272 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5758_6
timestamp 1730814361
transform 1 0 2264 0 -1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5756_6
timestamp 1730814361
transform 1 0 2384 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5759_6
timestamp 1730814361
transform 1 0 2408 0 -1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5756_6
timestamp 1730814361
transform 1 0 2384 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5759_6
timestamp 1730814361
transform 1 0 2408 0 -1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5757_6
timestamp 1730814361
transform 1 0 2496 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5760_6
timestamp 1730814361
transform 1 0 2552 0 -1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5757_6
timestamp 1730814361
transform 1 0 2496 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5760_6
timestamp 1730814361
transform 1 0 2552 0 -1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5482_6
timestamp 1730814361
transform 1 0 2608 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5482_6
timestamp 1730814361
transform 1 0 2608 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5483_6
timestamp 1730814361
transform 1 0 2728 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5486_6
timestamp 1730814361
transform 1 0 2688 0 -1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5483_6
timestamp 1730814361
transform 1 0 2728 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5486_6
timestamp 1730814361
transform 1 0 2688 0 -1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5484_6
timestamp 1730814361
transform 1 0 2848 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5487_6
timestamp 1730814361
transform 1 0 2832 0 -1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5484_6
timestamp 1730814361
transform 1 0 2848 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5487_6
timestamp 1730814361
transform 1 0 2832 0 -1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5469_6
timestamp 1730814361
transform 1 0 2976 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5488_6
timestamp 1730814361
transform 1 0 2976 0 -1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5469_6
timestamp 1730814361
transform 1 0 2976 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5488_6
timestamp 1730814361
transform 1 0 2976 0 -1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5493_6
timestamp 1730814361
transform 1 0 3104 0 1 1496
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5493_6
timestamp 1730814361
transform 1 0 3104 0 1 1496
box 7 3 20 38
use welltap_svt  __well_tap__185
timestamp 1730814361
transform 1 0 3184 0 1 1500
box 8 4 12 24
use welltap_svt  __well_tap__187
timestamp 1730814361
transform 1 0 3184 0 -1 1580
box 8 4 12 24
use welltap_svt  __well_tap__185
timestamp 1730814361
transform 1 0 3184 0 1 1500
box 8 4 12 24
use welltap_svt  __well_tap__187
timestamp 1730814361
transform 1 0 3184 0 -1 1580
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5713_6
timestamp 1730814361
transform 1 0 128 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5715_6
timestamp 1730814361
transform 1 0 128 0 -1 1652
box 7 3 20 38
use welltap_svt  __well_tap__60
timestamp 1730814361
transform 1 0 104 0 1 1568
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5713_6
timestamp 1730814361
transform 1 0 128 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5715_6
timestamp 1730814361
transform 1 0 128 0 -1 1652
box 7 3 20 38
use welltap_svt  __well_tap__60
timestamp 1730814361
transform 1 0 104 0 1 1568
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5716_6
timestamp 1730814361
transform 1 0 240 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5716_6
timestamp 1730814361
transform 1 0 240 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5714_6
timestamp 1730814361
transform 1 0 296 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5714_6
timestamp 1730814361
transform 1 0 296 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5717_6
timestamp 1730814361
transform 1 0 376 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5717_6
timestamp 1730814361
transform 1 0 376 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5711_6
timestamp 1730814361
transform 1 0 496 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5711_6
timestamp 1730814361
transform 1 0 496 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5718_6
timestamp 1730814361
transform 1 0 528 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5718_6
timestamp 1730814361
transform 1 0 528 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5712_6
timestamp 1730814361
transform 1 0 688 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5712_6
timestamp 1730814361
transform 1 0 688 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5955_6
timestamp 1730814361
transform 1 0 704 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5955_6
timestamp 1730814361
transform 1 0 704 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5953_6
timestamp 1730814361
transform 1 0 880 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5956_6
timestamp 1730814361
transform 1 0 912 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5953_6
timestamp 1730814361
transform 1 0 880 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5956_6
timestamp 1730814361
transform 1 0 912 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5875_6
timestamp 1730814361
transform 1 0 1056 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5875_6
timestamp 1730814361
transform 1 0 1056 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5957_6
timestamp 1730814361
transform 1 0 1136 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5957_6
timestamp 1730814361
transform 1 0 1136 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5951_6
timestamp 1730814361
transform 1 0 1232 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5951_6
timestamp 1730814361
transform 1 0 1232 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5952_6
timestamp 1730814361
transform 1 0 1408 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5958_6
timestamp 1730814361
transform 1 0 1376 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5952_6
timestamp 1730814361
transform 1 0 1408 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5958_6
timestamp 1730814361
transform 1 0 1376 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5762_6
timestamp 1730814361
transform 1 0 1584 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5763_6
timestamp 1730814361
transform 1 0 1592 0 -1 1652
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5762_6
timestamp 1730814361
transform 1 0 1584 0 1 1564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5763_6
timestamp 1730814361
transform 1 0 1592 0 -1 1652
box 7 3 20 38
use welltap_svt  __well_tap__61
timestamp 1730814361
transform 1 0 1624 0 1 1568
box 8 4 12 24
use welltap_svt  __well_tap__188
timestamp 1730814361
transform 1 0 1664 0 1 1588
box 8 4 12 24
use welltap_svt  __well_tap__61
timestamp 1730814361
transform 1 0 1624 0 1 1568
box 8 4 12 24
use welltap_svt  __well_tap__188
timestamp 1730814361
transform 1 0 1664 0 1 1588
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5494_6
timestamp 1730814361
transform 1 0 2312 0 1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5494_6
timestamp 1730814361
transform 1 0 2312 0 1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5489_6
timestamp 1730814361
transform 1 0 2512 0 1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5489_6
timestamp 1730814361
transform 1 0 2512 0 1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5490_6
timestamp 1730814361
transform 1 0 2704 0 1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5490_6
timestamp 1730814361
transform 1 0 2704 0 1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5491_6
timestamp 1730814361
transform 1 0 2904 0 1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5491_6
timestamp 1730814361
transform 1 0 2904 0 1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5295_6
timestamp 1730814361
transform 1 0 3104 0 1 1584
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5295_6
timestamp 1730814361
transform 1 0 3104 0 1 1584
box 7 3 20 38
use welltap_svt  __well_tap__189
timestamp 1730814361
transform 1 0 3184 0 1 1588
box 8 4 12 24
use welltap_svt  __well_tap__189
timestamp 1730814361
transform 1 0 3184 0 1 1588
box 8 4 12 24
use welltap_svt  __well_tap__62
timestamp 1730814361
transform 1 0 104 0 -1 1648
box 8 4 12 24
use welltap_svt  __well_tap__64
timestamp 1730814361
transform 1 0 104 0 1 1668
box 8 4 12 24
use welltap_svt  __well_tap__62
timestamp 1730814361
transform 1 0 104 0 -1 1648
box 8 4 12 24
use welltap_svt  __well_tap__64
timestamp 1730814361
transform 1 0 104 0 1 1668
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5547_6
timestamp 1730814361
transform 1 0 216 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5547_6
timestamp 1730814361
transform 1 0 216 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5532_6
timestamp 1730814361
transform 1 0 344 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5532_6
timestamp 1730814361
transform 1 0 344 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5533_6
timestamp 1730814361
transform 1 0 464 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5533_6
timestamp 1730814361
transform 1 0 464 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5534_6
timestamp 1730814361
transform 1 0 584 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5534_6
timestamp 1730814361
transform 1 0 584 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5959_6
timestamp 1730814361
transform 1 0 704 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5959_6
timestamp 1730814361
transform 1 0 704 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5960_6
timestamp 1730814361
transform 1 0 816 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5960_6
timestamp 1730814361
transform 1 0 816 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5961_6
timestamp 1730814361
transform 1 0 936 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5961_6
timestamp 1730814361
transform 1 0 936 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5962_6
timestamp 1730814361
transform 1 0 1056 0 1 1664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5962_6
timestamp 1730814361
transform 1 0 1056 0 1 1664
box 7 3 20 38
use welltap_svt  __well_tap__63
timestamp 1730814361
transform 1 0 1624 0 -1 1648
box 8 4 12 24
use welltap_svt  __well_tap__65
timestamp 1730814361
transform 1 0 1624 0 1 1668
box 8 4 12 24
use welltap_svt  __well_tap__190
timestamp 1730814361
transform 1 0 1664 0 -1 1664
box 8 4 12 24
use welltap_svt  __well_tap__192
timestamp 1730814361
transform 1 0 1664 0 1 1672
box 8 4 12 24
use welltap_svt  __well_tap__63
timestamp 1730814361
transform 1 0 1624 0 -1 1648
box 8 4 12 24
use welltap_svt  __well_tap__65
timestamp 1730814361
transform 1 0 1624 0 1 1668
box 8 4 12 24
use welltap_svt  __well_tap__190
timestamp 1730814361
transform 1 0 1664 0 -1 1664
box 8 4 12 24
use welltap_svt  __well_tap__192
timestamp 1730814361
transform 1 0 1664 0 1 1672
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5764_6
timestamp 1730814361
transform 1 0 1688 0 -1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5767_6
timestamp 1730814361
transform 1 0 1728 0 1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5764_6
timestamp 1730814361
transform 1 0 1688 0 -1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5767_6
timestamp 1730814361
transform 1 0 1728 0 1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5765_6
timestamp 1730814361
transform 1 0 1888 0 -1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5768_6
timestamp 1730814361
transform 1 0 1872 0 1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5765_6
timestamp 1730814361
transform 1 0 1888 0 -1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5768_6
timestamp 1730814361
transform 1 0 1872 0 1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5769_6
timestamp 1730814361
transform 1 0 2016 0 1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5769_6
timestamp 1730814361
transform 1 0 2016 0 1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5496_6
timestamp 1730814361
transform 1 0 2160 0 1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5813_6
timestamp 1730814361
transform 1 0 2120 0 -1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5496_6
timestamp 1730814361
transform 1 0 2160 0 1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5813_6
timestamp 1730814361
transform 1 0 2120 0 -1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5497_6
timestamp 1730814361
transform 1 0 2304 0 1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5497_6
timestamp 1730814361
transform 1 0 2304 0 1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5761_6
timestamp 1730814361
transform 1 0 2360 0 -1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5761_6
timestamp 1730814361
transform 1 0 2360 0 -1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5498_6
timestamp 1730814361
transform 1 0 2456 0 1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5498_6
timestamp 1730814361
transform 1 0 2456 0 1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5495_6
timestamp 1730814361
transform 1 0 2608 0 -1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5495_6
timestamp 1730814361
transform 1 0 2608 0 -1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5492_6
timestamp 1730814361
transform 1 0 2864 0 -1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5492_6
timestamp 1730814361
transform 1 0 2864 0 -1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5296_6
timestamp 1730814361
transform 1 0 3128 0 -1 1668
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5296_6
timestamp 1730814361
transform 1 0 3128 0 -1 1668
box 7 3 20 38
use welltap_svt  __well_tap__191
timestamp 1730814361
transform 1 0 3184 0 -1 1664
box 8 4 12 24
use welltap_svt  __well_tap__193
timestamp 1730814361
transform 1 0 3184 0 1 1672
box 8 4 12 24
use welltap_svt  __well_tap__191
timestamp 1730814361
transform 1 0 3184 0 -1 1664
box 8 4 12 24
use welltap_svt  __well_tap__193
timestamp 1730814361
transform 1 0 3184 0 1 1672
box 8 4 12 24
use welltap_svt  __well_tap__66
timestamp 1730814361
transform 1 0 104 0 -1 1752
box 8 4 12 24
use welltap_svt  __well_tap__66
timestamp 1730814361
transform 1 0 104 0 -1 1752
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5535_6
timestamp 1730814361
transform 1 0 320 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5535_6
timestamp 1730814361
transform 1 0 320 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5536_6
timestamp 1730814361
transform 1 0 448 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5536_6
timestamp 1730814361
transform 1 0 448 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5537_6
timestamp 1730814361
transform 1 0 568 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5537_6
timestamp 1730814361
transform 1 0 568 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5538_6
timestamp 1730814361
transform 1 0 688 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5538_6
timestamp 1730814361
transform 1 0 688 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5963_6
timestamp 1730814361
transform 1 0 808 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5963_6
timestamp 1730814361
transform 1 0 808 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5964_6
timestamp 1730814361
transform 1 0 920 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5964_6
timestamp 1730814361
transform 1 0 920 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5965_6
timestamp 1730814361
transform 1 0 1032 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5965_6
timestamp 1730814361
transform 1 0 1032 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5966_6
timestamp 1730814361
transform 1 0 1152 0 -1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5966_6
timestamp 1730814361
transform 1 0 1152 0 -1 1756
box 7 3 20 38
use welltap_svt  __well_tap__67
timestamp 1730814361
transform 1 0 1624 0 -1 1752
box 8 4 12 24
use welltap_svt  __well_tap__194
timestamp 1730814361
transform 1 0 1664 0 -1 1744
box 8 4 12 24
use welltap_svt  __well_tap__67
timestamp 1730814361
transform 1 0 1624 0 -1 1752
box 8 4 12 24
use welltap_svt  __well_tap__194
timestamp 1730814361
transform 1 0 1664 0 -1 1744
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5770_6
timestamp 1730814361
transform 1 0 1808 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5770_6
timestamp 1730814361
transform 1 0 1808 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5771_6
timestamp 1730814361
transform 1 0 1960 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5771_6
timestamp 1730814361
transform 1 0 1960 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5772_6
timestamp 1730814361
transform 1 0 2120 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5772_6
timestamp 1730814361
transform 1 0 2120 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5499_6
timestamp 1730814361
transform 1 0 2296 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5499_6
timestamp 1730814361
transform 1 0 2296 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5454_6
timestamp 1730814361
transform 1 0 2496 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5454_6
timestamp 1730814361
transform 1 0 2496 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5439_6
timestamp 1730814361
transform 1 0 2704 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5439_6
timestamp 1730814361
transform 1 0 2704 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5440_6
timestamp 1730814361
transform 1 0 2928 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5440_6
timestamp 1730814361
transform 1 0 2928 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5281_6
timestamp 1730814361
transform 1 0 3152 0 -1 1748
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5281_6
timestamp 1730814361
transform 1 0 3152 0 -1 1748
box 7 3 20 38
use welltap_svt  __well_tap__195
timestamp 1730814361
transform 1 0 3184 0 -1 1744
box 8 4 12 24
use welltap_svt  __well_tap__195
timestamp 1730814361
transform 1 0 3184 0 -1 1744
box 8 4 12 24
use welltap_svt  __well_tap__68
timestamp 1730814361
transform 1 0 104 0 1 1772
box 8 4 12 24
use welltap_svt  __well_tap__68
timestamp 1730814361
transform 1 0 104 0 1 1772
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5539_6
timestamp 1730814361
transform 1 0 416 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5539_6
timestamp 1730814361
transform 1 0 416 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5540_6
timestamp 1730814361
transform 1 0 544 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5540_6
timestamp 1730814361
transform 1 0 544 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5541_6
timestamp 1730814361
transform 1 0 672 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5541_6
timestamp 1730814361
transform 1 0 672 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5542_6
timestamp 1730814361
transform 1 0 792 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5542_6
timestamp 1730814361
transform 1 0 792 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5967_6
timestamp 1730814361
transform 1 0 912 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5967_6
timestamp 1730814361
transform 1 0 912 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5968_6
timestamp 1730814361
transform 1 0 1024 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5968_6
timestamp 1730814361
transform 1 0 1024 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5797_6
timestamp 1730814361
transform 1 0 1136 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5797_6
timestamp 1730814361
transform 1 0 1136 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5782_6
timestamp 1730814361
transform 1 0 1256 0 1 1768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5782_6
timestamp 1730814361
transform 1 0 1256 0 1 1768
box 7 3 20 38
use welltap_svt  __well_tap__69
timestamp 1730814361
transform 1 0 1624 0 1 1772
box 8 4 12 24
use welltap_svt  __well_tap__196
timestamp 1730814361
transform 1 0 1664 0 1 1760
box 8 4 12 24
use welltap_svt  __well_tap__69
timestamp 1730814361
transform 1 0 1624 0 1 1772
box 8 4 12 24
use welltap_svt  __well_tap__196
timestamp 1730814361
transform 1 0 1664 0 1 1760
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5773_6
timestamp 1730814361
transform 1 0 1896 0 1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5773_6
timestamp 1730814361
transform 1 0 1896 0 1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5776_6
timestamp 1730814361
transform 1 0 1976 0 -1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5776_6
timestamp 1730814361
transform 1 0 1976 0 -1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5774_6
timestamp 1730814361
transform 1 0 2072 0 1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5774_6
timestamp 1730814361
transform 1 0 2072 0 1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5777_6
timestamp 1730814361
transform 1 0 2128 0 -1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5777_6
timestamp 1730814361
transform 1 0 2128 0 -1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5775_6
timestamp 1730814361
transform 1 0 2264 0 1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5778_6
timestamp 1730814361
transform 1 0 2280 0 -1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5775_6
timestamp 1730814361
transform 1 0 2264 0 1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5778_6
timestamp 1730814361
transform 1 0 2280 0 -1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5444_6
timestamp 1730814361
transform 1 0 2424 0 -1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5444_6
timestamp 1730814361
transform 1 0 2424 0 -1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5441_6
timestamp 1730814361
transform 1 0 2480 0 1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5441_6
timestamp 1730814361
transform 1 0 2480 0 1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5445_6
timestamp 1730814361
transform 1 0 2576 0 -1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5445_6
timestamp 1730814361
transform 1 0 2576 0 -1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5442_6
timestamp 1730814361
transform 1 0 2704 0 1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5446_6
timestamp 1730814361
transform 1 0 2728 0 -1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5442_6
timestamp 1730814361
transform 1 0 2704 0 1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5446_6
timestamp 1730814361
transform 1 0 2728 0 -1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5443_6
timestamp 1730814361
transform 1 0 2936 0 1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5443_6
timestamp 1730814361
transform 1 0 2936 0 1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5298_6
timestamp 1730814361
transform 1 0 3152 0 1 1756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5298_6
timestamp 1730814361
transform 1 0 3152 0 1 1756
box 7 3 20 38
use welltap_svt  __well_tap__197
timestamp 1730814361
transform 1 0 3184 0 1 1760
box 8 4 12 24
use welltap_svt  __well_tap__197
timestamp 1730814361
transform 1 0 3184 0 1 1760
box 8 4 12 24
use welltap_svt  __well_tap__70
timestamp 1730814361
transform 1 0 104 0 -1 1852
box 8 4 12 24
use welltap_svt  __well_tap__70
timestamp 1730814361
transform 1 0 104 0 -1 1852
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5543_6
timestamp 1730814361
transform 1 0 520 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5543_6
timestamp 1730814361
transform 1 0 520 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5544_6
timestamp 1730814361
transform 1 0 648 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5544_6
timestamp 1730814361
transform 1 0 648 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5545_6
timestamp 1730814361
transform 1 0 768 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5545_6
timestamp 1730814361
transform 1 0 768 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5546_6
timestamp 1730814361
transform 1 0 888 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5546_6
timestamp 1730814361
transform 1 0 888 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5783_6
timestamp 1730814361
transform 1 0 1008 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5783_6
timestamp 1730814361
transform 1 0 1008 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5784_6
timestamp 1730814361
transform 1 0 1120 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5784_6
timestamp 1730814361
transform 1 0 1120 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5785_6
timestamp 1730814361
transform 1 0 1240 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5785_6
timestamp 1730814361
transform 1 0 1240 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5786_6
timestamp 1730814361
transform 1 0 1360 0 -1 1856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5786_6
timestamp 1730814361
transform 1 0 1360 0 -1 1856
box 7 3 20 38
use welltap_svt  __well_tap__71
timestamp 1730814361
transform 1 0 1624 0 -1 1852
box 8 4 12 24
use welltap_svt  __well_tap__198
timestamp 1730814361
transform 1 0 1664 0 -1 1832
box 8 4 12 24
use welltap_svt  __well_tap__200
timestamp 1730814361
transform 1 0 1664 0 1 1840
box 8 4 12 24
use welltap_svt  __well_tap__71
timestamp 1730814361
transform 1 0 1624 0 -1 1852
box 8 4 12 24
use welltap_svt  __well_tap__198
timestamp 1730814361
transform 1 0 1664 0 -1 1832
box 8 4 12 24
use welltap_svt  __well_tap__200
timestamp 1730814361
transform 1 0 1664 0 1 1840
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5779_6
timestamp 1730814361
transform 1 0 2064 0 1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5779_6
timestamp 1730814361
transform 1 0 2064 0 1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5780_6
timestamp 1730814361
transform 1 0 2232 0 1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5780_6
timestamp 1730814361
transform 1 0 2232 0 1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5860_6
timestamp 1730814361
transform 1 0 2408 0 1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5860_6
timestamp 1730814361
transform 1 0 2408 0 1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5447_6
timestamp 1730814361
transform 1 0 2592 0 1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5447_6
timestamp 1730814361
transform 1 0 2592 0 1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5448_6
timestamp 1730814361
transform 1 0 2784 0 1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5448_6
timestamp 1730814361
transform 1 0 2784 0 1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5449_6
timestamp 1730814361
transform 1 0 2976 0 1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5449_6
timestamp 1730814361
transform 1 0 2976 0 1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5299_6
timestamp 1730814361
transform 1 0 3152 0 1 1836
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5299_6
timestamp 1730814361
transform 1 0 3152 0 1 1836
box 7 3 20 38
use welltap_svt  __well_tap__199
timestamp 1730814361
transform 1 0 3184 0 -1 1832
box 8 4 12 24
use welltap_svt  __well_tap__201
timestamp 1730814361
transform 1 0 3184 0 1 1840
box 8 4 12 24
use welltap_svt  __well_tap__199
timestamp 1730814361
transform 1 0 3184 0 -1 1832
box 8 4 12 24
use welltap_svt  __well_tap__201
timestamp 1730814361
transform 1 0 3184 0 1 1840
box 8 4 12 24
use welltap_svt  __well_tap__72
timestamp 1730814361
transform 1 0 104 0 1 1872
box 8 4 12 24
use welltap_svt  __well_tap__72
timestamp 1730814361
transform 1 0 104 0 1 1872
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5531_6
timestamp 1730814361
transform 1 0 624 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5531_6
timestamp 1730814361
transform 1 0 624 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5548_6
timestamp 1730814361
transform 1 0 752 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5551_6
timestamp 1730814361
transform 1 0 720 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5548_6
timestamp 1730814361
transform 1 0 752 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5551_6
timestamp 1730814361
transform 1 0 720 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5549_6
timestamp 1730814361
transform 1 0 872 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5552_6
timestamp 1730814361
transform 1 0 848 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5549_6
timestamp 1730814361
transform 1 0 872 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5552_6
timestamp 1730814361
transform 1 0 848 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5550_6
timestamp 1730814361
transform 1 0 992 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5553_6
timestamp 1730814361
transform 1 0 976 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5550_6
timestamp 1730814361
transform 1 0 992 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5553_6
timestamp 1730814361
transform 1 0 976 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5554_6
timestamp 1730814361
transform 1 0 1096 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5787_6
timestamp 1730814361
transform 1 0 1112 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5554_6
timestamp 1730814361
transform 1 0 1096 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5787_6
timestamp 1730814361
transform 1 0 1112 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5788_6
timestamp 1730814361
transform 1 0 1224 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5791_6
timestamp 1730814361
transform 1 0 1216 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5788_6
timestamp 1730814361
transform 1 0 1224 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5791_6
timestamp 1730814361
transform 1 0 1216 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5789_6
timestamp 1730814361
transform 1 0 1336 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5792_6
timestamp 1730814361
transform 1 0 1328 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5789_6
timestamp 1730814361
transform 1 0 1336 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5792_6
timestamp 1730814361
transform 1 0 1328 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5790_6
timestamp 1730814361
transform 1 0 1456 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5793_6
timestamp 1730814361
transform 1 0 1440 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5790_6
timestamp 1730814361
transform 1 0 1456 0 1 1868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5793_6
timestamp 1730814361
transform 1 0 1440 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5794_6
timestamp 1730814361
transform 1 0 1560 0 -1 1960
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5794_6
timestamp 1730814361
transform 1 0 1560 0 -1 1960
box 7 3 20 38
use welltap_svt  __well_tap__73
timestamp 1730814361
transform 1 0 1624 0 1 1872
box 8 4 12 24
use welltap_svt  __well_tap__202
timestamp 1730814361
transform 1 0 1664 0 -1 1916
box 8 4 12 24
use welltap_svt  __well_tap__73
timestamp 1730814361
transform 1 0 1624 0 1 1872
box 8 4 12 24
use welltap_svt  __well_tap__202
timestamp 1730814361
transform 1 0 1664 0 -1 1916
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5845_6
timestamp 1730814361
transform 1 0 2144 0 -1 1920
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5845_6
timestamp 1730814361
transform 1 0 2144 0 -1 1920
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5848_6
timestamp 1730814361
transform 1 0 2232 0 1 1924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5848_6
timestamp 1730814361
transform 1 0 2232 0 1 1924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5846_6
timestamp 1730814361
transform 1 0 2304 0 -1 1920
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5846_6
timestamp 1730814361
transform 1 0 2304 0 -1 1920
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5849_6
timestamp 1730814361
transform 1 0 2384 0 1 1924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5849_6
timestamp 1730814361
transform 1 0 2384 0 1 1924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5847_6
timestamp 1730814361
transform 1 0 2464 0 -1 1920
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5847_6
timestamp 1730814361
transform 1 0 2464 0 -1 1920
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5850_6
timestamp 1730814361
transform 1 0 2536 0 1 1924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5850_6
timestamp 1730814361
transform 1 0 2536 0 1 1924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5450_6
timestamp 1730814361
transform 1 0 2632 0 -1 1920
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5450_6
timestamp 1730814361
transform 1 0 2632 0 -1 1920
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5453_6
timestamp 1730814361
transform 1 0 2688 0 1 1924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5453_6
timestamp 1730814361
transform 1 0 2688 0 1 1924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5375_6
timestamp 1730814361
transform 1 0 2840 0 1 1924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5451_6
timestamp 1730814361
transform 1 0 2808 0 -1 1920
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5375_6
timestamp 1730814361
transform 1 0 2840 0 1 1924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5451_6
timestamp 1730814361
transform 1 0 2808 0 -1 1920
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5452_6
timestamp 1730814361
transform 1 0 2992 0 -1 1920
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5455_6
timestamp 1730814361
transform 1 0 2992 0 1 1924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5452_6
timestamp 1730814361
transform 1 0 2992 0 -1 1920
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5455_6
timestamp 1730814361
transform 1 0 2992 0 1 1924
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5300_6
timestamp 1730814361
transform 1 0 3152 0 -1 1920
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5300_6
timestamp 1730814361
transform 1 0 3152 0 -1 1920
box 7 3 20 38
use welltap_svt  __well_tap__203
timestamp 1730814361
transform 1 0 3184 0 -1 1916
box 8 4 12 24
use welltap_svt  __well_tap__203
timestamp 1730814361
transform 1 0 3184 0 -1 1916
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5855_6
timestamp 1730814361
transform 1 0 128 0 1 1968
box 7 3 20 38
use welltap_svt  __well_tap__74
timestamp 1730814361
transform 1 0 104 0 -1 1956
box 8 4 12 24
use welltap_svt  __well_tap__76
timestamp 1730814361
transform 1 0 104 0 1 1972
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5855_6
timestamp 1730814361
transform 1 0 128 0 1 1968
box 7 3 20 38
use welltap_svt  __well_tap__74
timestamp 1730814361
transform 1 0 104 0 -1 1956
box 8 4 12 24
use welltap_svt  __well_tap__76
timestamp 1730814361
transform 1 0 104 0 1 1972
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5856_6
timestamp 1730814361
transform 1 0 224 0 1 1968
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5856_6
timestamp 1730814361
transform 1 0 224 0 1 1968
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5857_6
timestamp 1730814361
transform 1 0 344 0 1 1968
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5857_6
timestamp 1730814361
transform 1 0 344 0 1 1968
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5858_6
timestamp 1730814361
transform 1 0 456 0 1 1968
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5858_6
timestamp 1730814361
transform 1 0 456 0 1 1968
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5131_6
timestamp 1730814361
transform 1 0 568 0 1 1968
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5131_6
timestamp 1730814361
transform 1 0 568 0 1 1968
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5132_6
timestamp 1730814361
transform 1 0 680 0 1 1968
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5132_6
timestamp 1730814361
transform 1 0 680 0 1 1968
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5133_6
timestamp 1730814361
transform 1 0 792 0 1 1968
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5133_6
timestamp 1730814361
transform 1 0 792 0 1 1968
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5134_6
timestamp 1730814361
transform 1 0 904 0 1 1968
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5134_6
timestamp 1730814361
transform 1 0 904 0 1 1968
box 7 3 20 38
use welltap_svt  __well_tap__75
timestamp 1730814361
transform 1 0 1624 0 -1 1956
box 8 4 12 24
use welltap_svt  __well_tap__77
timestamp 1730814361
transform 1 0 1624 0 1 1972
box 8 4 12 24
use welltap_svt  __well_tap__204
timestamp 1730814361
transform 1 0 1664 0 1 1928
box 8 4 12 24
use welltap_svt  __well_tap__206
timestamp 1730814361
transform 1 0 1664 0 -1 2000
box 8 4 12 24
use welltap_svt  __well_tap__75
timestamp 1730814361
transform 1 0 1624 0 -1 1956
box 8 4 12 24
use welltap_svt  __well_tap__77
timestamp 1730814361
transform 1 0 1624 0 1 1972
box 8 4 12 24
use welltap_svt  __well_tap__204
timestamp 1730814361
transform 1 0 1664 0 1 1928
box 8 4 12 24
use welltap_svt  __well_tap__206
timestamp 1730814361
transform 1 0 1664 0 -1 2000
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5851_6
timestamp 1730814361
transform 1 0 2256 0 -1 2004
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5851_6
timestamp 1730814361
transform 1 0 2256 0 -1 2004
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5852_6
timestamp 1730814361
transform 1 0 2408 0 -1 2004
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5852_6
timestamp 1730814361
transform 1 0 2408 0 -1 2004
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5853_6
timestamp 1730814361
transform 1 0 2552 0 -1 2004
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5853_6
timestamp 1730814361
transform 1 0 2552 0 -1 2004
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5458_6
timestamp 1730814361
transform 1 0 2696 0 -1 2004
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5458_6
timestamp 1730814361
transform 1 0 2696 0 -1 2004
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5456_6
timestamp 1730814361
transform 1 0 2832 0 -1 2004
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5456_6
timestamp 1730814361
transform 1 0 2832 0 -1 2004
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5457_6
timestamp 1730814361
transform 1 0 2968 0 -1 2004
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5457_6
timestamp 1730814361
transform 1 0 2968 0 -1 2004
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5462_6
timestamp 1730814361
transform 1 0 3104 0 -1 2004
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5462_6
timestamp 1730814361
transform 1 0 3104 0 -1 2004
box 7 3 20 38
use welltap_svt  __well_tap__205
timestamp 1730814361
transform 1 0 3184 0 1 1928
box 8 4 12 24
use welltap_svt  __well_tap__207
timestamp 1730814361
transform 1 0 3184 0 -1 2000
box 8 4 12 24
use welltap_svt  __well_tap__205
timestamp 1730814361
transform 1 0 3184 0 1 1928
box 8 4 12 24
use welltap_svt  __well_tap__207
timestamp 1730814361
transform 1 0 3184 0 -1 2000
box 8 4 12 24
use welltap_svt  __well_tap__78
timestamp 1730814361
transform 1 0 104 0 -1 2044
box 8 4 12 24
use welltap_svt  __well_tap__78
timestamp 1730814361
transform 1 0 104 0 -1 2044
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5859_6
timestamp 1730814361
transform 1 0 168 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5859_6
timestamp 1730814361
transform 1 0 168 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5844_6
timestamp 1730814361
transform 1 0 360 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5844_6
timestamp 1730814361
transform 1 0 360 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5861_6
timestamp 1730814361
transform 1 0 552 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5861_6
timestamp 1730814361
transform 1 0 552 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5135_6
timestamp 1730814361
transform 1 0 752 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5135_6
timestamp 1730814361
transform 1 0 752 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5136_6
timestamp 1730814361
transform 1 0 960 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5136_6
timestamp 1730814361
transform 1 0 960 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5137_6
timestamp 1730814361
transform 1 0 1176 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5137_6
timestamp 1730814361
transform 1 0 1176 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5224_6
timestamp 1730814361
transform 1 0 1392 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5224_6
timestamp 1730814361
transform 1 0 1392 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5225_6
timestamp 1730814361
transform 1 0 1592 0 -1 2048
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5225_6
timestamp 1730814361
transform 1 0 1592 0 -1 2048
box 7 3 20 38
use welltap_svt  __well_tap__79
timestamp 1730814361
transform 1 0 1624 0 -1 2044
box 8 4 12 24
use welltap_svt  __well_tap__208
timestamp 1730814361
transform 1 0 1664 0 1 2016
box 8 4 12 24
use welltap_svt  __well_tap__79
timestamp 1730814361
transform 1 0 1624 0 -1 2044
box 8 4 12 24
use welltap_svt  __well_tap__208
timestamp 1730814361
transform 1 0 1664 0 1 2016
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5226_6
timestamp 1730814361
transform 1 0 1688 0 1 2012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5227_6
timestamp 1730814361
transform 1 0 1688 0 -1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5226_6
timestamp 1730814361
transform 1 0 1688 0 1 2012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5227_6
timestamp 1730814361
transform 1 0 1688 0 -1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5228_6
timestamp 1730814361
transform 1 0 1816 0 -1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5228_6
timestamp 1730814361
transform 1 0 1816 0 -1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5229_6
timestamp 1730814361
transform 1 0 1960 0 -1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5229_6
timestamp 1730814361
transform 1 0 1960 0 -1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5459_6
timestamp 1730814361
transform 1 0 2032 0 1 2012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5459_6
timestamp 1730814361
transform 1 0 2032 0 1 2012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5854_6
timestamp 1730814361
transform 1 0 2104 0 -1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5854_6
timestamp 1730814361
transform 1 0 2104 0 -1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5301_6
timestamp 1730814361
transform 1 0 2248 0 -1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5301_6
timestamp 1730814361
transform 1 0 2248 0 -1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5302_6
timestamp 1730814361
transform 1 0 2400 0 -1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5460_6
timestamp 1730814361
transform 1 0 2400 0 1 2012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5302_6
timestamp 1730814361
transform 1 0 2400 0 -1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5460_6
timestamp 1730814361
transform 1 0 2400 0 1 2012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5461_6
timestamp 1730814361
transform 1 0 2760 0 1 2012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5461_6
timestamp 1730814361
transform 1 0 2760 0 1 2012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5328_6
timestamp 1730814361
transform 1 0 3128 0 1 2012
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5328_6
timestamp 1730814361
transform 1 0 3128 0 1 2012
box 7 3 20 38
use welltap_svt  __well_tap__209
timestamp 1730814361
transform 1 0 3184 0 1 2016
box 8 4 12 24
use welltap_svt  __well_tap__209
timestamp 1730814361
transform 1 0 3184 0 1 2016
box 8 4 12 24
use welltap_svt  __well_tap__80
timestamp 1730814361
transform 1 0 104 0 1 2060
box 8 4 12 24
use welltap_svt  __well_tap__80
timestamp 1730814361
transform 1 0 104 0 1 2060
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5862_6
timestamp 1730814361
transform 1 0 240 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5862_6
timestamp 1730814361
transform 1 0 240 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5863_6
timestamp 1730814361
transform 1 0 368 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5866_6
timestamp 1730814361
transform 1 0 344 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5863_6
timestamp 1730814361
transform 1 0 368 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5866_6
timestamp 1730814361
transform 1 0 344 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5864_6
timestamp 1730814361
transform 1 0 496 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5867_6
timestamp 1730814361
transform 1 0 472 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5864_6
timestamp 1730814361
transform 1 0 496 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5867_6
timestamp 1730814361
transform 1 0 472 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5865_6
timestamp 1730814361
transform 1 0 616 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5868_6
timestamp 1730814361
transform 1 0 592 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5865_6
timestamp 1730814361
transform 1 0 616 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5868_6
timestamp 1730814361
transform 1 0 592 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5138_6
timestamp 1730814361
transform 1 0 736 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5869_6
timestamp 1730814361
transform 1 0 712 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5138_6
timestamp 1730814361
transform 1 0 736 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5869_6
timestamp 1730814361
transform 1 0 712 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5139_6
timestamp 1730814361
transform 1 0 848 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5142_6
timestamp 1730814361
transform 1 0 832 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5139_6
timestamp 1730814361
transform 1 0 848 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5142_6
timestamp 1730814361
transform 1 0 832 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5140_6
timestamp 1730814361
transform 1 0 960 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5143_6
timestamp 1730814361
transform 1 0 944 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5140_6
timestamp 1730814361
transform 1 0 960 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5143_6
timestamp 1730814361
transform 1 0 944 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5144_6
timestamp 1730814361
transform 1 0 1056 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5144_6
timestamp 1730814361
transform 1 0 1056 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5188_6
timestamp 1730814361
transform 1 0 1080 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5188_6
timestamp 1730814361
transform 1 0 1080 0 1 2056
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5145_6
timestamp 1730814361
transform 1 0 1176 0 -1 2148
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5145_6
timestamp 1730814361
transform 1 0 1176 0 -1 2148
box 7 3 20 38
use welltap_svt  __well_tap__81
timestamp 1730814361
transform 1 0 1624 0 1 2060
box 8 4 12 24
use welltap_svt  __well_tap__210
timestamp 1730814361
transform 1 0 1664 0 -1 2088
box 8 4 12 24
use welltap_svt  __well_tap__212
timestamp 1730814361
transform 1 0 1664 0 1 2096
box 8 4 12 24
use welltap_svt  __well_tap__81
timestamp 1730814361
transform 1 0 1624 0 1 2060
box 8 4 12 24
use welltap_svt  __well_tap__210
timestamp 1730814361
transform 1 0 1664 0 -1 2088
box 8 4 12 24
use welltap_svt  __well_tap__212
timestamp 1730814361
transform 1 0 1664 0 1 2096
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5230_6
timestamp 1730814361
transform 1 0 1752 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5230_6
timestamp 1730814361
transform 1 0 1752 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5231_6
timestamp 1730814361
transform 1 0 1904 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5231_6
timestamp 1730814361
transform 1 0 1904 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5232_6
timestamp 1730814361
transform 1 0 2064 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5232_6
timestamp 1730814361
transform 1 0 2064 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5303_6
timestamp 1730814361
transform 1 0 2248 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5303_6
timestamp 1730814361
transform 1 0 2248 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5304_6
timestamp 1730814361
transform 1 0 2456 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5304_6
timestamp 1730814361
transform 1 0 2456 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5305_6
timestamp 1730814361
transform 1 0 2680 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5305_6
timestamp 1730814361
transform 1 0 2680 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5306_6
timestamp 1730814361
transform 1 0 2920 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5306_6
timestamp 1730814361
transform 1 0 2920 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_50_6
timestamp 1730814361
transform 1 0 3152 0 1 2092
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_50_6
timestamp 1730814361
transform 1 0 3152 0 1 2092
box 7 3 20 38
use welltap_svt  __well_tap__211
timestamp 1730814361
transform 1 0 3184 0 -1 2088
box 8 4 12 24
use welltap_svt  __well_tap__213
timestamp 1730814361
transform 1 0 3184 0 1 2096
box 8 4 12 24
use welltap_svt  __well_tap__211
timestamp 1730814361
transform 1 0 3184 0 -1 2088
box 8 4 12 24
use welltap_svt  __well_tap__213
timestamp 1730814361
transform 1 0 3184 0 1 2096
box 8 4 12 24
use welltap_svt  __well_tap__82
timestamp 1730814361
transform 1 0 104 0 -1 2144
box 8 4 12 24
use welltap_svt  __well_tap__84
timestamp 1730814361
transform 1 0 104 0 1 2164
box 8 4 12 24
use welltap_svt  __well_tap__82
timestamp 1730814361
transform 1 0 104 0 -1 2144
box 8 4 12 24
use welltap_svt  __well_tap__84
timestamp 1730814361
transform 1 0 104 0 1 2164
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5870_6
timestamp 1730814361
transform 1 0 448 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5870_6
timestamp 1730814361
transform 1 0 448 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5871_6
timestamp 1730814361
transform 1 0 576 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5871_6
timestamp 1730814361
transform 1 0 576 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5872_6
timestamp 1730814361
transform 1 0 696 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5872_6
timestamp 1730814361
transform 1 0 696 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5873_6
timestamp 1730814361
transform 1 0 816 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5873_6
timestamp 1730814361
transform 1 0 816 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5146_6
timestamp 1730814361
transform 1 0 936 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5146_6
timestamp 1730814361
transform 1 0 936 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5147_6
timestamp 1730814361
transform 1 0 1048 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5147_6
timestamp 1730814361
transform 1 0 1048 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5148_6
timestamp 1730814361
transform 1 0 1160 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5148_6
timestamp 1730814361
transform 1 0 1160 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5149_6
timestamp 1730814361
transform 1 0 1280 0 1 2160
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5149_6
timestamp 1730814361
transform 1 0 1280 0 1 2160
box 7 3 20 38
use welltap_svt  __well_tap__83
timestamp 1730814361
transform 1 0 1624 0 -1 2144
box 8 4 12 24
use welltap_svt  __well_tap__85
timestamp 1730814361
transform 1 0 1624 0 1 2164
box 8 4 12 24
use welltap_svt  __well_tap__214
timestamp 1730814361
transform 1 0 1664 0 -1 2172
box 8 4 12 24
use welltap_svt  __well_tap__83
timestamp 1730814361
transform 1 0 1624 0 -1 2144
box 8 4 12 24
use welltap_svt  __well_tap__85
timestamp 1730814361
transform 1 0 1624 0 1 2164
box 8 4 12 24
use welltap_svt  __well_tap__214
timestamp 1730814361
transform 1 0 1664 0 -1 2172
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5233_6
timestamp 1730814361
transform 1 0 1840 0 -1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5233_6
timestamp 1730814361
transform 1 0 1840 0 -1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5236_6
timestamp 1730814361
transform 1 0 1920 0 1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5236_6
timestamp 1730814361
transform 1 0 1920 0 1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5234_6
timestamp 1730814361
transform 1 0 1992 0 -1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5234_6
timestamp 1730814361
transform 1 0 1992 0 -1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5237_6
timestamp 1730814361
transform 1 0 2096 0 1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5237_6
timestamp 1730814361
transform 1 0 2096 0 1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5219_6
timestamp 1730814361
transform 1 0 2144 0 -1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5219_6
timestamp 1730814361
transform 1 0 2144 0 -1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5238_6
timestamp 1730814361
transform 1 0 2288 0 1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5307_6
timestamp 1730814361
transform 1 0 2288 0 -1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5238_6
timestamp 1730814361
transform 1 0 2288 0 1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5307_6
timestamp 1730814361
transform 1 0 2288 0 -1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5308_6
timestamp 1730814361
transform 1 0 2440 0 -1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5308_6
timestamp 1730814361
transform 1 0 2440 0 -1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5310_6
timestamp 1730814361
transform 1 0 2496 0 1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5310_6
timestamp 1730814361
transform 1 0 2496 0 1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5309_6
timestamp 1730814361
transform 1 0 2592 0 -1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5309_6
timestamp 1730814361
transform 1 0 2592 0 -1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5311_6
timestamp 1730814361
transform 1 0 2712 0 1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5311_6
timestamp 1730814361
transform 1 0 2712 0 1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5312_6
timestamp 1730814361
transform 1 0 2944 0 1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5312_6
timestamp 1730814361
transform 1 0 2944 0 1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5330_6
timestamp 1730814361
transform 1 0 3152 0 1 2176
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5330_6
timestamp 1730814361
transform 1 0 3152 0 1 2176
box 7 3 20 38
use welltap_svt  __well_tap__215
timestamp 1730814361
transform 1 0 3184 0 -1 2172
box 8 4 12 24
use welltap_svt  __well_tap__215
timestamp 1730814361
transform 1 0 3184 0 -1 2172
box 8 4 12 24
use welltap_svt  __well_tap__86
timestamp 1730814361
transform 1 0 104 0 -1 2244
box 8 4 12 24
use welltap_svt  __well_tap__86
timestamp 1730814361
transform 1 0 104 0 -1 2244
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5874_6
timestamp 1730814361
transform 1 0 544 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5874_6
timestamp 1730814361
transform 1 0 544 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5829_6
timestamp 1730814361
transform 1 0 672 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5829_6
timestamp 1730814361
transform 1 0 672 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5814_6
timestamp 1730814361
transform 1 0 800 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5814_6
timestamp 1730814361
transform 1 0 800 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5815_6
timestamp 1730814361
transform 1 0 920 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5815_6
timestamp 1730814361
transform 1 0 920 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5150_6
timestamp 1730814361
transform 1 0 1040 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5150_6
timestamp 1730814361
transform 1 0 1040 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5151_6
timestamp 1730814361
transform 1 0 1152 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5151_6
timestamp 1730814361
transform 1 0 1152 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5152_6
timestamp 1730814361
transform 1 0 1264 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5152_6
timestamp 1730814361
transform 1 0 1264 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5153_6
timestamp 1730814361
transform 1 0 1384 0 -1 2248
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5153_6
timestamp 1730814361
transform 1 0 1384 0 -1 2248
box 7 3 20 38
use welltap_svt  __well_tap__87
timestamp 1730814361
transform 1 0 1624 0 -1 2244
box 8 4 12 24
use welltap_svt  __well_tap__216
timestamp 1730814361
transform 1 0 1664 0 1 2180
box 8 4 12 24
use welltap_svt  __well_tap__218
timestamp 1730814361
transform 1 0 1664 0 -1 2256
box 8 4 12 24
use welltap_svt  __well_tap__87
timestamp 1730814361
transform 1 0 1624 0 -1 2244
box 8 4 12 24
use welltap_svt  __well_tap__216
timestamp 1730814361
transform 1 0 1664 0 1 2180
box 8 4 12 24
use welltap_svt  __well_tap__218
timestamp 1730814361
transform 1 0 1664 0 -1 2256
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5239_6
timestamp 1730814361
transform 1 0 2008 0 -1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5239_6
timestamp 1730814361
transform 1 0 2008 0 -1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5240_6
timestamp 1730814361
transform 1 0 2160 0 -1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5240_6
timestamp 1730814361
transform 1 0 2160 0 -1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5241_6
timestamp 1730814361
transform 1 0 2312 0 -1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5241_6
timestamp 1730814361
transform 1 0 2312 0 -1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5266_6
timestamp 1730814361
transform 1 0 2456 0 -1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5266_6
timestamp 1730814361
transform 1 0 2456 0 -1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5251_6
timestamp 1730814361
transform 1 0 2600 0 -1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5251_6
timestamp 1730814361
transform 1 0 2600 0 -1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5252_6
timestamp 1730814361
transform 1 0 2752 0 -1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5252_6
timestamp 1730814361
transform 1 0 2752 0 -1 2260
box 7 3 20 38
use welltap_svt  __well_tap__217
timestamp 1730814361
transform 1 0 3184 0 1 2180
box 8 4 12 24
use welltap_svt  __well_tap__219
timestamp 1730814361
transform 1 0 3184 0 -1 2256
box 8 4 12 24
use welltap_svt  __well_tap__217
timestamp 1730814361
transform 1 0 3184 0 1 2180
box 8 4 12 24
use welltap_svt  __well_tap__219
timestamp 1730814361
transform 1 0 3184 0 -1 2256
box 8 4 12 24
use welltap_svt  __well_tap__88
timestamp 1730814361
transform 1 0 104 0 1 2264
box 8 4 12 24
use welltap_svt  __well_tap__88
timestamp 1730814361
transform 1 0 104 0 1 2264
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5816_6
timestamp 1730814361
transform 1 0 648 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5816_6
timestamp 1730814361
transform 1 0 648 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5817_6
timestamp 1730814361
transform 1 0 776 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5817_6
timestamp 1730814361
transform 1 0 776 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5818_6
timestamp 1730814361
transform 1 0 896 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5818_6
timestamp 1730814361
transform 1 0 896 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5819_6
timestamp 1730814361
transform 1 0 1016 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5819_6
timestamp 1730814361
transform 1 0 1016 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5154_6
timestamp 1730814361
transform 1 0 1136 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5154_6
timestamp 1730814361
transform 1 0 1136 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5155_6
timestamp 1730814361
transform 1 0 1248 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5155_6
timestamp 1730814361
transform 1 0 1248 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5235_6
timestamp 1730814361
transform 1 0 1360 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5235_6
timestamp 1730814361
transform 1 0 1360 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5220_6
timestamp 1730814361
transform 1 0 1480 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5220_6
timestamp 1730814361
transform 1 0 1480 0 1 2260
box 7 3 20 38
use welltap_svt  __well_tap__89
timestamp 1730814361
transform 1 0 1624 0 1 2264
box 8 4 12 24
use welltap_svt  __well_tap__220
timestamp 1730814361
transform 1 0 1664 0 1 2264
box 8 4 12 24
use welltap_svt  __well_tap__89
timestamp 1730814361
transform 1 0 1624 0 1 2264
box 8 4 12 24
use welltap_svt  __well_tap__220
timestamp 1730814361
transform 1 0 1664 0 1 2264
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5242_6
timestamp 1730814361
transform 1 0 2088 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5242_6
timestamp 1730814361
transform 1 0 2088 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5243_6
timestamp 1730814361
transform 1 0 2256 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5243_6
timestamp 1730814361
transform 1 0 2256 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5244_6
timestamp 1730814361
transform 1 0 2424 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5244_6
timestamp 1730814361
transform 1 0 2424 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5253_6
timestamp 1730814361
transform 1 0 2600 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5253_6
timestamp 1730814361
transform 1 0 2600 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5254_6
timestamp 1730814361
transform 1 0 2784 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5254_6
timestamp 1730814361
transform 1 0 2784 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5255_6
timestamp 1730814361
transform 1 0 2976 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5255_6
timestamp 1730814361
transform 1 0 2976 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5331_6
timestamp 1730814361
transform 1 0 3152 0 1 2260
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5331_6
timestamp 1730814361
transform 1 0 3152 0 1 2260
box 7 3 20 38
use welltap_svt  __well_tap__221
timestamp 1730814361
transform 1 0 3184 0 1 2264
box 8 4 12 24
use welltap_svt  __well_tap__221
timestamp 1730814361
transform 1 0 3184 0 1 2264
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5823_6
timestamp 1730814361
transform 1 0 128 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5824_6
timestamp 1730814361
transform 1 0 128 0 1 2360
box 7 3 20 38
use welltap_svt  __well_tap__90
timestamp 1730814361
transform 1 0 104 0 -1 2348
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5823_6
timestamp 1730814361
transform 1 0 128 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5824_6
timestamp 1730814361
transform 1 0 128 0 1 2360
box 7 3 20 38
use welltap_svt  __well_tap__90
timestamp 1730814361
transform 1 0 104 0 -1 2348
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5825_6
timestamp 1730814361
transform 1 0 232 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5825_6
timestamp 1730814361
transform 1 0 232 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5820_6
timestamp 1730814361
transform 1 0 336 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5826_6
timestamp 1730814361
transform 1 0 352 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5820_6
timestamp 1730814361
transform 1 0 336 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5826_6
timestamp 1730814361
transform 1 0 352 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5827_6
timestamp 1730814361
transform 1 0 472 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5827_6
timestamp 1730814361
transform 1 0 472 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5821_6
timestamp 1730814361
transform 1 0 560 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5821_6
timestamp 1730814361
transform 1 0 560 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5193_6
timestamp 1730814361
transform 1 0 584 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5193_6
timestamp 1730814361
transform 1 0 584 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5194_6
timestamp 1730814361
transform 1 0 696 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5194_6
timestamp 1730814361
transform 1 0 696 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5195_6
timestamp 1730814361
transform 1 0 808 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5822_6
timestamp 1730814361
transform 1 0 768 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5195_6
timestamp 1730814361
transform 1 0 808 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5822_6
timestamp 1730814361
transform 1 0 768 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5196_6
timestamp 1730814361
transform 1 0 928 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5196_6
timestamp 1730814361
transform 1 0 928 0 1 2360
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5192_6
timestamp 1730814361
transform 1 0 968 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5192_6
timestamp 1730814361
transform 1 0 968 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5221_6
timestamp 1730814361
transform 1 0 1168 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5221_6
timestamp 1730814361
transform 1 0 1168 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5222_6
timestamp 1730814361
transform 1 0 1360 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5222_6
timestamp 1730814361
transform 1 0 1360 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5223_6
timestamp 1730814361
transform 1 0 1560 0 -1 2352
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5223_6
timestamp 1730814361
transform 1 0 1560 0 -1 2352
box 7 3 20 38
use welltap_svt  __well_tap__91
timestamp 1730814361
transform 1 0 1624 0 -1 2348
box 8 4 12 24
use welltap_svt  __well_tap__222
timestamp 1730814361
transform 1 0 1664 0 -1 2340
box 8 4 12 24
use welltap_svt  __well_tap__224
timestamp 1730814361
transform 1 0 1664 0 1 2348
box 8 4 12 24
use welltap_svt  __well_tap__91
timestamp 1730814361
transform 1 0 1624 0 -1 2348
box 8 4 12 24
use welltap_svt  __well_tap__222
timestamp 1730814361
transform 1 0 1664 0 -1 2340
box 8 4 12 24
use welltap_svt  __well_tap__224
timestamp 1730814361
transform 1 0 1664 0 1 2348
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5245_6
timestamp 1730814361
transform 1 0 2176 0 -1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5248_6
timestamp 1730814361
transform 1 0 2136 0 1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5245_6
timestamp 1730814361
transform 1 0 2176 0 -1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5248_6
timestamp 1730814361
transform 1 0 2136 0 1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5249_6
timestamp 1730814361
transform 1 0 2304 0 1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5249_6
timestamp 1730814361
transform 1 0 2304 0 1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5246_6
timestamp 1730814361
transform 1 0 2328 0 -1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5246_6
timestamp 1730814361
transform 1 0 2328 0 -1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5204_6
timestamp 1730814361
transform 1 0 2472 0 1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5247_6
timestamp 1730814361
transform 1 0 2472 0 -1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5204_6
timestamp 1730814361
transform 1 0 2472 0 1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5247_6
timestamp 1730814361
transform 1 0 2472 0 -1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5256_6
timestamp 1730814361
transform 1 0 2616 0 -1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5259_6
timestamp 1730814361
transform 1 0 2648 0 1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5256_6
timestamp 1730814361
transform 1 0 2616 0 -1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5259_6
timestamp 1730814361
transform 1 0 2648 0 1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5257_6
timestamp 1730814361
transform 1 0 2760 0 -1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5257_6
timestamp 1730814361
transform 1 0 2760 0 -1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5260_6
timestamp 1730814361
transform 1 0 2824 0 1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5260_6
timestamp 1730814361
transform 1 0 2824 0 1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5258_6
timestamp 1730814361
transform 1 0 2912 0 -1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5258_6
timestamp 1730814361
transform 1 0 2912 0 -1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5261_6
timestamp 1730814361
transform 1 0 3000 0 1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5261_6
timestamp 1730814361
transform 1 0 3000 0 1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5332_6
timestamp 1730814361
transform 1 0 3152 0 1 2344
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5332_6
timestamp 1730814361
transform 1 0 3152 0 1 2344
box 7 3 20 38
use welltap_svt  __well_tap__223
timestamp 1730814361
transform 1 0 3184 0 -1 2340
box 8 4 12 24
use welltap_svt  __well_tap__225
timestamp 1730814361
transform 1 0 3184 0 1 2348
box 8 4 12 24
use welltap_svt  __well_tap__223
timestamp 1730814361
transform 1 0 3184 0 -1 2340
box 8 4 12 24
use welltap_svt  __well_tap__225
timestamp 1730814361
transform 1 0 3184 0 1 2348
box 8 4 12 24
use welltap_svt  __well_tap__92
timestamp 1730814361
transform 1 0 104 0 1 2364
box 8 4 12 24
use welltap_svt  __well_tap__92
timestamp 1730814361
transform 1 0 104 0 1 2364
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5828_6
timestamp 1730814361
transform 1 0 192 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5828_6
timestamp 1730814361
transform 1 0 192 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5500_6
timestamp 1730814361
transform 1 0 320 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5500_6
timestamp 1730814361
transform 1 0 320 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5830_6
timestamp 1730814361
transform 1 0 448 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5830_6
timestamp 1730814361
transform 1 0 448 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5831_6
timestamp 1730814361
transform 1 0 592 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5831_6
timestamp 1730814361
transform 1 0 592 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5197_6
timestamp 1730814361
transform 1 0 760 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5197_6
timestamp 1730814361
transform 1 0 760 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5198_6
timestamp 1730814361
transform 1 0 944 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5198_6
timestamp 1730814361
transform 1 0 944 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5199_6
timestamp 1730814361
transform 1 0 1152 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5199_6
timestamp 1730814361
transform 1 0 1152 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5200_6
timestamp 1730814361
transform 1 0 1368 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5200_6
timestamp 1730814361
transform 1 0 1368 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_51_6
timestamp 1730814361
transform 1 0 1584 0 -1 2456
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_51_6
timestamp 1730814361
transform 1 0 1584 0 -1 2456
box 7 3 20 38
use welltap_svt  __well_tap__93
timestamp 1730814361
transform 1 0 1624 0 1 2364
box 8 4 12 24
use welltap_svt  __well_tap__226
timestamp 1730814361
transform 1 0 1664 0 -1 2428
box 8 4 12 24
use welltap_svt  __well_tap__93
timestamp 1730814361
transform 1 0 1624 0 1 2364
box 8 4 12 24
use welltap_svt  __well_tap__226
timestamp 1730814361
transform 1 0 1664 0 -1 2428
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5189_6
timestamp 1730814361
transform 1 0 2224 0 -1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5189_6
timestamp 1730814361
transform 1 0 2224 0 -1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5190_6
timestamp 1730814361
transform 1 0 2384 0 -1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5190_6
timestamp 1730814361
transform 1 0 2384 0 -1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5191_6
timestamp 1730814361
transform 1 0 2536 0 -1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5191_6
timestamp 1730814361
transform 1 0 2536 0 -1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5262_6
timestamp 1730814361
transform 1 0 2680 0 -1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5262_6
timestamp 1730814361
transform 1 0 2680 0 -1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5263_6
timestamp 1730814361
transform 1 0 2816 0 -1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5263_6
timestamp 1730814361
transform 1 0 2816 0 -1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5264_6
timestamp 1730814361
transform 1 0 2960 0 -1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5264_6
timestamp 1730814361
transform 1 0 2960 0 -1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5333_6
timestamp 1730814361
transform 1 0 3104 0 -1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5333_6
timestamp 1730814361
transform 1 0 3104 0 -1 2432
box 7 3 20 38
use welltap_svt  __well_tap__227
timestamp 1730814361
transform 1 0 3184 0 -1 2428
box 8 4 12 24
use welltap_svt  __well_tap__227
timestamp 1730814361
transform 1 0 3184 0 -1 2428
box 8 4 12 24
use welltap_svt  __well_tap__94
timestamp 1730814361
transform 1 0 104 0 -1 2452
box 8 4 12 24
use welltap_svt  __well_tap__96
timestamp 1730814361
transform 1 0 104 0 1 2464
box 8 4 12 24
use welltap_svt  __well_tap__94
timestamp 1730814361
transform 1 0 104 0 -1 2452
box 8 4 12 24
use welltap_svt  __well_tap__96
timestamp 1730814361
transform 1 0 104 0 1 2464
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5832_6
timestamp 1730814361
transform 1 0 296 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5832_6
timestamp 1730814361
transform 1 0 296 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5833_6
timestamp 1730814361
transform 1 0 424 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5833_6
timestamp 1730814361
transform 1 0 424 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5834_6
timestamp 1730814361
transform 1 0 552 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5834_6
timestamp 1730814361
transform 1 0 552 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5835_6
timestamp 1730814361
transform 1 0 696 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5835_6
timestamp 1730814361
transform 1 0 696 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5201_6
timestamp 1730814361
transform 1 0 856 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5201_6
timestamp 1730814361
transform 1 0 856 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5202_6
timestamp 1730814361
transform 1 0 1032 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5202_6
timestamp 1730814361
transform 1 0 1032 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5203_6
timestamp 1730814361
transform 1 0 1216 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5203_6
timestamp 1730814361
transform 1 0 1216 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5125_6
timestamp 1730814361
transform 1 0 1416 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5125_6
timestamp 1730814361
transform 1 0 1416 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_52_6
timestamp 1730814361
transform 1 0 1592 0 1 2460
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_52_6
timestamp 1730814361
transform 1 0 1592 0 1 2460
box 7 3 20 38
use welltap_svt  __well_tap__95
timestamp 1730814361
transform 1 0 1624 0 -1 2452
box 8 4 12 24
use welltap_svt  __well_tap__97
timestamp 1730814361
transform 1 0 1624 0 1 2464
box 8 4 12 24
use welltap_svt  __well_tap__228
timestamp 1730814361
transform 1 0 1664 0 1 2436
box 8 4 12 24
use welltap_svt  __well_tap__95
timestamp 1730814361
transform 1 0 1624 0 -1 2452
box 8 4 12 24
use welltap_svt  __well_tap__97
timestamp 1730814361
transform 1 0 1624 0 1 2464
box 8 4 12 24
use welltap_svt  __well_tap__228
timestamp 1730814361
transform 1 0 1664 0 1 2436
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_53_6
timestamp 1730814361
transform 1 0 1688 0 -1 2520
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_53_6
timestamp 1730814361
transform 1 0 1688 0 -1 2520
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_54_6
timestamp 1730814361
transform 1 0 1856 0 -1 2520
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_54_6
timestamp 1730814361
transform 1 0 1856 0 -1 2520
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_55_6
timestamp 1730814361
transform 1 0 2072 0 -1 2520
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_55_6
timestamp 1730814361
transform 1 0 2072 0 -1 2520
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5267_6
timestamp 1730814361
transform 1 0 2312 0 1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5269_6
timestamp 1730814361
transform 1 0 2312 0 -1 2520
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5267_6
timestamp 1730814361
transform 1 0 2312 0 1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5269_6
timestamp 1730814361
transform 1 0 2312 0 -1 2520
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5268_6
timestamp 1730814361
transform 1 0 2560 0 1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5270_6
timestamp 1730814361
transform 1 0 2576 0 -1 2520
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5268_6
timestamp 1730814361
transform 1 0 2560 0 1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5270_6
timestamp 1730814361
transform 1 0 2576 0 -1 2520
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5265_6
timestamp 1730814361
transform 1 0 2816 0 1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5271_6
timestamp 1730814361
transform 1 0 2848 0 -1 2520
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5265_6
timestamp 1730814361
transform 1 0 2816 0 1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5271_6
timestamp 1730814361
transform 1 0 2848 0 -1 2520
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5313_6
timestamp 1730814361
transform 1 0 3072 0 1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5313_6
timestamp 1730814361
transform 1 0 3072 0 1 2432
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5334_6
timestamp 1730814361
transform 1 0 3128 0 -1 2520
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5334_6
timestamp 1730814361
transform 1 0 3128 0 -1 2520
box 7 3 20 38
use welltap_svt  __well_tap__229
timestamp 1730814361
transform 1 0 3184 0 1 2436
box 8 4 12 24
use welltap_svt  __well_tap__229
timestamp 1730814361
transform 1 0 3184 0 1 2436
box 8 4 12 24
use welltap_svt  __well_tap__98
timestamp 1730814361
transform 1 0 104 0 -1 2548
box 8 4 12 24
use welltap_svt  __well_tap__98
timestamp 1730814361
transform 1 0 104 0 -1 2548
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5836_6
timestamp 1730814361
transform 1 0 392 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5836_6
timestamp 1730814361
transform 1 0 392 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5837_6
timestamp 1730814361
transform 1 0 520 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5837_6
timestamp 1730814361
transform 1 0 520 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5838_6
timestamp 1730814361
transform 1 0 648 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5838_6
timestamp 1730814361
transform 1 0 648 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5839_6
timestamp 1730814361
transform 1 0 768 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5839_6
timestamp 1730814361
transform 1 0 768 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5205_6
timestamp 1730814361
transform 1 0 888 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5205_6
timestamp 1730814361
transform 1 0 888 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5206_6
timestamp 1730814361
transform 1 0 1000 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5206_6
timestamp 1730814361
transform 1 0 1000 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5207_6
timestamp 1730814361
transform 1 0 1112 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5207_6
timestamp 1730814361
transform 1 0 1112 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5208_6
timestamp 1730814361
transform 1 0 1232 0 -1 2552
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5208_6
timestamp 1730814361
transform 1 0 1232 0 -1 2552
box 7 3 20 38
use welltap_svt  __well_tap__99
timestamp 1730814361
transform 1 0 1624 0 -1 2548
box 8 4 12 24
use welltap_svt  __well_tap__230
timestamp 1730814361
transform 1 0 1664 0 -1 2516
box 8 4 12 24
use welltap_svt  __well_tap__232
timestamp 1730814361
transform 1 0 1664 0 1 2528
box 8 4 12 24
use welltap_svt  __well_tap__99
timestamp 1730814361
transform 1 0 1624 0 -1 2548
box 8 4 12 24
use welltap_svt  __well_tap__230
timestamp 1730814361
transform 1 0 1664 0 -1 2516
box 8 4 12 24
use welltap_svt  __well_tap__232
timestamp 1730814361
transform 1 0 1664 0 1 2528
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_56_6
timestamp 1730814361
transform 1 0 1728 0 1 2524
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_56_6
timestamp 1730814361
transform 1 0 1728 0 1 2524
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_57_6
timestamp 1730814361
transform 1 0 1888 0 1 2524
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_57_6
timestamp 1730814361
transform 1 0 1888 0 1 2524
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_58_6
timestamp 1730814361
transform 1 0 2048 0 1 2524
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_58_6
timestamp 1730814361
transform 1 0 2048 0 1 2524
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5272_6
timestamp 1730814361
transform 1 0 2208 0 1 2524
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5272_6
timestamp 1730814361
transform 1 0 2208 0 1 2524
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5273_6
timestamp 1730814361
transform 1 0 2368 0 1 2524
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5273_6
timestamp 1730814361
transform 1 0 2368 0 1 2524
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5274_6
timestamp 1730814361
transform 1 0 2528 0 1 2524
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5274_6
timestamp 1730814361
transform 1 0 2528 0 1 2524
box 7 3 20 38
use welltap_svt  __well_tap__231
timestamp 1730814361
transform 1 0 3184 0 -1 2516
box 8 4 12 24
use welltap_svt  __well_tap__233
timestamp 1730814361
transform 1 0 3184 0 1 2528
box 8 4 12 24
use welltap_svt  __well_tap__231
timestamp 1730814361
transform 1 0 3184 0 -1 2516
box 8 4 12 24
use welltap_svt  __well_tap__233
timestamp 1730814361
transform 1 0 3184 0 1 2528
box 8 4 12 24
use welltap_svt  __well_tap__100
timestamp 1730814361
transform 1 0 104 0 1 2568
box 8 4 12 24
use welltap_svt  __well_tap__100
timestamp 1730814361
transform 1 0 104 0 1 2568
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5840_6
timestamp 1730814361
transform 1 0 496 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5840_6
timestamp 1730814361
transform 1 0 496 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5841_6
timestamp 1730814361
transform 1 0 624 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5841_6
timestamp 1730814361
transform 1 0 624 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5842_6
timestamp 1730814361
transform 1 0 744 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5842_6
timestamp 1730814361
transform 1 0 744 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5843_6
timestamp 1730814361
transform 1 0 864 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5843_6
timestamp 1730814361
transform 1 0 864 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5209_6
timestamp 1730814361
transform 1 0 984 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5209_6
timestamp 1730814361
transform 1 0 984 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5210_6
timestamp 1730814361
transform 1 0 1096 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5210_6
timestamp 1730814361
transform 1 0 1096 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5211_6
timestamp 1730814361
transform 1 0 1208 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5211_6
timestamp 1730814361
transform 1 0 1208 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5212_6
timestamp 1730814361
transform 1 0 1328 0 1 2564
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5212_6
timestamp 1730814361
transform 1 0 1328 0 1 2564
box 7 3 20 38
use welltap_svt  __well_tap__101
timestamp 1730814361
transform 1 0 1624 0 1 2568
box 8 4 12 24
use welltap_svt  __well_tap__234
timestamp 1730814361
transform 1 0 1664 0 -1 2604
box 8 4 12 24
use welltap_svt  __well_tap__101
timestamp 1730814361
transform 1 0 1624 0 1 2568
box 8 4 12 24
use welltap_svt  __well_tap__234
timestamp 1730814361
transform 1 0 1664 0 -1 2604
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_59_6
timestamp 1730814361
transform 1 0 1816 0 -1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_59_6
timestamp 1730814361
transform 1 0 1816 0 -1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_512_6
timestamp 1730814361
transform 1 0 1904 0 1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_512_6
timestamp 1730814361
transform 1 0 1904 0 1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_510_6
timestamp 1730814361
transform 1 0 2008 0 -1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_510_6
timestamp 1730814361
transform 1 0 2008 0 -1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_513_6
timestamp 1730814361
transform 1 0 2096 0 1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_513_6
timestamp 1730814361
transform 1 0 2096 0 1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_511_6
timestamp 1730814361
transform 1 0 2208 0 -1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_511_6
timestamp 1730814361
transform 1 0 2208 0 -1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_514_6
timestamp 1730814361
transform 1 0 2288 0 1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_514_6
timestamp 1730814361
transform 1 0 2288 0 1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5275_6
timestamp 1730814361
transform 1 0 2432 0 -1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5278_6
timestamp 1730814361
transform 1 0 2480 0 1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5275_6
timestamp 1730814361
transform 1 0 2432 0 -1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5278_6
timestamp 1730814361
transform 1 0 2480 0 1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5276_6
timestamp 1730814361
transform 1 0 2664 0 -1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5276_6
timestamp 1730814361
transform 1 0 2664 0 -1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5279_6
timestamp 1730814361
transform 1 0 2680 0 1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5279_6
timestamp 1730814361
transform 1 0 2680 0 1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5277_6
timestamp 1730814361
transform 1 0 2912 0 -1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5277_6
timestamp 1730814361
transform 1 0 2912 0 -1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5335_6
timestamp 1730814361
transform 1 0 3152 0 -1 2608
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5335_6
timestamp 1730814361
transform 1 0 3152 0 -1 2608
box 7 3 20 38
use welltap_svt  __well_tap__235
timestamp 1730814361
transform 1 0 3184 0 -1 2604
box 8 4 12 24
use welltap_svt  __well_tap__235
timestamp 1730814361
transform 1 0 3184 0 -1 2604
box 8 4 12 24
use welltap_svt  __well_tap__102
timestamp 1730814361
transform 1 0 104 0 -1 2652
box 8 4 12 24
use welltap_svt  __well_tap__104
timestamp 1730814361
transform 1 0 104 0 1 2668
box 8 4 12 24
use welltap_svt  __well_tap__102
timestamp 1730814361
transform 1 0 104 0 -1 2652
box 8 4 12 24
use welltap_svt  __well_tap__104
timestamp 1730814361
transform 1 0 104 0 1 2668
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5172_6
timestamp 1730814361
transform 1 0 600 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5172_6
timestamp 1730814361
transform 1 0 600 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5157_6
timestamp 1730814361
transform 1 0 728 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5160_6
timestamp 1730814361
transform 1 0 696 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5157_6
timestamp 1730814361
transform 1 0 728 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5160_6
timestamp 1730814361
transform 1 0 696 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5158_6
timestamp 1730814361
transform 1 0 848 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5161_6
timestamp 1730814361
transform 1 0 824 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5158_6
timestamp 1730814361
transform 1 0 848 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5161_6
timestamp 1730814361
transform 1 0 824 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5159_6
timestamp 1730814361
transform 1 0 968 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5162_6
timestamp 1730814361
transform 1 0 952 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5159_6
timestamp 1730814361
transform 1 0 968 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5162_6
timestamp 1730814361
transform 1 0 952 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5163_6
timestamp 1730814361
transform 1 0 1072 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5213_6
timestamp 1730814361
transform 1 0 1088 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5163_6
timestamp 1730814361
transform 1 0 1072 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5213_6
timestamp 1730814361
transform 1 0 1088 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5214_6
timestamp 1730814361
transform 1 0 1200 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5217_6
timestamp 1730814361
transform 1 0 1192 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5214_6
timestamp 1730814361
transform 1 0 1200 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5217_6
timestamp 1730814361
transform 1 0 1192 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5215_6
timestamp 1730814361
transform 1 0 1312 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5218_6
timestamp 1730814361
transform 1 0 1304 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5215_6
timestamp 1730814361
transform 1 0 1312 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5218_6
timestamp 1730814361
transform 1 0 1304 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_547_6
timestamp 1730814361
transform 1 0 1416 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5216_6
timestamp 1730814361
transform 1 0 1432 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_547_6
timestamp 1730814361
transform 1 0 1416 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5216_6
timestamp 1730814361
transform 1 0 1432 0 -1 2656
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_532_6
timestamp 1730814361
transform 1 0 1536 0 1 2664
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_532_6
timestamp 1730814361
transform 1 0 1536 0 1 2664
box 7 3 20 38
use welltap_svt  __well_tap__103
timestamp 1730814361
transform 1 0 1624 0 -1 2652
box 8 4 12 24
use welltap_svt  __well_tap__105
timestamp 1730814361
transform 1 0 1624 0 1 2668
box 8 4 12 24
use welltap_svt  __well_tap__236
timestamp 1730814361
transform 1 0 1664 0 1 2612
box 8 4 12 24
use welltap_svt  __well_tap__238
timestamp 1730814361
transform 1 0 1664 0 -1 2684
box 8 4 12 24
use welltap_svt  __well_tap__103
timestamp 1730814361
transform 1 0 1624 0 -1 2652
box 8 4 12 24
use welltap_svt  __well_tap__105
timestamp 1730814361
transform 1 0 1624 0 1 2668
box 8 4 12 24
use welltap_svt  __well_tap__236
timestamp 1730814361
transform 1 0 1664 0 1 2612
box 8 4 12 24
use welltap_svt  __well_tap__238
timestamp 1730814361
transform 1 0 1664 0 -1 2684
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_515_6
timestamp 1730814361
transform 1 0 1992 0 -1 2688
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_515_6
timestamp 1730814361
transform 1 0 1992 0 -1 2688
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_563_6
timestamp 1730814361
transform 1 0 2168 0 -1 2688
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_563_6
timestamp 1730814361
transform 1 0 2168 0 -1 2688
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_517_6
timestamp 1730814361
transform 1 0 2352 0 -1 2688
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_517_6
timestamp 1730814361
transform 1 0 2352 0 -1 2688
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5280_6
timestamp 1730814361
transform 1 0 2544 0 -1 2688
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5280_6
timestamp 1730814361
transform 1 0 2544 0 -1 2688
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5360_6
timestamp 1730814361
transform 1 0 2752 0 -1 2688
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5360_6
timestamp 1730814361
transform 1 0 2752 0 -1 2688
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5345_6
timestamp 1730814361
transform 1 0 2960 0 -1 2688
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5345_6
timestamp 1730814361
transform 1 0 2960 0 -1 2688
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5336_6
timestamp 1730814361
transform 1 0 3152 0 -1 2688
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5336_6
timestamp 1730814361
transform 1 0 3152 0 -1 2688
box 7 3 20 38
use welltap_svt  __well_tap__237
timestamp 1730814361
transform 1 0 3184 0 1 2612
box 8 4 12 24
use welltap_svt  __well_tap__239
timestamp 1730814361
transform 1 0 3184 0 -1 2684
box 8 4 12 24
use welltap_svt  __well_tap__237
timestamp 1730814361
transform 1 0 3184 0 1 2612
box 8 4 12 24
use welltap_svt  __well_tap__239
timestamp 1730814361
transform 1 0 3184 0 -1 2684
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5165_6
timestamp 1730814361
transform 1 0 128 0 -1 2756
box 7 3 20 38
use welltap_svt  __well_tap__106
timestamp 1730814361
transform 1 0 104 0 -1 2752
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5165_6
timestamp 1730814361
transform 1 0 128 0 -1 2756
box 7 3 20 38
use welltap_svt  __well_tap__106
timestamp 1730814361
transform 1 0 104 0 -1 2752
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5166_6
timestamp 1730814361
transform 1 0 256 0 -1 2756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5166_6
timestamp 1730814361
transform 1 0 256 0 -1 2756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5167_6
timestamp 1730814361
transform 1 0 424 0 -1 2756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5167_6
timestamp 1730814361
transform 1 0 424 0 -1 2756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5164_6
timestamp 1730814361
transform 1 0 616 0 -1 2756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5164_6
timestamp 1730814361
transform 1 0 616 0 -1 2756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_534_6
timestamp 1730814361
transform 1 0 832 0 -1 2756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_534_6
timestamp 1730814361
transform 1 0 832 0 -1 2756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_535_6
timestamp 1730814361
transform 1 0 1064 0 -1 2756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_535_6
timestamp 1730814361
transform 1 0 1064 0 -1 2756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_536_6
timestamp 1730814361
transform 1 0 1312 0 -1 2756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_536_6
timestamp 1730814361
transform 1 0 1312 0 -1 2756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_533_6
timestamp 1730814361
transform 1 0 1560 0 -1 2756
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_533_6
timestamp 1730814361
transform 1 0 1560 0 -1 2756
box 7 3 20 38
use welltap_svt  __well_tap__107
timestamp 1730814361
transform 1 0 1624 0 -1 2752
box 8 4 12 24
use welltap_svt  __well_tap__240
timestamp 1730814361
transform 1 0 1664 0 1 2700
box 8 4 12 24
use welltap_svt  __well_tap__107
timestamp 1730814361
transform 1 0 1624 0 -1 2752
box 8 4 12 24
use welltap_svt  __well_tap__240
timestamp 1730814361
transform 1 0 1664 0 1 2700
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_520_6
timestamp 1730814361
transform 1 0 2008 0 1 2696
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_520_6
timestamp 1730814361
transform 1 0 2008 0 1 2696
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_518_6
timestamp 1730814361
transform 1 0 2192 0 1 2696
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_518_6
timestamp 1730814361
transform 1 0 2192 0 1 2696
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_519_6
timestamp 1730814361
transform 1 0 2376 0 1 2696
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_519_6
timestamp 1730814361
transform 1 0 2376 0 1 2696
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5348_6
timestamp 1730814361
transform 1 0 2568 0 1 2696
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5348_6
timestamp 1730814361
transform 1 0 2568 0 1 2696
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5346_6
timestamp 1730814361
transform 1 0 2768 0 1 2696
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5346_6
timestamp 1730814361
transform 1 0 2768 0 1 2696
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5347_6
timestamp 1730814361
transform 1 0 2968 0 1 2696
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5347_6
timestamp 1730814361
transform 1 0 2968 0 1 2696
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5337_6
timestamp 1730814361
transform 1 0 3152 0 1 2696
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5337_6
timestamp 1730814361
transform 1 0 3152 0 1 2696
box 7 3 20 38
use welltap_svt  __well_tap__241
timestamp 1730814361
transform 1 0 3184 0 1 2700
box 8 4 12 24
use welltap_svt  __well_tap__241
timestamp 1730814361
transform 1 0 3184 0 1 2700
box 8 4 12 24
use welltap_svt  __well_tap__108
timestamp 1730814361
transform 1 0 104 0 1 2772
box 8 4 12 24
use welltap_svt  __well_tap__108
timestamp 1730814361
transform 1 0 104 0 1 2772
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5168_6
timestamp 1730814361
transform 1 0 144 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5168_6
timestamp 1730814361
transform 1 0 144 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5169_6
timestamp 1730814361
transform 1 0 272 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5169_6
timestamp 1730814361
transform 1 0 272 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5170_6
timestamp 1730814361
transform 1 0 392 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5170_6
timestamp 1730814361
transform 1 0 392 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5171_6
timestamp 1730814361
transform 1 0 512 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5171_6
timestamp 1730814361
transform 1 0 512 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_537_6
timestamp 1730814361
transform 1 0 632 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_537_6
timestamp 1730814361
transform 1 0 632 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_538_6
timestamp 1730814361
transform 1 0 744 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_538_6
timestamp 1730814361
transform 1 0 744 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_539_6
timestamp 1730814361
transform 1 0 856 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_539_6
timestamp 1730814361
transform 1 0 856 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_540_6
timestamp 1730814361
transform 1 0 976 0 1 2768
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_540_6
timestamp 1730814361
transform 1 0 976 0 1 2768
box 7 3 20 38
use welltap_svt  __well_tap__109
timestamp 1730814361
transform 1 0 1624 0 1 2772
box 8 4 12 24
use welltap_svt  __well_tap__242
timestamp 1730814361
transform 1 0 1664 0 -1 2776
box 8 4 12 24
use welltap_svt  __well_tap__244
timestamp 1730814361
transform 1 0 1664 0 1 2784
box 8 4 12 24
use welltap_svt  __well_tap__109
timestamp 1730814361
transform 1 0 1624 0 1 2772
box 8 4 12 24
use welltap_svt  __well_tap__242
timestamp 1730814361
transform 1 0 1664 0 -1 2776
box 8 4 12 24
use welltap_svt  __well_tap__244
timestamp 1730814361
transform 1 0 1664 0 1 2784
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_521_6
timestamp 1730814361
transform 1 0 2032 0 -1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_521_6
timestamp 1730814361
transform 1 0 2032 0 -1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_524_6
timestamp 1730814361
transform 1 0 2120 0 1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_524_6
timestamp 1730814361
transform 1 0 2120 0 1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_522_6
timestamp 1730814361
transform 1 0 2200 0 -1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_522_6
timestamp 1730814361
transform 1 0 2200 0 -1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_525_6
timestamp 1730814361
transform 1 0 2296 0 1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_525_6
timestamp 1730814361
transform 1 0 2296 0 1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_523_6
timestamp 1730814361
transform 1 0 2368 0 -1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_523_6
timestamp 1730814361
transform 1 0 2368 0 -1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_526_6
timestamp 1730814361
transform 1 0 2472 0 1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_526_6
timestamp 1730814361
transform 1 0 2472 0 1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5349_6
timestamp 1730814361
transform 1 0 2528 0 -1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5349_6
timestamp 1730814361
transform 1 0 2528 0 -1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5352_6
timestamp 1730814361
transform 1 0 2648 0 1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5352_6
timestamp 1730814361
transform 1 0 2648 0 1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5350_6
timestamp 1730814361
transform 1 0 2696 0 -1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5350_6
timestamp 1730814361
transform 1 0 2696 0 -1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5353_6
timestamp 1730814361
transform 1 0 2824 0 1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5353_6
timestamp 1730814361
transform 1 0 2824 0 1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5351_6
timestamp 1730814361
transform 1 0 2864 0 -1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5351_6
timestamp 1730814361
transform 1 0 2864 0 -1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5354_6
timestamp 1730814361
transform 1 0 3000 0 1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5354_6
timestamp 1730814361
transform 1 0 3000 0 1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5338_6
timestamp 1730814361
transform 1 0 3152 0 1 2780
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5338_6
timestamp 1730814361
transform 1 0 3152 0 1 2780
box 7 3 20 38
use welltap_svt  __well_tap__243
timestamp 1730814361
transform 1 0 3184 0 -1 2776
box 8 4 12 24
use welltap_svt  __well_tap__245
timestamp 1730814361
transform 1 0 3184 0 1 2784
box 8 4 12 24
use welltap_svt  __well_tap__243
timestamp 1730814361
transform 1 0 3184 0 -1 2776
box 8 4 12 24
use welltap_svt  __well_tap__245
timestamp 1730814361
transform 1 0 3184 0 1 2784
box 8 4 12 24
use welltap_svt  __well_tap__110
timestamp 1730814361
transform 1 0 104 0 -1 2852
box 8 4 12 24
use welltap_svt  __well_tap__110
timestamp 1730814361
transform 1 0 104 0 -1 2852
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5156_6
timestamp 1730814361
transform 1 0 248 0 -1 2856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5156_6
timestamp 1730814361
transform 1 0 248 0 -1 2856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5173_6
timestamp 1730814361
transform 1 0 408 0 -1 2856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5173_6
timestamp 1730814361
transform 1 0 408 0 -1 2856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5174_6
timestamp 1730814361
transform 1 0 552 0 -1 2856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5174_6
timestamp 1730814361
transform 1 0 552 0 -1 2856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_541_6
timestamp 1730814361
transform 1 0 688 0 -1 2856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_541_6
timestamp 1730814361
transform 1 0 688 0 -1 2856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_542_6
timestamp 1730814361
transform 1 0 816 0 -1 2856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_542_6
timestamp 1730814361
transform 1 0 816 0 -1 2856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_543_6
timestamp 1730814361
transform 1 0 944 0 -1 2856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_543_6
timestamp 1730814361
transform 1 0 944 0 -1 2856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_544_6
timestamp 1730814361
transform 1 0 1080 0 -1 2856
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_544_6
timestamp 1730814361
transform 1 0 1080 0 -1 2856
box 7 3 20 38
use welltap_svt  __well_tap__111
timestamp 1730814361
transform 1 0 1624 0 -1 2852
box 8 4 12 24
use welltap_svt  __well_tap__246
timestamp 1730814361
transform 1 0 1664 0 -1 2864
box 8 4 12 24
use welltap_svt  __well_tap__111
timestamp 1730814361
transform 1 0 1624 0 -1 2852
box 8 4 12 24
use welltap_svt  __well_tap__246
timestamp 1730814361
transform 1 0 1664 0 -1 2864
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_527_6
timestamp 1730814361
transform 1 0 2200 0 -1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_527_6
timestamp 1730814361
transform 1 0 2200 0 -1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_528_6
timestamp 1730814361
transform 1 0 2368 0 -1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_528_6
timestamp 1730814361
transform 1 0 2368 0 -1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_529_6
timestamp 1730814361
transform 1 0 2528 0 -1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_529_6
timestamp 1730814361
transform 1 0 2528 0 -1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5355_6
timestamp 1730814361
transform 1 0 2672 0 -1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5355_6
timestamp 1730814361
transform 1 0 2672 0 -1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5356_6
timestamp 1730814361
transform 1 0 2816 0 -1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5356_6
timestamp 1730814361
transform 1 0 2816 0 -1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5357_6
timestamp 1730814361
transform 1 0 2960 0 -1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5357_6
timestamp 1730814361
transform 1 0 2960 0 -1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5359_6
timestamp 1730814361
transform 1 0 3104 0 -1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5359_6
timestamp 1730814361
transform 1 0 3104 0 -1 2868
box 7 3 20 38
use welltap_svt  __well_tap__247
timestamp 1730814361
transform 1 0 3184 0 -1 2864
box 8 4 12 24
use welltap_svt  __well_tap__247
timestamp 1730814361
transform 1 0 3184 0 -1 2864
box 8 4 12 24
use welltap_svt  __well_tap__112
timestamp 1730814361
transform 1 0 104 0 1 2868
box 8 4 12 24
use welltap_svt  __well_tap__114
timestamp 1730814361
transform 1 0 104 0 -1 2940
box 8 4 12 24
use welltap_svt  __well_tap__112
timestamp 1730814361
transform 1 0 104 0 1 2868
box 8 4 12 24
use welltap_svt  __well_tap__114
timestamp 1730814361
transform 1 0 104 0 -1 2940
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5175_6
timestamp 1730814361
transform 1 0 328 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5175_6
timestamp 1730814361
transform 1 0 328 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5179_6
timestamp 1730814361
transform 1 0 432 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5179_6
timestamp 1730814361
transform 1 0 432 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5176_6
timestamp 1730814361
transform 1 0 464 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5176_6
timestamp 1730814361
transform 1 0 464 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5177_6
timestamp 1730814361
transform 1 0 616 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5180_6
timestamp 1730814361
transform 1 0 592 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5177_6
timestamp 1730814361
transform 1 0 616 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5180_6
timestamp 1730814361
transform 1 0 592 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5181_6
timestamp 1730814361
transform 1 0 752 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5181_6
timestamp 1730814361
transform 1 0 752 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5178_6
timestamp 1730814361
transform 1 0 784 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5178_6
timestamp 1730814361
transform 1 0 784 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_548_6
timestamp 1730814361
transform 1 0 920 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_548_6
timestamp 1730814361
transform 1 0 920 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_545_6
timestamp 1730814361
transform 1 0 968 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_545_6
timestamp 1730814361
transform 1 0 968 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_549_6
timestamp 1730814361
transform 1 0 1088 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_549_6
timestamp 1730814361
transform 1 0 1088 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_546_6
timestamp 1730814361
transform 1 0 1168 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_546_6
timestamp 1730814361
transform 1 0 1168 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_550_6
timestamp 1730814361
transform 1 0 1256 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_550_6
timestamp 1730814361
transform 1 0 1256 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_531_6
timestamp 1730814361
transform 1 0 1376 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_551_6
timestamp 1730814361
transform 1 0 1432 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_531_6
timestamp 1730814361
transform 1 0 1376 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_551_6
timestamp 1730814361
transform 1 0 1432 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_595_6
timestamp 1730814361
transform 1 0 1592 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5110_6
timestamp 1730814361
transform 1 0 1584 0 1 2864
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_595_6
timestamp 1730814361
transform 1 0 1592 0 -1 2944
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5110_6
timestamp 1730814361
transform 1 0 1584 0 1 2864
box 7 3 20 38
use welltap_svt  __well_tap__113
timestamp 1730814361
transform 1 0 1624 0 1 2868
box 8 4 12 24
use welltap_svt  __well_tap__115
timestamp 1730814361
transform 1 0 1624 0 -1 2940
box 8 4 12 24
use welltap_svt  __well_tap__248
timestamp 1730814361
transform 1 0 1664 0 1 2872
box 8 4 12 24
use welltap_svt  __well_tap__250
timestamp 1730814361
transform 1 0 1664 0 -1 2944
box 8 4 12 24
use welltap_svt  __well_tap__113
timestamp 1730814361
transform 1 0 1624 0 1 2868
box 8 4 12 24
use welltap_svt  __well_tap__115
timestamp 1730814361
transform 1 0 1624 0 -1 2940
box 8 4 12 24
use welltap_svt  __well_tap__248
timestamp 1730814361
transform 1 0 1664 0 1 2872
box 8 4 12 24
use welltap_svt  __well_tap__250
timestamp 1730814361
transform 1 0 1664 0 -1 2944
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_596_6
timestamp 1730814361
transform 1 0 1688 0 -1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_596_6
timestamp 1730814361
transform 1 0 1688 0 -1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_597_6
timestamp 1730814361
transform 1 0 1928 0 -1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_597_6
timestamp 1730814361
transform 1 0 1928 0 -1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5362_6
timestamp 1730814361
transform 1 0 2216 0 -1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5362_6
timestamp 1730814361
transform 1 0 2216 0 -1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_530_6
timestamp 1730814361
transform 1 0 2288 0 1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_530_6
timestamp 1730814361
transform 1 0 2288 0 1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5344_6
timestamp 1730814361
transform 1 0 2544 0 1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5363_6
timestamp 1730814361
transform 1 0 2512 0 -1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5344_6
timestamp 1730814361
transform 1 0 2544 0 1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5363_6
timestamp 1730814361
transform 1 0 2512 0 -1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5361_6
timestamp 1730814361
transform 1 0 2808 0 1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5364_6
timestamp 1730814361
transform 1 0 2816 0 -1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5361_6
timestamp 1730814361
transform 1 0 2808 0 1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5364_6
timestamp 1730814361
transform 1 0 2816 0 -1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5358_6
timestamp 1730814361
transform 1 0 3072 0 1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5358_6
timestamp 1730814361
transform 1 0 3072 0 1 2868
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5339_6
timestamp 1730814361
transform 1 0 3128 0 -1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5339_6
timestamp 1730814361
transform 1 0 3128 0 -1 2948
box 7 3 20 38
use welltap_svt  __well_tap__249
timestamp 1730814361
transform 1 0 3184 0 1 2872
box 8 4 12 24
use welltap_svt  __well_tap__251
timestamp 1730814361
transform 1 0 3184 0 -1 2944
box 8 4 12 24
use welltap_svt  __well_tap__249
timestamp 1730814361
transform 1 0 3184 0 1 2872
box 8 4 12 24
use welltap_svt  __well_tap__251
timestamp 1730814361
transform 1 0 3184 0 -1 2944
box 8 4 12 24
use welltap_svt  __well_tap__116
timestamp 1730814361
transform 1 0 104 0 1 2956
box 8 4 12 24
use welltap_svt  __well_tap__116
timestamp 1730814361
transform 1 0 104 0 1 2956
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5182_6
timestamp 1730814361
transform 1 0 512 0 1 2952
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5182_6
timestamp 1730814361
transform 1 0 512 0 1 2952
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5183_6
timestamp 1730814361
transform 1 0 640 0 1 2952
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5183_6
timestamp 1730814361
transform 1 0 640 0 1 2952
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5184_6
timestamp 1730814361
transform 1 0 776 0 1 2952
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5184_6
timestamp 1730814361
transform 1 0 776 0 1 2952
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5185_6
timestamp 1730814361
transform 1 0 912 0 1 2952
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5185_6
timestamp 1730814361
transform 1 0 912 0 1 2952
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_552_6
timestamp 1730814361
transform 1 0 1048 0 1 2952
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_552_6
timestamp 1730814361
transform 1 0 1048 0 1 2952
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_553_6
timestamp 1730814361
transform 1 0 1184 0 1 2952
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_553_6
timestamp 1730814361
transform 1 0 1184 0 1 2952
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_554_6
timestamp 1730814361
transform 1 0 1328 0 1 2952
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_554_6
timestamp 1730814361
transform 1 0 1328 0 1 2952
box 7 3 20 38
use welltap_svt  __well_tap__117
timestamp 1730814361
transform 1 0 1624 0 1 2956
box 8 4 12 24
use welltap_svt  __well_tap__252
timestamp 1730814361
transform 1 0 1664 0 1 2952
box 8 4 12 24
use welltap_svt  __well_tap__117
timestamp 1730814361
transform 1 0 1624 0 1 2956
box 8 4 12 24
use welltap_svt  __well_tap__252
timestamp 1730814361
transform 1 0 1664 0 1 2952
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_598_6
timestamp 1730814361
transform 1 0 1696 0 1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_598_6
timestamp 1730814361
transform 1 0 1696 0 1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_599_6
timestamp 1730814361
transform 1 0 1896 0 1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_599_6
timestamp 1730814361
transform 1 0 1896 0 1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5100_6
timestamp 1730814361
transform 1 0 2120 0 1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5100_6
timestamp 1730814361
transform 1 0 2120 0 1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5365_6
timestamp 1730814361
transform 1 0 2360 0 1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5365_6
timestamp 1730814361
transform 1 0 2360 0 1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5366_6
timestamp 1730814361
transform 1 0 2616 0 1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5366_6
timestamp 1730814361
transform 1 0 2616 0 1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5367_6
timestamp 1730814361
transform 1 0 2880 0 1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5367_6
timestamp 1730814361
transform 1 0 2880 0 1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5340_6
timestamp 1730814361
transform 1 0 3152 0 1 2948
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5340_6
timestamp 1730814361
transform 1 0 3152 0 1 2948
box 7 3 20 38
use welltap_svt  __well_tap__253
timestamp 1730814361
transform 1 0 3184 0 1 2952
box 8 4 12 24
use welltap_svt  __well_tap__253
timestamp 1730814361
transform 1 0 3184 0 1 2952
box 8 4 12 24
use welltap_svt  __well_tap__118
timestamp 1730814361
transform 1 0 104 0 -1 3032
box 8 4 12 24
use welltap_svt  __well_tap__118
timestamp 1730814361
transform 1 0 104 0 -1 3032
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5186_6
timestamp 1730814361
transform 1 0 616 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5186_6
timestamp 1730814361
transform 1 0 616 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5126_6
timestamp 1730814361
transform 1 0 696 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5126_6
timestamp 1730814361
transform 1 0 696 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5187_6
timestamp 1730814361
transform 1 0 776 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5187_6
timestamp 1730814361
transform 1 0 776 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5127_6
timestamp 1730814361
transform 1 0 824 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5127_6
timestamp 1730814361
transform 1 0 824 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5141_6
timestamp 1730814361
transform 1 0 920 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5141_6
timestamp 1730814361
transform 1 0 920 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5128_6
timestamp 1730814361
transform 1 0 952 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5128_6
timestamp 1730814361
transform 1 0 952 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_555_6
timestamp 1730814361
transform 1 0 1056 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_555_6
timestamp 1730814361
transform 1 0 1056 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5129_6
timestamp 1730814361
transform 1 0 1072 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5129_6
timestamp 1730814361
transform 1 0 1072 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_556_6
timestamp 1730814361
transform 1 0 1184 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_556_6
timestamp 1730814361
transform 1 0 1184 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_559_6
timestamp 1730814361
transform 1 0 1192 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_559_6
timestamp 1730814361
transform 1 0 1192 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_557_6
timestamp 1730814361
transform 1 0 1304 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_560_6
timestamp 1730814361
transform 1 0 1304 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_557_6
timestamp 1730814361
transform 1 0 1304 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_560_6
timestamp 1730814361
transform 1 0 1304 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_558_6
timestamp 1730814361
transform 1 0 1432 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_561_6
timestamp 1730814361
transform 1 0 1416 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_558_6
timestamp 1730814361
transform 1 0 1432 0 -1 3036
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_561_6
timestamp 1730814361
transform 1 0 1416 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_562_6
timestamp 1730814361
transform 1 0 1536 0 1 3044
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_562_6
timestamp 1730814361
transform 1 0 1536 0 1 3044
box 7 3 20 38
use welltap_svt  __well_tap__119
timestamp 1730814361
transform 1 0 1624 0 -1 3032
box 8 4 12 24
use welltap_svt  __well_tap__254
timestamp 1730814361
transform 1 0 1664 0 -1 3024
box 8 4 12 24
use welltap_svt  __well_tap__256
timestamp 1730814361
transform 1 0 1664 0 1 3032
box 8 4 12 24
use welltap_svt  __well_tap__119
timestamp 1730814361
transform 1 0 1624 0 -1 3032
box 8 4 12 24
use welltap_svt  __well_tap__254
timestamp 1730814361
transform 1 0 1664 0 -1 3024
box 8 4 12 24
use welltap_svt  __well_tap__256
timestamp 1730814361
transform 1 0 1664 0 1 3032
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5101_6
timestamp 1730814361
transform 1 0 1784 0 -1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5101_6
timestamp 1730814361
transform 1 0 1784 0 -1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5104_6
timestamp 1730814361
transform 1 0 1864 0 1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5104_6
timestamp 1730814361
transform 1 0 1864 0 1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5102_6
timestamp 1730814361
transform 1 0 1952 0 -1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5102_6
timestamp 1730814361
transform 1 0 1952 0 -1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5105_6
timestamp 1730814361
transform 1 0 2104 0 1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5105_6
timestamp 1730814361
transform 1 0 2104 0 1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5103_6
timestamp 1730814361
transform 1 0 2120 0 -1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5103_6
timestamp 1730814361
transform 1 0 2120 0 -1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5368_6
timestamp 1730814361
transform 1 0 2280 0 -1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5368_6
timestamp 1730814361
transform 1 0 2280 0 -1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5106_6
timestamp 1730814361
transform 1 0 2360 0 1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5106_6
timestamp 1730814361
transform 1 0 2360 0 1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5369_6
timestamp 1730814361
transform 1 0 2448 0 -1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5369_6
timestamp 1730814361
transform 1 0 2448 0 -1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5370_6
timestamp 1730814361
transform 1 0 2616 0 -1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5371_6
timestamp 1730814361
transform 1 0 2624 0 1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5370_6
timestamp 1730814361
transform 1 0 2616 0 -1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5371_6
timestamp 1730814361
transform 1 0 2624 0 1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5372_6
timestamp 1730814361
transform 1 0 2896 0 1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5372_6
timestamp 1730814361
transform 1 0 2896 0 1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5341_6
timestamp 1730814361
transform 1 0 3152 0 1 3028
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5341_6
timestamp 1730814361
transform 1 0 3152 0 1 3028
box 7 3 20 38
use welltap_svt  __well_tap__255
timestamp 1730814361
transform 1 0 3184 0 -1 3024
box 8 4 12 24
use welltap_svt  __well_tap__257
timestamp 1730814361
transform 1 0 3184 0 1 3032
box 8 4 12 24
use welltap_svt  __well_tap__255
timestamp 1730814361
transform 1 0 3184 0 -1 3024
box 8 4 12 24
use welltap_svt  __well_tap__257
timestamp 1730814361
transform 1 0 3184 0 1 3032
box 8 4 12 24
use welltap_svt  __well_tap__120
timestamp 1730814361
transform 1 0 104 0 1 3048
box 8 4 12 24
use welltap_svt  __well_tap__122
timestamp 1730814361
transform 1 0 104 0 -1 3124
box 8 4 12 24
use welltap_svt  __well_tap__120
timestamp 1730814361
transform 1 0 104 0 1 3048
box 8 4 12 24
use welltap_svt  __well_tap__122
timestamp 1730814361
transform 1 0 104 0 -1 3124
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5130_6
timestamp 1730814361
transform 1 0 800 0 -1 3128
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5130_6
timestamp 1730814361
transform 1 0 800 0 -1 3128
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_516_6
timestamp 1730814361
transform 1 0 1072 0 -1 3128
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_516_6
timestamp 1730814361
transform 1 0 1072 0 -1 3128
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5109_6
timestamp 1730814361
transform 1 0 1344 0 -1 3128
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5109_6
timestamp 1730814361
transform 1 0 1344 0 -1 3128
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_594_6
timestamp 1730814361
transform 1 0 1592 0 -1 3128
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_594_6
timestamp 1730814361
transform 1 0 1592 0 -1 3128
box 7 3 20 38
use welltap_svt  __well_tap__121
timestamp 1730814361
transform 1 0 1624 0 1 3048
box 8 4 12 24
use welltap_svt  __well_tap__123
timestamp 1730814361
transform 1 0 1624 0 -1 3124
box 8 4 12 24
use welltap_svt  __well_tap__258
timestamp 1730814361
transform 1 0 1664 0 -1 3104
box 8 4 12 24
use welltap_svt  __well_tap__121
timestamp 1730814361
transform 1 0 1624 0 1 3048
box 8 4 12 24
use welltap_svt  __well_tap__123
timestamp 1730814361
transform 1 0 1624 0 -1 3124
box 8 4 12 24
use welltap_svt  __well_tap__258
timestamp 1730814361
transform 1 0 1664 0 -1 3104
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5107_6
timestamp 1730814361
transform 1 0 1952 0 -1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5107_6
timestamp 1730814361
transform 1 0 1952 0 -1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5108_6
timestamp 1730814361
transform 1 0 2176 0 -1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5108_6
timestamp 1730814361
transform 1 0 2176 0 -1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5329_6
timestamp 1730814361
transform 1 0 2408 0 -1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5329_6
timestamp 1730814361
transform 1 0 2408 0 -1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5373_6
timestamp 1730814361
transform 1 0 2648 0 -1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5373_6
timestamp 1730814361
transform 1 0 2648 0 -1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5374_6
timestamp 1730814361
transform 1 0 2896 0 -1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5374_6
timestamp 1730814361
transform 1 0 2896 0 -1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5342_6
timestamp 1730814361
transform 1 0 3152 0 -1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5342_6
timestamp 1730814361
transform 1 0 3152 0 -1 3108
box 7 3 20 38
use welltap_svt  __well_tap__259
timestamp 1730814361
transform 1 0 3184 0 -1 3104
box 8 4 12 24
use welltap_svt  __well_tap__259
timestamp 1730814361
transform 1 0 3184 0 -1 3104
box 8 4 12 24
use welltap_svt  __well_tap__260
timestamp 1730814361
transform 1 0 1664 0 1 3112
box 8 4 12 24
use welltap_svt  __well_tap__262
timestamp 1730814361
transform 1 0 1664 0 -1 3184
box 8 4 12 24
use welltap_svt  __well_tap__260
timestamp 1730814361
transform 1 0 1664 0 1 3112
box 8 4 12 24
use welltap_svt  __well_tap__262
timestamp 1730814361
transform 1 0 1664 0 -1 3184
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5111_6
timestamp 1730814361
transform 1 0 1688 0 1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5111_6
timestamp 1730814361
transform 1 0 1688 0 1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5112_6
timestamp 1730814361
transform 1 0 1856 0 1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5114_6
timestamp 1730814361
transform 1 0 1840 0 -1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5112_6
timestamp 1730814361
transform 1 0 1856 0 1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5114_6
timestamp 1730814361
transform 1 0 1840 0 -1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5113_6
timestamp 1730814361
transform 1 0 2016 0 1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5115_6
timestamp 1730814361
transform 1 0 2032 0 -1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5113_6
timestamp 1730814361
transform 1 0 2016 0 1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5115_6
timestamp 1730814361
transform 1 0 2032 0 -1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5314_6
timestamp 1730814361
transform 1 0 2176 0 1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5314_6
timestamp 1730814361
transform 1 0 2176 0 1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5116_6
timestamp 1730814361
transform 1 0 2240 0 -1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5116_6
timestamp 1730814361
transform 1 0 2240 0 -1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5315_6
timestamp 1730814361
transform 1 0 2336 0 1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5315_6
timestamp 1730814361
transform 1 0 2336 0 1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5317_6
timestamp 1730814361
transform 1 0 2456 0 -1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5317_6
timestamp 1730814361
transform 1 0 2456 0 -1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5316_6
timestamp 1730814361
transform 1 0 2504 0 1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5316_6
timestamp 1730814361
transform 1 0 2504 0 1 3108
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5318_6
timestamp 1730814361
transform 1 0 2688 0 -1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5318_6
timestamp 1730814361
transform 1 0 2688 0 -1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5319_6
timestamp 1730814361
transform 1 0 2928 0 -1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5319_6
timestamp 1730814361
transform 1 0 2928 0 -1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5343_6
timestamp 1730814361
transform 1 0 3152 0 -1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5343_6
timestamp 1730814361
transform 1 0 3152 0 -1 3188
box 7 3 20 38
use welltap_svt  __well_tap__261
timestamp 1730814361
transform 1 0 3184 0 1 3112
box 8 4 12 24
use welltap_svt  __well_tap__263
timestamp 1730814361
transform 1 0 3184 0 -1 3184
box 8 4 12 24
use welltap_svt  __well_tap__261
timestamp 1730814361
transform 1 0 3184 0 1 3112
box 8 4 12 24
use welltap_svt  __well_tap__263
timestamp 1730814361
transform 1 0 3184 0 -1 3184
box 8 4 12 24
use welltap_svt  __well_tap__264
timestamp 1730814361
transform 1 0 1664 0 1 3192
box 8 4 12 24
use welltap_svt  __well_tap__264
timestamp 1730814361
transform 1 0 1664 0 1 3192
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5117_6
timestamp 1730814361
transform 1 0 1992 0 1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5117_6
timestamp 1730814361
transform 1 0 1992 0 1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5118_6
timestamp 1730814361
transform 1 0 2168 0 1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5120_6
timestamp 1730814361
transform 1 0 2144 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5118_6
timestamp 1730814361
transform 1 0 2168 0 1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5120_6
timestamp 1730814361
transform 1 0 2144 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5121_6
timestamp 1730814361
transform 1 0 2280 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5121_6
timestamp 1730814361
transform 1 0 2280 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5119_6
timestamp 1730814361
transform 1 0 2352 0 1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5119_6
timestamp 1730814361
transform 1 0 2352 0 1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5122_6
timestamp 1730814361
transform 1 0 2416 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5122_6
timestamp 1730814361
transform 1 0 2416 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5320_6
timestamp 1730814361
transform 1 0 2536 0 1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5320_6
timestamp 1730814361
transform 1 0 2536 0 1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5123_6
timestamp 1730814361
transform 1 0 2560 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5123_6
timestamp 1730814361
transform 1 0 2560 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5321_6
timestamp 1730814361
transform 1 0 2720 0 1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5323_6
timestamp 1730814361
transform 1 0 2704 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5321_6
timestamp 1730814361
transform 1 0 2720 0 1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5323_6
timestamp 1730814361
transform 1 0 2704 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5324_6
timestamp 1730814361
transform 1 0 2848 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5324_6
timestamp 1730814361
transform 1 0 2848 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5322_6
timestamp 1730814361
transform 1 0 2912 0 1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5322_6
timestamp 1730814361
transform 1 0 2912 0 1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5325_6
timestamp 1730814361
transform 1 0 2992 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5325_6
timestamp 1730814361
transform 1 0 2992 0 -1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5327_6
timestamp 1730814361
transform 1 0 3104 0 1 3188
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5327_6
timestamp 1730814361
transform 1 0 3104 0 1 3188
box 7 3 20 38
use welltap_svt  __well_tap__265
timestamp 1730814361
transform 1 0 3184 0 1 3192
box 8 4 12 24
use welltap_svt  __well_tap__265
timestamp 1730814361
transform 1 0 3184 0 1 3192
box 8 4 12 24
use welltap_svt  __well_tap__266
timestamp 1730814361
transform 1 0 1664 0 -1 3264
box 8 4 12 24
use welltap_svt  __well_tap__268
timestamp 1730814361
transform 1 0 1664 0 1 3272
box 8 4 12 24
use welltap_svt  __well_tap__266
timestamp 1730814361
transform 1 0 1664 0 -1 3264
box 8 4 12 24
use welltap_svt  __well_tap__268
timestamp 1730814361
transform 1 0 1664 0 1 3272
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  tielo_5326_6
timestamp 1730814361
transform 1 0 3048 0 1 3268
box 7 3 20 38
use _0_0std_0_0cells_0_0TIELOX1  tielo_5326_6
timestamp 1730814361
transform 1 0 3048 0 1 3268
box 7 3 20 38
use welltap_svt  __well_tap__267
timestamp 1730814361
transform 1 0 3184 0 -1 3264
box 8 4 12 24
use welltap_svt  __well_tap__269
timestamp 1730814361
transform 1 0 3184 0 1 3272
box 8 4 12 24
use welltap_svt  __well_tap__267
timestamp 1730814361
transform 1 0 3184 0 -1 3264
box 8 4 12 24
use welltap_svt  __well_tap__269
timestamp 1730814361
transform 1 0 3184 0 1 3272
box 8 4 12 24
<< end >>
