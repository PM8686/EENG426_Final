magic
tech sky130l
timestamp 1730768254
<< m1 >>
rect 832 1359 836 1399
rect 1560 1359 1564 1399
rect 944 1291 948 1331
rect 928 915 932 955
rect 928 695 932 735
rect 424 619 428 659
rect 264 455 268 495
rect 944 455 948 495
<< m2c >>
rect 232 1729 236 1733
rect 368 1729 372 1733
rect 504 1729 508 1733
rect 640 1729 644 1733
rect 776 1729 780 1733
rect 111 1725 115 1729
rect 1719 1725 1723 1729
rect 111 1707 115 1711
rect 1719 1707 1723 1711
rect 111 1641 115 1645
rect 1719 1641 1723 1645
rect 111 1623 115 1627
rect 1719 1623 1723 1627
rect 312 1619 316 1623
rect 448 1619 452 1623
rect 584 1619 588 1623
rect 720 1619 724 1623
rect 856 1619 860 1623
rect 696 1505 700 1509
rect 832 1505 836 1509
rect 968 1505 972 1509
rect 1112 1505 1116 1509
rect 1256 1505 1260 1509
rect 1400 1505 1404 1509
rect 1536 1505 1540 1509
rect 1672 1505 1676 1509
rect 111 1501 115 1505
rect 1719 1501 1723 1505
rect 111 1483 115 1487
rect 1719 1483 1723 1487
rect 111 1421 115 1425
rect 1719 1421 1723 1425
rect 111 1403 115 1407
rect 1719 1403 1723 1407
rect 672 1399 676 1403
rect 808 1399 812 1403
rect 832 1399 836 1403
rect 952 1399 956 1403
rect 1096 1399 1100 1403
rect 1240 1399 1244 1403
rect 1392 1399 1396 1403
rect 1536 1399 1540 1403
rect 1560 1399 1564 1403
rect 1672 1399 1676 1403
rect 832 1355 836 1359
rect 1560 1355 1564 1359
rect 944 1331 948 1335
rect 232 1285 236 1289
rect 400 1285 404 1289
rect 616 1285 620 1289
rect 848 1285 852 1289
rect 944 1287 948 1291
rect 1096 1285 1100 1289
rect 1352 1285 1356 1289
rect 1616 1285 1620 1289
rect 111 1281 115 1285
rect 1719 1281 1723 1285
rect 111 1263 115 1267
rect 1719 1263 1723 1267
rect 111 1193 115 1197
rect 1719 1193 1723 1197
rect 111 1175 115 1179
rect 1719 1175 1723 1179
rect 232 1171 236 1175
rect 472 1171 476 1175
rect 744 1171 748 1175
rect 1032 1171 1036 1175
rect 1328 1171 1332 1175
rect 1624 1171 1628 1175
rect 288 1073 292 1077
rect 512 1073 516 1077
rect 768 1073 772 1077
rect 1048 1073 1052 1077
rect 1344 1073 1348 1077
rect 1640 1073 1644 1077
rect 111 1069 115 1073
rect 1719 1069 1723 1073
rect 111 1051 115 1055
rect 1719 1051 1723 1055
rect 111 977 115 981
rect 1719 977 1723 981
rect 111 959 115 963
rect 1719 959 1723 963
rect 584 955 588 959
rect 736 955 740 959
rect 904 955 908 959
rect 928 955 932 959
rect 1080 955 1084 959
rect 1272 955 1276 959
rect 1472 955 1476 959
rect 1672 955 1676 959
rect 928 911 932 915
rect 856 845 860 849
rect 1008 845 1012 849
rect 1168 845 1172 849
rect 1336 845 1340 849
rect 1504 845 1508 849
rect 1672 845 1676 849
rect 111 841 115 845
rect 1719 841 1723 845
rect 111 823 115 827
rect 1719 823 1723 827
rect 111 757 115 761
rect 1719 757 1723 761
rect 111 739 115 743
rect 1719 739 1723 743
rect 768 735 772 739
rect 904 735 908 739
rect 928 735 932 739
rect 1048 735 1052 739
rect 1192 735 1196 739
rect 1344 735 1348 739
rect 1504 735 1508 739
rect 1672 735 1676 739
rect 928 691 932 695
rect 424 659 428 663
rect 344 613 348 617
rect 424 615 428 619
rect 528 613 532 617
rect 728 613 732 617
rect 944 613 948 617
rect 1176 613 1180 617
rect 1416 613 1420 617
rect 1656 613 1660 617
rect 111 609 115 613
rect 1719 609 1723 613
rect 111 591 115 595
rect 1719 591 1723 595
rect 111 517 115 521
rect 1719 517 1723 521
rect 111 499 115 503
rect 1719 499 1723 503
rect 232 495 236 499
rect 264 495 268 499
rect 416 495 420 499
rect 648 495 652 499
rect 904 495 908 499
rect 944 495 948 499
rect 1168 495 1172 499
rect 1440 495 1444 499
rect 264 451 268 455
rect 944 451 948 455
rect 296 385 300 389
rect 512 385 516 389
rect 728 385 732 389
rect 952 385 956 389
rect 1184 385 1188 389
rect 1424 385 1428 389
rect 1672 385 1676 389
rect 111 381 115 385
rect 1719 381 1723 385
rect 111 363 115 367
rect 1719 363 1723 367
rect 111 301 115 305
rect 1719 301 1723 305
rect 111 283 115 287
rect 1719 283 1723 287
rect 632 279 636 283
rect 832 279 836 283
rect 1040 279 1044 283
rect 1256 279 1260 283
rect 1472 279 1476 283
rect 1672 279 1676 283
rect 584 169 588 173
rect 720 169 724 173
rect 856 169 860 173
rect 992 169 996 173
rect 1128 169 1132 173
rect 1264 169 1268 173
rect 1400 169 1404 173
rect 1672 169 1676 173
rect 111 165 115 169
rect 1719 165 1723 169
rect 111 147 115 151
rect 1719 147 1723 151
<< m2 >>
rect 250 1779 256 1780
rect 250 1775 251 1779
rect 255 1778 256 1779
rect 386 1779 392 1780
rect 255 1776 273 1778
rect 255 1775 256 1776
rect 250 1774 256 1775
rect 386 1775 387 1779
rect 391 1778 392 1779
rect 522 1779 528 1780
rect 391 1776 409 1778
rect 391 1775 392 1776
rect 386 1774 392 1775
rect 522 1775 523 1779
rect 527 1778 528 1779
rect 658 1779 664 1780
rect 527 1776 545 1778
rect 527 1775 528 1776
rect 522 1774 528 1775
rect 658 1775 659 1779
rect 663 1778 664 1779
rect 663 1776 681 1778
rect 663 1775 664 1776
rect 658 1774 664 1775
rect 231 1733 237 1734
rect 110 1729 116 1730
rect 110 1725 111 1729
rect 115 1725 116 1729
rect 231 1729 232 1733
rect 236 1732 237 1733
rect 250 1733 256 1734
rect 250 1732 251 1733
rect 236 1730 251 1732
rect 236 1729 237 1730
rect 231 1728 237 1729
rect 250 1729 251 1730
rect 255 1729 256 1733
rect 250 1728 256 1729
rect 367 1733 373 1734
rect 367 1729 368 1733
rect 372 1732 373 1733
rect 386 1733 392 1734
rect 386 1732 387 1733
rect 372 1730 387 1732
rect 372 1729 373 1730
rect 367 1728 373 1729
rect 386 1729 387 1730
rect 391 1729 392 1733
rect 386 1728 392 1729
rect 503 1733 509 1734
rect 503 1729 504 1733
rect 508 1732 509 1733
rect 522 1733 528 1734
rect 522 1732 523 1733
rect 508 1730 523 1732
rect 508 1729 509 1730
rect 503 1728 509 1729
rect 522 1729 523 1730
rect 527 1729 528 1733
rect 522 1728 528 1729
rect 639 1733 645 1734
rect 639 1729 640 1733
rect 644 1732 645 1733
rect 658 1733 664 1734
rect 658 1732 659 1733
rect 644 1730 659 1732
rect 644 1729 645 1730
rect 639 1728 645 1729
rect 658 1729 659 1730
rect 663 1729 664 1733
rect 658 1728 664 1729
rect 774 1733 781 1734
rect 774 1729 775 1733
rect 780 1729 781 1733
rect 774 1728 781 1729
rect 1718 1729 1724 1730
rect 110 1724 116 1725
rect 134 1727 140 1728
rect 134 1723 135 1727
rect 139 1723 140 1727
rect 134 1722 140 1723
rect 270 1727 276 1728
rect 270 1723 271 1727
rect 275 1723 276 1727
rect 270 1722 276 1723
rect 406 1727 412 1728
rect 406 1723 407 1727
rect 411 1723 412 1727
rect 406 1722 412 1723
rect 542 1727 548 1728
rect 542 1723 543 1727
rect 547 1723 548 1727
rect 542 1722 548 1723
rect 678 1727 684 1728
rect 678 1723 679 1727
rect 683 1723 684 1727
rect 1718 1725 1719 1729
rect 1723 1725 1724 1729
rect 1718 1724 1724 1725
rect 678 1722 684 1723
rect 158 1712 164 1713
rect 110 1711 116 1712
rect 110 1707 111 1711
rect 115 1707 116 1711
rect 158 1708 159 1712
rect 163 1708 164 1712
rect 158 1707 164 1708
rect 294 1712 300 1713
rect 294 1708 295 1712
rect 299 1708 300 1712
rect 294 1707 300 1708
rect 430 1712 436 1713
rect 430 1708 431 1712
rect 435 1708 436 1712
rect 430 1707 436 1708
rect 566 1712 572 1713
rect 566 1708 567 1712
rect 571 1708 572 1712
rect 566 1707 572 1708
rect 702 1712 708 1713
rect 702 1708 703 1712
rect 707 1708 708 1712
rect 702 1707 708 1708
rect 1718 1711 1724 1712
rect 1718 1707 1719 1711
rect 1723 1707 1724 1711
rect 110 1706 116 1707
rect 1718 1706 1724 1707
rect 306 1675 312 1676
rect 306 1671 307 1675
rect 311 1674 312 1675
rect 774 1675 780 1676
rect 774 1674 775 1675
rect 311 1672 775 1674
rect 311 1671 312 1672
rect 306 1670 312 1671
rect 774 1671 775 1672
rect 779 1671 780 1675
rect 774 1670 780 1671
rect 110 1645 116 1646
rect 1718 1645 1724 1646
rect 110 1641 111 1645
rect 115 1641 116 1645
rect 110 1640 116 1641
rect 238 1644 244 1645
rect 238 1640 239 1644
rect 243 1640 244 1644
rect 238 1639 244 1640
rect 374 1644 380 1645
rect 374 1640 375 1644
rect 379 1640 380 1644
rect 374 1639 380 1640
rect 510 1644 516 1645
rect 510 1640 511 1644
rect 515 1640 516 1644
rect 510 1639 516 1640
rect 646 1644 652 1645
rect 646 1640 647 1644
rect 651 1640 652 1644
rect 646 1639 652 1640
rect 782 1644 788 1645
rect 782 1640 783 1644
rect 787 1640 788 1644
rect 1718 1641 1719 1645
rect 1723 1641 1724 1645
rect 1718 1640 1724 1641
rect 782 1639 788 1640
rect 214 1629 220 1630
rect 110 1627 116 1628
rect 110 1623 111 1627
rect 115 1623 116 1627
rect 214 1625 215 1629
rect 219 1625 220 1629
rect 214 1624 220 1625
rect 350 1629 356 1630
rect 350 1625 351 1629
rect 355 1625 356 1629
rect 350 1624 356 1625
rect 486 1629 492 1630
rect 486 1625 487 1629
rect 491 1625 492 1629
rect 486 1624 492 1625
rect 622 1629 628 1630
rect 622 1625 623 1629
rect 627 1625 628 1629
rect 622 1624 628 1625
rect 758 1629 764 1630
rect 758 1625 759 1629
rect 763 1625 764 1629
rect 758 1624 764 1625
rect 1718 1627 1724 1628
rect 110 1622 116 1623
rect 311 1623 317 1624
rect 311 1619 312 1623
rect 316 1622 317 1623
rect 330 1623 336 1624
rect 330 1622 331 1623
rect 316 1620 331 1622
rect 316 1619 317 1620
rect 311 1618 317 1619
rect 330 1619 331 1620
rect 335 1619 336 1623
rect 330 1618 336 1619
rect 447 1623 453 1624
rect 447 1619 448 1623
rect 452 1622 453 1623
rect 466 1623 472 1624
rect 466 1622 467 1623
rect 452 1620 467 1622
rect 452 1619 453 1620
rect 447 1618 453 1619
rect 466 1619 467 1620
rect 471 1619 472 1623
rect 466 1618 472 1619
rect 583 1623 589 1624
rect 583 1619 584 1623
rect 588 1620 589 1623
rect 719 1623 725 1624
rect 588 1619 592 1620
rect 583 1618 587 1619
rect 584 1616 587 1618
rect 586 1615 587 1616
rect 591 1615 592 1619
rect 719 1619 720 1623
rect 724 1622 725 1623
rect 738 1623 744 1624
rect 738 1622 739 1623
rect 724 1620 739 1622
rect 724 1619 725 1620
rect 719 1618 725 1619
rect 738 1619 739 1620
rect 743 1619 744 1623
rect 855 1623 861 1624
rect 855 1622 856 1623
rect 738 1618 744 1619
rect 748 1620 856 1622
rect 586 1614 592 1615
rect 690 1615 696 1616
rect 690 1611 691 1615
rect 695 1614 696 1615
rect 748 1614 750 1620
rect 855 1619 856 1620
rect 860 1619 861 1623
rect 1718 1623 1719 1627
rect 1723 1623 1724 1627
rect 1718 1622 1724 1623
rect 855 1618 861 1619
rect 695 1612 750 1614
rect 695 1611 696 1612
rect 690 1610 696 1611
rect 306 1579 312 1580
rect 306 1575 307 1579
rect 311 1575 312 1579
rect 306 1574 312 1575
rect 330 1579 336 1580
rect 330 1575 331 1579
rect 335 1578 336 1579
rect 466 1579 472 1580
rect 335 1576 353 1578
rect 335 1575 336 1576
rect 330 1574 336 1575
rect 466 1575 467 1579
rect 471 1578 472 1579
rect 586 1579 592 1580
rect 471 1576 489 1578
rect 471 1575 472 1576
rect 466 1574 472 1575
rect 586 1575 587 1579
rect 591 1578 592 1579
rect 738 1579 744 1580
rect 591 1576 625 1578
rect 591 1575 592 1576
rect 586 1574 592 1575
rect 738 1575 739 1579
rect 743 1578 744 1579
rect 743 1576 761 1578
rect 743 1575 744 1576
rect 738 1574 744 1575
rect 690 1555 696 1556
rect 690 1551 691 1555
rect 695 1551 696 1555
rect 690 1550 696 1551
rect 714 1555 720 1556
rect 714 1551 715 1555
rect 719 1554 720 1555
rect 862 1555 868 1556
rect 719 1552 737 1554
rect 719 1551 720 1552
rect 714 1550 720 1551
rect 862 1551 863 1555
rect 867 1554 868 1555
rect 970 1555 976 1556
rect 867 1552 873 1554
rect 867 1551 868 1552
rect 862 1550 868 1551
rect 970 1551 971 1555
rect 975 1554 976 1555
rect 1114 1555 1120 1556
rect 975 1552 1017 1554
rect 975 1551 976 1552
rect 970 1550 976 1551
rect 1114 1551 1115 1555
rect 1119 1554 1120 1555
rect 1418 1555 1424 1556
rect 1119 1552 1161 1554
rect 1119 1551 1120 1552
rect 1114 1550 1120 1551
rect 1394 1551 1400 1552
rect 1394 1547 1395 1551
rect 1399 1547 1400 1551
rect 1418 1551 1419 1555
rect 1423 1554 1424 1555
rect 1554 1555 1560 1556
rect 1423 1552 1441 1554
rect 1423 1551 1424 1552
rect 1418 1550 1424 1551
rect 1554 1551 1555 1555
rect 1559 1554 1560 1555
rect 1559 1552 1577 1554
rect 1559 1551 1560 1552
rect 1554 1550 1560 1551
rect 1394 1546 1400 1547
rect 862 1511 868 1512
rect 862 1510 863 1511
rect 695 1509 701 1510
rect 110 1505 116 1506
rect 110 1501 111 1505
rect 115 1501 116 1505
rect 695 1505 696 1509
rect 700 1508 701 1509
rect 714 1509 720 1510
rect 714 1508 715 1509
rect 700 1506 715 1508
rect 700 1505 701 1506
rect 695 1504 701 1505
rect 714 1505 715 1506
rect 719 1505 720 1509
rect 714 1504 720 1505
rect 831 1509 837 1510
rect 831 1505 832 1509
rect 836 1508 837 1509
rect 848 1508 863 1510
rect 836 1506 850 1508
rect 862 1507 863 1508
rect 867 1507 868 1511
rect 862 1506 868 1507
rect 967 1509 976 1510
rect 836 1505 837 1506
rect 831 1504 837 1505
rect 967 1505 968 1509
rect 975 1505 976 1509
rect 967 1504 976 1505
rect 1111 1509 1120 1510
rect 1111 1505 1112 1509
rect 1119 1505 1120 1509
rect 1111 1504 1120 1505
rect 1242 1509 1248 1510
rect 1242 1505 1243 1509
rect 1247 1508 1248 1509
rect 1255 1509 1261 1510
rect 1255 1508 1256 1509
rect 1247 1506 1256 1508
rect 1247 1505 1248 1506
rect 1242 1504 1248 1505
rect 1255 1505 1256 1506
rect 1260 1505 1261 1509
rect 1255 1504 1261 1505
rect 1399 1509 1405 1510
rect 1399 1505 1400 1509
rect 1404 1508 1405 1509
rect 1418 1509 1424 1510
rect 1418 1508 1419 1509
rect 1404 1506 1419 1508
rect 1404 1505 1405 1506
rect 1399 1504 1405 1505
rect 1418 1505 1419 1506
rect 1423 1505 1424 1509
rect 1418 1504 1424 1505
rect 1535 1509 1541 1510
rect 1535 1505 1536 1509
rect 1540 1508 1541 1509
rect 1554 1509 1560 1510
rect 1554 1508 1555 1509
rect 1540 1506 1555 1508
rect 1540 1505 1541 1506
rect 1535 1504 1541 1505
rect 1554 1505 1555 1506
rect 1559 1505 1560 1509
rect 1554 1504 1560 1505
rect 1666 1509 1677 1510
rect 1666 1505 1667 1509
rect 1671 1505 1672 1509
rect 1676 1505 1677 1509
rect 1666 1504 1677 1505
rect 1718 1505 1724 1506
rect 110 1500 116 1501
rect 598 1503 604 1504
rect 598 1499 599 1503
rect 603 1499 604 1503
rect 598 1498 604 1499
rect 734 1503 740 1504
rect 734 1499 735 1503
rect 739 1499 740 1503
rect 734 1498 740 1499
rect 870 1503 876 1504
rect 870 1499 871 1503
rect 875 1499 876 1503
rect 870 1498 876 1499
rect 1014 1503 1020 1504
rect 1014 1499 1015 1503
rect 1019 1499 1020 1503
rect 1014 1498 1020 1499
rect 1158 1503 1164 1504
rect 1158 1499 1159 1503
rect 1163 1499 1164 1503
rect 1158 1498 1164 1499
rect 1302 1503 1308 1504
rect 1302 1499 1303 1503
rect 1307 1499 1308 1503
rect 1302 1498 1308 1499
rect 1438 1503 1444 1504
rect 1438 1499 1439 1503
rect 1443 1499 1444 1503
rect 1438 1498 1444 1499
rect 1574 1503 1580 1504
rect 1574 1499 1575 1503
rect 1579 1499 1580 1503
rect 1718 1501 1719 1505
rect 1723 1501 1724 1505
rect 1718 1500 1724 1501
rect 1574 1498 1580 1499
rect 622 1488 628 1489
rect 110 1487 116 1488
rect 110 1483 111 1487
rect 115 1483 116 1487
rect 622 1484 623 1488
rect 627 1484 628 1488
rect 622 1483 628 1484
rect 758 1488 764 1489
rect 758 1484 759 1488
rect 763 1484 764 1488
rect 758 1483 764 1484
rect 894 1488 900 1489
rect 894 1484 895 1488
rect 899 1484 900 1488
rect 894 1483 900 1484
rect 1038 1488 1044 1489
rect 1038 1484 1039 1488
rect 1043 1484 1044 1488
rect 1038 1483 1044 1484
rect 1182 1488 1188 1489
rect 1182 1484 1183 1488
rect 1187 1484 1188 1488
rect 1182 1483 1188 1484
rect 1326 1488 1332 1489
rect 1326 1484 1327 1488
rect 1331 1484 1332 1488
rect 1326 1483 1332 1484
rect 1462 1488 1468 1489
rect 1462 1484 1463 1488
rect 1467 1484 1468 1488
rect 1462 1483 1468 1484
rect 1598 1488 1604 1489
rect 1598 1484 1599 1488
rect 1603 1484 1604 1488
rect 1598 1483 1604 1484
rect 1718 1487 1724 1488
rect 1718 1483 1719 1487
rect 1723 1483 1724 1487
rect 110 1482 116 1483
rect 1718 1482 1724 1483
rect 110 1425 116 1426
rect 1718 1425 1724 1426
rect 110 1421 111 1425
rect 115 1421 116 1425
rect 110 1420 116 1421
rect 598 1424 604 1425
rect 598 1420 599 1424
rect 603 1420 604 1424
rect 598 1419 604 1420
rect 734 1424 740 1425
rect 734 1420 735 1424
rect 739 1420 740 1424
rect 734 1419 740 1420
rect 878 1424 884 1425
rect 878 1420 879 1424
rect 883 1420 884 1424
rect 878 1419 884 1420
rect 1022 1424 1028 1425
rect 1022 1420 1023 1424
rect 1027 1420 1028 1424
rect 1022 1419 1028 1420
rect 1166 1424 1172 1425
rect 1166 1420 1167 1424
rect 1171 1420 1172 1424
rect 1166 1419 1172 1420
rect 1318 1424 1324 1425
rect 1318 1420 1319 1424
rect 1323 1420 1324 1424
rect 1318 1419 1324 1420
rect 1462 1424 1468 1425
rect 1462 1420 1463 1424
rect 1467 1420 1468 1424
rect 1462 1419 1468 1420
rect 1598 1424 1604 1425
rect 1598 1420 1599 1424
rect 1603 1420 1604 1424
rect 1718 1421 1719 1425
rect 1723 1421 1724 1425
rect 1718 1420 1724 1421
rect 1598 1419 1604 1420
rect 574 1409 580 1410
rect 110 1407 116 1408
rect 110 1403 111 1407
rect 115 1403 116 1407
rect 574 1405 575 1409
rect 579 1405 580 1409
rect 574 1404 580 1405
rect 710 1409 716 1410
rect 710 1405 711 1409
rect 715 1405 716 1409
rect 710 1404 716 1405
rect 854 1409 860 1410
rect 854 1405 855 1409
rect 859 1405 860 1409
rect 854 1404 860 1405
rect 998 1409 1004 1410
rect 998 1405 999 1409
rect 1003 1405 1004 1409
rect 998 1404 1004 1405
rect 1142 1409 1148 1410
rect 1142 1405 1143 1409
rect 1147 1405 1148 1409
rect 1142 1404 1148 1405
rect 1294 1409 1300 1410
rect 1294 1405 1295 1409
rect 1299 1405 1300 1409
rect 1294 1404 1300 1405
rect 1438 1409 1444 1410
rect 1438 1405 1439 1409
rect 1443 1405 1444 1409
rect 1438 1404 1444 1405
rect 1574 1409 1580 1410
rect 1574 1405 1575 1409
rect 1579 1405 1580 1409
rect 1574 1404 1580 1405
rect 1718 1407 1724 1408
rect 110 1402 116 1403
rect 671 1403 677 1404
rect 671 1399 672 1403
rect 676 1402 677 1403
rect 690 1403 696 1404
rect 690 1402 691 1403
rect 676 1400 691 1402
rect 676 1399 677 1400
rect 671 1398 677 1399
rect 690 1399 691 1400
rect 695 1399 696 1403
rect 690 1398 696 1399
rect 807 1403 813 1404
rect 807 1399 808 1403
rect 812 1402 813 1403
rect 831 1403 837 1404
rect 831 1402 832 1403
rect 812 1400 832 1402
rect 812 1399 813 1400
rect 807 1398 813 1399
rect 831 1399 832 1400
rect 836 1399 837 1403
rect 831 1398 837 1399
rect 951 1403 960 1404
rect 951 1399 952 1403
rect 959 1399 960 1403
rect 1095 1403 1101 1404
rect 1095 1402 1096 1403
rect 951 1398 960 1399
rect 964 1400 1096 1402
rect 666 1395 672 1396
rect 666 1391 667 1395
rect 671 1394 672 1395
rect 964 1394 966 1400
rect 1095 1399 1096 1400
rect 1100 1399 1101 1403
rect 1095 1398 1101 1399
rect 1118 1403 1124 1404
rect 1118 1399 1119 1403
rect 1123 1402 1124 1403
rect 1239 1403 1245 1404
rect 1239 1402 1240 1403
rect 1123 1400 1240 1402
rect 1123 1399 1124 1400
rect 1118 1398 1124 1399
rect 1239 1399 1240 1400
rect 1244 1399 1245 1403
rect 1239 1398 1245 1399
rect 1391 1403 1400 1404
rect 1391 1399 1392 1403
rect 1399 1399 1400 1403
rect 1391 1398 1400 1399
rect 1534 1403 1541 1404
rect 1534 1399 1535 1403
rect 1540 1399 1541 1403
rect 1534 1398 1541 1399
rect 1559 1403 1565 1404
rect 1559 1399 1560 1403
rect 1564 1402 1565 1403
rect 1671 1403 1677 1404
rect 1671 1402 1672 1403
rect 1564 1400 1672 1402
rect 1564 1399 1565 1400
rect 1559 1398 1565 1399
rect 1671 1399 1672 1400
rect 1676 1399 1677 1403
rect 1718 1403 1719 1407
rect 1723 1403 1724 1407
rect 1718 1402 1724 1403
rect 1671 1398 1677 1399
rect 671 1392 966 1394
rect 671 1391 672 1392
rect 666 1390 672 1391
rect 666 1359 672 1360
rect 666 1355 667 1359
rect 671 1355 672 1359
rect 666 1354 672 1355
rect 690 1359 696 1360
rect 690 1355 691 1359
rect 695 1358 696 1359
rect 831 1359 837 1360
rect 695 1356 713 1358
rect 695 1355 696 1356
rect 690 1354 696 1355
rect 831 1355 832 1359
rect 836 1358 837 1359
rect 1118 1359 1124 1360
rect 1118 1358 1119 1359
rect 836 1356 857 1358
rect 1093 1356 1119 1358
rect 836 1355 837 1356
rect 831 1354 837 1355
rect 1118 1355 1119 1356
rect 1123 1355 1124 1359
rect 1242 1359 1248 1360
rect 1242 1358 1243 1359
rect 1237 1356 1243 1358
rect 1118 1354 1124 1355
rect 1242 1355 1243 1356
rect 1247 1355 1248 1359
rect 1242 1354 1248 1355
rect 1350 1359 1356 1360
rect 1350 1355 1351 1359
rect 1355 1355 1356 1359
rect 1559 1359 1565 1360
rect 1559 1358 1560 1359
rect 1533 1356 1560 1358
rect 1350 1354 1356 1355
rect 1559 1355 1560 1356
rect 1564 1355 1565 1359
rect 1559 1354 1565 1355
rect 1666 1359 1672 1360
rect 1666 1355 1667 1359
rect 1671 1355 1672 1359
rect 1666 1354 1672 1355
rect 294 1335 300 1336
rect 294 1334 295 1335
rect 229 1332 295 1334
rect 294 1331 295 1332
rect 299 1331 300 1335
rect 510 1335 516 1336
rect 510 1334 511 1335
rect 397 1332 511 1334
rect 294 1330 300 1331
rect 510 1331 511 1332
rect 515 1331 516 1335
rect 730 1335 736 1336
rect 730 1334 731 1335
rect 613 1332 731 1334
rect 510 1330 516 1331
rect 730 1331 731 1332
rect 735 1331 736 1335
rect 943 1335 949 1336
rect 943 1334 944 1335
rect 845 1332 944 1334
rect 730 1330 736 1331
rect 943 1331 944 1332
rect 948 1331 949 1335
rect 943 1330 949 1331
rect 954 1335 960 1336
rect 954 1331 955 1335
rect 959 1334 960 1335
rect 1326 1335 1332 1336
rect 959 1332 1001 1334
rect 959 1331 960 1332
rect 954 1330 960 1331
rect 1326 1331 1327 1335
rect 1331 1331 1332 1335
rect 1326 1330 1332 1331
rect 1534 1335 1540 1336
rect 1534 1331 1535 1335
rect 1539 1331 1540 1335
rect 1534 1330 1540 1331
rect 294 1291 300 1292
rect 226 1289 237 1290
rect 110 1285 116 1286
rect 110 1281 111 1285
rect 115 1281 116 1285
rect 226 1285 227 1289
rect 231 1285 232 1289
rect 236 1285 237 1289
rect 294 1287 295 1291
rect 299 1290 300 1291
rect 510 1291 516 1292
rect 299 1288 382 1290
rect 399 1289 405 1290
rect 399 1288 400 1289
rect 299 1287 300 1288
rect 294 1286 300 1287
rect 380 1286 400 1288
rect 226 1284 237 1285
rect 399 1285 400 1286
rect 404 1285 405 1289
rect 510 1287 511 1291
rect 515 1290 516 1291
rect 730 1291 736 1292
rect 515 1288 598 1290
rect 615 1289 621 1290
rect 615 1288 616 1289
rect 515 1287 516 1288
rect 510 1286 516 1287
rect 596 1286 616 1288
rect 399 1284 405 1285
rect 615 1285 616 1286
rect 620 1285 621 1289
rect 730 1287 731 1291
rect 735 1290 736 1291
rect 943 1291 949 1292
rect 735 1288 830 1290
rect 847 1289 853 1290
rect 847 1288 848 1289
rect 735 1287 736 1288
rect 730 1286 736 1287
rect 828 1286 848 1288
rect 615 1284 621 1285
rect 847 1285 848 1286
rect 852 1285 853 1289
rect 943 1287 944 1291
rect 948 1290 949 1291
rect 948 1288 1078 1290
rect 1095 1289 1101 1290
rect 1095 1288 1096 1289
rect 948 1287 949 1288
rect 943 1286 949 1287
rect 1076 1286 1096 1288
rect 847 1284 853 1285
rect 1095 1285 1096 1286
rect 1100 1285 1101 1289
rect 1095 1284 1101 1285
rect 1350 1289 1357 1290
rect 1350 1285 1351 1289
rect 1356 1285 1357 1289
rect 1350 1284 1357 1285
rect 1614 1289 1621 1290
rect 1614 1285 1615 1289
rect 1620 1285 1621 1289
rect 1614 1284 1621 1285
rect 1718 1285 1724 1286
rect 110 1280 116 1281
rect 134 1283 140 1284
rect 134 1279 135 1283
rect 139 1279 140 1283
rect 134 1278 140 1279
rect 302 1283 308 1284
rect 302 1279 303 1283
rect 307 1279 308 1283
rect 302 1278 308 1279
rect 518 1283 524 1284
rect 518 1279 519 1283
rect 523 1279 524 1283
rect 518 1278 524 1279
rect 750 1283 756 1284
rect 750 1279 751 1283
rect 755 1279 756 1283
rect 750 1278 756 1279
rect 998 1283 1004 1284
rect 998 1279 999 1283
rect 1003 1279 1004 1283
rect 998 1278 1004 1279
rect 1254 1283 1260 1284
rect 1254 1279 1255 1283
rect 1259 1279 1260 1283
rect 1254 1278 1260 1279
rect 1518 1283 1524 1284
rect 1518 1279 1519 1283
rect 1523 1279 1524 1283
rect 1718 1281 1719 1285
rect 1723 1281 1724 1285
rect 1718 1280 1724 1281
rect 1518 1278 1524 1279
rect 158 1268 164 1269
rect 110 1267 116 1268
rect 110 1263 111 1267
rect 115 1263 116 1267
rect 158 1264 159 1268
rect 163 1264 164 1268
rect 158 1263 164 1264
rect 326 1268 332 1269
rect 326 1264 327 1268
rect 331 1264 332 1268
rect 326 1263 332 1264
rect 542 1268 548 1269
rect 542 1264 543 1268
rect 547 1264 548 1268
rect 542 1263 548 1264
rect 774 1268 780 1269
rect 774 1264 775 1268
rect 779 1264 780 1268
rect 774 1263 780 1264
rect 1022 1268 1028 1269
rect 1022 1264 1023 1268
rect 1027 1264 1028 1268
rect 1022 1263 1028 1264
rect 1278 1268 1284 1269
rect 1278 1264 1279 1268
rect 1283 1264 1284 1268
rect 1278 1263 1284 1264
rect 1542 1268 1548 1269
rect 1542 1264 1543 1268
rect 1547 1264 1548 1268
rect 1542 1263 1548 1264
rect 1718 1267 1724 1268
rect 1718 1263 1719 1267
rect 1723 1263 1724 1267
rect 110 1262 116 1263
rect 1718 1262 1724 1263
rect 110 1197 116 1198
rect 1718 1197 1724 1198
rect 110 1193 111 1197
rect 115 1193 116 1197
rect 110 1192 116 1193
rect 158 1196 164 1197
rect 158 1192 159 1196
rect 163 1192 164 1196
rect 158 1191 164 1192
rect 398 1196 404 1197
rect 398 1192 399 1196
rect 403 1192 404 1196
rect 398 1191 404 1192
rect 670 1196 676 1197
rect 670 1192 671 1196
rect 675 1192 676 1196
rect 670 1191 676 1192
rect 958 1196 964 1197
rect 958 1192 959 1196
rect 963 1192 964 1196
rect 958 1191 964 1192
rect 1254 1196 1260 1197
rect 1254 1192 1255 1196
rect 1259 1192 1260 1196
rect 1254 1191 1260 1192
rect 1550 1196 1556 1197
rect 1550 1192 1551 1196
rect 1555 1192 1556 1196
rect 1718 1193 1719 1197
rect 1723 1193 1724 1197
rect 1718 1192 1724 1193
rect 1550 1191 1556 1192
rect 134 1181 140 1182
rect 110 1179 116 1180
rect 110 1175 111 1179
rect 115 1175 116 1179
rect 134 1177 135 1181
rect 139 1177 140 1181
rect 134 1176 140 1177
rect 374 1181 380 1182
rect 374 1177 375 1181
rect 379 1177 380 1181
rect 374 1176 380 1177
rect 646 1181 652 1182
rect 646 1177 647 1181
rect 651 1177 652 1181
rect 646 1176 652 1177
rect 934 1181 940 1182
rect 934 1177 935 1181
rect 939 1177 940 1181
rect 934 1176 940 1177
rect 1230 1181 1236 1182
rect 1230 1177 1231 1181
rect 1235 1177 1236 1181
rect 1230 1176 1236 1177
rect 1526 1181 1532 1182
rect 1526 1177 1527 1181
rect 1531 1177 1532 1181
rect 1526 1176 1532 1177
rect 1718 1179 1724 1180
rect 110 1174 116 1175
rect 231 1175 240 1176
rect 231 1171 232 1175
rect 239 1171 240 1175
rect 231 1170 240 1171
rect 471 1175 480 1176
rect 471 1171 472 1175
rect 479 1171 480 1175
rect 471 1170 480 1171
rect 743 1175 749 1176
rect 743 1171 744 1175
rect 748 1174 749 1175
rect 802 1175 808 1176
rect 802 1174 803 1175
rect 748 1172 803 1174
rect 748 1171 749 1172
rect 743 1170 749 1171
rect 802 1171 803 1172
rect 807 1171 808 1175
rect 802 1170 808 1171
rect 918 1175 924 1176
rect 918 1171 919 1175
rect 923 1174 924 1175
rect 1031 1175 1037 1176
rect 1031 1174 1032 1175
rect 923 1172 1032 1174
rect 923 1171 924 1172
rect 918 1170 924 1171
rect 1031 1171 1032 1172
rect 1036 1171 1037 1175
rect 1031 1170 1037 1171
rect 1326 1175 1333 1176
rect 1326 1171 1327 1175
rect 1332 1171 1333 1175
rect 1326 1170 1333 1171
rect 1622 1175 1629 1176
rect 1622 1171 1623 1175
rect 1628 1171 1629 1175
rect 1718 1175 1719 1179
rect 1723 1175 1724 1179
rect 1718 1174 1724 1175
rect 1622 1170 1629 1171
rect 282 1155 288 1156
rect 282 1151 283 1155
rect 287 1154 288 1155
rect 918 1155 924 1156
rect 918 1154 919 1155
rect 287 1152 919 1154
rect 287 1151 288 1152
rect 282 1150 288 1151
rect 918 1151 919 1152
rect 923 1151 924 1155
rect 918 1150 924 1151
rect 226 1131 232 1132
rect 226 1127 227 1131
rect 231 1127 232 1131
rect 226 1126 232 1127
rect 234 1131 240 1132
rect 234 1127 235 1131
rect 239 1130 240 1131
rect 474 1131 480 1132
rect 239 1128 377 1130
rect 239 1127 240 1128
rect 234 1126 240 1127
rect 474 1127 475 1131
rect 479 1130 480 1131
rect 802 1131 808 1132
rect 479 1128 649 1130
rect 479 1127 480 1128
rect 474 1126 480 1127
rect 802 1127 803 1131
rect 807 1130 808 1131
rect 1410 1131 1416 1132
rect 1410 1130 1411 1131
rect 807 1128 937 1130
rect 1325 1128 1411 1130
rect 807 1127 808 1128
rect 802 1126 808 1127
rect 1410 1127 1411 1128
rect 1415 1127 1416 1131
rect 1410 1126 1416 1127
rect 1614 1131 1620 1132
rect 1614 1127 1615 1131
rect 1619 1127 1620 1131
rect 1614 1126 1620 1127
rect 282 1123 288 1124
rect 282 1119 283 1123
rect 287 1119 288 1123
rect 282 1118 288 1119
rect 290 1123 296 1124
rect 290 1119 291 1123
rect 295 1122 296 1123
rect 530 1123 536 1124
rect 295 1120 417 1122
rect 295 1119 296 1120
rect 290 1118 296 1119
rect 530 1119 531 1123
rect 535 1122 536 1123
rect 786 1123 792 1124
rect 535 1120 673 1122
rect 535 1119 536 1120
rect 530 1118 536 1119
rect 786 1119 787 1123
rect 791 1122 792 1123
rect 1066 1123 1072 1124
rect 791 1120 953 1122
rect 791 1119 792 1120
rect 786 1118 792 1119
rect 1066 1119 1067 1123
rect 1071 1122 1072 1123
rect 1622 1123 1628 1124
rect 1071 1120 1249 1122
rect 1071 1119 1072 1120
rect 1066 1118 1072 1119
rect 1622 1119 1623 1123
rect 1627 1119 1628 1123
rect 1622 1118 1628 1119
rect 287 1077 296 1078
rect 110 1073 116 1074
rect 110 1069 111 1073
rect 115 1069 116 1073
rect 287 1073 288 1077
rect 295 1073 296 1077
rect 287 1072 296 1073
rect 511 1077 517 1078
rect 511 1073 512 1077
rect 516 1076 517 1077
rect 530 1077 536 1078
rect 530 1076 531 1077
rect 516 1074 531 1076
rect 516 1073 517 1074
rect 511 1072 517 1073
rect 530 1073 531 1074
rect 535 1073 536 1077
rect 530 1072 536 1073
rect 767 1077 773 1078
rect 767 1073 768 1077
rect 772 1076 773 1077
rect 786 1077 792 1078
rect 786 1076 787 1077
rect 772 1074 787 1076
rect 772 1073 773 1074
rect 767 1072 773 1073
rect 786 1073 787 1074
rect 791 1073 792 1077
rect 786 1072 792 1073
rect 1047 1077 1053 1078
rect 1047 1073 1048 1077
rect 1052 1076 1053 1077
rect 1066 1077 1072 1078
rect 1066 1076 1067 1077
rect 1052 1074 1067 1076
rect 1052 1073 1053 1074
rect 1047 1072 1053 1073
rect 1066 1073 1067 1074
rect 1071 1073 1072 1077
rect 1066 1072 1072 1073
rect 1342 1077 1349 1078
rect 1342 1073 1343 1077
rect 1348 1073 1349 1077
rect 1342 1072 1349 1073
rect 1638 1077 1645 1078
rect 1638 1073 1639 1077
rect 1644 1073 1645 1077
rect 1638 1072 1645 1073
rect 1718 1073 1724 1074
rect 110 1068 116 1069
rect 190 1071 196 1072
rect 190 1067 191 1071
rect 195 1067 196 1071
rect 190 1066 196 1067
rect 414 1071 420 1072
rect 414 1067 415 1071
rect 419 1067 420 1071
rect 414 1066 420 1067
rect 670 1071 676 1072
rect 670 1067 671 1071
rect 675 1067 676 1071
rect 670 1066 676 1067
rect 950 1071 956 1072
rect 950 1067 951 1071
rect 955 1067 956 1071
rect 950 1066 956 1067
rect 1246 1071 1252 1072
rect 1246 1067 1247 1071
rect 1251 1067 1252 1071
rect 1246 1066 1252 1067
rect 1542 1071 1548 1072
rect 1542 1067 1543 1071
rect 1547 1067 1548 1071
rect 1718 1069 1719 1073
rect 1723 1069 1724 1073
rect 1718 1068 1724 1069
rect 1542 1066 1548 1067
rect 214 1056 220 1057
rect 110 1055 116 1056
rect 110 1051 111 1055
rect 115 1051 116 1055
rect 214 1052 215 1056
rect 219 1052 220 1056
rect 214 1051 220 1052
rect 438 1056 444 1057
rect 438 1052 439 1056
rect 443 1052 444 1056
rect 438 1051 444 1052
rect 694 1056 700 1057
rect 694 1052 695 1056
rect 699 1052 700 1056
rect 694 1051 700 1052
rect 974 1056 980 1057
rect 974 1052 975 1056
rect 979 1052 980 1056
rect 974 1051 980 1052
rect 1270 1056 1276 1057
rect 1270 1052 1271 1056
rect 1275 1052 1276 1056
rect 1270 1051 1276 1052
rect 1566 1056 1572 1057
rect 1566 1052 1567 1056
rect 1571 1052 1572 1056
rect 1566 1051 1572 1052
rect 1718 1055 1724 1056
rect 1718 1051 1719 1055
rect 1723 1051 1724 1055
rect 110 1050 116 1051
rect 1718 1050 1724 1051
rect 110 981 116 982
rect 1718 981 1724 982
rect 110 977 111 981
rect 115 977 116 981
rect 110 976 116 977
rect 510 980 516 981
rect 510 976 511 980
rect 515 976 516 980
rect 510 975 516 976
rect 662 980 668 981
rect 662 976 663 980
rect 667 976 668 980
rect 662 975 668 976
rect 830 980 836 981
rect 830 976 831 980
rect 835 976 836 980
rect 830 975 836 976
rect 1006 980 1012 981
rect 1006 976 1007 980
rect 1011 976 1012 980
rect 1006 975 1012 976
rect 1198 980 1204 981
rect 1198 976 1199 980
rect 1203 976 1204 980
rect 1198 975 1204 976
rect 1398 980 1404 981
rect 1398 976 1399 980
rect 1403 976 1404 980
rect 1398 975 1404 976
rect 1598 980 1604 981
rect 1598 976 1599 980
rect 1603 976 1604 980
rect 1718 977 1719 981
rect 1723 977 1724 981
rect 1718 976 1724 977
rect 1598 975 1604 976
rect 486 965 492 966
rect 110 963 116 964
rect 110 959 111 963
rect 115 959 116 963
rect 486 961 487 965
rect 491 961 492 965
rect 486 960 492 961
rect 638 965 644 966
rect 638 961 639 965
rect 643 961 644 965
rect 638 960 644 961
rect 806 965 812 966
rect 806 961 807 965
rect 811 961 812 965
rect 806 960 812 961
rect 982 965 988 966
rect 982 961 983 965
rect 987 961 988 965
rect 982 960 988 961
rect 1174 965 1180 966
rect 1174 961 1175 965
rect 1179 961 1180 965
rect 1174 960 1180 961
rect 1374 965 1380 966
rect 1374 961 1375 965
rect 1379 961 1380 965
rect 1374 960 1380 961
rect 1574 965 1580 966
rect 1574 961 1575 965
rect 1579 961 1580 965
rect 1574 960 1580 961
rect 1718 963 1724 964
rect 110 958 116 959
rect 583 959 592 960
rect 583 955 584 959
rect 591 955 592 959
rect 583 954 592 955
rect 735 959 744 960
rect 735 955 736 959
rect 743 955 744 959
rect 735 954 744 955
rect 903 959 909 960
rect 903 955 904 959
rect 908 958 909 959
rect 927 959 933 960
rect 927 958 928 959
rect 908 956 928 958
rect 908 955 909 956
rect 903 954 909 955
rect 927 955 928 956
rect 932 955 933 959
rect 927 954 933 955
rect 1079 959 1085 960
rect 1079 955 1080 959
rect 1084 958 1085 959
rect 1118 959 1124 960
rect 1118 958 1119 959
rect 1084 956 1119 958
rect 1084 955 1085 956
rect 1079 954 1085 955
rect 1118 955 1119 956
rect 1123 955 1124 959
rect 1118 954 1124 955
rect 1158 959 1164 960
rect 1158 955 1159 959
rect 1163 958 1164 959
rect 1271 959 1277 960
rect 1271 958 1272 959
rect 1163 956 1272 958
rect 1163 955 1164 956
rect 1158 954 1164 955
rect 1271 955 1272 956
rect 1276 955 1277 959
rect 1271 954 1277 955
rect 1410 959 1416 960
rect 1410 955 1411 959
rect 1415 958 1416 959
rect 1471 959 1477 960
rect 1471 958 1472 959
rect 1415 956 1472 958
rect 1415 955 1416 956
rect 1410 954 1416 955
rect 1471 955 1472 956
rect 1476 955 1477 959
rect 1471 954 1477 955
rect 1666 959 1677 960
rect 1666 955 1667 959
rect 1671 955 1672 959
rect 1676 955 1677 959
rect 1718 959 1719 963
rect 1723 959 1724 963
rect 1718 958 1724 959
rect 1666 954 1677 955
rect 578 951 584 952
rect 578 947 579 951
rect 583 950 584 951
rect 1342 951 1348 952
rect 1342 950 1343 951
rect 583 948 1343 950
rect 583 947 584 948
rect 578 946 584 947
rect 1342 947 1343 948
rect 1347 947 1348 951
rect 1342 946 1348 947
rect 578 915 584 916
rect 578 911 579 915
rect 583 911 584 915
rect 578 910 584 911
rect 586 915 592 916
rect 586 911 587 915
rect 591 914 592 915
rect 738 915 744 916
rect 591 912 641 914
rect 591 911 592 912
rect 586 910 592 911
rect 738 911 739 915
rect 743 914 744 915
rect 927 915 933 916
rect 743 912 809 914
rect 743 911 744 912
rect 738 910 744 911
rect 927 911 928 915
rect 932 914 933 915
rect 1118 915 1124 916
rect 932 912 985 914
rect 932 911 933 912
rect 927 910 933 911
rect 1118 911 1119 915
rect 1123 914 1124 915
rect 1638 915 1644 916
rect 1123 912 1177 914
rect 1123 911 1124 912
rect 1118 910 1124 911
rect 1456 910 1458 913
rect 1494 911 1500 912
rect 1494 910 1495 911
rect 1456 908 1495 910
rect 1494 907 1495 908
rect 1499 907 1500 911
rect 1638 911 1639 915
rect 1643 911 1644 915
rect 1638 910 1644 911
rect 1494 906 1500 907
rect 1158 903 1164 904
rect 1158 902 1159 903
rect 848 900 1159 902
rect 848 893 850 900
rect 1158 899 1159 900
rect 1163 899 1164 903
rect 1158 898 1164 899
rect 858 895 864 896
rect 858 891 859 895
rect 863 894 864 895
rect 1010 895 1016 896
rect 863 892 913 894
rect 863 891 864 892
rect 858 890 864 891
rect 1010 891 1011 895
rect 1015 894 1016 895
rect 1182 895 1188 896
rect 1015 892 1073 894
rect 1015 891 1016 892
rect 1010 890 1016 891
rect 1182 891 1183 895
rect 1187 894 1188 895
rect 1338 895 1344 896
rect 1187 892 1241 894
rect 1187 891 1188 892
rect 1182 890 1188 891
rect 1338 891 1339 895
rect 1343 894 1344 895
rect 1666 895 1672 896
rect 1343 892 1409 894
rect 1343 891 1344 892
rect 1338 890 1344 891
rect 1666 891 1667 895
rect 1671 891 1672 895
rect 1666 890 1672 891
rect 1338 851 1344 852
rect 1338 850 1339 851
rect 855 849 864 850
rect 110 845 116 846
rect 110 841 111 845
rect 115 841 116 845
rect 855 845 856 849
rect 863 845 864 849
rect 855 844 864 845
rect 1007 849 1016 850
rect 1007 845 1008 849
rect 1015 845 1016 849
rect 1007 844 1016 845
rect 1167 849 1173 850
rect 1167 845 1168 849
rect 1172 848 1173 849
rect 1182 849 1188 850
rect 1182 848 1183 849
rect 1172 846 1183 848
rect 1172 845 1173 846
rect 1167 844 1173 845
rect 1182 845 1183 846
rect 1187 845 1188 849
rect 1182 844 1188 845
rect 1335 849 1339 850
rect 1335 845 1336 849
rect 1343 847 1344 851
rect 1340 846 1344 847
rect 1378 851 1384 852
rect 1378 847 1379 851
rect 1383 850 1384 851
rect 1383 848 1486 850
rect 1503 849 1509 850
rect 1503 848 1504 849
rect 1383 847 1384 848
rect 1378 846 1384 847
rect 1484 846 1504 848
rect 1340 845 1341 846
rect 1335 844 1341 845
rect 1503 845 1504 846
rect 1508 845 1509 849
rect 1503 844 1509 845
rect 1666 849 1677 850
rect 1666 845 1667 849
rect 1671 845 1672 849
rect 1676 845 1677 849
rect 1666 844 1677 845
rect 1718 845 1724 846
rect 110 840 116 841
rect 758 843 764 844
rect 758 839 759 843
rect 763 839 764 843
rect 758 838 764 839
rect 910 843 916 844
rect 910 839 911 843
rect 915 839 916 843
rect 910 838 916 839
rect 1070 843 1076 844
rect 1070 839 1071 843
rect 1075 839 1076 843
rect 1070 838 1076 839
rect 1238 843 1244 844
rect 1238 839 1239 843
rect 1243 839 1244 843
rect 1238 838 1244 839
rect 1406 843 1412 844
rect 1406 839 1407 843
rect 1411 839 1412 843
rect 1406 838 1412 839
rect 1574 843 1580 844
rect 1574 839 1575 843
rect 1579 839 1580 843
rect 1718 841 1719 845
rect 1723 841 1724 845
rect 1718 840 1724 841
rect 1574 838 1580 839
rect 782 828 788 829
rect 110 827 116 828
rect 110 823 111 827
rect 115 823 116 827
rect 782 824 783 828
rect 787 824 788 828
rect 782 823 788 824
rect 934 828 940 829
rect 934 824 935 828
rect 939 824 940 828
rect 934 823 940 824
rect 1094 828 1100 829
rect 1094 824 1095 828
rect 1099 824 1100 828
rect 1094 823 1100 824
rect 1262 828 1268 829
rect 1262 824 1263 828
rect 1267 824 1268 828
rect 1262 823 1268 824
rect 1430 828 1436 829
rect 1430 824 1431 828
rect 1435 824 1436 828
rect 1430 823 1436 824
rect 1598 828 1604 829
rect 1598 824 1599 828
rect 1603 824 1604 828
rect 1598 823 1604 824
rect 1718 827 1724 828
rect 1718 823 1719 827
rect 1723 823 1724 827
rect 110 822 116 823
rect 1718 822 1724 823
rect 110 761 116 762
rect 1718 761 1724 762
rect 110 757 111 761
rect 115 757 116 761
rect 110 756 116 757
rect 694 760 700 761
rect 694 756 695 760
rect 699 756 700 760
rect 694 755 700 756
rect 830 760 836 761
rect 830 756 831 760
rect 835 756 836 760
rect 830 755 836 756
rect 974 760 980 761
rect 974 756 975 760
rect 979 756 980 760
rect 974 755 980 756
rect 1118 760 1124 761
rect 1118 756 1119 760
rect 1123 756 1124 760
rect 1118 755 1124 756
rect 1270 760 1276 761
rect 1270 756 1271 760
rect 1275 756 1276 760
rect 1270 755 1276 756
rect 1430 760 1436 761
rect 1430 756 1431 760
rect 1435 756 1436 760
rect 1430 755 1436 756
rect 1598 760 1604 761
rect 1598 756 1599 760
rect 1603 756 1604 760
rect 1718 757 1719 761
rect 1723 757 1724 761
rect 1718 756 1724 757
rect 1598 755 1604 756
rect 670 745 676 746
rect 110 743 116 744
rect 110 739 111 743
rect 115 739 116 743
rect 670 741 671 745
rect 675 741 676 745
rect 670 740 676 741
rect 806 745 812 746
rect 806 741 807 745
rect 811 741 812 745
rect 806 740 812 741
rect 950 745 956 746
rect 950 741 951 745
rect 955 741 956 745
rect 950 740 956 741
rect 1094 745 1100 746
rect 1094 741 1095 745
rect 1099 741 1100 745
rect 1094 740 1100 741
rect 1246 745 1252 746
rect 1246 741 1247 745
rect 1251 741 1252 745
rect 1246 740 1252 741
rect 1406 745 1412 746
rect 1406 741 1407 745
rect 1411 741 1412 745
rect 1406 740 1412 741
rect 1574 745 1580 746
rect 1574 741 1575 745
rect 1579 741 1580 745
rect 1574 740 1580 741
rect 1718 743 1724 744
rect 110 738 116 739
rect 767 739 773 740
rect 767 735 768 739
rect 772 738 773 739
rect 790 739 796 740
rect 790 738 791 739
rect 772 736 791 738
rect 772 735 773 736
rect 767 734 773 735
rect 790 735 791 736
rect 795 735 796 739
rect 790 734 796 735
rect 903 739 909 740
rect 903 735 904 739
rect 908 738 909 739
rect 927 739 933 740
rect 927 738 928 739
rect 908 736 928 738
rect 908 735 909 736
rect 903 734 909 735
rect 927 735 928 736
rect 932 735 933 739
rect 927 734 933 735
rect 1047 739 1056 740
rect 1047 735 1048 739
rect 1055 735 1056 739
rect 1191 739 1197 740
rect 1191 738 1192 739
rect 1047 734 1056 735
rect 1060 736 1192 738
rect 762 731 768 732
rect 762 727 763 731
rect 767 730 768 731
rect 1060 730 1062 736
rect 1191 735 1192 736
rect 1196 735 1197 739
rect 1191 734 1197 735
rect 1218 739 1224 740
rect 1218 735 1219 739
rect 1223 738 1224 739
rect 1343 739 1349 740
rect 1343 738 1344 739
rect 1223 736 1344 738
rect 1223 735 1224 736
rect 1218 734 1224 735
rect 1343 735 1344 736
rect 1348 735 1349 739
rect 1343 734 1349 735
rect 1494 739 1500 740
rect 1494 735 1495 739
rect 1499 738 1500 739
rect 1503 739 1509 740
rect 1503 738 1504 739
rect 1499 736 1504 738
rect 1499 735 1500 736
rect 1494 734 1500 735
rect 1503 735 1504 736
rect 1508 735 1509 739
rect 1503 734 1509 735
rect 1650 739 1656 740
rect 1650 735 1651 739
rect 1655 738 1656 739
rect 1671 739 1677 740
rect 1671 738 1672 739
rect 1655 736 1672 738
rect 1655 735 1656 736
rect 1650 734 1656 735
rect 1671 735 1672 736
rect 1676 735 1677 739
rect 1718 739 1719 743
rect 1723 739 1724 743
rect 1718 738 1724 739
rect 1671 734 1677 735
rect 767 728 1062 730
rect 767 727 768 728
rect 762 726 768 727
rect 762 695 768 696
rect 762 691 763 695
rect 767 691 768 695
rect 762 690 768 691
rect 790 695 796 696
rect 790 691 791 695
rect 795 694 796 695
rect 927 695 933 696
rect 795 692 809 694
rect 795 691 796 692
rect 790 690 796 691
rect 927 691 928 695
rect 932 694 933 695
rect 1218 695 1224 696
rect 1218 694 1219 695
rect 932 692 953 694
rect 1189 692 1219 694
rect 932 691 933 692
rect 927 690 933 691
rect 1218 691 1219 692
rect 1223 691 1224 695
rect 1378 695 1384 696
rect 1378 694 1379 695
rect 1341 692 1379 694
rect 1218 690 1224 691
rect 1378 691 1379 692
rect 1383 691 1384 695
rect 1378 690 1384 691
rect 1414 695 1420 696
rect 1414 691 1415 695
rect 1419 691 1420 695
rect 1414 690 1420 691
rect 1666 695 1672 696
rect 1666 691 1667 695
rect 1671 691 1672 695
rect 1666 690 1672 691
rect 423 663 429 664
rect 423 662 424 663
rect 341 660 424 662
rect 423 659 424 660
rect 428 659 429 663
rect 622 663 628 664
rect 622 662 623 663
rect 525 660 623 662
rect 423 658 429 659
rect 622 659 623 660
rect 627 659 628 663
rect 838 663 844 664
rect 838 662 839 663
rect 725 660 839 662
rect 622 658 628 659
rect 838 659 839 660
rect 843 659 844 663
rect 1042 663 1048 664
rect 1042 662 1043 663
rect 941 660 1043 662
rect 838 658 844 659
rect 1042 659 1043 660
rect 1047 659 1048 663
rect 1042 658 1048 659
rect 1050 663 1056 664
rect 1050 659 1051 663
rect 1055 662 1056 663
rect 1434 663 1440 664
rect 1434 662 1435 663
rect 1055 660 1081 662
rect 1413 660 1435 662
rect 1055 659 1056 660
rect 1050 658 1056 659
rect 1434 659 1435 660
rect 1439 659 1440 663
rect 1434 658 1440 659
rect 1650 663 1656 664
rect 1650 659 1651 663
rect 1655 659 1656 663
rect 1650 658 1656 659
rect 258 619 264 620
rect 258 615 259 619
rect 263 618 264 619
rect 423 619 429 620
rect 263 616 326 618
rect 343 617 349 618
rect 343 616 344 617
rect 263 615 264 616
rect 258 614 264 615
rect 324 614 344 616
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 343 613 344 614
rect 348 613 349 617
rect 423 615 424 619
rect 428 618 429 619
rect 622 619 628 620
rect 428 616 510 618
rect 527 617 533 618
rect 527 616 528 617
rect 428 615 429 616
rect 423 614 429 615
rect 508 614 528 616
rect 343 612 349 613
rect 527 613 528 614
rect 532 613 533 617
rect 622 615 623 619
rect 627 618 628 619
rect 838 619 844 620
rect 627 616 710 618
rect 727 617 733 618
rect 727 616 728 617
rect 627 615 628 616
rect 622 614 628 615
rect 708 614 728 616
rect 527 612 533 613
rect 727 613 728 614
rect 732 613 733 617
rect 838 615 839 619
rect 843 618 844 619
rect 1042 619 1048 620
rect 843 616 926 618
rect 943 617 949 618
rect 943 616 944 617
rect 843 615 844 616
rect 838 614 844 615
rect 924 614 944 616
rect 727 612 733 613
rect 943 613 944 614
rect 948 613 949 617
rect 1042 615 1043 619
rect 1047 618 1048 619
rect 1047 616 1158 618
rect 1175 617 1181 618
rect 1175 616 1176 617
rect 1047 615 1048 616
rect 1042 614 1048 615
rect 1156 614 1176 616
rect 943 612 949 613
rect 1175 613 1176 614
rect 1180 613 1181 617
rect 1175 612 1181 613
rect 1414 617 1421 618
rect 1414 613 1415 617
rect 1420 613 1421 617
rect 1414 612 1421 613
rect 1654 617 1661 618
rect 1654 613 1655 617
rect 1660 613 1661 617
rect 1654 612 1661 613
rect 1718 613 1724 614
rect 110 608 116 609
rect 246 611 252 612
rect 246 607 247 611
rect 251 607 252 611
rect 246 606 252 607
rect 430 611 436 612
rect 430 607 431 611
rect 435 607 436 611
rect 430 606 436 607
rect 630 611 636 612
rect 630 607 631 611
rect 635 607 636 611
rect 630 606 636 607
rect 846 611 852 612
rect 846 607 847 611
rect 851 607 852 611
rect 846 606 852 607
rect 1078 611 1084 612
rect 1078 607 1079 611
rect 1083 607 1084 611
rect 1078 606 1084 607
rect 1318 611 1324 612
rect 1318 607 1319 611
rect 1323 607 1324 611
rect 1318 606 1324 607
rect 1558 611 1564 612
rect 1558 607 1559 611
rect 1563 607 1564 611
rect 1718 609 1719 613
rect 1723 609 1724 613
rect 1718 608 1724 609
rect 1558 606 1564 607
rect 270 596 276 597
rect 110 595 116 596
rect 110 591 111 595
rect 115 591 116 595
rect 270 592 271 596
rect 275 592 276 596
rect 270 591 276 592
rect 454 596 460 597
rect 454 592 455 596
rect 459 592 460 596
rect 454 591 460 592
rect 654 596 660 597
rect 654 592 655 596
rect 659 592 660 596
rect 654 591 660 592
rect 870 596 876 597
rect 870 592 871 596
rect 875 592 876 596
rect 870 591 876 592
rect 1102 596 1108 597
rect 1102 592 1103 596
rect 1107 592 1108 596
rect 1102 591 1108 592
rect 1342 596 1348 597
rect 1342 592 1343 596
rect 1347 592 1348 596
rect 1342 591 1348 592
rect 1582 596 1588 597
rect 1582 592 1583 596
rect 1587 592 1588 596
rect 1582 591 1588 592
rect 1718 595 1724 596
rect 1718 591 1719 595
rect 1723 591 1724 595
rect 110 590 116 591
rect 1718 590 1724 591
rect 110 521 116 522
rect 1718 521 1724 522
rect 110 517 111 521
rect 115 517 116 521
rect 110 516 116 517
rect 158 520 164 521
rect 158 516 159 520
rect 163 516 164 520
rect 158 515 164 516
rect 342 520 348 521
rect 342 516 343 520
rect 347 516 348 520
rect 342 515 348 516
rect 574 520 580 521
rect 574 516 575 520
rect 579 516 580 520
rect 574 515 580 516
rect 830 520 836 521
rect 830 516 831 520
rect 835 516 836 520
rect 830 515 836 516
rect 1094 520 1100 521
rect 1094 516 1095 520
rect 1099 516 1100 520
rect 1094 515 1100 516
rect 1366 520 1372 521
rect 1366 516 1367 520
rect 1371 516 1372 520
rect 1718 517 1719 521
rect 1723 517 1724 521
rect 1718 516 1724 517
rect 1366 515 1372 516
rect 134 505 140 506
rect 110 503 116 504
rect 110 499 111 503
rect 115 499 116 503
rect 134 501 135 505
rect 139 501 140 505
rect 134 500 140 501
rect 318 505 324 506
rect 318 501 319 505
rect 323 501 324 505
rect 318 500 324 501
rect 550 505 556 506
rect 550 501 551 505
rect 555 501 556 505
rect 550 500 556 501
rect 806 505 812 506
rect 806 501 807 505
rect 811 501 812 505
rect 806 500 812 501
rect 1070 505 1076 506
rect 1070 501 1071 505
rect 1075 501 1076 505
rect 1070 500 1076 501
rect 1342 505 1348 506
rect 1342 501 1343 505
rect 1347 501 1348 505
rect 1342 500 1348 501
rect 1718 503 1724 504
rect 110 498 116 499
rect 231 499 237 500
rect 231 495 232 499
rect 236 498 237 499
rect 263 499 269 500
rect 263 498 264 499
rect 236 496 264 498
rect 236 495 237 496
rect 231 494 237 495
rect 263 495 264 496
rect 268 495 269 499
rect 263 494 269 495
rect 415 499 424 500
rect 415 495 416 499
rect 423 495 424 499
rect 415 494 424 495
rect 647 499 656 500
rect 647 495 648 499
rect 655 495 656 499
rect 647 494 656 495
rect 903 499 909 500
rect 903 495 904 499
rect 908 498 909 499
rect 943 499 949 500
rect 943 498 944 499
rect 908 496 944 498
rect 908 495 909 496
rect 903 494 909 495
rect 943 495 944 496
rect 948 495 949 499
rect 1167 499 1173 500
rect 1167 498 1168 499
rect 943 494 949 495
rect 952 496 1168 498
rect 290 491 296 492
rect 290 487 291 491
rect 295 490 296 491
rect 952 490 954 496
rect 1167 495 1168 496
rect 1172 495 1173 499
rect 1167 494 1173 495
rect 1434 499 1445 500
rect 1434 495 1435 499
rect 1439 495 1440 499
rect 1444 495 1445 499
rect 1718 499 1719 503
rect 1723 499 1724 503
rect 1718 498 1724 499
rect 1434 494 1445 495
rect 295 488 954 490
rect 295 487 296 488
rect 290 486 296 487
rect 254 455 260 456
rect 254 454 255 455
rect 229 452 255 454
rect 254 451 255 452
rect 259 451 260 455
rect 254 450 260 451
rect 263 455 269 456
rect 263 451 264 455
rect 268 454 269 455
rect 418 455 424 456
rect 268 452 321 454
rect 268 451 269 452
rect 263 450 269 451
rect 418 451 419 455
rect 423 454 424 455
rect 650 455 656 456
rect 423 452 553 454
rect 423 451 424 452
rect 418 450 424 451
rect 650 451 651 455
rect 655 454 656 455
rect 943 455 949 456
rect 655 452 809 454
rect 655 451 656 452
rect 650 450 656 451
rect 943 451 944 455
rect 948 454 949 455
rect 1422 455 1428 456
rect 948 452 1073 454
rect 948 451 949 452
rect 943 450 949 451
rect 1422 451 1423 455
rect 1427 451 1428 455
rect 1422 450 1428 451
rect 290 435 296 436
rect 290 431 291 435
rect 295 431 296 435
rect 290 430 296 431
rect 298 435 304 436
rect 298 431 299 435
rect 303 434 304 435
rect 530 435 536 436
rect 303 432 417 434
rect 303 431 304 432
rect 298 430 304 431
rect 530 431 531 435
rect 535 434 536 435
rect 730 435 736 436
rect 535 432 633 434
rect 535 431 536 432
rect 530 430 536 431
rect 730 431 731 435
rect 735 434 736 435
rect 1174 435 1180 436
rect 735 432 857 434
rect 735 431 736 432
rect 730 430 736 431
rect 1174 431 1175 435
rect 1179 431 1180 435
rect 1174 430 1180 431
rect 1186 435 1192 436
rect 1186 431 1187 435
rect 1191 434 1192 435
rect 1654 435 1660 436
rect 1191 432 1329 434
rect 1191 431 1192 432
rect 1186 430 1192 431
rect 1654 431 1655 435
rect 1659 431 1660 435
rect 1654 430 1660 431
rect 295 389 304 390
rect 110 385 116 386
rect 110 381 111 385
rect 115 381 116 385
rect 295 385 296 389
rect 303 385 304 389
rect 295 384 304 385
rect 511 389 517 390
rect 511 385 512 389
rect 516 388 517 389
rect 530 389 536 390
rect 530 388 531 389
rect 516 386 531 388
rect 516 385 517 386
rect 511 384 517 385
rect 530 385 531 386
rect 535 385 536 389
rect 530 384 536 385
rect 727 389 736 390
rect 727 385 728 389
rect 735 385 736 389
rect 727 384 736 385
rect 950 389 957 390
rect 950 385 951 389
rect 956 385 957 389
rect 950 384 957 385
rect 1183 389 1192 390
rect 1183 385 1184 389
rect 1191 385 1192 389
rect 1183 384 1192 385
rect 1422 389 1429 390
rect 1422 385 1423 389
rect 1428 385 1429 389
rect 1422 384 1429 385
rect 1671 389 1680 390
rect 1671 385 1672 389
rect 1679 385 1680 389
rect 1671 384 1680 385
rect 1718 385 1724 386
rect 110 380 116 381
rect 198 383 204 384
rect 198 379 199 383
rect 203 379 204 383
rect 198 378 204 379
rect 414 383 420 384
rect 414 379 415 383
rect 419 379 420 383
rect 414 378 420 379
rect 630 383 636 384
rect 630 379 631 383
rect 635 379 636 383
rect 630 378 636 379
rect 854 383 860 384
rect 854 379 855 383
rect 859 379 860 383
rect 854 378 860 379
rect 1086 383 1092 384
rect 1086 379 1087 383
rect 1091 379 1092 383
rect 1086 378 1092 379
rect 1326 383 1332 384
rect 1326 379 1327 383
rect 1331 379 1332 383
rect 1326 378 1332 379
rect 1574 383 1580 384
rect 1574 379 1575 383
rect 1579 379 1580 383
rect 1718 381 1719 385
rect 1723 381 1724 385
rect 1718 380 1724 381
rect 1574 378 1580 379
rect 222 368 228 369
rect 110 367 116 368
rect 110 363 111 367
rect 115 363 116 367
rect 222 364 223 368
rect 227 364 228 368
rect 222 363 228 364
rect 438 368 444 369
rect 438 364 439 368
rect 443 364 444 368
rect 438 363 444 364
rect 654 368 660 369
rect 654 364 655 368
rect 659 364 660 368
rect 654 363 660 364
rect 878 368 884 369
rect 878 364 879 368
rect 883 364 884 368
rect 878 363 884 364
rect 1110 368 1116 369
rect 1110 364 1111 368
rect 1115 364 1116 368
rect 1110 363 1116 364
rect 1350 368 1356 369
rect 1350 364 1351 368
rect 1355 364 1356 368
rect 1350 363 1356 364
rect 1598 368 1604 369
rect 1598 364 1599 368
rect 1603 364 1604 368
rect 1598 363 1604 364
rect 1718 367 1724 368
rect 1718 363 1719 367
rect 1723 363 1724 367
rect 110 362 116 363
rect 1718 362 1724 363
rect 110 305 116 306
rect 1718 305 1724 306
rect 110 301 111 305
rect 115 301 116 305
rect 110 300 116 301
rect 558 304 564 305
rect 558 300 559 304
rect 563 300 564 304
rect 558 299 564 300
rect 758 304 764 305
rect 758 300 759 304
rect 763 300 764 304
rect 758 299 764 300
rect 966 304 972 305
rect 966 300 967 304
rect 971 300 972 304
rect 966 299 972 300
rect 1182 304 1188 305
rect 1182 300 1183 304
rect 1187 300 1188 304
rect 1182 299 1188 300
rect 1398 304 1404 305
rect 1398 300 1399 304
rect 1403 300 1404 304
rect 1398 299 1404 300
rect 1598 304 1604 305
rect 1598 300 1599 304
rect 1603 300 1604 304
rect 1718 301 1719 305
rect 1723 301 1724 305
rect 1718 300 1724 301
rect 1598 299 1604 300
rect 534 289 540 290
rect 110 287 116 288
rect 110 283 111 287
rect 115 283 116 287
rect 534 285 535 289
rect 539 285 540 289
rect 534 284 540 285
rect 734 289 740 290
rect 734 285 735 289
rect 739 285 740 289
rect 734 284 740 285
rect 942 289 948 290
rect 942 285 943 289
rect 947 285 948 289
rect 942 284 948 285
rect 1158 289 1164 290
rect 1158 285 1159 289
rect 1163 285 1164 289
rect 1158 284 1164 285
rect 1374 289 1380 290
rect 1374 285 1375 289
rect 1379 285 1380 289
rect 1374 284 1380 285
rect 1574 289 1580 290
rect 1574 285 1575 289
rect 1579 285 1580 289
rect 1574 284 1580 285
rect 1718 287 1724 288
rect 110 282 116 283
rect 578 283 584 284
rect 578 279 579 283
rect 583 282 584 283
rect 631 283 637 284
rect 631 282 632 283
rect 583 280 632 282
rect 583 279 584 280
rect 578 278 584 279
rect 631 279 632 280
rect 636 279 637 283
rect 631 278 637 279
rect 654 283 660 284
rect 654 279 655 283
rect 659 282 660 283
rect 831 283 837 284
rect 831 282 832 283
rect 659 280 832 282
rect 659 279 660 280
rect 654 278 660 279
rect 831 279 832 280
rect 836 279 837 283
rect 831 278 837 279
rect 886 283 892 284
rect 886 279 887 283
rect 891 282 892 283
rect 1039 283 1045 284
rect 1039 282 1040 283
rect 891 280 1040 282
rect 891 279 892 280
rect 886 278 892 279
rect 1039 279 1040 280
rect 1044 279 1045 283
rect 1039 278 1045 279
rect 1174 283 1180 284
rect 1174 279 1175 283
rect 1179 282 1180 283
rect 1255 283 1261 284
rect 1255 282 1256 283
rect 1179 280 1256 282
rect 1179 279 1180 280
rect 1174 278 1180 279
rect 1255 279 1256 280
rect 1260 279 1261 283
rect 1255 278 1261 279
rect 1314 283 1320 284
rect 1314 279 1315 283
rect 1319 282 1320 283
rect 1471 283 1477 284
rect 1471 282 1472 283
rect 1319 280 1472 282
rect 1319 279 1320 280
rect 1314 278 1320 279
rect 1471 279 1472 280
rect 1476 279 1477 283
rect 1471 278 1477 279
rect 1666 283 1677 284
rect 1666 279 1667 283
rect 1671 279 1672 283
rect 1676 279 1677 283
rect 1718 283 1719 287
rect 1723 283 1724 287
rect 1718 282 1724 283
rect 1666 278 1677 279
rect 654 239 660 240
rect 654 238 655 239
rect 629 236 655 238
rect 654 235 655 236
rect 659 235 660 239
rect 886 239 892 240
rect 886 238 887 239
rect 829 236 887 238
rect 654 234 660 235
rect 886 235 887 236
rect 891 235 892 239
rect 886 234 892 235
rect 950 239 956 240
rect 950 235 951 239
rect 955 235 956 239
rect 1314 239 1320 240
rect 1314 238 1315 239
rect 1253 236 1315 238
rect 950 234 956 235
rect 1314 235 1315 236
rect 1319 235 1320 239
rect 1314 234 1320 235
rect 1398 239 1404 240
rect 1398 235 1399 239
rect 1403 235 1404 239
rect 1674 239 1680 240
rect 1674 238 1675 239
rect 1669 236 1675 238
rect 1398 234 1404 235
rect 1674 235 1675 236
rect 1679 235 1680 239
rect 1674 234 1680 235
rect 578 219 584 220
rect 578 215 579 219
rect 583 215 584 219
rect 578 214 584 215
rect 586 219 592 220
rect 586 215 587 219
rect 591 218 592 219
rect 722 219 728 220
rect 591 216 625 218
rect 591 215 592 216
rect 586 214 592 215
rect 722 215 723 219
rect 727 218 728 219
rect 874 219 880 220
rect 727 216 761 218
rect 727 215 728 216
rect 722 214 728 215
rect 874 215 875 219
rect 879 218 880 219
rect 1010 219 1016 220
rect 879 216 897 218
rect 879 215 880 216
rect 874 214 880 215
rect 1010 215 1011 219
rect 1015 218 1016 219
rect 1130 219 1136 220
rect 1015 216 1033 218
rect 1015 215 1016 216
rect 1010 214 1016 215
rect 1130 215 1131 219
rect 1135 218 1136 219
rect 1282 219 1288 220
rect 1135 216 1169 218
rect 1135 215 1136 216
rect 1130 214 1136 215
rect 1282 215 1283 219
rect 1287 218 1288 219
rect 1666 219 1672 220
rect 1287 216 1305 218
rect 1287 215 1288 216
rect 1282 214 1288 215
rect 1530 215 1536 216
rect 1530 211 1531 215
rect 1535 211 1536 215
rect 1666 215 1667 219
rect 1671 215 1672 219
rect 1666 214 1672 215
rect 1530 210 1536 211
rect 1530 175 1536 176
rect 583 173 592 174
rect 110 169 116 170
rect 110 165 111 169
rect 115 165 116 169
rect 583 169 584 173
rect 591 169 592 173
rect 583 168 592 169
rect 719 173 728 174
rect 719 169 720 173
rect 727 169 728 173
rect 719 168 728 169
rect 855 173 861 174
rect 855 169 856 173
rect 860 172 861 173
rect 874 173 880 174
rect 874 172 875 173
rect 860 170 875 172
rect 860 169 861 170
rect 855 168 861 169
rect 874 169 875 170
rect 879 169 880 173
rect 874 168 880 169
rect 991 173 997 174
rect 991 169 992 173
rect 996 172 997 173
rect 1010 173 1016 174
rect 1010 172 1011 173
rect 996 170 1011 172
rect 996 169 997 170
rect 991 168 997 169
rect 1010 169 1011 170
rect 1015 169 1016 173
rect 1010 168 1016 169
rect 1127 173 1136 174
rect 1127 169 1128 173
rect 1135 169 1136 173
rect 1127 168 1136 169
rect 1263 173 1269 174
rect 1263 169 1264 173
rect 1268 172 1269 173
rect 1282 173 1288 174
rect 1282 172 1283 173
rect 1268 170 1283 172
rect 1268 169 1269 170
rect 1263 168 1269 169
rect 1282 169 1283 170
rect 1287 169 1288 173
rect 1282 168 1288 169
rect 1398 173 1405 174
rect 1398 169 1399 173
rect 1404 169 1405 173
rect 1530 171 1531 175
rect 1535 174 1536 175
rect 1535 172 1654 174
rect 1671 173 1677 174
rect 1671 172 1672 173
rect 1535 171 1536 172
rect 1530 170 1536 171
rect 1652 170 1672 172
rect 1398 168 1405 169
rect 1671 169 1672 170
rect 1676 169 1677 173
rect 1671 168 1677 169
rect 1718 169 1724 170
rect 110 164 116 165
rect 486 167 492 168
rect 486 163 487 167
rect 491 163 492 167
rect 486 162 492 163
rect 622 167 628 168
rect 622 163 623 167
rect 627 163 628 167
rect 622 162 628 163
rect 758 167 764 168
rect 758 163 759 167
rect 763 163 764 167
rect 758 162 764 163
rect 894 167 900 168
rect 894 163 895 167
rect 899 163 900 167
rect 894 162 900 163
rect 1030 167 1036 168
rect 1030 163 1031 167
rect 1035 163 1036 167
rect 1030 162 1036 163
rect 1166 167 1172 168
rect 1166 163 1167 167
rect 1171 163 1172 167
rect 1166 162 1172 163
rect 1302 167 1308 168
rect 1302 163 1303 167
rect 1307 163 1308 167
rect 1302 162 1308 163
rect 1438 167 1444 168
rect 1438 163 1439 167
rect 1443 163 1444 167
rect 1438 162 1444 163
rect 1574 167 1580 168
rect 1574 163 1575 167
rect 1579 163 1580 167
rect 1718 165 1719 169
rect 1723 165 1724 169
rect 1718 164 1724 165
rect 1574 162 1580 163
rect 510 152 516 153
rect 110 151 116 152
rect 110 147 111 151
rect 115 147 116 151
rect 510 148 511 152
rect 515 148 516 152
rect 510 147 516 148
rect 646 152 652 153
rect 646 148 647 152
rect 651 148 652 152
rect 646 147 652 148
rect 782 152 788 153
rect 782 148 783 152
rect 787 148 788 152
rect 782 147 788 148
rect 918 152 924 153
rect 918 148 919 152
rect 923 148 924 152
rect 918 147 924 148
rect 1054 152 1060 153
rect 1054 148 1055 152
rect 1059 148 1060 152
rect 1054 147 1060 148
rect 1190 152 1196 153
rect 1190 148 1191 152
rect 1195 148 1196 152
rect 1190 147 1196 148
rect 1326 152 1332 153
rect 1326 148 1327 152
rect 1331 148 1332 152
rect 1326 147 1332 148
rect 1462 152 1468 153
rect 1462 148 1463 152
rect 1467 148 1468 152
rect 1462 147 1468 148
rect 1598 152 1604 153
rect 1598 148 1599 152
rect 1603 148 1604 152
rect 1598 147 1604 148
rect 1718 151 1724 152
rect 1718 147 1719 151
rect 1723 147 1724 151
rect 110 146 116 147
rect 1718 146 1724 147
<< m3c >>
rect 251 1775 255 1779
rect 387 1775 391 1779
rect 523 1775 527 1779
rect 659 1775 663 1779
rect 111 1725 115 1729
rect 251 1729 255 1733
rect 387 1729 391 1733
rect 523 1729 527 1733
rect 659 1729 663 1733
rect 775 1729 776 1733
rect 776 1729 779 1733
rect 135 1723 139 1727
rect 271 1723 275 1727
rect 407 1723 411 1727
rect 543 1723 547 1727
rect 679 1723 683 1727
rect 1719 1725 1723 1729
rect 111 1707 115 1711
rect 159 1708 163 1712
rect 295 1708 299 1712
rect 431 1708 435 1712
rect 567 1708 571 1712
rect 703 1708 707 1712
rect 1719 1707 1723 1711
rect 307 1671 311 1675
rect 775 1671 779 1675
rect 111 1641 115 1645
rect 239 1640 243 1644
rect 375 1640 379 1644
rect 511 1640 515 1644
rect 647 1640 651 1644
rect 783 1640 787 1644
rect 1719 1641 1723 1645
rect 111 1623 115 1627
rect 215 1625 219 1629
rect 351 1625 355 1629
rect 487 1625 491 1629
rect 623 1625 627 1629
rect 759 1625 763 1629
rect 331 1619 335 1623
rect 467 1619 471 1623
rect 587 1615 591 1619
rect 739 1619 743 1623
rect 691 1611 695 1615
rect 1719 1623 1723 1627
rect 307 1575 311 1579
rect 331 1575 335 1579
rect 467 1575 471 1579
rect 587 1575 591 1579
rect 739 1575 743 1579
rect 691 1551 695 1555
rect 715 1551 719 1555
rect 863 1551 867 1555
rect 971 1551 975 1555
rect 1115 1551 1119 1555
rect 1395 1547 1399 1551
rect 1419 1551 1423 1555
rect 1555 1551 1559 1555
rect 111 1501 115 1505
rect 715 1505 719 1509
rect 863 1507 867 1511
rect 971 1505 972 1509
rect 972 1505 975 1509
rect 1115 1505 1116 1509
rect 1116 1505 1119 1509
rect 1243 1505 1247 1509
rect 1419 1505 1423 1509
rect 1555 1505 1559 1509
rect 1667 1505 1671 1509
rect 599 1499 603 1503
rect 735 1499 739 1503
rect 871 1499 875 1503
rect 1015 1499 1019 1503
rect 1159 1499 1163 1503
rect 1303 1499 1307 1503
rect 1439 1499 1443 1503
rect 1575 1499 1579 1503
rect 1719 1501 1723 1505
rect 111 1483 115 1487
rect 623 1484 627 1488
rect 759 1484 763 1488
rect 895 1484 899 1488
rect 1039 1484 1043 1488
rect 1183 1484 1187 1488
rect 1327 1484 1331 1488
rect 1463 1484 1467 1488
rect 1599 1484 1603 1488
rect 1719 1483 1723 1487
rect 111 1421 115 1425
rect 599 1420 603 1424
rect 735 1420 739 1424
rect 879 1420 883 1424
rect 1023 1420 1027 1424
rect 1167 1420 1171 1424
rect 1319 1420 1323 1424
rect 1463 1420 1467 1424
rect 1599 1420 1603 1424
rect 1719 1421 1723 1425
rect 111 1403 115 1407
rect 575 1405 579 1409
rect 711 1405 715 1409
rect 855 1405 859 1409
rect 999 1405 1003 1409
rect 1143 1405 1147 1409
rect 1295 1405 1299 1409
rect 1439 1405 1443 1409
rect 1575 1405 1579 1409
rect 691 1399 695 1403
rect 955 1399 956 1403
rect 956 1399 959 1403
rect 667 1391 671 1395
rect 1119 1399 1123 1403
rect 1395 1399 1396 1403
rect 1396 1399 1399 1403
rect 1535 1399 1536 1403
rect 1536 1399 1539 1403
rect 1719 1403 1723 1407
rect 667 1355 671 1359
rect 691 1355 695 1359
rect 1119 1355 1123 1359
rect 1243 1355 1247 1359
rect 1351 1355 1355 1359
rect 1667 1355 1671 1359
rect 295 1331 299 1335
rect 511 1331 515 1335
rect 731 1331 735 1335
rect 955 1331 959 1335
rect 1327 1331 1331 1335
rect 1535 1331 1539 1335
rect 111 1281 115 1285
rect 227 1285 231 1289
rect 295 1287 299 1291
rect 511 1287 515 1291
rect 731 1287 735 1291
rect 1351 1285 1352 1289
rect 1352 1285 1355 1289
rect 1615 1285 1616 1289
rect 1616 1285 1619 1289
rect 135 1279 139 1283
rect 303 1279 307 1283
rect 519 1279 523 1283
rect 751 1279 755 1283
rect 999 1279 1003 1283
rect 1255 1279 1259 1283
rect 1519 1279 1523 1283
rect 1719 1281 1723 1285
rect 111 1263 115 1267
rect 159 1264 163 1268
rect 327 1264 331 1268
rect 543 1264 547 1268
rect 775 1264 779 1268
rect 1023 1264 1027 1268
rect 1279 1264 1283 1268
rect 1543 1264 1547 1268
rect 1719 1263 1723 1267
rect 111 1193 115 1197
rect 159 1192 163 1196
rect 399 1192 403 1196
rect 671 1192 675 1196
rect 959 1192 963 1196
rect 1255 1192 1259 1196
rect 1551 1192 1555 1196
rect 1719 1193 1723 1197
rect 111 1175 115 1179
rect 135 1177 139 1181
rect 375 1177 379 1181
rect 647 1177 651 1181
rect 935 1177 939 1181
rect 1231 1177 1235 1181
rect 1527 1177 1531 1181
rect 235 1171 236 1175
rect 236 1171 239 1175
rect 475 1171 476 1175
rect 476 1171 479 1175
rect 803 1171 807 1175
rect 919 1171 923 1175
rect 1327 1171 1328 1175
rect 1328 1171 1331 1175
rect 1623 1171 1624 1175
rect 1624 1171 1627 1175
rect 1719 1175 1723 1179
rect 283 1151 287 1155
rect 919 1151 923 1155
rect 227 1127 231 1131
rect 235 1127 239 1131
rect 475 1127 479 1131
rect 803 1127 807 1131
rect 1411 1127 1415 1131
rect 1615 1127 1619 1131
rect 283 1119 287 1123
rect 291 1119 295 1123
rect 531 1119 535 1123
rect 787 1119 791 1123
rect 1067 1119 1071 1123
rect 1623 1119 1627 1123
rect 111 1069 115 1073
rect 291 1073 292 1077
rect 292 1073 295 1077
rect 531 1073 535 1077
rect 787 1073 791 1077
rect 1067 1073 1071 1077
rect 1343 1073 1344 1077
rect 1344 1073 1347 1077
rect 1639 1073 1640 1077
rect 1640 1073 1643 1077
rect 191 1067 195 1071
rect 415 1067 419 1071
rect 671 1067 675 1071
rect 951 1067 955 1071
rect 1247 1067 1251 1071
rect 1543 1067 1547 1071
rect 1719 1069 1723 1073
rect 111 1051 115 1055
rect 215 1052 219 1056
rect 439 1052 443 1056
rect 695 1052 699 1056
rect 975 1052 979 1056
rect 1271 1052 1275 1056
rect 1567 1052 1571 1056
rect 1719 1051 1723 1055
rect 111 977 115 981
rect 511 976 515 980
rect 663 976 667 980
rect 831 976 835 980
rect 1007 976 1011 980
rect 1199 976 1203 980
rect 1399 976 1403 980
rect 1599 976 1603 980
rect 1719 977 1723 981
rect 111 959 115 963
rect 487 961 491 965
rect 639 961 643 965
rect 807 961 811 965
rect 983 961 987 965
rect 1175 961 1179 965
rect 1375 961 1379 965
rect 1575 961 1579 965
rect 587 955 588 959
rect 588 955 591 959
rect 739 955 740 959
rect 740 955 743 959
rect 1119 955 1123 959
rect 1159 955 1163 959
rect 1411 955 1415 959
rect 1667 955 1671 959
rect 1719 959 1723 963
rect 579 947 583 951
rect 1343 947 1347 951
rect 579 911 583 915
rect 587 911 591 915
rect 739 911 743 915
rect 1119 911 1123 915
rect 1495 907 1499 911
rect 1639 911 1643 915
rect 1159 899 1163 903
rect 859 891 863 895
rect 1011 891 1015 895
rect 1183 891 1187 895
rect 1339 891 1343 895
rect 1667 891 1671 895
rect 111 841 115 845
rect 859 845 860 849
rect 860 845 863 849
rect 1011 845 1012 849
rect 1012 845 1015 849
rect 1183 845 1187 849
rect 1339 849 1343 851
rect 1339 847 1340 849
rect 1340 847 1343 849
rect 1379 847 1383 851
rect 1667 845 1671 849
rect 759 839 763 843
rect 911 839 915 843
rect 1071 839 1075 843
rect 1239 839 1243 843
rect 1407 839 1411 843
rect 1575 839 1579 843
rect 1719 841 1723 845
rect 111 823 115 827
rect 783 824 787 828
rect 935 824 939 828
rect 1095 824 1099 828
rect 1263 824 1267 828
rect 1431 824 1435 828
rect 1599 824 1603 828
rect 1719 823 1723 827
rect 111 757 115 761
rect 695 756 699 760
rect 831 756 835 760
rect 975 756 979 760
rect 1119 756 1123 760
rect 1271 756 1275 760
rect 1431 756 1435 760
rect 1599 756 1603 760
rect 1719 757 1723 761
rect 111 739 115 743
rect 671 741 675 745
rect 807 741 811 745
rect 951 741 955 745
rect 1095 741 1099 745
rect 1247 741 1251 745
rect 1407 741 1411 745
rect 1575 741 1579 745
rect 791 735 795 739
rect 1051 735 1052 739
rect 1052 735 1055 739
rect 763 727 767 731
rect 1219 735 1223 739
rect 1495 735 1499 739
rect 1651 735 1655 739
rect 1719 739 1723 743
rect 763 691 767 695
rect 791 691 795 695
rect 1219 691 1223 695
rect 1379 691 1383 695
rect 1415 691 1419 695
rect 1667 691 1671 695
rect 623 659 627 663
rect 839 659 843 663
rect 1043 659 1047 663
rect 1051 659 1055 663
rect 1435 659 1439 663
rect 1651 659 1655 663
rect 259 615 263 619
rect 111 609 115 613
rect 623 615 627 619
rect 839 615 843 619
rect 1043 615 1047 619
rect 1415 613 1416 617
rect 1416 613 1419 617
rect 1655 613 1656 617
rect 1656 613 1659 617
rect 247 607 251 611
rect 431 607 435 611
rect 631 607 635 611
rect 847 607 851 611
rect 1079 607 1083 611
rect 1319 607 1323 611
rect 1559 607 1563 611
rect 1719 609 1723 613
rect 111 591 115 595
rect 271 592 275 596
rect 455 592 459 596
rect 655 592 659 596
rect 871 592 875 596
rect 1103 592 1107 596
rect 1343 592 1347 596
rect 1583 592 1587 596
rect 1719 591 1723 595
rect 111 517 115 521
rect 159 516 163 520
rect 343 516 347 520
rect 575 516 579 520
rect 831 516 835 520
rect 1095 516 1099 520
rect 1367 516 1371 520
rect 1719 517 1723 521
rect 111 499 115 503
rect 135 501 139 505
rect 319 501 323 505
rect 551 501 555 505
rect 807 501 811 505
rect 1071 501 1075 505
rect 1343 501 1347 505
rect 419 495 420 499
rect 420 495 423 499
rect 651 495 652 499
rect 652 495 655 499
rect 291 487 295 491
rect 1435 495 1439 499
rect 1719 499 1723 503
rect 255 451 259 455
rect 419 451 423 455
rect 651 451 655 455
rect 1423 451 1427 455
rect 291 431 295 435
rect 299 431 303 435
rect 531 431 535 435
rect 731 431 735 435
rect 1175 431 1179 435
rect 1187 431 1191 435
rect 1655 431 1659 435
rect 111 381 115 385
rect 299 385 300 389
rect 300 385 303 389
rect 531 385 535 389
rect 731 385 732 389
rect 732 385 735 389
rect 951 385 952 389
rect 952 385 955 389
rect 1187 385 1188 389
rect 1188 385 1191 389
rect 1423 385 1424 389
rect 1424 385 1427 389
rect 1675 385 1676 389
rect 1676 385 1679 389
rect 199 379 203 383
rect 415 379 419 383
rect 631 379 635 383
rect 855 379 859 383
rect 1087 379 1091 383
rect 1327 379 1331 383
rect 1575 379 1579 383
rect 1719 381 1723 385
rect 111 363 115 367
rect 223 364 227 368
rect 439 364 443 368
rect 655 364 659 368
rect 879 364 883 368
rect 1111 364 1115 368
rect 1351 364 1355 368
rect 1599 364 1603 368
rect 1719 363 1723 367
rect 111 301 115 305
rect 559 300 563 304
rect 759 300 763 304
rect 967 300 971 304
rect 1183 300 1187 304
rect 1399 300 1403 304
rect 1599 300 1603 304
rect 1719 301 1723 305
rect 111 283 115 287
rect 535 285 539 289
rect 735 285 739 289
rect 943 285 947 289
rect 1159 285 1163 289
rect 1375 285 1379 289
rect 1575 285 1579 289
rect 579 279 583 283
rect 655 279 659 283
rect 887 279 891 283
rect 1175 279 1179 283
rect 1315 279 1319 283
rect 1667 279 1671 283
rect 1719 283 1723 287
rect 655 235 659 239
rect 887 235 891 239
rect 951 235 955 239
rect 1315 235 1319 239
rect 1399 235 1403 239
rect 1675 235 1679 239
rect 579 215 583 219
rect 587 215 591 219
rect 723 215 727 219
rect 875 215 879 219
rect 1011 215 1015 219
rect 1131 215 1135 219
rect 1283 215 1287 219
rect 1531 211 1535 215
rect 1667 215 1671 219
rect 111 165 115 169
rect 587 169 588 173
rect 588 169 591 173
rect 723 169 724 173
rect 724 169 727 173
rect 875 169 879 173
rect 1011 169 1015 173
rect 1131 169 1132 173
rect 1132 169 1135 173
rect 1283 169 1287 173
rect 1399 169 1400 173
rect 1400 169 1403 173
rect 1531 171 1535 175
rect 487 163 491 167
rect 623 163 627 167
rect 759 163 763 167
rect 895 163 899 167
rect 1031 163 1035 167
rect 1167 163 1171 167
rect 1303 163 1307 167
rect 1439 163 1443 167
rect 1575 163 1579 167
rect 1719 165 1723 169
rect 111 147 115 151
rect 511 148 515 152
rect 647 148 651 152
rect 783 148 787 152
rect 919 148 923 152
rect 1055 148 1059 152
rect 1191 148 1195 152
rect 1327 148 1331 152
rect 1463 148 1467 152
rect 1599 148 1603 152
rect 1719 147 1723 151
<< m3 >>
rect 111 1782 115 1783
rect 111 1777 115 1778
rect 135 1782 139 1783
rect 271 1782 275 1783
rect 135 1777 139 1778
rect 250 1779 256 1780
rect 112 1730 114 1777
rect 110 1729 116 1730
rect 110 1725 111 1729
rect 115 1725 116 1729
rect 136 1728 138 1777
rect 250 1775 251 1779
rect 255 1775 256 1779
rect 407 1782 411 1783
rect 271 1777 275 1778
rect 386 1779 392 1780
rect 250 1774 256 1775
rect 252 1734 254 1774
rect 250 1733 256 1734
rect 250 1729 251 1733
rect 255 1729 256 1733
rect 250 1728 256 1729
rect 272 1728 274 1777
rect 386 1775 387 1779
rect 391 1775 392 1779
rect 543 1782 547 1783
rect 407 1777 411 1778
rect 522 1779 528 1780
rect 386 1774 392 1775
rect 388 1734 390 1774
rect 386 1733 392 1734
rect 386 1729 387 1733
rect 391 1729 392 1733
rect 386 1728 392 1729
rect 408 1728 410 1777
rect 522 1775 523 1779
rect 527 1775 528 1779
rect 679 1782 683 1783
rect 543 1777 547 1778
rect 658 1779 664 1780
rect 522 1774 528 1775
rect 524 1734 526 1774
rect 522 1733 528 1734
rect 522 1729 523 1733
rect 527 1729 528 1733
rect 522 1728 528 1729
rect 544 1728 546 1777
rect 658 1775 659 1779
rect 663 1775 664 1779
rect 679 1777 683 1778
rect 1719 1782 1723 1783
rect 1719 1777 1723 1778
rect 658 1774 664 1775
rect 660 1734 662 1774
rect 658 1733 664 1734
rect 658 1729 659 1733
rect 663 1729 664 1733
rect 658 1728 664 1729
rect 680 1728 682 1777
rect 774 1733 780 1734
rect 774 1729 775 1733
rect 779 1729 780 1733
rect 1720 1730 1722 1777
rect 774 1728 780 1729
rect 1718 1729 1724 1730
rect 110 1724 116 1725
rect 134 1727 140 1728
rect 134 1723 135 1727
rect 139 1723 140 1727
rect 134 1722 140 1723
rect 270 1727 276 1728
rect 270 1723 271 1727
rect 275 1723 276 1727
rect 270 1722 276 1723
rect 406 1727 412 1728
rect 406 1723 407 1727
rect 411 1723 412 1727
rect 406 1722 412 1723
rect 542 1727 548 1728
rect 542 1723 543 1727
rect 547 1723 548 1727
rect 542 1722 548 1723
rect 678 1727 684 1728
rect 678 1723 679 1727
rect 683 1723 684 1727
rect 678 1722 684 1723
rect 158 1712 164 1713
rect 110 1711 116 1712
rect 110 1707 111 1711
rect 115 1707 116 1711
rect 158 1708 159 1712
rect 163 1708 164 1712
rect 158 1707 164 1708
rect 294 1712 300 1713
rect 294 1708 295 1712
rect 299 1708 300 1712
rect 294 1707 300 1708
rect 430 1712 436 1713
rect 430 1708 431 1712
rect 435 1708 436 1712
rect 430 1707 436 1708
rect 566 1712 572 1713
rect 566 1708 567 1712
rect 571 1708 572 1712
rect 566 1707 572 1708
rect 702 1712 708 1713
rect 702 1708 703 1712
rect 707 1708 708 1712
rect 702 1707 708 1708
rect 110 1706 116 1707
rect 112 1675 114 1706
rect 160 1675 162 1707
rect 296 1675 298 1707
rect 306 1675 312 1676
rect 432 1675 434 1707
rect 568 1675 570 1707
rect 704 1675 706 1707
rect 776 1676 778 1728
rect 1718 1725 1719 1729
rect 1723 1725 1724 1729
rect 1718 1724 1724 1725
rect 1718 1711 1724 1712
rect 1718 1707 1719 1711
rect 1723 1707 1724 1711
rect 1718 1706 1724 1707
rect 774 1675 780 1676
rect 1720 1675 1722 1706
rect 111 1674 115 1675
rect 111 1669 115 1670
rect 159 1674 163 1675
rect 159 1669 163 1670
rect 239 1674 243 1675
rect 239 1669 243 1670
rect 295 1674 299 1675
rect 306 1671 307 1675
rect 311 1671 312 1675
rect 306 1670 312 1671
rect 375 1674 379 1675
rect 295 1669 299 1670
rect 112 1646 114 1669
rect 110 1645 116 1646
rect 240 1645 242 1669
rect 110 1641 111 1645
rect 115 1641 116 1645
rect 110 1640 116 1641
rect 238 1644 244 1645
rect 238 1640 239 1644
rect 243 1640 244 1644
rect 238 1639 244 1640
rect 214 1629 220 1630
rect 110 1627 116 1628
rect 110 1623 111 1627
rect 115 1623 116 1627
rect 214 1625 215 1629
rect 219 1625 220 1629
rect 214 1624 220 1625
rect 110 1622 116 1623
rect 112 1559 114 1622
rect 216 1559 218 1624
rect 308 1580 310 1670
rect 375 1669 379 1670
rect 431 1674 435 1675
rect 431 1669 435 1670
rect 511 1674 515 1675
rect 511 1669 515 1670
rect 567 1674 571 1675
rect 567 1669 571 1670
rect 647 1674 651 1675
rect 647 1669 651 1670
rect 703 1674 707 1675
rect 774 1671 775 1675
rect 779 1671 780 1675
rect 774 1670 780 1671
rect 783 1674 787 1675
rect 703 1669 707 1670
rect 783 1669 787 1670
rect 1719 1674 1723 1675
rect 1719 1669 1723 1670
rect 376 1645 378 1669
rect 512 1645 514 1669
rect 648 1645 650 1669
rect 784 1645 786 1669
rect 1720 1646 1722 1669
rect 1718 1645 1724 1646
rect 374 1644 380 1645
rect 374 1640 375 1644
rect 379 1640 380 1644
rect 374 1639 380 1640
rect 510 1644 516 1645
rect 510 1640 511 1644
rect 515 1640 516 1644
rect 510 1639 516 1640
rect 646 1644 652 1645
rect 646 1640 647 1644
rect 651 1640 652 1644
rect 646 1639 652 1640
rect 782 1644 788 1645
rect 782 1640 783 1644
rect 787 1640 788 1644
rect 1718 1641 1719 1645
rect 1723 1641 1724 1645
rect 1718 1640 1724 1641
rect 782 1639 788 1640
rect 350 1629 356 1630
rect 350 1625 351 1629
rect 355 1625 356 1629
rect 350 1624 356 1625
rect 486 1629 492 1630
rect 486 1625 487 1629
rect 491 1625 492 1629
rect 486 1624 492 1625
rect 622 1629 628 1630
rect 622 1625 623 1629
rect 627 1625 628 1629
rect 622 1624 628 1625
rect 758 1629 764 1630
rect 758 1625 759 1629
rect 763 1625 764 1629
rect 758 1624 764 1625
rect 1718 1627 1724 1628
rect 330 1623 336 1624
rect 330 1619 331 1623
rect 335 1619 336 1623
rect 330 1618 336 1619
rect 332 1580 334 1618
rect 306 1579 312 1580
rect 306 1575 307 1579
rect 311 1575 312 1579
rect 306 1574 312 1575
rect 330 1579 336 1580
rect 330 1575 331 1579
rect 335 1575 336 1579
rect 330 1574 336 1575
rect 352 1559 354 1624
rect 466 1623 472 1624
rect 466 1619 467 1623
rect 471 1619 472 1623
rect 466 1618 472 1619
rect 468 1580 470 1618
rect 466 1579 472 1580
rect 466 1575 467 1579
rect 471 1575 472 1579
rect 466 1574 472 1575
rect 488 1559 490 1624
rect 586 1619 592 1620
rect 586 1615 587 1619
rect 591 1615 592 1619
rect 586 1614 592 1615
rect 588 1580 590 1614
rect 586 1579 592 1580
rect 586 1575 587 1579
rect 591 1575 592 1579
rect 586 1574 592 1575
rect 624 1559 626 1624
rect 738 1623 744 1624
rect 738 1619 739 1623
rect 743 1619 744 1623
rect 738 1618 744 1619
rect 690 1615 696 1616
rect 690 1611 691 1615
rect 695 1611 696 1615
rect 690 1610 696 1611
rect 111 1558 115 1559
rect 111 1553 115 1554
rect 215 1558 219 1559
rect 215 1553 219 1554
rect 351 1558 355 1559
rect 351 1553 355 1554
rect 487 1558 491 1559
rect 487 1553 491 1554
rect 599 1558 603 1559
rect 599 1553 603 1554
rect 623 1558 627 1559
rect 692 1556 694 1610
rect 740 1580 742 1618
rect 738 1579 744 1580
rect 738 1575 739 1579
rect 743 1575 744 1579
rect 738 1574 744 1575
rect 760 1559 762 1624
rect 1718 1623 1719 1627
rect 1723 1623 1724 1627
rect 1718 1622 1724 1623
rect 1720 1559 1722 1622
rect 735 1558 739 1559
rect 623 1553 627 1554
rect 690 1555 696 1556
rect 112 1506 114 1553
rect 110 1505 116 1506
rect 110 1501 111 1505
rect 115 1501 116 1505
rect 600 1504 602 1553
rect 690 1551 691 1555
rect 695 1551 696 1555
rect 690 1550 696 1551
rect 714 1555 720 1556
rect 714 1551 715 1555
rect 719 1551 720 1555
rect 735 1553 739 1554
rect 759 1558 763 1559
rect 871 1558 875 1559
rect 759 1553 763 1554
rect 862 1555 868 1556
rect 714 1550 720 1551
rect 716 1510 718 1550
rect 714 1509 720 1510
rect 714 1505 715 1509
rect 719 1505 720 1509
rect 714 1504 720 1505
rect 736 1504 738 1553
rect 862 1551 863 1555
rect 867 1551 868 1555
rect 1015 1558 1019 1559
rect 871 1553 875 1554
rect 970 1555 976 1556
rect 862 1550 868 1551
rect 864 1512 866 1550
rect 862 1511 868 1512
rect 862 1507 863 1511
rect 867 1507 868 1511
rect 862 1506 868 1507
rect 872 1504 874 1553
rect 970 1551 971 1555
rect 975 1551 976 1555
rect 1159 1558 1163 1559
rect 1015 1553 1019 1554
rect 1114 1555 1120 1556
rect 970 1550 976 1551
rect 972 1510 974 1550
rect 970 1509 976 1510
rect 970 1505 971 1509
rect 975 1505 976 1509
rect 970 1504 976 1505
rect 1016 1504 1018 1553
rect 1114 1551 1115 1555
rect 1119 1551 1120 1555
rect 1159 1553 1163 1554
rect 1303 1558 1307 1559
rect 1439 1558 1443 1559
rect 1303 1553 1307 1554
rect 1418 1555 1424 1556
rect 1114 1550 1120 1551
rect 1116 1510 1118 1550
rect 1114 1509 1120 1510
rect 1114 1505 1115 1509
rect 1119 1505 1120 1509
rect 1114 1504 1120 1505
rect 1160 1504 1162 1553
rect 1242 1509 1248 1510
rect 1242 1505 1243 1509
rect 1247 1505 1248 1509
rect 1242 1504 1248 1505
rect 1304 1504 1306 1553
rect 1394 1551 1400 1552
rect 1394 1547 1395 1551
rect 1399 1547 1400 1551
rect 1418 1551 1419 1555
rect 1423 1551 1424 1555
rect 1575 1558 1579 1559
rect 1439 1553 1443 1554
rect 1554 1555 1560 1556
rect 1418 1550 1424 1551
rect 1394 1546 1400 1547
rect 110 1500 116 1501
rect 598 1503 604 1504
rect 598 1499 599 1503
rect 603 1499 604 1503
rect 598 1498 604 1499
rect 734 1503 740 1504
rect 734 1499 735 1503
rect 739 1499 740 1503
rect 734 1498 740 1499
rect 870 1503 876 1504
rect 870 1499 871 1503
rect 875 1499 876 1503
rect 870 1498 876 1499
rect 1014 1503 1020 1504
rect 1014 1499 1015 1503
rect 1019 1499 1020 1503
rect 1014 1498 1020 1499
rect 1158 1503 1164 1504
rect 1158 1499 1159 1503
rect 1163 1499 1164 1503
rect 1158 1498 1164 1499
rect 622 1488 628 1489
rect 110 1487 116 1488
rect 110 1483 111 1487
rect 115 1483 116 1487
rect 622 1484 623 1488
rect 627 1484 628 1488
rect 622 1483 628 1484
rect 758 1488 764 1489
rect 758 1484 759 1488
rect 763 1484 764 1488
rect 758 1483 764 1484
rect 894 1488 900 1489
rect 894 1484 895 1488
rect 899 1484 900 1488
rect 894 1483 900 1484
rect 1038 1488 1044 1489
rect 1038 1484 1039 1488
rect 1043 1484 1044 1488
rect 1038 1483 1044 1484
rect 1182 1488 1188 1489
rect 1182 1484 1183 1488
rect 1187 1484 1188 1488
rect 1182 1483 1188 1484
rect 110 1482 116 1483
rect 112 1455 114 1482
rect 624 1455 626 1483
rect 760 1455 762 1483
rect 896 1455 898 1483
rect 1040 1455 1042 1483
rect 1184 1455 1186 1483
rect 111 1454 115 1455
rect 111 1449 115 1450
rect 599 1454 603 1455
rect 599 1449 603 1450
rect 623 1454 627 1455
rect 623 1449 627 1450
rect 735 1454 739 1455
rect 735 1449 739 1450
rect 759 1454 763 1455
rect 759 1449 763 1450
rect 879 1454 883 1455
rect 879 1449 883 1450
rect 895 1454 899 1455
rect 895 1449 899 1450
rect 1023 1454 1027 1455
rect 1023 1449 1027 1450
rect 1039 1454 1043 1455
rect 1039 1449 1043 1450
rect 1167 1454 1171 1455
rect 1167 1449 1171 1450
rect 1183 1454 1187 1455
rect 1183 1449 1187 1450
rect 112 1426 114 1449
rect 110 1425 116 1426
rect 600 1425 602 1449
rect 736 1425 738 1449
rect 880 1425 882 1449
rect 1024 1425 1026 1449
rect 1168 1425 1170 1449
rect 110 1421 111 1425
rect 115 1421 116 1425
rect 110 1420 116 1421
rect 598 1424 604 1425
rect 598 1420 599 1424
rect 603 1420 604 1424
rect 598 1419 604 1420
rect 734 1424 740 1425
rect 734 1420 735 1424
rect 739 1420 740 1424
rect 734 1419 740 1420
rect 878 1424 884 1425
rect 878 1420 879 1424
rect 883 1420 884 1424
rect 878 1419 884 1420
rect 1022 1424 1028 1425
rect 1022 1420 1023 1424
rect 1027 1420 1028 1424
rect 1022 1419 1028 1420
rect 1166 1424 1172 1425
rect 1166 1420 1167 1424
rect 1171 1420 1172 1424
rect 1166 1419 1172 1420
rect 574 1409 580 1410
rect 110 1407 116 1408
rect 110 1403 111 1407
rect 115 1403 116 1407
rect 574 1405 575 1409
rect 579 1405 580 1409
rect 574 1404 580 1405
rect 710 1409 716 1410
rect 710 1405 711 1409
rect 715 1405 716 1409
rect 710 1404 716 1405
rect 854 1409 860 1410
rect 854 1405 855 1409
rect 859 1405 860 1409
rect 854 1404 860 1405
rect 998 1409 1004 1410
rect 998 1405 999 1409
rect 1003 1405 1004 1409
rect 998 1404 1004 1405
rect 1142 1409 1148 1410
rect 1142 1405 1143 1409
rect 1147 1405 1148 1409
rect 1142 1404 1148 1405
rect 110 1402 116 1403
rect 112 1339 114 1402
rect 576 1339 578 1404
rect 690 1403 696 1404
rect 690 1399 691 1403
rect 695 1399 696 1403
rect 690 1398 696 1399
rect 666 1395 672 1396
rect 666 1391 667 1395
rect 671 1391 672 1395
rect 666 1390 672 1391
rect 668 1360 670 1390
rect 692 1360 694 1398
rect 666 1359 672 1360
rect 666 1355 667 1359
rect 671 1355 672 1359
rect 666 1354 672 1355
rect 690 1359 696 1360
rect 690 1355 691 1359
rect 695 1355 696 1359
rect 690 1354 696 1355
rect 712 1339 714 1404
rect 856 1339 858 1404
rect 954 1403 960 1404
rect 954 1399 955 1403
rect 959 1399 960 1403
rect 954 1398 960 1399
rect 111 1338 115 1339
rect 111 1333 115 1334
rect 135 1338 139 1339
rect 303 1338 307 1339
rect 135 1333 139 1334
rect 294 1335 300 1336
rect 112 1286 114 1333
rect 110 1285 116 1286
rect 110 1281 111 1285
rect 115 1281 116 1285
rect 136 1284 138 1333
rect 294 1331 295 1335
rect 299 1331 300 1335
rect 519 1338 523 1339
rect 303 1333 307 1334
rect 510 1335 516 1336
rect 294 1330 300 1331
rect 296 1292 298 1330
rect 294 1291 300 1292
rect 226 1289 232 1290
rect 226 1285 227 1289
rect 231 1285 232 1289
rect 294 1287 295 1291
rect 299 1287 300 1291
rect 294 1286 300 1287
rect 226 1284 232 1285
rect 304 1284 306 1333
rect 510 1331 511 1335
rect 515 1331 516 1335
rect 519 1333 523 1334
rect 575 1338 579 1339
rect 575 1333 579 1334
rect 711 1338 715 1339
rect 751 1338 755 1339
rect 711 1333 715 1334
rect 730 1335 736 1336
rect 510 1330 516 1331
rect 512 1292 514 1330
rect 510 1291 516 1292
rect 510 1287 511 1291
rect 515 1287 516 1291
rect 510 1286 516 1287
rect 520 1284 522 1333
rect 730 1331 731 1335
rect 735 1331 736 1335
rect 751 1333 755 1334
rect 855 1338 859 1339
rect 956 1336 958 1398
rect 1000 1339 1002 1404
rect 1118 1403 1124 1404
rect 1118 1399 1119 1403
rect 1123 1399 1124 1403
rect 1118 1398 1124 1399
rect 1120 1360 1122 1398
rect 1118 1359 1124 1360
rect 1118 1355 1119 1359
rect 1123 1355 1124 1359
rect 1118 1354 1124 1355
rect 1144 1339 1146 1404
rect 1244 1360 1246 1504
rect 1302 1503 1308 1504
rect 1302 1499 1303 1503
rect 1307 1499 1308 1503
rect 1302 1498 1308 1499
rect 1326 1488 1332 1489
rect 1326 1484 1327 1488
rect 1331 1484 1332 1488
rect 1326 1483 1332 1484
rect 1328 1455 1330 1483
rect 1319 1454 1323 1455
rect 1319 1449 1323 1450
rect 1327 1454 1331 1455
rect 1327 1449 1331 1450
rect 1320 1425 1322 1449
rect 1318 1424 1324 1425
rect 1318 1420 1319 1424
rect 1323 1420 1324 1424
rect 1318 1419 1324 1420
rect 1294 1409 1300 1410
rect 1294 1405 1295 1409
rect 1299 1405 1300 1409
rect 1294 1404 1300 1405
rect 1396 1404 1398 1546
rect 1420 1510 1422 1550
rect 1418 1509 1424 1510
rect 1418 1505 1419 1509
rect 1423 1505 1424 1509
rect 1418 1504 1424 1505
rect 1440 1504 1442 1553
rect 1554 1551 1555 1555
rect 1559 1551 1560 1555
rect 1575 1553 1579 1554
rect 1719 1558 1723 1559
rect 1719 1553 1723 1554
rect 1554 1550 1560 1551
rect 1556 1510 1558 1550
rect 1554 1509 1560 1510
rect 1554 1505 1555 1509
rect 1559 1505 1560 1509
rect 1554 1504 1560 1505
rect 1576 1504 1578 1553
rect 1666 1509 1672 1510
rect 1666 1505 1667 1509
rect 1671 1505 1672 1509
rect 1720 1506 1722 1553
rect 1666 1504 1672 1505
rect 1718 1505 1724 1506
rect 1438 1503 1444 1504
rect 1438 1499 1439 1503
rect 1443 1499 1444 1503
rect 1438 1498 1444 1499
rect 1574 1503 1580 1504
rect 1574 1499 1575 1503
rect 1579 1499 1580 1503
rect 1574 1498 1580 1499
rect 1462 1488 1468 1489
rect 1462 1484 1463 1488
rect 1467 1484 1468 1488
rect 1462 1483 1468 1484
rect 1598 1488 1604 1489
rect 1598 1484 1599 1488
rect 1603 1484 1604 1488
rect 1598 1483 1604 1484
rect 1464 1455 1466 1483
rect 1600 1455 1602 1483
rect 1463 1454 1467 1455
rect 1463 1449 1467 1450
rect 1599 1454 1603 1455
rect 1599 1449 1603 1450
rect 1464 1425 1466 1449
rect 1600 1425 1602 1449
rect 1462 1424 1468 1425
rect 1462 1420 1463 1424
rect 1467 1420 1468 1424
rect 1462 1419 1468 1420
rect 1598 1424 1604 1425
rect 1598 1420 1599 1424
rect 1603 1420 1604 1424
rect 1598 1419 1604 1420
rect 1438 1409 1444 1410
rect 1438 1405 1439 1409
rect 1443 1405 1444 1409
rect 1438 1404 1444 1405
rect 1574 1409 1580 1410
rect 1574 1405 1575 1409
rect 1579 1405 1580 1409
rect 1574 1404 1580 1405
rect 1242 1359 1248 1360
rect 1242 1355 1243 1359
rect 1247 1355 1248 1359
rect 1242 1354 1248 1355
rect 1296 1339 1298 1404
rect 1394 1403 1400 1404
rect 1394 1399 1395 1403
rect 1399 1399 1400 1403
rect 1394 1398 1400 1399
rect 1350 1359 1356 1360
rect 1350 1355 1351 1359
rect 1355 1355 1356 1359
rect 1350 1354 1356 1355
rect 999 1338 1003 1339
rect 855 1333 859 1334
rect 954 1335 960 1336
rect 730 1330 736 1331
rect 732 1292 734 1330
rect 730 1291 736 1292
rect 730 1287 731 1291
rect 735 1287 736 1291
rect 730 1286 736 1287
rect 752 1284 754 1333
rect 954 1331 955 1335
rect 959 1331 960 1335
rect 999 1333 1003 1334
rect 1143 1338 1147 1339
rect 1143 1333 1147 1334
rect 1255 1338 1259 1339
rect 1255 1333 1259 1334
rect 1295 1338 1299 1339
rect 1295 1333 1299 1334
rect 1326 1335 1332 1336
rect 954 1330 960 1331
rect 1000 1284 1002 1333
rect 1256 1284 1258 1333
rect 1326 1331 1327 1335
rect 1331 1331 1332 1335
rect 1326 1330 1332 1331
rect 110 1280 116 1281
rect 134 1283 140 1284
rect 134 1279 135 1283
rect 139 1279 140 1283
rect 134 1278 140 1279
rect 158 1268 164 1269
rect 110 1267 116 1268
rect 110 1263 111 1267
rect 115 1263 116 1267
rect 158 1264 159 1268
rect 163 1264 164 1268
rect 158 1263 164 1264
rect 110 1262 116 1263
rect 112 1227 114 1262
rect 160 1227 162 1263
rect 111 1226 115 1227
rect 111 1221 115 1222
rect 159 1226 163 1227
rect 159 1221 163 1222
rect 112 1198 114 1221
rect 110 1197 116 1198
rect 160 1197 162 1221
rect 110 1193 111 1197
rect 115 1193 116 1197
rect 110 1192 116 1193
rect 158 1196 164 1197
rect 158 1192 159 1196
rect 163 1192 164 1196
rect 158 1191 164 1192
rect 134 1181 140 1182
rect 110 1179 116 1180
rect 110 1175 111 1179
rect 115 1175 116 1179
rect 134 1177 135 1181
rect 139 1177 140 1181
rect 134 1176 140 1177
rect 110 1174 116 1175
rect 112 1127 114 1174
rect 136 1127 138 1176
rect 228 1132 230 1284
rect 302 1283 308 1284
rect 302 1279 303 1283
rect 307 1279 308 1283
rect 302 1278 308 1279
rect 518 1283 524 1284
rect 518 1279 519 1283
rect 523 1279 524 1283
rect 518 1278 524 1279
rect 750 1283 756 1284
rect 750 1279 751 1283
rect 755 1279 756 1283
rect 750 1278 756 1279
rect 998 1283 1004 1284
rect 998 1279 999 1283
rect 1003 1279 1004 1283
rect 998 1278 1004 1279
rect 1254 1283 1260 1284
rect 1254 1279 1255 1283
rect 1259 1279 1260 1283
rect 1254 1278 1260 1279
rect 326 1268 332 1269
rect 326 1264 327 1268
rect 331 1264 332 1268
rect 326 1263 332 1264
rect 542 1268 548 1269
rect 542 1264 543 1268
rect 547 1264 548 1268
rect 542 1263 548 1264
rect 774 1268 780 1269
rect 774 1264 775 1268
rect 779 1264 780 1268
rect 774 1263 780 1264
rect 1022 1268 1028 1269
rect 1022 1264 1023 1268
rect 1027 1264 1028 1268
rect 1022 1263 1028 1264
rect 1278 1268 1284 1269
rect 1278 1264 1279 1268
rect 1283 1264 1284 1268
rect 1278 1263 1284 1264
rect 328 1227 330 1263
rect 544 1227 546 1263
rect 776 1227 778 1263
rect 1024 1227 1026 1263
rect 1280 1227 1282 1263
rect 327 1226 331 1227
rect 327 1221 331 1222
rect 399 1226 403 1227
rect 399 1221 403 1222
rect 543 1226 547 1227
rect 543 1221 547 1222
rect 671 1226 675 1227
rect 671 1221 675 1222
rect 775 1226 779 1227
rect 775 1221 779 1222
rect 959 1226 963 1227
rect 959 1221 963 1222
rect 1023 1226 1027 1227
rect 1023 1221 1027 1222
rect 1255 1226 1259 1227
rect 1255 1221 1259 1222
rect 1279 1226 1283 1227
rect 1279 1221 1283 1222
rect 400 1197 402 1221
rect 672 1197 674 1221
rect 960 1197 962 1221
rect 1256 1197 1258 1221
rect 398 1196 404 1197
rect 398 1192 399 1196
rect 403 1192 404 1196
rect 398 1191 404 1192
rect 670 1196 676 1197
rect 670 1192 671 1196
rect 675 1192 676 1196
rect 670 1191 676 1192
rect 958 1196 964 1197
rect 958 1192 959 1196
rect 963 1192 964 1196
rect 958 1191 964 1192
rect 1254 1196 1260 1197
rect 1254 1192 1255 1196
rect 1259 1192 1260 1196
rect 1254 1191 1260 1192
rect 374 1181 380 1182
rect 374 1177 375 1181
rect 379 1177 380 1181
rect 374 1176 380 1177
rect 646 1181 652 1182
rect 646 1177 647 1181
rect 651 1177 652 1181
rect 646 1176 652 1177
rect 934 1181 940 1182
rect 934 1177 935 1181
rect 939 1177 940 1181
rect 934 1176 940 1177
rect 1230 1181 1236 1182
rect 1230 1177 1231 1181
rect 1235 1177 1236 1181
rect 1230 1176 1236 1177
rect 1328 1176 1330 1330
rect 1352 1290 1354 1354
rect 1440 1339 1442 1404
rect 1534 1403 1540 1404
rect 1534 1399 1535 1403
rect 1539 1399 1540 1403
rect 1534 1398 1540 1399
rect 1439 1338 1443 1339
rect 1439 1333 1443 1334
rect 1519 1338 1523 1339
rect 1536 1336 1538 1398
rect 1576 1339 1578 1404
rect 1668 1360 1670 1504
rect 1718 1501 1719 1505
rect 1723 1501 1724 1505
rect 1718 1500 1724 1501
rect 1718 1487 1724 1488
rect 1718 1483 1719 1487
rect 1723 1483 1724 1487
rect 1718 1482 1724 1483
rect 1720 1455 1722 1482
rect 1719 1454 1723 1455
rect 1719 1449 1723 1450
rect 1720 1426 1722 1449
rect 1718 1425 1724 1426
rect 1718 1421 1719 1425
rect 1723 1421 1724 1425
rect 1718 1420 1724 1421
rect 1718 1407 1724 1408
rect 1718 1403 1719 1407
rect 1723 1403 1724 1407
rect 1718 1402 1724 1403
rect 1666 1359 1672 1360
rect 1666 1355 1667 1359
rect 1671 1355 1672 1359
rect 1666 1354 1672 1355
rect 1720 1339 1722 1402
rect 1575 1338 1579 1339
rect 1519 1333 1523 1334
rect 1534 1335 1540 1336
rect 1350 1289 1356 1290
rect 1350 1285 1351 1289
rect 1355 1285 1356 1289
rect 1350 1284 1356 1285
rect 1520 1284 1522 1333
rect 1534 1331 1535 1335
rect 1539 1331 1540 1335
rect 1575 1333 1579 1334
rect 1719 1338 1723 1339
rect 1719 1333 1723 1334
rect 1534 1330 1540 1331
rect 1614 1289 1620 1290
rect 1614 1285 1615 1289
rect 1619 1285 1620 1289
rect 1720 1286 1722 1333
rect 1614 1284 1620 1285
rect 1718 1285 1724 1286
rect 1518 1283 1524 1284
rect 1518 1279 1519 1283
rect 1523 1279 1524 1283
rect 1518 1278 1524 1279
rect 1542 1268 1548 1269
rect 1542 1264 1543 1268
rect 1547 1264 1548 1268
rect 1542 1263 1548 1264
rect 1544 1227 1546 1263
rect 1543 1226 1547 1227
rect 1543 1221 1547 1222
rect 1551 1226 1555 1227
rect 1551 1221 1555 1222
rect 1552 1197 1554 1221
rect 1550 1196 1556 1197
rect 1550 1192 1551 1196
rect 1555 1192 1556 1196
rect 1550 1191 1556 1192
rect 1526 1181 1532 1182
rect 1526 1177 1527 1181
rect 1531 1177 1532 1181
rect 1526 1176 1532 1177
rect 234 1175 240 1176
rect 234 1171 235 1175
rect 239 1171 240 1175
rect 234 1170 240 1171
rect 236 1132 238 1170
rect 282 1155 288 1156
rect 282 1151 283 1155
rect 287 1151 288 1155
rect 282 1150 288 1151
rect 226 1131 232 1132
rect 226 1127 227 1131
rect 231 1127 232 1131
rect 111 1126 115 1127
rect 111 1121 115 1122
rect 135 1126 139 1127
rect 135 1121 139 1122
rect 191 1126 195 1127
rect 226 1126 232 1127
rect 234 1131 240 1132
rect 234 1127 235 1131
rect 239 1127 240 1131
rect 234 1126 240 1127
rect 284 1124 286 1150
rect 376 1127 378 1176
rect 474 1175 480 1176
rect 474 1171 475 1175
rect 479 1171 480 1175
rect 474 1170 480 1171
rect 476 1132 478 1170
rect 474 1131 480 1132
rect 474 1127 475 1131
rect 479 1127 480 1131
rect 648 1127 650 1176
rect 802 1175 808 1176
rect 802 1171 803 1175
rect 807 1171 808 1175
rect 802 1170 808 1171
rect 918 1175 924 1176
rect 918 1171 919 1175
rect 923 1171 924 1175
rect 918 1170 924 1171
rect 804 1132 806 1170
rect 920 1156 922 1170
rect 918 1155 924 1156
rect 918 1151 919 1155
rect 923 1151 924 1155
rect 918 1150 924 1151
rect 802 1131 808 1132
rect 802 1127 803 1131
rect 807 1127 808 1131
rect 936 1127 938 1176
rect 1232 1127 1234 1176
rect 1326 1175 1332 1176
rect 1326 1171 1327 1175
rect 1331 1171 1332 1175
rect 1326 1170 1332 1171
rect 1410 1131 1416 1132
rect 1410 1127 1411 1131
rect 1415 1127 1416 1131
rect 1528 1127 1530 1176
rect 1616 1132 1618 1284
rect 1718 1281 1719 1285
rect 1723 1281 1724 1285
rect 1718 1280 1724 1281
rect 1718 1267 1724 1268
rect 1718 1263 1719 1267
rect 1723 1263 1724 1267
rect 1718 1262 1724 1263
rect 1720 1227 1722 1262
rect 1719 1226 1723 1227
rect 1719 1221 1723 1222
rect 1720 1198 1722 1221
rect 1718 1197 1724 1198
rect 1718 1193 1719 1197
rect 1723 1193 1724 1197
rect 1718 1192 1724 1193
rect 1718 1179 1724 1180
rect 1622 1175 1628 1176
rect 1622 1171 1623 1175
rect 1627 1171 1628 1175
rect 1718 1175 1719 1179
rect 1723 1175 1724 1179
rect 1718 1174 1724 1175
rect 1622 1170 1628 1171
rect 1614 1131 1620 1132
rect 1614 1127 1615 1131
rect 1619 1127 1620 1131
rect 375 1126 379 1127
rect 191 1121 195 1122
rect 282 1123 288 1124
rect 112 1074 114 1121
rect 110 1073 116 1074
rect 110 1069 111 1073
rect 115 1069 116 1073
rect 192 1072 194 1121
rect 282 1119 283 1123
rect 287 1119 288 1123
rect 282 1118 288 1119
rect 290 1123 296 1124
rect 290 1119 291 1123
rect 295 1119 296 1123
rect 375 1121 379 1122
rect 415 1126 419 1127
rect 474 1126 480 1127
rect 647 1126 651 1127
rect 415 1121 419 1122
rect 530 1123 536 1124
rect 290 1118 296 1119
rect 292 1078 294 1118
rect 290 1077 296 1078
rect 290 1073 291 1077
rect 295 1073 296 1077
rect 290 1072 296 1073
rect 416 1072 418 1121
rect 530 1119 531 1123
rect 535 1119 536 1123
rect 647 1121 651 1122
rect 671 1126 675 1127
rect 802 1126 808 1127
rect 935 1126 939 1127
rect 671 1121 675 1122
rect 786 1123 792 1124
rect 530 1118 536 1119
rect 532 1078 534 1118
rect 530 1077 536 1078
rect 530 1073 531 1077
rect 535 1073 536 1077
rect 530 1072 536 1073
rect 672 1072 674 1121
rect 786 1119 787 1123
rect 791 1119 792 1123
rect 935 1121 939 1122
rect 951 1126 955 1127
rect 1231 1126 1235 1127
rect 951 1121 955 1122
rect 1066 1123 1072 1124
rect 786 1118 792 1119
rect 788 1078 790 1118
rect 786 1077 792 1078
rect 786 1073 787 1077
rect 791 1073 792 1077
rect 786 1072 792 1073
rect 952 1072 954 1121
rect 1066 1119 1067 1123
rect 1071 1119 1072 1123
rect 1231 1121 1235 1122
rect 1247 1126 1251 1127
rect 1410 1126 1416 1127
rect 1527 1126 1531 1127
rect 1247 1121 1251 1122
rect 1066 1118 1072 1119
rect 1068 1078 1070 1118
rect 1066 1077 1072 1078
rect 1066 1073 1067 1077
rect 1071 1073 1072 1077
rect 1066 1072 1072 1073
rect 1248 1072 1250 1121
rect 1342 1077 1348 1078
rect 1342 1073 1343 1077
rect 1347 1073 1348 1077
rect 1342 1072 1348 1073
rect 110 1068 116 1069
rect 190 1071 196 1072
rect 190 1067 191 1071
rect 195 1067 196 1071
rect 190 1066 196 1067
rect 414 1071 420 1072
rect 414 1067 415 1071
rect 419 1067 420 1071
rect 414 1066 420 1067
rect 670 1071 676 1072
rect 670 1067 671 1071
rect 675 1067 676 1071
rect 670 1066 676 1067
rect 950 1071 956 1072
rect 950 1067 951 1071
rect 955 1067 956 1071
rect 950 1066 956 1067
rect 1246 1071 1252 1072
rect 1246 1067 1247 1071
rect 1251 1067 1252 1071
rect 1246 1066 1252 1067
rect 214 1056 220 1057
rect 110 1055 116 1056
rect 110 1051 111 1055
rect 115 1051 116 1055
rect 214 1052 215 1056
rect 219 1052 220 1056
rect 214 1051 220 1052
rect 438 1056 444 1057
rect 438 1052 439 1056
rect 443 1052 444 1056
rect 438 1051 444 1052
rect 694 1056 700 1057
rect 694 1052 695 1056
rect 699 1052 700 1056
rect 694 1051 700 1052
rect 974 1056 980 1057
rect 974 1052 975 1056
rect 979 1052 980 1056
rect 974 1051 980 1052
rect 1270 1056 1276 1057
rect 1270 1052 1271 1056
rect 1275 1052 1276 1056
rect 1270 1051 1276 1052
rect 110 1050 116 1051
rect 112 1011 114 1050
rect 216 1011 218 1051
rect 440 1011 442 1051
rect 696 1011 698 1051
rect 976 1011 978 1051
rect 1272 1011 1274 1051
rect 111 1010 115 1011
rect 111 1005 115 1006
rect 215 1010 219 1011
rect 215 1005 219 1006
rect 439 1010 443 1011
rect 439 1005 443 1006
rect 511 1010 515 1011
rect 511 1005 515 1006
rect 663 1010 667 1011
rect 663 1005 667 1006
rect 695 1010 699 1011
rect 695 1005 699 1006
rect 831 1010 835 1011
rect 831 1005 835 1006
rect 975 1010 979 1011
rect 975 1005 979 1006
rect 1007 1010 1011 1011
rect 1007 1005 1011 1006
rect 1199 1010 1203 1011
rect 1199 1005 1203 1006
rect 1271 1010 1275 1011
rect 1271 1005 1275 1006
rect 112 982 114 1005
rect 110 981 116 982
rect 512 981 514 1005
rect 664 981 666 1005
rect 832 981 834 1005
rect 1008 981 1010 1005
rect 1200 981 1202 1005
rect 110 977 111 981
rect 115 977 116 981
rect 110 976 116 977
rect 510 980 516 981
rect 510 976 511 980
rect 515 976 516 980
rect 510 975 516 976
rect 662 980 668 981
rect 662 976 663 980
rect 667 976 668 980
rect 662 975 668 976
rect 830 980 836 981
rect 830 976 831 980
rect 835 976 836 980
rect 830 975 836 976
rect 1006 980 1012 981
rect 1006 976 1007 980
rect 1011 976 1012 980
rect 1006 975 1012 976
rect 1198 980 1204 981
rect 1198 976 1199 980
rect 1203 976 1204 980
rect 1198 975 1204 976
rect 486 965 492 966
rect 110 963 116 964
rect 110 959 111 963
rect 115 959 116 963
rect 486 961 487 965
rect 491 961 492 965
rect 486 960 492 961
rect 638 965 644 966
rect 638 961 639 965
rect 643 961 644 965
rect 638 960 644 961
rect 806 965 812 966
rect 806 961 807 965
rect 811 961 812 965
rect 806 960 812 961
rect 982 965 988 966
rect 982 961 983 965
rect 987 961 988 965
rect 982 960 988 961
rect 1174 965 1180 966
rect 1174 961 1175 965
rect 1179 961 1180 965
rect 1174 960 1180 961
rect 110 958 116 959
rect 112 899 114 958
rect 488 899 490 960
rect 586 959 592 960
rect 586 955 587 959
rect 591 955 592 959
rect 586 954 592 955
rect 578 951 584 952
rect 578 947 579 951
rect 583 947 584 951
rect 578 946 584 947
rect 580 916 582 946
rect 588 916 590 954
rect 578 915 584 916
rect 578 911 579 915
rect 583 911 584 915
rect 578 910 584 911
rect 586 915 592 916
rect 586 911 587 915
rect 591 911 592 915
rect 586 910 592 911
rect 640 899 642 960
rect 738 959 744 960
rect 738 955 739 959
rect 743 955 744 959
rect 738 954 744 955
rect 740 916 742 954
rect 738 915 744 916
rect 738 911 739 915
rect 743 911 744 915
rect 738 910 744 911
rect 808 899 810 960
rect 984 899 986 960
rect 1118 959 1124 960
rect 1118 955 1119 959
rect 1123 955 1124 959
rect 1118 954 1124 955
rect 1158 959 1164 960
rect 1158 955 1159 959
rect 1163 955 1164 959
rect 1158 954 1164 955
rect 1120 916 1122 954
rect 1118 915 1124 916
rect 1118 911 1119 915
rect 1123 911 1124 915
rect 1118 910 1124 911
rect 1160 904 1162 954
rect 1158 903 1164 904
rect 1158 899 1159 903
rect 1163 899 1164 903
rect 1176 899 1178 960
rect 1344 952 1346 1072
rect 1399 1010 1403 1011
rect 1399 1005 1403 1006
rect 1400 981 1402 1005
rect 1398 980 1404 981
rect 1398 976 1399 980
rect 1403 976 1404 980
rect 1398 975 1404 976
rect 1374 965 1380 966
rect 1374 961 1375 965
rect 1379 961 1380 965
rect 1374 960 1380 961
rect 1412 960 1414 1126
rect 1527 1121 1531 1122
rect 1543 1126 1547 1127
rect 1614 1126 1620 1127
rect 1624 1124 1626 1170
rect 1720 1127 1722 1174
rect 1719 1126 1723 1127
rect 1543 1121 1547 1122
rect 1622 1123 1628 1124
rect 1544 1072 1546 1121
rect 1622 1119 1623 1123
rect 1627 1119 1628 1123
rect 1719 1121 1723 1122
rect 1622 1118 1628 1119
rect 1638 1077 1644 1078
rect 1638 1073 1639 1077
rect 1643 1073 1644 1077
rect 1720 1074 1722 1121
rect 1638 1072 1644 1073
rect 1718 1073 1724 1074
rect 1542 1071 1548 1072
rect 1542 1067 1543 1071
rect 1547 1067 1548 1071
rect 1542 1066 1548 1067
rect 1566 1056 1572 1057
rect 1566 1052 1567 1056
rect 1571 1052 1572 1056
rect 1566 1051 1572 1052
rect 1568 1011 1570 1051
rect 1567 1010 1571 1011
rect 1567 1005 1571 1006
rect 1599 1010 1603 1011
rect 1599 1005 1603 1006
rect 1600 981 1602 1005
rect 1598 980 1604 981
rect 1598 976 1599 980
rect 1603 976 1604 980
rect 1598 975 1604 976
rect 1574 965 1580 966
rect 1574 961 1575 965
rect 1579 961 1580 965
rect 1574 960 1580 961
rect 1342 951 1348 952
rect 1342 947 1343 951
rect 1347 947 1348 951
rect 1342 946 1348 947
rect 1376 899 1378 960
rect 1410 959 1416 960
rect 1410 955 1411 959
rect 1415 955 1416 959
rect 1410 954 1416 955
rect 1494 911 1500 912
rect 1494 907 1495 911
rect 1499 907 1500 911
rect 1494 906 1500 907
rect 111 898 115 899
rect 111 893 115 894
rect 487 898 491 899
rect 487 893 491 894
rect 639 898 643 899
rect 639 893 643 894
rect 759 898 763 899
rect 759 893 763 894
rect 807 898 811 899
rect 911 898 915 899
rect 807 893 811 894
rect 858 895 864 896
rect 112 846 114 893
rect 110 845 116 846
rect 110 841 111 845
rect 115 841 116 845
rect 760 844 762 893
rect 858 891 859 895
rect 863 891 864 895
rect 911 893 915 894
rect 983 898 987 899
rect 1071 898 1075 899
rect 1158 898 1164 899
rect 1175 898 1179 899
rect 983 893 987 894
rect 1010 895 1016 896
rect 858 890 864 891
rect 860 850 862 890
rect 858 849 864 850
rect 858 845 859 849
rect 863 845 864 849
rect 858 844 864 845
rect 912 844 914 893
rect 1010 891 1011 895
rect 1015 891 1016 895
rect 1071 893 1075 894
rect 1239 898 1243 899
rect 1175 893 1179 894
rect 1182 895 1188 896
rect 1010 890 1016 891
rect 1012 850 1014 890
rect 1010 849 1016 850
rect 1010 845 1011 849
rect 1015 845 1016 849
rect 1010 844 1016 845
rect 1072 844 1074 893
rect 1182 891 1183 895
rect 1187 891 1188 895
rect 1375 898 1379 899
rect 1239 893 1243 894
rect 1338 895 1344 896
rect 1182 890 1188 891
rect 1184 850 1186 890
rect 1182 849 1188 850
rect 1182 845 1183 849
rect 1187 845 1188 849
rect 1182 844 1188 845
rect 1240 844 1242 893
rect 1338 891 1339 895
rect 1343 891 1344 895
rect 1375 893 1379 894
rect 1407 898 1411 899
rect 1407 893 1411 894
rect 1338 890 1344 891
rect 1340 852 1342 890
rect 1338 851 1344 852
rect 1338 847 1339 851
rect 1343 847 1344 851
rect 1338 846 1344 847
rect 1378 851 1384 852
rect 1378 847 1379 851
rect 1383 847 1384 851
rect 1378 846 1384 847
rect 110 840 116 841
rect 758 843 764 844
rect 758 839 759 843
rect 763 839 764 843
rect 758 838 764 839
rect 910 843 916 844
rect 910 839 911 843
rect 915 839 916 843
rect 910 838 916 839
rect 1070 843 1076 844
rect 1070 839 1071 843
rect 1075 839 1076 843
rect 1070 838 1076 839
rect 1238 843 1244 844
rect 1238 839 1239 843
rect 1243 839 1244 843
rect 1238 838 1244 839
rect 782 828 788 829
rect 110 827 116 828
rect 110 823 111 827
rect 115 823 116 827
rect 782 824 783 828
rect 787 824 788 828
rect 782 823 788 824
rect 934 828 940 829
rect 934 824 935 828
rect 939 824 940 828
rect 934 823 940 824
rect 1094 828 1100 829
rect 1094 824 1095 828
rect 1099 824 1100 828
rect 1094 823 1100 824
rect 1262 828 1268 829
rect 1262 824 1263 828
rect 1267 824 1268 828
rect 1262 823 1268 824
rect 110 822 116 823
rect 112 791 114 822
rect 784 791 786 823
rect 936 791 938 823
rect 1096 791 1098 823
rect 1264 791 1266 823
rect 111 790 115 791
rect 111 785 115 786
rect 695 790 699 791
rect 695 785 699 786
rect 783 790 787 791
rect 783 785 787 786
rect 831 790 835 791
rect 831 785 835 786
rect 935 790 939 791
rect 935 785 939 786
rect 975 790 979 791
rect 975 785 979 786
rect 1095 790 1099 791
rect 1095 785 1099 786
rect 1119 790 1123 791
rect 1119 785 1123 786
rect 1263 790 1267 791
rect 1263 785 1267 786
rect 1271 790 1275 791
rect 1271 785 1275 786
rect 112 762 114 785
rect 110 761 116 762
rect 696 761 698 785
rect 832 761 834 785
rect 976 761 978 785
rect 1120 761 1122 785
rect 1272 761 1274 785
rect 110 757 111 761
rect 115 757 116 761
rect 110 756 116 757
rect 694 760 700 761
rect 694 756 695 760
rect 699 756 700 760
rect 694 755 700 756
rect 830 760 836 761
rect 830 756 831 760
rect 835 756 836 760
rect 830 755 836 756
rect 974 760 980 761
rect 974 756 975 760
rect 979 756 980 760
rect 974 755 980 756
rect 1118 760 1124 761
rect 1118 756 1119 760
rect 1123 756 1124 760
rect 1118 755 1124 756
rect 1270 760 1276 761
rect 1270 756 1271 760
rect 1275 756 1276 760
rect 1270 755 1276 756
rect 670 745 676 746
rect 110 743 116 744
rect 110 739 111 743
rect 115 739 116 743
rect 670 741 671 745
rect 675 741 676 745
rect 670 740 676 741
rect 806 745 812 746
rect 806 741 807 745
rect 811 741 812 745
rect 806 740 812 741
rect 950 745 956 746
rect 950 741 951 745
rect 955 741 956 745
rect 950 740 956 741
rect 1094 745 1100 746
rect 1094 741 1095 745
rect 1099 741 1100 745
rect 1094 740 1100 741
rect 1246 745 1252 746
rect 1246 741 1247 745
rect 1251 741 1252 745
rect 1246 740 1252 741
rect 110 738 116 739
rect 112 667 114 738
rect 672 667 674 740
rect 790 739 796 740
rect 790 735 791 739
rect 795 735 796 739
rect 790 734 796 735
rect 762 731 768 732
rect 762 727 763 731
rect 767 727 768 731
rect 762 726 768 727
rect 764 696 766 726
rect 792 696 794 734
rect 762 695 768 696
rect 762 691 763 695
rect 767 691 768 695
rect 762 690 768 691
rect 790 695 796 696
rect 790 691 791 695
rect 795 691 796 695
rect 790 690 796 691
rect 808 667 810 740
rect 952 667 954 740
rect 1050 739 1056 740
rect 1050 735 1051 739
rect 1055 735 1056 739
rect 1050 734 1056 735
rect 111 666 115 667
rect 111 661 115 662
rect 247 666 251 667
rect 247 661 251 662
rect 431 666 435 667
rect 631 666 635 667
rect 431 661 435 662
rect 622 663 628 664
rect 112 614 114 661
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 248 612 250 661
rect 258 619 264 620
rect 258 615 259 619
rect 263 615 264 619
rect 258 614 264 615
rect 110 608 116 609
rect 246 611 252 612
rect 246 607 247 611
rect 251 607 252 611
rect 246 606 252 607
rect 110 595 116 596
rect 110 591 111 595
rect 115 591 116 595
rect 110 590 116 591
rect 112 551 114 590
rect 111 550 115 551
rect 111 545 115 546
rect 159 550 163 551
rect 159 545 163 546
rect 112 522 114 545
rect 110 521 116 522
rect 160 521 162 545
rect 110 517 111 521
rect 115 517 116 521
rect 110 516 116 517
rect 158 520 164 521
rect 158 516 159 520
rect 163 516 164 520
rect 158 515 164 516
rect 134 505 140 506
rect 110 503 116 504
rect 110 499 111 503
rect 115 499 116 503
rect 134 501 135 505
rect 139 501 140 505
rect 134 500 140 501
rect 110 498 116 499
rect 112 439 114 498
rect 136 439 138 500
rect 260 467 262 614
rect 432 612 434 661
rect 622 659 623 663
rect 627 659 628 663
rect 631 661 635 662
rect 671 666 675 667
rect 671 661 675 662
rect 807 666 811 667
rect 847 666 851 667
rect 807 661 811 662
rect 838 663 844 664
rect 622 658 628 659
rect 624 620 626 658
rect 622 619 628 620
rect 622 615 623 619
rect 627 615 628 619
rect 622 614 628 615
rect 632 612 634 661
rect 838 659 839 663
rect 843 659 844 663
rect 847 661 851 662
rect 951 666 955 667
rect 1052 664 1054 734
rect 1096 667 1098 740
rect 1218 739 1224 740
rect 1218 735 1219 739
rect 1223 735 1224 739
rect 1218 734 1224 735
rect 1220 696 1222 734
rect 1218 695 1224 696
rect 1218 691 1219 695
rect 1223 691 1224 695
rect 1218 690 1224 691
rect 1248 667 1250 740
rect 1380 696 1382 846
rect 1408 844 1410 893
rect 1406 843 1412 844
rect 1406 839 1407 843
rect 1411 839 1412 843
rect 1406 838 1412 839
rect 1430 828 1436 829
rect 1430 824 1431 828
rect 1435 824 1436 828
rect 1430 823 1436 824
rect 1432 791 1434 823
rect 1431 790 1435 791
rect 1431 785 1435 786
rect 1432 761 1434 785
rect 1430 760 1436 761
rect 1430 756 1431 760
rect 1435 756 1436 760
rect 1430 755 1436 756
rect 1406 745 1412 746
rect 1406 741 1407 745
rect 1411 741 1412 745
rect 1406 740 1412 741
rect 1496 740 1498 906
rect 1576 899 1578 960
rect 1640 916 1642 1072
rect 1718 1069 1719 1073
rect 1723 1069 1724 1073
rect 1718 1068 1724 1069
rect 1718 1055 1724 1056
rect 1718 1051 1719 1055
rect 1723 1051 1724 1055
rect 1718 1050 1724 1051
rect 1720 1011 1722 1050
rect 1719 1010 1723 1011
rect 1719 1005 1723 1006
rect 1720 982 1722 1005
rect 1718 981 1724 982
rect 1718 977 1719 981
rect 1723 977 1724 981
rect 1718 976 1724 977
rect 1718 963 1724 964
rect 1666 959 1672 960
rect 1666 955 1667 959
rect 1671 955 1672 959
rect 1718 959 1719 963
rect 1723 959 1724 963
rect 1718 958 1724 959
rect 1666 954 1672 955
rect 1638 915 1644 916
rect 1638 911 1639 915
rect 1643 911 1644 915
rect 1638 910 1644 911
rect 1575 898 1579 899
rect 1668 896 1670 954
rect 1720 899 1722 958
rect 1719 898 1723 899
rect 1575 893 1579 894
rect 1666 895 1672 896
rect 1576 844 1578 893
rect 1666 891 1667 895
rect 1671 891 1672 895
rect 1719 893 1723 894
rect 1666 890 1672 891
rect 1666 849 1672 850
rect 1666 845 1667 849
rect 1671 845 1672 849
rect 1720 846 1722 893
rect 1666 844 1672 845
rect 1718 845 1724 846
rect 1574 843 1580 844
rect 1574 839 1575 843
rect 1579 839 1580 843
rect 1574 838 1580 839
rect 1598 828 1604 829
rect 1598 824 1599 828
rect 1603 824 1604 828
rect 1598 823 1604 824
rect 1600 791 1602 823
rect 1599 790 1603 791
rect 1599 785 1603 786
rect 1600 761 1602 785
rect 1598 760 1604 761
rect 1598 756 1599 760
rect 1603 756 1604 760
rect 1598 755 1604 756
rect 1574 745 1580 746
rect 1574 741 1575 745
rect 1579 741 1580 745
rect 1574 740 1580 741
rect 1378 695 1384 696
rect 1378 691 1379 695
rect 1383 691 1384 695
rect 1378 690 1384 691
rect 1408 667 1410 740
rect 1494 739 1500 740
rect 1494 735 1495 739
rect 1499 735 1500 739
rect 1494 734 1500 735
rect 1414 695 1420 696
rect 1414 691 1415 695
rect 1419 691 1420 695
rect 1414 690 1420 691
rect 1079 666 1083 667
rect 951 661 955 662
rect 1042 663 1048 664
rect 838 658 844 659
rect 840 620 842 658
rect 838 619 844 620
rect 838 615 839 619
rect 843 615 844 619
rect 838 614 844 615
rect 848 612 850 661
rect 1042 659 1043 663
rect 1047 659 1048 663
rect 1042 658 1048 659
rect 1050 663 1056 664
rect 1050 659 1051 663
rect 1055 659 1056 663
rect 1079 661 1083 662
rect 1095 666 1099 667
rect 1095 661 1099 662
rect 1247 666 1251 667
rect 1247 661 1251 662
rect 1319 666 1323 667
rect 1319 661 1323 662
rect 1407 666 1411 667
rect 1407 661 1411 662
rect 1050 658 1056 659
rect 1044 620 1046 658
rect 1042 619 1048 620
rect 1042 615 1043 619
rect 1047 615 1048 619
rect 1042 614 1048 615
rect 1080 612 1082 661
rect 1320 612 1322 661
rect 1416 618 1418 690
rect 1576 667 1578 740
rect 1650 739 1656 740
rect 1650 735 1651 739
rect 1655 735 1656 739
rect 1650 734 1656 735
rect 1559 666 1563 667
rect 1434 663 1440 664
rect 1434 659 1435 663
rect 1439 659 1440 663
rect 1559 661 1563 662
rect 1575 666 1579 667
rect 1652 664 1654 734
rect 1668 696 1670 844
rect 1718 841 1719 845
rect 1723 841 1724 845
rect 1718 840 1724 841
rect 1718 827 1724 828
rect 1718 823 1719 827
rect 1723 823 1724 827
rect 1718 822 1724 823
rect 1720 791 1722 822
rect 1719 790 1723 791
rect 1719 785 1723 786
rect 1720 762 1722 785
rect 1718 761 1724 762
rect 1718 757 1719 761
rect 1723 757 1724 761
rect 1718 756 1724 757
rect 1718 743 1724 744
rect 1718 739 1719 743
rect 1723 739 1724 743
rect 1718 738 1724 739
rect 1666 695 1672 696
rect 1666 691 1667 695
rect 1671 691 1672 695
rect 1666 690 1672 691
rect 1720 667 1722 738
rect 1719 666 1723 667
rect 1575 661 1579 662
rect 1650 663 1656 664
rect 1434 658 1440 659
rect 1414 617 1420 618
rect 1414 613 1415 617
rect 1419 613 1420 617
rect 1414 612 1420 613
rect 430 611 436 612
rect 430 607 431 611
rect 435 607 436 611
rect 430 606 436 607
rect 630 611 636 612
rect 630 607 631 611
rect 635 607 636 611
rect 630 606 636 607
rect 846 611 852 612
rect 846 607 847 611
rect 851 607 852 611
rect 846 606 852 607
rect 1078 611 1084 612
rect 1078 607 1079 611
rect 1083 607 1084 611
rect 1078 606 1084 607
rect 1318 611 1324 612
rect 1318 607 1319 611
rect 1323 607 1324 611
rect 1318 606 1324 607
rect 270 596 276 597
rect 270 592 271 596
rect 275 592 276 596
rect 270 591 276 592
rect 454 596 460 597
rect 454 592 455 596
rect 459 592 460 596
rect 454 591 460 592
rect 654 596 660 597
rect 654 592 655 596
rect 659 592 660 596
rect 654 591 660 592
rect 870 596 876 597
rect 870 592 871 596
rect 875 592 876 596
rect 870 591 876 592
rect 1102 596 1108 597
rect 1102 592 1103 596
rect 1107 592 1108 596
rect 1102 591 1108 592
rect 1342 596 1348 597
rect 1342 592 1343 596
rect 1347 592 1348 596
rect 1342 591 1348 592
rect 272 551 274 591
rect 456 551 458 591
rect 656 551 658 591
rect 872 551 874 591
rect 1104 551 1106 591
rect 1344 551 1346 591
rect 271 550 275 551
rect 271 545 275 546
rect 343 550 347 551
rect 343 545 347 546
rect 455 550 459 551
rect 455 545 459 546
rect 575 550 579 551
rect 575 545 579 546
rect 655 550 659 551
rect 655 545 659 546
rect 831 550 835 551
rect 831 545 835 546
rect 871 550 875 551
rect 871 545 875 546
rect 1095 550 1099 551
rect 1095 545 1099 546
rect 1103 550 1107 551
rect 1103 545 1107 546
rect 1343 550 1347 551
rect 1343 545 1347 546
rect 1367 550 1371 551
rect 1367 545 1371 546
rect 344 521 346 545
rect 576 521 578 545
rect 832 521 834 545
rect 1096 521 1098 545
rect 1368 521 1370 545
rect 342 520 348 521
rect 342 516 343 520
rect 347 516 348 520
rect 342 515 348 516
rect 574 520 580 521
rect 574 516 575 520
rect 579 516 580 520
rect 574 515 580 516
rect 830 520 836 521
rect 830 516 831 520
rect 835 516 836 520
rect 830 515 836 516
rect 1094 520 1100 521
rect 1094 516 1095 520
rect 1099 516 1100 520
rect 1094 515 1100 516
rect 1366 520 1372 521
rect 1366 516 1367 520
rect 1371 516 1372 520
rect 1366 515 1372 516
rect 318 505 324 506
rect 318 501 319 505
rect 323 501 324 505
rect 318 500 324 501
rect 550 505 556 506
rect 550 501 551 505
rect 555 501 556 505
rect 550 500 556 501
rect 806 505 812 506
rect 806 501 807 505
rect 811 501 812 505
rect 806 500 812 501
rect 1070 505 1076 506
rect 1070 501 1071 505
rect 1075 501 1076 505
rect 1070 500 1076 501
rect 1342 505 1348 506
rect 1342 501 1343 505
rect 1347 501 1348 505
rect 1342 500 1348 501
rect 1436 500 1438 658
rect 1560 612 1562 661
rect 1650 659 1651 663
rect 1655 659 1656 663
rect 1719 661 1723 662
rect 1650 658 1656 659
rect 1654 617 1660 618
rect 1654 613 1655 617
rect 1659 613 1660 617
rect 1720 614 1722 661
rect 1654 612 1660 613
rect 1718 613 1724 614
rect 1558 611 1564 612
rect 1558 607 1559 611
rect 1563 607 1564 611
rect 1558 606 1564 607
rect 1582 596 1588 597
rect 1582 592 1583 596
rect 1587 592 1588 596
rect 1582 591 1588 592
rect 1584 551 1586 591
rect 1583 550 1587 551
rect 1583 545 1587 546
rect 290 491 296 492
rect 290 487 291 491
rect 295 487 296 491
rect 290 486 296 487
rect 256 465 262 467
rect 256 456 258 465
rect 254 455 260 456
rect 254 451 255 455
rect 259 451 260 455
rect 254 450 260 451
rect 111 438 115 439
rect 111 433 115 434
rect 135 438 139 439
rect 135 433 139 434
rect 199 438 203 439
rect 292 436 294 486
rect 320 439 322 500
rect 418 499 424 500
rect 418 495 419 499
rect 423 495 424 499
rect 418 494 424 495
rect 420 456 422 494
rect 418 455 424 456
rect 418 451 419 455
rect 423 451 424 455
rect 418 450 424 451
rect 552 439 554 500
rect 650 499 656 500
rect 650 495 651 499
rect 655 495 656 499
rect 650 494 656 495
rect 652 456 654 494
rect 650 455 656 456
rect 650 451 651 455
rect 655 451 656 455
rect 650 450 656 451
rect 808 439 810 500
rect 1072 439 1074 500
rect 1344 439 1346 500
rect 1434 499 1440 500
rect 1434 495 1435 499
rect 1439 495 1440 499
rect 1434 494 1440 495
rect 1422 455 1428 456
rect 1422 451 1423 455
rect 1427 451 1428 455
rect 1422 450 1428 451
rect 319 438 323 439
rect 199 433 203 434
rect 290 435 296 436
rect 112 386 114 433
rect 110 385 116 386
rect 110 381 111 385
rect 115 381 116 385
rect 200 384 202 433
rect 290 431 291 435
rect 295 431 296 435
rect 290 430 296 431
rect 298 435 304 436
rect 298 431 299 435
rect 303 431 304 435
rect 319 433 323 434
rect 415 438 419 439
rect 551 438 555 439
rect 415 433 419 434
rect 530 435 536 436
rect 298 430 304 431
rect 300 390 302 430
rect 298 389 304 390
rect 298 385 299 389
rect 303 385 304 389
rect 298 384 304 385
rect 416 384 418 433
rect 530 431 531 435
rect 535 431 536 435
rect 551 433 555 434
rect 631 438 635 439
rect 807 438 811 439
rect 631 433 635 434
rect 730 435 736 436
rect 530 430 536 431
rect 532 390 534 430
rect 530 389 536 390
rect 530 385 531 389
rect 535 385 536 389
rect 530 384 536 385
rect 632 384 634 433
rect 730 431 731 435
rect 735 431 736 435
rect 807 433 811 434
rect 855 438 859 439
rect 855 433 859 434
rect 1071 438 1075 439
rect 1071 433 1075 434
rect 1087 438 1091 439
rect 1327 438 1331 439
rect 1087 433 1091 434
rect 1174 435 1180 436
rect 730 430 736 431
rect 732 390 734 430
rect 730 389 736 390
rect 730 385 731 389
rect 735 385 736 389
rect 730 384 736 385
rect 856 384 858 433
rect 950 389 956 390
rect 950 385 951 389
rect 955 385 956 389
rect 950 384 956 385
rect 1088 384 1090 433
rect 1174 431 1175 435
rect 1179 431 1180 435
rect 1174 430 1180 431
rect 1186 435 1192 436
rect 1186 431 1187 435
rect 1191 431 1192 435
rect 1327 433 1331 434
rect 1343 438 1347 439
rect 1343 433 1347 434
rect 1186 430 1192 431
rect 110 380 116 381
rect 198 383 204 384
rect 198 379 199 383
rect 203 379 204 383
rect 198 378 204 379
rect 414 383 420 384
rect 414 379 415 383
rect 419 379 420 383
rect 414 378 420 379
rect 630 383 636 384
rect 630 379 631 383
rect 635 379 636 383
rect 630 378 636 379
rect 854 383 860 384
rect 854 379 855 383
rect 859 379 860 383
rect 854 378 860 379
rect 222 368 228 369
rect 110 367 116 368
rect 110 363 111 367
rect 115 363 116 367
rect 222 364 223 368
rect 227 364 228 368
rect 222 363 228 364
rect 438 368 444 369
rect 438 364 439 368
rect 443 364 444 368
rect 438 363 444 364
rect 654 368 660 369
rect 654 364 655 368
rect 659 364 660 368
rect 654 363 660 364
rect 878 368 884 369
rect 878 364 879 368
rect 883 364 884 368
rect 878 363 884 364
rect 110 362 116 363
rect 112 335 114 362
rect 224 335 226 363
rect 440 335 442 363
rect 656 335 658 363
rect 880 335 882 363
rect 111 334 115 335
rect 111 329 115 330
rect 223 334 227 335
rect 223 329 227 330
rect 439 334 443 335
rect 439 329 443 330
rect 559 334 563 335
rect 559 329 563 330
rect 655 334 659 335
rect 655 329 659 330
rect 759 334 763 335
rect 759 329 763 330
rect 879 334 883 335
rect 879 329 883 330
rect 112 306 114 329
rect 110 305 116 306
rect 560 305 562 329
rect 760 305 762 329
rect 110 301 111 305
rect 115 301 116 305
rect 110 300 116 301
rect 558 304 564 305
rect 558 300 559 304
rect 563 300 564 304
rect 558 299 564 300
rect 758 304 764 305
rect 758 300 759 304
rect 763 300 764 304
rect 758 299 764 300
rect 534 289 540 290
rect 110 287 116 288
rect 110 283 111 287
rect 115 283 116 287
rect 534 285 535 289
rect 539 285 540 289
rect 534 284 540 285
rect 734 289 740 290
rect 734 285 735 289
rect 739 285 740 289
rect 734 284 740 285
rect 942 289 948 290
rect 942 285 943 289
rect 947 285 948 289
rect 942 284 948 285
rect 110 282 116 283
rect 112 223 114 282
rect 536 223 538 284
rect 578 283 584 284
rect 578 279 579 283
rect 583 279 584 283
rect 578 278 584 279
rect 654 283 660 284
rect 654 279 655 283
rect 659 279 660 283
rect 654 278 660 279
rect 111 222 115 223
rect 111 217 115 218
rect 487 222 491 223
rect 487 217 491 218
rect 535 222 539 223
rect 580 220 582 278
rect 656 240 658 278
rect 654 239 660 240
rect 654 235 655 239
rect 659 235 660 239
rect 654 234 660 235
rect 736 223 738 284
rect 886 283 892 284
rect 886 279 887 283
rect 891 279 892 283
rect 886 278 892 279
rect 888 240 890 278
rect 886 239 892 240
rect 886 235 887 239
rect 891 235 892 239
rect 886 234 892 235
rect 944 223 946 284
rect 952 240 954 384
rect 1086 383 1092 384
rect 1086 379 1087 383
rect 1091 379 1092 383
rect 1086 378 1092 379
rect 1110 368 1116 369
rect 1110 364 1111 368
rect 1115 364 1116 368
rect 1110 363 1116 364
rect 1112 335 1114 363
rect 967 334 971 335
rect 967 329 971 330
rect 1111 334 1115 335
rect 1111 329 1115 330
rect 968 305 970 329
rect 966 304 972 305
rect 966 300 967 304
rect 971 300 972 304
rect 966 299 972 300
rect 1158 289 1164 290
rect 1158 285 1159 289
rect 1163 285 1164 289
rect 1158 284 1164 285
rect 1176 284 1178 430
rect 1188 390 1190 430
rect 1186 389 1192 390
rect 1186 385 1187 389
rect 1191 385 1192 389
rect 1186 384 1192 385
rect 1328 384 1330 433
rect 1424 390 1426 450
rect 1575 438 1579 439
rect 1656 436 1658 612
rect 1718 609 1719 613
rect 1723 609 1724 613
rect 1718 608 1724 609
rect 1718 595 1724 596
rect 1718 591 1719 595
rect 1723 591 1724 595
rect 1718 590 1724 591
rect 1720 551 1722 590
rect 1719 550 1723 551
rect 1719 545 1723 546
rect 1720 522 1722 545
rect 1718 521 1724 522
rect 1718 517 1719 521
rect 1723 517 1724 521
rect 1718 516 1724 517
rect 1718 503 1724 504
rect 1718 499 1719 503
rect 1723 499 1724 503
rect 1718 498 1724 499
rect 1720 439 1722 498
rect 1719 438 1723 439
rect 1575 433 1579 434
rect 1654 435 1660 436
rect 1422 389 1428 390
rect 1422 385 1423 389
rect 1427 385 1428 389
rect 1422 384 1428 385
rect 1576 384 1578 433
rect 1654 431 1655 435
rect 1659 431 1660 435
rect 1719 433 1723 434
rect 1654 430 1660 431
rect 1674 389 1680 390
rect 1674 385 1675 389
rect 1679 385 1680 389
rect 1720 386 1722 433
rect 1674 384 1680 385
rect 1718 385 1724 386
rect 1326 383 1332 384
rect 1326 379 1327 383
rect 1331 379 1332 383
rect 1326 378 1332 379
rect 1574 383 1580 384
rect 1574 379 1575 383
rect 1579 379 1580 383
rect 1574 378 1580 379
rect 1350 368 1356 369
rect 1350 364 1351 368
rect 1355 364 1356 368
rect 1350 363 1356 364
rect 1598 368 1604 369
rect 1598 364 1599 368
rect 1603 364 1604 368
rect 1598 363 1604 364
rect 1352 335 1354 363
rect 1600 335 1602 363
rect 1183 334 1187 335
rect 1183 329 1187 330
rect 1351 334 1355 335
rect 1351 329 1355 330
rect 1399 334 1403 335
rect 1399 329 1403 330
rect 1599 334 1603 335
rect 1599 329 1603 330
rect 1184 305 1186 329
rect 1400 305 1402 329
rect 1600 305 1602 329
rect 1182 304 1188 305
rect 1182 300 1183 304
rect 1187 300 1188 304
rect 1182 299 1188 300
rect 1398 304 1404 305
rect 1398 300 1399 304
rect 1403 300 1404 304
rect 1398 299 1404 300
rect 1598 304 1604 305
rect 1598 300 1599 304
rect 1603 300 1604 304
rect 1598 299 1604 300
rect 1374 289 1380 290
rect 1374 285 1375 289
rect 1379 285 1380 289
rect 1374 284 1380 285
rect 1574 289 1580 290
rect 1574 285 1575 289
rect 1579 285 1580 289
rect 1574 284 1580 285
rect 950 239 956 240
rect 950 235 951 239
rect 955 235 956 239
rect 950 234 956 235
rect 1160 223 1162 284
rect 1174 283 1180 284
rect 1174 279 1175 283
rect 1179 279 1180 283
rect 1174 278 1180 279
rect 1314 283 1320 284
rect 1314 279 1315 283
rect 1319 279 1320 283
rect 1314 278 1320 279
rect 1316 240 1318 278
rect 1314 239 1320 240
rect 1314 235 1315 239
rect 1319 235 1320 239
rect 1314 234 1320 235
rect 1376 223 1378 284
rect 1398 239 1404 240
rect 1398 235 1399 239
rect 1403 235 1404 239
rect 1398 234 1404 235
rect 623 222 627 223
rect 535 217 539 218
rect 578 219 584 220
rect 112 170 114 217
rect 110 169 116 170
rect 110 165 111 169
rect 115 165 116 169
rect 488 168 490 217
rect 578 215 579 219
rect 583 215 584 219
rect 578 214 584 215
rect 586 219 592 220
rect 586 215 587 219
rect 591 215 592 219
rect 735 222 739 223
rect 623 217 627 218
rect 722 219 728 220
rect 586 214 592 215
rect 588 174 590 214
rect 586 173 592 174
rect 586 169 587 173
rect 591 169 592 173
rect 586 168 592 169
rect 624 168 626 217
rect 722 215 723 219
rect 727 215 728 219
rect 735 217 739 218
rect 759 222 763 223
rect 895 222 899 223
rect 759 217 763 218
rect 874 219 880 220
rect 722 214 728 215
rect 724 174 726 214
rect 722 173 728 174
rect 722 169 723 173
rect 727 169 728 173
rect 722 168 728 169
rect 760 168 762 217
rect 874 215 875 219
rect 879 215 880 219
rect 895 217 899 218
rect 943 222 947 223
rect 1031 222 1035 223
rect 943 217 947 218
rect 1010 219 1016 220
rect 874 214 880 215
rect 876 174 878 214
rect 874 173 880 174
rect 874 169 875 173
rect 879 169 880 173
rect 874 168 880 169
rect 896 168 898 217
rect 1010 215 1011 219
rect 1015 215 1016 219
rect 1159 222 1163 223
rect 1031 217 1035 218
rect 1130 219 1136 220
rect 1010 214 1016 215
rect 1012 174 1014 214
rect 1010 173 1016 174
rect 1010 169 1011 173
rect 1015 169 1016 173
rect 1010 168 1016 169
rect 1032 168 1034 217
rect 1130 215 1131 219
rect 1135 215 1136 219
rect 1159 217 1163 218
rect 1167 222 1171 223
rect 1303 222 1307 223
rect 1167 217 1171 218
rect 1282 219 1288 220
rect 1130 214 1136 215
rect 1132 174 1134 214
rect 1130 173 1136 174
rect 1130 169 1131 173
rect 1135 169 1136 173
rect 1130 168 1136 169
rect 1168 168 1170 217
rect 1282 215 1283 219
rect 1287 215 1288 219
rect 1303 217 1307 218
rect 1375 222 1379 223
rect 1375 217 1379 218
rect 1282 214 1288 215
rect 1284 174 1286 214
rect 1282 173 1288 174
rect 1282 169 1283 173
rect 1287 169 1288 173
rect 1282 168 1288 169
rect 1304 168 1306 217
rect 1400 174 1402 234
rect 1576 223 1578 284
rect 1666 283 1672 284
rect 1666 279 1667 283
rect 1671 279 1672 283
rect 1666 278 1672 279
rect 1439 222 1443 223
rect 1439 217 1443 218
rect 1575 222 1579 223
rect 1668 220 1670 278
rect 1676 240 1678 384
rect 1718 381 1719 385
rect 1723 381 1724 385
rect 1718 380 1724 381
rect 1718 367 1724 368
rect 1718 363 1719 367
rect 1723 363 1724 367
rect 1718 362 1724 363
rect 1720 335 1722 362
rect 1719 334 1723 335
rect 1719 329 1723 330
rect 1720 306 1722 329
rect 1718 305 1724 306
rect 1718 301 1719 305
rect 1723 301 1724 305
rect 1718 300 1724 301
rect 1718 287 1724 288
rect 1718 283 1719 287
rect 1723 283 1724 287
rect 1718 282 1724 283
rect 1674 239 1680 240
rect 1674 235 1675 239
rect 1679 235 1680 239
rect 1674 234 1680 235
rect 1720 223 1722 282
rect 1719 222 1723 223
rect 1575 217 1579 218
rect 1666 219 1672 220
rect 1398 173 1404 174
rect 1398 169 1399 173
rect 1403 169 1404 173
rect 1398 168 1404 169
rect 1440 168 1442 217
rect 1530 215 1536 216
rect 1530 211 1531 215
rect 1535 211 1536 215
rect 1530 210 1536 211
rect 1532 176 1534 210
rect 1530 175 1536 176
rect 1530 171 1531 175
rect 1535 171 1536 175
rect 1530 170 1536 171
rect 1576 168 1578 217
rect 1666 215 1667 219
rect 1671 215 1672 219
rect 1719 217 1723 218
rect 1666 214 1672 215
rect 1720 170 1722 217
rect 1718 169 1724 170
rect 110 164 116 165
rect 486 167 492 168
rect 486 163 487 167
rect 491 163 492 167
rect 486 162 492 163
rect 622 167 628 168
rect 622 163 623 167
rect 627 163 628 167
rect 622 162 628 163
rect 758 167 764 168
rect 758 163 759 167
rect 763 163 764 167
rect 758 162 764 163
rect 894 167 900 168
rect 894 163 895 167
rect 899 163 900 167
rect 894 162 900 163
rect 1030 167 1036 168
rect 1030 163 1031 167
rect 1035 163 1036 167
rect 1030 162 1036 163
rect 1166 167 1172 168
rect 1166 163 1167 167
rect 1171 163 1172 167
rect 1166 162 1172 163
rect 1302 167 1308 168
rect 1302 163 1303 167
rect 1307 163 1308 167
rect 1302 162 1308 163
rect 1438 167 1444 168
rect 1438 163 1439 167
rect 1443 163 1444 167
rect 1438 162 1444 163
rect 1574 167 1580 168
rect 1574 163 1575 167
rect 1579 163 1580 167
rect 1718 165 1719 169
rect 1723 165 1724 169
rect 1718 164 1724 165
rect 1574 162 1580 163
rect 510 152 516 153
rect 110 151 116 152
rect 110 147 111 151
rect 115 147 116 151
rect 510 148 511 152
rect 515 148 516 152
rect 510 147 516 148
rect 646 152 652 153
rect 646 148 647 152
rect 651 148 652 152
rect 646 147 652 148
rect 782 152 788 153
rect 782 148 783 152
rect 787 148 788 152
rect 782 147 788 148
rect 918 152 924 153
rect 918 148 919 152
rect 923 148 924 152
rect 918 147 924 148
rect 1054 152 1060 153
rect 1054 148 1055 152
rect 1059 148 1060 152
rect 1054 147 1060 148
rect 1190 152 1196 153
rect 1190 148 1191 152
rect 1195 148 1196 152
rect 1190 147 1196 148
rect 1326 152 1332 153
rect 1326 148 1327 152
rect 1331 148 1332 152
rect 1326 147 1332 148
rect 1462 152 1468 153
rect 1462 148 1463 152
rect 1467 148 1468 152
rect 1462 147 1468 148
rect 1598 152 1604 153
rect 1598 148 1599 152
rect 1603 148 1604 152
rect 1598 147 1604 148
rect 1718 151 1724 152
rect 1718 147 1719 151
rect 1723 147 1724 151
rect 110 146 116 147
rect 112 123 114 146
rect 512 123 514 147
rect 648 123 650 147
rect 784 123 786 147
rect 920 123 922 147
rect 1056 123 1058 147
rect 1192 123 1194 147
rect 1328 123 1330 147
rect 1464 123 1466 147
rect 1600 123 1602 147
rect 1718 146 1724 147
rect 1720 123 1722 146
rect 111 122 115 123
rect 111 117 115 118
rect 511 122 515 123
rect 511 117 515 118
rect 647 122 651 123
rect 647 117 651 118
rect 783 122 787 123
rect 783 117 787 118
rect 919 122 923 123
rect 919 117 923 118
rect 1055 122 1059 123
rect 1055 117 1059 118
rect 1191 122 1195 123
rect 1191 117 1195 118
rect 1327 122 1331 123
rect 1327 117 1331 118
rect 1463 122 1467 123
rect 1463 117 1467 118
rect 1599 122 1603 123
rect 1599 117 1603 118
rect 1719 122 1723 123
rect 1719 117 1723 118
<< m4c >>
rect 111 1778 115 1782
rect 135 1778 139 1782
rect 271 1778 275 1782
rect 407 1778 411 1782
rect 543 1778 547 1782
rect 679 1778 683 1782
rect 1719 1778 1723 1782
rect 111 1670 115 1674
rect 159 1670 163 1674
rect 239 1670 243 1674
rect 295 1670 299 1674
rect 375 1670 379 1674
rect 431 1670 435 1674
rect 511 1670 515 1674
rect 567 1670 571 1674
rect 647 1670 651 1674
rect 703 1670 707 1674
rect 783 1670 787 1674
rect 1719 1670 1723 1674
rect 111 1554 115 1558
rect 215 1554 219 1558
rect 351 1554 355 1558
rect 487 1554 491 1558
rect 599 1554 603 1558
rect 623 1554 627 1558
rect 735 1554 739 1558
rect 759 1554 763 1558
rect 871 1554 875 1558
rect 1015 1554 1019 1558
rect 1159 1554 1163 1558
rect 1303 1554 1307 1558
rect 1439 1554 1443 1558
rect 111 1450 115 1454
rect 599 1450 603 1454
rect 623 1450 627 1454
rect 735 1450 739 1454
rect 759 1450 763 1454
rect 879 1450 883 1454
rect 895 1450 899 1454
rect 1023 1450 1027 1454
rect 1039 1450 1043 1454
rect 1167 1450 1171 1454
rect 1183 1450 1187 1454
rect 111 1334 115 1338
rect 135 1334 139 1338
rect 303 1334 307 1338
rect 519 1334 523 1338
rect 575 1334 579 1338
rect 711 1334 715 1338
rect 751 1334 755 1338
rect 855 1334 859 1338
rect 1319 1450 1323 1454
rect 1327 1450 1331 1454
rect 1575 1554 1579 1558
rect 1719 1554 1723 1558
rect 1463 1450 1467 1454
rect 1599 1450 1603 1454
rect 999 1334 1003 1338
rect 1143 1334 1147 1338
rect 1255 1334 1259 1338
rect 1295 1334 1299 1338
rect 111 1222 115 1226
rect 159 1222 163 1226
rect 327 1222 331 1226
rect 399 1222 403 1226
rect 543 1222 547 1226
rect 671 1222 675 1226
rect 775 1222 779 1226
rect 959 1222 963 1226
rect 1023 1222 1027 1226
rect 1255 1222 1259 1226
rect 1279 1222 1283 1226
rect 1439 1334 1443 1338
rect 1519 1334 1523 1338
rect 1719 1450 1723 1454
rect 1575 1334 1579 1338
rect 1719 1334 1723 1338
rect 1543 1222 1547 1226
rect 1551 1222 1555 1226
rect 111 1122 115 1126
rect 135 1122 139 1126
rect 191 1122 195 1126
rect 1719 1222 1723 1226
rect 375 1122 379 1126
rect 415 1122 419 1126
rect 647 1122 651 1126
rect 671 1122 675 1126
rect 935 1122 939 1126
rect 951 1122 955 1126
rect 1231 1122 1235 1126
rect 1247 1122 1251 1126
rect 111 1006 115 1010
rect 215 1006 219 1010
rect 439 1006 443 1010
rect 511 1006 515 1010
rect 663 1006 667 1010
rect 695 1006 699 1010
rect 831 1006 835 1010
rect 975 1006 979 1010
rect 1007 1006 1011 1010
rect 1199 1006 1203 1010
rect 1271 1006 1275 1010
rect 1399 1006 1403 1010
rect 1527 1122 1531 1126
rect 1543 1122 1547 1126
rect 1719 1122 1723 1126
rect 1567 1006 1571 1010
rect 1599 1006 1603 1010
rect 111 894 115 898
rect 487 894 491 898
rect 639 894 643 898
rect 759 894 763 898
rect 807 894 811 898
rect 911 894 915 898
rect 983 894 987 898
rect 1071 894 1075 898
rect 1175 894 1179 898
rect 1239 894 1243 898
rect 1375 894 1379 898
rect 1407 894 1411 898
rect 111 786 115 790
rect 695 786 699 790
rect 783 786 787 790
rect 831 786 835 790
rect 935 786 939 790
rect 975 786 979 790
rect 1095 786 1099 790
rect 1119 786 1123 790
rect 1263 786 1267 790
rect 1271 786 1275 790
rect 111 662 115 666
rect 247 662 251 666
rect 431 662 435 666
rect 111 546 115 550
rect 159 546 163 550
rect 631 662 635 666
rect 671 662 675 666
rect 807 662 811 666
rect 847 662 851 666
rect 951 662 955 666
rect 1431 786 1435 790
rect 1719 1006 1723 1010
rect 1575 894 1579 898
rect 1719 894 1723 898
rect 1599 786 1603 790
rect 1079 662 1083 666
rect 1095 662 1099 666
rect 1247 662 1251 666
rect 1319 662 1323 666
rect 1407 662 1411 666
rect 1559 662 1563 666
rect 1575 662 1579 666
rect 1719 786 1723 790
rect 271 546 275 550
rect 343 546 347 550
rect 455 546 459 550
rect 575 546 579 550
rect 655 546 659 550
rect 831 546 835 550
rect 871 546 875 550
rect 1095 546 1099 550
rect 1103 546 1107 550
rect 1343 546 1347 550
rect 1367 546 1371 550
rect 1719 662 1723 666
rect 1583 546 1587 550
rect 111 434 115 438
rect 135 434 139 438
rect 199 434 203 438
rect 319 434 323 438
rect 415 434 419 438
rect 551 434 555 438
rect 631 434 635 438
rect 807 434 811 438
rect 855 434 859 438
rect 1071 434 1075 438
rect 1087 434 1091 438
rect 1327 434 1331 438
rect 1343 434 1347 438
rect 111 330 115 334
rect 223 330 227 334
rect 439 330 443 334
rect 559 330 563 334
rect 655 330 659 334
rect 759 330 763 334
rect 879 330 883 334
rect 111 218 115 222
rect 487 218 491 222
rect 535 218 539 222
rect 967 330 971 334
rect 1111 330 1115 334
rect 1575 434 1579 438
rect 1719 546 1723 550
rect 1719 434 1723 438
rect 1183 330 1187 334
rect 1351 330 1355 334
rect 1399 330 1403 334
rect 1599 330 1603 334
rect 623 218 627 222
rect 735 218 739 222
rect 759 218 763 222
rect 895 218 899 222
rect 943 218 947 222
rect 1031 218 1035 222
rect 1159 218 1163 222
rect 1167 218 1171 222
rect 1303 218 1307 222
rect 1375 218 1379 222
rect 1439 218 1443 222
rect 1575 218 1579 222
rect 1719 330 1723 334
rect 1719 218 1723 222
rect 111 118 115 122
rect 511 118 515 122
rect 647 118 651 122
rect 783 118 787 122
rect 919 118 923 122
rect 1055 118 1059 122
rect 1191 118 1195 122
rect 1327 118 1331 122
rect 1463 118 1467 122
rect 1599 118 1603 122
rect 1719 118 1723 122
<< m4 >>
rect 96 1777 97 1783
rect 103 1782 1755 1783
rect 103 1778 111 1782
rect 115 1778 135 1782
rect 139 1778 271 1782
rect 275 1778 407 1782
rect 411 1778 543 1782
rect 547 1778 679 1782
rect 683 1778 1719 1782
rect 1723 1778 1755 1782
rect 103 1777 1755 1778
rect 1761 1777 1762 1783
rect 84 1669 85 1675
rect 91 1674 1743 1675
rect 91 1670 111 1674
rect 115 1670 159 1674
rect 163 1670 239 1674
rect 243 1670 295 1674
rect 299 1670 375 1674
rect 379 1670 431 1674
rect 435 1670 511 1674
rect 515 1670 567 1674
rect 571 1670 647 1674
rect 651 1670 703 1674
rect 707 1670 783 1674
rect 787 1670 1719 1674
rect 1723 1670 1743 1674
rect 91 1669 1743 1670
rect 1749 1669 1750 1675
rect 96 1553 97 1559
rect 103 1558 1755 1559
rect 103 1554 111 1558
rect 115 1554 215 1558
rect 219 1554 351 1558
rect 355 1554 487 1558
rect 491 1554 599 1558
rect 603 1554 623 1558
rect 627 1554 735 1558
rect 739 1554 759 1558
rect 763 1554 871 1558
rect 875 1554 1015 1558
rect 1019 1554 1159 1558
rect 1163 1554 1303 1558
rect 1307 1554 1439 1558
rect 1443 1554 1575 1558
rect 1579 1554 1719 1558
rect 1723 1554 1755 1558
rect 103 1553 1755 1554
rect 1761 1553 1762 1559
rect 84 1449 85 1455
rect 91 1454 1743 1455
rect 91 1450 111 1454
rect 115 1450 599 1454
rect 603 1450 623 1454
rect 627 1450 735 1454
rect 739 1450 759 1454
rect 763 1450 879 1454
rect 883 1450 895 1454
rect 899 1450 1023 1454
rect 1027 1450 1039 1454
rect 1043 1450 1167 1454
rect 1171 1450 1183 1454
rect 1187 1450 1319 1454
rect 1323 1450 1327 1454
rect 1331 1450 1463 1454
rect 1467 1450 1599 1454
rect 1603 1450 1719 1454
rect 1723 1450 1743 1454
rect 91 1449 1743 1450
rect 1749 1449 1750 1455
rect 96 1333 97 1339
rect 103 1338 1755 1339
rect 103 1334 111 1338
rect 115 1334 135 1338
rect 139 1334 303 1338
rect 307 1334 519 1338
rect 523 1334 575 1338
rect 579 1334 711 1338
rect 715 1334 751 1338
rect 755 1334 855 1338
rect 859 1334 999 1338
rect 1003 1334 1143 1338
rect 1147 1334 1255 1338
rect 1259 1334 1295 1338
rect 1299 1334 1439 1338
rect 1443 1334 1519 1338
rect 1523 1334 1575 1338
rect 1579 1334 1719 1338
rect 1723 1334 1755 1338
rect 103 1333 1755 1334
rect 1761 1333 1762 1339
rect 84 1221 85 1227
rect 91 1226 1743 1227
rect 91 1222 111 1226
rect 115 1222 159 1226
rect 163 1222 327 1226
rect 331 1222 399 1226
rect 403 1222 543 1226
rect 547 1222 671 1226
rect 675 1222 775 1226
rect 779 1222 959 1226
rect 963 1222 1023 1226
rect 1027 1222 1255 1226
rect 1259 1222 1279 1226
rect 1283 1222 1543 1226
rect 1547 1222 1551 1226
rect 1555 1222 1719 1226
rect 1723 1222 1743 1226
rect 91 1221 1743 1222
rect 1749 1221 1750 1227
rect 96 1121 97 1127
rect 103 1126 1755 1127
rect 103 1122 111 1126
rect 115 1122 135 1126
rect 139 1122 191 1126
rect 195 1122 375 1126
rect 379 1122 415 1126
rect 419 1122 647 1126
rect 651 1122 671 1126
rect 675 1122 935 1126
rect 939 1122 951 1126
rect 955 1122 1231 1126
rect 1235 1122 1247 1126
rect 1251 1122 1527 1126
rect 1531 1122 1543 1126
rect 1547 1122 1719 1126
rect 1723 1122 1755 1126
rect 103 1121 1755 1122
rect 1761 1121 1762 1127
rect 84 1005 85 1011
rect 91 1010 1743 1011
rect 91 1006 111 1010
rect 115 1006 215 1010
rect 219 1006 439 1010
rect 443 1006 511 1010
rect 515 1006 663 1010
rect 667 1006 695 1010
rect 699 1006 831 1010
rect 835 1006 975 1010
rect 979 1006 1007 1010
rect 1011 1006 1199 1010
rect 1203 1006 1271 1010
rect 1275 1006 1399 1010
rect 1403 1006 1567 1010
rect 1571 1006 1599 1010
rect 1603 1006 1719 1010
rect 1723 1006 1743 1010
rect 91 1005 1743 1006
rect 1749 1005 1750 1011
rect 96 893 97 899
rect 103 898 1755 899
rect 103 894 111 898
rect 115 894 487 898
rect 491 894 639 898
rect 643 894 759 898
rect 763 894 807 898
rect 811 894 911 898
rect 915 894 983 898
rect 987 894 1071 898
rect 1075 894 1175 898
rect 1179 894 1239 898
rect 1243 894 1375 898
rect 1379 894 1407 898
rect 1411 894 1575 898
rect 1579 894 1719 898
rect 1723 894 1755 898
rect 103 893 1755 894
rect 1761 893 1762 899
rect 84 785 85 791
rect 91 790 1743 791
rect 91 786 111 790
rect 115 786 695 790
rect 699 786 783 790
rect 787 786 831 790
rect 835 786 935 790
rect 939 786 975 790
rect 979 786 1095 790
rect 1099 786 1119 790
rect 1123 786 1263 790
rect 1267 786 1271 790
rect 1275 786 1431 790
rect 1435 786 1599 790
rect 1603 786 1719 790
rect 1723 786 1743 790
rect 91 785 1743 786
rect 1749 785 1750 791
rect 96 661 97 667
rect 103 666 1755 667
rect 103 662 111 666
rect 115 662 247 666
rect 251 662 431 666
rect 435 662 631 666
rect 635 662 671 666
rect 675 662 807 666
rect 811 662 847 666
rect 851 662 951 666
rect 955 662 1079 666
rect 1083 662 1095 666
rect 1099 662 1247 666
rect 1251 662 1319 666
rect 1323 662 1407 666
rect 1411 662 1559 666
rect 1563 662 1575 666
rect 1579 662 1719 666
rect 1723 662 1755 666
rect 103 661 1755 662
rect 1761 661 1762 667
rect 84 545 85 551
rect 91 550 1743 551
rect 91 546 111 550
rect 115 546 159 550
rect 163 546 271 550
rect 275 546 343 550
rect 347 546 455 550
rect 459 546 575 550
rect 579 546 655 550
rect 659 546 831 550
rect 835 546 871 550
rect 875 546 1095 550
rect 1099 546 1103 550
rect 1107 546 1343 550
rect 1347 546 1367 550
rect 1371 546 1583 550
rect 1587 546 1719 550
rect 1723 546 1743 550
rect 91 545 1743 546
rect 1749 545 1750 551
rect 96 433 97 439
rect 103 438 1755 439
rect 103 434 111 438
rect 115 434 135 438
rect 139 434 199 438
rect 203 434 319 438
rect 323 434 415 438
rect 419 434 551 438
rect 555 434 631 438
rect 635 434 807 438
rect 811 434 855 438
rect 859 434 1071 438
rect 1075 434 1087 438
rect 1091 434 1327 438
rect 1331 434 1343 438
rect 1347 434 1575 438
rect 1579 434 1719 438
rect 1723 434 1755 438
rect 103 433 1755 434
rect 1761 433 1762 439
rect 84 329 85 335
rect 91 334 1743 335
rect 91 330 111 334
rect 115 330 223 334
rect 227 330 439 334
rect 443 330 559 334
rect 563 330 655 334
rect 659 330 759 334
rect 763 330 879 334
rect 883 330 967 334
rect 971 330 1111 334
rect 1115 330 1183 334
rect 1187 330 1351 334
rect 1355 330 1399 334
rect 1403 330 1599 334
rect 1603 330 1719 334
rect 1723 330 1743 334
rect 91 329 1743 330
rect 1749 329 1750 335
rect 96 217 97 223
rect 103 222 1755 223
rect 103 218 111 222
rect 115 218 487 222
rect 491 218 535 222
rect 539 218 623 222
rect 627 218 735 222
rect 739 218 759 222
rect 763 218 895 222
rect 899 218 943 222
rect 947 218 1031 222
rect 1035 218 1159 222
rect 1163 218 1167 222
rect 1171 218 1303 222
rect 1307 218 1375 222
rect 1379 218 1439 222
rect 1443 218 1575 222
rect 1579 218 1719 222
rect 1723 218 1755 222
rect 103 217 1755 218
rect 1761 217 1762 223
rect 84 117 85 123
rect 91 122 1743 123
rect 91 118 111 122
rect 115 118 511 122
rect 515 118 647 122
rect 651 118 783 122
rect 787 118 919 122
rect 923 118 1055 122
rect 1059 118 1191 122
rect 1195 118 1327 122
rect 1331 118 1463 122
rect 1467 118 1599 122
rect 1603 118 1719 122
rect 1723 118 1743 122
rect 91 117 1743 118
rect 1749 117 1750 123
<< m5c >>
rect 97 1777 103 1783
rect 1755 1777 1761 1783
rect 85 1669 91 1675
rect 1743 1669 1749 1675
rect 97 1553 103 1559
rect 1755 1553 1761 1559
rect 85 1449 91 1455
rect 1743 1449 1749 1455
rect 97 1333 103 1339
rect 1755 1333 1761 1339
rect 85 1221 91 1227
rect 1743 1221 1749 1227
rect 97 1121 103 1127
rect 1755 1121 1761 1127
rect 85 1005 91 1011
rect 1743 1005 1749 1011
rect 97 893 103 899
rect 1755 893 1761 899
rect 85 785 91 791
rect 1743 785 1749 791
rect 97 661 103 667
rect 1755 661 1761 667
rect 85 545 91 551
rect 1743 545 1749 551
rect 97 433 103 439
rect 1755 433 1761 439
rect 85 329 91 335
rect 1743 329 1749 335
rect 97 217 103 223
rect 1755 217 1761 223
rect 85 117 91 123
rect 1743 117 1749 123
<< m5 >>
rect 84 1675 92 1800
rect 84 1669 85 1675
rect 91 1669 92 1675
rect 84 1455 92 1669
rect 84 1449 85 1455
rect 91 1449 92 1455
rect 84 1227 92 1449
rect 84 1221 85 1227
rect 91 1221 92 1227
rect 84 1011 92 1221
rect 84 1005 85 1011
rect 91 1005 92 1011
rect 84 791 92 1005
rect 84 785 85 791
rect 91 785 92 791
rect 84 551 92 785
rect 84 545 85 551
rect 91 545 92 551
rect 84 335 92 545
rect 84 329 85 335
rect 91 329 92 335
rect 84 123 92 329
rect 84 117 85 123
rect 91 117 92 123
rect 84 72 92 117
rect 96 1783 104 1800
rect 96 1777 97 1783
rect 103 1777 104 1783
rect 96 1559 104 1777
rect 96 1553 97 1559
rect 103 1553 104 1559
rect 96 1339 104 1553
rect 96 1333 97 1339
rect 103 1333 104 1339
rect 96 1127 104 1333
rect 96 1121 97 1127
rect 103 1121 104 1127
rect 96 899 104 1121
rect 96 893 97 899
rect 103 893 104 899
rect 96 667 104 893
rect 96 661 97 667
rect 103 661 104 667
rect 96 439 104 661
rect 96 433 97 439
rect 103 433 104 439
rect 96 223 104 433
rect 96 217 97 223
rect 103 217 104 223
rect 96 72 104 217
rect 1742 1675 1750 1800
rect 1742 1669 1743 1675
rect 1749 1669 1750 1675
rect 1742 1455 1750 1669
rect 1742 1449 1743 1455
rect 1749 1449 1750 1455
rect 1742 1227 1750 1449
rect 1742 1221 1743 1227
rect 1749 1221 1750 1227
rect 1742 1011 1750 1221
rect 1742 1005 1743 1011
rect 1749 1005 1750 1011
rect 1742 791 1750 1005
rect 1742 785 1743 791
rect 1749 785 1750 791
rect 1742 551 1750 785
rect 1742 545 1743 551
rect 1749 545 1750 551
rect 1742 335 1750 545
rect 1742 329 1743 335
rect 1749 329 1750 335
rect 1742 123 1750 329
rect 1742 117 1743 123
rect 1749 117 1750 123
rect 1742 72 1750 117
rect 1754 1783 1762 1800
rect 1754 1777 1755 1783
rect 1761 1777 1762 1783
rect 1754 1559 1762 1777
rect 1754 1553 1755 1559
rect 1761 1553 1762 1559
rect 1754 1339 1762 1553
rect 1754 1333 1755 1339
rect 1761 1333 1762 1339
rect 1754 1127 1762 1333
rect 1754 1121 1755 1127
rect 1761 1121 1762 1127
rect 1754 899 1762 1121
rect 1754 893 1755 899
rect 1761 893 1762 899
rect 1754 667 1762 893
rect 1754 661 1755 667
rect 1761 661 1762 667
rect 1754 439 1762 661
rect 1754 433 1755 439
rect 1761 433 1762 439
rect 1754 223 1762 433
rect 1754 217 1755 223
rect 1761 217 1762 223
rect 1754 72 1762 217
use welltap_svt  __well_tap__0
timestamp 1730768254
transform 1 0 104 0 1 144
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__0
timestamp 1730768254
transform 1 0 104 0 1 144
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0FAX1  fax_566_6
timestamp 1730768254
transform 1 0 480 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_566_6
timestamp 1730768254
transform 1 0 480 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_567_6
timestamp 1730768254
transform 1 0 616 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_567_6
timestamp 1730768254
transform 1 0 616 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_568_6
timestamp 1730768254
transform 1 0 752 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_568_6
timestamp 1730768254
transform 1 0 752 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_569_6
timestamp 1730768254
transform 1 0 888 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_569_6
timestamp 1730768254
transform 1 0 888 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_570_6
timestamp 1730768254
transform 1 0 1024 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_570_6
timestamp 1730768254
transform 1 0 1024 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_571_6
timestamp 1730768254
transform 1 0 1160 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_571_6
timestamp 1730768254
transform 1 0 1160 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_572_6
timestamp 1730768254
transform 1 0 1296 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_572_6
timestamp 1730768254
transform 1 0 1296 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_599_6
timestamp 1730768254
transform 1 0 1432 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_599_6
timestamp 1730768254
transform 1 0 1432 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_598_6
timestamp 1730768254
transform 1 0 1568 0 1 120
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_598_6
timestamp 1730768254
transform 1 0 1568 0 1 120
box 8 5 126 98
use welltap_svt  __well_tap__1
timestamp 1730768254
transform 1 0 1712 0 1 144
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730768254
transform 1 0 1712 0 1 144
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_565_6
timestamp 1730768254
transform 1 0 528 0 -1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_565_6
timestamp 1730768254
transform 1 0 528 0 -1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_564_6
timestamp 1730768254
transform 1 0 728 0 -1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_564_6
timestamp 1730768254
transform 1 0 728 0 -1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_563_6
timestamp 1730768254
transform 1 0 936 0 -1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_563_6
timestamp 1730768254
transform 1 0 936 0 -1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_574_6
timestamp 1730768254
transform 1 0 1152 0 -1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_574_6
timestamp 1730768254
transform 1 0 1152 0 -1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_573_6
timestamp 1730768254
transform 1 0 1368 0 -1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_573_6
timestamp 1730768254
transform 1 0 1368 0 -1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_597_6
timestamp 1730768254
transform 1 0 1568 0 -1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_597_6
timestamp 1730768254
transform 1 0 1568 0 -1 332
box 8 5 126 98
use welltap_svt  __well_tap__2
timestamp 1730768254
transform 1 0 104 0 -1 308
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730768254
transform 1 0 104 0 -1 308
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_559_6
timestamp 1730768254
transform 1 0 192 0 1 336
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_559_6
timestamp 1730768254
transform 1 0 192 0 1 336
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_560_6
timestamp 1730768254
transform 1 0 408 0 1 336
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_560_6
timestamp 1730768254
transform 1 0 408 0 1 336
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_561_6
timestamp 1730768254
transform 1 0 624 0 1 336
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_561_6
timestamp 1730768254
transform 1 0 624 0 1 336
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_562_6
timestamp 1730768254
transform 1 0 848 0 1 336
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_562_6
timestamp 1730768254
transform 1 0 848 0 1 336
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_575_6
timestamp 1730768254
transform 1 0 1080 0 1 336
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_575_6
timestamp 1730768254
transform 1 0 1080 0 1 336
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_576_6
timestamp 1730768254
transform 1 0 1320 0 1 336
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_576_6
timestamp 1730768254
transform 1 0 1320 0 1 336
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_596_6
timestamp 1730768254
transform 1 0 1568 0 1 336
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_596_6
timestamp 1730768254
transform 1 0 1568 0 1 336
box 8 5 126 98
use welltap_svt  __well_tap__3
timestamp 1730768254
transform 1 0 1712 0 -1 308
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730768254
transform 1 0 1712 0 -1 308
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730768254
transform 1 0 104 0 1 360
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730768254
transform 1 0 104 0 1 360
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730768254
transform 1 0 1712 0 1 360
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730768254
transform 1 0 1712 0 1 360
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_554_6
timestamp 1730768254
transform 1 0 128 0 -1 548
box 8 5 126 98
use welltap_svt  __well_tap__6
timestamp 1730768254
transform 1 0 104 0 -1 524
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_554_6
timestamp 1730768254
transform 1 0 128 0 -1 548
box 8 5 126 98
use welltap_svt  __well_tap__6
timestamp 1730768254
transform 1 0 104 0 -1 524
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_555_6
timestamp 1730768254
transform 1 0 312 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_555_6
timestamp 1730768254
transform 1 0 312 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_556_6
timestamp 1730768254
transform 1 0 544 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_556_6
timestamp 1730768254
transform 1 0 544 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_557_6
timestamp 1730768254
transform 1 0 800 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_557_6
timestamp 1730768254
transform 1 0 800 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_558_6
timestamp 1730768254
transform 1 0 1064 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_558_6
timestamp 1730768254
transform 1 0 1064 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_577_6
timestamp 1730768254
transform 1 0 1336 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_577_6
timestamp 1730768254
transform 1 0 1336 0 -1 548
box 8 5 126 98
use welltap_svt  __well_tap__7
timestamp 1730768254
transform 1 0 1712 0 -1 524
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730768254
transform 1 0 1712 0 -1 524
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730768254
transform 1 0 104 0 1 588
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730768254
transform 1 0 104 0 1 588
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_553_6
timestamp 1730768254
transform 1 0 240 0 1 564
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_553_6
timestamp 1730768254
transform 1 0 240 0 1 564
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_552_6
timestamp 1730768254
transform 1 0 424 0 1 564
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_552_6
timestamp 1730768254
transform 1 0 424 0 1 564
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_551_6
timestamp 1730768254
transform 1 0 624 0 1 564
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_551_6
timestamp 1730768254
transform 1 0 624 0 1 564
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_550_6
timestamp 1730768254
transform 1 0 840 0 1 564
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_550_6
timestamp 1730768254
transform 1 0 840 0 1 564
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_549_6
timestamp 1730768254
transform 1 0 1072 0 1 564
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_549_6
timestamp 1730768254
transform 1 0 1072 0 1 564
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_578_6
timestamp 1730768254
transform 1 0 1312 0 1 564
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_578_6
timestamp 1730768254
transform 1 0 1312 0 1 564
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_595_6
timestamp 1730768254
transform 1 0 1552 0 1 564
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_595_6
timestamp 1730768254
transform 1 0 1552 0 1 564
box 8 5 126 98
use welltap_svt  __well_tap__9
timestamp 1730768254
transform 1 0 1712 0 1 588
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730768254
transform 1 0 1712 0 1 588
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_546_6
timestamp 1730768254
transform 1 0 664 0 -1 788
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_546_6
timestamp 1730768254
transform 1 0 664 0 -1 788
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_547_6
timestamp 1730768254
transform 1 0 800 0 -1 788
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_547_6
timestamp 1730768254
transform 1 0 800 0 -1 788
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_548_6
timestamp 1730768254
transform 1 0 944 0 -1 788
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_548_6
timestamp 1730768254
transform 1 0 944 0 -1 788
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_545_6
timestamp 1730768254
transform 1 0 1088 0 -1 788
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_545_6
timestamp 1730768254
transform 1 0 1088 0 -1 788
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_544_6
timestamp 1730768254
transform 1 0 1240 0 -1 788
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_544_6
timestamp 1730768254
transform 1 0 1240 0 -1 788
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_579_6
timestamp 1730768254
transform 1 0 1400 0 -1 788
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_579_6
timestamp 1730768254
transform 1 0 1400 0 -1 788
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_594_6
timestamp 1730768254
transform 1 0 1568 0 -1 788
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_594_6
timestamp 1730768254
transform 1 0 1568 0 -1 788
box 8 5 126 98
use welltap_svt  __well_tap__10
timestamp 1730768254
transform 1 0 104 0 -1 764
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730768254
transform 1 0 104 0 -1 764
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_539_6
timestamp 1730768254
transform 1 0 752 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_539_6
timestamp 1730768254
transform 1 0 752 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_540_6
timestamp 1730768254
transform 1 0 904 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_540_6
timestamp 1730768254
transform 1 0 904 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_541_6
timestamp 1730768254
transform 1 0 1064 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_541_6
timestamp 1730768254
transform 1 0 1064 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_542_6
timestamp 1730768254
transform 1 0 1232 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_542_6
timestamp 1730768254
transform 1 0 1232 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_543_6
timestamp 1730768254
transform 1 0 1400 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_543_6
timestamp 1730768254
transform 1 0 1400 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_593_6
timestamp 1730768254
transform 1 0 1568 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_593_6
timestamp 1730768254
transform 1 0 1568 0 1 796
box 8 5 126 98
use welltap_svt  __well_tap__11
timestamp 1730768254
transform 1 0 1712 0 -1 764
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730768254
transform 1 0 1712 0 -1 764
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730768254
transform 1 0 104 0 1 820
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730768254
transform 1 0 104 0 1 820
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_534_6
timestamp 1730768254
transform 1 0 480 0 -1 1008
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_534_6
timestamp 1730768254
transform 1 0 480 0 -1 1008
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_535_6
timestamp 1730768254
transform 1 0 632 0 -1 1008
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_535_6
timestamp 1730768254
transform 1 0 632 0 -1 1008
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_536_6
timestamp 1730768254
transform 1 0 800 0 -1 1008
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_536_6
timestamp 1730768254
transform 1 0 800 0 -1 1008
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_537_6
timestamp 1730768254
transform 1 0 976 0 -1 1008
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_537_6
timestamp 1730768254
transform 1 0 976 0 -1 1008
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_538_6
timestamp 1730768254
transform 1 0 1168 0 -1 1008
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_538_6
timestamp 1730768254
transform 1 0 1168 0 -1 1008
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_580_6
timestamp 1730768254
transform 1 0 1368 0 -1 1008
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_580_6
timestamp 1730768254
transform 1 0 1368 0 -1 1008
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_592_6
timestamp 1730768254
transform 1 0 1568 0 -1 1008
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_592_6
timestamp 1730768254
transform 1 0 1568 0 -1 1008
box 8 5 126 98
use welltap_svt  __well_tap__13
timestamp 1730768254
transform 1 0 1712 0 1 820
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730768254
transform 1 0 1712 0 1 820
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730768254
transform 1 0 104 0 -1 984
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730768254
transform 1 0 104 0 -1 984
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730768254
transform 1 0 1712 0 -1 984
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730768254
transform 1 0 1712 0 -1 984
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_529_6
timestamp 1730768254
transform 1 0 184 0 1 1024
box 8 5 126 98
use welltap_svt  __well_tap__16
timestamp 1730768254
transform 1 0 104 0 1 1048
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_529_6
timestamp 1730768254
transform 1 0 184 0 1 1024
box 8 5 126 98
use welltap_svt  __well_tap__16
timestamp 1730768254
transform 1 0 104 0 1 1048
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_530_6
timestamp 1730768254
transform 1 0 408 0 1 1024
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_530_6
timestamp 1730768254
transform 1 0 408 0 1 1024
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_531_6
timestamp 1730768254
transform 1 0 664 0 1 1024
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_531_6
timestamp 1730768254
transform 1 0 664 0 1 1024
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_532_6
timestamp 1730768254
transform 1 0 944 0 1 1024
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_532_6
timestamp 1730768254
transform 1 0 944 0 1 1024
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_533_6
timestamp 1730768254
transform 1 0 1240 0 1 1024
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_533_6
timestamp 1730768254
transform 1 0 1240 0 1 1024
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_591_6
timestamp 1730768254
transform 1 0 1536 0 1 1024
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_591_6
timestamp 1730768254
transform 1 0 1536 0 1 1024
box 8 5 126 98
use welltap_svt  __well_tap__17
timestamp 1730768254
transform 1 0 1712 0 1 1048
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730768254
transform 1 0 1712 0 1 1048
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_525_6
timestamp 1730768254
transform 1 0 128 0 -1 1224
box 8 5 126 98
use welltap_svt  __well_tap__18
timestamp 1730768254
transform 1 0 104 0 -1 1200
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_525_6
timestamp 1730768254
transform 1 0 128 0 -1 1224
box 8 5 126 98
use welltap_svt  __well_tap__18
timestamp 1730768254
transform 1 0 104 0 -1 1200
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_526_6
timestamp 1730768254
transform 1 0 368 0 -1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_526_6
timestamp 1730768254
transform 1 0 368 0 -1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_527_6
timestamp 1730768254
transform 1 0 640 0 -1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_527_6
timestamp 1730768254
transform 1 0 640 0 -1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_528_6
timestamp 1730768254
transform 1 0 928 0 -1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_528_6
timestamp 1730768254
transform 1 0 928 0 -1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_581_6
timestamp 1730768254
transform 1 0 1224 0 -1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_581_6
timestamp 1730768254
transform 1 0 1224 0 -1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_590_6
timestamp 1730768254
transform 1 0 1520 0 -1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_590_6
timestamp 1730768254
transform 1 0 1520 0 -1 1224
box 8 5 126 98
use welltap_svt  __well_tap__19
timestamp 1730768254
transform 1 0 1712 0 -1 1200
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730768254
transform 1 0 1712 0 -1 1200
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_524_6
timestamp 1730768254
transform 1 0 128 0 1 1236
box 8 5 126 98
use welltap_svt  __well_tap__20
timestamp 1730768254
transform 1 0 104 0 1 1260
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_524_6
timestamp 1730768254
transform 1 0 128 0 1 1236
box 8 5 126 98
use welltap_svt  __well_tap__20
timestamp 1730768254
transform 1 0 104 0 1 1260
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_523_6
timestamp 1730768254
transform 1 0 296 0 1 1236
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_523_6
timestamp 1730768254
transform 1 0 296 0 1 1236
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_522_6
timestamp 1730768254
transform 1 0 512 0 1 1236
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_522_6
timestamp 1730768254
transform 1 0 512 0 1 1236
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_521_6
timestamp 1730768254
transform 1 0 744 0 1 1236
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_521_6
timestamp 1730768254
transform 1 0 744 0 1 1236
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_520_6
timestamp 1730768254
transform 1 0 992 0 1 1236
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_520_6
timestamp 1730768254
transform 1 0 992 0 1 1236
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_582_6
timestamp 1730768254
transform 1 0 1248 0 1 1236
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_582_6
timestamp 1730768254
transform 1 0 1248 0 1 1236
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_589_6
timestamp 1730768254
transform 1 0 1512 0 1 1236
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_589_6
timestamp 1730768254
transform 1 0 1512 0 1 1236
box 8 5 126 98
use welltap_svt  __well_tap__21
timestamp 1730768254
transform 1 0 1712 0 1 1260
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730768254
transform 1 0 1712 0 1 1260
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_517_6
timestamp 1730768254
transform 1 0 568 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_517_6
timestamp 1730768254
transform 1 0 568 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_518_6
timestamp 1730768254
transform 1 0 704 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_518_6
timestamp 1730768254
transform 1 0 704 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_519_6
timestamp 1730768254
transform 1 0 848 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_519_6
timestamp 1730768254
transform 1 0 848 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_516_6
timestamp 1730768254
transform 1 0 992 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_516_6
timestamp 1730768254
transform 1 0 992 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_515_6
timestamp 1730768254
transform 1 0 1136 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_515_6
timestamp 1730768254
transform 1 0 1136 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_583_6
timestamp 1730768254
transform 1 0 1288 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_583_6
timestamp 1730768254
transform 1 0 1288 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_588_6
timestamp 1730768254
transform 1 0 1432 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_588_6
timestamp 1730768254
transform 1 0 1432 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_587_6
timestamp 1730768254
transform 1 0 1568 0 -1 1452
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_587_6
timestamp 1730768254
transform 1 0 1568 0 -1 1452
box 8 5 126 98
use welltap_svt  __well_tap__22
timestamp 1730768254
transform 1 0 104 0 -1 1428
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730768254
transform 1 0 104 0 -1 1428
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_510_6
timestamp 1730768254
transform 1 0 592 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_510_6
timestamp 1730768254
transform 1 0 592 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_511_6
timestamp 1730768254
transform 1 0 728 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_511_6
timestamp 1730768254
transform 1 0 728 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_512_6
timestamp 1730768254
transform 1 0 864 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_512_6
timestamp 1730768254
transform 1 0 864 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_513_6
timestamp 1730768254
transform 1 0 1008 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_513_6
timestamp 1730768254
transform 1 0 1008 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_514_6
timestamp 1730768254
transform 1 0 1152 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_514_6
timestamp 1730768254
transform 1 0 1152 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_584_6
timestamp 1730768254
transform 1 0 1296 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_584_6
timestamp 1730768254
transform 1 0 1296 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_585_6
timestamp 1730768254
transform 1 0 1432 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_585_6
timestamp 1730768254
transform 1 0 1432 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_586_6
timestamp 1730768254
transform 1 0 1568 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_586_6
timestamp 1730768254
transform 1 0 1568 0 1 1456
box 8 5 126 98
use welltap_svt  __well_tap__23
timestamp 1730768254
transform 1 0 1712 0 -1 1428
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730768254
transform 1 0 1712 0 -1 1428
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730768254
transform 1 0 104 0 1 1480
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730768254
transform 1 0 104 0 1 1480
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_55_6
timestamp 1730768254
transform 1 0 208 0 -1 1672
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_55_6
timestamp 1730768254
transform 1 0 208 0 -1 1672
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_56_6
timestamp 1730768254
transform 1 0 344 0 -1 1672
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_56_6
timestamp 1730768254
transform 1 0 344 0 -1 1672
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_57_6
timestamp 1730768254
transform 1 0 480 0 -1 1672
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_57_6
timestamp 1730768254
transform 1 0 480 0 -1 1672
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_58_6
timestamp 1730768254
transform 1 0 616 0 -1 1672
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_58_6
timestamp 1730768254
transform 1 0 616 0 -1 1672
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_59_6
timestamp 1730768254
transform 1 0 752 0 -1 1672
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_59_6
timestamp 1730768254
transform 1 0 752 0 -1 1672
box 8 5 126 98
use welltap_svt  __well_tap__25
timestamp 1730768254
transform 1 0 1712 0 1 1480
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730768254
transform 1 0 1712 0 1 1480
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730768254
transform 1 0 104 0 -1 1648
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730768254
transform 1 0 104 0 -1 1648
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730768254
transform 1 0 1712 0 -1 1648
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730768254
transform 1 0 1712 0 -1 1648
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_50_6
timestamp 1730768254
transform 1 0 128 0 1 1680
box 8 5 126 98
use welltap_svt  __well_tap__28
timestamp 1730768254
transform 1 0 104 0 1 1704
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_50_6
timestamp 1730768254
transform 1 0 128 0 1 1680
box 8 5 126 98
use welltap_svt  __well_tap__28
timestamp 1730768254
transform 1 0 104 0 1 1704
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_51_6
timestamp 1730768254
transform 1 0 264 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_51_6
timestamp 1730768254
transform 1 0 264 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_52_6
timestamp 1730768254
transform 1 0 400 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_52_6
timestamp 1730768254
transform 1 0 400 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_53_6
timestamp 1730768254
transform 1 0 536 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_53_6
timestamp 1730768254
transform 1 0 536 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_54_6
timestamp 1730768254
transform 1 0 672 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_54_6
timestamp 1730768254
transform 1 0 672 0 1 1680
box 8 5 126 98
use welltap_svt  __well_tap__29
timestamp 1730768254
transform 1 0 1712 0 1 1704
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1730768254
transform 1 0 1712 0 1 1704
box 8 4 12 24
<< end >>
