magic
tech sky130l
timestamp 1731220339
<< m2 >>
rect 2070 3992 2076 3993
rect 2046 3989 2052 3990
rect 2046 3985 2047 3989
rect 2051 3985 2052 3989
rect 2070 3988 2071 3992
rect 2075 3988 2076 3992
rect 2070 3987 2076 3988
rect 2326 3992 2332 3993
rect 2326 3988 2327 3992
rect 2331 3988 2332 3992
rect 2326 3987 2332 3988
rect 2590 3992 2596 3993
rect 2590 3988 2591 3992
rect 2595 3988 2596 3992
rect 2590 3987 2596 3988
rect 2838 3992 2844 3993
rect 2838 3988 2839 3992
rect 2843 3988 2844 3992
rect 2838 3987 2844 3988
rect 3086 3992 3092 3993
rect 3086 3988 3087 3992
rect 3091 3988 3092 3992
rect 3086 3987 3092 3988
rect 3342 3992 3348 3993
rect 3342 3988 3343 3992
rect 3347 3988 3348 3992
rect 3342 3987 3348 3988
rect 3942 3989 3948 3990
rect 2046 3984 2052 3985
rect 3942 3985 3943 3989
rect 3947 3985 3948 3989
rect 3942 3984 3948 3985
rect 2070 3973 2076 3974
rect 310 3972 316 3973
rect 110 3969 116 3970
rect 110 3965 111 3969
rect 115 3965 116 3969
rect 310 3968 311 3972
rect 315 3968 316 3972
rect 310 3967 316 3968
rect 510 3972 516 3973
rect 510 3968 511 3972
rect 515 3968 516 3972
rect 510 3967 516 3968
rect 702 3972 708 3973
rect 702 3968 703 3972
rect 707 3968 708 3972
rect 702 3967 708 3968
rect 886 3972 892 3973
rect 886 3968 887 3972
rect 891 3968 892 3972
rect 886 3967 892 3968
rect 1062 3972 1068 3973
rect 1062 3968 1063 3972
rect 1067 3968 1068 3972
rect 1062 3967 1068 3968
rect 1230 3972 1236 3973
rect 1230 3968 1231 3972
rect 1235 3968 1236 3972
rect 1230 3967 1236 3968
rect 1382 3972 1388 3973
rect 1382 3968 1383 3972
rect 1387 3968 1388 3972
rect 1382 3967 1388 3968
rect 1518 3972 1524 3973
rect 1518 3968 1519 3972
rect 1523 3968 1524 3972
rect 1518 3967 1524 3968
rect 1654 3972 1660 3973
rect 1654 3968 1655 3972
rect 1659 3968 1660 3972
rect 1654 3967 1660 3968
rect 1790 3972 1796 3973
rect 1790 3968 1791 3972
rect 1795 3968 1796 3972
rect 1790 3967 1796 3968
rect 1902 3972 1908 3973
rect 1902 3968 1903 3972
rect 1907 3968 1908 3972
rect 2046 3972 2052 3973
rect 1902 3967 1908 3968
rect 2006 3969 2012 3970
rect 110 3964 116 3965
rect 2006 3965 2007 3969
rect 2011 3965 2012 3969
rect 2046 3968 2047 3972
rect 2051 3968 2052 3972
rect 2070 3969 2071 3973
rect 2075 3969 2076 3973
rect 2070 3968 2076 3969
rect 2326 3973 2332 3974
rect 2326 3969 2327 3973
rect 2331 3969 2332 3973
rect 2326 3968 2332 3969
rect 2590 3973 2596 3974
rect 2590 3969 2591 3973
rect 2595 3969 2596 3973
rect 2590 3968 2596 3969
rect 2838 3973 2844 3974
rect 2838 3969 2839 3973
rect 2843 3969 2844 3973
rect 2838 3968 2844 3969
rect 3086 3973 3092 3974
rect 3086 3969 3087 3973
rect 3091 3969 3092 3973
rect 3086 3968 3092 3969
rect 3342 3973 3348 3974
rect 3342 3969 3343 3973
rect 3347 3969 3348 3973
rect 3342 3968 3348 3969
rect 3942 3972 3948 3973
rect 3942 3968 3943 3972
rect 3947 3968 3948 3972
rect 2046 3967 2052 3968
rect 3942 3967 3948 3968
rect 2006 3964 2012 3965
rect 310 3953 316 3954
rect 110 3952 116 3953
rect 110 3948 111 3952
rect 115 3948 116 3952
rect 310 3949 311 3953
rect 315 3949 316 3953
rect 310 3948 316 3949
rect 510 3953 516 3954
rect 510 3949 511 3953
rect 515 3949 516 3953
rect 510 3948 516 3949
rect 702 3953 708 3954
rect 702 3949 703 3953
rect 707 3949 708 3953
rect 702 3948 708 3949
rect 886 3953 892 3954
rect 886 3949 887 3953
rect 891 3949 892 3953
rect 886 3948 892 3949
rect 1062 3953 1068 3954
rect 1062 3949 1063 3953
rect 1067 3949 1068 3953
rect 1062 3948 1068 3949
rect 1230 3953 1236 3954
rect 1230 3949 1231 3953
rect 1235 3949 1236 3953
rect 1230 3948 1236 3949
rect 1382 3953 1388 3954
rect 1382 3949 1383 3953
rect 1387 3949 1388 3953
rect 1382 3948 1388 3949
rect 1518 3953 1524 3954
rect 1518 3949 1519 3953
rect 1523 3949 1524 3953
rect 1518 3948 1524 3949
rect 1654 3953 1660 3954
rect 1654 3949 1655 3953
rect 1659 3949 1660 3953
rect 1654 3948 1660 3949
rect 1790 3953 1796 3954
rect 1790 3949 1791 3953
rect 1795 3949 1796 3953
rect 1790 3948 1796 3949
rect 1902 3953 1908 3954
rect 1902 3949 1903 3953
rect 1907 3949 1908 3953
rect 1902 3948 1908 3949
rect 2006 3952 2012 3953
rect 2006 3948 2007 3952
rect 2011 3948 2012 3952
rect 110 3947 116 3948
rect 2006 3947 2012 3948
rect 2046 3920 2052 3921
rect 3942 3920 3948 3921
rect 2046 3916 2047 3920
rect 2051 3916 2052 3920
rect 2046 3915 2052 3916
rect 2126 3919 2132 3920
rect 2126 3915 2127 3919
rect 2131 3915 2132 3919
rect 2126 3914 2132 3915
rect 2270 3919 2276 3920
rect 2270 3915 2271 3919
rect 2275 3915 2276 3919
rect 2270 3914 2276 3915
rect 2438 3919 2444 3920
rect 2438 3915 2439 3919
rect 2443 3915 2444 3919
rect 2438 3914 2444 3915
rect 2614 3919 2620 3920
rect 2614 3915 2615 3919
rect 2619 3915 2620 3919
rect 2614 3914 2620 3915
rect 2798 3919 2804 3920
rect 2798 3915 2799 3919
rect 2803 3915 2804 3919
rect 2798 3914 2804 3915
rect 2982 3919 2988 3920
rect 2982 3915 2983 3919
rect 2987 3915 2988 3919
rect 2982 3914 2988 3915
rect 3174 3919 3180 3920
rect 3174 3915 3175 3919
rect 3179 3915 3180 3919
rect 3174 3914 3180 3915
rect 3366 3919 3372 3920
rect 3366 3915 3367 3919
rect 3371 3915 3372 3919
rect 3366 3914 3372 3915
rect 3558 3919 3564 3920
rect 3558 3915 3559 3919
rect 3563 3915 3564 3919
rect 3942 3916 3943 3920
rect 3947 3916 3948 3920
rect 3942 3915 3948 3916
rect 3558 3914 3564 3915
rect 2046 3903 2052 3904
rect 110 3900 116 3901
rect 2006 3900 2012 3901
rect 110 3896 111 3900
rect 115 3896 116 3900
rect 110 3895 116 3896
rect 278 3899 284 3900
rect 278 3895 279 3899
rect 283 3895 284 3899
rect 278 3894 284 3895
rect 414 3899 420 3900
rect 414 3895 415 3899
rect 419 3895 420 3899
rect 414 3894 420 3895
rect 566 3899 572 3900
rect 566 3895 567 3899
rect 571 3895 572 3899
rect 566 3894 572 3895
rect 734 3899 740 3900
rect 734 3895 735 3899
rect 739 3895 740 3899
rect 734 3894 740 3895
rect 910 3899 916 3900
rect 910 3895 911 3899
rect 915 3895 916 3899
rect 910 3894 916 3895
rect 1094 3899 1100 3900
rect 1094 3895 1095 3899
rect 1099 3895 1100 3899
rect 1094 3894 1100 3895
rect 1286 3899 1292 3900
rect 1286 3895 1287 3899
rect 1291 3895 1292 3899
rect 1286 3894 1292 3895
rect 1478 3899 1484 3900
rect 1478 3895 1479 3899
rect 1483 3895 1484 3899
rect 1478 3894 1484 3895
rect 1678 3899 1684 3900
rect 1678 3895 1679 3899
rect 1683 3895 1684 3899
rect 2006 3896 2007 3900
rect 2011 3896 2012 3900
rect 2046 3899 2047 3903
rect 2051 3899 2052 3903
rect 3942 3903 3948 3904
rect 2046 3898 2052 3899
rect 2126 3900 2132 3901
rect 2006 3895 2012 3896
rect 2126 3896 2127 3900
rect 2131 3896 2132 3900
rect 2126 3895 2132 3896
rect 2270 3900 2276 3901
rect 2270 3896 2271 3900
rect 2275 3896 2276 3900
rect 2270 3895 2276 3896
rect 2438 3900 2444 3901
rect 2438 3896 2439 3900
rect 2443 3896 2444 3900
rect 2438 3895 2444 3896
rect 2614 3900 2620 3901
rect 2614 3896 2615 3900
rect 2619 3896 2620 3900
rect 2614 3895 2620 3896
rect 2798 3900 2804 3901
rect 2798 3896 2799 3900
rect 2803 3896 2804 3900
rect 2798 3895 2804 3896
rect 2982 3900 2988 3901
rect 2982 3896 2983 3900
rect 2987 3896 2988 3900
rect 2982 3895 2988 3896
rect 3174 3900 3180 3901
rect 3174 3896 3175 3900
rect 3179 3896 3180 3900
rect 3174 3895 3180 3896
rect 3366 3900 3372 3901
rect 3366 3896 3367 3900
rect 3371 3896 3372 3900
rect 3366 3895 3372 3896
rect 3558 3900 3564 3901
rect 3558 3896 3559 3900
rect 3563 3896 3564 3900
rect 3942 3899 3943 3903
rect 3947 3899 3948 3903
rect 3942 3898 3948 3899
rect 3558 3895 3564 3896
rect 1678 3894 1684 3895
rect 110 3883 116 3884
rect 110 3879 111 3883
rect 115 3879 116 3883
rect 2006 3883 2012 3884
rect 110 3878 116 3879
rect 278 3880 284 3881
rect 278 3876 279 3880
rect 283 3876 284 3880
rect 278 3875 284 3876
rect 414 3880 420 3881
rect 414 3876 415 3880
rect 419 3876 420 3880
rect 414 3875 420 3876
rect 566 3880 572 3881
rect 566 3876 567 3880
rect 571 3876 572 3880
rect 566 3875 572 3876
rect 734 3880 740 3881
rect 734 3876 735 3880
rect 739 3876 740 3880
rect 734 3875 740 3876
rect 910 3880 916 3881
rect 910 3876 911 3880
rect 915 3876 916 3880
rect 910 3875 916 3876
rect 1094 3880 1100 3881
rect 1094 3876 1095 3880
rect 1099 3876 1100 3880
rect 1094 3875 1100 3876
rect 1286 3880 1292 3881
rect 1286 3876 1287 3880
rect 1291 3876 1292 3880
rect 1286 3875 1292 3876
rect 1478 3880 1484 3881
rect 1478 3876 1479 3880
rect 1483 3876 1484 3880
rect 1478 3875 1484 3876
rect 1678 3880 1684 3881
rect 1678 3876 1679 3880
rect 1683 3876 1684 3880
rect 2006 3879 2007 3883
rect 2011 3879 2012 3883
rect 2006 3878 2012 3879
rect 1678 3875 1684 3876
rect 2262 3840 2268 3841
rect 2046 3837 2052 3838
rect 2046 3833 2047 3837
rect 2051 3833 2052 3837
rect 2262 3836 2263 3840
rect 2267 3836 2268 3840
rect 2262 3835 2268 3836
rect 2374 3840 2380 3841
rect 2374 3836 2375 3840
rect 2379 3836 2380 3840
rect 2374 3835 2380 3836
rect 2494 3840 2500 3841
rect 2494 3836 2495 3840
rect 2499 3836 2500 3840
rect 2494 3835 2500 3836
rect 2630 3840 2636 3841
rect 2630 3836 2631 3840
rect 2635 3836 2636 3840
rect 2630 3835 2636 3836
rect 2774 3840 2780 3841
rect 2774 3836 2775 3840
rect 2779 3836 2780 3840
rect 2774 3835 2780 3836
rect 2918 3840 2924 3841
rect 2918 3836 2919 3840
rect 2923 3836 2924 3840
rect 2918 3835 2924 3836
rect 3062 3840 3068 3841
rect 3062 3836 3063 3840
rect 3067 3836 3068 3840
rect 3062 3835 3068 3836
rect 3206 3840 3212 3841
rect 3206 3836 3207 3840
rect 3211 3836 3212 3840
rect 3206 3835 3212 3836
rect 3342 3840 3348 3841
rect 3342 3836 3343 3840
rect 3347 3836 3348 3840
rect 3342 3835 3348 3836
rect 3470 3840 3476 3841
rect 3470 3836 3471 3840
rect 3475 3836 3476 3840
rect 3470 3835 3476 3836
rect 3598 3840 3604 3841
rect 3598 3836 3599 3840
rect 3603 3836 3604 3840
rect 3598 3835 3604 3836
rect 3726 3840 3732 3841
rect 3726 3836 3727 3840
rect 3731 3836 3732 3840
rect 3726 3835 3732 3836
rect 3838 3840 3844 3841
rect 3838 3836 3839 3840
rect 3843 3836 3844 3840
rect 3838 3835 3844 3836
rect 3942 3837 3948 3838
rect 2046 3832 2052 3833
rect 3942 3833 3943 3837
rect 3947 3833 3948 3837
rect 3942 3832 3948 3833
rect 2262 3821 2268 3822
rect 2046 3820 2052 3821
rect 2046 3816 2047 3820
rect 2051 3816 2052 3820
rect 2262 3817 2263 3821
rect 2267 3817 2268 3821
rect 2262 3816 2268 3817
rect 2374 3821 2380 3822
rect 2374 3817 2375 3821
rect 2379 3817 2380 3821
rect 2374 3816 2380 3817
rect 2494 3821 2500 3822
rect 2494 3817 2495 3821
rect 2499 3817 2500 3821
rect 2494 3816 2500 3817
rect 2630 3821 2636 3822
rect 2630 3817 2631 3821
rect 2635 3817 2636 3821
rect 2630 3816 2636 3817
rect 2774 3821 2780 3822
rect 2774 3817 2775 3821
rect 2779 3817 2780 3821
rect 2774 3816 2780 3817
rect 2918 3821 2924 3822
rect 2918 3817 2919 3821
rect 2923 3817 2924 3821
rect 2918 3816 2924 3817
rect 3062 3821 3068 3822
rect 3062 3817 3063 3821
rect 3067 3817 3068 3821
rect 3062 3816 3068 3817
rect 3206 3821 3212 3822
rect 3206 3817 3207 3821
rect 3211 3817 3212 3821
rect 3206 3816 3212 3817
rect 3342 3821 3348 3822
rect 3342 3817 3343 3821
rect 3347 3817 3348 3821
rect 3342 3816 3348 3817
rect 3470 3821 3476 3822
rect 3470 3817 3471 3821
rect 3475 3817 3476 3821
rect 3470 3816 3476 3817
rect 3598 3821 3604 3822
rect 3598 3817 3599 3821
rect 3603 3817 3604 3821
rect 3598 3816 3604 3817
rect 3726 3821 3732 3822
rect 3726 3817 3727 3821
rect 3731 3817 3732 3821
rect 3726 3816 3732 3817
rect 3838 3821 3844 3822
rect 3838 3817 3839 3821
rect 3843 3817 3844 3821
rect 3838 3816 3844 3817
rect 3942 3820 3948 3821
rect 3942 3816 3943 3820
rect 3947 3816 3948 3820
rect 2046 3815 2052 3816
rect 3942 3815 3948 3816
rect 230 3812 236 3813
rect 110 3809 116 3810
rect 110 3805 111 3809
rect 115 3805 116 3809
rect 230 3808 231 3812
rect 235 3808 236 3812
rect 230 3807 236 3808
rect 334 3812 340 3813
rect 334 3808 335 3812
rect 339 3808 340 3812
rect 334 3807 340 3808
rect 438 3812 444 3813
rect 438 3808 439 3812
rect 443 3808 444 3812
rect 438 3807 444 3808
rect 534 3812 540 3813
rect 534 3808 535 3812
rect 539 3808 540 3812
rect 534 3807 540 3808
rect 630 3812 636 3813
rect 630 3808 631 3812
rect 635 3808 636 3812
rect 630 3807 636 3808
rect 726 3812 732 3813
rect 726 3808 727 3812
rect 731 3808 732 3812
rect 726 3807 732 3808
rect 830 3812 836 3813
rect 830 3808 831 3812
rect 835 3808 836 3812
rect 830 3807 836 3808
rect 934 3812 940 3813
rect 934 3808 935 3812
rect 939 3808 940 3812
rect 934 3807 940 3808
rect 1038 3812 1044 3813
rect 1038 3808 1039 3812
rect 1043 3808 1044 3812
rect 1038 3807 1044 3808
rect 1150 3812 1156 3813
rect 1150 3808 1151 3812
rect 1155 3808 1156 3812
rect 1150 3807 1156 3808
rect 1262 3812 1268 3813
rect 1262 3808 1263 3812
rect 1267 3808 1268 3812
rect 1262 3807 1268 3808
rect 1382 3812 1388 3813
rect 1382 3808 1383 3812
rect 1387 3808 1388 3812
rect 1382 3807 1388 3808
rect 1502 3812 1508 3813
rect 1502 3808 1503 3812
rect 1507 3808 1508 3812
rect 1502 3807 1508 3808
rect 1630 3812 1636 3813
rect 1630 3808 1631 3812
rect 1635 3808 1636 3812
rect 1630 3807 1636 3808
rect 2006 3809 2012 3810
rect 110 3804 116 3805
rect 2006 3805 2007 3809
rect 2011 3805 2012 3809
rect 2006 3804 2012 3805
rect 230 3793 236 3794
rect 110 3792 116 3793
rect 110 3788 111 3792
rect 115 3788 116 3792
rect 230 3789 231 3793
rect 235 3789 236 3793
rect 230 3788 236 3789
rect 334 3793 340 3794
rect 334 3789 335 3793
rect 339 3789 340 3793
rect 334 3788 340 3789
rect 438 3793 444 3794
rect 438 3789 439 3793
rect 443 3789 444 3793
rect 438 3788 444 3789
rect 534 3793 540 3794
rect 534 3789 535 3793
rect 539 3789 540 3793
rect 534 3788 540 3789
rect 630 3793 636 3794
rect 630 3789 631 3793
rect 635 3789 636 3793
rect 630 3788 636 3789
rect 726 3793 732 3794
rect 726 3789 727 3793
rect 731 3789 732 3793
rect 726 3788 732 3789
rect 830 3793 836 3794
rect 830 3789 831 3793
rect 835 3789 836 3793
rect 830 3788 836 3789
rect 934 3793 940 3794
rect 934 3789 935 3793
rect 939 3789 940 3793
rect 934 3788 940 3789
rect 1038 3793 1044 3794
rect 1038 3789 1039 3793
rect 1043 3789 1044 3793
rect 1038 3788 1044 3789
rect 1150 3793 1156 3794
rect 1150 3789 1151 3793
rect 1155 3789 1156 3793
rect 1150 3788 1156 3789
rect 1262 3793 1268 3794
rect 1262 3789 1263 3793
rect 1267 3789 1268 3793
rect 1262 3788 1268 3789
rect 1382 3793 1388 3794
rect 1382 3789 1383 3793
rect 1387 3789 1388 3793
rect 1382 3788 1388 3789
rect 1502 3793 1508 3794
rect 1502 3789 1503 3793
rect 1507 3789 1508 3793
rect 1502 3788 1508 3789
rect 1630 3793 1636 3794
rect 1630 3789 1631 3793
rect 1635 3789 1636 3793
rect 1630 3788 1636 3789
rect 2006 3792 2012 3793
rect 2006 3788 2007 3792
rect 2011 3788 2012 3792
rect 110 3787 116 3788
rect 2006 3787 2012 3788
rect 2046 3752 2052 3753
rect 3942 3752 3948 3753
rect 2046 3748 2047 3752
rect 2051 3748 2052 3752
rect 2046 3747 2052 3748
rect 2070 3751 2076 3752
rect 2070 3747 2071 3751
rect 2075 3747 2076 3751
rect 2070 3746 2076 3747
rect 2182 3751 2188 3752
rect 2182 3747 2183 3751
rect 2187 3747 2188 3751
rect 2182 3746 2188 3747
rect 2326 3751 2332 3752
rect 2326 3747 2327 3751
rect 2331 3747 2332 3751
rect 2326 3746 2332 3747
rect 2478 3751 2484 3752
rect 2478 3747 2479 3751
rect 2483 3747 2484 3751
rect 2478 3746 2484 3747
rect 2638 3751 2644 3752
rect 2638 3747 2639 3751
rect 2643 3747 2644 3751
rect 2638 3746 2644 3747
rect 2806 3751 2812 3752
rect 2806 3747 2807 3751
rect 2811 3747 2812 3751
rect 2806 3746 2812 3747
rect 2982 3751 2988 3752
rect 2982 3747 2983 3751
rect 2987 3747 2988 3751
rect 2982 3746 2988 3747
rect 3158 3751 3164 3752
rect 3158 3747 3159 3751
rect 3163 3747 3164 3751
rect 3158 3746 3164 3747
rect 3334 3751 3340 3752
rect 3334 3747 3335 3751
rect 3339 3747 3340 3751
rect 3334 3746 3340 3747
rect 3510 3751 3516 3752
rect 3510 3747 3511 3751
rect 3515 3747 3516 3751
rect 3510 3746 3516 3747
rect 3686 3751 3692 3752
rect 3686 3747 3687 3751
rect 3691 3747 3692 3751
rect 3686 3746 3692 3747
rect 3838 3751 3844 3752
rect 3838 3747 3839 3751
rect 3843 3747 3844 3751
rect 3942 3748 3943 3752
rect 3947 3748 3948 3752
rect 3942 3747 3948 3748
rect 3838 3746 3844 3747
rect 110 3740 116 3741
rect 2006 3740 2012 3741
rect 110 3736 111 3740
rect 115 3736 116 3740
rect 110 3735 116 3736
rect 158 3739 164 3740
rect 158 3735 159 3739
rect 163 3735 164 3739
rect 158 3734 164 3735
rect 350 3739 356 3740
rect 350 3735 351 3739
rect 355 3735 356 3739
rect 350 3734 356 3735
rect 550 3739 556 3740
rect 550 3735 551 3739
rect 555 3735 556 3739
rect 550 3734 556 3735
rect 750 3739 756 3740
rect 750 3735 751 3739
rect 755 3735 756 3739
rect 750 3734 756 3735
rect 958 3739 964 3740
rect 958 3735 959 3739
rect 963 3735 964 3739
rect 958 3734 964 3735
rect 1166 3739 1172 3740
rect 1166 3735 1167 3739
rect 1171 3735 1172 3739
rect 1166 3734 1172 3735
rect 1382 3739 1388 3740
rect 1382 3735 1383 3739
rect 1387 3735 1388 3739
rect 1382 3734 1388 3735
rect 1606 3739 1612 3740
rect 1606 3735 1607 3739
rect 1611 3735 1612 3739
rect 2006 3736 2007 3740
rect 2011 3736 2012 3740
rect 2006 3735 2012 3736
rect 2046 3735 2052 3736
rect 1606 3734 1612 3735
rect 2046 3731 2047 3735
rect 2051 3731 2052 3735
rect 3942 3735 3948 3736
rect 2046 3730 2052 3731
rect 2070 3732 2076 3733
rect 2070 3728 2071 3732
rect 2075 3728 2076 3732
rect 2070 3727 2076 3728
rect 2182 3732 2188 3733
rect 2182 3728 2183 3732
rect 2187 3728 2188 3732
rect 2182 3727 2188 3728
rect 2326 3732 2332 3733
rect 2326 3728 2327 3732
rect 2331 3728 2332 3732
rect 2326 3727 2332 3728
rect 2478 3732 2484 3733
rect 2478 3728 2479 3732
rect 2483 3728 2484 3732
rect 2478 3727 2484 3728
rect 2638 3732 2644 3733
rect 2638 3728 2639 3732
rect 2643 3728 2644 3732
rect 2638 3727 2644 3728
rect 2806 3732 2812 3733
rect 2806 3728 2807 3732
rect 2811 3728 2812 3732
rect 2806 3727 2812 3728
rect 2982 3732 2988 3733
rect 2982 3728 2983 3732
rect 2987 3728 2988 3732
rect 2982 3727 2988 3728
rect 3158 3732 3164 3733
rect 3158 3728 3159 3732
rect 3163 3728 3164 3732
rect 3158 3727 3164 3728
rect 3334 3732 3340 3733
rect 3334 3728 3335 3732
rect 3339 3728 3340 3732
rect 3334 3727 3340 3728
rect 3510 3732 3516 3733
rect 3510 3728 3511 3732
rect 3515 3728 3516 3732
rect 3510 3727 3516 3728
rect 3686 3732 3692 3733
rect 3686 3728 3687 3732
rect 3691 3728 3692 3732
rect 3686 3727 3692 3728
rect 3838 3732 3844 3733
rect 3838 3728 3839 3732
rect 3843 3728 3844 3732
rect 3942 3731 3943 3735
rect 3947 3731 3948 3735
rect 3942 3730 3948 3731
rect 3838 3727 3844 3728
rect 110 3723 116 3724
rect 110 3719 111 3723
rect 115 3719 116 3723
rect 2006 3723 2012 3724
rect 110 3718 116 3719
rect 158 3720 164 3721
rect 158 3716 159 3720
rect 163 3716 164 3720
rect 158 3715 164 3716
rect 350 3720 356 3721
rect 350 3716 351 3720
rect 355 3716 356 3720
rect 350 3715 356 3716
rect 550 3720 556 3721
rect 550 3716 551 3720
rect 555 3716 556 3720
rect 550 3715 556 3716
rect 750 3720 756 3721
rect 750 3716 751 3720
rect 755 3716 756 3720
rect 750 3715 756 3716
rect 958 3720 964 3721
rect 958 3716 959 3720
rect 963 3716 964 3720
rect 958 3715 964 3716
rect 1166 3720 1172 3721
rect 1166 3716 1167 3720
rect 1171 3716 1172 3720
rect 1166 3715 1172 3716
rect 1382 3720 1388 3721
rect 1382 3716 1383 3720
rect 1387 3716 1388 3720
rect 1382 3715 1388 3716
rect 1606 3720 1612 3721
rect 1606 3716 1607 3720
rect 1611 3716 1612 3720
rect 2006 3719 2007 3723
rect 2011 3719 2012 3723
rect 2006 3718 2012 3719
rect 1606 3715 1612 3716
rect 2070 3660 2076 3661
rect 2046 3657 2052 3658
rect 2046 3653 2047 3657
rect 2051 3653 2052 3657
rect 2070 3656 2071 3660
rect 2075 3656 2076 3660
rect 2070 3655 2076 3656
rect 2198 3660 2204 3661
rect 2198 3656 2199 3660
rect 2203 3656 2204 3660
rect 2198 3655 2204 3656
rect 2366 3660 2372 3661
rect 2366 3656 2367 3660
rect 2371 3656 2372 3660
rect 2366 3655 2372 3656
rect 2550 3660 2556 3661
rect 2550 3656 2551 3660
rect 2555 3656 2556 3660
rect 2550 3655 2556 3656
rect 2734 3660 2740 3661
rect 2734 3656 2735 3660
rect 2739 3656 2740 3660
rect 2734 3655 2740 3656
rect 2926 3660 2932 3661
rect 2926 3656 2927 3660
rect 2931 3656 2932 3660
rect 2926 3655 2932 3656
rect 3110 3660 3116 3661
rect 3110 3656 3111 3660
rect 3115 3656 3116 3660
rect 3110 3655 3116 3656
rect 3294 3660 3300 3661
rect 3294 3656 3295 3660
rect 3299 3656 3300 3660
rect 3294 3655 3300 3656
rect 3478 3660 3484 3661
rect 3478 3656 3479 3660
rect 3483 3656 3484 3660
rect 3478 3655 3484 3656
rect 3670 3660 3676 3661
rect 3670 3656 3671 3660
rect 3675 3656 3676 3660
rect 3670 3655 3676 3656
rect 3838 3660 3844 3661
rect 3838 3656 3839 3660
rect 3843 3656 3844 3660
rect 3838 3655 3844 3656
rect 3942 3657 3948 3658
rect 150 3652 156 3653
rect 110 3649 116 3650
rect 110 3645 111 3649
rect 115 3645 116 3649
rect 150 3648 151 3652
rect 155 3648 156 3652
rect 150 3647 156 3648
rect 382 3652 388 3653
rect 382 3648 383 3652
rect 387 3648 388 3652
rect 382 3647 388 3648
rect 614 3652 620 3653
rect 614 3648 615 3652
rect 619 3648 620 3652
rect 614 3647 620 3648
rect 838 3652 844 3653
rect 838 3648 839 3652
rect 843 3648 844 3652
rect 838 3647 844 3648
rect 1054 3652 1060 3653
rect 1054 3648 1055 3652
rect 1059 3648 1060 3652
rect 1054 3647 1060 3648
rect 1262 3652 1268 3653
rect 1262 3648 1263 3652
rect 1267 3648 1268 3652
rect 1262 3647 1268 3648
rect 1478 3652 1484 3653
rect 1478 3648 1479 3652
rect 1483 3648 1484 3652
rect 1478 3647 1484 3648
rect 1694 3652 1700 3653
rect 2046 3652 2052 3653
rect 3942 3653 3943 3657
rect 3947 3653 3948 3657
rect 3942 3652 3948 3653
rect 1694 3648 1695 3652
rect 1699 3648 1700 3652
rect 1694 3647 1700 3648
rect 2006 3649 2012 3650
rect 110 3644 116 3645
rect 2006 3645 2007 3649
rect 2011 3645 2012 3649
rect 2006 3644 2012 3645
rect 2070 3641 2076 3642
rect 2046 3640 2052 3641
rect 2046 3636 2047 3640
rect 2051 3636 2052 3640
rect 2070 3637 2071 3641
rect 2075 3637 2076 3641
rect 2070 3636 2076 3637
rect 2198 3641 2204 3642
rect 2198 3637 2199 3641
rect 2203 3637 2204 3641
rect 2198 3636 2204 3637
rect 2366 3641 2372 3642
rect 2366 3637 2367 3641
rect 2371 3637 2372 3641
rect 2366 3636 2372 3637
rect 2550 3641 2556 3642
rect 2550 3637 2551 3641
rect 2555 3637 2556 3641
rect 2550 3636 2556 3637
rect 2734 3641 2740 3642
rect 2734 3637 2735 3641
rect 2739 3637 2740 3641
rect 2734 3636 2740 3637
rect 2926 3641 2932 3642
rect 2926 3637 2927 3641
rect 2931 3637 2932 3641
rect 2926 3636 2932 3637
rect 3110 3641 3116 3642
rect 3110 3637 3111 3641
rect 3115 3637 3116 3641
rect 3110 3636 3116 3637
rect 3294 3641 3300 3642
rect 3294 3637 3295 3641
rect 3299 3637 3300 3641
rect 3294 3636 3300 3637
rect 3478 3641 3484 3642
rect 3478 3637 3479 3641
rect 3483 3637 3484 3641
rect 3478 3636 3484 3637
rect 3670 3641 3676 3642
rect 3670 3637 3671 3641
rect 3675 3637 3676 3641
rect 3670 3636 3676 3637
rect 3838 3641 3844 3642
rect 3838 3637 3839 3641
rect 3843 3637 3844 3641
rect 3838 3636 3844 3637
rect 3942 3640 3948 3641
rect 3942 3636 3943 3640
rect 3947 3636 3948 3640
rect 2046 3635 2052 3636
rect 3942 3635 3948 3636
rect 150 3633 156 3634
rect 110 3632 116 3633
rect 110 3628 111 3632
rect 115 3628 116 3632
rect 150 3629 151 3633
rect 155 3629 156 3633
rect 150 3628 156 3629
rect 382 3633 388 3634
rect 382 3629 383 3633
rect 387 3629 388 3633
rect 382 3628 388 3629
rect 614 3633 620 3634
rect 614 3629 615 3633
rect 619 3629 620 3633
rect 614 3628 620 3629
rect 838 3633 844 3634
rect 838 3629 839 3633
rect 843 3629 844 3633
rect 838 3628 844 3629
rect 1054 3633 1060 3634
rect 1054 3629 1055 3633
rect 1059 3629 1060 3633
rect 1054 3628 1060 3629
rect 1262 3633 1268 3634
rect 1262 3629 1263 3633
rect 1267 3629 1268 3633
rect 1262 3628 1268 3629
rect 1478 3633 1484 3634
rect 1478 3629 1479 3633
rect 1483 3629 1484 3633
rect 1478 3628 1484 3629
rect 1694 3633 1700 3634
rect 1694 3629 1695 3633
rect 1699 3629 1700 3633
rect 1694 3628 1700 3629
rect 2006 3632 2012 3633
rect 2006 3628 2007 3632
rect 2011 3628 2012 3632
rect 110 3627 116 3628
rect 2006 3627 2012 3628
rect 2046 3584 2052 3585
rect 3942 3584 3948 3585
rect 2046 3580 2047 3584
rect 2051 3580 2052 3584
rect 2046 3579 2052 3580
rect 2102 3583 2108 3584
rect 2102 3579 2103 3583
rect 2107 3579 2108 3583
rect 2102 3578 2108 3579
rect 2278 3583 2284 3584
rect 2278 3579 2279 3583
rect 2283 3579 2284 3583
rect 2278 3578 2284 3579
rect 2470 3583 2476 3584
rect 2470 3579 2471 3583
rect 2475 3579 2476 3583
rect 2470 3578 2476 3579
rect 2670 3583 2676 3584
rect 2670 3579 2671 3583
rect 2675 3579 2676 3583
rect 2670 3578 2676 3579
rect 2870 3583 2876 3584
rect 2870 3579 2871 3583
rect 2875 3579 2876 3583
rect 2870 3578 2876 3579
rect 3062 3583 3068 3584
rect 3062 3579 3063 3583
rect 3067 3579 3068 3583
rect 3062 3578 3068 3579
rect 3254 3583 3260 3584
rect 3254 3579 3255 3583
rect 3259 3579 3260 3583
rect 3254 3578 3260 3579
rect 3446 3583 3452 3584
rect 3446 3579 3447 3583
rect 3451 3579 3452 3583
rect 3446 3578 3452 3579
rect 3638 3583 3644 3584
rect 3638 3579 3639 3583
rect 3643 3579 3644 3583
rect 3638 3578 3644 3579
rect 3838 3583 3844 3584
rect 3838 3579 3839 3583
rect 3843 3579 3844 3583
rect 3942 3580 3943 3584
rect 3947 3580 3948 3584
rect 3942 3579 3948 3580
rect 3838 3578 3844 3579
rect 110 3576 116 3577
rect 2006 3576 2012 3577
rect 110 3572 111 3576
rect 115 3572 116 3576
rect 110 3571 116 3572
rect 166 3575 172 3576
rect 166 3571 167 3575
rect 171 3571 172 3575
rect 166 3570 172 3571
rect 358 3575 364 3576
rect 358 3571 359 3575
rect 363 3571 364 3575
rect 358 3570 364 3571
rect 558 3575 564 3576
rect 558 3571 559 3575
rect 563 3571 564 3575
rect 558 3570 564 3571
rect 774 3575 780 3576
rect 774 3571 775 3575
rect 779 3571 780 3575
rect 774 3570 780 3571
rect 990 3575 996 3576
rect 990 3571 991 3575
rect 995 3571 996 3575
rect 990 3570 996 3571
rect 1214 3575 1220 3576
rect 1214 3571 1215 3575
rect 1219 3571 1220 3575
rect 1214 3570 1220 3571
rect 1446 3575 1452 3576
rect 1446 3571 1447 3575
rect 1451 3571 1452 3575
rect 1446 3570 1452 3571
rect 1686 3575 1692 3576
rect 1686 3571 1687 3575
rect 1691 3571 1692 3575
rect 2006 3572 2007 3576
rect 2011 3572 2012 3576
rect 2006 3571 2012 3572
rect 1686 3570 1692 3571
rect 2046 3567 2052 3568
rect 2046 3563 2047 3567
rect 2051 3563 2052 3567
rect 3942 3567 3948 3568
rect 2046 3562 2052 3563
rect 2102 3564 2108 3565
rect 2102 3560 2103 3564
rect 2107 3560 2108 3564
rect 110 3559 116 3560
rect 110 3555 111 3559
rect 115 3555 116 3559
rect 2006 3559 2012 3560
rect 2102 3559 2108 3560
rect 2278 3564 2284 3565
rect 2278 3560 2279 3564
rect 2283 3560 2284 3564
rect 2278 3559 2284 3560
rect 2470 3564 2476 3565
rect 2470 3560 2471 3564
rect 2475 3560 2476 3564
rect 2470 3559 2476 3560
rect 2670 3564 2676 3565
rect 2670 3560 2671 3564
rect 2675 3560 2676 3564
rect 2670 3559 2676 3560
rect 2870 3564 2876 3565
rect 2870 3560 2871 3564
rect 2875 3560 2876 3564
rect 2870 3559 2876 3560
rect 3062 3564 3068 3565
rect 3062 3560 3063 3564
rect 3067 3560 3068 3564
rect 3062 3559 3068 3560
rect 3254 3564 3260 3565
rect 3254 3560 3255 3564
rect 3259 3560 3260 3564
rect 3254 3559 3260 3560
rect 3446 3564 3452 3565
rect 3446 3560 3447 3564
rect 3451 3560 3452 3564
rect 3446 3559 3452 3560
rect 3638 3564 3644 3565
rect 3638 3560 3639 3564
rect 3643 3560 3644 3564
rect 3638 3559 3644 3560
rect 3838 3564 3844 3565
rect 3838 3560 3839 3564
rect 3843 3560 3844 3564
rect 3942 3563 3943 3567
rect 3947 3563 3948 3567
rect 3942 3562 3948 3563
rect 3838 3559 3844 3560
rect 110 3554 116 3555
rect 166 3556 172 3557
rect 166 3552 167 3556
rect 171 3552 172 3556
rect 166 3551 172 3552
rect 358 3556 364 3557
rect 358 3552 359 3556
rect 363 3552 364 3556
rect 358 3551 364 3552
rect 558 3556 564 3557
rect 558 3552 559 3556
rect 563 3552 564 3556
rect 558 3551 564 3552
rect 774 3556 780 3557
rect 774 3552 775 3556
rect 779 3552 780 3556
rect 774 3551 780 3552
rect 990 3556 996 3557
rect 990 3552 991 3556
rect 995 3552 996 3556
rect 990 3551 996 3552
rect 1214 3556 1220 3557
rect 1214 3552 1215 3556
rect 1219 3552 1220 3556
rect 1214 3551 1220 3552
rect 1446 3556 1452 3557
rect 1446 3552 1447 3556
rect 1451 3552 1452 3556
rect 1446 3551 1452 3552
rect 1686 3556 1692 3557
rect 1686 3552 1687 3556
rect 1691 3552 1692 3556
rect 2006 3555 2007 3559
rect 2011 3555 2012 3559
rect 2006 3554 2012 3555
rect 1686 3551 1692 3552
rect 2326 3500 2332 3501
rect 2046 3497 2052 3498
rect 2046 3493 2047 3497
rect 2051 3493 2052 3497
rect 2326 3496 2327 3500
rect 2331 3496 2332 3500
rect 2326 3495 2332 3496
rect 2446 3500 2452 3501
rect 2446 3496 2447 3500
rect 2451 3496 2452 3500
rect 2446 3495 2452 3496
rect 2582 3500 2588 3501
rect 2582 3496 2583 3500
rect 2587 3496 2588 3500
rect 2582 3495 2588 3496
rect 2734 3500 2740 3501
rect 2734 3496 2735 3500
rect 2739 3496 2740 3500
rect 2734 3495 2740 3496
rect 2910 3500 2916 3501
rect 2910 3496 2911 3500
rect 2915 3496 2916 3500
rect 2910 3495 2916 3496
rect 3110 3500 3116 3501
rect 3110 3496 3111 3500
rect 3115 3496 3116 3500
rect 3110 3495 3116 3496
rect 3334 3500 3340 3501
rect 3334 3496 3335 3500
rect 3339 3496 3340 3500
rect 3334 3495 3340 3496
rect 3566 3500 3572 3501
rect 3566 3496 3567 3500
rect 3571 3496 3572 3500
rect 3566 3495 3572 3496
rect 3806 3500 3812 3501
rect 3806 3496 3807 3500
rect 3811 3496 3812 3500
rect 3806 3495 3812 3496
rect 3942 3497 3948 3498
rect 2046 3492 2052 3493
rect 3942 3493 3943 3497
rect 3947 3493 3948 3497
rect 3942 3492 3948 3493
rect 294 3488 300 3489
rect 110 3485 116 3486
rect 110 3481 111 3485
rect 115 3481 116 3485
rect 294 3484 295 3488
rect 299 3484 300 3488
rect 294 3483 300 3484
rect 430 3488 436 3489
rect 430 3484 431 3488
rect 435 3484 436 3488
rect 430 3483 436 3484
rect 582 3488 588 3489
rect 582 3484 583 3488
rect 587 3484 588 3488
rect 582 3483 588 3484
rect 742 3488 748 3489
rect 742 3484 743 3488
rect 747 3484 748 3488
rect 742 3483 748 3484
rect 910 3488 916 3489
rect 910 3484 911 3488
rect 915 3484 916 3488
rect 910 3483 916 3484
rect 1078 3488 1084 3489
rect 1078 3484 1079 3488
rect 1083 3484 1084 3488
rect 1078 3483 1084 3484
rect 1246 3488 1252 3489
rect 1246 3484 1247 3488
rect 1251 3484 1252 3488
rect 1246 3483 1252 3484
rect 1422 3488 1428 3489
rect 1422 3484 1423 3488
rect 1427 3484 1428 3488
rect 1422 3483 1428 3484
rect 1598 3488 1604 3489
rect 1598 3484 1599 3488
rect 1603 3484 1604 3488
rect 1598 3483 1604 3484
rect 1774 3488 1780 3489
rect 1774 3484 1775 3488
rect 1779 3484 1780 3488
rect 1774 3483 1780 3484
rect 2006 3485 2012 3486
rect 110 3480 116 3481
rect 2006 3481 2007 3485
rect 2011 3481 2012 3485
rect 2326 3481 2332 3482
rect 2006 3480 2012 3481
rect 2046 3480 2052 3481
rect 2046 3476 2047 3480
rect 2051 3476 2052 3480
rect 2326 3477 2327 3481
rect 2331 3477 2332 3481
rect 2326 3476 2332 3477
rect 2446 3481 2452 3482
rect 2446 3477 2447 3481
rect 2451 3477 2452 3481
rect 2446 3476 2452 3477
rect 2582 3481 2588 3482
rect 2582 3477 2583 3481
rect 2587 3477 2588 3481
rect 2582 3476 2588 3477
rect 2734 3481 2740 3482
rect 2734 3477 2735 3481
rect 2739 3477 2740 3481
rect 2734 3476 2740 3477
rect 2910 3481 2916 3482
rect 2910 3477 2911 3481
rect 2915 3477 2916 3481
rect 2910 3476 2916 3477
rect 3110 3481 3116 3482
rect 3110 3477 3111 3481
rect 3115 3477 3116 3481
rect 3110 3476 3116 3477
rect 3334 3481 3340 3482
rect 3334 3477 3335 3481
rect 3339 3477 3340 3481
rect 3334 3476 3340 3477
rect 3566 3481 3572 3482
rect 3566 3477 3567 3481
rect 3571 3477 3572 3481
rect 3566 3476 3572 3477
rect 3806 3481 3812 3482
rect 3806 3477 3807 3481
rect 3811 3477 3812 3481
rect 3806 3476 3812 3477
rect 3942 3480 3948 3481
rect 3942 3476 3943 3480
rect 3947 3476 3948 3480
rect 2046 3475 2052 3476
rect 3942 3475 3948 3476
rect 294 3469 300 3470
rect 110 3468 116 3469
rect 110 3464 111 3468
rect 115 3464 116 3468
rect 294 3465 295 3469
rect 299 3465 300 3469
rect 294 3464 300 3465
rect 430 3469 436 3470
rect 430 3465 431 3469
rect 435 3465 436 3469
rect 430 3464 436 3465
rect 582 3469 588 3470
rect 582 3465 583 3469
rect 587 3465 588 3469
rect 582 3464 588 3465
rect 742 3469 748 3470
rect 742 3465 743 3469
rect 747 3465 748 3469
rect 742 3464 748 3465
rect 910 3469 916 3470
rect 910 3465 911 3469
rect 915 3465 916 3469
rect 910 3464 916 3465
rect 1078 3469 1084 3470
rect 1078 3465 1079 3469
rect 1083 3465 1084 3469
rect 1078 3464 1084 3465
rect 1246 3469 1252 3470
rect 1246 3465 1247 3469
rect 1251 3465 1252 3469
rect 1246 3464 1252 3465
rect 1422 3469 1428 3470
rect 1422 3465 1423 3469
rect 1427 3465 1428 3469
rect 1422 3464 1428 3465
rect 1598 3469 1604 3470
rect 1598 3465 1599 3469
rect 1603 3465 1604 3469
rect 1598 3464 1604 3465
rect 1774 3469 1780 3470
rect 1774 3465 1775 3469
rect 1779 3465 1780 3469
rect 1774 3464 1780 3465
rect 2006 3468 2012 3469
rect 2006 3464 2007 3468
rect 2011 3464 2012 3468
rect 110 3463 116 3464
rect 2006 3463 2012 3464
rect 2046 3428 2052 3429
rect 3942 3428 3948 3429
rect 2046 3424 2047 3428
rect 2051 3424 2052 3428
rect 2046 3423 2052 3424
rect 2446 3427 2452 3428
rect 2446 3423 2447 3427
rect 2451 3423 2452 3427
rect 2446 3422 2452 3423
rect 2550 3427 2556 3428
rect 2550 3423 2551 3427
rect 2555 3423 2556 3427
rect 2550 3422 2556 3423
rect 2662 3427 2668 3428
rect 2662 3423 2663 3427
rect 2667 3423 2668 3427
rect 2662 3422 2668 3423
rect 2774 3427 2780 3428
rect 2774 3423 2775 3427
rect 2779 3423 2780 3427
rect 2774 3422 2780 3423
rect 2902 3427 2908 3428
rect 2902 3423 2903 3427
rect 2907 3423 2908 3427
rect 2902 3422 2908 3423
rect 3046 3427 3052 3428
rect 3046 3423 3047 3427
rect 3051 3423 3052 3427
rect 3046 3422 3052 3423
rect 3206 3427 3212 3428
rect 3206 3423 3207 3427
rect 3211 3423 3212 3427
rect 3206 3422 3212 3423
rect 3382 3427 3388 3428
rect 3382 3423 3383 3427
rect 3387 3423 3388 3427
rect 3382 3422 3388 3423
rect 3566 3427 3572 3428
rect 3566 3423 3567 3427
rect 3571 3423 3572 3427
rect 3566 3422 3572 3423
rect 3750 3427 3756 3428
rect 3750 3423 3751 3427
rect 3755 3423 3756 3427
rect 3942 3424 3943 3428
rect 3947 3424 3948 3428
rect 3942 3423 3948 3424
rect 3750 3422 3756 3423
rect 2046 3411 2052 3412
rect 2046 3407 2047 3411
rect 2051 3407 2052 3411
rect 3942 3411 3948 3412
rect 2046 3406 2052 3407
rect 2446 3408 2452 3409
rect 2446 3404 2447 3408
rect 2451 3404 2452 3408
rect 2446 3403 2452 3404
rect 2550 3408 2556 3409
rect 2550 3404 2551 3408
rect 2555 3404 2556 3408
rect 2550 3403 2556 3404
rect 2662 3408 2668 3409
rect 2662 3404 2663 3408
rect 2667 3404 2668 3408
rect 2662 3403 2668 3404
rect 2774 3408 2780 3409
rect 2774 3404 2775 3408
rect 2779 3404 2780 3408
rect 2774 3403 2780 3404
rect 2902 3408 2908 3409
rect 2902 3404 2903 3408
rect 2907 3404 2908 3408
rect 2902 3403 2908 3404
rect 3046 3408 3052 3409
rect 3046 3404 3047 3408
rect 3051 3404 3052 3408
rect 3046 3403 3052 3404
rect 3206 3408 3212 3409
rect 3206 3404 3207 3408
rect 3211 3404 3212 3408
rect 3206 3403 3212 3404
rect 3382 3408 3388 3409
rect 3382 3404 3383 3408
rect 3387 3404 3388 3408
rect 3382 3403 3388 3404
rect 3566 3408 3572 3409
rect 3566 3404 3567 3408
rect 3571 3404 3572 3408
rect 3566 3403 3572 3404
rect 3750 3408 3756 3409
rect 3750 3404 3751 3408
rect 3755 3404 3756 3408
rect 3942 3407 3943 3411
rect 3947 3407 3948 3411
rect 3942 3406 3948 3407
rect 3750 3403 3756 3404
rect 110 3396 116 3397
rect 2006 3396 2012 3397
rect 110 3392 111 3396
rect 115 3392 116 3396
rect 110 3391 116 3392
rect 494 3395 500 3396
rect 494 3391 495 3395
rect 499 3391 500 3395
rect 494 3390 500 3391
rect 646 3395 652 3396
rect 646 3391 647 3395
rect 651 3391 652 3395
rect 646 3390 652 3391
rect 798 3395 804 3396
rect 798 3391 799 3395
rect 803 3391 804 3395
rect 798 3390 804 3391
rect 958 3395 964 3396
rect 958 3391 959 3395
rect 963 3391 964 3395
rect 958 3390 964 3391
rect 1126 3395 1132 3396
rect 1126 3391 1127 3395
rect 1131 3391 1132 3395
rect 1126 3390 1132 3391
rect 1294 3395 1300 3396
rect 1294 3391 1295 3395
rect 1299 3391 1300 3395
rect 1294 3390 1300 3391
rect 1462 3395 1468 3396
rect 1462 3391 1463 3395
rect 1467 3391 1468 3395
rect 1462 3390 1468 3391
rect 1638 3395 1644 3396
rect 1638 3391 1639 3395
rect 1643 3391 1644 3395
rect 1638 3390 1644 3391
rect 1814 3395 1820 3396
rect 1814 3391 1815 3395
rect 1819 3391 1820 3395
rect 2006 3392 2007 3396
rect 2011 3392 2012 3396
rect 2006 3391 2012 3392
rect 1814 3390 1820 3391
rect 110 3379 116 3380
rect 110 3375 111 3379
rect 115 3375 116 3379
rect 2006 3379 2012 3380
rect 110 3374 116 3375
rect 494 3376 500 3377
rect 494 3372 495 3376
rect 499 3372 500 3376
rect 494 3371 500 3372
rect 646 3376 652 3377
rect 646 3372 647 3376
rect 651 3372 652 3376
rect 646 3371 652 3372
rect 798 3376 804 3377
rect 798 3372 799 3376
rect 803 3372 804 3376
rect 798 3371 804 3372
rect 958 3376 964 3377
rect 958 3372 959 3376
rect 963 3372 964 3376
rect 958 3371 964 3372
rect 1126 3376 1132 3377
rect 1126 3372 1127 3376
rect 1131 3372 1132 3376
rect 1126 3371 1132 3372
rect 1294 3376 1300 3377
rect 1294 3372 1295 3376
rect 1299 3372 1300 3376
rect 1294 3371 1300 3372
rect 1462 3376 1468 3377
rect 1462 3372 1463 3376
rect 1467 3372 1468 3376
rect 1462 3371 1468 3372
rect 1638 3376 1644 3377
rect 1638 3372 1639 3376
rect 1643 3372 1644 3376
rect 1638 3371 1644 3372
rect 1814 3376 1820 3377
rect 1814 3372 1815 3376
rect 1819 3372 1820 3376
rect 2006 3375 2007 3379
rect 2011 3375 2012 3379
rect 2006 3374 2012 3375
rect 1814 3371 1820 3372
rect 2566 3336 2572 3337
rect 2046 3333 2052 3334
rect 2046 3329 2047 3333
rect 2051 3329 2052 3333
rect 2566 3332 2567 3336
rect 2571 3332 2572 3336
rect 2566 3331 2572 3332
rect 2718 3336 2724 3337
rect 2718 3332 2719 3336
rect 2723 3332 2724 3336
rect 2718 3331 2724 3332
rect 2870 3336 2876 3337
rect 2870 3332 2871 3336
rect 2875 3332 2876 3336
rect 2870 3331 2876 3332
rect 3022 3336 3028 3337
rect 3022 3332 3023 3336
rect 3027 3332 3028 3336
rect 3022 3331 3028 3332
rect 3174 3336 3180 3337
rect 3174 3332 3175 3336
rect 3179 3332 3180 3336
rect 3174 3331 3180 3332
rect 3326 3336 3332 3337
rect 3326 3332 3327 3336
rect 3331 3332 3332 3336
rect 3326 3331 3332 3332
rect 3478 3336 3484 3337
rect 3478 3332 3479 3336
rect 3483 3332 3484 3336
rect 3478 3331 3484 3332
rect 3630 3336 3636 3337
rect 3630 3332 3631 3336
rect 3635 3332 3636 3336
rect 3630 3331 3636 3332
rect 3782 3336 3788 3337
rect 3782 3332 3783 3336
rect 3787 3332 3788 3336
rect 3782 3331 3788 3332
rect 3942 3333 3948 3334
rect 2046 3328 2052 3329
rect 3942 3329 3943 3333
rect 3947 3329 3948 3333
rect 3942 3328 3948 3329
rect 2566 3317 2572 3318
rect 2046 3316 2052 3317
rect 2046 3312 2047 3316
rect 2051 3312 2052 3316
rect 2566 3313 2567 3317
rect 2571 3313 2572 3317
rect 2566 3312 2572 3313
rect 2718 3317 2724 3318
rect 2718 3313 2719 3317
rect 2723 3313 2724 3317
rect 2718 3312 2724 3313
rect 2870 3317 2876 3318
rect 2870 3313 2871 3317
rect 2875 3313 2876 3317
rect 2870 3312 2876 3313
rect 3022 3317 3028 3318
rect 3022 3313 3023 3317
rect 3027 3313 3028 3317
rect 3022 3312 3028 3313
rect 3174 3317 3180 3318
rect 3174 3313 3175 3317
rect 3179 3313 3180 3317
rect 3174 3312 3180 3313
rect 3326 3317 3332 3318
rect 3326 3313 3327 3317
rect 3331 3313 3332 3317
rect 3326 3312 3332 3313
rect 3478 3317 3484 3318
rect 3478 3313 3479 3317
rect 3483 3313 3484 3317
rect 3478 3312 3484 3313
rect 3630 3317 3636 3318
rect 3630 3313 3631 3317
rect 3635 3313 3636 3317
rect 3630 3312 3636 3313
rect 3782 3317 3788 3318
rect 3782 3313 3783 3317
rect 3787 3313 3788 3317
rect 3782 3312 3788 3313
rect 3942 3316 3948 3317
rect 3942 3312 3943 3316
rect 3947 3312 3948 3316
rect 2046 3311 2052 3312
rect 3942 3311 3948 3312
rect 134 3304 140 3305
rect 110 3301 116 3302
rect 110 3297 111 3301
rect 115 3297 116 3301
rect 134 3300 135 3304
rect 139 3300 140 3304
rect 134 3299 140 3300
rect 294 3304 300 3305
rect 294 3300 295 3304
rect 299 3300 300 3304
rect 294 3299 300 3300
rect 478 3304 484 3305
rect 478 3300 479 3304
rect 483 3300 484 3304
rect 478 3299 484 3300
rect 670 3304 676 3305
rect 670 3300 671 3304
rect 675 3300 676 3304
rect 670 3299 676 3300
rect 862 3304 868 3305
rect 862 3300 863 3304
rect 867 3300 868 3304
rect 862 3299 868 3300
rect 1054 3304 1060 3305
rect 1054 3300 1055 3304
rect 1059 3300 1060 3304
rect 1054 3299 1060 3300
rect 1246 3304 1252 3305
rect 1246 3300 1247 3304
rect 1251 3300 1252 3304
rect 1246 3299 1252 3300
rect 1438 3304 1444 3305
rect 1438 3300 1439 3304
rect 1443 3300 1444 3304
rect 1438 3299 1444 3300
rect 1630 3304 1636 3305
rect 1630 3300 1631 3304
rect 1635 3300 1636 3304
rect 1630 3299 1636 3300
rect 1822 3304 1828 3305
rect 1822 3300 1823 3304
rect 1827 3300 1828 3304
rect 1822 3299 1828 3300
rect 2006 3301 2012 3302
rect 110 3296 116 3297
rect 2006 3297 2007 3301
rect 2011 3297 2012 3301
rect 2006 3296 2012 3297
rect 134 3285 140 3286
rect 110 3284 116 3285
rect 110 3280 111 3284
rect 115 3280 116 3284
rect 134 3281 135 3285
rect 139 3281 140 3285
rect 134 3280 140 3281
rect 294 3285 300 3286
rect 294 3281 295 3285
rect 299 3281 300 3285
rect 294 3280 300 3281
rect 478 3285 484 3286
rect 478 3281 479 3285
rect 483 3281 484 3285
rect 478 3280 484 3281
rect 670 3285 676 3286
rect 670 3281 671 3285
rect 675 3281 676 3285
rect 670 3280 676 3281
rect 862 3285 868 3286
rect 862 3281 863 3285
rect 867 3281 868 3285
rect 862 3280 868 3281
rect 1054 3285 1060 3286
rect 1054 3281 1055 3285
rect 1059 3281 1060 3285
rect 1054 3280 1060 3281
rect 1246 3285 1252 3286
rect 1246 3281 1247 3285
rect 1251 3281 1252 3285
rect 1246 3280 1252 3281
rect 1438 3285 1444 3286
rect 1438 3281 1439 3285
rect 1443 3281 1444 3285
rect 1438 3280 1444 3281
rect 1630 3285 1636 3286
rect 1630 3281 1631 3285
rect 1635 3281 1636 3285
rect 1630 3280 1636 3281
rect 1822 3285 1828 3286
rect 1822 3281 1823 3285
rect 1827 3281 1828 3285
rect 1822 3280 1828 3281
rect 2006 3284 2012 3285
rect 2006 3280 2007 3284
rect 2011 3280 2012 3284
rect 110 3279 116 3280
rect 2006 3279 2012 3280
rect 2046 3260 2052 3261
rect 3942 3260 3948 3261
rect 2046 3256 2047 3260
rect 2051 3256 2052 3260
rect 2046 3255 2052 3256
rect 2414 3259 2420 3260
rect 2414 3255 2415 3259
rect 2419 3255 2420 3259
rect 2414 3254 2420 3255
rect 2550 3259 2556 3260
rect 2550 3255 2551 3259
rect 2555 3255 2556 3259
rect 2550 3254 2556 3255
rect 2686 3259 2692 3260
rect 2686 3255 2687 3259
rect 2691 3255 2692 3259
rect 2686 3254 2692 3255
rect 2830 3259 2836 3260
rect 2830 3255 2831 3259
rect 2835 3255 2836 3259
rect 2830 3254 2836 3255
rect 2974 3259 2980 3260
rect 2974 3255 2975 3259
rect 2979 3255 2980 3259
rect 2974 3254 2980 3255
rect 3118 3259 3124 3260
rect 3118 3255 3119 3259
rect 3123 3255 3124 3259
rect 3118 3254 3124 3255
rect 3254 3259 3260 3260
rect 3254 3255 3255 3259
rect 3259 3255 3260 3259
rect 3254 3254 3260 3255
rect 3382 3259 3388 3260
rect 3382 3255 3383 3259
rect 3387 3255 3388 3259
rect 3382 3254 3388 3255
rect 3502 3259 3508 3260
rect 3502 3255 3503 3259
rect 3507 3255 3508 3259
rect 3502 3254 3508 3255
rect 3622 3259 3628 3260
rect 3622 3255 3623 3259
rect 3627 3255 3628 3259
rect 3622 3254 3628 3255
rect 3742 3259 3748 3260
rect 3742 3255 3743 3259
rect 3747 3255 3748 3259
rect 3742 3254 3748 3255
rect 3838 3259 3844 3260
rect 3838 3255 3839 3259
rect 3843 3255 3844 3259
rect 3942 3256 3943 3260
rect 3947 3256 3948 3260
rect 3942 3255 3948 3256
rect 3838 3254 3844 3255
rect 2046 3243 2052 3244
rect 2046 3239 2047 3243
rect 2051 3239 2052 3243
rect 3942 3243 3948 3244
rect 2046 3238 2052 3239
rect 2414 3240 2420 3241
rect 2414 3236 2415 3240
rect 2419 3236 2420 3240
rect 2414 3235 2420 3236
rect 2550 3240 2556 3241
rect 2550 3236 2551 3240
rect 2555 3236 2556 3240
rect 2550 3235 2556 3236
rect 2686 3240 2692 3241
rect 2686 3236 2687 3240
rect 2691 3236 2692 3240
rect 2686 3235 2692 3236
rect 2830 3240 2836 3241
rect 2830 3236 2831 3240
rect 2835 3236 2836 3240
rect 2830 3235 2836 3236
rect 2974 3240 2980 3241
rect 2974 3236 2975 3240
rect 2979 3236 2980 3240
rect 2974 3235 2980 3236
rect 3118 3240 3124 3241
rect 3118 3236 3119 3240
rect 3123 3236 3124 3240
rect 3118 3235 3124 3236
rect 3254 3240 3260 3241
rect 3254 3236 3255 3240
rect 3259 3236 3260 3240
rect 3254 3235 3260 3236
rect 3382 3240 3388 3241
rect 3382 3236 3383 3240
rect 3387 3236 3388 3240
rect 3382 3235 3388 3236
rect 3502 3240 3508 3241
rect 3502 3236 3503 3240
rect 3507 3236 3508 3240
rect 3502 3235 3508 3236
rect 3622 3240 3628 3241
rect 3622 3236 3623 3240
rect 3627 3236 3628 3240
rect 3622 3235 3628 3236
rect 3742 3240 3748 3241
rect 3742 3236 3743 3240
rect 3747 3236 3748 3240
rect 3742 3235 3748 3236
rect 3838 3240 3844 3241
rect 3838 3236 3839 3240
rect 3843 3236 3844 3240
rect 3942 3239 3943 3243
rect 3947 3239 3948 3243
rect 3942 3238 3948 3239
rect 3838 3235 3844 3236
rect 110 3228 116 3229
rect 2006 3228 2012 3229
rect 110 3224 111 3228
rect 115 3224 116 3228
rect 110 3223 116 3224
rect 134 3227 140 3228
rect 134 3223 135 3227
rect 139 3223 140 3227
rect 134 3222 140 3223
rect 318 3227 324 3228
rect 318 3223 319 3227
rect 323 3223 324 3227
rect 318 3222 324 3223
rect 518 3227 524 3228
rect 518 3223 519 3227
rect 523 3223 524 3227
rect 518 3222 524 3223
rect 718 3227 724 3228
rect 718 3223 719 3227
rect 723 3223 724 3227
rect 718 3222 724 3223
rect 910 3227 916 3228
rect 910 3223 911 3227
rect 915 3223 916 3227
rect 910 3222 916 3223
rect 1094 3227 1100 3228
rect 1094 3223 1095 3227
rect 1099 3223 1100 3227
rect 1094 3222 1100 3223
rect 1270 3227 1276 3228
rect 1270 3223 1271 3227
rect 1275 3223 1276 3227
rect 1270 3222 1276 3223
rect 1446 3227 1452 3228
rect 1446 3223 1447 3227
rect 1451 3223 1452 3227
rect 1446 3222 1452 3223
rect 1622 3227 1628 3228
rect 1622 3223 1623 3227
rect 1627 3223 1628 3227
rect 1622 3222 1628 3223
rect 1798 3227 1804 3228
rect 1798 3223 1799 3227
rect 1803 3223 1804 3227
rect 2006 3224 2007 3228
rect 2011 3224 2012 3228
rect 2006 3223 2012 3224
rect 1798 3222 1804 3223
rect 110 3211 116 3212
rect 110 3207 111 3211
rect 115 3207 116 3211
rect 2006 3211 2012 3212
rect 110 3206 116 3207
rect 134 3208 140 3209
rect 134 3204 135 3208
rect 139 3204 140 3208
rect 134 3203 140 3204
rect 318 3208 324 3209
rect 318 3204 319 3208
rect 323 3204 324 3208
rect 318 3203 324 3204
rect 518 3208 524 3209
rect 518 3204 519 3208
rect 523 3204 524 3208
rect 518 3203 524 3204
rect 718 3208 724 3209
rect 718 3204 719 3208
rect 723 3204 724 3208
rect 718 3203 724 3204
rect 910 3208 916 3209
rect 910 3204 911 3208
rect 915 3204 916 3208
rect 910 3203 916 3204
rect 1094 3208 1100 3209
rect 1094 3204 1095 3208
rect 1099 3204 1100 3208
rect 1094 3203 1100 3204
rect 1270 3208 1276 3209
rect 1270 3204 1271 3208
rect 1275 3204 1276 3208
rect 1270 3203 1276 3204
rect 1446 3208 1452 3209
rect 1446 3204 1447 3208
rect 1451 3204 1452 3208
rect 1446 3203 1452 3204
rect 1622 3208 1628 3209
rect 1622 3204 1623 3208
rect 1627 3204 1628 3208
rect 1622 3203 1628 3204
rect 1798 3208 1804 3209
rect 1798 3204 1799 3208
rect 1803 3204 1804 3208
rect 2006 3207 2007 3211
rect 2011 3207 2012 3211
rect 2006 3206 2012 3207
rect 1798 3203 1804 3204
rect 2246 3168 2252 3169
rect 2046 3165 2052 3166
rect 2046 3161 2047 3165
rect 2051 3161 2052 3165
rect 2246 3164 2247 3168
rect 2251 3164 2252 3168
rect 2246 3163 2252 3164
rect 2398 3168 2404 3169
rect 2398 3164 2399 3168
rect 2403 3164 2404 3168
rect 2398 3163 2404 3164
rect 2558 3168 2564 3169
rect 2558 3164 2559 3168
rect 2563 3164 2564 3168
rect 2558 3163 2564 3164
rect 2726 3168 2732 3169
rect 2726 3164 2727 3168
rect 2731 3164 2732 3168
rect 2726 3163 2732 3164
rect 2902 3168 2908 3169
rect 2902 3164 2903 3168
rect 2907 3164 2908 3168
rect 2902 3163 2908 3164
rect 3078 3168 3084 3169
rect 3078 3164 3079 3168
rect 3083 3164 3084 3168
rect 3078 3163 3084 3164
rect 3262 3168 3268 3169
rect 3262 3164 3263 3168
rect 3267 3164 3268 3168
rect 3262 3163 3268 3164
rect 3446 3168 3452 3169
rect 3446 3164 3447 3168
rect 3451 3164 3452 3168
rect 3446 3163 3452 3164
rect 3630 3168 3636 3169
rect 3630 3164 3631 3168
rect 3635 3164 3636 3168
rect 3630 3163 3636 3164
rect 3814 3168 3820 3169
rect 3814 3164 3815 3168
rect 3819 3164 3820 3168
rect 3814 3163 3820 3164
rect 3942 3165 3948 3166
rect 2046 3160 2052 3161
rect 3942 3161 3943 3165
rect 3947 3161 3948 3165
rect 3942 3160 3948 3161
rect 2246 3149 2252 3150
rect 2046 3148 2052 3149
rect 2046 3144 2047 3148
rect 2051 3144 2052 3148
rect 2246 3145 2247 3149
rect 2251 3145 2252 3149
rect 2246 3144 2252 3145
rect 2398 3149 2404 3150
rect 2398 3145 2399 3149
rect 2403 3145 2404 3149
rect 2398 3144 2404 3145
rect 2558 3149 2564 3150
rect 2558 3145 2559 3149
rect 2563 3145 2564 3149
rect 2558 3144 2564 3145
rect 2726 3149 2732 3150
rect 2726 3145 2727 3149
rect 2731 3145 2732 3149
rect 2726 3144 2732 3145
rect 2902 3149 2908 3150
rect 2902 3145 2903 3149
rect 2907 3145 2908 3149
rect 2902 3144 2908 3145
rect 3078 3149 3084 3150
rect 3078 3145 3079 3149
rect 3083 3145 3084 3149
rect 3078 3144 3084 3145
rect 3262 3149 3268 3150
rect 3262 3145 3263 3149
rect 3267 3145 3268 3149
rect 3262 3144 3268 3145
rect 3446 3149 3452 3150
rect 3446 3145 3447 3149
rect 3451 3145 3452 3149
rect 3446 3144 3452 3145
rect 3630 3149 3636 3150
rect 3630 3145 3631 3149
rect 3635 3145 3636 3149
rect 3630 3144 3636 3145
rect 3814 3149 3820 3150
rect 3814 3145 3815 3149
rect 3819 3145 3820 3149
rect 3814 3144 3820 3145
rect 3942 3148 3948 3149
rect 3942 3144 3943 3148
rect 3947 3144 3948 3148
rect 2046 3143 2052 3144
rect 3942 3143 3948 3144
rect 142 3140 148 3141
rect 110 3137 116 3138
rect 110 3133 111 3137
rect 115 3133 116 3137
rect 142 3136 143 3140
rect 147 3136 148 3140
rect 142 3135 148 3136
rect 342 3140 348 3141
rect 342 3136 343 3140
rect 347 3136 348 3140
rect 342 3135 348 3136
rect 542 3140 548 3141
rect 542 3136 543 3140
rect 547 3136 548 3140
rect 542 3135 548 3136
rect 742 3140 748 3141
rect 742 3136 743 3140
rect 747 3136 748 3140
rect 742 3135 748 3136
rect 926 3140 932 3141
rect 926 3136 927 3140
rect 931 3136 932 3140
rect 926 3135 932 3136
rect 1102 3140 1108 3141
rect 1102 3136 1103 3140
rect 1107 3136 1108 3140
rect 1102 3135 1108 3136
rect 1262 3140 1268 3141
rect 1262 3136 1263 3140
rect 1267 3136 1268 3140
rect 1262 3135 1268 3136
rect 1422 3140 1428 3141
rect 1422 3136 1423 3140
rect 1427 3136 1428 3140
rect 1422 3135 1428 3136
rect 1574 3140 1580 3141
rect 1574 3136 1575 3140
rect 1579 3136 1580 3140
rect 1574 3135 1580 3136
rect 1734 3140 1740 3141
rect 1734 3136 1735 3140
rect 1739 3136 1740 3140
rect 1734 3135 1740 3136
rect 2006 3137 2012 3138
rect 110 3132 116 3133
rect 2006 3133 2007 3137
rect 2011 3133 2012 3137
rect 2006 3132 2012 3133
rect 142 3121 148 3122
rect 110 3120 116 3121
rect 110 3116 111 3120
rect 115 3116 116 3120
rect 142 3117 143 3121
rect 147 3117 148 3121
rect 142 3116 148 3117
rect 342 3121 348 3122
rect 342 3117 343 3121
rect 347 3117 348 3121
rect 342 3116 348 3117
rect 542 3121 548 3122
rect 542 3117 543 3121
rect 547 3117 548 3121
rect 542 3116 548 3117
rect 742 3121 748 3122
rect 742 3117 743 3121
rect 747 3117 748 3121
rect 742 3116 748 3117
rect 926 3121 932 3122
rect 926 3117 927 3121
rect 931 3117 932 3121
rect 926 3116 932 3117
rect 1102 3121 1108 3122
rect 1102 3117 1103 3121
rect 1107 3117 1108 3121
rect 1102 3116 1108 3117
rect 1262 3121 1268 3122
rect 1262 3117 1263 3121
rect 1267 3117 1268 3121
rect 1262 3116 1268 3117
rect 1422 3121 1428 3122
rect 1422 3117 1423 3121
rect 1427 3117 1428 3121
rect 1422 3116 1428 3117
rect 1574 3121 1580 3122
rect 1574 3117 1575 3121
rect 1579 3117 1580 3121
rect 1574 3116 1580 3117
rect 1734 3121 1740 3122
rect 1734 3117 1735 3121
rect 1739 3117 1740 3121
rect 1734 3116 1740 3117
rect 2006 3120 2012 3121
rect 2006 3116 2007 3120
rect 2011 3116 2012 3120
rect 110 3115 116 3116
rect 2006 3115 2012 3116
rect 2046 3092 2052 3093
rect 3942 3092 3948 3093
rect 2046 3088 2047 3092
rect 2051 3088 2052 3092
rect 2046 3087 2052 3088
rect 2078 3091 2084 3092
rect 2078 3087 2079 3091
rect 2083 3087 2084 3091
rect 2078 3086 2084 3087
rect 2222 3091 2228 3092
rect 2222 3087 2223 3091
rect 2227 3087 2228 3091
rect 2222 3086 2228 3087
rect 2374 3091 2380 3092
rect 2374 3087 2375 3091
rect 2379 3087 2380 3091
rect 2374 3086 2380 3087
rect 2526 3091 2532 3092
rect 2526 3087 2527 3091
rect 2531 3087 2532 3091
rect 2526 3086 2532 3087
rect 2686 3091 2692 3092
rect 2686 3087 2687 3091
rect 2691 3087 2692 3091
rect 2686 3086 2692 3087
rect 2854 3091 2860 3092
rect 2854 3087 2855 3091
rect 2859 3087 2860 3091
rect 2854 3086 2860 3087
rect 3038 3091 3044 3092
rect 3038 3087 3039 3091
rect 3043 3087 3044 3091
rect 3038 3086 3044 3087
rect 3230 3091 3236 3092
rect 3230 3087 3231 3091
rect 3235 3087 3236 3091
rect 3230 3086 3236 3087
rect 3430 3091 3436 3092
rect 3430 3087 3431 3091
rect 3435 3087 3436 3091
rect 3430 3086 3436 3087
rect 3638 3091 3644 3092
rect 3638 3087 3639 3091
rect 3643 3087 3644 3091
rect 3638 3086 3644 3087
rect 3838 3091 3844 3092
rect 3838 3087 3839 3091
rect 3843 3087 3844 3091
rect 3942 3088 3943 3092
rect 3947 3088 3948 3092
rect 3942 3087 3948 3088
rect 3838 3086 3844 3087
rect 2046 3075 2052 3076
rect 2046 3071 2047 3075
rect 2051 3071 2052 3075
rect 3942 3075 3948 3076
rect 2046 3070 2052 3071
rect 2078 3072 2084 3073
rect 110 3068 116 3069
rect 2006 3068 2012 3069
rect 110 3064 111 3068
rect 115 3064 116 3068
rect 110 3063 116 3064
rect 262 3067 268 3068
rect 262 3063 263 3067
rect 267 3063 268 3067
rect 262 3062 268 3063
rect 438 3067 444 3068
rect 438 3063 439 3067
rect 443 3063 444 3067
rect 438 3062 444 3063
rect 614 3067 620 3068
rect 614 3063 615 3067
rect 619 3063 620 3067
rect 614 3062 620 3063
rect 798 3067 804 3068
rect 798 3063 799 3067
rect 803 3063 804 3067
rect 798 3062 804 3063
rect 974 3067 980 3068
rect 974 3063 975 3067
rect 979 3063 980 3067
rect 974 3062 980 3063
rect 1142 3067 1148 3068
rect 1142 3063 1143 3067
rect 1147 3063 1148 3067
rect 1142 3062 1148 3063
rect 1302 3067 1308 3068
rect 1302 3063 1303 3067
rect 1307 3063 1308 3067
rect 1302 3062 1308 3063
rect 1454 3067 1460 3068
rect 1454 3063 1455 3067
rect 1459 3063 1460 3067
rect 1454 3062 1460 3063
rect 1606 3067 1612 3068
rect 1606 3063 1607 3067
rect 1611 3063 1612 3067
rect 1606 3062 1612 3063
rect 1766 3067 1772 3068
rect 1766 3063 1767 3067
rect 1771 3063 1772 3067
rect 2006 3064 2007 3068
rect 2011 3064 2012 3068
rect 2078 3068 2079 3072
rect 2083 3068 2084 3072
rect 2078 3067 2084 3068
rect 2222 3072 2228 3073
rect 2222 3068 2223 3072
rect 2227 3068 2228 3072
rect 2222 3067 2228 3068
rect 2374 3072 2380 3073
rect 2374 3068 2375 3072
rect 2379 3068 2380 3072
rect 2374 3067 2380 3068
rect 2526 3072 2532 3073
rect 2526 3068 2527 3072
rect 2531 3068 2532 3072
rect 2526 3067 2532 3068
rect 2686 3072 2692 3073
rect 2686 3068 2687 3072
rect 2691 3068 2692 3072
rect 2686 3067 2692 3068
rect 2854 3072 2860 3073
rect 2854 3068 2855 3072
rect 2859 3068 2860 3072
rect 2854 3067 2860 3068
rect 3038 3072 3044 3073
rect 3038 3068 3039 3072
rect 3043 3068 3044 3072
rect 3038 3067 3044 3068
rect 3230 3072 3236 3073
rect 3230 3068 3231 3072
rect 3235 3068 3236 3072
rect 3230 3067 3236 3068
rect 3430 3072 3436 3073
rect 3430 3068 3431 3072
rect 3435 3068 3436 3072
rect 3430 3067 3436 3068
rect 3638 3072 3644 3073
rect 3638 3068 3639 3072
rect 3643 3068 3644 3072
rect 3638 3067 3644 3068
rect 3838 3072 3844 3073
rect 3838 3068 3839 3072
rect 3843 3068 3844 3072
rect 3942 3071 3943 3075
rect 3947 3071 3948 3075
rect 3942 3070 3948 3071
rect 3838 3067 3844 3068
rect 2006 3063 2012 3064
rect 1766 3062 1772 3063
rect 110 3051 116 3052
rect 110 3047 111 3051
rect 115 3047 116 3051
rect 2006 3051 2012 3052
rect 110 3046 116 3047
rect 262 3048 268 3049
rect 262 3044 263 3048
rect 267 3044 268 3048
rect 262 3043 268 3044
rect 438 3048 444 3049
rect 438 3044 439 3048
rect 443 3044 444 3048
rect 438 3043 444 3044
rect 614 3048 620 3049
rect 614 3044 615 3048
rect 619 3044 620 3048
rect 614 3043 620 3044
rect 798 3048 804 3049
rect 798 3044 799 3048
rect 803 3044 804 3048
rect 798 3043 804 3044
rect 974 3048 980 3049
rect 974 3044 975 3048
rect 979 3044 980 3048
rect 974 3043 980 3044
rect 1142 3048 1148 3049
rect 1142 3044 1143 3048
rect 1147 3044 1148 3048
rect 1142 3043 1148 3044
rect 1302 3048 1308 3049
rect 1302 3044 1303 3048
rect 1307 3044 1308 3048
rect 1302 3043 1308 3044
rect 1454 3048 1460 3049
rect 1454 3044 1455 3048
rect 1459 3044 1460 3048
rect 1454 3043 1460 3044
rect 1606 3048 1612 3049
rect 1606 3044 1607 3048
rect 1611 3044 1612 3048
rect 1606 3043 1612 3044
rect 1766 3048 1772 3049
rect 1766 3044 1767 3048
rect 1771 3044 1772 3048
rect 2006 3047 2007 3051
rect 2011 3047 2012 3051
rect 2006 3046 2012 3047
rect 1766 3043 1772 3044
rect 2070 3004 2076 3005
rect 2046 3001 2052 3002
rect 2046 2997 2047 3001
rect 2051 2997 2052 3001
rect 2070 3000 2071 3004
rect 2075 3000 2076 3004
rect 2070 2999 2076 3000
rect 2182 3004 2188 3005
rect 2182 3000 2183 3004
rect 2187 3000 2188 3004
rect 2182 2999 2188 3000
rect 2326 3004 2332 3005
rect 2326 3000 2327 3004
rect 2331 3000 2332 3004
rect 2326 2999 2332 3000
rect 2478 3004 2484 3005
rect 2478 3000 2479 3004
rect 2483 3000 2484 3004
rect 2478 2999 2484 3000
rect 2654 3004 2660 3005
rect 2654 3000 2655 3004
rect 2659 3000 2660 3004
rect 2654 2999 2660 3000
rect 2854 3004 2860 3005
rect 2854 3000 2855 3004
rect 2859 3000 2860 3004
rect 2854 2999 2860 3000
rect 3086 3004 3092 3005
rect 3086 3000 3087 3004
rect 3091 3000 3092 3004
rect 3086 2999 3092 3000
rect 3334 3004 3340 3005
rect 3334 3000 3335 3004
rect 3339 3000 3340 3004
rect 3334 2999 3340 3000
rect 3598 3004 3604 3005
rect 3598 3000 3599 3004
rect 3603 3000 3604 3004
rect 3598 2999 3604 3000
rect 3838 3004 3844 3005
rect 3838 3000 3839 3004
rect 3843 3000 3844 3004
rect 3838 2999 3844 3000
rect 3942 3001 3948 3002
rect 2046 2996 2052 2997
rect 3942 2997 3943 3001
rect 3947 2997 3948 3001
rect 3942 2996 3948 2997
rect 2070 2985 2076 2986
rect 2046 2984 2052 2985
rect 2046 2980 2047 2984
rect 2051 2980 2052 2984
rect 2070 2981 2071 2985
rect 2075 2981 2076 2985
rect 2070 2980 2076 2981
rect 2182 2985 2188 2986
rect 2182 2981 2183 2985
rect 2187 2981 2188 2985
rect 2182 2980 2188 2981
rect 2326 2985 2332 2986
rect 2326 2981 2327 2985
rect 2331 2981 2332 2985
rect 2326 2980 2332 2981
rect 2478 2985 2484 2986
rect 2478 2981 2479 2985
rect 2483 2981 2484 2985
rect 2478 2980 2484 2981
rect 2654 2985 2660 2986
rect 2654 2981 2655 2985
rect 2659 2981 2660 2985
rect 2654 2980 2660 2981
rect 2854 2985 2860 2986
rect 2854 2981 2855 2985
rect 2859 2981 2860 2985
rect 2854 2980 2860 2981
rect 3086 2985 3092 2986
rect 3086 2981 3087 2985
rect 3091 2981 3092 2985
rect 3086 2980 3092 2981
rect 3334 2985 3340 2986
rect 3334 2981 3335 2985
rect 3339 2981 3340 2985
rect 3334 2980 3340 2981
rect 3598 2985 3604 2986
rect 3598 2981 3599 2985
rect 3603 2981 3604 2985
rect 3598 2980 3604 2981
rect 3838 2985 3844 2986
rect 3838 2981 3839 2985
rect 3843 2981 3844 2985
rect 3838 2980 3844 2981
rect 3942 2984 3948 2985
rect 3942 2980 3943 2984
rect 3947 2980 3948 2984
rect 2046 2979 2052 2980
rect 3942 2979 3948 2980
rect 342 2964 348 2965
rect 110 2961 116 2962
rect 110 2957 111 2961
rect 115 2957 116 2961
rect 342 2960 343 2964
rect 347 2960 348 2964
rect 342 2959 348 2960
rect 438 2964 444 2965
rect 438 2960 439 2964
rect 443 2960 444 2964
rect 438 2959 444 2960
rect 542 2964 548 2965
rect 542 2960 543 2964
rect 547 2960 548 2964
rect 542 2959 548 2960
rect 654 2964 660 2965
rect 654 2960 655 2964
rect 659 2960 660 2964
rect 654 2959 660 2960
rect 782 2964 788 2965
rect 782 2960 783 2964
rect 787 2960 788 2964
rect 782 2959 788 2960
rect 934 2964 940 2965
rect 934 2960 935 2964
rect 939 2960 940 2964
rect 934 2959 940 2960
rect 1102 2964 1108 2965
rect 1102 2960 1103 2964
rect 1107 2960 1108 2964
rect 1102 2959 1108 2960
rect 1294 2964 1300 2965
rect 1294 2960 1295 2964
rect 1299 2960 1300 2964
rect 1294 2959 1300 2960
rect 1494 2964 1500 2965
rect 1494 2960 1495 2964
rect 1499 2960 1500 2964
rect 1494 2959 1500 2960
rect 1710 2964 1716 2965
rect 1710 2960 1711 2964
rect 1715 2960 1716 2964
rect 1710 2959 1716 2960
rect 1902 2964 1908 2965
rect 1902 2960 1903 2964
rect 1907 2960 1908 2964
rect 1902 2959 1908 2960
rect 2006 2961 2012 2962
rect 110 2956 116 2957
rect 2006 2957 2007 2961
rect 2011 2957 2012 2961
rect 2006 2956 2012 2957
rect 342 2945 348 2946
rect 110 2944 116 2945
rect 110 2940 111 2944
rect 115 2940 116 2944
rect 342 2941 343 2945
rect 347 2941 348 2945
rect 342 2940 348 2941
rect 438 2945 444 2946
rect 438 2941 439 2945
rect 443 2941 444 2945
rect 438 2940 444 2941
rect 542 2945 548 2946
rect 542 2941 543 2945
rect 547 2941 548 2945
rect 542 2940 548 2941
rect 654 2945 660 2946
rect 654 2941 655 2945
rect 659 2941 660 2945
rect 654 2940 660 2941
rect 782 2945 788 2946
rect 782 2941 783 2945
rect 787 2941 788 2945
rect 782 2940 788 2941
rect 934 2945 940 2946
rect 934 2941 935 2945
rect 939 2941 940 2945
rect 934 2940 940 2941
rect 1102 2945 1108 2946
rect 1102 2941 1103 2945
rect 1107 2941 1108 2945
rect 1102 2940 1108 2941
rect 1294 2945 1300 2946
rect 1294 2941 1295 2945
rect 1299 2941 1300 2945
rect 1294 2940 1300 2941
rect 1494 2945 1500 2946
rect 1494 2941 1495 2945
rect 1499 2941 1500 2945
rect 1494 2940 1500 2941
rect 1710 2945 1716 2946
rect 1710 2941 1711 2945
rect 1715 2941 1716 2945
rect 1710 2940 1716 2941
rect 1902 2945 1908 2946
rect 1902 2941 1903 2945
rect 1907 2941 1908 2945
rect 1902 2940 1908 2941
rect 2006 2944 2012 2945
rect 2006 2940 2007 2944
rect 2011 2940 2012 2944
rect 110 2939 116 2940
rect 2006 2939 2012 2940
rect 2046 2928 2052 2929
rect 3942 2928 3948 2929
rect 2046 2924 2047 2928
rect 2051 2924 2052 2928
rect 2046 2923 2052 2924
rect 2070 2927 2076 2928
rect 2070 2923 2071 2927
rect 2075 2923 2076 2927
rect 2070 2922 2076 2923
rect 2262 2927 2268 2928
rect 2262 2923 2263 2927
rect 2267 2923 2268 2927
rect 2262 2922 2268 2923
rect 2486 2927 2492 2928
rect 2486 2923 2487 2927
rect 2491 2923 2492 2927
rect 2486 2922 2492 2923
rect 2734 2927 2740 2928
rect 2734 2923 2735 2927
rect 2739 2923 2740 2927
rect 2734 2922 2740 2923
rect 2998 2927 3004 2928
rect 2998 2923 2999 2927
rect 3003 2923 3004 2927
rect 2998 2922 3004 2923
rect 3278 2927 3284 2928
rect 3278 2923 3279 2927
rect 3283 2923 3284 2927
rect 3278 2922 3284 2923
rect 3566 2927 3572 2928
rect 3566 2923 3567 2927
rect 3571 2923 3572 2927
rect 3566 2922 3572 2923
rect 3838 2927 3844 2928
rect 3838 2923 3839 2927
rect 3843 2923 3844 2927
rect 3942 2924 3943 2928
rect 3947 2924 3948 2928
rect 3942 2923 3948 2924
rect 3838 2922 3844 2923
rect 2046 2911 2052 2912
rect 2046 2907 2047 2911
rect 2051 2907 2052 2911
rect 3942 2911 3948 2912
rect 2046 2906 2052 2907
rect 2070 2908 2076 2909
rect 2070 2904 2071 2908
rect 2075 2904 2076 2908
rect 2070 2903 2076 2904
rect 2262 2908 2268 2909
rect 2262 2904 2263 2908
rect 2267 2904 2268 2908
rect 2262 2903 2268 2904
rect 2486 2908 2492 2909
rect 2486 2904 2487 2908
rect 2491 2904 2492 2908
rect 2486 2903 2492 2904
rect 2734 2908 2740 2909
rect 2734 2904 2735 2908
rect 2739 2904 2740 2908
rect 2734 2903 2740 2904
rect 2998 2908 3004 2909
rect 2998 2904 2999 2908
rect 3003 2904 3004 2908
rect 2998 2903 3004 2904
rect 3278 2908 3284 2909
rect 3278 2904 3279 2908
rect 3283 2904 3284 2908
rect 3278 2903 3284 2904
rect 3566 2908 3572 2909
rect 3566 2904 3567 2908
rect 3571 2904 3572 2908
rect 3566 2903 3572 2904
rect 3838 2908 3844 2909
rect 3838 2904 3839 2908
rect 3843 2904 3844 2908
rect 3942 2907 3943 2911
rect 3947 2907 3948 2911
rect 3942 2906 3948 2907
rect 3838 2903 3844 2904
rect 110 2892 116 2893
rect 2006 2892 2012 2893
rect 110 2888 111 2892
rect 115 2888 116 2892
rect 110 2887 116 2888
rect 206 2891 212 2892
rect 206 2887 207 2891
rect 211 2887 212 2891
rect 206 2886 212 2887
rect 326 2891 332 2892
rect 326 2887 327 2891
rect 331 2887 332 2891
rect 326 2886 332 2887
rect 446 2891 452 2892
rect 446 2887 447 2891
rect 451 2887 452 2891
rect 446 2886 452 2887
rect 574 2891 580 2892
rect 574 2887 575 2891
rect 579 2887 580 2891
rect 574 2886 580 2887
rect 702 2891 708 2892
rect 702 2887 703 2891
rect 707 2887 708 2891
rect 702 2886 708 2887
rect 846 2891 852 2892
rect 846 2887 847 2891
rect 851 2887 852 2891
rect 846 2886 852 2887
rect 998 2891 1004 2892
rect 998 2887 999 2891
rect 1003 2887 1004 2891
rect 998 2886 1004 2887
rect 1166 2891 1172 2892
rect 1166 2887 1167 2891
rect 1171 2887 1172 2891
rect 1166 2886 1172 2887
rect 1350 2891 1356 2892
rect 1350 2887 1351 2891
rect 1355 2887 1356 2891
rect 1350 2886 1356 2887
rect 1534 2891 1540 2892
rect 1534 2887 1535 2891
rect 1539 2887 1540 2891
rect 1534 2886 1540 2887
rect 1726 2891 1732 2892
rect 1726 2887 1727 2891
rect 1731 2887 1732 2891
rect 1726 2886 1732 2887
rect 1902 2891 1908 2892
rect 1902 2887 1903 2891
rect 1907 2887 1908 2891
rect 2006 2888 2007 2892
rect 2011 2888 2012 2892
rect 2006 2887 2012 2888
rect 1902 2886 1908 2887
rect 110 2875 116 2876
rect 110 2871 111 2875
rect 115 2871 116 2875
rect 2006 2875 2012 2876
rect 110 2870 116 2871
rect 206 2872 212 2873
rect 206 2868 207 2872
rect 211 2868 212 2872
rect 206 2867 212 2868
rect 326 2872 332 2873
rect 326 2868 327 2872
rect 331 2868 332 2872
rect 326 2867 332 2868
rect 446 2872 452 2873
rect 446 2868 447 2872
rect 451 2868 452 2872
rect 446 2867 452 2868
rect 574 2872 580 2873
rect 574 2868 575 2872
rect 579 2868 580 2872
rect 574 2867 580 2868
rect 702 2872 708 2873
rect 702 2868 703 2872
rect 707 2868 708 2872
rect 702 2867 708 2868
rect 846 2872 852 2873
rect 846 2868 847 2872
rect 851 2868 852 2872
rect 846 2867 852 2868
rect 998 2872 1004 2873
rect 998 2868 999 2872
rect 1003 2868 1004 2872
rect 998 2867 1004 2868
rect 1166 2872 1172 2873
rect 1166 2868 1167 2872
rect 1171 2868 1172 2872
rect 1166 2867 1172 2868
rect 1350 2872 1356 2873
rect 1350 2868 1351 2872
rect 1355 2868 1356 2872
rect 1350 2867 1356 2868
rect 1534 2872 1540 2873
rect 1534 2868 1535 2872
rect 1539 2868 1540 2872
rect 1534 2867 1540 2868
rect 1726 2872 1732 2873
rect 1726 2868 1727 2872
rect 1731 2868 1732 2872
rect 1726 2867 1732 2868
rect 1902 2872 1908 2873
rect 1902 2868 1903 2872
rect 1907 2868 1908 2872
rect 2006 2871 2007 2875
rect 2011 2871 2012 2875
rect 2006 2870 2012 2871
rect 1902 2867 1908 2868
rect 2670 2840 2676 2841
rect 2046 2837 2052 2838
rect 2046 2833 2047 2837
rect 2051 2833 2052 2837
rect 2670 2836 2671 2840
rect 2675 2836 2676 2840
rect 2670 2835 2676 2836
rect 2886 2840 2892 2841
rect 2886 2836 2887 2840
rect 2891 2836 2892 2840
rect 2886 2835 2892 2836
rect 3094 2840 3100 2841
rect 3094 2836 3095 2840
rect 3099 2836 3100 2840
rect 3094 2835 3100 2836
rect 3286 2840 3292 2841
rect 3286 2836 3287 2840
rect 3291 2836 3292 2840
rect 3286 2835 3292 2836
rect 3478 2840 3484 2841
rect 3478 2836 3479 2840
rect 3483 2836 3484 2840
rect 3478 2835 3484 2836
rect 3670 2840 3676 2841
rect 3670 2836 3671 2840
rect 3675 2836 3676 2840
rect 3670 2835 3676 2836
rect 3838 2840 3844 2841
rect 3838 2836 3839 2840
rect 3843 2836 3844 2840
rect 3838 2835 3844 2836
rect 3942 2837 3948 2838
rect 2046 2832 2052 2833
rect 3942 2833 3943 2837
rect 3947 2833 3948 2837
rect 3942 2832 3948 2833
rect 2670 2821 2676 2822
rect 2046 2820 2052 2821
rect 2046 2816 2047 2820
rect 2051 2816 2052 2820
rect 2670 2817 2671 2821
rect 2675 2817 2676 2821
rect 2670 2816 2676 2817
rect 2886 2821 2892 2822
rect 2886 2817 2887 2821
rect 2891 2817 2892 2821
rect 2886 2816 2892 2817
rect 3094 2821 3100 2822
rect 3094 2817 3095 2821
rect 3099 2817 3100 2821
rect 3094 2816 3100 2817
rect 3286 2821 3292 2822
rect 3286 2817 3287 2821
rect 3291 2817 3292 2821
rect 3286 2816 3292 2817
rect 3478 2821 3484 2822
rect 3478 2817 3479 2821
rect 3483 2817 3484 2821
rect 3478 2816 3484 2817
rect 3670 2821 3676 2822
rect 3670 2817 3671 2821
rect 3675 2817 3676 2821
rect 3670 2816 3676 2817
rect 3838 2821 3844 2822
rect 3838 2817 3839 2821
rect 3843 2817 3844 2821
rect 3838 2816 3844 2817
rect 3942 2820 3948 2821
rect 3942 2816 3943 2820
rect 3947 2816 3948 2820
rect 2046 2815 2052 2816
rect 3942 2815 3948 2816
rect 134 2808 140 2809
rect 110 2805 116 2806
rect 110 2801 111 2805
rect 115 2801 116 2805
rect 134 2804 135 2808
rect 139 2804 140 2808
rect 134 2803 140 2804
rect 246 2808 252 2809
rect 246 2804 247 2808
rect 251 2804 252 2808
rect 246 2803 252 2804
rect 398 2808 404 2809
rect 398 2804 399 2808
rect 403 2804 404 2808
rect 398 2803 404 2804
rect 550 2808 556 2809
rect 550 2804 551 2808
rect 555 2804 556 2808
rect 550 2803 556 2804
rect 710 2808 716 2809
rect 710 2804 711 2808
rect 715 2804 716 2808
rect 710 2803 716 2804
rect 878 2808 884 2809
rect 878 2804 879 2808
rect 883 2804 884 2808
rect 878 2803 884 2804
rect 1046 2808 1052 2809
rect 1046 2804 1047 2808
rect 1051 2804 1052 2808
rect 1046 2803 1052 2804
rect 1222 2808 1228 2809
rect 1222 2804 1223 2808
rect 1227 2804 1228 2808
rect 1222 2803 1228 2804
rect 1398 2808 1404 2809
rect 1398 2804 1399 2808
rect 1403 2804 1404 2808
rect 1398 2803 1404 2804
rect 1574 2808 1580 2809
rect 1574 2804 1575 2808
rect 1579 2804 1580 2808
rect 1574 2803 1580 2804
rect 1750 2808 1756 2809
rect 1750 2804 1751 2808
rect 1755 2804 1756 2808
rect 1750 2803 1756 2804
rect 1902 2808 1908 2809
rect 1902 2804 1903 2808
rect 1907 2804 1908 2808
rect 1902 2803 1908 2804
rect 2006 2805 2012 2806
rect 110 2800 116 2801
rect 2006 2801 2007 2805
rect 2011 2801 2012 2805
rect 2006 2800 2012 2801
rect 134 2789 140 2790
rect 110 2788 116 2789
rect 110 2784 111 2788
rect 115 2784 116 2788
rect 134 2785 135 2789
rect 139 2785 140 2789
rect 134 2784 140 2785
rect 246 2789 252 2790
rect 246 2785 247 2789
rect 251 2785 252 2789
rect 246 2784 252 2785
rect 398 2789 404 2790
rect 398 2785 399 2789
rect 403 2785 404 2789
rect 398 2784 404 2785
rect 550 2789 556 2790
rect 550 2785 551 2789
rect 555 2785 556 2789
rect 550 2784 556 2785
rect 710 2789 716 2790
rect 710 2785 711 2789
rect 715 2785 716 2789
rect 710 2784 716 2785
rect 878 2789 884 2790
rect 878 2785 879 2789
rect 883 2785 884 2789
rect 878 2784 884 2785
rect 1046 2789 1052 2790
rect 1046 2785 1047 2789
rect 1051 2785 1052 2789
rect 1046 2784 1052 2785
rect 1222 2789 1228 2790
rect 1222 2785 1223 2789
rect 1227 2785 1228 2789
rect 1222 2784 1228 2785
rect 1398 2789 1404 2790
rect 1398 2785 1399 2789
rect 1403 2785 1404 2789
rect 1398 2784 1404 2785
rect 1574 2789 1580 2790
rect 1574 2785 1575 2789
rect 1579 2785 1580 2789
rect 1574 2784 1580 2785
rect 1750 2789 1756 2790
rect 1750 2785 1751 2789
rect 1755 2785 1756 2789
rect 1750 2784 1756 2785
rect 1902 2789 1908 2790
rect 1902 2785 1903 2789
rect 1907 2785 1908 2789
rect 1902 2784 1908 2785
rect 2006 2788 2012 2789
rect 2006 2784 2007 2788
rect 2011 2784 2012 2788
rect 110 2783 116 2784
rect 2006 2783 2012 2784
rect 2046 2768 2052 2769
rect 3942 2768 3948 2769
rect 2046 2764 2047 2768
rect 2051 2764 2052 2768
rect 2046 2763 2052 2764
rect 2070 2767 2076 2768
rect 2070 2763 2071 2767
rect 2075 2763 2076 2767
rect 2070 2762 2076 2763
rect 2198 2767 2204 2768
rect 2198 2763 2199 2767
rect 2203 2763 2204 2767
rect 2198 2762 2204 2763
rect 2342 2767 2348 2768
rect 2342 2763 2343 2767
rect 2347 2763 2348 2767
rect 2342 2762 2348 2763
rect 2478 2767 2484 2768
rect 2478 2763 2479 2767
rect 2483 2763 2484 2767
rect 2478 2762 2484 2763
rect 2606 2767 2612 2768
rect 2606 2763 2607 2767
rect 2611 2763 2612 2767
rect 2606 2762 2612 2763
rect 2726 2767 2732 2768
rect 2726 2763 2727 2767
rect 2731 2763 2732 2767
rect 2726 2762 2732 2763
rect 2838 2767 2844 2768
rect 2838 2763 2839 2767
rect 2843 2763 2844 2767
rect 2838 2762 2844 2763
rect 2942 2767 2948 2768
rect 2942 2763 2943 2767
rect 2947 2763 2948 2767
rect 2942 2762 2948 2763
rect 3046 2767 3052 2768
rect 3046 2763 3047 2767
rect 3051 2763 3052 2767
rect 3046 2762 3052 2763
rect 3142 2767 3148 2768
rect 3142 2763 3143 2767
rect 3147 2763 3148 2767
rect 3142 2762 3148 2763
rect 3238 2767 3244 2768
rect 3238 2763 3239 2767
rect 3243 2763 3244 2767
rect 3238 2762 3244 2763
rect 3342 2767 3348 2768
rect 3342 2763 3343 2767
rect 3347 2763 3348 2767
rect 3342 2762 3348 2763
rect 3446 2767 3452 2768
rect 3446 2763 3447 2767
rect 3451 2763 3452 2767
rect 3446 2762 3452 2763
rect 3550 2767 3556 2768
rect 3550 2763 3551 2767
rect 3555 2763 3556 2767
rect 3550 2762 3556 2763
rect 3646 2767 3652 2768
rect 3646 2763 3647 2767
rect 3651 2763 3652 2767
rect 3646 2762 3652 2763
rect 3742 2767 3748 2768
rect 3742 2763 3743 2767
rect 3747 2763 3748 2767
rect 3742 2762 3748 2763
rect 3838 2767 3844 2768
rect 3838 2763 3839 2767
rect 3843 2763 3844 2767
rect 3942 2764 3943 2768
rect 3947 2764 3948 2768
rect 3942 2763 3948 2764
rect 3838 2762 3844 2763
rect 2046 2751 2052 2752
rect 2046 2747 2047 2751
rect 2051 2747 2052 2751
rect 3942 2751 3948 2752
rect 2046 2746 2052 2747
rect 2070 2748 2076 2749
rect 2070 2744 2071 2748
rect 2075 2744 2076 2748
rect 2070 2743 2076 2744
rect 2198 2748 2204 2749
rect 2198 2744 2199 2748
rect 2203 2744 2204 2748
rect 2198 2743 2204 2744
rect 2342 2748 2348 2749
rect 2342 2744 2343 2748
rect 2347 2744 2348 2748
rect 2342 2743 2348 2744
rect 2478 2748 2484 2749
rect 2478 2744 2479 2748
rect 2483 2744 2484 2748
rect 2478 2743 2484 2744
rect 2606 2748 2612 2749
rect 2606 2744 2607 2748
rect 2611 2744 2612 2748
rect 2606 2743 2612 2744
rect 2726 2748 2732 2749
rect 2726 2744 2727 2748
rect 2731 2744 2732 2748
rect 2726 2743 2732 2744
rect 2838 2748 2844 2749
rect 2838 2744 2839 2748
rect 2843 2744 2844 2748
rect 2838 2743 2844 2744
rect 2942 2748 2948 2749
rect 2942 2744 2943 2748
rect 2947 2744 2948 2748
rect 2942 2743 2948 2744
rect 3046 2748 3052 2749
rect 3046 2744 3047 2748
rect 3051 2744 3052 2748
rect 3046 2743 3052 2744
rect 3142 2748 3148 2749
rect 3142 2744 3143 2748
rect 3147 2744 3148 2748
rect 3142 2743 3148 2744
rect 3238 2748 3244 2749
rect 3238 2744 3239 2748
rect 3243 2744 3244 2748
rect 3238 2743 3244 2744
rect 3342 2748 3348 2749
rect 3342 2744 3343 2748
rect 3347 2744 3348 2748
rect 3342 2743 3348 2744
rect 3446 2748 3452 2749
rect 3446 2744 3447 2748
rect 3451 2744 3452 2748
rect 3446 2743 3452 2744
rect 3550 2748 3556 2749
rect 3550 2744 3551 2748
rect 3555 2744 3556 2748
rect 3550 2743 3556 2744
rect 3646 2748 3652 2749
rect 3646 2744 3647 2748
rect 3651 2744 3652 2748
rect 3646 2743 3652 2744
rect 3742 2748 3748 2749
rect 3742 2744 3743 2748
rect 3747 2744 3748 2748
rect 3742 2743 3748 2744
rect 3838 2748 3844 2749
rect 3838 2744 3839 2748
rect 3843 2744 3844 2748
rect 3942 2747 3943 2751
rect 3947 2747 3948 2751
rect 3942 2746 3948 2747
rect 3838 2743 3844 2744
rect 110 2728 116 2729
rect 2006 2728 2012 2729
rect 110 2724 111 2728
rect 115 2724 116 2728
rect 110 2723 116 2724
rect 134 2727 140 2728
rect 134 2723 135 2727
rect 139 2723 140 2727
rect 134 2722 140 2723
rect 254 2727 260 2728
rect 254 2723 255 2727
rect 259 2723 260 2727
rect 254 2722 260 2723
rect 406 2727 412 2728
rect 406 2723 407 2727
rect 411 2723 412 2727
rect 406 2722 412 2723
rect 574 2727 580 2728
rect 574 2723 575 2727
rect 579 2723 580 2727
rect 574 2722 580 2723
rect 742 2727 748 2728
rect 742 2723 743 2727
rect 747 2723 748 2727
rect 742 2722 748 2723
rect 918 2727 924 2728
rect 918 2723 919 2727
rect 923 2723 924 2727
rect 918 2722 924 2723
rect 1086 2727 1092 2728
rect 1086 2723 1087 2727
rect 1091 2723 1092 2727
rect 1086 2722 1092 2723
rect 1254 2727 1260 2728
rect 1254 2723 1255 2727
rect 1259 2723 1260 2727
rect 1254 2722 1260 2723
rect 1422 2727 1428 2728
rect 1422 2723 1423 2727
rect 1427 2723 1428 2727
rect 1422 2722 1428 2723
rect 1598 2727 1604 2728
rect 1598 2723 1599 2727
rect 1603 2723 1604 2727
rect 2006 2724 2007 2728
rect 2011 2724 2012 2728
rect 2006 2723 2012 2724
rect 1598 2722 1604 2723
rect 110 2711 116 2712
rect 110 2707 111 2711
rect 115 2707 116 2711
rect 2006 2711 2012 2712
rect 110 2706 116 2707
rect 134 2708 140 2709
rect 134 2704 135 2708
rect 139 2704 140 2708
rect 134 2703 140 2704
rect 254 2708 260 2709
rect 254 2704 255 2708
rect 259 2704 260 2708
rect 254 2703 260 2704
rect 406 2708 412 2709
rect 406 2704 407 2708
rect 411 2704 412 2708
rect 406 2703 412 2704
rect 574 2708 580 2709
rect 574 2704 575 2708
rect 579 2704 580 2708
rect 574 2703 580 2704
rect 742 2708 748 2709
rect 742 2704 743 2708
rect 747 2704 748 2708
rect 742 2703 748 2704
rect 918 2708 924 2709
rect 918 2704 919 2708
rect 923 2704 924 2708
rect 918 2703 924 2704
rect 1086 2708 1092 2709
rect 1086 2704 1087 2708
rect 1091 2704 1092 2708
rect 1086 2703 1092 2704
rect 1254 2708 1260 2709
rect 1254 2704 1255 2708
rect 1259 2704 1260 2708
rect 1254 2703 1260 2704
rect 1422 2708 1428 2709
rect 1422 2704 1423 2708
rect 1427 2704 1428 2708
rect 1422 2703 1428 2704
rect 1598 2708 1604 2709
rect 1598 2704 1599 2708
rect 1603 2704 1604 2708
rect 2006 2707 2007 2711
rect 2011 2707 2012 2711
rect 2006 2706 2012 2707
rect 1598 2703 1604 2704
rect 2094 2668 2100 2669
rect 2046 2665 2052 2666
rect 2046 2661 2047 2665
rect 2051 2661 2052 2665
rect 2094 2664 2095 2668
rect 2099 2664 2100 2668
rect 2094 2663 2100 2664
rect 2262 2668 2268 2669
rect 2262 2664 2263 2668
rect 2267 2664 2268 2668
rect 2262 2663 2268 2664
rect 2438 2668 2444 2669
rect 2438 2664 2439 2668
rect 2443 2664 2444 2668
rect 2438 2663 2444 2664
rect 2614 2668 2620 2669
rect 2614 2664 2615 2668
rect 2619 2664 2620 2668
rect 2614 2663 2620 2664
rect 2782 2668 2788 2669
rect 2782 2664 2783 2668
rect 2787 2664 2788 2668
rect 2782 2663 2788 2664
rect 2942 2668 2948 2669
rect 2942 2664 2943 2668
rect 2947 2664 2948 2668
rect 2942 2663 2948 2664
rect 3094 2668 3100 2669
rect 3094 2664 3095 2668
rect 3099 2664 3100 2668
rect 3094 2663 3100 2664
rect 3238 2668 3244 2669
rect 3238 2664 3239 2668
rect 3243 2664 3244 2668
rect 3238 2663 3244 2664
rect 3382 2668 3388 2669
rect 3382 2664 3383 2668
rect 3387 2664 3388 2668
rect 3382 2663 3388 2664
rect 3534 2668 3540 2669
rect 3534 2664 3535 2668
rect 3539 2664 3540 2668
rect 3534 2663 3540 2664
rect 3942 2665 3948 2666
rect 2046 2660 2052 2661
rect 3942 2661 3943 2665
rect 3947 2661 3948 2665
rect 3942 2660 3948 2661
rect 2094 2649 2100 2650
rect 166 2648 172 2649
rect 110 2645 116 2646
rect 110 2641 111 2645
rect 115 2641 116 2645
rect 166 2644 167 2648
rect 171 2644 172 2648
rect 166 2643 172 2644
rect 358 2648 364 2649
rect 358 2644 359 2648
rect 363 2644 364 2648
rect 358 2643 364 2644
rect 558 2648 564 2649
rect 558 2644 559 2648
rect 563 2644 564 2648
rect 558 2643 564 2644
rect 758 2648 764 2649
rect 758 2644 759 2648
rect 763 2644 764 2648
rect 758 2643 764 2644
rect 950 2648 956 2649
rect 950 2644 951 2648
rect 955 2644 956 2648
rect 950 2643 956 2644
rect 1142 2648 1148 2649
rect 1142 2644 1143 2648
rect 1147 2644 1148 2648
rect 1142 2643 1148 2644
rect 1326 2648 1332 2649
rect 1326 2644 1327 2648
rect 1331 2644 1332 2648
rect 1326 2643 1332 2644
rect 1510 2648 1516 2649
rect 1510 2644 1511 2648
rect 1515 2644 1516 2648
rect 1510 2643 1516 2644
rect 1702 2648 1708 2649
rect 1702 2644 1703 2648
rect 1707 2644 1708 2648
rect 2046 2648 2052 2649
rect 1702 2643 1708 2644
rect 2006 2645 2012 2646
rect 110 2640 116 2641
rect 2006 2641 2007 2645
rect 2011 2641 2012 2645
rect 2046 2644 2047 2648
rect 2051 2644 2052 2648
rect 2094 2645 2095 2649
rect 2099 2645 2100 2649
rect 2094 2644 2100 2645
rect 2262 2649 2268 2650
rect 2262 2645 2263 2649
rect 2267 2645 2268 2649
rect 2262 2644 2268 2645
rect 2438 2649 2444 2650
rect 2438 2645 2439 2649
rect 2443 2645 2444 2649
rect 2438 2644 2444 2645
rect 2614 2649 2620 2650
rect 2614 2645 2615 2649
rect 2619 2645 2620 2649
rect 2614 2644 2620 2645
rect 2782 2649 2788 2650
rect 2782 2645 2783 2649
rect 2787 2645 2788 2649
rect 2782 2644 2788 2645
rect 2942 2649 2948 2650
rect 2942 2645 2943 2649
rect 2947 2645 2948 2649
rect 2942 2644 2948 2645
rect 3094 2649 3100 2650
rect 3094 2645 3095 2649
rect 3099 2645 3100 2649
rect 3094 2644 3100 2645
rect 3238 2649 3244 2650
rect 3238 2645 3239 2649
rect 3243 2645 3244 2649
rect 3238 2644 3244 2645
rect 3382 2649 3388 2650
rect 3382 2645 3383 2649
rect 3387 2645 3388 2649
rect 3382 2644 3388 2645
rect 3534 2649 3540 2650
rect 3534 2645 3535 2649
rect 3539 2645 3540 2649
rect 3534 2644 3540 2645
rect 3942 2648 3948 2649
rect 3942 2644 3943 2648
rect 3947 2644 3948 2648
rect 2046 2643 2052 2644
rect 3942 2643 3948 2644
rect 2006 2640 2012 2641
rect 166 2629 172 2630
rect 110 2628 116 2629
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 166 2625 167 2629
rect 171 2625 172 2629
rect 166 2624 172 2625
rect 358 2629 364 2630
rect 358 2625 359 2629
rect 363 2625 364 2629
rect 358 2624 364 2625
rect 558 2629 564 2630
rect 558 2625 559 2629
rect 563 2625 564 2629
rect 558 2624 564 2625
rect 758 2629 764 2630
rect 758 2625 759 2629
rect 763 2625 764 2629
rect 758 2624 764 2625
rect 950 2629 956 2630
rect 950 2625 951 2629
rect 955 2625 956 2629
rect 950 2624 956 2625
rect 1142 2629 1148 2630
rect 1142 2625 1143 2629
rect 1147 2625 1148 2629
rect 1142 2624 1148 2625
rect 1326 2629 1332 2630
rect 1326 2625 1327 2629
rect 1331 2625 1332 2629
rect 1326 2624 1332 2625
rect 1510 2629 1516 2630
rect 1510 2625 1511 2629
rect 1515 2625 1516 2629
rect 1510 2624 1516 2625
rect 1702 2629 1708 2630
rect 1702 2625 1703 2629
rect 1707 2625 1708 2629
rect 1702 2624 1708 2625
rect 2006 2628 2012 2629
rect 2006 2624 2007 2628
rect 2011 2624 2012 2628
rect 110 2623 116 2624
rect 2006 2623 2012 2624
rect 2046 2588 2052 2589
rect 3942 2588 3948 2589
rect 2046 2584 2047 2588
rect 2051 2584 2052 2588
rect 2046 2583 2052 2584
rect 2214 2587 2220 2588
rect 2214 2583 2215 2587
rect 2219 2583 2220 2587
rect 2214 2582 2220 2583
rect 2366 2587 2372 2588
rect 2366 2583 2367 2587
rect 2371 2583 2372 2587
rect 2366 2582 2372 2583
rect 2518 2587 2524 2588
rect 2518 2583 2519 2587
rect 2523 2583 2524 2587
rect 2518 2582 2524 2583
rect 2670 2587 2676 2588
rect 2670 2583 2671 2587
rect 2675 2583 2676 2587
rect 2670 2582 2676 2583
rect 2814 2587 2820 2588
rect 2814 2583 2815 2587
rect 2819 2583 2820 2587
rect 2814 2582 2820 2583
rect 2950 2587 2956 2588
rect 2950 2583 2951 2587
rect 2955 2583 2956 2587
rect 2950 2582 2956 2583
rect 3086 2587 3092 2588
rect 3086 2583 3087 2587
rect 3091 2583 3092 2587
rect 3086 2582 3092 2583
rect 3222 2587 3228 2588
rect 3222 2583 3223 2587
rect 3227 2583 3228 2587
rect 3222 2582 3228 2583
rect 3366 2587 3372 2588
rect 3366 2583 3367 2587
rect 3371 2583 3372 2587
rect 3942 2584 3943 2588
rect 3947 2584 3948 2588
rect 3942 2583 3948 2584
rect 3366 2582 3372 2583
rect 2046 2571 2052 2572
rect 2046 2567 2047 2571
rect 2051 2567 2052 2571
rect 3942 2571 3948 2572
rect 2046 2566 2052 2567
rect 2214 2568 2220 2569
rect 2214 2564 2215 2568
rect 2219 2564 2220 2568
rect 2214 2563 2220 2564
rect 2366 2568 2372 2569
rect 2366 2564 2367 2568
rect 2371 2564 2372 2568
rect 2366 2563 2372 2564
rect 2518 2568 2524 2569
rect 2518 2564 2519 2568
rect 2523 2564 2524 2568
rect 2518 2563 2524 2564
rect 2670 2568 2676 2569
rect 2670 2564 2671 2568
rect 2675 2564 2676 2568
rect 2670 2563 2676 2564
rect 2814 2568 2820 2569
rect 2814 2564 2815 2568
rect 2819 2564 2820 2568
rect 2814 2563 2820 2564
rect 2950 2568 2956 2569
rect 2950 2564 2951 2568
rect 2955 2564 2956 2568
rect 2950 2563 2956 2564
rect 3086 2568 3092 2569
rect 3086 2564 3087 2568
rect 3091 2564 3092 2568
rect 3086 2563 3092 2564
rect 3222 2568 3228 2569
rect 3222 2564 3223 2568
rect 3227 2564 3228 2568
rect 3222 2563 3228 2564
rect 3366 2568 3372 2569
rect 3366 2564 3367 2568
rect 3371 2564 3372 2568
rect 3942 2567 3943 2571
rect 3947 2567 3948 2571
rect 3942 2566 3948 2567
rect 3366 2563 3372 2564
rect 110 2560 116 2561
rect 2006 2560 2012 2561
rect 110 2556 111 2560
rect 115 2556 116 2560
rect 110 2555 116 2556
rect 574 2559 580 2560
rect 574 2555 575 2559
rect 579 2555 580 2559
rect 574 2554 580 2555
rect 686 2559 692 2560
rect 686 2555 687 2559
rect 691 2555 692 2559
rect 686 2554 692 2555
rect 806 2559 812 2560
rect 806 2555 807 2559
rect 811 2555 812 2559
rect 806 2554 812 2555
rect 934 2559 940 2560
rect 934 2555 935 2559
rect 939 2555 940 2559
rect 934 2554 940 2555
rect 1070 2559 1076 2560
rect 1070 2555 1071 2559
rect 1075 2555 1076 2559
rect 1070 2554 1076 2555
rect 1206 2559 1212 2560
rect 1206 2555 1207 2559
rect 1211 2555 1212 2559
rect 1206 2554 1212 2555
rect 1350 2559 1356 2560
rect 1350 2555 1351 2559
rect 1355 2555 1356 2559
rect 1350 2554 1356 2555
rect 1494 2559 1500 2560
rect 1494 2555 1495 2559
rect 1499 2555 1500 2559
rect 1494 2554 1500 2555
rect 1646 2559 1652 2560
rect 1646 2555 1647 2559
rect 1651 2555 1652 2559
rect 1646 2554 1652 2555
rect 1798 2559 1804 2560
rect 1798 2555 1799 2559
rect 1803 2555 1804 2559
rect 2006 2556 2007 2560
rect 2011 2556 2012 2560
rect 2006 2555 2012 2556
rect 1798 2554 1804 2555
rect 110 2543 116 2544
rect 110 2539 111 2543
rect 115 2539 116 2543
rect 2006 2543 2012 2544
rect 110 2538 116 2539
rect 574 2540 580 2541
rect 574 2536 575 2540
rect 579 2536 580 2540
rect 574 2535 580 2536
rect 686 2540 692 2541
rect 686 2536 687 2540
rect 691 2536 692 2540
rect 686 2535 692 2536
rect 806 2540 812 2541
rect 806 2536 807 2540
rect 811 2536 812 2540
rect 806 2535 812 2536
rect 934 2540 940 2541
rect 934 2536 935 2540
rect 939 2536 940 2540
rect 934 2535 940 2536
rect 1070 2540 1076 2541
rect 1070 2536 1071 2540
rect 1075 2536 1076 2540
rect 1070 2535 1076 2536
rect 1206 2540 1212 2541
rect 1206 2536 1207 2540
rect 1211 2536 1212 2540
rect 1206 2535 1212 2536
rect 1350 2540 1356 2541
rect 1350 2536 1351 2540
rect 1355 2536 1356 2540
rect 1350 2535 1356 2536
rect 1494 2540 1500 2541
rect 1494 2536 1495 2540
rect 1499 2536 1500 2540
rect 1494 2535 1500 2536
rect 1646 2540 1652 2541
rect 1646 2536 1647 2540
rect 1651 2536 1652 2540
rect 1646 2535 1652 2536
rect 1798 2540 1804 2541
rect 1798 2536 1799 2540
rect 1803 2536 1804 2540
rect 2006 2539 2007 2543
rect 2011 2539 2012 2543
rect 2006 2538 2012 2539
rect 1798 2535 1804 2536
rect 2094 2504 2100 2505
rect 2046 2501 2052 2502
rect 2046 2497 2047 2501
rect 2051 2497 2052 2501
rect 2094 2500 2095 2504
rect 2099 2500 2100 2504
rect 2094 2499 2100 2500
rect 2214 2504 2220 2505
rect 2214 2500 2215 2504
rect 2219 2500 2220 2504
rect 2214 2499 2220 2500
rect 2342 2504 2348 2505
rect 2342 2500 2343 2504
rect 2347 2500 2348 2504
rect 2342 2499 2348 2500
rect 2470 2504 2476 2505
rect 2470 2500 2471 2504
rect 2475 2500 2476 2504
rect 2470 2499 2476 2500
rect 2598 2504 2604 2505
rect 2598 2500 2599 2504
rect 2603 2500 2604 2504
rect 2598 2499 2604 2500
rect 2718 2504 2724 2505
rect 2718 2500 2719 2504
rect 2723 2500 2724 2504
rect 2718 2499 2724 2500
rect 2838 2504 2844 2505
rect 2838 2500 2839 2504
rect 2843 2500 2844 2504
rect 2838 2499 2844 2500
rect 2966 2504 2972 2505
rect 2966 2500 2967 2504
rect 2971 2500 2972 2504
rect 2966 2499 2972 2500
rect 3094 2504 3100 2505
rect 3094 2500 3095 2504
rect 3099 2500 3100 2504
rect 3094 2499 3100 2500
rect 3222 2504 3228 2505
rect 3222 2500 3223 2504
rect 3227 2500 3228 2504
rect 3222 2499 3228 2500
rect 3942 2501 3948 2502
rect 2046 2496 2052 2497
rect 3942 2497 3943 2501
rect 3947 2497 3948 2501
rect 3942 2496 3948 2497
rect 2094 2485 2100 2486
rect 2046 2484 2052 2485
rect 2046 2480 2047 2484
rect 2051 2480 2052 2484
rect 2094 2481 2095 2485
rect 2099 2481 2100 2485
rect 2094 2480 2100 2481
rect 2214 2485 2220 2486
rect 2214 2481 2215 2485
rect 2219 2481 2220 2485
rect 2214 2480 2220 2481
rect 2342 2485 2348 2486
rect 2342 2481 2343 2485
rect 2347 2481 2348 2485
rect 2342 2480 2348 2481
rect 2470 2485 2476 2486
rect 2470 2481 2471 2485
rect 2475 2481 2476 2485
rect 2470 2480 2476 2481
rect 2598 2485 2604 2486
rect 2598 2481 2599 2485
rect 2603 2481 2604 2485
rect 2598 2480 2604 2481
rect 2718 2485 2724 2486
rect 2718 2481 2719 2485
rect 2723 2481 2724 2485
rect 2718 2480 2724 2481
rect 2838 2485 2844 2486
rect 2838 2481 2839 2485
rect 2843 2481 2844 2485
rect 2838 2480 2844 2481
rect 2966 2485 2972 2486
rect 2966 2481 2967 2485
rect 2971 2481 2972 2485
rect 2966 2480 2972 2481
rect 3094 2485 3100 2486
rect 3094 2481 3095 2485
rect 3099 2481 3100 2485
rect 3094 2480 3100 2481
rect 3222 2485 3228 2486
rect 3222 2481 3223 2485
rect 3227 2481 3228 2485
rect 3222 2480 3228 2481
rect 3942 2484 3948 2485
rect 3942 2480 3943 2484
rect 3947 2480 3948 2484
rect 2046 2479 2052 2480
rect 3942 2479 3948 2480
rect 502 2476 508 2477
rect 110 2473 116 2474
rect 110 2469 111 2473
rect 115 2469 116 2473
rect 502 2472 503 2476
rect 507 2472 508 2476
rect 502 2471 508 2472
rect 606 2476 612 2477
rect 606 2472 607 2476
rect 611 2472 612 2476
rect 606 2471 612 2472
rect 718 2476 724 2477
rect 718 2472 719 2476
rect 723 2472 724 2476
rect 718 2471 724 2472
rect 846 2476 852 2477
rect 846 2472 847 2476
rect 851 2472 852 2476
rect 846 2471 852 2472
rect 982 2476 988 2477
rect 982 2472 983 2476
rect 987 2472 988 2476
rect 982 2471 988 2472
rect 1126 2476 1132 2477
rect 1126 2472 1127 2476
rect 1131 2472 1132 2476
rect 1126 2471 1132 2472
rect 1278 2476 1284 2477
rect 1278 2472 1279 2476
rect 1283 2472 1284 2476
rect 1278 2471 1284 2472
rect 1430 2476 1436 2477
rect 1430 2472 1431 2476
rect 1435 2472 1436 2476
rect 1430 2471 1436 2472
rect 1582 2476 1588 2477
rect 1582 2472 1583 2476
rect 1587 2472 1588 2476
rect 1582 2471 1588 2472
rect 1742 2476 1748 2477
rect 1742 2472 1743 2476
rect 1747 2472 1748 2476
rect 1742 2471 1748 2472
rect 1902 2476 1908 2477
rect 1902 2472 1903 2476
rect 1907 2472 1908 2476
rect 1902 2471 1908 2472
rect 2006 2473 2012 2474
rect 110 2468 116 2469
rect 2006 2469 2007 2473
rect 2011 2469 2012 2473
rect 2006 2468 2012 2469
rect 502 2457 508 2458
rect 110 2456 116 2457
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 502 2453 503 2457
rect 507 2453 508 2457
rect 502 2452 508 2453
rect 606 2457 612 2458
rect 606 2453 607 2457
rect 611 2453 612 2457
rect 606 2452 612 2453
rect 718 2457 724 2458
rect 718 2453 719 2457
rect 723 2453 724 2457
rect 718 2452 724 2453
rect 846 2457 852 2458
rect 846 2453 847 2457
rect 851 2453 852 2457
rect 846 2452 852 2453
rect 982 2457 988 2458
rect 982 2453 983 2457
rect 987 2453 988 2457
rect 982 2452 988 2453
rect 1126 2457 1132 2458
rect 1126 2453 1127 2457
rect 1131 2453 1132 2457
rect 1126 2452 1132 2453
rect 1278 2457 1284 2458
rect 1278 2453 1279 2457
rect 1283 2453 1284 2457
rect 1278 2452 1284 2453
rect 1430 2457 1436 2458
rect 1430 2453 1431 2457
rect 1435 2453 1436 2457
rect 1430 2452 1436 2453
rect 1582 2457 1588 2458
rect 1582 2453 1583 2457
rect 1587 2453 1588 2457
rect 1582 2452 1588 2453
rect 1742 2457 1748 2458
rect 1742 2453 1743 2457
rect 1747 2453 1748 2457
rect 1742 2452 1748 2453
rect 1902 2457 1908 2458
rect 1902 2453 1903 2457
rect 1907 2453 1908 2457
rect 1902 2452 1908 2453
rect 2006 2456 2012 2457
rect 2006 2452 2007 2456
rect 2011 2452 2012 2456
rect 110 2451 116 2452
rect 2006 2451 2012 2452
rect 2046 2420 2052 2421
rect 3942 2420 3948 2421
rect 2046 2416 2047 2420
rect 2051 2416 2052 2420
rect 2046 2415 2052 2416
rect 2070 2419 2076 2420
rect 2070 2415 2071 2419
rect 2075 2415 2076 2419
rect 2070 2414 2076 2415
rect 2190 2419 2196 2420
rect 2190 2415 2191 2419
rect 2195 2415 2196 2419
rect 2190 2414 2196 2415
rect 2318 2419 2324 2420
rect 2318 2415 2319 2419
rect 2323 2415 2324 2419
rect 2318 2414 2324 2415
rect 2438 2419 2444 2420
rect 2438 2415 2439 2419
rect 2443 2415 2444 2419
rect 2438 2414 2444 2415
rect 2558 2419 2564 2420
rect 2558 2415 2559 2419
rect 2563 2415 2564 2419
rect 2558 2414 2564 2415
rect 2678 2419 2684 2420
rect 2678 2415 2679 2419
rect 2683 2415 2684 2419
rect 2678 2414 2684 2415
rect 2790 2419 2796 2420
rect 2790 2415 2791 2419
rect 2795 2415 2796 2419
rect 2790 2414 2796 2415
rect 2910 2419 2916 2420
rect 2910 2415 2911 2419
rect 2915 2415 2916 2419
rect 2910 2414 2916 2415
rect 3030 2419 3036 2420
rect 3030 2415 3031 2419
rect 3035 2415 3036 2419
rect 3030 2414 3036 2415
rect 3150 2419 3156 2420
rect 3150 2415 3151 2419
rect 3155 2415 3156 2419
rect 3942 2416 3943 2420
rect 3947 2416 3948 2420
rect 3942 2415 3948 2416
rect 3150 2414 3156 2415
rect 2046 2403 2052 2404
rect 2046 2399 2047 2403
rect 2051 2399 2052 2403
rect 3942 2403 3948 2404
rect 2046 2398 2052 2399
rect 2070 2400 2076 2401
rect 2070 2396 2071 2400
rect 2075 2396 2076 2400
rect 2070 2395 2076 2396
rect 2190 2400 2196 2401
rect 2190 2396 2191 2400
rect 2195 2396 2196 2400
rect 2190 2395 2196 2396
rect 2318 2400 2324 2401
rect 2318 2396 2319 2400
rect 2323 2396 2324 2400
rect 2318 2395 2324 2396
rect 2438 2400 2444 2401
rect 2438 2396 2439 2400
rect 2443 2396 2444 2400
rect 2438 2395 2444 2396
rect 2558 2400 2564 2401
rect 2558 2396 2559 2400
rect 2563 2396 2564 2400
rect 2558 2395 2564 2396
rect 2678 2400 2684 2401
rect 2678 2396 2679 2400
rect 2683 2396 2684 2400
rect 2678 2395 2684 2396
rect 2790 2400 2796 2401
rect 2790 2396 2791 2400
rect 2795 2396 2796 2400
rect 2790 2395 2796 2396
rect 2910 2400 2916 2401
rect 2910 2396 2911 2400
rect 2915 2396 2916 2400
rect 2910 2395 2916 2396
rect 3030 2400 3036 2401
rect 3030 2396 3031 2400
rect 3035 2396 3036 2400
rect 3030 2395 3036 2396
rect 3150 2400 3156 2401
rect 3150 2396 3151 2400
rect 3155 2396 3156 2400
rect 3942 2399 3943 2403
rect 3947 2399 3948 2403
rect 3942 2398 3948 2399
rect 3150 2395 3156 2396
rect 110 2388 116 2389
rect 2006 2388 2012 2389
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 110 2383 116 2384
rect 534 2387 540 2388
rect 534 2383 535 2387
rect 539 2383 540 2387
rect 534 2382 540 2383
rect 670 2387 676 2388
rect 670 2383 671 2387
rect 675 2383 676 2387
rect 670 2382 676 2383
rect 814 2387 820 2388
rect 814 2383 815 2387
rect 819 2383 820 2387
rect 814 2382 820 2383
rect 958 2387 964 2388
rect 958 2383 959 2387
rect 963 2383 964 2387
rect 958 2382 964 2383
rect 1102 2387 1108 2388
rect 1102 2383 1103 2387
rect 1107 2383 1108 2387
rect 1102 2382 1108 2383
rect 1246 2387 1252 2388
rect 1246 2383 1247 2387
rect 1251 2383 1252 2387
rect 1246 2382 1252 2383
rect 1390 2387 1396 2388
rect 1390 2383 1391 2387
rect 1395 2383 1396 2387
rect 1390 2382 1396 2383
rect 1526 2387 1532 2388
rect 1526 2383 1527 2387
rect 1531 2383 1532 2387
rect 1526 2382 1532 2383
rect 1654 2387 1660 2388
rect 1654 2383 1655 2387
rect 1659 2383 1660 2387
rect 1654 2382 1660 2383
rect 1790 2387 1796 2388
rect 1790 2383 1791 2387
rect 1795 2383 1796 2387
rect 1790 2382 1796 2383
rect 1902 2387 1908 2388
rect 1902 2383 1903 2387
rect 1907 2383 1908 2387
rect 2006 2384 2007 2388
rect 2011 2384 2012 2388
rect 2006 2383 2012 2384
rect 1902 2382 1908 2383
rect 110 2371 116 2372
rect 110 2367 111 2371
rect 115 2367 116 2371
rect 2006 2371 2012 2372
rect 110 2366 116 2367
rect 534 2368 540 2369
rect 534 2364 535 2368
rect 539 2364 540 2368
rect 534 2363 540 2364
rect 670 2368 676 2369
rect 670 2364 671 2368
rect 675 2364 676 2368
rect 670 2363 676 2364
rect 814 2368 820 2369
rect 814 2364 815 2368
rect 819 2364 820 2368
rect 814 2363 820 2364
rect 958 2368 964 2369
rect 958 2364 959 2368
rect 963 2364 964 2368
rect 958 2363 964 2364
rect 1102 2368 1108 2369
rect 1102 2364 1103 2368
rect 1107 2364 1108 2368
rect 1102 2363 1108 2364
rect 1246 2368 1252 2369
rect 1246 2364 1247 2368
rect 1251 2364 1252 2368
rect 1246 2363 1252 2364
rect 1390 2368 1396 2369
rect 1390 2364 1391 2368
rect 1395 2364 1396 2368
rect 1390 2363 1396 2364
rect 1526 2368 1532 2369
rect 1526 2364 1527 2368
rect 1531 2364 1532 2368
rect 1526 2363 1532 2364
rect 1654 2368 1660 2369
rect 1654 2364 1655 2368
rect 1659 2364 1660 2368
rect 1654 2363 1660 2364
rect 1790 2368 1796 2369
rect 1790 2364 1791 2368
rect 1795 2364 1796 2368
rect 1790 2363 1796 2364
rect 1902 2368 1908 2369
rect 1902 2364 1903 2368
rect 1907 2364 1908 2368
rect 2006 2367 2007 2371
rect 2011 2367 2012 2371
rect 2006 2366 2012 2367
rect 1902 2363 1908 2364
rect 2166 2336 2172 2337
rect 2046 2333 2052 2334
rect 2046 2329 2047 2333
rect 2051 2329 2052 2333
rect 2166 2332 2167 2336
rect 2171 2332 2172 2336
rect 2166 2331 2172 2332
rect 2358 2336 2364 2337
rect 2358 2332 2359 2336
rect 2363 2332 2364 2336
rect 2358 2331 2364 2332
rect 2534 2336 2540 2337
rect 2534 2332 2535 2336
rect 2539 2332 2540 2336
rect 2534 2331 2540 2332
rect 2702 2336 2708 2337
rect 2702 2332 2703 2336
rect 2707 2332 2708 2336
rect 2702 2331 2708 2332
rect 2870 2336 2876 2337
rect 2870 2332 2871 2336
rect 2875 2332 2876 2336
rect 2870 2331 2876 2332
rect 3030 2336 3036 2337
rect 3030 2332 3031 2336
rect 3035 2332 3036 2336
rect 3030 2331 3036 2332
rect 3198 2336 3204 2337
rect 3198 2332 3199 2336
rect 3203 2332 3204 2336
rect 3198 2331 3204 2332
rect 3942 2333 3948 2334
rect 2046 2328 2052 2329
rect 3942 2329 3943 2333
rect 3947 2329 3948 2333
rect 3942 2328 3948 2329
rect 2166 2317 2172 2318
rect 2046 2316 2052 2317
rect 2046 2312 2047 2316
rect 2051 2312 2052 2316
rect 2166 2313 2167 2317
rect 2171 2313 2172 2317
rect 2166 2312 2172 2313
rect 2358 2317 2364 2318
rect 2358 2313 2359 2317
rect 2363 2313 2364 2317
rect 2358 2312 2364 2313
rect 2534 2317 2540 2318
rect 2534 2313 2535 2317
rect 2539 2313 2540 2317
rect 2534 2312 2540 2313
rect 2702 2317 2708 2318
rect 2702 2313 2703 2317
rect 2707 2313 2708 2317
rect 2702 2312 2708 2313
rect 2870 2317 2876 2318
rect 2870 2313 2871 2317
rect 2875 2313 2876 2317
rect 2870 2312 2876 2313
rect 3030 2317 3036 2318
rect 3030 2313 3031 2317
rect 3035 2313 3036 2317
rect 3030 2312 3036 2313
rect 3198 2317 3204 2318
rect 3198 2313 3199 2317
rect 3203 2313 3204 2317
rect 3198 2312 3204 2313
rect 3942 2316 3948 2317
rect 3942 2312 3943 2316
rect 3947 2312 3948 2316
rect 2046 2311 2052 2312
rect 3942 2311 3948 2312
rect 534 2304 540 2305
rect 110 2301 116 2302
rect 110 2297 111 2301
rect 115 2297 116 2301
rect 534 2300 535 2304
rect 539 2300 540 2304
rect 534 2299 540 2300
rect 646 2304 652 2305
rect 646 2300 647 2304
rect 651 2300 652 2304
rect 646 2299 652 2300
rect 766 2304 772 2305
rect 766 2300 767 2304
rect 771 2300 772 2304
rect 766 2299 772 2300
rect 894 2304 900 2305
rect 894 2300 895 2304
rect 899 2300 900 2304
rect 894 2299 900 2300
rect 1030 2304 1036 2305
rect 1030 2300 1031 2304
rect 1035 2300 1036 2304
rect 1030 2299 1036 2300
rect 1166 2304 1172 2305
rect 1166 2300 1167 2304
rect 1171 2300 1172 2304
rect 1166 2299 1172 2300
rect 1294 2304 1300 2305
rect 1294 2300 1295 2304
rect 1299 2300 1300 2304
rect 1294 2299 1300 2300
rect 1422 2304 1428 2305
rect 1422 2300 1423 2304
rect 1427 2300 1428 2304
rect 1422 2299 1428 2300
rect 1550 2304 1556 2305
rect 1550 2300 1551 2304
rect 1555 2300 1556 2304
rect 1550 2299 1556 2300
rect 1670 2304 1676 2305
rect 1670 2300 1671 2304
rect 1675 2300 1676 2304
rect 1670 2299 1676 2300
rect 1798 2304 1804 2305
rect 1798 2300 1799 2304
rect 1803 2300 1804 2304
rect 1798 2299 1804 2300
rect 1902 2304 1908 2305
rect 1902 2300 1903 2304
rect 1907 2300 1908 2304
rect 1902 2299 1908 2300
rect 2006 2301 2012 2302
rect 110 2296 116 2297
rect 2006 2297 2007 2301
rect 2011 2297 2012 2301
rect 2006 2296 2012 2297
rect 534 2285 540 2286
rect 110 2284 116 2285
rect 110 2280 111 2284
rect 115 2280 116 2284
rect 534 2281 535 2285
rect 539 2281 540 2285
rect 534 2280 540 2281
rect 646 2285 652 2286
rect 646 2281 647 2285
rect 651 2281 652 2285
rect 646 2280 652 2281
rect 766 2285 772 2286
rect 766 2281 767 2285
rect 771 2281 772 2285
rect 766 2280 772 2281
rect 894 2285 900 2286
rect 894 2281 895 2285
rect 899 2281 900 2285
rect 894 2280 900 2281
rect 1030 2285 1036 2286
rect 1030 2281 1031 2285
rect 1035 2281 1036 2285
rect 1030 2280 1036 2281
rect 1166 2285 1172 2286
rect 1166 2281 1167 2285
rect 1171 2281 1172 2285
rect 1166 2280 1172 2281
rect 1294 2285 1300 2286
rect 1294 2281 1295 2285
rect 1299 2281 1300 2285
rect 1294 2280 1300 2281
rect 1422 2285 1428 2286
rect 1422 2281 1423 2285
rect 1427 2281 1428 2285
rect 1422 2280 1428 2281
rect 1550 2285 1556 2286
rect 1550 2281 1551 2285
rect 1555 2281 1556 2285
rect 1550 2280 1556 2281
rect 1670 2285 1676 2286
rect 1670 2281 1671 2285
rect 1675 2281 1676 2285
rect 1670 2280 1676 2281
rect 1798 2285 1804 2286
rect 1798 2281 1799 2285
rect 1803 2281 1804 2285
rect 1798 2280 1804 2281
rect 1902 2285 1908 2286
rect 1902 2281 1903 2285
rect 1907 2281 1908 2285
rect 1902 2280 1908 2281
rect 2006 2284 2012 2285
rect 2006 2280 2007 2284
rect 2011 2280 2012 2284
rect 110 2279 116 2280
rect 2006 2279 2012 2280
rect 2046 2264 2052 2265
rect 3942 2264 3948 2265
rect 2046 2260 2047 2264
rect 2051 2260 2052 2264
rect 2046 2259 2052 2260
rect 2070 2263 2076 2264
rect 2070 2259 2071 2263
rect 2075 2259 2076 2263
rect 2070 2258 2076 2259
rect 2166 2263 2172 2264
rect 2166 2259 2167 2263
rect 2171 2259 2172 2263
rect 2166 2258 2172 2259
rect 2286 2263 2292 2264
rect 2286 2259 2287 2263
rect 2291 2259 2292 2263
rect 2286 2258 2292 2259
rect 2422 2263 2428 2264
rect 2422 2259 2423 2263
rect 2427 2259 2428 2263
rect 2422 2258 2428 2259
rect 2558 2263 2564 2264
rect 2558 2259 2559 2263
rect 2563 2259 2564 2263
rect 2558 2258 2564 2259
rect 2702 2263 2708 2264
rect 2702 2259 2703 2263
rect 2707 2259 2708 2263
rect 2702 2258 2708 2259
rect 2838 2263 2844 2264
rect 2838 2259 2839 2263
rect 2843 2259 2844 2263
rect 2838 2258 2844 2259
rect 2982 2263 2988 2264
rect 2982 2259 2983 2263
rect 2987 2259 2988 2263
rect 2982 2258 2988 2259
rect 3126 2263 3132 2264
rect 3126 2259 3127 2263
rect 3131 2259 3132 2263
rect 3126 2258 3132 2259
rect 3270 2263 3276 2264
rect 3270 2259 3271 2263
rect 3275 2259 3276 2263
rect 3942 2260 3943 2264
rect 3947 2260 3948 2264
rect 3942 2259 3948 2260
rect 3270 2258 3276 2259
rect 2046 2247 2052 2248
rect 2046 2243 2047 2247
rect 2051 2243 2052 2247
rect 3942 2247 3948 2248
rect 2046 2242 2052 2243
rect 2070 2244 2076 2245
rect 2070 2240 2071 2244
rect 2075 2240 2076 2244
rect 2070 2239 2076 2240
rect 2166 2244 2172 2245
rect 2166 2240 2167 2244
rect 2171 2240 2172 2244
rect 2166 2239 2172 2240
rect 2286 2244 2292 2245
rect 2286 2240 2287 2244
rect 2291 2240 2292 2244
rect 2286 2239 2292 2240
rect 2422 2244 2428 2245
rect 2422 2240 2423 2244
rect 2427 2240 2428 2244
rect 2422 2239 2428 2240
rect 2558 2244 2564 2245
rect 2558 2240 2559 2244
rect 2563 2240 2564 2244
rect 2558 2239 2564 2240
rect 2702 2244 2708 2245
rect 2702 2240 2703 2244
rect 2707 2240 2708 2244
rect 2702 2239 2708 2240
rect 2838 2244 2844 2245
rect 2838 2240 2839 2244
rect 2843 2240 2844 2244
rect 2838 2239 2844 2240
rect 2982 2244 2988 2245
rect 2982 2240 2983 2244
rect 2987 2240 2988 2244
rect 2982 2239 2988 2240
rect 3126 2244 3132 2245
rect 3126 2240 3127 2244
rect 3131 2240 3132 2244
rect 3126 2239 3132 2240
rect 3270 2244 3276 2245
rect 3270 2240 3271 2244
rect 3275 2240 3276 2244
rect 3942 2243 3943 2247
rect 3947 2243 3948 2247
rect 3942 2242 3948 2243
rect 3270 2239 3276 2240
rect 110 2228 116 2229
rect 2006 2228 2012 2229
rect 110 2224 111 2228
rect 115 2224 116 2228
rect 110 2223 116 2224
rect 414 2227 420 2228
rect 414 2223 415 2227
rect 419 2223 420 2227
rect 414 2222 420 2223
rect 534 2227 540 2228
rect 534 2223 535 2227
rect 539 2223 540 2227
rect 534 2222 540 2223
rect 670 2227 676 2228
rect 670 2223 671 2227
rect 675 2223 676 2227
rect 670 2222 676 2223
rect 822 2227 828 2228
rect 822 2223 823 2227
rect 827 2223 828 2227
rect 822 2222 828 2223
rect 990 2227 996 2228
rect 990 2223 991 2227
rect 995 2223 996 2227
rect 990 2222 996 2223
rect 1174 2227 1180 2228
rect 1174 2223 1175 2227
rect 1179 2223 1180 2227
rect 1174 2222 1180 2223
rect 1366 2227 1372 2228
rect 1366 2223 1367 2227
rect 1371 2223 1372 2227
rect 1366 2222 1372 2223
rect 1566 2227 1572 2228
rect 1566 2223 1567 2227
rect 1571 2223 1572 2227
rect 1566 2222 1572 2223
rect 1766 2227 1772 2228
rect 1766 2223 1767 2227
rect 1771 2223 1772 2227
rect 2006 2224 2007 2228
rect 2011 2224 2012 2228
rect 2006 2223 2012 2224
rect 1766 2222 1772 2223
rect 110 2211 116 2212
rect 110 2207 111 2211
rect 115 2207 116 2211
rect 2006 2211 2012 2212
rect 110 2206 116 2207
rect 414 2208 420 2209
rect 414 2204 415 2208
rect 419 2204 420 2208
rect 414 2203 420 2204
rect 534 2208 540 2209
rect 534 2204 535 2208
rect 539 2204 540 2208
rect 534 2203 540 2204
rect 670 2208 676 2209
rect 670 2204 671 2208
rect 675 2204 676 2208
rect 670 2203 676 2204
rect 822 2208 828 2209
rect 822 2204 823 2208
rect 827 2204 828 2208
rect 822 2203 828 2204
rect 990 2208 996 2209
rect 990 2204 991 2208
rect 995 2204 996 2208
rect 990 2203 996 2204
rect 1174 2208 1180 2209
rect 1174 2204 1175 2208
rect 1179 2204 1180 2208
rect 1174 2203 1180 2204
rect 1366 2208 1372 2209
rect 1366 2204 1367 2208
rect 1371 2204 1372 2208
rect 1366 2203 1372 2204
rect 1566 2208 1572 2209
rect 1566 2204 1567 2208
rect 1571 2204 1572 2208
rect 1566 2203 1572 2204
rect 1766 2208 1772 2209
rect 1766 2204 1767 2208
rect 1771 2204 1772 2208
rect 2006 2207 2007 2211
rect 2011 2207 2012 2211
rect 2006 2206 2012 2207
rect 1766 2203 1772 2204
rect 2070 2184 2076 2185
rect 2046 2181 2052 2182
rect 2046 2177 2047 2181
rect 2051 2177 2052 2181
rect 2070 2180 2071 2184
rect 2075 2180 2076 2184
rect 2070 2179 2076 2180
rect 2294 2184 2300 2185
rect 2294 2180 2295 2184
rect 2299 2180 2300 2184
rect 2294 2179 2300 2180
rect 2502 2184 2508 2185
rect 2502 2180 2503 2184
rect 2507 2180 2508 2184
rect 2502 2179 2508 2180
rect 2686 2184 2692 2185
rect 2686 2180 2687 2184
rect 2691 2180 2692 2184
rect 2686 2179 2692 2180
rect 2862 2184 2868 2185
rect 2862 2180 2863 2184
rect 2867 2180 2868 2184
rect 2862 2179 2868 2180
rect 3022 2184 3028 2185
rect 3022 2180 3023 2184
rect 3027 2180 3028 2184
rect 3022 2179 3028 2180
rect 3174 2184 3180 2185
rect 3174 2180 3175 2184
rect 3179 2180 3180 2184
rect 3174 2179 3180 2180
rect 3318 2184 3324 2185
rect 3318 2180 3319 2184
rect 3323 2180 3324 2184
rect 3318 2179 3324 2180
rect 3470 2184 3476 2185
rect 3470 2180 3471 2184
rect 3475 2180 3476 2184
rect 3470 2179 3476 2180
rect 3942 2181 3948 2182
rect 2046 2176 2052 2177
rect 3942 2177 3943 2181
rect 3947 2177 3948 2181
rect 3942 2176 3948 2177
rect 2070 2165 2076 2166
rect 2046 2164 2052 2165
rect 2046 2160 2047 2164
rect 2051 2160 2052 2164
rect 2070 2161 2071 2165
rect 2075 2161 2076 2165
rect 2070 2160 2076 2161
rect 2294 2165 2300 2166
rect 2294 2161 2295 2165
rect 2299 2161 2300 2165
rect 2294 2160 2300 2161
rect 2502 2165 2508 2166
rect 2502 2161 2503 2165
rect 2507 2161 2508 2165
rect 2502 2160 2508 2161
rect 2686 2165 2692 2166
rect 2686 2161 2687 2165
rect 2691 2161 2692 2165
rect 2686 2160 2692 2161
rect 2862 2165 2868 2166
rect 2862 2161 2863 2165
rect 2867 2161 2868 2165
rect 2862 2160 2868 2161
rect 3022 2165 3028 2166
rect 3022 2161 3023 2165
rect 3027 2161 3028 2165
rect 3022 2160 3028 2161
rect 3174 2165 3180 2166
rect 3174 2161 3175 2165
rect 3179 2161 3180 2165
rect 3174 2160 3180 2161
rect 3318 2165 3324 2166
rect 3318 2161 3319 2165
rect 3323 2161 3324 2165
rect 3318 2160 3324 2161
rect 3470 2165 3476 2166
rect 3470 2161 3471 2165
rect 3475 2161 3476 2165
rect 3470 2160 3476 2161
rect 3942 2164 3948 2165
rect 3942 2160 3943 2164
rect 3947 2160 3948 2164
rect 2046 2159 2052 2160
rect 3942 2159 3948 2160
rect 134 2140 140 2141
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 134 2136 135 2140
rect 139 2136 140 2140
rect 134 2135 140 2136
rect 246 2140 252 2141
rect 246 2136 247 2140
rect 251 2136 252 2140
rect 246 2135 252 2136
rect 390 2140 396 2141
rect 390 2136 391 2140
rect 395 2136 396 2140
rect 390 2135 396 2136
rect 550 2140 556 2141
rect 550 2136 551 2140
rect 555 2136 556 2140
rect 550 2135 556 2136
rect 710 2140 716 2141
rect 710 2136 711 2140
rect 715 2136 716 2140
rect 710 2135 716 2136
rect 870 2140 876 2141
rect 870 2136 871 2140
rect 875 2136 876 2140
rect 870 2135 876 2136
rect 1030 2140 1036 2141
rect 1030 2136 1031 2140
rect 1035 2136 1036 2140
rect 1030 2135 1036 2136
rect 1190 2140 1196 2141
rect 1190 2136 1191 2140
rect 1195 2136 1196 2140
rect 1190 2135 1196 2136
rect 1350 2140 1356 2141
rect 1350 2136 1351 2140
rect 1355 2136 1356 2140
rect 1350 2135 1356 2136
rect 1510 2140 1516 2141
rect 1510 2136 1511 2140
rect 1515 2136 1516 2140
rect 1510 2135 1516 2136
rect 1678 2140 1684 2141
rect 1678 2136 1679 2140
rect 1683 2136 1684 2140
rect 1678 2135 1684 2136
rect 2006 2137 2012 2138
rect 110 2132 116 2133
rect 2006 2133 2007 2137
rect 2011 2133 2012 2137
rect 2006 2132 2012 2133
rect 134 2121 140 2122
rect 110 2120 116 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 134 2117 135 2121
rect 139 2117 140 2121
rect 134 2116 140 2117
rect 246 2121 252 2122
rect 246 2117 247 2121
rect 251 2117 252 2121
rect 246 2116 252 2117
rect 390 2121 396 2122
rect 390 2117 391 2121
rect 395 2117 396 2121
rect 390 2116 396 2117
rect 550 2121 556 2122
rect 550 2117 551 2121
rect 555 2117 556 2121
rect 550 2116 556 2117
rect 710 2121 716 2122
rect 710 2117 711 2121
rect 715 2117 716 2121
rect 710 2116 716 2117
rect 870 2121 876 2122
rect 870 2117 871 2121
rect 875 2117 876 2121
rect 870 2116 876 2117
rect 1030 2121 1036 2122
rect 1030 2117 1031 2121
rect 1035 2117 1036 2121
rect 1030 2116 1036 2117
rect 1190 2121 1196 2122
rect 1190 2117 1191 2121
rect 1195 2117 1196 2121
rect 1190 2116 1196 2117
rect 1350 2121 1356 2122
rect 1350 2117 1351 2121
rect 1355 2117 1356 2121
rect 1350 2116 1356 2117
rect 1510 2121 1516 2122
rect 1510 2117 1511 2121
rect 1515 2117 1516 2121
rect 1510 2116 1516 2117
rect 1678 2121 1684 2122
rect 1678 2117 1679 2121
rect 1683 2117 1684 2121
rect 1678 2116 1684 2117
rect 2006 2120 2012 2121
rect 2006 2116 2007 2120
rect 2011 2116 2012 2120
rect 110 2115 116 2116
rect 2006 2115 2012 2116
rect 2046 2088 2052 2089
rect 3942 2088 3948 2089
rect 2046 2084 2047 2088
rect 2051 2084 2052 2088
rect 2046 2083 2052 2084
rect 2398 2087 2404 2088
rect 2398 2083 2399 2087
rect 2403 2083 2404 2087
rect 2398 2082 2404 2083
rect 2494 2087 2500 2088
rect 2494 2083 2495 2087
rect 2499 2083 2500 2087
rect 2494 2082 2500 2083
rect 2590 2087 2596 2088
rect 2590 2083 2591 2087
rect 2595 2083 2596 2087
rect 2590 2082 2596 2083
rect 2686 2087 2692 2088
rect 2686 2083 2687 2087
rect 2691 2083 2692 2087
rect 2686 2082 2692 2083
rect 2782 2087 2788 2088
rect 2782 2083 2783 2087
rect 2787 2083 2788 2087
rect 2782 2082 2788 2083
rect 2878 2087 2884 2088
rect 2878 2083 2879 2087
rect 2883 2083 2884 2087
rect 2878 2082 2884 2083
rect 2974 2087 2980 2088
rect 2974 2083 2975 2087
rect 2979 2083 2980 2087
rect 2974 2082 2980 2083
rect 3070 2087 3076 2088
rect 3070 2083 3071 2087
rect 3075 2083 3076 2087
rect 3070 2082 3076 2083
rect 3166 2087 3172 2088
rect 3166 2083 3167 2087
rect 3171 2083 3172 2087
rect 3166 2082 3172 2083
rect 3262 2087 3268 2088
rect 3262 2083 3263 2087
rect 3267 2083 3268 2087
rect 3262 2082 3268 2083
rect 3358 2087 3364 2088
rect 3358 2083 3359 2087
rect 3363 2083 3364 2087
rect 3358 2082 3364 2083
rect 3454 2087 3460 2088
rect 3454 2083 3455 2087
rect 3459 2083 3460 2087
rect 3454 2082 3460 2083
rect 3550 2087 3556 2088
rect 3550 2083 3551 2087
rect 3555 2083 3556 2087
rect 3550 2082 3556 2083
rect 3646 2087 3652 2088
rect 3646 2083 3647 2087
rect 3651 2083 3652 2087
rect 3646 2082 3652 2083
rect 3742 2087 3748 2088
rect 3742 2083 3743 2087
rect 3747 2083 3748 2087
rect 3742 2082 3748 2083
rect 3838 2087 3844 2088
rect 3838 2083 3839 2087
rect 3843 2083 3844 2087
rect 3942 2084 3943 2088
rect 3947 2084 3948 2088
rect 3942 2083 3948 2084
rect 3838 2082 3844 2083
rect 2046 2071 2052 2072
rect 2046 2067 2047 2071
rect 2051 2067 2052 2071
rect 3942 2071 3948 2072
rect 2046 2066 2052 2067
rect 2398 2068 2404 2069
rect 2398 2064 2399 2068
rect 2403 2064 2404 2068
rect 2398 2063 2404 2064
rect 2494 2068 2500 2069
rect 2494 2064 2495 2068
rect 2499 2064 2500 2068
rect 2494 2063 2500 2064
rect 2590 2068 2596 2069
rect 2590 2064 2591 2068
rect 2595 2064 2596 2068
rect 2590 2063 2596 2064
rect 2686 2068 2692 2069
rect 2686 2064 2687 2068
rect 2691 2064 2692 2068
rect 2686 2063 2692 2064
rect 2782 2068 2788 2069
rect 2782 2064 2783 2068
rect 2787 2064 2788 2068
rect 2782 2063 2788 2064
rect 2878 2068 2884 2069
rect 2878 2064 2879 2068
rect 2883 2064 2884 2068
rect 2878 2063 2884 2064
rect 2974 2068 2980 2069
rect 2974 2064 2975 2068
rect 2979 2064 2980 2068
rect 2974 2063 2980 2064
rect 3070 2068 3076 2069
rect 3070 2064 3071 2068
rect 3075 2064 3076 2068
rect 3070 2063 3076 2064
rect 3166 2068 3172 2069
rect 3166 2064 3167 2068
rect 3171 2064 3172 2068
rect 3166 2063 3172 2064
rect 3262 2068 3268 2069
rect 3262 2064 3263 2068
rect 3267 2064 3268 2068
rect 3262 2063 3268 2064
rect 3358 2068 3364 2069
rect 3358 2064 3359 2068
rect 3363 2064 3364 2068
rect 3358 2063 3364 2064
rect 3454 2068 3460 2069
rect 3454 2064 3455 2068
rect 3459 2064 3460 2068
rect 3454 2063 3460 2064
rect 3550 2068 3556 2069
rect 3550 2064 3551 2068
rect 3555 2064 3556 2068
rect 3550 2063 3556 2064
rect 3646 2068 3652 2069
rect 3646 2064 3647 2068
rect 3651 2064 3652 2068
rect 3646 2063 3652 2064
rect 3742 2068 3748 2069
rect 3742 2064 3743 2068
rect 3747 2064 3748 2068
rect 3742 2063 3748 2064
rect 3838 2068 3844 2069
rect 3838 2064 3839 2068
rect 3843 2064 3844 2068
rect 3942 2067 3943 2071
rect 3947 2067 3948 2071
rect 3942 2066 3948 2067
rect 3838 2063 3844 2064
rect 110 2060 116 2061
rect 2006 2060 2012 2061
rect 110 2056 111 2060
rect 115 2056 116 2060
rect 110 2055 116 2056
rect 134 2059 140 2060
rect 134 2055 135 2059
rect 139 2055 140 2059
rect 134 2054 140 2055
rect 246 2059 252 2060
rect 246 2055 247 2059
rect 251 2055 252 2059
rect 246 2054 252 2055
rect 398 2059 404 2060
rect 398 2055 399 2059
rect 403 2055 404 2059
rect 398 2054 404 2055
rect 550 2059 556 2060
rect 550 2055 551 2059
rect 555 2055 556 2059
rect 550 2054 556 2055
rect 702 2059 708 2060
rect 702 2055 703 2059
rect 707 2055 708 2059
rect 702 2054 708 2055
rect 846 2059 852 2060
rect 846 2055 847 2059
rect 851 2055 852 2059
rect 846 2054 852 2055
rect 990 2059 996 2060
rect 990 2055 991 2059
rect 995 2055 996 2059
rect 990 2054 996 2055
rect 1126 2059 1132 2060
rect 1126 2055 1127 2059
rect 1131 2055 1132 2059
rect 1126 2054 1132 2055
rect 1254 2059 1260 2060
rect 1254 2055 1255 2059
rect 1259 2055 1260 2059
rect 1254 2054 1260 2055
rect 1382 2059 1388 2060
rect 1382 2055 1383 2059
rect 1387 2055 1388 2059
rect 1382 2054 1388 2055
rect 1518 2059 1524 2060
rect 1518 2055 1519 2059
rect 1523 2055 1524 2059
rect 2006 2056 2007 2060
rect 2011 2056 2012 2060
rect 2006 2055 2012 2056
rect 1518 2054 1524 2055
rect 110 2043 116 2044
rect 110 2039 111 2043
rect 115 2039 116 2043
rect 2006 2043 2012 2044
rect 110 2038 116 2039
rect 134 2040 140 2041
rect 134 2036 135 2040
rect 139 2036 140 2040
rect 134 2035 140 2036
rect 246 2040 252 2041
rect 246 2036 247 2040
rect 251 2036 252 2040
rect 246 2035 252 2036
rect 398 2040 404 2041
rect 398 2036 399 2040
rect 403 2036 404 2040
rect 398 2035 404 2036
rect 550 2040 556 2041
rect 550 2036 551 2040
rect 555 2036 556 2040
rect 550 2035 556 2036
rect 702 2040 708 2041
rect 702 2036 703 2040
rect 707 2036 708 2040
rect 702 2035 708 2036
rect 846 2040 852 2041
rect 846 2036 847 2040
rect 851 2036 852 2040
rect 846 2035 852 2036
rect 990 2040 996 2041
rect 990 2036 991 2040
rect 995 2036 996 2040
rect 990 2035 996 2036
rect 1126 2040 1132 2041
rect 1126 2036 1127 2040
rect 1131 2036 1132 2040
rect 1126 2035 1132 2036
rect 1254 2040 1260 2041
rect 1254 2036 1255 2040
rect 1259 2036 1260 2040
rect 1254 2035 1260 2036
rect 1382 2040 1388 2041
rect 1382 2036 1383 2040
rect 1387 2036 1388 2040
rect 1382 2035 1388 2036
rect 1518 2040 1524 2041
rect 1518 2036 1519 2040
rect 1523 2036 1524 2040
rect 2006 2039 2007 2043
rect 2011 2039 2012 2043
rect 2006 2038 2012 2039
rect 1518 2035 1524 2036
rect 2190 2008 2196 2009
rect 2046 2005 2052 2006
rect 2046 2001 2047 2005
rect 2051 2001 2052 2005
rect 2190 2004 2191 2008
rect 2195 2004 2196 2008
rect 2190 2003 2196 2004
rect 2398 2008 2404 2009
rect 2398 2004 2399 2008
rect 2403 2004 2404 2008
rect 2398 2003 2404 2004
rect 2646 2008 2652 2009
rect 2646 2004 2647 2008
rect 2651 2004 2652 2008
rect 2646 2003 2652 2004
rect 2918 2008 2924 2009
rect 2918 2004 2919 2008
rect 2923 2004 2924 2008
rect 2918 2003 2924 2004
rect 3214 2008 3220 2009
rect 3214 2004 3215 2008
rect 3219 2004 3220 2008
rect 3214 2003 3220 2004
rect 3526 2008 3532 2009
rect 3526 2004 3527 2008
rect 3531 2004 3532 2008
rect 3526 2003 3532 2004
rect 3838 2008 3844 2009
rect 3838 2004 3839 2008
rect 3843 2004 3844 2008
rect 3838 2003 3844 2004
rect 3942 2005 3948 2006
rect 2046 2000 2052 2001
rect 3942 2001 3943 2005
rect 3947 2001 3948 2005
rect 3942 2000 3948 2001
rect 2190 1989 2196 1990
rect 2046 1988 2052 1989
rect 2046 1984 2047 1988
rect 2051 1984 2052 1988
rect 2190 1985 2191 1989
rect 2195 1985 2196 1989
rect 2190 1984 2196 1985
rect 2398 1989 2404 1990
rect 2398 1985 2399 1989
rect 2403 1985 2404 1989
rect 2398 1984 2404 1985
rect 2646 1989 2652 1990
rect 2646 1985 2647 1989
rect 2651 1985 2652 1989
rect 2646 1984 2652 1985
rect 2918 1989 2924 1990
rect 2918 1985 2919 1989
rect 2923 1985 2924 1989
rect 2918 1984 2924 1985
rect 3214 1989 3220 1990
rect 3214 1985 3215 1989
rect 3219 1985 3220 1989
rect 3214 1984 3220 1985
rect 3526 1989 3532 1990
rect 3526 1985 3527 1989
rect 3531 1985 3532 1989
rect 3526 1984 3532 1985
rect 3838 1989 3844 1990
rect 3838 1985 3839 1989
rect 3843 1985 3844 1989
rect 3838 1984 3844 1985
rect 3942 1988 3948 1989
rect 3942 1984 3943 1988
rect 3947 1984 3948 1988
rect 2046 1983 2052 1984
rect 3942 1983 3948 1984
rect 230 1964 236 1965
rect 110 1961 116 1962
rect 110 1957 111 1961
rect 115 1957 116 1961
rect 230 1960 231 1964
rect 235 1960 236 1964
rect 230 1959 236 1960
rect 390 1964 396 1965
rect 390 1960 391 1964
rect 395 1960 396 1964
rect 390 1959 396 1960
rect 566 1964 572 1965
rect 566 1960 567 1964
rect 571 1960 572 1964
rect 566 1959 572 1960
rect 750 1964 756 1965
rect 750 1960 751 1964
rect 755 1960 756 1964
rect 750 1959 756 1960
rect 942 1964 948 1965
rect 942 1960 943 1964
rect 947 1960 948 1964
rect 942 1959 948 1960
rect 1134 1964 1140 1965
rect 1134 1960 1135 1964
rect 1139 1960 1140 1964
rect 1134 1959 1140 1960
rect 1334 1964 1340 1965
rect 1334 1960 1335 1964
rect 1339 1960 1340 1964
rect 1334 1959 1340 1960
rect 1542 1964 1548 1965
rect 1542 1960 1543 1964
rect 1547 1960 1548 1964
rect 1542 1959 1548 1960
rect 2006 1961 2012 1962
rect 110 1956 116 1957
rect 2006 1957 2007 1961
rect 2011 1957 2012 1961
rect 2006 1956 2012 1957
rect 230 1945 236 1946
rect 110 1944 116 1945
rect 110 1940 111 1944
rect 115 1940 116 1944
rect 230 1941 231 1945
rect 235 1941 236 1945
rect 230 1940 236 1941
rect 390 1945 396 1946
rect 390 1941 391 1945
rect 395 1941 396 1945
rect 390 1940 396 1941
rect 566 1945 572 1946
rect 566 1941 567 1945
rect 571 1941 572 1945
rect 566 1940 572 1941
rect 750 1945 756 1946
rect 750 1941 751 1945
rect 755 1941 756 1945
rect 750 1940 756 1941
rect 942 1945 948 1946
rect 942 1941 943 1945
rect 947 1941 948 1945
rect 942 1940 948 1941
rect 1134 1945 1140 1946
rect 1134 1941 1135 1945
rect 1139 1941 1140 1945
rect 1134 1940 1140 1941
rect 1334 1945 1340 1946
rect 1334 1941 1335 1945
rect 1339 1941 1340 1945
rect 1334 1940 1340 1941
rect 1542 1945 1548 1946
rect 1542 1941 1543 1945
rect 1547 1941 1548 1945
rect 1542 1940 1548 1941
rect 2006 1944 2012 1945
rect 2006 1940 2007 1944
rect 2011 1940 2012 1944
rect 110 1939 116 1940
rect 2006 1939 2012 1940
rect 2046 1924 2052 1925
rect 3942 1924 3948 1925
rect 2046 1920 2047 1924
rect 2051 1920 2052 1924
rect 2046 1919 2052 1920
rect 2070 1923 2076 1924
rect 2070 1919 2071 1923
rect 2075 1919 2076 1923
rect 2070 1918 2076 1919
rect 2238 1923 2244 1924
rect 2238 1919 2239 1923
rect 2243 1919 2244 1923
rect 2238 1918 2244 1919
rect 2446 1923 2452 1924
rect 2446 1919 2447 1923
rect 2451 1919 2452 1923
rect 2446 1918 2452 1919
rect 2670 1923 2676 1924
rect 2670 1919 2671 1923
rect 2675 1919 2676 1923
rect 2670 1918 2676 1919
rect 2894 1923 2900 1924
rect 2894 1919 2895 1923
rect 2899 1919 2900 1923
rect 2894 1918 2900 1919
rect 3126 1923 3132 1924
rect 3126 1919 3127 1923
rect 3131 1919 3132 1923
rect 3126 1918 3132 1919
rect 3358 1923 3364 1924
rect 3358 1919 3359 1923
rect 3363 1919 3364 1923
rect 3358 1918 3364 1919
rect 3590 1923 3596 1924
rect 3590 1919 3591 1923
rect 3595 1919 3596 1923
rect 3590 1918 3596 1919
rect 3830 1923 3836 1924
rect 3830 1919 3831 1923
rect 3835 1919 3836 1923
rect 3942 1920 3943 1924
rect 3947 1920 3948 1924
rect 3942 1919 3948 1920
rect 3830 1918 3836 1919
rect 2046 1907 2052 1908
rect 2046 1903 2047 1907
rect 2051 1903 2052 1907
rect 3942 1907 3948 1908
rect 2046 1902 2052 1903
rect 2070 1904 2076 1905
rect 2070 1900 2071 1904
rect 2075 1900 2076 1904
rect 2070 1899 2076 1900
rect 2238 1904 2244 1905
rect 2238 1900 2239 1904
rect 2243 1900 2244 1904
rect 2238 1899 2244 1900
rect 2446 1904 2452 1905
rect 2446 1900 2447 1904
rect 2451 1900 2452 1904
rect 2446 1899 2452 1900
rect 2670 1904 2676 1905
rect 2670 1900 2671 1904
rect 2675 1900 2676 1904
rect 2670 1899 2676 1900
rect 2894 1904 2900 1905
rect 2894 1900 2895 1904
rect 2899 1900 2900 1904
rect 2894 1899 2900 1900
rect 3126 1904 3132 1905
rect 3126 1900 3127 1904
rect 3131 1900 3132 1904
rect 3126 1899 3132 1900
rect 3358 1904 3364 1905
rect 3358 1900 3359 1904
rect 3363 1900 3364 1904
rect 3358 1899 3364 1900
rect 3590 1904 3596 1905
rect 3590 1900 3591 1904
rect 3595 1900 3596 1904
rect 3590 1899 3596 1900
rect 3830 1904 3836 1905
rect 3830 1900 3831 1904
rect 3835 1900 3836 1904
rect 3942 1903 3943 1907
rect 3947 1903 3948 1907
rect 3942 1902 3948 1903
rect 3830 1899 3836 1900
rect 110 1892 116 1893
rect 2006 1892 2012 1893
rect 110 1888 111 1892
rect 115 1888 116 1892
rect 110 1887 116 1888
rect 510 1891 516 1892
rect 510 1887 511 1891
rect 515 1887 516 1891
rect 510 1886 516 1887
rect 622 1891 628 1892
rect 622 1887 623 1891
rect 627 1887 628 1891
rect 622 1886 628 1887
rect 742 1891 748 1892
rect 742 1887 743 1891
rect 747 1887 748 1891
rect 742 1886 748 1887
rect 862 1891 868 1892
rect 862 1887 863 1891
rect 867 1887 868 1891
rect 862 1886 868 1887
rect 982 1891 988 1892
rect 982 1887 983 1891
rect 987 1887 988 1891
rect 982 1886 988 1887
rect 1102 1891 1108 1892
rect 1102 1887 1103 1891
rect 1107 1887 1108 1891
rect 1102 1886 1108 1887
rect 1222 1891 1228 1892
rect 1222 1887 1223 1891
rect 1227 1887 1228 1891
rect 1222 1886 1228 1887
rect 1334 1891 1340 1892
rect 1334 1887 1335 1891
rect 1339 1887 1340 1891
rect 1334 1886 1340 1887
rect 1454 1891 1460 1892
rect 1454 1887 1455 1891
rect 1459 1887 1460 1891
rect 1454 1886 1460 1887
rect 1574 1891 1580 1892
rect 1574 1887 1575 1891
rect 1579 1887 1580 1891
rect 1574 1886 1580 1887
rect 1694 1891 1700 1892
rect 1694 1887 1695 1891
rect 1699 1887 1700 1891
rect 2006 1888 2007 1892
rect 2011 1888 2012 1892
rect 2006 1887 2012 1888
rect 1694 1886 1700 1887
rect 110 1875 116 1876
rect 110 1871 111 1875
rect 115 1871 116 1875
rect 2006 1875 2012 1876
rect 110 1870 116 1871
rect 510 1872 516 1873
rect 510 1868 511 1872
rect 515 1868 516 1872
rect 510 1867 516 1868
rect 622 1872 628 1873
rect 622 1868 623 1872
rect 627 1868 628 1872
rect 622 1867 628 1868
rect 742 1872 748 1873
rect 742 1868 743 1872
rect 747 1868 748 1872
rect 742 1867 748 1868
rect 862 1872 868 1873
rect 862 1868 863 1872
rect 867 1868 868 1872
rect 862 1867 868 1868
rect 982 1872 988 1873
rect 982 1868 983 1872
rect 987 1868 988 1872
rect 982 1867 988 1868
rect 1102 1872 1108 1873
rect 1102 1868 1103 1872
rect 1107 1868 1108 1872
rect 1102 1867 1108 1868
rect 1222 1872 1228 1873
rect 1222 1868 1223 1872
rect 1227 1868 1228 1872
rect 1222 1867 1228 1868
rect 1334 1872 1340 1873
rect 1334 1868 1335 1872
rect 1339 1868 1340 1872
rect 1334 1867 1340 1868
rect 1454 1872 1460 1873
rect 1454 1868 1455 1872
rect 1459 1868 1460 1872
rect 1454 1867 1460 1868
rect 1574 1872 1580 1873
rect 1574 1868 1575 1872
rect 1579 1868 1580 1872
rect 1574 1867 1580 1868
rect 1694 1872 1700 1873
rect 1694 1868 1695 1872
rect 1699 1868 1700 1872
rect 2006 1871 2007 1875
rect 2011 1871 2012 1875
rect 2006 1870 2012 1871
rect 1694 1867 1700 1868
rect 2070 1844 2076 1845
rect 2046 1841 2052 1842
rect 2046 1837 2047 1841
rect 2051 1837 2052 1841
rect 2070 1840 2071 1844
rect 2075 1840 2076 1844
rect 2070 1839 2076 1840
rect 2198 1844 2204 1845
rect 2198 1840 2199 1844
rect 2203 1840 2204 1844
rect 2198 1839 2204 1840
rect 2366 1844 2372 1845
rect 2366 1840 2367 1844
rect 2371 1840 2372 1844
rect 2366 1839 2372 1840
rect 2542 1844 2548 1845
rect 2542 1840 2543 1844
rect 2547 1840 2548 1844
rect 2542 1839 2548 1840
rect 2718 1844 2724 1845
rect 2718 1840 2719 1844
rect 2723 1840 2724 1844
rect 2718 1839 2724 1840
rect 2886 1844 2892 1845
rect 2886 1840 2887 1844
rect 2891 1840 2892 1844
rect 2886 1839 2892 1840
rect 3038 1844 3044 1845
rect 3038 1840 3039 1844
rect 3043 1840 3044 1844
rect 3038 1839 3044 1840
rect 3182 1844 3188 1845
rect 3182 1840 3183 1844
rect 3187 1840 3188 1844
rect 3182 1839 3188 1840
rect 3318 1844 3324 1845
rect 3318 1840 3319 1844
rect 3323 1840 3324 1844
rect 3318 1839 3324 1840
rect 3454 1844 3460 1845
rect 3454 1840 3455 1844
rect 3459 1840 3460 1844
rect 3454 1839 3460 1840
rect 3582 1844 3588 1845
rect 3582 1840 3583 1844
rect 3587 1840 3588 1844
rect 3582 1839 3588 1840
rect 3710 1844 3716 1845
rect 3710 1840 3711 1844
rect 3715 1840 3716 1844
rect 3710 1839 3716 1840
rect 3838 1844 3844 1845
rect 3838 1840 3839 1844
rect 3843 1840 3844 1844
rect 3838 1839 3844 1840
rect 3942 1841 3948 1842
rect 2046 1836 2052 1837
rect 3942 1837 3943 1841
rect 3947 1837 3948 1841
rect 3942 1836 3948 1837
rect 2070 1825 2076 1826
rect 2046 1824 2052 1825
rect 2046 1820 2047 1824
rect 2051 1820 2052 1824
rect 2070 1821 2071 1825
rect 2075 1821 2076 1825
rect 2070 1820 2076 1821
rect 2198 1825 2204 1826
rect 2198 1821 2199 1825
rect 2203 1821 2204 1825
rect 2198 1820 2204 1821
rect 2366 1825 2372 1826
rect 2366 1821 2367 1825
rect 2371 1821 2372 1825
rect 2366 1820 2372 1821
rect 2542 1825 2548 1826
rect 2542 1821 2543 1825
rect 2547 1821 2548 1825
rect 2542 1820 2548 1821
rect 2718 1825 2724 1826
rect 2718 1821 2719 1825
rect 2723 1821 2724 1825
rect 2718 1820 2724 1821
rect 2886 1825 2892 1826
rect 2886 1821 2887 1825
rect 2891 1821 2892 1825
rect 2886 1820 2892 1821
rect 3038 1825 3044 1826
rect 3038 1821 3039 1825
rect 3043 1821 3044 1825
rect 3038 1820 3044 1821
rect 3182 1825 3188 1826
rect 3182 1821 3183 1825
rect 3187 1821 3188 1825
rect 3182 1820 3188 1821
rect 3318 1825 3324 1826
rect 3318 1821 3319 1825
rect 3323 1821 3324 1825
rect 3318 1820 3324 1821
rect 3454 1825 3460 1826
rect 3454 1821 3455 1825
rect 3459 1821 3460 1825
rect 3454 1820 3460 1821
rect 3582 1825 3588 1826
rect 3582 1821 3583 1825
rect 3587 1821 3588 1825
rect 3582 1820 3588 1821
rect 3710 1825 3716 1826
rect 3710 1821 3711 1825
rect 3715 1821 3716 1825
rect 3710 1820 3716 1821
rect 3838 1825 3844 1826
rect 3838 1821 3839 1825
rect 3843 1821 3844 1825
rect 3838 1820 3844 1821
rect 3942 1824 3948 1825
rect 3942 1820 3943 1824
rect 3947 1820 3948 1824
rect 2046 1819 2052 1820
rect 3942 1819 3948 1820
rect 614 1804 620 1805
rect 110 1801 116 1802
rect 110 1797 111 1801
rect 115 1797 116 1801
rect 614 1800 615 1804
rect 619 1800 620 1804
rect 614 1799 620 1800
rect 710 1804 716 1805
rect 710 1800 711 1804
rect 715 1800 716 1804
rect 710 1799 716 1800
rect 814 1804 820 1805
rect 814 1800 815 1804
rect 819 1800 820 1804
rect 814 1799 820 1800
rect 926 1804 932 1805
rect 926 1800 927 1804
rect 931 1800 932 1804
rect 926 1799 932 1800
rect 1038 1804 1044 1805
rect 1038 1800 1039 1804
rect 1043 1800 1044 1804
rect 1038 1799 1044 1800
rect 1158 1804 1164 1805
rect 1158 1800 1159 1804
rect 1163 1800 1164 1804
rect 1158 1799 1164 1800
rect 1278 1804 1284 1805
rect 1278 1800 1279 1804
rect 1283 1800 1284 1804
rect 1278 1799 1284 1800
rect 1398 1804 1404 1805
rect 1398 1800 1399 1804
rect 1403 1800 1404 1804
rect 1398 1799 1404 1800
rect 1518 1804 1524 1805
rect 1518 1800 1519 1804
rect 1523 1800 1524 1804
rect 1518 1799 1524 1800
rect 1638 1804 1644 1805
rect 1638 1800 1639 1804
rect 1643 1800 1644 1804
rect 1638 1799 1644 1800
rect 2006 1801 2012 1802
rect 110 1796 116 1797
rect 2006 1797 2007 1801
rect 2011 1797 2012 1801
rect 2006 1796 2012 1797
rect 614 1785 620 1786
rect 110 1784 116 1785
rect 110 1780 111 1784
rect 115 1780 116 1784
rect 614 1781 615 1785
rect 619 1781 620 1785
rect 614 1780 620 1781
rect 710 1785 716 1786
rect 710 1781 711 1785
rect 715 1781 716 1785
rect 710 1780 716 1781
rect 814 1785 820 1786
rect 814 1781 815 1785
rect 819 1781 820 1785
rect 814 1780 820 1781
rect 926 1785 932 1786
rect 926 1781 927 1785
rect 931 1781 932 1785
rect 926 1780 932 1781
rect 1038 1785 1044 1786
rect 1038 1781 1039 1785
rect 1043 1781 1044 1785
rect 1038 1780 1044 1781
rect 1158 1785 1164 1786
rect 1158 1781 1159 1785
rect 1163 1781 1164 1785
rect 1158 1780 1164 1781
rect 1278 1785 1284 1786
rect 1278 1781 1279 1785
rect 1283 1781 1284 1785
rect 1278 1780 1284 1781
rect 1398 1785 1404 1786
rect 1398 1781 1399 1785
rect 1403 1781 1404 1785
rect 1398 1780 1404 1781
rect 1518 1785 1524 1786
rect 1518 1781 1519 1785
rect 1523 1781 1524 1785
rect 1518 1780 1524 1781
rect 1638 1785 1644 1786
rect 1638 1781 1639 1785
rect 1643 1781 1644 1785
rect 1638 1780 1644 1781
rect 2006 1784 2012 1785
rect 2006 1780 2007 1784
rect 2011 1780 2012 1784
rect 110 1779 116 1780
rect 2006 1779 2012 1780
rect 2046 1768 2052 1769
rect 3942 1768 3948 1769
rect 2046 1764 2047 1768
rect 2051 1764 2052 1768
rect 2046 1763 2052 1764
rect 2070 1767 2076 1768
rect 2070 1763 2071 1767
rect 2075 1763 2076 1767
rect 2070 1762 2076 1763
rect 2182 1767 2188 1768
rect 2182 1763 2183 1767
rect 2187 1763 2188 1767
rect 2182 1762 2188 1763
rect 2326 1767 2332 1768
rect 2326 1763 2327 1767
rect 2331 1763 2332 1767
rect 2326 1762 2332 1763
rect 2486 1767 2492 1768
rect 2486 1763 2487 1767
rect 2491 1763 2492 1767
rect 2486 1762 2492 1763
rect 2654 1767 2660 1768
rect 2654 1763 2655 1767
rect 2659 1763 2660 1767
rect 2654 1762 2660 1763
rect 2830 1767 2836 1768
rect 2830 1763 2831 1767
rect 2835 1763 2836 1767
rect 2830 1762 2836 1763
rect 3022 1767 3028 1768
rect 3022 1763 3023 1767
rect 3027 1763 3028 1767
rect 3022 1762 3028 1763
rect 3222 1767 3228 1768
rect 3222 1763 3223 1767
rect 3227 1763 3228 1767
rect 3222 1762 3228 1763
rect 3430 1767 3436 1768
rect 3430 1763 3431 1767
rect 3435 1763 3436 1767
rect 3430 1762 3436 1763
rect 3646 1767 3652 1768
rect 3646 1763 3647 1767
rect 3651 1763 3652 1767
rect 3646 1762 3652 1763
rect 3838 1767 3844 1768
rect 3838 1763 3839 1767
rect 3843 1763 3844 1767
rect 3942 1764 3943 1768
rect 3947 1764 3948 1768
rect 3942 1763 3948 1764
rect 3838 1762 3844 1763
rect 2046 1751 2052 1752
rect 2046 1747 2047 1751
rect 2051 1747 2052 1751
rect 3942 1751 3948 1752
rect 2046 1746 2052 1747
rect 2070 1748 2076 1749
rect 2070 1744 2071 1748
rect 2075 1744 2076 1748
rect 2070 1743 2076 1744
rect 2182 1748 2188 1749
rect 2182 1744 2183 1748
rect 2187 1744 2188 1748
rect 2182 1743 2188 1744
rect 2326 1748 2332 1749
rect 2326 1744 2327 1748
rect 2331 1744 2332 1748
rect 2326 1743 2332 1744
rect 2486 1748 2492 1749
rect 2486 1744 2487 1748
rect 2491 1744 2492 1748
rect 2486 1743 2492 1744
rect 2654 1748 2660 1749
rect 2654 1744 2655 1748
rect 2659 1744 2660 1748
rect 2654 1743 2660 1744
rect 2830 1748 2836 1749
rect 2830 1744 2831 1748
rect 2835 1744 2836 1748
rect 2830 1743 2836 1744
rect 3022 1748 3028 1749
rect 3022 1744 3023 1748
rect 3027 1744 3028 1748
rect 3022 1743 3028 1744
rect 3222 1748 3228 1749
rect 3222 1744 3223 1748
rect 3227 1744 3228 1748
rect 3222 1743 3228 1744
rect 3430 1748 3436 1749
rect 3430 1744 3431 1748
rect 3435 1744 3436 1748
rect 3430 1743 3436 1744
rect 3646 1748 3652 1749
rect 3646 1744 3647 1748
rect 3651 1744 3652 1748
rect 3646 1743 3652 1744
rect 3838 1748 3844 1749
rect 3838 1744 3839 1748
rect 3843 1744 3844 1748
rect 3942 1747 3943 1751
rect 3947 1747 3948 1751
rect 3942 1746 3948 1747
rect 3838 1743 3844 1744
rect 110 1732 116 1733
rect 2006 1732 2012 1733
rect 110 1728 111 1732
rect 115 1728 116 1732
rect 110 1727 116 1728
rect 366 1731 372 1732
rect 366 1727 367 1731
rect 371 1727 372 1731
rect 366 1726 372 1727
rect 494 1731 500 1732
rect 494 1727 495 1731
rect 499 1727 500 1731
rect 494 1726 500 1727
rect 638 1731 644 1732
rect 638 1727 639 1731
rect 643 1727 644 1731
rect 638 1726 644 1727
rect 798 1731 804 1732
rect 798 1727 799 1731
rect 803 1727 804 1731
rect 798 1726 804 1727
rect 966 1731 972 1732
rect 966 1727 967 1731
rect 971 1727 972 1731
rect 966 1726 972 1727
rect 1142 1731 1148 1732
rect 1142 1727 1143 1731
rect 1147 1727 1148 1731
rect 1142 1726 1148 1727
rect 1326 1731 1332 1732
rect 1326 1727 1327 1731
rect 1331 1727 1332 1731
rect 1326 1726 1332 1727
rect 1510 1731 1516 1732
rect 1510 1727 1511 1731
rect 1515 1727 1516 1731
rect 1510 1726 1516 1727
rect 1702 1731 1708 1732
rect 1702 1727 1703 1731
rect 1707 1727 1708 1731
rect 2006 1728 2007 1732
rect 2011 1728 2012 1732
rect 2006 1727 2012 1728
rect 1702 1726 1708 1727
rect 110 1715 116 1716
rect 110 1711 111 1715
rect 115 1711 116 1715
rect 2006 1715 2012 1716
rect 110 1710 116 1711
rect 366 1712 372 1713
rect 366 1708 367 1712
rect 371 1708 372 1712
rect 366 1707 372 1708
rect 494 1712 500 1713
rect 494 1708 495 1712
rect 499 1708 500 1712
rect 494 1707 500 1708
rect 638 1712 644 1713
rect 638 1708 639 1712
rect 643 1708 644 1712
rect 638 1707 644 1708
rect 798 1712 804 1713
rect 798 1708 799 1712
rect 803 1708 804 1712
rect 798 1707 804 1708
rect 966 1712 972 1713
rect 966 1708 967 1712
rect 971 1708 972 1712
rect 966 1707 972 1708
rect 1142 1712 1148 1713
rect 1142 1708 1143 1712
rect 1147 1708 1148 1712
rect 1142 1707 1148 1708
rect 1326 1712 1332 1713
rect 1326 1708 1327 1712
rect 1331 1708 1332 1712
rect 1326 1707 1332 1708
rect 1510 1712 1516 1713
rect 1510 1708 1511 1712
rect 1515 1708 1516 1712
rect 1510 1707 1516 1708
rect 1702 1712 1708 1713
rect 1702 1708 1703 1712
rect 1707 1708 1708 1712
rect 2006 1711 2007 1715
rect 2011 1711 2012 1715
rect 2006 1710 2012 1711
rect 1702 1707 1708 1708
rect 2222 1680 2228 1681
rect 2046 1677 2052 1678
rect 2046 1673 2047 1677
rect 2051 1673 2052 1677
rect 2222 1676 2223 1680
rect 2227 1676 2228 1680
rect 2222 1675 2228 1676
rect 2326 1680 2332 1681
rect 2326 1676 2327 1680
rect 2331 1676 2332 1680
rect 2326 1675 2332 1676
rect 2438 1680 2444 1681
rect 2438 1676 2439 1680
rect 2443 1676 2444 1680
rect 2438 1675 2444 1676
rect 2558 1680 2564 1681
rect 2558 1676 2559 1680
rect 2563 1676 2564 1680
rect 2558 1675 2564 1676
rect 2686 1680 2692 1681
rect 2686 1676 2687 1680
rect 2691 1676 2692 1680
rect 2686 1675 2692 1676
rect 2822 1680 2828 1681
rect 2822 1676 2823 1680
rect 2827 1676 2828 1680
rect 2822 1675 2828 1676
rect 2966 1680 2972 1681
rect 2966 1676 2967 1680
rect 2971 1676 2972 1680
rect 2966 1675 2972 1676
rect 3126 1680 3132 1681
rect 3126 1676 3127 1680
rect 3131 1676 3132 1680
rect 3126 1675 3132 1676
rect 3302 1680 3308 1681
rect 3302 1676 3303 1680
rect 3307 1676 3308 1680
rect 3302 1675 3308 1676
rect 3486 1680 3492 1681
rect 3486 1676 3487 1680
rect 3491 1676 3492 1680
rect 3486 1675 3492 1676
rect 3670 1680 3676 1681
rect 3670 1676 3671 1680
rect 3675 1676 3676 1680
rect 3670 1675 3676 1676
rect 3838 1680 3844 1681
rect 3838 1676 3839 1680
rect 3843 1676 3844 1680
rect 3838 1675 3844 1676
rect 3942 1677 3948 1678
rect 2046 1672 2052 1673
rect 3942 1673 3943 1677
rect 3947 1673 3948 1677
rect 3942 1672 3948 1673
rect 2222 1661 2228 1662
rect 2046 1660 2052 1661
rect 2046 1656 2047 1660
rect 2051 1656 2052 1660
rect 2222 1657 2223 1661
rect 2227 1657 2228 1661
rect 2222 1656 2228 1657
rect 2326 1661 2332 1662
rect 2326 1657 2327 1661
rect 2331 1657 2332 1661
rect 2326 1656 2332 1657
rect 2438 1661 2444 1662
rect 2438 1657 2439 1661
rect 2443 1657 2444 1661
rect 2438 1656 2444 1657
rect 2558 1661 2564 1662
rect 2558 1657 2559 1661
rect 2563 1657 2564 1661
rect 2558 1656 2564 1657
rect 2686 1661 2692 1662
rect 2686 1657 2687 1661
rect 2691 1657 2692 1661
rect 2686 1656 2692 1657
rect 2822 1661 2828 1662
rect 2822 1657 2823 1661
rect 2827 1657 2828 1661
rect 2822 1656 2828 1657
rect 2966 1661 2972 1662
rect 2966 1657 2967 1661
rect 2971 1657 2972 1661
rect 2966 1656 2972 1657
rect 3126 1661 3132 1662
rect 3126 1657 3127 1661
rect 3131 1657 3132 1661
rect 3126 1656 3132 1657
rect 3302 1661 3308 1662
rect 3302 1657 3303 1661
rect 3307 1657 3308 1661
rect 3302 1656 3308 1657
rect 3486 1661 3492 1662
rect 3486 1657 3487 1661
rect 3491 1657 3492 1661
rect 3486 1656 3492 1657
rect 3670 1661 3676 1662
rect 3670 1657 3671 1661
rect 3675 1657 3676 1661
rect 3670 1656 3676 1657
rect 3838 1661 3844 1662
rect 3838 1657 3839 1661
rect 3843 1657 3844 1661
rect 3838 1656 3844 1657
rect 3942 1660 3948 1661
rect 3942 1656 3943 1660
rect 3947 1656 3948 1660
rect 2046 1655 2052 1656
rect 3942 1655 3948 1656
rect 134 1648 140 1649
rect 110 1645 116 1646
rect 110 1641 111 1645
rect 115 1641 116 1645
rect 134 1644 135 1648
rect 139 1644 140 1648
rect 134 1643 140 1644
rect 246 1648 252 1649
rect 246 1644 247 1648
rect 251 1644 252 1648
rect 246 1643 252 1644
rect 398 1648 404 1649
rect 398 1644 399 1648
rect 403 1644 404 1648
rect 398 1643 404 1644
rect 566 1648 572 1649
rect 566 1644 567 1648
rect 571 1644 572 1648
rect 566 1643 572 1644
rect 742 1648 748 1649
rect 742 1644 743 1648
rect 747 1644 748 1648
rect 742 1643 748 1644
rect 934 1648 940 1649
rect 934 1644 935 1648
rect 939 1644 940 1648
rect 934 1643 940 1644
rect 1134 1648 1140 1649
rect 1134 1644 1135 1648
rect 1139 1644 1140 1648
rect 1134 1643 1140 1644
rect 1342 1648 1348 1649
rect 1342 1644 1343 1648
rect 1347 1644 1348 1648
rect 1342 1643 1348 1644
rect 1550 1648 1556 1649
rect 1550 1644 1551 1648
rect 1555 1644 1556 1648
rect 1550 1643 1556 1644
rect 1766 1648 1772 1649
rect 1766 1644 1767 1648
rect 1771 1644 1772 1648
rect 1766 1643 1772 1644
rect 2006 1645 2012 1646
rect 110 1640 116 1641
rect 2006 1641 2007 1645
rect 2011 1641 2012 1645
rect 2006 1640 2012 1641
rect 134 1629 140 1630
rect 110 1628 116 1629
rect 110 1624 111 1628
rect 115 1624 116 1628
rect 134 1625 135 1629
rect 139 1625 140 1629
rect 134 1624 140 1625
rect 246 1629 252 1630
rect 246 1625 247 1629
rect 251 1625 252 1629
rect 246 1624 252 1625
rect 398 1629 404 1630
rect 398 1625 399 1629
rect 403 1625 404 1629
rect 398 1624 404 1625
rect 566 1629 572 1630
rect 566 1625 567 1629
rect 571 1625 572 1629
rect 566 1624 572 1625
rect 742 1629 748 1630
rect 742 1625 743 1629
rect 747 1625 748 1629
rect 742 1624 748 1625
rect 934 1629 940 1630
rect 934 1625 935 1629
rect 939 1625 940 1629
rect 934 1624 940 1625
rect 1134 1629 1140 1630
rect 1134 1625 1135 1629
rect 1139 1625 1140 1629
rect 1134 1624 1140 1625
rect 1342 1629 1348 1630
rect 1342 1625 1343 1629
rect 1347 1625 1348 1629
rect 1342 1624 1348 1625
rect 1550 1629 1556 1630
rect 1550 1625 1551 1629
rect 1555 1625 1556 1629
rect 1550 1624 1556 1625
rect 1766 1629 1772 1630
rect 1766 1625 1767 1629
rect 1771 1625 1772 1629
rect 1766 1624 1772 1625
rect 2006 1628 2012 1629
rect 2006 1624 2007 1628
rect 2011 1624 2012 1628
rect 110 1623 116 1624
rect 2006 1623 2012 1624
rect 2046 1604 2052 1605
rect 3942 1604 3948 1605
rect 2046 1600 2047 1604
rect 2051 1600 2052 1604
rect 2046 1599 2052 1600
rect 2390 1603 2396 1604
rect 2390 1599 2391 1603
rect 2395 1599 2396 1603
rect 2390 1598 2396 1599
rect 2502 1603 2508 1604
rect 2502 1599 2503 1603
rect 2507 1599 2508 1603
rect 2502 1598 2508 1599
rect 2614 1603 2620 1604
rect 2614 1599 2615 1603
rect 2619 1599 2620 1603
rect 2614 1598 2620 1599
rect 2734 1603 2740 1604
rect 2734 1599 2735 1603
rect 2739 1599 2740 1603
rect 2734 1598 2740 1599
rect 2854 1603 2860 1604
rect 2854 1599 2855 1603
rect 2859 1599 2860 1603
rect 2854 1598 2860 1599
rect 2974 1603 2980 1604
rect 2974 1599 2975 1603
rect 2979 1599 2980 1603
rect 2974 1598 2980 1599
rect 3094 1603 3100 1604
rect 3094 1599 3095 1603
rect 3099 1599 3100 1603
rect 3094 1598 3100 1599
rect 3214 1603 3220 1604
rect 3214 1599 3215 1603
rect 3219 1599 3220 1603
rect 3214 1598 3220 1599
rect 3334 1603 3340 1604
rect 3334 1599 3335 1603
rect 3339 1599 3340 1603
rect 3334 1598 3340 1599
rect 3454 1603 3460 1604
rect 3454 1599 3455 1603
rect 3459 1599 3460 1603
rect 3942 1600 3943 1604
rect 3947 1600 3948 1604
rect 3942 1599 3948 1600
rect 3454 1598 3460 1599
rect 2046 1587 2052 1588
rect 2046 1583 2047 1587
rect 2051 1583 2052 1587
rect 3942 1587 3948 1588
rect 2046 1582 2052 1583
rect 2390 1584 2396 1585
rect 2390 1580 2391 1584
rect 2395 1580 2396 1584
rect 2390 1579 2396 1580
rect 2502 1584 2508 1585
rect 2502 1580 2503 1584
rect 2507 1580 2508 1584
rect 2502 1579 2508 1580
rect 2614 1584 2620 1585
rect 2614 1580 2615 1584
rect 2619 1580 2620 1584
rect 2614 1579 2620 1580
rect 2734 1584 2740 1585
rect 2734 1580 2735 1584
rect 2739 1580 2740 1584
rect 2734 1579 2740 1580
rect 2854 1584 2860 1585
rect 2854 1580 2855 1584
rect 2859 1580 2860 1584
rect 2854 1579 2860 1580
rect 2974 1584 2980 1585
rect 2974 1580 2975 1584
rect 2979 1580 2980 1584
rect 2974 1579 2980 1580
rect 3094 1584 3100 1585
rect 3094 1580 3095 1584
rect 3099 1580 3100 1584
rect 3094 1579 3100 1580
rect 3214 1584 3220 1585
rect 3214 1580 3215 1584
rect 3219 1580 3220 1584
rect 3214 1579 3220 1580
rect 3334 1584 3340 1585
rect 3334 1580 3335 1584
rect 3339 1580 3340 1584
rect 3334 1579 3340 1580
rect 3454 1584 3460 1585
rect 3454 1580 3455 1584
rect 3459 1580 3460 1584
rect 3942 1583 3943 1587
rect 3947 1583 3948 1587
rect 3942 1582 3948 1583
rect 3454 1579 3460 1580
rect 110 1572 116 1573
rect 2006 1572 2012 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 110 1567 116 1568
rect 134 1571 140 1572
rect 134 1567 135 1571
rect 139 1567 140 1571
rect 134 1566 140 1567
rect 254 1571 260 1572
rect 254 1567 255 1571
rect 259 1567 260 1571
rect 254 1566 260 1567
rect 422 1571 428 1572
rect 422 1567 423 1571
rect 427 1567 428 1571
rect 422 1566 428 1567
rect 614 1571 620 1572
rect 614 1567 615 1571
rect 619 1567 620 1571
rect 614 1566 620 1567
rect 830 1571 836 1572
rect 830 1567 831 1571
rect 835 1567 836 1571
rect 830 1566 836 1567
rect 1062 1571 1068 1572
rect 1062 1567 1063 1571
rect 1067 1567 1068 1571
rect 1062 1566 1068 1567
rect 1310 1571 1316 1572
rect 1310 1567 1311 1571
rect 1315 1567 1316 1571
rect 1310 1566 1316 1567
rect 1566 1571 1572 1572
rect 1566 1567 1567 1571
rect 1571 1567 1572 1571
rect 1566 1566 1572 1567
rect 1830 1571 1836 1572
rect 1830 1567 1831 1571
rect 1835 1567 1836 1571
rect 2006 1568 2007 1572
rect 2011 1568 2012 1572
rect 2006 1567 2012 1568
rect 1830 1566 1836 1567
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 2006 1555 2012 1556
rect 110 1550 116 1551
rect 134 1552 140 1553
rect 134 1548 135 1552
rect 139 1548 140 1552
rect 134 1547 140 1548
rect 254 1552 260 1553
rect 254 1548 255 1552
rect 259 1548 260 1552
rect 254 1547 260 1548
rect 422 1552 428 1553
rect 422 1548 423 1552
rect 427 1548 428 1552
rect 422 1547 428 1548
rect 614 1552 620 1553
rect 614 1548 615 1552
rect 619 1548 620 1552
rect 614 1547 620 1548
rect 830 1552 836 1553
rect 830 1548 831 1552
rect 835 1548 836 1552
rect 830 1547 836 1548
rect 1062 1552 1068 1553
rect 1062 1548 1063 1552
rect 1067 1548 1068 1552
rect 1062 1547 1068 1548
rect 1310 1552 1316 1553
rect 1310 1548 1311 1552
rect 1315 1548 1316 1552
rect 1310 1547 1316 1548
rect 1566 1552 1572 1553
rect 1566 1548 1567 1552
rect 1571 1548 1572 1552
rect 1566 1547 1572 1548
rect 1830 1552 1836 1553
rect 1830 1548 1831 1552
rect 1835 1548 1836 1552
rect 2006 1551 2007 1555
rect 2011 1551 2012 1555
rect 2006 1550 2012 1551
rect 1830 1547 1836 1548
rect 2542 1524 2548 1525
rect 2046 1521 2052 1522
rect 2046 1517 2047 1521
rect 2051 1517 2052 1521
rect 2542 1520 2543 1524
rect 2547 1520 2548 1524
rect 2542 1519 2548 1520
rect 2670 1524 2676 1525
rect 2670 1520 2671 1524
rect 2675 1520 2676 1524
rect 2670 1519 2676 1520
rect 2798 1524 2804 1525
rect 2798 1520 2799 1524
rect 2803 1520 2804 1524
rect 2798 1519 2804 1520
rect 2934 1524 2940 1525
rect 2934 1520 2935 1524
rect 2939 1520 2940 1524
rect 2934 1519 2940 1520
rect 3070 1524 3076 1525
rect 3070 1520 3071 1524
rect 3075 1520 3076 1524
rect 3070 1519 3076 1520
rect 3206 1524 3212 1525
rect 3206 1520 3207 1524
rect 3211 1520 3212 1524
rect 3206 1519 3212 1520
rect 3334 1524 3340 1525
rect 3334 1520 3335 1524
rect 3339 1520 3340 1524
rect 3334 1519 3340 1520
rect 3462 1524 3468 1525
rect 3462 1520 3463 1524
rect 3467 1520 3468 1524
rect 3462 1519 3468 1520
rect 3590 1524 3596 1525
rect 3590 1520 3591 1524
rect 3595 1520 3596 1524
rect 3590 1519 3596 1520
rect 3726 1524 3732 1525
rect 3726 1520 3727 1524
rect 3731 1520 3732 1524
rect 3726 1519 3732 1520
rect 3838 1524 3844 1525
rect 3838 1520 3839 1524
rect 3843 1520 3844 1524
rect 3838 1519 3844 1520
rect 3942 1521 3948 1522
rect 2046 1516 2052 1517
rect 3942 1517 3943 1521
rect 3947 1517 3948 1521
rect 3942 1516 3948 1517
rect 2542 1505 2548 1506
rect 2046 1504 2052 1505
rect 2046 1500 2047 1504
rect 2051 1500 2052 1504
rect 2542 1501 2543 1505
rect 2547 1501 2548 1505
rect 2542 1500 2548 1501
rect 2670 1505 2676 1506
rect 2670 1501 2671 1505
rect 2675 1501 2676 1505
rect 2670 1500 2676 1501
rect 2798 1505 2804 1506
rect 2798 1501 2799 1505
rect 2803 1501 2804 1505
rect 2798 1500 2804 1501
rect 2934 1505 2940 1506
rect 2934 1501 2935 1505
rect 2939 1501 2940 1505
rect 2934 1500 2940 1501
rect 3070 1505 3076 1506
rect 3070 1501 3071 1505
rect 3075 1501 3076 1505
rect 3070 1500 3076 1501
rect 3206 1505 3212 1506
rect 3206 1501 3207 1505
rect 3211 1501 3212 1505
rect 3206 1500 3212 1501
rect 3334 1505 3340 1506
rect 3334 1501 3335 1505
rect 3339 1501 3340 1505
rect 3334 1500 3340 1501
rect 3462 1505 3468 1506
rect 3462 1501 3463 1505
rect 3467 1501 3468 1505
rect 3462 1500 3468 1501
rect 3590 1505 3596 1506
rect 3590 1501 3591 1505
rect 3595 1501 3596 1505
rect 3590 1500 3596 1501
rect 3726 1505 3732 1506
rect 3726 1501 3727 1505
rect 3731 1501 3732 1505
rect 3726 1500 3732 1501
rect 3838 1505 3844 1506
rect 3838 1501 3839 1505
rect 3843 1501 3844 1505
rect 3838 1500 3844 1501
rect 3942 1504 3948 1505
rect 3942 1500 3943 1504
rect 3947 1500 3948 1504
rect 2046 1499 2052 1500
rect 3942 1499 3948 1500
rect 238 1488 244 1489
rect 110 1485 116 1486
rect 110 1481 111 1485
rect 115 1481 116 1485
rect 238 1484 239 1488
rect 243 1484 244 1488
rect 238 1483 244 1484
rect 406 1488 412 1489
rect 406 1484 407 1488
rect 411 1484 412 1488
rect 406 1483 412 1484
rect 582 1488 588 1489
rect 582 1484 583 1488
rect 587 1484 588 1488
rect 582 1483 588 1484
rect 774 1488 780 1489
rect 774 1484 775 1488
rect 779 1484 780 1488
rect 774 1483 780 1484
rect 966 1488 972 1489
rect 966 1484 967 1488
rect 971 1484 972 1488
rect 966 1483 972 1484
rect 1158 1488 1164 1489
rect 1158 1484 1159 1488
rect 1163 1484 1164 1488
rect 1158 1483 1164 1484
rect 1350 1488 1356 1489
rect 1350 1484 1351 1488
rect 1355 1484 1356 1488
rect 1350 1483 1356 1484
rect 1542 1488 1548 1489
rect 1542 1484 1543 1488
rect 1547 1484 1548 1488
rect 1542 1483 1548 1484
rect 1734 1488 1740 1489
rect 1734 1484 1735 1488
rect 1739 1484 1740 1488
rect 1734 1483 1740 1484
rect 1902 1488 1908 1489
rect 1902 1484 1903 1488
rect 1907 1484 1908 1488
rect 1902 1483 1908 1484
rect 2006 1485 2012 1486
rect 110 1480 116 1481
rect 2006 1481 2007 1485
rect 2011 1481 2012 1485
rect 2006 1480 2012 1481
rect 238 1469 244 1470
rect 110 1468 116 1469
rect 110 1464 111 1468
rect 115 1464 116 1468
rect 238 1465 239 1469
rect 243 1465 244 1469
rect 238 1464 244 1465
rect 406 1469 412 1470
rect 406 1465 407 1469
rect 411 1465 412 1469
rect 406 1464 412 1465
rect 582 1469 588 1470
rect 582 1465 583 1469
rect 587 1465 588 1469
rect 582 1464 588 1465
rect 774 1469 780 1470
rect 774 1465 775 1469
rect 779 1465 780 1469
rect 774 1464 780 1465
rect 966 1469 972 1470
rect 966 1465 967 1469
rect 971 1465 972 1469
rect 966 1464 972 1465
rect 1158 1469 1164 1470
rect 1158 1465 1159 1469
rect 1163 1465 1164 1469
rect 1158 1464 1164 1465
rect 1350 1469 1356 1470
rect 1350 1465 1351 1469
rect 1355 1465 1356 1469
rect 1350 1464 1356 1465
rect 1542 1469 1548 1470
rect 1542 1465 1543 1469
rect 1547 1465 1548 1469
rect 1542 1464 1548 1465
rect 1734 1469 1740 1470
rect 1734 1465 1735 1469
rect 1739 1465 1740 1469
rect 1734 1464 1740 1465
rect 1902 1469 1908 1470
rect 1902 1465 1903 1469
rect 1907 1465 1908 1469
rect 1902 1464 1908 1465
rect 2006 1468 2012 1469
rect 2006 1464 2007 1468
rect 2011 1464 2012 1468
rect 110 1463 116 1464
rect 2006 1463 2012 1464
rect 2046 1440 2052 1441
rect 3942 1440 3948 1441
rect 2046 1436 2047 1440
rect 2051 1436 2052 1440
rect 2046 1435 2052 1436
rect 2518 1439 2524 1440
rect 2518 1435 2519 1439
rect 2523 1435 2524 1439
rect 2518 1434 2524 1435
rect 2630 1439 2636 1440
rect 2630 1435 2631 1439
rect 2635 1435 2636 1439
rect 2630 1434 2636 1435
rect 2758 1439 2764 1440
rect 2758 1435 2759 1439
rect 2763 1435 2764 1439
rect 2758 1434 2764 1435
rect 2894 1439 2900 1440
rect 2894 1435 2895 1439
rect 2899 1435 2900 1439
rect 2894 1434 2900 1435
rect 3030 1439 3036 1440
rect 3030 1435 3031 1439
rect 3035 1435 3036 1439
rect 3030 1434 3036 1435
rect 3174 1439 3180 1440
rect 3174 1435 3175 1439
rect 3179 1435 3180 1439
rect 3174 1434 3180 1435
rect 3310 1439 3316 1440
rect 3310 1435 3311 1439
rect 3315 1435 3316 1439
rect 3310 1434 3316 1435
rect 3446 1439 3452 1440
rect 3446 1435 3447 1439
rect 3451 1435 3452 1439
rect 3446 1434 3452 1435
rect 3582 1439 3588 1440
rect 3582 1435 3583 1439
rect 3587 1435 3588 1439
rect 3582 1434 3588 1435
rect 3718 1439 3724 1440
rect 3718 1435 3719 1439
rect 3723 1435 3724 1439
rect 3718 1434 3724 1435
rect 3838 1439 3844 1440
rect 3838 1435 3839 1439
rect 3843 1435 3844 1439
rect 3942 1436 3943 1440
rect 3947 1436 3948 1440
rect 3942 1435 3948 1436
rect 3838 1434 3844 1435
rect 2046 1423 2052 1424
rect 2046 1419 2047 1423
rect 2051 1419 2052 1423
rect 3942 1423 3948 1424
rect 2046 1418 2052 1419
rect 2518 1420 2524 1421
rect 2518 1416 2519 1420
rect 2523 1416 2524 1420
rect 2518 1415 2524 1416
rect 2630 1420 2636 1421
rect 2630 1416 2631 1420
rect 2635 1416 2636 1420
rect 2630 1415 2636 1416
rect 2758 1420 2764 1421
rect 2758 1416 2759 1420
rect 2763 1416 2764 1420
rect 2758 1415 2764 1416
rect 2894 1420 2900 1421
rect 2894 1416 2895 1420
rect 2899 1416 2900 1420
rect 2894 1415 2900 1416
rect 3030 1420 3036 1421
rect 3030 1416 3031 1420
rect 3035 1416 3036 1420
rect 3030 1415 3036 1416
rect 3174 1420 3180 1421
rect 3174 1416 3175 1420
rect 3179 1416 3180 1420
rect 3174 1415 3180 1416
rect 3310 1420 3316 1421
rect 3310 1416 3311 1420
rect 3315 1416 3316 1420
rect 3310 1415 3316 1416
rect 3446 1420 3452 1421
rect 3446 1416 3447 1420
rect 3451 1416 3452 1420
rect 3446 1415 3452 1416
rect 3582 1420 3588 1421
rect 3582 1416 3583 1420
rect 3587 1416 3588 1420
rect 3582 1415 3588 1416
rect 3718 1420 3724 1421
rect 3718 1416 3719 1420
rect 3723 1416 3724 1420
rect 3718 1415 3724 1416
rect 3838 1420 3844 1421
rect 3838 1416 3839 1420
rect 3843 1416 3844 1420
rect 3942 1419 3943 1423
rect 3947 1419 3948 1423
rect 3942 1418 3948 1419
rect 3838 1415 3844 1416
rect 110 1408 116 1409
rect 2006 1408 2012 1409
rect 110 1404 111 1408
rect 115 1404 116 1408
rect 110 1403 116 1404
rect 462 1407 468 1408
rect 462 1403 463 1407
rect 467 1403 468 1407
rect 462 1402 468 1403
rect 582 1407 588 1408
rect 582 1403 583 1407
rect 587 1403 588 1407
rect 582 1402 588 1403
rect 710 1407 716 1408
rect 710 1403 711 1407
rect 715 1403 716 1407
rect 710 1402 716 1403
rect 854 1407 860 1408
rect 854 1403 855 1407
rect 859 1403 860 1407
rect 854 1402 860 1403
rect 1006 1407 1012 1408
rect 1006 1403 1007 1407
rect 1011 1403 1012 1407
rect 1006 1402 1012 1403
rect 1166 1407 1172 1408
rect 1166 1403 1167 1407
rect 1171 1403 1172 1407
rect 1166 1402 1172 1403
rect 1334 1407 1340 1408
rect 1334 1403 1335 1407
rect 1339 1403 1340 1407
rect 1334 1402 1340 1403
rect 1510 1407 1516 1408
rect 1510 1403 1511 1407
rect 1515 1403 1516 1407
rect 1510 1402 1516 1403
rect 1686 1407 1692 1408
rect 1686 1403 1687 1407
rect 1691 1403 1692 1407
rect 1686 1402 1692 1403
rect 1870 1407 1876 1408
rect 1870 1403 1871 1407
rect 1875 1403 1876 1407
rect 2006 1404 2007 1408
rect 2011 1404 2012 1408
rect 2006 1403 2012 1404
rect 1870 1402 1876 1403
rect 110 1391 116 1392
rect 110 1387 111 1391
rect 115 1387 116 1391
rect 2006 1391 2012 1392
rect 110 1386 116 1387
rect 462 1388 468 1389
rect 462 1384 463 1388
rect 467 1384 468 1388
rect 462 1383 468 1384
rect 582 1388 588 1389
rect 582 1384 583 1388
rect 587 1384 588 1388
rect 582 1383 588 1384
rect 710 1388 716 1389
rect 710 1384 711 1388
rect 715 1384 716 1388
rect 710 1383 716 1384
rect 854 1388 860 1389
rect 854 1384 855 1388
rect 859 1384 860 1388
rect 854 1383 860 1384
rect 1006 1388 1012 1389
rect 1006 1384 1007 1388
rect 1011 1384 1012 1388
rect 1006 1383 1012 1384
rect 1166 1388 1172 1389
rect 1166 1384 1167 1388
rect 1171 1384 1172 1388
rect 1166 1383 1172 1384
rect 1334 1388 1340 1389
rect 1334 1384 1335 1388
rect 1339 1384 1340 1388
rect 1334 1383 1340 1384
rect 1510 1388 1516 1389
rect 1510 1384 1511 1388
rect 1515 1384 1516 1388
rect 1510 1383 1516 1384
rect 1686 1388 1692 1389
rect 1686 1384 1687 1388
rect 1691 1384 1692 1388
rect 1686 1383 1692 1384
rect 1870 1388 1876 1389
rect 1870 1384 1871 1388
rect 1875 1384 1876 1388
rect 2006 1387 2007 1391
rect 2011 1387 2012 1391
rect 2006 1386 2012 1387
rect 1870 1383 1876 1384
rect 2398 1360 2404 1361
rect 2046 1357 2052 1358
rect 2046 1353 2047 1357
rect 2051 1353 2052 1357
rect 2398 1356 2399 1360
rect 2403 1356 2404 1360
rect 2398 1355 2404 1356
rect 2534 1360 2540 1361
rect 2534 1356 2535 1360
rect 2539 1356 2540 1360
rect 2534 1355 2540 1356
rect 2678 1360 2684 1361
rect 2678 1356 2679 1360
rect 2683 1356 2684 1360
rect 2678 1355 2684 1356
rect 2822 1360 2828 1361
rect 2822 1356 2823 1360
rect 2827 1356 2828 1360
rect 2822 1355 2828 1356
rect 2966 1360 2972 1361
rect 2966 1356 2967 1360
rect 2971 1356 2972 1360
rect 2966 1355 2972 1356
rect 3110 1360 3116 1361
rect 3110 1356 3111 1360
rect 3115 1356 3116 1360
rect 3110 1355 3116 1356
rect 3254 1360 3260 1361
rect 3254 1356 3255 1360
rect 3259 1356 3260 1360
rect 3254 1355 3260 1356
rect 3406 1360 3412 1361
rect 3406 1356 3407 1360
rect 3411 1356 3412 1360
rect 3406 1355 3412 1356
rect 3558 1360 3564 1361
rect 3558 1356 3559 1360
rect 3563 1356 3564 1360
rect 3558 1355 3564 1356
rect 3710 1360 3716 1361
rect 3710 1356 3711 1360
rect 3715 1356 3716 1360
rect 3710 1355 3716 1356
rect 3838 1360 3844 1361
rect 3838 1356 3839 1360
rect 3843 1356 3844 1360
rect 3838 1355 3844 1356
rect 3942 1357 3948 1358
rect 2046 1352 2052 1353
rect 3942 1353 3943 1357
rect 3947 1353 3948 1357
rect 3942 1352 3948 1353
rect 2398 1341 2404 1342
rect 2046 1340 2052 1341
rect 2046 1336 2047 1340
rect 2051 1336 2052 1340
rect 2398 1337 2399 1341
rect 2403 1337 2404 1341
rect 2398 1336 2404 1337
rect 2534 1341 2540 1342
rect 2534 1337 2535 1341
rect 2539 1337 2540 1341
rect 2534 1336 2540 1337
rect 2678 1341 2684 1342
rect 2678 1337 2679 1341
rect 2683 1337 2684 1341
rect 2678 1336 2684 1337
rect 2822 1341 2828 1342
rect 2822 1337 2823 1341
rect 2827 1337 2828 1341
rect 2822 1336 2828 1337
rect 2966 1341 2972 1342
rect 2966 1337 2967 1341
rect 2971 1337 2972 1341
rect 2966 1336 2972 1337
rect 3110 1341 3116 1342
rect 3110 1337 3111 1341
rect 3115 1337 3116 1341
rect 3110 1336 3116 1337
rect 3254 1341 3260 1342
rect 3254 1337 3255 1341
rect 3259 1337 3260 1341
rect 3254 1336 3260 1337
rect 3406 1341 3412 1342
rect 3406 1337 3407 1341
rect 3411 1337 3412 1341
rect 3406 1336 3412 1337
rect 3558 1341 3564 1342
rect 3558 1337 3559 1341
rect 3563 1337 3564 1341
rect 3558 1336 3564 1337
rect 3710 1341 3716 1342
rect 3710 1337 3711 1341
rect 3715 1337 3716 1341
rect 3710 1336 3716 1337
rect 3838 1341 3844 1342
rect 3838 1337 3839 1341
rect 3843 1337 3844 1341
rect 3838 1336 3844 1337
rect 3942 1340 3948 1341
rect 3942 1336 3943 1340
rect 3947 1336 3948 1340
rect 2046 1335 2052 1336
rect 3942 1335 3948 1336
rect 654 1328 660 1329
rect 110 1325 116 1326
rect 110 1321 111 1325
rect 115 1321 116 1325
rect 654 1324 655 1328
rect 659 1324 660 1328
rect 654 1323 660 1324
rect 766 1328 772 1329
rect 766 1324 767 1328
rect 771 1324 772 1328
rect 766 1323 772 1324
rect 886 1328 892 1329
rect 886 1324 887 1328
rect 891 1324 892 1328
rect 886 1323 892 1324
rect 1014 1328 1020 1329
rect 1014 1324 1015 1328
rect 1019 1324 1020 1328
rect 1014 1323 1020 1324
rect 1142 1328 1148 1329
rect 1142 1324 1143 1328
rect 1147 1324 1148 1328
rect 1142 1323 1148 1324
rect 1278 1328 1284 1329
rect 1278 1324 1279 1328
rect 1283 1324 1284 1328
rect 1278 1323 1284 1324
rect 1414 1328 1420 1329
rect 1414 1324 1415 1328
rect 1419 1324 1420 1328
rect 1414 1323 1420 1324
rect 1558 1328 1564 1329
rect 1558 1324 1559 1328
rect 1563 1324 1564 1328
rect 1558 1323 1564 1324
rect 1702 1328 1708 1329
rect 1702 1324 1703 1328
rect 1707 1324 1708 1328
rect 1702 1323 1708 1324
rect 1846 1328 1852 1329
rect 1846 1324 1847 1328
rect 1851 1324 1852 1328
rect 1846 1323 1852 1324
rect 2006 1325 2012 1326
rect 110 1320 116 1321
rect 2006 1321 2007 1325
rect 2011 1321 2012 1325
rect 2006 1320 2012 1321
rect 654 1309 660 1310
rect 110 1308 116 1309
rect 110 1304 111 1308
rect 115 1304 116 1308
rect 654 1305 655 1309
rect 659 1305 660 1309
rect 654 1304 660 1305
rect 766 1309 772 1310
rect 766 1305 767 1309
rect 771 1305 772 1309
rect 766 1304 772 1305
rect 886 1309 892 1310
rect 886 1305 887 1309
rect 891 1305 892 1309
rect 886 1304 892 1305
rect 1014 1309 1020 1310
rect 1014 1305 1015 1309
rect 1019 1305 1020 1309
rect 1014 1304 1020 1305
rect 1142 1309 1148 1310
rect 1142 1305 1143 1309
rect 1147 1305 1148 1309
rect 1142 1304 1148 1305
rect 1278 1309 1284 1310
rect 1278 1305 1279 1309
rect 1283 1305 1284 1309
rect 1278 1304 1284 1305
rect 1414 1309 1420 1310
rect 1414 1305 1415 1309
rect 1419 1305 1420 1309
rect 1414 1304 1420 1305
rect 1558 1309 1564 1310
rect 1558 1305 1559 1309
rect 1563 1305 1564 1309
rect 1558 1304 1564 1305
rect 1702 1309 1708 1310
rect 1702 1305 1703 1309
rect 1707 1305 1708 1309
rect 1702 1304 1708 1305
rect 1846 1309 1852 1310
rect 1846 1305 1847 1309
rect 1851 1305 1852 1309
rect 1846 1304 1852 1305
rect 2006 1308 2012 1309
rect 2006 1304 2007 1308
rect 2011 1304 2012 1308
rect 110 1303 116 1304
rect 2006 1303 2012 1304
rect 2046 1284 2052 1285
rect 3942 1284 3948 1285
rect 2046 1280 2047 1284
rect 2051 1280 2052 1284
rect 2046 1279 2052 1280
rect 2246 1283 2252 1284
rect 2246 1279 2247 1283
rect 2251 1279 2252 1283
rect 2246 1278 2252 1279
rect 2374 1283 2380 1284
rect 2374 1279 2375 1283
rect 2379 1279 2380 1283
rect 2374 1278 2380 1279
rect 2510 1283 2516 1284
rect 2510 1279 2511 1283
rect 2515 1279 2516 1283
rect 2510 1278 2516 1279
rect 2646 1283 2652 1284
rect 2646 1279 2647 1283
rect 2651 1279 2652 1283
rect 2646 1278 2652 1279
rect 2790 1283 2796 1284
rect 2790 1279 2791 1283
rect 2795 1279 2796 1283
rect 2790 1278 2796 1279
rect 2942 1283 2948 1284
rect 2942 1279 2943 1283
rect 2947 1279 2948 1283
rect 2942 1278 2948 1279
rect 3110 1283 3116 1284
rect 3110 1279 3111 1283
rect 3115 1279 3116 1283
rect 3110 1278 3116 1279
rect 3286 1283 3292 1284
rect 3286 1279 3287 1283
rect 3291 1279 3292 1283
rect 3286 1278 3292 1279
rect 3470 1283 3476 1284
rect 3470 1279 3471 1283
rect 3475 1279 3476 1283
rect 3470 1278 3476 1279
rect 3662 1283 3668 1284
rect 3662 1279 3663 1283
rect 3667 1279 3668 1283
rect 3662 1278 3668 1279
rect 3838 1283 3844 1284
rect 3838 1279 3839 1283
rect 3843 1279 3844 1283
rect 3942 1280 3943 1284
rect 3947 1280 3948 1284
rect 3942 1279 3948 1280
rect 3838 1278 3844 1279
rect 2046 1267 2052 1268
rect 2046 1263 2047 1267
rect 2051 1263 2052 1267
rect 3942 1267 3948 1268
rect 2046 1262 2052 1263
rect 2246 1264 2252 1265
rect 2246 1260 2247 1264
rect 2251 1260 2252 1264
rect 2246 1259 2252 1260
rect 2374 1264 2380 1265
rect 2374 1260 2375 1264
rect 2379 1260 2380 1264
rect 2374 1259 2380 1260
rect 2510 1264 2516 1265
rect 2510 1260 2511 1264
rect 2515 1260 2516 1264
rect 2510 1259 2516 1260
rect 2646 1264 2652 1265
rect 2646 1260 2647 1264
rect 2651 1260 2652 1264
rect 2646 1259 2652 1260
rect 2790 1264 2796 1265
rect 2790 1260 2791 1264
rect 2795 1260 2796 1264
rect 2790 1259 2796 1260
rect 2942 1264 2948 1265
rect 2942 1260 2943 1264
rect 2947 1260 2948 1264
rect 2942 1259 2948 1260
rect 3110 1264 3116 1265
rect 3110 1260 3111 1264
rect 3115 1260 3116 1264
rect 3110 1259 3116 1260
rect 3286 1264 3292 1265
rect 3286 1260 3287 1264
rect 3291 1260 3292 1264
rect 3286 1259 3292 1260
rect 3470 1264 3476 1265
rect 3470 1260 3471 1264
rect 3475 1260 3476 1264
rect 3470 1259 3476 1260
rect 3662 1264 3668 1265
rect 3662 1260 3663 1264
rect 3667 1260 3668 1264
rect 3662 1259 3668 1260
rect 3838 1264 3844 1265
rect 3838 1260 3839 1264
rect 3843 1260 3844 1264
rect 3942 1263 3943 1267
rect 3947 1263 3948 1267
rect 3942 1262 3948 1263
rect 3838 1259 3844 1260
rect 110 1252 116 1253
rect 2006 1252 2012 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 438 1251 444 1252
rect 438 1247 439 1251
rect 443 1247 444 1251
rect 438 1246 444 1247
rect 550 1251 556 1252
rect 550 1247 551 1251
rect 555 1247 556 1251
rect 550 1246 556 1247
rect 670 1251 676 1252
rect 670 1247 671 1251
rect 675 1247 676 1251
rect 670 1246 676 1247
rect 798 1251 804 1252
rect 798 1247 799 1251
rect 803 1247 804 1251
rect 798 1246 804 1247
rect 934 1251 940 1252
rect 934 1247 935 1251
rect 939 1247 940 1251
rect 934 1246 940 1247
rect 1078 1251 1084 1252
rect 1078 1247 1079 1251
rect 1083 1247 1084 1251
rect 1078 1246 1084 1247
rect 1230 1251 1236 1252
rect 1230 1247 1231 1251
rect 1235 1247 1236 1251
rect 1230 1246 1236 1247
rect 1390 1251 1396 1252
rect 1390 1247 1391 1251
rect 1395 1247 1396 1251
rect 1390 1246 1396 1247
rect 1550 1251 1556 1252
rect 1550 1247 1551 1251
rect 1555 1247 1556 1251
rect 1550 1246 1556 1247
rect 1718 1251 1724 1252
rect 1718 1247 1719 1251
rect 1723 1247 1724 1251
rect 2006 1248 2007 1252
rect 2011 1248 2012 1252
rect 2006 1247 2012 1248
rect 1718 1246 1724 1247
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 2006 1235 2012 1236
rect 110 1230 116 1231
rect 438 1232 444 1233
rect 438 1228 439 1232
rect 443 1228 444 1232
rect 438 1227 444 1228
rect 550 1232 556 1233
rect 550 1228 551 1232
rect 555 1228 556 1232
rect 550 1227 556 1228
rect 670 1232 676 1233
rect 670 1228 671 1232
rect 675 1228 676 1232
rect 670 1227 676 1228
rect 798 1232 804 1233
rect 798 1228 799 1232
rect 803 1228 804 1232
rect 798 1227 804 1228
rect 934 1232 940 1233
rect 934 1228 935 1232
rect 939 1228 940 1232
rect 934 1227 940 1228
rect 1078 1232 1084 1233
rect 1078 1228 1079 1232
rect 1083 1228 1084 1232
rect 1078 1227 1084 1228
rect 1230 1232 1236 1233
rect 1230 1228 1231 1232
rect 1235 1228 1236 1232
rect 1230 1227 1236 1228
rect 1390 1232 1396 1233
rect 1390 1228 1391 1232
rect 1395 1228 1396 1232
rect 1390 1227 1396 1228
rect 1550 1232 1556 1233
rect 1550 1228 1551 1232
rect 1555 1228 1556 1232
rect 1550 1227 1556 1228
rect 1718 1232 1724 1233
rect 1718 1228 1719 1232
rect 1723 1228 1724 1232
rect 2006 1231 2007 1235
rect 2011 1231 2012 1235
rect 2006 1230 2012 1231
rect 1718 1227 1724 1228
rect 2070 1200 2076 1201
rect 2046 1197 2052 1198
rect 2046 1193 2047 1197
rect 2051 1193 2052 1197
rect 2070 1196 2071 1200
rect 2075 1196 2076 1200
rect 2070 1195 2076 1196
rect 2182 1200 2188 1201
rect 2182 1196 2183 1200
rect 2187 1196 2188 1200
rect 2182 1195 2188 1196
rect 2302 1200 2308 1201
rect 2302 1196 2303 1200
rect 2307 1196 2308 1200
rect 2302 1195 2308 1196
rect 2430 1200 2436 1201
rect 2430 1196 2431 1200
rect 2435 1196 2436 1200
rect 2430 1195 2436 1196
rect 2558 1200 2564 1201
rect 2558 1196 2559 1200
rect 2563 1196 2564 1200
rect 2558 1195 2564 1196
rect 2710 1200 2716 1201
rect 2710 1196 2711 1200
rect 2715 1196 2716 1200
rect 2710 1195 2716 1196
rect 2886 1200 2892 1201
rect 2886 1196 2887 1200
rect 2891 1196 2892 1200
rect 2886 1195 2892 1196
rect 3086 1200 3092 1201
rect 3086 1196 3087 1200
rect 3091 1196 3092 1200
rect 3086 1195 3092 1196
rect 3310 1200 3316 1201
rect 3310 1196 3311 1200
rect 3315 1196 3316 1200
rect 3310 1195 3316 1196
rect 3542 1200 3548 1201
rect 3542 1196 3543 1200
rect 3547 1196 3548 1200
rect 3542 1195 3548 1196
rect 3782 1200 3788 1201
rect 3782 1196 3783 1200
rect 3787 1196 3788 1200
rect 3782 1195 3788 1196
rect 3942 1197 3948 1198
rect 2046 1192 2052 1193
rect 3942 1193 3943 1197
rect 3947 1193 3948 1197
rect 3942 1192 3948 1193
rect 2070 1181 2076 1182
rect 2046 1180 2052 1181
rect 2046 1176 2047 1180
rect 2051 1176 2052 1180
rect 2070 1177 2071 1181
rect 2075 1177 2076 1181
rect 2070 1176 2076 1177
rect 2182 1181 2188 1182
rect 2182 1177 2183 1181
rect 2187 1177 2188 1181
rect 2182 1176 2188 1177
rect 2302 1181 2308 1182
rect 2302 1177 2303 1181
rect 2307 1177 2308 1181
rect 2302 1176 2308 1177
rect 2430 1181 2436 1182
rect 2430 1177 2431 1181
rect 2435 1177 2436 1181
rect 2430 1176 2436 1177
rect 2558 1181 2564 1182
rect 2558 1177 2559 1181
rect 2563 1177 2564 1181
rect 2558 1176 2564 1177
rect 2710 1181 2716 1182
rect 2710 1177 2711 1181
rect 2715 1177 2716 1181
rect 2710 1176 2716 1177
rect 2886 1181 2892 1182
rect 2886 1177 2887 1181
rect 2891 1177 2892 1181
rect 2886 1176 2892 1177
rect 3086 1181 3092 1182
rect 3086 1177 3087 1181
rect 3091 1177 3092 1181
rect 3086 1176 3092 1177
rect 3310 1181 3316 1182
rect 3310 1177 3311 1181
rect 3315 1177 3316 1181
rect 3310 1176 3316 1177
rect 3542 1181 3548 1182
rect 3542 1177 3543 1181
rect 3547 1177 3548 1181
rect 3542 1176 3548 1177
rect 3782 1181 3788 1182
rect 3782 1177 3783 1181
rect 3787 1177 3788 1181
rect 3782 1176 3788 1177
rect 3942 1180 3948 1181
rect 3942 1176 3943 1180
rect 3947 1176 3948 1180
rect 2046 1175 2052 1176
rect 3942 1175 3948 1176
rect 166 1172 172 1173
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 166 1168 167 1172
rect 171 1168 172 1172
rect 166 1167 172 1168
rect 302 1172 308 1173
rect 302 1168 303 1172
rect 307 1168 308 1172
rect 302 1167 308 1168
rect 462 1172 468 1173
rect 462 1168 463 1172
rect 467 1168 468 1172
rect 462 1167 468 1168
rect 630 1172 636 1173
rect 630 1168 631 1172
rect 635 1168 636 1172
rect 630 1167 636 1168
rect 806 1172 812 1173
rect 806 1168 807 1172
rect 811 1168 812 1172
rect 806 1167 812 1168
rect 982 1172 988 1173
rect 982 1168 983 1172
rect 987 1168 988 1172
rect 982 1167 988 1168
rect 1158 1172 1164 1173
rect 1158 1168 1159 1172
rect 1163 1168 1164 1172
rect 1158 1167 1164 1168
rect 1334 1172 1340 1173
rect 1334 1168 1335 1172
rect 1339 1168 1340 1172
rect 1334 1167 1340 1168
rect 1510 1172 1516 1173
rect 1510 1168 1511 1172
rect 1515 1168 1516 1172
rect 1510 1167 1516 1168
rect 1694 1172 1700 1173
rect 1694 1168 1695 1172
rect 1699 1168 1700 1172
rect 1694 1167 1700 1168
rect 2006 1169 2012 1170
rect 110 1164 116 1165
rect 2006 1165 2007 1169
rect 2011 1165 2012 1169
rect 2006 1164 2012 1165
rect 166 1153 172 1154
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 166 1149 167 1153
rect 171 1149 172 1153
rect 166 1148 172 1149
rect 302 1153 308 1154
rect 302 1149 303 1153
rect 307 1149 308 1153
rect 302 1148 308 1149
rect 462 1153 468 1154
rect 462 1149 463 1153
rect 467 1149 468 1153
rect 462 1148 468 1149
rect 630 1153 636 1154
rect 630 1149 631 1153
rect 635 1149 636 1153
rect 630 1148 636 1149
rect 806 1153 812 1154
rect 806 1149 807 1153
rect 811 1149 812 1153
rect 806 1148 812 1149
rect 982 1153 988 1154
rect 982 1149 983 1153
rect 987 1149 988 1153
rect 982 1148 988 1149
rect 1158 1153 1164 1154
rect 1158 1149 1159 1153
rect 1163 1149 1164 1153
rect 1158 1148 1164 1149
rect 1334 1153 1340 1154
rect 1334 1149 1335 1153
rect 1339 1149 1340 1153
rect 1334 1148 1340 1149
rect 1510 1153 1516 1154
rect 1510 1149 1511 1153
rect 1515 1149 1516 1153
rect 1510 1148 1516 1149
rect 1694 1153 1700 1154
rect 1694 1149 1695 1153
rect 1699 1149 1700 1153
rect 1694 1148 1700 1149
rect 2006 1152 2012 1153
rect 2006 1148 2007 1152
rect 2011 1148 2012 1152
rect 110 1147 116 1148
rect 2006 1147 2012 1148
rect 2046 1124 2052 1125
rect 3942 1124 3948 1125
rect 2046 1120 2047 1124
rect 2051 1120 2052 1124
rect 2046 1119 2052 1120
rect 2070 1123 2076 1124
rect 2070 1119 2071 1123
rect 2075 1119 2076 1123
rect 2070 1118 2076 1119
rect 2198 1123 2204 1124
rect 2198 1119 2199 1123
rect 2203 1119 2204 1123
rect 2198 1118 2204 1119
rect 2350 1123 2356 1124
rect 2350 1119 2351 1123
rect 2355 1119 2356 1123
rect 2350 1118 2356 1119
rect 2510 1123 2516 1124
rect 2510 1119 2511 1123
rect 2515 1119 2516 1123
rect 2510 1118 2516 1119
rect 2678 1123 2684 1124
rect 2678 1119 2679 1123
rect 2683 1119 2684 1123
rect 2678 1118 2684 1119
rect 2870 1123 2876 1124
rect 2870 1119 2871 1123
rect 2875 1119 2876 1123
rect 2870 1118 2876 1119
rect 3086 1123 3092 1124
rect 3086 1119 3087 1123
rect 3091 1119 3092 1123
rect 3086 1118 3092 1119
rect 3318 1123 3324 1124
rect 3318 1119 3319 1123
rect 3323 1119 3324 1123
rect 3318 1118 3324 1119
rect 3558 1123 3564 1124
rect 3558 1119 3559 1123
rect 3563 1119 3564 1123
rect 3558 1118 3564 1119
rect 3806 1123 3812 1124
rect 3806 1119 3807 1123
rect 3811 1119 3812 1123
rect 3942 1120 3943 1124
rect 3947 1120 3948 1124
rect 3942 1119 3948 1120
rect 3806 1118 3812 1119
rect 2046 1107 2052 1108
rect 2046 1103 2047 1107
rect 2051 1103 2052 1107
rect 3942 1107 3948 1108
rect 2046 1102 2052 1103
rect 2070 1104 2076 1105
rect 2070 1100 2071 1104
rect 2075 1100 2076 1104
rect 2070 1099 2076 1100
rect 2198 1104 2204 1105
rect 2198 1100 2199 1104
rect 2203 1100 2204 1104
rect 2198 1099 2204 1100
rect 2350 1104 2356 1105
rect 2350 1100 2351 1104
rect 2355 1100 2356 1104
rect 2350 1099 2356 1100
rect 2510 1104 2516 1105
rect 2510 1100 2511 1104
rect 2515 1100 2516 1104
rect 2510 1099 2516 1100
rect 2678 1104 2684 1105
rect 2678 1100 2679 1104
rect 2683 1100 2684 1104
rect 2678 1099 2684 1100
rect 2870 1104 2876 1105
rect 2870 1100 2871 1104
rect 2875 1100 2876 1104
rect 2870 1099 2876 1100
rect 3086 1104 3092 1105
rect 3086 1100 3087 1104
rect 3091 1100 3092 1104
rect 3086 1099 3092 1100
rect 3318 1104 3324 1105
rect 3318 1100 3319 1104
rect 3323 1100 3324 1104
rect 3318 1099 3324 1100
rect 3558 1104 3564 1105
rect 3558 1100 3559 1104
rect 3563 1100 3564 1104
rect 3558 1099 3564 1100
rect 3806 1104 3812 1105
rect 3806 1100 3807 1104
rect 3811 1100 3812 1104
rect 3942 1103 3943 1107
rect 3947 1103 3948 1107
rect 3942 1102 3948 1103
rect 3806 1099 3812 1100
rect 110 1096 116 1097
rect 2006 1096 2012 1097
rect 110 1092 111 1096
rect 115 1092 116 1096
rect 110 1091 116 1092
rect 134 1095 140 1096
rect 134 1091 135 1095
rect 139 1091 140 1095
rect 134 1090 140 1091
rect 238 1095 244 1096
rect 238 1091 239 1095
rect 243 1091 244 1095
rect 238 1090 244 1091
rect 374 1095 380 1096
rect 374 1091 375 1095
rect 379 1091 380 1095
rect 374 1090 380 1091
rect 526 1095 532 1096
rect 526 1091 527 1095
rect 531 1091 532 1095
rect 526 1090 532 1091
rect 694 1095 700 1096
rect 694 1091 695 1095
rect 699 1091 700 1095
rect 694 1090 700 1091
rect 862 1095 868 1096
rect 862 1091 863 1095
rect 867 1091 868 1095
rect 862 1090 868 1091
rect 1038 1095 1044 1096
rect 1038 1091 1039 1095
rect 1043 1091 1044 1095
rect 1038 1090 1044 1091
rect 1214 1095 1220 1096
rect 1214 1091 1215 1095
rect 1219 1091 1220 1095
rect 1214 1090 1220 1091
rect 1390 1095 1396 1096
rect 1390 1091 1391 1095
rect 1395 1091 1396 1095
rect 1390 1090 1396 1091
rect 1566 1095 1572 1096
rect 1566 1091 1567 1095
rect 1571 1091 1572 1095
rect 1566 1090 1572 1091
rect 1742 1095 1748 1096
rect 1742 1091 1743 1095
rect 1747 1091 1748 1095
rect 1742 1090 1748 1091
rect 1902 1095 1908 1096
rect 1902 1091 1903 1095
rect 1907 1091 1908 1095
rect 2006 1092 2007 1096
rect 2011 1092 2012 1096
rect 2006 1091 2012 1092
rect 1902 1090 1908 1091
rect 110 1079 116 1080
rect 110 1075 111 1079
rect 115 1075 116 1079
rect 2006 1079 2012 1080
rect 110 1074 116 1075
rect 134 1076 140 1077
rect 134 1072 135 1076
rect 139 1072 140 1076
rect 134 1071 140 1072
rect 238 1076 244 1077
rect 238 1072 239 1076
rect 243 1072 244 1076
rect 238 1071 244 1072
rect 374 1076 380 1077
rect 374 1072 375 1076
rect 379 1072 380 1076
rect 374 1071 380 1072
rect 526 1076 532 1077
rect 526 1072 527 1076
rect 531 1072 532 1076
rect 526 1071 532 1072
rect 694 1076 700 1077
rect 694 1072 695 1076
rect 699 1072 700 1076
rect 694 1071 700 1072
rect 862 1076 868 1077
rect 862 1072 863 1076
rect 867 1072 868 1076
rect 862 1071 868 1072
rect 1038 1076 1044 1077
rect 1038 1072 1039 1076
rect 1043 1072 1044 1076
rect 1038 1071 1044 1072
rect 1214 1076 1220 1077
rect 1214 1072 1215 1076
rect 1219 1072 1220 1076
rect 1214 1071 1220 1072
rect 1390 1076 1396 1077
rect 1390 1072 1391 1076
rect 1395 1072 1396 1076
rect 1390 1071 1396 1072
rect 1566 1076 1572 1077
rect 1566 1072 1567 1076
rect 1571 1072 1572 1076
rect 1566 1071 1572 1072
rect 1742 1076 1748 1077
rect 1742 1072 1743 1076
rect 1747 1072 1748 1076
rect 1742 1071 1748 1072
rect 1902 1076 1908 1077
rect 1902 1072 1903 1076
rect 1907 1072 1908 1076
rect 2006 1075 2007 1079
rect 2011 1075 2012 1079
rect 2006 1074 2012 1075
rect 1902 1071 1908 1072
rect 2070 1032 2076 1033
rect 2046 1029 2052 1030
rect 2046 1025 2047 1029
rect 2051 1025 2052 1029
rect 2070 1028 2071 1032
rect 2075 1028 2076 1032
rect 2070 1027 2076 1028
rect 2262 1032 2268 1033
rect 2262 1028 2263 1032
rect 2267 1028 2268 1032
rect 2262 1027 2268 1028
rect 2486 1032 2492 1033
rect 2486 1028 2487 1032
rect 2491 1028 2492 1032
rect 2486 1027 2492 1028
rect 2702 1032 2708 1033
rect 2702 1028 2703 1032
rect 2707 1028 2708 1032
rect 2702 1027 2708 1028
rect 2918 1032 2924 1033
rect 2918 1028 2919 1032
rect 2923 1028 2924 1032
rect 2918 1027 2924 1028
rect 3118 1032 3124 1033
rect 3118 1028 3119 1032
rect 3123 1028 3124 1032
rect 3118 1027 3124 1028
rect 3310 1032 3316 1033
rect 3310 1028 3311 1032
rect 3315 1028 3316 1032
rect 3310 1027 3316 1028
rect 3494 1032 3500 1033
rect 3494 1028 3495 1032
rect 3499 1028 3500 1032
rect 3494 1027 3500 1028
rect 3678 1032 3684 1033
rect 3678 1028 3679 1032
rect 3683 1028 3684 1032
rect 3678 1027 3684 1028
rect 3838 1032 3844 1033
rect 3838 1028 3839 1032
rect 3843 1028 3844 1032
rect 3838 1027 3844 1028
rect 3942 1029 3948 1030
rect 2046 1024 2052 1025
rect 3942 1025 3943 1029
rect 3947 1025 3948 1029
rect 3942 1024 3948 1025
rect 134 1016 140 1017
rect 110 1013 116 1014
rect 110 1009 111 1013
rect 115 1009 116 1013
rect 134 1012 135 1016
rect 139 1012 140 1016
rect 134 1011 140 1012
rect 286 1016 292 1017
rect 286 1012 287 1016
rect 291 1012 292 1016
rect 286 1011 292 1012
rect 470 1016 476 1017
rect 470 1012 471 1016
rect 475 1012 476 1016
rect 470 1011 476 1012
rect 654 1016 660 1017
rect 654 1012 655 1016
rect 659 1012 660 1016
rect 654 1011 660 1012
rect 838 1016 844 1017
rect 838 1012 839 1016
rect 843 1012 844 1016
rect 838 1011 844 1012
rect 1014 1016 1020 1017
rect 1014 1012 1015 1016
rect 1019 1012 1020 1016
rect 1014 1011 1020 1012
rect 1198 1016 1204 1017
rect 1198 1012 1199 1016
rect 1203 1012 1204 1016
rect 1198 1011 1204 1012
rect 1382 1016 1388 1017
rect 1382 1012 1383 1016
rect 1387 1012 1388 1016
rect 1382 1011 1388 1012
rect 1566 1016 1572 1017
rect 1566 1012 1567 1016
rect 1571 1012 1572 1016
rect 1566 1011 1572 1012
rect 2006 1013 2012 1014
rect 2070 1013 2076 1014
rect 110 1008 116 1009
rect 2006 1009 2007 1013
rect 2011 1009 2012 1013
rect 2006 1008 2012 1009
rect 2046 1012 2052 1013
rect 2046 1008 2047 1012
rect 2051 1008 2052 1012
rect 2070 1009 2071 1013
rect 2075 1009 2076 1013
rect 2070 1008 2076 1009
rect 2262 1013 2268 1014
rect 2262 1009 2263 1013
rect 2267 1009 2268 1013
rect 2262 1008 2268 1009
rect 2486 1013 2492 1014
rect 2486 1009 2487 1013
rect 2491 1009 2492 1013
rect 2486 1008 2492 1009
rect 2702 1013 2708 1014
rect 2702 1009 2703 1013
rect 2707 1009 2708 1013
rect 2702 1008 2708 1009
rect 2918 1013 2924 1014
rect 2918 1009 2919 1013
rect 2923 1009 2924 1013
rect 2918 1008 2924 1009
rect 3118 1013 3124 1014
rect 3118 1009 3119 1013
rect 3123 1009 3124 1013
rect 3118 1008 3124 1009
rect 3310 1013 3316 1014
rect 3310 1009 3311 1013
rect 3315 1009 3316 1013
rect 3310 1008 3316 1009
rect 3494 1013 3500 1014
rect 3494 1009 3495 1013
rect 3499 1009 3500 1013
rect 3494 1008 3500 1009
rect 3678 1013 3684 1014
rect 3678 1009 3679 1013
rect 3683 1009 3684 1013
rect 3678 1008 3684 1009
rect 3838 1013 3844 1014
rect 3838 1009 3839 1013
rect 3843 1009 3844 1013
rect 3838 1008 3844 1009
rect 3942 1012 3948 1013
rect 3942 1008 3943 1012
rect 3947 1008 3948 1012
rect 2046 1007 2052 1008
rect 3942 1007 3948 1008
rect 134 997 140 998
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 134 993 135 997
rect 139 993 140 997
rect 134 992 140 993
rect 286 997 292 998
rect 286 993 287 997
rect 291 993 292 997
rect 286 992 292 993
rect 470 997 476 998
rect 470 993 471 997
rect 475 993 476 997
rect 470 992 476 993
rect 654 997 660 998
rect 654 993 655 997
rect 659 993 660 997
rect 654 992 660 993
rect 838 997 844 998
rect 838 993 839 997
rect 843 993 844 997
rect 838 992 844 993
rect 1014 997 1020 998
rect 1014 993 1015 997
rect 1019 993 1020 997
rect 1014 992 1020 993
rect 1198 997 1204 998
rect 1198 993 1199 997
rect 1203 993 1204 997
rect 1198 992 1204 993
rect 1382 997 1388 998
rect 1382 993 1383 997
rect 1387 993 1388 997
rect 1382 992 1388 993
rect 1566 997 1572 998
rect 1566 993 1567 997
rect 1571 993 1572 997
rect 1566 992 1572 993
rect 2006 996 2012 997
rect 2006 992 2007 996
rect 2011 992 2012 996
rect 110 991 116 992
rect 2006 991 2012 992
rect 2046 956 2052 957
rect 3942 956 3948 957
rect 2046 952 2047 956
rect 2051 952 2052 956
rect 2046 951 2052 952
rect 2302 955 2308 956
rect 2302 951 2303 955
rect 2307 951 2308 955
rect 2302 950 2308 951
rect 2454 955 2460 956
rect 2454 951 2455 955
rect 2459 951 2460 955
rect 2454 950 2460 951
rect 2614 955 2620 956
rect 2614 951 2615 955
rect 2619 951 2620 955
rect 2614 950 2620 951
rect 2782 955 2788 956
rect 2782 951 2783 955
rect 2787 951 2788 955
rect 2782 950 2788 951
rect 2950 955 2956 956
rect 2950 951 2951 955
rect 2955 951 2956 955
rect 2950 950 2956 951
rect 3110 955 3116 956
rect 3110 951 3111 955
rect 3115 951 3116 955
rect 3110 950 3116 951
rect 3262 955 3268 956
rect 3262 951 3263 955
rect 3267 951 3268 955
rect 3262 950 3268 951
rect 3414 955 3420 956
rect 3414 951 3415 955
rect 3419 951 3420 955
rect 3414 950 3420 951
rect 3558 955 3564 956
rect 3558 951 3559 955
rect 3563 951 3564 955
rect 3558 950 3564 951
rect 3710 955 3716 956
rect 3710 951 3711 955
rect 3715 951 3716 955
rect 3710 950 3716 951
rect 3838 955 3844 956
rect 3838 951 3839 955
rect 3843 951 3844 955
rect 3942 952 3943 956
rect 3947 952 3948 956
rect 3942 951 3948 952
rect 3838 950 3844 951
rect 110 940 116 941
rect 2006 940 2012 941
rect 110 936 111 940
rect 115 936 116 940
rect 110 935 116 936
rect 134 939 140 940
rect 134 935 135 939
rect 139 935 140 939
rect 134 934 140 935
rect 294 939 300 940
rect 294 935 295 939
rect 299 935 300 939
rect 294 934 300 935
rect 470 939 476 940
rect 470 935 471 939
rect 475 935 476 939
rect 470 934 476 935
rect 638 939 644 940
rect 638 935 639 939
rect 643 935 644 939
rect 638 934 644 935
rect 798 939 804 940
rect 798 935 799 939
rect 803 935 804 939
rect 798 934 804 935
rect 950 939 956 940
rect 950 935 951 939
rect 955 935 956 939
rect 950 934 956 935
rect 1086 939 1092 940
rect 1086 935 1087 939
rect 1091 935 1092 939
rect 1086 934 1092 935
rect 1222 939 1228 940
rect 1222 935 1223 939
rect 1227 935 1228 939
rect 1222 934 1228 935
rect 1358 939 1364 940
rect 1358 935 1359 939
rect 1363 935 1364 939
rect 1358 934 1364 935
rect 1494 939 1500 940
rect 1494 935 1495 939
rect 1499 935 1500 939
rect 2006 936 2007 940
rect 2011 936 2012 940
rect 2006 935 2012 936
rect 2046 939 2052 940
rect 2046 935 2047 939
rect 2051 935 2052 939
rect 3942 939 3948 940
rect 1494 934 1500 935
rect 2046 934 2052 935
rect 2302 936 2308 937
rect 2302 932 2303 936
rect 2307 932 2308 936
rect 2302 931 2308 932
rect 2454 936 2460 937
rect 2454 932 2455 936
rect 2459 932 2460 936
rect 2454 931 2460 932
rect 2614 936 2620 937
rect 2614 932 2615 936
rect 2619 932 2620 936
rect 2614 931 2620 932
rect 2782 936 2788 937
rect 2782 932 2783 936
rect 2787 932 2788 936
rect 2782 931 2788 932
rect 2950 936 2956 937
rect 2950 932 2951 936
rect 2955 932 2956 936
rect 2950 931 2956 932
rect 3110 936 3116 937
rect 3110 932 3111 936
rect 3115 932 3116 936
rect 3110 931 3116 932
rect 3262 936 3268 937
rect 3262 932 3263 936
rect 3267 932 3268 936
rect 3262 931 3268 932
rect 3414 936 3420 937
rect 3414 932 3415 936
rect 3419 932 3420 936
rect 3414 931 3420 932
rect 3558 936 3564 937
rect 3558 932 3559 936
rect 3563 932 3564 936
rect 3558 931 3564 932
rect 3710 936 3716 937
rect 3710 932 3711 936
rect 3715 932 3716 936
rect 3710 931 3716 932
rect 3838 936 3844 937
rect 3838 932 3839 936
rect 3843 932 3844 936
rect 3942 935 3943 939
rect 3947 935 3948 939
rect 3942 934 3948 935
rect 3838 931 3844 932
rect 110 923 116 924
rect 110 919 111 923
rect 115 919 116 923
rect 2006 923 2012 924
rect 110 918 116 919
rect 134 920 140 921
rect 134 916 135 920
rect 139 916 140 920
rect 134 915 140 916
rect 294 920 300 921
rect 294 916 295 920
rect 299 916 300 920
rect 294 915 300 916
rect 470 920 476 921
rect 470 916 471 920
rect 475 916 476 920
rect 470 915 476 916
rect 638 920 644 921
rect 638 916 639 920
rect 643 916 644 920
rect 638 915 644 916
rect 798 920 804 921
rect 798 916 799 920
rect 803 916 804 920
rect 798 915 804 916
rect 950 920 956 921
rect 950 916 951 920
rect 955 916 956 920
rect 950 915 956 916
rect 1086 920 1092 921
rect 1086 916 1087 920
rect 1091 916 1092 920
rect 1086 915 1092 916
rect 1222 920 1228 921
rect 1222 916 1223 920
rect 1227 916 1228 920
rect 1222 915 1228 916
rect 1358 920 1364 921
rect 1358 916 1359 920
rect 1363 916 1364 920
rect 1358 915 1364 916
rect 1494 920 1500 921
rect 1494 916 1495 920
rect 1499 916 1500 920
rect 2006 919 2007 923
rect 2011 919 2012 923
rect 2006 918 2012 919
rect 1494 915 1500 916
rect 2558 872 2564 873
rect 2046 869 2052 870
rect 2046 865 2047 869
rect 2051 865 2052 869
rect 2558 868 2559 872
rect 2563 868 2564 872
rect 2558 867 2564 868
rect 2678 872 2684 873
rect 2678 868 2679 872
rect 2683 868 2684 872
rect 2678 867 2684 868
rect 2806 872 2812 873
rect 2806 868 2807 872
rect 2811 868 2812 872
rect 2806 867 2812 868
rect 2942 872 2948 873
rect 2942 868 2943 872
rect 2947 868 2948 872
rect 2942 867 2948 868
rect 3078 872 3084 873
rect 3078 868 3079 872
rect 3083 868 3084 872
rect 3078 867 3084 868
rect 3206 872 3212 873
rect 3206 868 3207 872
rect 3211 868 3212 872
rect 3206 867 3212 868
rect 3334 872 3340 873
rect 3334 868 3335 872
rect 3339 868 3340 872
rect 3334 867 3340 868
rect 3462 872 3468 873
rect 3462 868 3463 872
rect 3467 868 3468 872
rect 3462 867 3468 868
rect 3590 872 3596 873
rect 3590 868 3591 872
rect 3595 868 3596 872
rect 3590 867 3596 868
rect 3726 872 3732 873
rect 3726 868 3727 872
rect 3731 868 3732 872
rect 3726 867 3732 868
rect 3838 872 3844 873
rect 3838 868 3839 872
rect 3843 868 3844 872
rect 3838 867 3844 868
rect 3942 869 3948 870
rect 2046 864 2052 865
rect 3942 865 3943 869
rect 3947 865 3948 869
rect 3942 864 3948 865
rect 158 860 164 861
rect 110 857 116 858
rect 110 853 111 857
rect 115 853 116 857
rect 158 856 159 860
rect 163 856 164 860
rect 158 855 164 856
rect 318 860 324 861
rect 318 856 319 860
rect 323 856 324 860
rect 318 855 324 856
rect 470 860 476 861
rect 470 856 471 860
rect 475 856 476 860
rect 470 855 476 856
rect 614 860 620 861
rect 614 856 615 860
rect 619 856 620 860
rect 614 855 620 856
rect 750 860 756 861
rect 750 856 751 860
rect 755 856 756 860
rect 750 855 756 856
rect 878 860 884 861
rect 878 856 879 860
rect 883 856 884 860
rect 878 855 884 856
rect 998 860 1004 861
rect 998 856 999 860
rect 1003 856 1004 860
rect 998 855 1004 856
rect 1110 860 1116 861
rect 1110 856 1111 860
rect 1115 856 1116 860
rect 1110 855 1116 856
rect 1230 860 1236 861
rect 1230 856 1231 860
rect 1235 856 1236 860
rect 1230 855 1236 856
rect 1350 860 1356 861
rect 1350 856 1351 860
rect 1355 856 1356 860
rect 1350 855 1356 856
rect 2006 857 2012 858
rect 110 852 116 853
rect 2006 853 2007 857
rect 2011 853 2012 857
rect 2558 853 2564 854
rect 2006 852 2012 853
rect 2046 852 2052 853
rect 2046 848 2047 852
rect 2051 848 2052 852
rect 2558 849 2559 853
rect 2563 849 2564 853
rect 2558 848 2564 849
rect 2678 853 2684 854
rect 2678 849 2679 853
rect 2683 849 2684 853
rect 2678 848 2684 849
rect 2806 853 2812 854
rect 2806 849 2807 853
rect 2811 849 2812 853
rect 2806 848 2812 849
rect 2942 853 2948 854
rect 2942 849 2943 853
rect 2947 849 2948 853
rect 2942 848 2948 849
rect 3078 853 3084 854
rect 3078 849 3079 853
rect 3083 849 3084 853
rect 3078 848 3084 849
rect 3206 853 3212 854
rect 3206 849 3207 853
rect 3211 849 3212 853
rect 3206 848 3212 849
rect 3334 853 3340 854
rect 3334 849 3335 853
rect 3339 849 3340 853
rect 3334 848 3340 849
rect 3462 853 3468 854
rect 3462 849 3463 853
rect 3467 849 3468 853
rect 3462 848 3468 849
rect 3590 853 3596 854
rect 3590 849 3591 853
rect 3595 849 3596 853
rect 3590 848 3596 849
rect 3726 853 3732 854
rect 3726 849 3727 853
rect 3731 849 3732 853
rect 3726 848 3732 849
rect 3838 853 3844 854
rect 3838 849 3839 853
rect 3843 849 3844 853
rect 3838 848 3844 849
rect 3942 852 3948 853
rect 3942 848 3943 852
rect 3947 848 3948 852
rect 2046 847 2052 848
rect 3942 847 3948 848
rect 158 841 164 842
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 158 837 159 841
rect 163 837 164 841
rect 158 836 164 837
rect 318 841 324 842
rect 318 837 319 841
rect 323 837 324 841
rect 318 836 324 837
rect 470 841 476 842
rect 470 837 471 841
rect 475 837 476 841
rect 470 836 476 837
rect 614 841 620 842
rect 614 837 615 841
rect 619 837 620 841
rect 614 836 620 837
rect 750 841 756 842
rect 750 837 751 841
rect 755 837 756 841
rect 750 836 756 837
rect 878 841 884 842
rect 878 837 879 841
rect 883 837 884 841
rect 878 836 884 837
rect 998 841 1004 842
rect 998 837 999 841
rect 1003 837 1004 841
rect 998 836 1004 837
rect 1110 841 1116 842
rect 1110 837 1111 841
rect 1115 837 1116 841
rect 1110 836 1116 837
rect 1230 841 1236 842
rect 1230 837 1231 841
rect 1235 837 1236 841
rect 1230 836 1236 837
rect 1350 841 1356 842
rect 1350 837 1351 841
rect 1355 837 1356 841
rect 1350 836 1356 837
rect 2006 840 2012 841
rect 2006 836 2007 840
rect 2011 836 2012 840
rect 110 835 116 836
rect 2006 835 2012 836
rect 2046 796 2052 797
rect 3942 796 3948 797
rect 2046 792 2047 796
rect 2051 792 2052 796
rect 2046 791 2052 792
rect 2334 795 2340 796
rect 2334 791 2335 795
rect 2339 791 2340 795
rect 2334 790 2340 791
rect 2470 795 2476 796
rect 2470 791 2471 795
rect 2475 791 2476 795
rect 2470 790 2476 791
rect 2614 795 2620 796
rect 2614 791 2615 795
rect 2619 791 2620 795
rect 2614 790 2620 791
rect 2766 795 2772 796
rect 2766 791 2767 795
rect 2771 791 2772 795
rect 2766 790 2772 791
rect 2918 795 2924 796
rect 2918 791 2919 795
rect 2923 791 2924 795
rect 2918 790 2924 791
rect 3078 795 3084 796
rect 3078 791 3079 795
rect 3083 791 3084 795
rect 3078 790 3084 791
rect 3238 795 3244 796
rect 3238 791 3239 795
rect 3243 791 3244 795
rect 3238 790 3244 791
rect 3390 795 3396 796
rect 3390 791 3391 795
rect 3395 791 3396 795
rect 3390 790 3396 791
rect 3542 795 3548 796
rect 3542 791 3543 795
rect 3547 791 3548 795
rect 3542 790 3548 791
rect 3702 795 3708 796
rect 3702 791 3703 795
rect 3707 791 3708 795
rect 3702 790 3708 791
rect 3838 795 3844 796
rect 3838 791 3839 795
rect 3843 791 3844 795
rect 3942 792 3943 796
rect 3947 792 3948 796
rect 3942 791 3948 792
rect 3838 790 3844 791
rect 110 788 116 789
rect 2006 788 2012 789
rect 110 784 111 788
rect 115 784 116 788
rect 110 783 116 784
rect 222 787 228 788
rect 222 783 223 787
rect 227 783 228 787
rect 222 782 228 783
rect 382 787 388 788
rect 382 783 383 787
rect 387 783 388 787
rect 382 782 388 783
rect 534 787 540 788
rect 534 783 535 787
rect 539 783 540 787
rect 534 782 540 783
rect 678 787 684 788
rect 678 783 679 787
rect 683 783 684 787
rect 678 782 684 783
rect 814 787 820 788
rect 814 783 815 787
rect 819 783 820 787
rect 814 782 820 783
rect 950 787 956 788
rect 950 783 951 787
rect 955 783 956 787
rect 950 782 956 783
rect 1078 787 1084 788
rect 1078 783 1079 787
rect 1083 783 1084 787
rect 1078 782 1084 783
rect 1198 787 1204 788
rect 1198 783 1199 787
rect 1203 783 1204 787
rect 1198 782 1204 783
rect 1326 787 1332 788
rect 1326 783 1327 787
rect 1331 783 1332 787
rect 1326 782 1332 783
rect 1454 787 1460 788
rect 1454 783 1455 787
rect 1459 783 1460 787
rect 2006 784 2007 788
rect 2011 784 2012 788
rect 2006 783 2012 784
rect 1454 782 1460 783
rect 2046 779 2052 780
rect 2046 775 2047 779
rect 2051 775 2052 779
rect 3942 779 3948 780
rect 2046 774 2052 775
rect 2334 776 2340 777
rect 2334 772 2335 776
rect 2339 772 2340 776
rect 110 771 116 772
rect 110 767 111 771
rect 115 767 116 771
rect 2006 771 2012 772
rect 2334 771 2340 772
rect 2470 776 2476 777
rect 2470 772 2471 776
rect 2475 772 2476 776
rect 2470 771 2476 772
rect 2614 776 2620 777
rect 2614 772 2615 776
rect 2619 772 2620 776
rect 2614 771 2620 772
rect 2766 776 2772 777
rect 2766 772 2767 776
rect 2771 772 2772 776
rect 2766 771 2772 772
rect 2918 776 2924 777
rect 2918 772 2919 776
rect 2923 772 2924 776
rect 2918 771 2924 772
rect 3078 776 3084 777
rect 3078 772 3079 776
rect 3083 772 3084 776
rect 3078 771 3084 772
rect 3238 776 3244 777
rect 3238 772 3239 776
rect 3243 772 3244 776
rect 3238 771 3244 772
rect 3390 776 3396 777
rect 3390 772 3391 776
rect 3395 772 3396 776
rect 3390 771 3396 772
rect 3542 776 3548 777
rect 3542 772 3543 776
rect 3547 772 3548 776
rect 3542 771 3548 772
rect 3702 776 3708 777
rect 3702 772 3703 776
rect 3707 772 3708 776
rect 3702 771 3708 772
rect 3838 776 3844 777
rect 3838 772 3839 776
rect 3843 772 3844 776
rect 3942 775 3943 779
rect 3947 775 3948 779
rect 3942 774 3948 775
rect 3838 771 3844 772
rect 110 766 116 767
rect 222 768 228 769
rect 222 764 223 768
rect 227 764 228 768
rect 222 763 228 764
rect 382 768 388 769
rect 382 764 383 768
rect 387 764 388 768
rect 382 763 388 764
rect 534 768 540 769
rect 534 764 535 768
rect 539 764 540 768
rect 534 763 540 764
rect 678 768 684 769
rect 678 764 679 768
rect 683 764 684 768
rect 678 763 684 764
rect 814 768 820 769
rect 814 764 815 768
rect 819 764 820 768
rect 814 763 820 764
rect 950 768 956 769
rect 950 764 951 768
rect 955 764 956 768
rect 950 763 956 764
rect 1078 768 1084 769
rect 1078 764 1079 768
rect 1083 764 1084 768
rect 1078 763 1084 764
rect 1198 768 1204 769
rect 1198 764 1199 768
rect 1203 764 1204 768
rect 1198 763 1204 764
rect 1326 768 1332 769
rect 1326 764 1327 768
rect 1331 764 1332 768
rect 1326 763 1332 764
rect 1454 768 1460 769
rect 1454 764 1455 768
rect 1459 764 1460 768
rect 2006 767 2007 771
rect 2011 767 2012 771
rect 2006 766 2012 767
rect 1454 763 1460 764
rect 2070 712 2076 713
rect 2046 709 2052 710
rect 2046 705 2047 709
rect 2051 705 2052 709
rect 2070 708 2071 712
rect 2075 708 2076 712
rect 2070 707 2076 708
rect 2182 712 2188 713
rect 2182 708 2183 712
rect 2187 708 2188 712
rect 2182 707 2188 708
rect 2334 712 2340 713
rect 2334 708 2335 712
rect 2339 708 2340 712
rect 2334 707 2340 708
rect 2486 712 2492 713
rect 2486 708 2487 712
rect 2491 708 2492 712
rect 2486 707 2492 708
rect 2638 712 2644 713
rect 2638 708 2639 712
rect 2643 708 2644 712
rect 2638 707 2644 708
rect 2806 712 2812 713
rect 2806 708 2807 712
rect 2811 708 2812 712
rect 2806 707 2812 708
rect 2982 712 2988 713
rect 2982 708 2983 712
rect 2987 708 2988 712
rect 2982 707 2988 708
rect 3166 712 3172 713
rect 3166 708 3167 712
rect 3171 708 3172 712
rect 3166 707 3172 708
rect 3366 712 3372 713
rect 3366 708 3367 712
rect 3371 708 3372 712
rect 3366 707 3372 708
rect 3574 712 3580 713
rect 3574 708 3575 712
rect 3579 708 3580 712
rect 3574 707 3580 708
rect 3782 712 3788 713
rect 3782 708 3783 712
rect 3787 708 3788 712
rect 3782 707 3788 708
rect 3942 709 3948 710
rect 310 704 316 705
rect 110 701 116 702
rect 110 697 111 701
rect 115 697 116 701
rect 310 700 311 704
rect 315 700 316 704
rect 310 699 316 700
rect 470 704 476 705
rect 470 700 471 704
rect 475 700 476 704
rect 470 699 476 700
rect 638 704 644 705
rect 638 700 639 704
rect 643 700 644 704
rect 638 699 644 700
rect 806 704 812 705
rect 806 700 807 704
rect 811 700 812 704
rect 806 699 812 700
rect 974 704 980 705
rect 974 700 975 704
rect 979 700 980 704
rect 974 699 980 700
rect 1134 704 1140 705
rect 1134 700 1135 704
rect 1139 700 1140 704
rect 1134 699 1140 700
rect 1294 704 1300 705
rect 1294 700 1295 704
rect 1299 700 1300 704
rect 1294 699 1300 700
rect 1454 704 1460 705
rect 1454 700 1455 704
rect 1459 700 1460 704
rect 1454 699 1460 700
rect 1606 704 1612 705
rect 1606 700 1607 704
rect 1611 700 1612 704
rect 1606 699 1612 700
rect 1766 704 1772 705
rect 1766 700 1767 704
rect 1771 700 1772 704
rect 1766 699 1772 700
rect 1902 704 1908 705
rect 2046 704 2052 705
rect 3942 705 3943 709
rect 3947 705 3948 709
rect 3942 704 3948 705
rect 1902 700 1903 704
rect 1907 700 1908 704
rect 1902 699 1908 700
rect 2006 701 2012 702
rect 110 696 116 697
rect 2006 697 2007 701
rect 2011 697 2012 701
rect 2006 696 2012 697
rect 2070 693 2076 694
rect 2046 692 2052 693
rect 2046 688 2047 692
rect 2051 688 2052 692
rect 2070 689 2071 693
rect 2075 689 2076 693
rect 2070 688 2076 689
rect 2182 693 2188 694
rect 2182 689 2183 693
rect 2187 689 2188 693
rect 2182 688 2188 689
rect 2334 693 2340 694
rect 2334 689 2335 693
rect 2339 689 2340 693
rect 2334 688 2340 689
rect 2486 693 2492 694
rect 2486 689 2487 693
rect 2491 689 2492 693
rect 2486 688 2492 689
rect 2638 693 2644 694
rect 2638 689 2639 693
rect 2643 689 2644 693
rect 2638 688 2644 689
rect 2806 693 2812 694
rect 2806 689 2807 693
rect 2811 689 2812 693
rect 2806 688 2812 689
rect 2982 693 2988 694
rect 2982 689 2983 693
rect 2987 689 2988 693
rect 2982 688 2988 689
rect 3166 693 3172 694
rect 3166 689 3167 693
rect 3171 689 3172 693
rect 3166 688 3172 689
rect 3366 693 3372 694
rect 3366 689 3367 693
rect 3371 689 3372 693
rect 3366 688 3372 689
rect 3574 693 3580 694
rect 3574 689 3575 693
rect 3579 689 3580 693
rect 3574 688 3580 689
rect 3782 693 3788 694
rect 3782 689 3783 693
rect 3787 689 3788 693
rect 3782 688 3788 689
rect 3942 692 3948 693
rect 3942 688 3943 692
rect 3947 688 3948 692
rect 2046 687 2052 688
rect 3942 687 3948 688
rect 310 685 316 686
rect 110 684 116 685
rect 110 680 111 684
rect 115 680 116 684
rect 310 681 311 685
rect 315 681 316 685
rect 310 680 316 681
rect 470 685 476 686
rect 470 681 471 685
rect 475 681 476 685
rect 470 680 476 681
rect 638 685 644 686
rect 638 681 639 685
rect 643 681 644 685
rect 638 680 644 681
rect 806 685 812 686
rect 806 681 807 685
rect 811 681 812 685
rect 806 680 812 681
rect 974 685 980 686
rect 974 681 975 685
rect 979 681 980 685
rect 974 680 980 681
rect 1134 685 1140 686
rect 1134 681 1135 685
rect 1139 681 1140 685
rect 1134 680 1140 681
rect 1294 685 1300 686
rect 1294 681 1295 685
rect 1299 681 1300 685
rect 1294 680 1300 681
rect 1454 685 1460 686
rect 1454 681 1455 685
rect 1459 681 1460 685
rect 1454 680 1460 681
rect 1606 685 1612 686
rect 1606 681 1607 685
rect 1611 681 1612 685
rect 1606 680 1612 681
rect 1766 685 1772 686
rect 1766 681 1767 685
rect 1771 681 1772 685
rect 1766 680 1772 681
rect 1902 685 1908 686
rect 1902 681 1903 685
rect 1907 681 1908 685
rect 1902 680 1908 681
rect 2006 684 2012 685
rect 2006 680 2007 684
rect 2011 680 2012 684
rect 110 679 116 680
rect 2006 679 2012 680
rect 110 632 116 633
rect 2006 632 2012 633
rect 110 628 111 632
rect 115 628 116 632
rect 110 627 116 628
rect 294 631 300 632
rect 294 627 295 631
rect 299 627 300 631
rect 294 626 300 627
rect 446 631 452 632
rect 446 627 447 631
rect 451 627 452 631
rect 446 626 452 627
rect 614 631 620 632
rect 614 627 615 631
rect 619 627 620 631
rect 614 626 620 627
rect 782 631 788 632
rect 782 627 783 631
rect 787 627 788 631
rect 782 626 788 627
rect 950 631 956 632
rect 950 627 951 631
rect 955 627 956 631
rect 950 626 956 627
rect 1110 631 1116 632
rect 1110 627 1111 631
rect 1115 627 1116 631
rect 1110 626 1116 627
rect 1262 631 1268 632
rect 1262 627 1263 631
rect 1267 627 1268 631
rect 1262 626 1268 627
rect 1398 631 1404 632
rect 1398 627 1399 631
rect 1403 627 1404 631
rect 1398 626 1404 627
rect 1534 631 1540 632
rect 1534 627 1535 631
rect 1539 627 1540 631
rect 1534 626 1540 627
rect 1662 631 1668 632
rect 1662 627 1663 631
rect 1667 627 1668 631
rect 1662 626 1668 627
rect 1790 631 1796 632
rect 1790 627 1791 631
rect 1795 627 1796 631
rect 1790 626 1796 627
rect 1902 631 1908 632
rect 1902 627 1903 631
rect 1907 627 1908 631
rect 2006 628 2007 632
rect 2011 628 2012 632
rect 2006 627 2012 628
rect 2046 628 2052 629
rect 3942 628 3948 629
rect 1902 626 1908 627
rect 2046 624 2047 628
rect 2051 624 2052 628
rect 2046 623 2052 624
rect 2070 627 2076 628
rect 2070 623 2071 627
rect 2075 623 2076 627
rect 2070 622 2076 623
rect 2238 627 2244 628
rect 2238 623 2239 627
rect 2243 623 2244 627
rect 2238 622 2244 623
rect 2422 627 2428 628
rect 2422 623 2423 627
rect 2427 623 2428 627
rect 2422 622 2428 623
rect 2622 627 2628 628
rect 2622 623 2623 627
rect 2627 623 2628 627
rect 2622 622 2628 623
rect 2838 627 2844 628
rect 2838 623 2839 627
rect 2843 623 2844 627
rect 2838 622 2844 623
rect 3070 627 3076 628
rect 3070 623 3071 627
rect 3075 623 3076 627
rect 3070 622 3076 623
rect 3318 627 3324 628
rect 3318 623 3319 627
rect 3323 623 3324 627
rect 3318 622 3324 623
rect 3574 627 3580 628
rect 3574 623 3575 627
rect 3579 623 3580 627
rect 3574 622 3580 623
rect 3838 627 3844 628
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3942 624 3943 628
rect 3947 624 3948 628
rect 3942 623 3948 624
rect 3838 622 3844 623
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 2006 615 2012 616
rect 110 610 116 611
rect 294 612 300 613
rect 294 608 295 612
rect 299 608 300 612
rect 294 607 300 608
rect 446 612 452 613
rect 446 608 447 612
rect 451 608 452 612
rect 446 607 452 608
rect 614 612 620 613
rect 614 608 615 612
rect 619 608 620 612
rect 614 607 620 608
rect 782 612 788 613
rect 782 608 783 612
rect 787 608 788 612
rect 782 607 788 608
rect 950 612 956 613
rect 950 608 951 612
rect 955 608 956 612
rect 950 607 956 608
rect 1110 612 1116 613
rect 1110 608 1111 612
rect 1115 608 1116 612
rect 1110 607 1116 608
rect 1262 612 1268 613
rect 1262 608 1263 612
rect 1267 608 1268 612
rect 1262 607 1268 608
rect 1398 612 1404 613
rect 1398 608 1399 612
rect 1403 608 1404 612
rect 1398 607 1404 608
rect 1534 612 1540 613
rect 1534 608 1535 612
rect 1539 608 1540 612
rect 1534 607 1540 608
rect 1662 612 1668 613
rect 1662 608 1663 612
rect 1667 608 1668 612
rect 1662 607 1668 608
rect 1790 612 1796 613
rect 1790 608 1791 612
rect 1795 608 1796 612
rect 1790 607 1796 608
rect 1902 612 1908 613
rect 1902 608 1903 612
rect 1907 608 1908 612
rect 2006 611 2007 615
rect 2011 611 2012 615
rect 2006 610 2012 611
rect 2046 611 2052 612
rect 1902 607 1908 608
rect 2046 607 2047 611
rect 2051 607 2052 611
rect 3942 611 3948 612
rect 2046 606 2052 607
rect 2070 608 2076 609
rect 2070 604 2071 608
rect 2075 604 2076 608
rect 2070 603 2076 604
rect 2238 608 2244 609
rect 2238 604 2239 608
rect 2243 604 2244 608
rect 2238 603 2244 604
rect 2422 608 2428 609
rect 2422 604 2423 608
rect 2427 604 2428 608
rect 2422 603 2428 604
rect 2622 608 2628 609
rect 2622 604 2623 608
rect 2627 604 2628 608
rect 2622 603 2628 604
rect 2838 608 2844 609
rect 2838 604 2839 608
rect 2843 604 2844 608
rect 2838 603 2844 604
rect 3070 608 3076 609
rect 3070 604 3071 608
rect 3075 604 3076 608
rect 3070 603 3076 604
rect 3318 608 3324 609
rect 3318 604 3319 608
rect 3323 604 3324 608
rect 3318 603 3324 604
rect 3574 608 3580 609
rect 3574 604 3575 608
rect 3579 604 3580 608
rect 3574 603 3580 604
rect 3838 608 3844 609
rect 3838 604 3839 608
rect 3843 604 3844 608
rect 3942 607 3943 611
rect 3947 607 3948 611
rect 3942 606 3948 607
rect 3838 603 3844 604
rect 238 548 244 549
rect 110 545 116 546
rect 110 541 111 545
rect 115 541 116 545
rect 238 544 239 548
rect 243 544 244 548
rect 238 543 244 544
rect 414 548 420 549
rect 414 544 415 548
rect 419 544 420 548
rect 414 543 420 544
rect 606 548 612 549
rect 606 544 607 548
rect 611 544 612 548
rect 606 543 612 544
rect 798 548 804 549
rect 798 544 799 548
rect 803 544 804 548
rect 798 543 804 544
rect 990 548 996 549
rect 990 544 991 548
rect 995 544 996 548
rect 990 543 996 544
rect 1174 548 1180 549
rect 1174 544 1175 548
rect 1179 544 1180 548
rect 1174 543 1180 544
rect 1350 548 1356 549
rect 1350 544 1351 548
rect 1355 544 1356 548
rect 1350 543 1356 544
rect 1518 548 1524 549
rect 1518 544 1519 548
rect 1523 544 1524 548
rect 1518 543 1524 544
rect 1686 548 1692 549
rect 1686 544 1687 548
rect 1691 544 1692 548
rect 1686 543 1692 544
rect 1862 548 1868 549
rect 1862 544 1863 548
rect 1867 544 1868 548
rect 2190 548 2196 549
rect 1862 543 1868 544
rect 2006 545 2012 546
rect 110 540 116 541
rect 2006 541 2007 545
rect 2011 541 2012 545
rect 2006 540 2012 541
rect 2046 545 2052 546
rect 2046 541 2047 545
rect 2051 541 2052 545
rect 2190 544 2191 548
rect 2195 544 2196 548
rect 2190 543 2196 544
rect 2286 548 2292 549
rect 2286 544 2287 548
rect 2291 544 2292 548
rect 2286 543 2292 544
rect 2382 548 2388 549
rect 2382 544 2383 548
rect 2387 544 2388 548
rect 2382 543 2388 544
rect 2478 548 2484 549
rect 2478 544 2479 548
rect 2483 544 2484 548
rect 2478 543 2484 544
rect 2582 548 2588 549
rect 2582 544 2583 548
rect 2587 544 2588 548
rect 2582 543 2588 544
rect 2710 548 2716 549
rect 2710 544 2711 548
rect 2715 544 2716 548
rect 2710 543 2716 544
rect 2870 548 2876 549
rect 2870 544 2871 548
rect 2875 544 2876 548
rect 2870 543 2876 544
rect 3070 548 3076 549
rect 3070 544 3071 548
rect 3075 544 3076 548
rect 3070 543 3076 544
rect 3302 548 3308 549
rect 3302 544 3303 548
rect 3307 544 3308 548
rect 3302 543 3308 544
rect 3550 548 3556 549
rect 3550 544 3551 548
rect 3555 544 3556 548
rect 3550 543 3556 544
rect 3806 548 3812 549
rect 3806 544 3807 548
rect 3811 544 3812 548
rect 3806 543 3812 544
rect 3942 545 3948 546
rect 2046 540 2052 541
rect 3942 541 3943 545
rect 3947 541 3948 545
rect 3942 540 3948 541
rect 238 529 244 530
rect 110 528 116 529
rect 110 524 111 528
rect 115 524 116 528
rect 238 525 239 529
rect 243 525 244 529
rect 238 524 244 525
rect 414 529 420 530
rect 414 525 415 529
rect 419 525 420 529
rect 414 524 420 525
rect 606 529 612 530
rect 606 525 607 529
rect 611 525 612 529
rect 606 524 612 525
rect 798 529 804 530
rect 798 525 799 529
rect 803 525 804 529
rect 798 524 804 525
rect 990 529 996 530
rect 990 525 991 529
rect 995 525 996 529
rect 990 524 996 525
rect 1174 529 1180 530
rect 1174 525 1175 529
rect 1179 525 1180 529
rect 1174 524 1180 525
rect 1350 529 1356 530
rect 1350 525 1351 529
rect 1355 525 1356 529
rect 1350 524 1356 525
rect 1518 529 1524 530
rect 1518 525 1519 529
rect 1523 525 1524 529
rect 1518 524 1524 525
rect 1686 529 1692 530
rect 1686 525 1687 529
rect 1691 525 1692 529
rect 1686 524 1692 525
rect 1862 529 1868 530
rect 2190 529 2196 530
rect 1862 525 1863 529
rect 1867 525 1868 529
rect 1862 524 1868 525
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 110 523 116 524
rect 2006 523 2012 524
rect 2046 528 2052 529
rect 2046 524 2047 528
rect 2051 524 2052 528
rect 2190 525 2191 529
rect 2195 525 2196 529
rect 2190 524 2196 525
rect 2286 529 2292 530
rect 2286 525 2287 529
rect 2291 525 2292 529
rect 2286 524 2292 525
rect 2382 529 2388 530
rect 2382 525 2383 529
rect 2387 525 2388 529
rect 2382 524 2388 525
rect 2478 529 2484 530
rect 2478 525 2479 529
rect 2483 525 2484 529
rect 2478 524 2484 525
rect 2582 529 2588 530
rect 2582 525 2583 529
rect 2587 525 2588 529
rect 2582 524 2588 525
rect 2710 529 2716 530
rect 2710 525 2711 529
rect 2715 525 2716 529
rect 2710 524 2716 525
rect 2870 529 2876 530
rect 2870 525 2871 529
rect 2875 525 2876 529
rect 2870 524 2876 525
rect 3070 529 3076 530
rect 3070 525 3071 529
rect 3075 525 3076 529
rect 3070 524 3076 525
rect 3302 529 3308 530
rect 3302 525 3303 529
rect 3307 525 3308 529
rect 3302 524 3308 525
rect 3550 529 3556 530
rect 3550 525 3551 529
rect 3555 525 3556 529
rect 3550 524 3556 525
rect 3806 529 3812 530
rect 3806 525 3807 529
rect 3811 525 3812 529
rect 3806 524 3812 525
rect 3942 528 3948 529
rect 3942 524 3943 528
rect 3947 524 3948 528
rect 2046 523 2052 524
rect 3942 523 3948 524
rect 110 476 116 477
rect 2006 476 2012 477
rect 110 472 111 476
rect 115 472 116 476
rect 110 471 116 472
rect 134 475 140 476
rect 134 471 135 475
rect 139 471 140 475
rect 134 470 140 471
rect 286 475 292 476
rect 286 471 287 475
rect 291 471 292 475
rect 286 470 292 471
rect 462 475 468 476
rect 462 471 463 475
rect 467 471 468 475
rect 462 470 468 471
rect 638 475 644 476
rect 638 471 639 475
rect 643 471 644 475
rect 638 470 644 471
rect 806 475 812 476
rect 806 471 807 475
rect 811 471 812 475
rect 806 470 812 471
rect 966 475 972 476
rect 966 471 967 475
rect 971 471 972 475
rect 966 470 972 471
rect 1118 475 1124 476
rect 1118 471 1119 475
rect 1123 471 1124 475
rect 1118 470 1124 471
rect 1270 475 1276 476
rect 1270 471 1271 475
rect 1275 471 1276 475
rect 1270 470 1276 471
rect 1414 475 1420 476
rect 1414 471 1415 475
rect 1419 471 1420 475
rect 1414 470 1420 471
rect 1566 475 1572 476
rect 1566 471 1567 475
rect 1571 471 1572 475
rect 2006 472 2007 476
rect 2011 472 2012 476
rect 2006 471 2012 472
rect 2046 476 2052 477
rect 3942 476 3948 477
rect 2046 472 2047 476
rect 2051 472 2052 476
rect 2046 471 2052 472
rect 2430 475 2436 476
rect 2430 471 2431 475
rect 2435 471 2436 475
rect 1566 470 1572 471
rect 2430 470 2436 471
rect 2526 475 2532 476
rect 2526 471 2527 475
rect 2531 471 2532 475
rect 2526 470 2532 471
rect 2622 475 2628 476
rect 2622 471 2623 475
rect 2627 471 2628 475
rect 2622 470 2628 471
rect 2726 475 2732 476
rect 2726 471 2727 475
rect 2731 471 2732 475
rect 2726 470 2732 471
rect 2846 475 2852 476
rect 2846 471 2847 475
rect 2851 471 2852 475
rect 2846 470 2852 471
rect 2998 475 3004 476
rect 2998 471 2999 475
rect 3003 471 3004 475
rect 2998 470 3004 471
rect 3174 475 3180 476
rect 3174 471 3175 475
rect 3179 471 3180 475
rect 3174 470 3180 471
rect 3374 475 3380 476
rect 3374 471 3375 475
rect 3379 471 3380 475
rect 3374 470 3380 471
rect 3590 475 3596 476
rect 3590 471 3591 475
rect 3595 471 3596 475
rect 3590 470 3596 471
rect 3806 475 3812 476
rect 3806 471 3807 475
rect 3811 471 3812 475
rect 3942 472 3943 476
rect 3947 472 3948 476
rect 3942 471 3948 472
rect 3806 470 3812 471
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 2006 459 2012 460
rect 110 454 116 455
rect 134 456 140 457
rect 134 452 135 456
rect 139 452 140 456
rect 134 451 140 452
rect 286 456 292 457
rect 286 452 287 456
rect 291 452 292 456
rect 286 451 292 452
rect 462 456 468 457
rect 462 452 463 456
rect 467 452 468 456
rect 462 451 468 452
rect 638 456 644 457
rect 638 452 639 456
rect 643 452 644 456
rect 638 451 644 452
rect 806 456 812 457
rect 806 452 807 456
rect 811 452 812 456
rect 806 451 812 452
rect 966 456 972 457
rect 966 452 967 456
rect 971 452 972 456
rect 966 451 972 452
rect 1118 456 1124 457
rect 1118 452 1119 456
rect 1123 452 1124 456
rect 1118 451 1124 452
rect 1270 456 1276 457
rect 1270 452 1271 456
rect 1275 452 1276 456
rect 1270 451 1276 452
rect 1414 456 1420 457
rect 1414 452 1415 456
rect 1419 452 1420 456
rect 1414 451 1420 452
rect 1566 456 1572 457
rect 1566 452 1567 456
rect 1571 452 1572 456
rect 2006 455 2007 459
rect 2011 455 2012 459
rect 2006 454 2012 455
rect 2046 459 2052 460
rect 2046 455 2047 459
rect 2051 455 2052 459
rect 3942 459 3948 460
rect 2046 454 2052 455
rect 2430 456 2436 457
rect 1566 451 1572 452
rect 2430 452 2431 456
rect 2435 452 2436 456
rect 2430 451 2436 452
rect 2526 456 2532 457
rect 2526 452 2527 456
rect 2531 452 2532 456
rect 2526 451 2532 452
rect 2622 456 2628 457
rect 2622 452 2623 456
rect 2627 452 2628 456
rect 2622 451 2628 452
rect 2726 456 2732 457
rect 2726 452 2727 456
rect 2731 452 2732 456
rect 2726 451 2732 452
rect 2846 456 2852 457
rect 2846 452 2847 456
rect 2851 452 2852 456
rect 2846 451 2852 452
rect 2998 456 3004 457
rect 2998 452 2999 456
rect 3003 452 3004 456
rect 2998 451 3004 452
rect 3174 456 3180 457
rect 3174 452 3175 456
rect 3179 452 3180 456
rect 3174 451 3180 452
rect 3374 456 3380 457
rect 3374 452 3375 456
rect 3379 452 3380 456
rect 3374 451 3380 452
rect 3590 456 3596 457
rect 3590 452 3591 456
rect 3595 452 3596 456
rect 3590 451 3596 452
rect 3806 456 3812 457
rect 3806 452 3807 456
rect 3811 452 3812 456
rect 3942 455 3943 459
rect 3947 455 3948 459
rect 3942 454 3948 455
rect 3806 451 3812 452
rect 2430 396 2436 397
rect 2046 393 2052 394
rect 134 392 140 393
rect 110 389 116 390
rect 110 385 111 389
rect 115 385 116 389
rect 134 388 135 392
rect 139 388 140 392
rect 134 387 140 388
rect 278 392 284 393
rect 278 388 279 392
rect 283 388 284 392
rect 278 387 284 388
rect 438 392 444 393
rect 438 388 439 392
rect 443 388 444 392
rect 438 387 444 388
rect 582 392 588 393
rect 582 388 583 392
rect 587 388 588 392
rect 582 387 588 388
rect 718 392 724 393
rect 718 388 719 392
rect 723 388 724 392
rect 718 387 724 388
rect 846 392 852 393
rect 846 388 847 392
rect 851 388 852 392
rect 846 387 852 388
rect 966 392 972 393
rect 966 388 967 392
rect 971 388 972 392
rect 966 387 972 388
rect 1086 392 1092 393
rect 1086 388 1087 392
rect 1091 388 1092 392
rect 1086 387 1092 388
rect 1206 392 1212 393
rect 1206 388 1207 392
rect 1211 388 1212 392
rect 1206 387 1212 388
rect 1326 392 1332 393
rect 1326 388 1327 392
rect 1331 388 1332 392
rect 1326 387 1332 388
rect 2006 389 2012 390
rect 110 384 116 385
rect 2006 385 2007 389
rect 2011 385 2012 389
rect 2046 389 2047 393
rect 2051 389 2052 393
rect 2430 392 2431 396
rect 2435 392 2436 396
rect 2430 391 2436 392
rect 2526 396 2532 397
rect 2526 392 2527 396
rect 2531 392 2532 396
rect 2526 391 2532 392
rect 2622 396 2628 397
rect 2622 392 2623 396
rect 2627 392 2628 396
rect 2622 391 2628 392
rect 2718 396 2724 397
rect 2718 392 2719 396
rect 2723 392 2724 396
rect 2718 391 2724 392
rect 2814 396 2820 397
rect 2814 392 2815 396
rect 2819 392 2820 396
rect 2814 391 2820 392
rect 2926 396 2932 397
rect 2926 392 2927 396
rect 2931 392 2932 396
rect 2926 391 2932 392
rect 3062 396 3068 397
rect 3062 392 3063 396
rect 3067 392 3068 396
rect 3062 391 3068 392
rect 3222 396 3228 397
rect 3222 392 3223 396
rect 3227 392 3228 396
rect 3222 391 3228 392
rect 3398 396 3404 397
rect 3398 392 3399 396
rect 3403 392 3404 396
rect 3398 391 3404 392
rect 3590 396 3596 397
rect 3590 392 3591 396
rect 3595 392 3596 396
rect 3590 391 3596 392
rect 3782 396 3788 397
rect 3782 392 3783 396
rect 3787 392 3788 396
rect 3782 391 3788 392
rect 3942 393 3948 394
rect 2046 388 2052 389
rect 3942 389 3943 393
rect 3947 389 3948 393
rect 3942 388 3948 389
rect 2006 384 2012 385
rect 2430 377 2436 378
rect 2046 376 2052 377
rect 134 373 140 374
rect 110 372 116 373
rect 110 368 111 372
rect 115 368 116 372
rect 134 369 135 373
rect 139 369 140 373
rect 134 368 140 369
rect 278 373 284 374
rect 278 369 279 373
rect 283 369 284 373
rect 278 368 284 369
rect 438 373 444 374
rect 438 369 439 373
rect 443 369 444 373
rect 438 368 444 369
rect 582 373 588 374
rect 582 369 583 373
rect 587 369 588 373
rect 582 368 588 369
rect 718 373 724 374
rect 718 369 719 373
rect 723 369 724 373
rect 718 368 724 369
rect 846 373 852 374
rect 846 369 847 373
rect 851 369 852 373
rect 846 368 852 369
rect 966 373 972 374
rect 966 369 967 373
rect 971 369 972 373
rect 966 368 972 369
rect 1086 373 1092 374
rect 1086 369 1087 373
rect 1091 369 1092 373
rect 1086 368 1092 369
rect 1206 373 1212 374
rect 1206 369 1207 373
rect 1211 369 1212 373
rect 1206 368 1212 369
rect 1326 373 1332 374
rect 1326 369 1327 373
rect 1331 369 1332 373
rect 1326 368 1332 369
rect 2006 372 2012 373
rect 2006 368 2007 372
rect 2011 368 2012 372
rect 2046 372 2047 376
rect 2051 372 2052 376
rect 2430 373 2431 377
rect 2435 373 2436 377
rect 2430 372 2436 373
rect 2526 377 2532 378
rect 2526 373 2527 377
rect 2531 373 2532 377
rect 2526 372 2532 373
rect 2622 377 2628 378
rect 2622 373 2623 377
rect 2627 373 2628 377
rect 2622 372 2628 373
rect 2718 377 2724 378
rect 2718 373 2719 377
rect 2723 373 2724 377
rect 2718 372 2724 373
rect 2814 377 2820 378
rect 2814 373 2815 377
rect 2819 373 2820 377
rect 2814 372 2820 373
rect 2926 377 2932 378
rect 2926 373 2927 377
rect 2931 373 2932 377
rect 2926 372 2932 373
rect 3062 377 3068 378
rect 3062 373 3063 377
rect 3067 373 3068 377
rect 3062 372 3068 373
rect 3222 377 3228 378
rect 3222 373 3223 377
rect 3227 373 3228 377
rect 3222 372 3228 373
rect 3398 377 3404 378
rect 3398 373 3399 377
rect 3403 373 3404 377
rect 3398 372 3404 373
rect 3590 377 3596 378
rect 3590 373 3591 377
rect 3595 373 3596 377
rect 3590 372 3596 373
rect 3782 377 3788 378
rect 3782 373 3783 377
rect 3787 373 3788 377
rect 3782 372 3788 373
rect 3942 376 3948 377
rect 3942 372 3943 376
rect 3947 372 3948 376
rect 2046 371 2052 372
rect 3942 371 3948 372
rect 110 367 116 368
rect 2006 367 2012 368
rect 110 320 116 321
rect 2006 320 2012 321
rect 110 316 111 320
rect 115 316 116 320
rect 110 315 116 316
rect 142 319 148 320
rect 142 315 143 319
rect 147 315 148 319
rect 142 314 148 315
rect 318 319 324 320
rect 318 315 319 319
rect 323 315 324 319
rect 318 314 324 315
rect 478 319 484 320
rect 478 315 479 319
rect 483 315 484 319
rect 478 314 484 315
rect 630 319 636 320
rect 630 315 631 319
rect 635 315 636 319
rect 630 314 636 315
rect 774 319 780 320
rect 774 315 775 319
rect 779 315 780 319
rect 774 314 780 315
rect 902 319 908 320
rect 902 315 903 319
rect 907 315 908 319
rect 902 314 908 315
rect 1030 319 1036 320
rect 1030 315 1031 319
rect 1035 315 1036 319
rect 1030 314 1036 315
rect 1150 319 1156 320
rect 1150 315 1151 319
rect 1155 315 1156 319
rect 1150 314 1156 315
rect 1270 319 1276 320
rect 1270 315 1271 319
rect 1275 315 1276 319
rect 1270 314 1276 315
rect 1390 319 1396 320
rect 1390 315 1391 319
rect 1395 315 1396 319
rect 2006 316 2007 320
rect 2011 316 2012 320
rect 2006 315 2012 316
rect 2046 320 2052 321
rect 3942 320 3948 321
rect 2046 316 2047 320
rect 2051 316 2052 320
rect 2046 315 2052 316
rect 2190 319 2196 320
rect 2190 315 2191 319
rect 2195 315 2196 319
rect 1390 314 1396 315
rect 2190 314 2196 315
rect 2326 319 2332 320
rect 2326 315 2327 319
rect 2331 315 2332 319
rect 2326 314 2332 315
rect 2470 319 2476 320
rect 2470 315 2471 319
rect 2475 315 2476 319
rect 2470 314 2476 315
rect 2622 319 2628 320
rect 2622 315 2623 319
rect 2627 315 2628 319
rect 2622 314 2628 315
rect 2782 319 2788 320
rect 2782 315 2783 319
rect 2787 315 2788 319
rect 2782 314 2788 315
rect 2950 319 2956 320
rect 2950 315 2951 319
rect 2955 315 2956 319
rect 2950 314 2956 315
rect 3118 319 3124 320
rect 3118 315 3119 319
rect 3123 315 3124 319
rect 3118 314 3124 315
rect 3294 319 3300 320
rect 3294 315 3295 319
rect 3299 315 3300 319
rect 3294 314 3300 315
rect 3470 319 3476 320
rect 3470 315 3471 319
rect 3475 315 3476 319
rect 3470 314 3476 315
rect 3654 319 3660 320
rect 3654 315 3655 319
rect 3659 315 3660 319
rect 3654 314 3660 315
rect 3838 319 3844 320
rect 3838 315 3839 319
rect 3843 315 3844 319
rect 3942 316 3943 320
rect 3947 316 3948 320
rect 3942 315 3948 316
rect 3838 314 3844 315
rect 110 303 116 304
rect 110 299 111 303
rect 115 299 116 303
rect 2006 303 2012 304
rect 110 298 116 299
rect 142 300 148 301
rect 142 296 143 300
rect 147 296 148 300
rect 142 295 148 296
rect 318 300 324 301
rect 318 296 319 300
rect 323 296 324 300
rect 318 295 324 296
rect 478 300 484 301
rect 478 296 479 300
rect 483 296 484 300
rect 478 295 484 296
rect 630 300 636 301
rect 630 296 631 300
rect 635 296 636 300
rect 630 295 636 296
rect 774 300 780 301
rect 774 296 775 300
rect 779 296 780 300
rect 774 295 780 296
rect 902 300 908 301
rect 902 296 903 300
rect 907 296 908 300
rect 902 295 908 296
rect 1030 300 1036 301
rect 1030 296 1031 300
rect 1035 296 1036 300
rect 1030 295 1036 296
rect 1150 300 1156 301
rect 1150 296 1151 300
rect 1155 296 1156 300
rect 1150 295 1156 296
rect 1270 300 1276 301
rect 1270 296 1271 300
rect 1275 296 1276 300
rect 1270 295 1276 296
rect 1390 300 1396 301
rect 1390 296 1391 300
rect 1395 296 1396 300
rect 2006 299 2007 303
rect 2011 299 2012 303
rect 2006 298 2012 299
rect 2046 303 2052 304
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 3942 303 3948 304
rect 2046 298 2052 299
rect 2190 300 2196 301
rect 1390 295 1396 296
rect 2190 296 2191 300
rect 2195 296 2196 300
rect 2190 295 2196 296
rect 2326 300 2332 301
rect 2326 296 2327 300
rect 2331 296 2332 300
rect 2326 295 2332 296
rect 2470 300 2476 301
rect 2470 296 2471 300
rect 2475 296 2476 300
rect 2470 295 2476 296
rect 2622 300 2628 301
rect 2622 296 2623 300
rect 2627 296 2628 300
rect 2622 295 2628 296
rect 2782 300 2788 301
rect 2782 296 2783 300
rect 2787 296 2788 300
rect 2782 295 2788 296
rect 2950 300 2956 301
rect 2950 296 2951 300
rect 2955 296 2956 300
rect 2950 295 2956 296
rect 3118 300 3124 301
rect 3118 296 3119 300
rect 3123 296 3124 300
rect 3118 295 3124 296
rect 3294 300 3300 301
rect 3294 296 3295 300
rect 3299 296 3300 300
rect 3294 295 3300 296
rect 3470 300 3476 301
rect 3470 296 3471 300
rect 3475 296 3476 300
rect 3470 295 3476 296
rect 3654 300 3660 301
rect 3654 296 3655 300
rect 3659 296 3660 300
rect 3654 295 3660 296
rect 3838 300 3844 301
rect 3838 296 3839 300
rect 3843 296 3844 300
rect 3942 299 3943 303
rect 3947 299 3948 303
rect 3942 298 3948 299
rect 3838 295 3844 296
rect 2070 240 2076 241
rect 2046 237 2052 238
rect 222 236 228 237
rect 110 233 116 234
rect 110 229 111 233
rect 115 229 116 233
rect 222 232 223 236
rect 227 232 228 236
rect 222 231 228 232
rect 390 236 396 237
rect 390 232 391 236
rect 395 232 396 236
rect 390 231 396 232
rect 558 236 564 237
rect 558 232 559 236
rect 563 232 564 236
rect 558 231 564 232
rect 734 236 740 237
rect 734 232 735 236
rect 739 232 740 236
rect 734 231 740 232
rect 902 236 908 237
rect 902 232 903 236
rect 907 232 908 236
rect 902 231 908 232
rect 1062 236 1068 237
rect 1062 232 1063 236
rect 1067 232 1068 236
rect 1062 231 1068 232
rect 1214 236 1220 237
rect 1214 232 1215 236
rect 1219 232 1220 236
rect 1214 231 1220 232
rect 1358 236 1364 237
rect 1358 232 1359 236
rect 1363 232 1364 236
rect 1358 231 1364 232
rect 1510 236 1516 237
rect 1510 232 1511 236
rect 1515 232 1516 236
rect 1510 231 1516 232
rect 1662 236 1668 237
rect 1662 232 1663 236
rect 1667 232 1668 236
rect 1662 231 1668 232
rect 2006 233 2012 234
rect 110 228 116 229
rect 2006 229 2007 233
rect 2011 229 2012 233
rect 2046 233 2047 237
rect 2051 233 2052 237
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2214 240 2220 241
rect 2214 236 2215 240
rect 2219 236 2220 240
rect 2214 235 2220 236
rect 2398 240 2404 241
rect 2398 236 2399 240
rect 2403 236 2404 240
rect 2398 235 2404 236
rect 2590 240 2596 241
rect 2590 236 2591 240
rect 2595 236 2596 240
rect 2590 235 2596 236
rect 2790 240 2796 241
rect 2790 236 2791 240
rect 2795 236 2796 240
rect 2790 235 2796 236
rect 2982 240 2988 241
rect 2982 236 2983 240
rect 2987 236 2988 240
rect 2982 235 2988 236
rect 3166 240 3172 241
rect 3166 236 3167 240
rect 3171 236 3172 240
rect 3166 235 3172 236
rect 3342 240 3348 241
rect 3342 236 3343 240
rect 3347 236 3348 240
rect 3342 235 3348 236
rect 3510 240 3516 241
rect 3510 236 3511 240
rect 3515 236 3516 240
rect 3510 235 3516 236
rect 3686 240 3692 241
rect 3686 236 3687 240
rect 3691 236 3692 240
rect 3686 235 3692 236
rect 3838 240 3844 241
rect 3838 236 3839 240
rect 3843 236 3844 240
rect 3838 235 3844 236
rect 3942 237 3948 238
rect 2046 232 2052 233
rect 3942 233 3943 237
rect 3947 233 3948 237
rect 3942 232 3948 233
rect 2006 228 2012 229
rect 2070 221 2076 222
rect 2046 220 2052 221
rect 222 217 228 218
rect 110 216 116 217
rect 110 212 111 216
rect 115 212 116 216
rect 222 213 223 217
rect 227 213 228 217
rect 222 212 228 213
rect 390 217 396 218
rect 390 213 391 217
rect 395 213 396 217
rect 390 212 396 213
rect 558 217 564 218
rect 558 213 559 217
rect 563 213 564 217
rect 558 212 564 213
rect 734 217 740 218
rect 734 213 735 217
rect 739 213 740 217
rect 734 212 740 213
rect 902 217 908 218
rect 902 213 903 217
rect 907 213 908 217
rect 902 212 908 213
rect 1062 217 1068 218
rect 1062 213 1063 217
rect 1067 213 1068 217
rect 1062 212 1068 213
rect 1214 217 1220 218
rect 1214 213 1215 217
rect 1219 213 1220 217
rect 1214 212 1220 213
rect 1358 217 1364 218
rect 1358 213 1359 217
rect 1363 213 1364 217
rect 1358 212 1364 213
rect 1510 217 1516 218
rect 1510 213 1511 217
rect 1515 213 1516 217
rect 1510 212 1516 213
rect 1662 217 1668 218
rect 1662 213 1663 217
rect 1667 213 1668 217
rect 1662 212 1668 213
rect 2006 216 2012 217
rect 2006 212 2007 216
rect 2011 212 2012 216
rect 2046 216 2047 220
rect 2051 216 2052 220
rect 2070 217 2071 221
rect 2075 217 2076 221
rect 2070 216 2076 217
rect 2214 221 2220 222
rect 2214 217 2215 221
rect 2219 217 2220 221
rect 2214 216 2220 217
rect 2398 221 2404 222
rect 2398 217 2399 221
rect 2403 217 2404 221
rect 2398 216 2404 217
rect 2590 221 2596 222
rect 2590 217 2591 221
rect 2595 217 2596 221
rect 2590 216 2596 217
rect 2790 221 2796 222
rect 2790 217 2791 221
rect 2795 217 2796 221
rect 2790 216 2796 217
rect 2982 221 2988 222
rect 2982 217 2983 221
rect 2987 217 2988 221
rect 2982 216 2988 217
rect 3166 221 3172 222
rect 3166 217 3167 221
rect 3171 217 3172 221
rect 3166 216 3172 217
rect 3342 221 3348 222
rect 3342 217 3343 221
rect 3347 217 3348 221
rect 3342 216 3348 217
rect 3510 221 3516 222
rect 3510 217 3511 221
rect 3515 217 3516 221
rect 3510 216 3516 217
rect 3686 221 3692 222
rect 3686 217 3687 221
rect 3691 217 3692 221
rect 3686 216 3692 217
rect 3838 221 3844 222
rect 3838 217 3839 221
rect 3843 217 3844 221
rect 3838 216 3844 217
rect 3942 220 3948 221
rect 3942 216 3943 220
rect 3947 216 3948 220
rect 2046 215 2052 216
rect 3942 215 3948 216
rect 110 211 116 212
rect 2006 211 2012 212
rect 2046 144 2052 145
rect 3942 144 3948 145
rect 2046 140 2047 144
rect 2051 140 2052 144
rect 2046 139 2052 140
rect 2070 143 2076 144
rect 2070 139 2071 143
rect 2075 139 2076 143
rect 2070 138 2076 139
rect 2190 143 2196 144
rect 2190 139 2191 143
rect 2195 139 2196 143
rect 2190 138 2196 139
rect 2342 143 2348 144
rect 2342 139 2343 143
rect 2347 139 2348 143
rect 2342 138 2348 139
rect 2494 143 2500 144
rect 2494 139 2495 143
rect 2499 139 2500 143
rect 2494 138 2500 139
rect 2646 143 2652 144
rect 2646 139 2647 143
rect 2651 139 2652 143
rect 2646 138 2652 139
rect 2798 143 2804 144
rect 2798 139 2799 143
rect 2803 139 2804 143
rect 2798 138 2804 139
rect 2942 143 2948 144
rect 2942 139 2943 143
rect 2947 139 2948 143
rect 2942 138 2948 139
rect 3070 143 3076 144
rect 3070 139 3071 143
rect 3075 139 3076 143
rect 3070 138 3076 139
rect 3190 143 3196 144
rect 3190 139 3191 143
rect 3195 139 3196 143
rect 3190 138 3196 139
rect 3310 143 3316 144
rect 3310 139 3311 143
rect 3315 139 3316 143
rect 3310 138 3316 139
rect 3422 143 3428 144
rect 3422 139 3423 143
rect 3427 139 3428 143
rect 3422 138 3428 139
rect 3526 143 3532 144
rect 3526 139 3527 143
rect 3531 139 3532 143
rect 3526 138 3532 139
rect 3638 143 3644 144
rect 3638 139 3639 143
rect 3643 139 3644 143
rect 3638 138 3644 139
rect 3742 143 3748 144
rect 3742 139 3743 143
rect 3747 139 3748 143
rect 3742 138 3748 139
rect 3838 143 3844 144
rect 3838 139 3839 143
rect 3843 139 3844 143
rect 3942 140 3943 144
rect 3947 140 3948 144
rect 3942 139 3948 140
rect 3838 138 3844 139
rect 110 132 116 133
rect 2006 132 2012 133
rect 110 128 111 132
rect 115 128 116 132
rect 110 127 116 128
rect 150 131 156 132
rect 150 127 151 131
rect 155 127 156 131
rect 150 126 156 127
rect 246 131 252 132
rect 246 127 247 131
rect 251 127 252 131
rect 246 126 252 127
rect 342 131 348 132
rect 342 127 343 131
rect 347 127 348 131
rect 342 126 348 127
rect 438 131 444 132
rect 438 127 439 131
rect 443 127 444 131
rect 438 126 444 127
rect 534 131 540 132
rect 534 127 535 131
rect 539 127 540 131
rect 534 126 540 127
rect 630 131 636 132
rect 630 127 631 131
rect 635 127 636 131
rect 630 126 636 127
rect 726 131 732 132
rect 726 127 727 131
rect 731 127 732 131
rect 726 126 732 127
rect 822 131 828 132
rect 822 127 823 131
rect 827 127 828 131
rect 822 126 828 127
rect 918 131 924 132
rect 918 127 919 131
rect 923 127 924 131
rect 918 126 924 127
rect 1014 131 1020 132
rect 1014 127 1015 131
rect 1019 127 1020 131
rect 1014 126 1020 127
rect 1110 131 1116 132
rect 1110 127 1111 131
rect 1115 127 1116 131
rect 1110 126 1116 127
rect 1206 131 1212 132
rect 1206 127 1207 131
rect 1211 127 1212 131
rect 1206 126 1212 127
rect 1302 131 1308 132
rect 1302 127 1303 131
rect 1307 127 1308 131
rect 1302 126 1308 127
rect 1406 131 1412 132
rect 1406 127 1407 131
rect 1411 127 1412 131
rect 1406 126 1412 127
rect 1510 131 1516 132
rect 1510 127 1511 131
rect 1515 127 1516 131
rect 1510 126 1516 127
rect 1614 131 1620 132
rect 1614 127 1615 131
rect 1619 127 1620 131
rect 1614 126 1620 127
rect 1710 131 1716 132
rect 1710 127 1711 131
rect 1715 127 1716 131
rect 1710 126 1716 127
rect 1806 131 1812 132
rect 1806 127 1807 131
rect 1811 127 1812 131
rect 1806 126 1812 127
rect 1902 131 1908 132
rect 1902 127 1903 131
rect 1907 127 1908 131
rect 2006 128 2007 132
rect 2011 128 2012 132
rect 2006 127 2012 128
rect 2046 127 2052 128
rect 1902 126 1908 127
rect 2046 123 2047 127
rect 2051 123 2052 127
rect 3942 127 3948 128
rect 2046 122 2052 123
rect 2070 124 2076 125
rect 2070 120 2071 124
rect 2075 120 2076 124
rect 2070 119 2076 120
rect 2190 124 2196 125
rect 2190 120 2191 124
rect 2195 120 2196 124
rect 2190 119 2196 120
rect 2342 124 2348 125
rect 2342 120 2343 124
rect 2347 120 2348 124
rect 2342 119 2348 120
rect 2494 124 2500 125
rect 2494 120 2495 124
rect 2499 120 2500 124
rect 2494 119 2500 120
rect 2646 124 2652 125
rect 2646 120 2647 124
rect 2651 120 2652 124
rect 2646 119 2652 120
rect 2798 124 2804 125
rect 2798 120 2799 124
rect 2803 120 2804 124
rect 2798 119 2804 120
rect 2942 124 2948 125
rect 2942 120 2943 124
rect 2947 120 2948 124
rect 2942 119 2948 120
rect 3070 124 3076 125
rect 3070 120 3071 124
rect 3075 120 3076 124
rect 3070 119 3076 120
rect 3190 124 3196 125
rect 3190 120 3191 124
rect 3195 120 3196 124
rect 3190 119 3196 120
rect 3310 124 3316 125
rect 3310 120 3311 124
rect 3315 120 3316 124
rect 3310 119 3316 120
rect 3422 124 3428 125
rect 3422 120 3423 124
rect 3427 120 3428 124
rect 3422 119 3428 120
rect 3526 124 3532 125
rect 3526 120 3527 124
rect 3531 120 3532 124
rect 3526 119 3532 120
rect 3638 124 3644 125
rect 3638 120 3639 124
rect 3643 120 3644 124
rect 3638 119 3644 120
rect 3742 124 3748 125
rect 3742 120 3743 124
rect 3747 120 3748 124
rect 3742 119 3748 120
rect 3838 124 3844 125
rect 3838 120 3839 124
rect 3843 120 3844 124
rect 3942 123 3943 127
rect 3947 123 3948 127
rect 3942 122 3948 123
rect 3838 119 3844 120
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 2006 115 2012 116
rect 110 110 116 111
rect 150 112 156 113
rect 150 108 151 112
rect 155 108 156 112
rect 150 107 156 108
rect 246 112 252 113
rect 246 108 247 112
rect 251 108 252 112
rect 246 107 252 108
rect 342 112 348 113
rect 342 108 343 112
rect 347 108 348 112
rect 342 107 348 108
rect 438 112 444 113
rect 438 108 439 112
rect 443 108 444 112
rect 438 107 444 108
rect 534 112 540 113
rect 534 108 535 112
rect 539 108 540 112
rect 534 107 540 108
rect 630 112 636 113
rect 630 108 631 112
rect 635 108 636 112
rect 630 107 636 108
rect 726 112 732 113
rect 726 108 727 112
rect 731 108 732 112
rect 726 107 732 108
rect 822 112 828 113
rect 822 108 823 112
rect 827 108 828 112
rect 822 107 828 108
rect 918 112 924 113
rect 918 108 919 112
rect 923 108 924 112
rect 918 107 924 108
rect 1014 112 1020 113
rect 1014 108 1015 112
rect 1019 108 1020 112
rect 1014 107 1020 108
rect 1110 112 1116 113
rect 1110 108 1111 112
rect 1115 108 1116 112
rect 1110 107 1116 108
rect 1206 112 1212 113
rect 1206 108 1207 112
rect 1211 108 1212 112
rect 1206 107 1212 108
rect 1302 112 1308 113
rect 1302 108 1303 112
rect 1307 108 1308 112
rect 1302 107 1308 108
rect 1406 112 1412 113
rect 1406 108 1407 112
rect 1411 108 1412 112
rect 1406 107 1412 108
rect 1510 112 1516 113
rect 1510 108 1511 112
rect 1515 108 1516 112
rect 1510 107 1516 108
rect 1614 112 1620 113
rect 1614 108 1615 112
rect 1619 108 1620 112
rect 1614 107 1620 108
rect 1710 112 1716 113
rect 1710 108 1711 112
rect 1715 108 1716 112
rect 1710 107 1716 108
rect 1806 112 1812 113
rect 1806 108 1807 112
rect 1811 108 1812 112
rect 1806 107 1812 108
rect 1902 112 1908 113
rect 1902 108 1903 112
rect 1907 108 1908 112
rect 2006 111 2007 115
rect 2011 111 2012 115
rect 2006 110 2012 111
rect 1902 107 1908 108
<< m3c >>
rect 2047 3985 2051 3989
rect 2071 3988 2075 3992
rect 2327 3988 2331 3992
rect 2591 3988 2595 3992
rect 2839 3988 2843 3992
rect 3087 3988 3091 3992
rect 3343 3988 3347 3992
rect 3943 3985 3947 3989
rect 111 3965 115 3969
rect 311 3968 315 3972
rect 511 3968 515 3972
rect 703 3968 707 3972
rect 887 3968 891 3972
rect 1063 3968 1067 3972
rect 1231 3968 1235 3972
rect 1383 3968 1387 3972
rect 1519 3968 1523 3972
rect 1655 3968 1659 3972
rect 1791 3968 1795 3972
rect 1903 3968 1907 3972
rect 2007 3965 2011 3969
rect 2047 3968 2051 3972
rect 2071 3969 2075 3973
rect 2327 3969 2331 3973
rect 2591 3969 2595 3973
rect 2839 3969 2843 3973
rect 3087 3969 3091 3973
rect 3343 3969 3347 3973
rect 3943 3968 3947 3972
rect 111 3948 115 3952
rect 311 3949 315 3953
rect 511 3949 515 3953
rect 703 3949 707 3953
rect 887 3949 891 3953
rect 1063 3949 1067 3953
rect 1231 3949 1235 3953
rect 1383 3949 1387 3953
rect 1519 3949 1523 3953
rect 1655 3949 1659 3953
rect 1791 3949 1795 3953
rect 1903 3949 1907 3953
rect 2007 3948 2011 3952
rect 2047 3916 2051 3920
rect 2127 3915 2131 3919
rect 2271 3915 2275 3919
rect 2439 3915 2443 3919
rect 2615 3915 2619 3919
rect 2799 3915 2803 3919
rect 2983 3915 2987 3919
rect 3175 3915 3179 3919
rect 3367 3915 3371 3919
rect 3559 3915 3563 3919
rect 3943 3916 3947 3920
rect 111 3896 115 3900
rect 279 3895 283 3899
rect 415 3895 419 3899
rect 567 3895 571 3899
rect 735 3895 739 3899
rect 911 3895 915 3899
rect 1095 3895 1099 3899
rect 1287 3895 1291 3899
rect 1479 3895 1483 3899
rect 1679 3895 1683 3899
rect 2007 3896 2011 3900
rect 2047 3899 2051 3903
rect 2127 3896 2131 3900
rect 2271 3896 2275 3900
rect 2439 3896 2443 3900
rect 2615 3896 2619 3900
rect 2799 3896 2803 3900
rect 2983 3896 2987 3900
rect 3175 3896 3179 3900
rect 3367 3896 3371 3900
rect 3559 3896 3563 3900
rect 3943 3899 3947 3903
rect 111 3879 115 3883
rect 279 3876 283 3880
rect 415 3876 419 3880
rect 567 3876 571 3880
rect 735 3876 739 3880
rect 911 3876 915 3880
rect 1095 3876 1099 3880
rect 1287 3876 1291 3880
rect 1479 3876 1483 3880
rect 1679 3876 1683 3880
rect 2007 3879 2011 3883
rect 2047 3833 2051 3837
rect 2263 3836 2267 3840
rect 2375 3836 2379 3840
rect 2495 3836 2499 3840
rect 2631 3836 2635 3840
rect 2775 3836 2779 3840
rect 2919 3836 2923 3840
rect 3063 3836 3067 3840
rect 3207 3836 3211 3840
rect 3343 3836 3347 3840
rect 3471 3836 3475 3840
rect 3599 3836 3603 3840
rect 3727 3836 3731 3840
rect 3839 3836 3843 3840
rect 3943 3833 3947 3837
rect 2047 3816 2051 3820
rect 2263 3817 2267 3821
rect 2375 3817 2379 3821
rect 2495 3817 2499 3821
rect 2631 3817 2635 3821
rect 2775 3817 2779 3821
rect 2919 3817 2923 3821
rect 3063 3817 3067 3821
rect 3207 3817 3211 3821
rect 3343 3817 3347 3821
rect 3471 3817 3475 3821
rect 3599 3817 3603 3821
rect 3727 3817 3731 3821
rect 3839 3817 3843 3821
rect 3943 3816 3947 3820
rect 111 3805 115 3809
rect 231 3808 235 3812
rect 335 3808 339 3812
rect 439 3808 443 3812
rect 535 3808 539 3812
rect 631 3808 635 3812
rect 727 3808 731 3812
rect 831 3808 835 3812
rect 935 3808 939 3812
rect 1039 3808 1043 3812
rect 1151 3808 1155 3812
rect 1263 3808 1267 3812
rect 1383 3808 1387 3812
rect 1503 3808 1507 3812
rect 1631 3808 1635 3812
rect 2007 3805 2011 3809
rect 111 3788 115 3792
rect 231 3789 235 3793
rect 335 3789 339 3793
rect 439 3789 443 3793
rect 535 3789 539 3793
rect 631 3789 635 3793
rect 727 3789 731 3793
rect 831 3789 835 3793
rect 935 3789 939 3793
rect 1039 3789 1043 3793
rect 1151 3789 1155 3793
rect 1263 3789 1267 3793
rect 1383 3789 1387 3793
rect 1503 3789 1507 3793
rect 1631 3789 1635 3793
rect 2007 3788 2011 3792
rect 2047 3748 2051 3752
rect 2071 3747 2075 3751
rect 2183 3747 2187 3751
rect 2327 3747 2331 3751
rect 2479 3747 2483 3751
rect 2639 3747 2643 3751
rect 2807 3747 2811 3751
rect 2983 3747 2987 3751
rect 3159 3747 3163 3751
rect 3335 3747 3339 3751
rect 3511 3747 3515 3751
rect 3687 3747 3691 3751
rect 3839 3747 3843 3751
rect 3943 3748 3947 3752
rect 111 3736 115 3740
rect 159 3735 163 3739
rect 351 3735 355 3739
rect 551 3735 555 3739
rect 751 3735 755 3739
rect 959 3735 963 3739
rect 1167 3735 1171 3739
rect 1383 3735 1387 3739
rect 1607 3735 1611 3739
rect 2007 3736 2011 3740
rect 2047 3731 2051 3735
rect 2071 3728 2075 3732
rect 2183 3728 2187 3732
rect 2327 3728 2331 3732
rect 2479 3728 2483 3732
rect 2639 3728 2643 3732
rect 2807 3728 2811 3732
rect 2983 3728 2987 3732
rect 3159 3728 3163 3732
rect 3335 3728 3339 3732
rect 3511 3728 3515 3732
rect 3687 3728 3691 3732
rect 3839 3728 3843 3732
rect 3943 3731 3947 3735
rect 111 3719 115 3723
rect 159 3716 163 3720
rect 351 3716 355 3720
rect 551 3716 555 3720
rect 751 3716 755 3720
rect 959 3716 963 3720
rect 1167 3716 1171 3720
rect 1383 3716 1387 3720
rect 1607 3716 1611 3720
rect 2007 3719 2011 3723
rect 2047 3653 2051 3657
rect 2071 3656 2075 3660
rect 2199 3656 2203 3660
rect 2367 3656 2371 3660
rect 2551 3656 2555 3660
rect 2735 3656 2739 3660
rect 2927 3656 2931 3660
rect 3111 3656 3115 3660
rect 3295 3656 3299 3660
rect 3479 3656 3483 3660
rect 3671 3656 3675 3660
rect 3839 3656 3843 3660
rect 111 3645 115 3649
rect 151 3648 155 3652
rect 383 3648 387 3652
rect 615 3648 619 3652
rect 839 3648 843 3652
rect 1055 3648 1059 3652
rect 1263 3648 1267 3652
rect 1479 3648 1483 3652
rect 3943 3653 3947 3657
rect 1695 3648 1699 3652
rect 2007 3645 2011 3649
rect 2047 3636 2051 3640
rect 2071 3637 2075 3641
rect 2199 3637 2203 3641
rect 2367 3637 2371 3641
rect 2551 3637 2555 3641
rect 2735 3637 2739 3641
rect 2927 3637 2931 3641
rect 3111 3637 3115 3641
rect 3295 3637 3299 3641
rect 3479 3637 3483 3641
rect 3671 3637 3675 3641
rect 3839 3637 3843 3641
rect 3943 3636 3947 3640
rect 111 3628 115 3632
rect 151 3629 155 3633
rect 383 3629 387 3633
rect 615 3629 619 3633
rect 839 3629 843 3633
rect 1055 3629 1059 3633
rect 1263 3629 1267 3633
rect 1479 3629 1483 3633
rect 1695 3629 1699 3633
rect 2007 3628 2011 3632
rect 2047 3580 2051 3584
rect 2103 3579 2107 3583
rect 2279 3579 2283 3583
rect 2471 3579 2475 3583
rect 2671 3579 2675 3583
rect 2871 3579 2875 3583
rect 3063 3579 3067 3583
rect 3255 3579 3259 3583
rect 3447 3579 3451 3583
rect 3639 3579 3643 3583
rect 3839 3579 3843 3583
rect 3943 3580 3947 3584
rect 111 3572 115 3576
rect 167 3571 171 3575
rect 359 3571 363 3575
rect 559 3571 563 3575
rect 775 3571 779 3575
rect 991 3571 995 3575
rect 1215 3571 1219 3575
rect 1447 3571 1451 3575
rect 1687 3571 1691 3575
rect 2007 3572 2011 3576
rect 2047 3563 2051 3567
rect 2103 3560 2107 3564
rect 111 3555 115 3559
rect 2279 3560 2283 3564
rect 2471 3560 2475 3564
rect 2671 3560 2675 3564
rect 2871 3560 2875 3564
rect 3063 3560 3067 3564
rect 3255 3560 3259 3564
rect 3447 3560 3451 3564
rect 3639 3560 3643 3564
rect 3839 3560 3843 3564
rect 3943 3563 3947 3567
rect 167 3552 171 3556
rect 359 3552 363 3556
rect 559 3552 563 3556
rect 775 3552 779 3556
rect 991 3552 995 3556
rect 1215 3552 1219 3556
rect 1447 3552 1451 3556
rect 1687 3552 1691 3556
rect 2007 3555 2011 3559
rect 2047 3493 2051 3497
rect 2327 3496 2331 3500
rect 2447 3496 2451 3500
rect 2583 3496 2587 3500
rect 2735 3496 2739 3500
rect 2911 3496 2915 3500
rect 3111 3496 3115 3500
rect 3335 3496 3339 3500
rect 3567 3496 3571 3500
rect 3807 3496 3811 3500
rect 3943 3493 3947 3497
rect 111 3481 115 3485
rect 295 3484 299 3488
rect 431 3484 435 3488
rect 583 3484 587 3488
rect 743 3484 747 3488
rect 911 3484 915 3488
rect 1079 3484 1083 3488
rect 1247 3484 1251 3488
rect 1423 3484 1427 3488
rect 1599 3484 1603 3488
rect 1775 3484 1779 3488
rect 2007 3481 2011 3485
rect 2047 3476 2051 3480
rect 2327 3477 2331 3481
rect 2447 3477 2451 3481
rect 2583 3477 2587 3481
rect 2735 3477 2739 3481
rect 2911 3477 2915 3481
rect 3111 3477 3115 3481
rect 3335 3477 3339 3481
rect 3567 3477 3571 3481
rect 3807 3477 3811 3481
rect 3943 3476 3947 3480
rect 111 3464 115 3468
rect 295 3465 299 3469
rect 431 3465 435 3469
rect 583 3465 587 3469
rect 743 3465 747 3469
rect 911 3465 915 3469
rect 1079 3465 1083 3469
rect 1247 3465 1251 3469
rect 1423 3465 1427 3469
rect 1599 3465 1603 3469
rect 1775 3465 1779 3469
rect 2007 3464 2011 3468
rect 2047 3424 2051 3428
rect 2447 3423 2451 3427
rect 2551 3423 2555 3427
rect 2663 3423 2667 3427
rect 2775 3423 2779 3427
rect 2903 3423 2907 3427
rect 3047 3423 3051 3427
rect 3207 3423 3211 3427
rect 3383 3423 3387 3427
rect 3567 3423 3571 3427
rect 3751 3423 3755 3427
rect 3943 3424 3947 3428
rect 2047 3407 2051 3411
rect 2447 3404 2451 3408
rect 2551 3404 2555 3408
rect 2663 3404 2667 3408
rect 2775 3404 2779 3408
rect 2903 3404 2907 3408
rect 3047 3404 3051 3408
rect 3207 3404 3211 3408
rect 3383 3404 3387 3408
rect 3567 3404 3571 3408
rect 3751 3404 3755 3408
rect 3943 3407 3947 3411
rect 111 3392 115 3396
rect 495 3391 499 3395
rect 647 3391 651 3395
rect 799 3391 803 3395
rect 959 3391 963 3395
rect 1127 3391 1131 3395
rect 1295 3391 1299 3395
rect 1463 3391 1467 3395
rect 1639 3391 1643 3395
rect 1815 3391 1819 3395
rect 2007 3392 2011 3396
rect 111 3375 115 3379
rect 495 3372 499 3376
rect 647 3372 651 3376
rect 799 3372 803 3376
rect 959 3372 963 3376
rect 1127 3372 1131 3376
rect 1295 3372 1299 3376
rect 1463 3372 1467 3376
rect 1639 3372 1643 3376
rect 1815 3372 1819 3376
rect 2007 3375 2011 3379
rect 2047 3329 2051 3333
rect 2567 3332 2571 3336
rect 2719 3332 2723 3336
rect 2871 3332 2875 3336
rect 3023 3332 3027 3336
rect 3175 3332 3179 3336
rect 3327 3332 3331 3336
rect 3479 3332 3483 3336
rect 3631 3332 3635 3336
rect 3783 3332 3787 3336
rect 3943 3329 3947 3333
rect 2047 3312 2051 3316
rect 2567 3313 2571 3317
rect 2719 3313 2723 3317
rect 2871 3313 2875 3317
rect 3023 3313 3027 3317
rect 3175 3313 3179 3317
rect 3327 3313 3331 3317
rect 3479 3313 3483 3317
rect 3631 3313 3635 3317
rect 3783 3313 3787 3317
rect 3943 3312 3947 3316
rect 111 3297 115 3301
rect 135 3300 139 3304
rect 295 3300 299 3304
rect 479 3300 483 3304
rect 671 3300 675 3304
rect 863 3300 867 3304
rect 1055 3300 1059 3304
rect 1247 3300 1251 3304
rect 1439 3300 1443 3304
rect 1631 3300 1635 3304
rect 1823 3300 1827 3304
rect 2007 3297 2011 3301
rect 111 3280 115 3284
rect 135 3281 139 3285
rect 295 3281 299 3285
rect 479 3281 483 3285
rect 671 3281 675 3285
rect 863 3281 867 3285
rect 1055 3281 1059 3285
rect 1247 3281 1251 3285
rect 1439 3281 1443 3285
rect 1631 3281 1635 3285
rect 1823 3281 1827 3285
rect 2007 3280 2011 3284
rect 2047 3256 2051 3260
rect 2415 3255 2419 3259
rect 2551 3255 2555 3259
rect 2687 3255 2691 3259
rect 2831 3255 2835 3259
rect 2975 3255 2979 3259
rect 3119 3255 3123 3259
rect 3255 3255 3259 3259
rect 3383 3255 3387 3259
rect 3503 3255 3507 3259
rect 3623 3255 3627 3259
rect 3743 3255 3747 3259
rect 3839 3255 3843 3259
rect 3943 3256 3947 3260
rect 2047 3239 2051 3243
rect 2415 3236 2419 3240
rect 2551 3236 2555 3240
rect 2687 3236 2691 3240
rect 2831 3236 2835 3240
rect 2975 3236 2979 3240
rect 3119 3236 3123 3240
rect 3255 3236 3259 3240
rect 3383 3236 3387 3240
rect 3503 3236 3507 3240
rect 3623 3236 3627 3240
rect 3743 3236 3747 3240
rect 3839 3236 3843 3240
rect 3943 3239 3947 3243
rect 111 3224 115 3228
rect 135 3223 139 3227
rect 319 3223 323 3227
rect 519 3223 523 3227
rect 719 3223 723 3227
rect 911 3223 915 3227
rect 1095 3223 1099 3227
rect 1271 3223 1275 3227
rect 1447 3223 1451 3227
rect 1623 3223 1627 3227
rect 1799 3223 1803 3227
rect 2007 3224 2011 3228
rect 111 3207 115 3211
rect 135 3204 139 3208
rect 319 3204 323 3208
rect 519 3204 523 3208
rect 719 3204 723 3208
rect 911 3204 915 3208
rect 1095 3204 1099 3208
rect 1271 3204 1275 3208
rect 1447 3204 1451 3208
rect 1623 3204 1627 3208
rect 1799 3204 1803 3208
rect 2007 3207 2011 3211
rect 2047 3161 2051 3165
rect 2247 3164 2251 3168
rect 2399 3164 2403 3168
rect 2559 3164 2563 3168
rect 2727 3164 2731 3168
rect 2903 3164 2907 3168
rect 3079 3164 3083 3168
rect 3263 3164 3267 3168
rect 3447 3164 3451 3168
rect 3631 3164 3635 3168
rect 3815 3164 3819 3168
rect 3943 3161 3947 3165
rect 2047 3144 2051 3148
rect 2247 3145 2251 3149
rect 2399 3145 2403 3149
rect 2559 3145 2563 3149
rect 2727 3145 2731 3149
rect 2903 3145 2907 3149
rect 3079 3145 3083 3149
rect 3263 3145 3267 3149
rect 3447 3145 3451 3149
rect 3631 3145 3635 3149
rect 3815 3145 3819 3149
rect 3943 3144 3947 3148
rect 111 3133 115 3137
rect 143 3136 147 3140
rect 343 3136 347 3140
rect 543 3136 547 3140
rect 743 3136 747 3140
rect 927 3136 931 3140
rect 1103 3136 1107 3140
rect 1263 3136 1267 3140
rect 1423 3136 1427 3140
rect 1575 3136 1579 3140
rect 1735 3136 1739 3140
rect 2007 3133 2011 3137
rect 111 3116 115 3120
rect 143 3117 147 3121
rect 343 3117 347 3121
rect 543 3117 547 3121
rect 743 3117 747 3121
rect 927 3117 931 3121
rect 1103 3117 1107 3121
rect 1263 3117 1267 3121
rect 1423 3117 1427 3121
rect 1575 3117 1579 3121
rect 1735 3117 1739 3121
rect 2007 3116 2011 3120
rect 2047 3088 2051 3092
rect 2079 3087 2083 3091
rect 2223 3087 2227 3091
rect 2375 3087 2379 3091
rect 2527 3087 2531 3091
rect 2687 3087 2691 3091
rect 2855 3087 2859 3091
rect 3039 3087 3043 3091
rect 3231 3087 3235 3091
rect 3431 3087 3435 3091
rect 3639 3087 3643 3091
rect 3839 3087 3843 3091
rect 3943 3088 3947 3092
rect 2047 3071 2051 3075
rect 111 3064 115 3068
rect 263 3063 267 3067
rect 439 3063 443 3067
rect 615 3063 619 3067
rect 799 3063 803 3067
rect 975 3063 979 3067
rect 1143 3063 1147 3067
rect 1303 3063 1307 3067
rect 1455 3063 1459 3067
rect 1607 3063 1611 3067
rect 1767 3063 1771 3067
rect 2007 3064 2011 3068
rect 2079 3068 2083 3072
rect 2223 3068 2227 3072
rect 2375 3068 2379 3072
rect 2527 3068 2531 3072
rect 2687 3068 2691 3072
rect 2855 3068 2859 3072
rect 3039 3068 3043 3072
rect 3231 3068 3235 3072
rect 3431 3068 3435 3072
rect 3639 3068 3643 3072
rect 3839 3068 3843 3072
rect 3943 3071 3947 3075
rect 111 3047 115 3051
rect 263 3044 267 3048
rect 439 3044 443 3048
rect 615 3044 619 3048
rect 799 3044 803 3048
rect 975 3044 979 3048
rect 1143 3044 1147 3048
rect 1303 3044 1307 3048
rect 1455 3044 1459 3048
rect 1607 3044 1611 3048
rect 1767 3044 1771 3048
rect 2007 3047 2011 3051
rect 2047 2997 2051 3001
rect 2071 3000 2075 3004
rect 2183 3000 2187 3004
rect 2327 3000 2331 3004
rect 2479 3000 2483 3004
rect 2655 3000 2659 3004
rect 2855 3000 2859 3004
rect 3087 3000 3091 3004
rect 3335 3000 3339 3004
rect 3599 3000 3603 3004
rect 3839 3000 3843 3004
rect 3943 2997 3947 3001
rect 2047 2980 2051 2984
rect 2071 2981 2075 2985
rect 2183 2981 2187 2985
rect 2327 2981 2331 2985
rect 2479 2981 2483 2985
rect 2655 2981 2659 2985
rect 2855 2981 2859 2985
rect 3087 2981 3091 2985
rect 3335 2981 3339 2985
rect 3599 2981 3603 2985
rect 3839 2981 3843 2985
rect 3943 2980 3947 2984
rect 111 2957 115 2961
rect 343 2960 347 2964
rect 439 2960 443 2964
rect 543 2960 547 2964
rect 655 2960 659 2964
rect 783 2960 787 2964
rect 935 2960 939 2964
rect 1103 2960 1107 2964
rect 1295 2960 1299 2964
rect 1495 2960 1499 2964
rect 1711 2960 1715 2964
rect 1903 2960 1907 2964
rect 2007 2957 2011 2961
rect 111 2940 115 2944
rect 343 2941 347 2945
rect 439 2941 443 2945
rect 543 2941 547 2945
rect 655 2941 659 2945
rect 783 2941 787 2945
rect 935 2941 939 2945
rect 1103 2941 1107 2945
rect 1295 2941 1299 2945
rect 1495 2941 1499 2945
rect 1711 2941 1715 2945
rect 1903 2941 1907 2945
rect 2007 2940 2011 2944
rect 2047 2924 2051 2928
rect 2071 2923 2075 2927
rect 2263 2923 2267 2927
rect 2487 2923 2491 2927
rect 2735 2923 2739 2927
rect 2999 2923 3003 2927
rect 3279 2923 3283 2927
rect 3567 2923 3571 2927
rect 3839 2923 3843 2927
rect 3943 2924 3947 2928
rect 2047 2907 2051 2911
rect 2071 2904 2075 2908
rect 2263 2904 2267 2908
rect 2487 2904 2491 2908
rect 2735 2904 2739 2908
rect 2999 2904 3003 2908
rect 3279 2904 3283 2908
rect 3567 2904 3571 2908
rect 3839 2904 3843 2908
rect 3943 2907 3947 2911
rect 111 2888 115 2892
rect 207 2887 211 2891
rect 327 2887 331 2891
rect 447 2887 451 2891
rect 575 2887 579 2891
rect 703 2887 707 2891
rect 847 2887 851 2891
rect 999 2887 1003 2891
rect 1167 2887 1171 2891
rect 1351 2887 1355 2891
rect 1535 2887 1539 2891
rect 1727 2887 1731 2891
rect 1903 2887 1907 2891
rect 2007 2888 2011 2892
rect 111 2871 115 2875
rect 207 2868 211 2872
rect 327 2868 331 2872
rect 447 2868 451 2872
rect 575 2868 579 2872
rect 703 2868 707 2872
rect 847 2868 851 2872
rect 999 2868 1003 2872
rect 1167 2868 1171 2872
rect 1351 2868 1355 2872
rect 1535 2868 1539 2872
rect 1727 2868 1731 2872
rect 1903 2868 1907 2872
rect 2007 2871 2011 2875
rect 2047 2833 2051 2837
rect 2671 2836 2675 2840
rect 2887 2836 2891 2840
rect 3095 2836 3099 2840
rect 3287 2836 3291 2840
rect 3479 2836 3483 2840
rect 3671 2836 3675 2840
rect 3839 2836 3843 2840
rect 3943 2833 3947 2837
rect 2047 2816 2051 2820
rect 2671 2817 2675 2821
rect 2887 2817 2891 2821
rect 3095 2817 3099 2821
rect 3287 2817 3291 2821
rect 3479 2817 3483 2821
rect 3671 2817 3675 2821
rect 3839 2817 3843 2821
rect 3943 2816 3947 2820
rect 111 2801 115 2805
rect 135 2804 139 2808
rect 247 2804 251 2808
rect 399 2804 403 2808
rect 551 2804 555 2808
rect 711 2804 715 2808
rect 879 2804 883 2808
rect 1047 2804 1051 2808
rect 1223 2804 1227 2808
rect 1399 2804 1403 2808
rect 1575 2804 1579 2808
rect 1751 2804 1755 2808
rect 1903 2804 1907 2808
rect 2007 2801 2011 2805
rect 111 2784 115 2788
rect 135 2785 139 2789
rect 247 2785 251 2789
rect 399 2785 403 2789
rect 551 2785 555 2789
rect 711 2785 715 2789
rect 879 2785 883 2789
rect 1047 2785 1051 2789
rect 1223 2785 1227 2789
rect 1399 2785 1403 2789
rect 1575 2785 1579 2789
rect 1751 2785 1755 2789
rect 1903 2785 1907 2789
rect 2007 2784 2011 2788
rect 2047 2764 2051 2768
rect 2071 2763 2075 2767
rect 2199 2763 2203 2767
rect 2343 2763 2347 2767
rect 2479 2763 2483 2767
rect 2607 2763 2611 2767
rect 2727 2763 2731 2767
rect 2839 2763 2843 2767
rect 2943 2763 2947 2767
rect 3047 2763 3051 2767
rect 3143 2763 3147 2767
rect 3239 2763 3243 2767
rect 3343 2763 3347 2767
rect 3447 2763 3451 2767
rect 3551 2763 3555 2767
rect 3647 2763 3651 2767
rect 3743 2763 3747 2767
rect 3839 2763 3843 2767
rect 3943 2764 3947 2768
rect 2047 2747 2051 2751
rect 2071 2744 2075 2748
rect 2199 2744 2203 2748
rect 2343 2744 2347 2748
rect 2479 2744 2483 2748
rect 2607 2744 2611 2748
rect 2727 2744 2731 2748
rect 2839 2744 2843 2748
rect 2943 2744 2947 2748
rect 3047 2744 3051 2748
rect 3143 2744 3147 2748
rect 3239 2744 3243 2748
rect 3343 2744 3347 2748
rect 3447 2744 3451 2748
rect 3551 2744 3555 2748
rect 3647 2744 3651 2748
rect 3743 2744 3747 2748
rect 3839 2744 3843 2748
rect 3943 2747 3947 2751
rect 111 2724 115 2728
rect 135 2723 139 2727
rect 255 2723 259 2727
rect 407 2723 411 2727
rect 575 2723 579 2727
rect 743 2723 747 2727
rect 919 2723 923 2727
rect 1087 2723 1091 2727
rect 1255 2723 1259 2727
rect 1423 2723 1427 2727
rect 1599 2723 1603 2727
rect 2007 2724 2011 2728
rect 111 2707 115 2711
rect 135 2704 139 2708
rect 255 2704 259 2708
rect 407 2704 411 2708
rect 575 2704 579 2708
rect 743 2704 747 2708
rect 919 2704 923 2708
rect 1087 2704 1091 2708
rect 1255 2704 1259 2708
rect 1423 2704 1427 2708
rect 1599 2704 1603 2708
rect 2007 2707 2011 2711
rect 2047 2661 2051 2665
rect 2095 2664 2099 2668
rect 2263 2664 2267 2668
rect 2439 2664 2443 2668
rect 2615 2664 2619 2668
rect 2783 2664 2787 2668
rect 2943 2664 2947 2668
rect 3095 2664 3099 2668
rect 3239 2664 3243 2668
rect 3383 2664 3387 2668
rect 3535 2664 3539 2668
rect 3943 2661 3947 2665
rect 111 2641 115 2645
rect 167 2644 171 2648
rect 359 2644 363 2648
rect 559 2644 563 2648
rect 759 2644 763 2648
rect 951 2644 955 2648
rect 1143 2644 1147 2648
rect 1327 2644 1331 2648
rect 1511 2644 1515 2648
rect 1703 2644 1707 2648
rect 2007 2641 2011 2645
rect 2047 2644 2051 2648
rect 2095 2645 2099 2649
rect 2263 2645 2267 2649
rect 2439 2645 2443 2649
rect 2615 2645 2619 2649
rect 2783 2645 2787 2649
rect 2943 2645 2947 2649
rect 3095 2645 3099 2649
rect 3239 2645 3243 2649
rect 3383 2645 3387 2649
rect 3535 2645 3539 2649
rect 3943 2644 3947 2648
rect 111 2624 115 2628
rect 167 2625 171 2629
rect 359 2625 363 2629
rect 559 2625 563 2629
rect 759 2625 763 2629
rect 951 2625 955 2629
rect 1143 2625 1147 2629
rect 1327 2625 1331 2629
rect 1511 2625 1515 2629
rect 1703 2625 1707 2629
rect 2007 2624 2011 2628
rect 2047 2584 2051 2588
rect 2215 2583 2219 2587
rect 2367 2583 2371 2587
rect 2519 2583 2523 2587
rect 2671 2583 2675 2587
rect 2815 2583 2819 2587
rect 2951 2583 2955 2587
rect 3087 2583 3091 2587
rect 3223 2583 3227 2587
rect 3367 2583 3371 2587
rect 3943 2584 3947 2588
rect 2047 2567 2051 2571
rect 2215 2564 2219 2568
rect 2367 2564 2371 2568
rect 2519 2564 2523 2568
rect 2671 2564 2675 2568
rect 2815 2564 2819 2568
rect 2951 2564 2955 2568
rect 3087 2564 3091 2568
rect 3223 2564 3227 2568
rect 3367 2564 3371 2568
rect 3943 2567 3947 2571
rect 111 2556 115 2560
rect 575 2555 579 2559
rect 687 2555 691 2559
rect 807 2555 811 2559
rect 935 2555 939 2559
rect 1071 2555 1075 2559
rect 1207 2555 1211 2559
rect 1351 2555 1355 2559
rect 1495 2555 1499 2559
rect 1647 2555 1651 2559
rect 1799 2555 1803 2559
rect 2007 2556 2011 2560
rect 111 2539 115 2543
rect 575 2536 579 2540
rect 687 2536 691 2540
rect 807 2536 811 2540
rect 935 2536 939 2540
rect 1071 2536 1075 2540
rect 1207 2536 1211 2540
rect 1351 2536 1355 2540
rect 1495 2536 1499 2540
rect 1647 2536 1651 2540
rect 1799 2536 1803 2540
rect 2007 2539 2011 2543
rect 2047 2497 2051 2501
rect 2095 2500 2099 2504
rect 2215 2500 2219 2504
rect 2343 2500 2347 2504
rect 2471 2500 2475 2504
rect 2599 2500 2603 2504
rect 2719 2500 2723 2504
rect 2839 2500 2843 2504
rect 2967 2500 2971 2504
rect 3095 2500 3099 2504
rect 3223 2500 3227 2504
rect 3943 2497 3947 2501
rect 2047 2480 2051 2484
rect 2095 2481 2099 2485
rect 2215 2481 2219 2485
rect 2343 2481 2347 2485
rect 2471 2481 2475 2485
rect 2599 2481 2603 2485
rect 2719 2481 2723 2485
rect 2839 2481 2843 2485
rect 2967 2481 2971 2485
rect 3095 2481 3099 2485
rect 3223 2481 3227 2485
rect 3943 2480 3947 2484
rect 111 2469 115 2473
rect 503 2472 507 2476
rect 607 2472 611 2476
rect 719 2472 723 2476
rect 847 2472 851 2476
rect 983 2472 987 2476
rect 1127 2472 1131 2476
rect 1279 2472 1283 2476
rect 1431 2472 1435 2476
rect 1583 2472 1587 2476
rect 1743 2472 1747 2476
rect 1903 2472 1907 2476
rect 2007 2469 2011 2473
rect 111 2452 115 2456
rect 503 2453 507 2457
rect 607 2453 611 2457
rect 719 2453 723 2457
rect 847 2453 851 2457
rect 983 2453 987 2457
rect 1127 2453 1131 2457
rect 1279 2453 1283 2457
rect 1431 2453 1435 2457
rect 1583 2453 1587 2457
rect 1743 2453 1747 2457
rect 1903 2453 1907 2457
rect 2007 2452 2011 2456
rect 2047 2416 2051 2420
rect 2071 2415 2075 2419
rect 2191 2415 2195 2419
rect 2319 2415 2323 2419
rect 2439 2415 2443 2419
rect 2559 2415 2563 2419
rect 2679 2415 2683 2419
rect 2791 2415 2795 2419
rect 2911 2415 2915 2419
rect 3031 2415 3035 2419
rect 3151 2415 3155 2419
rect 3943 2416 3947 2420
rect 2047 2399 2051 2403
rect 2071 2396 2075 2400
rect 2191 2396 2195 2400
rect 2319 2396 2323 2400
rect 2439 2396 2443 2400
rect 2559 2396 2563 2400
rect 2679 2396 2683 2400
rect 2791 2396 2795 2400
rect 2911 2396 2915 2400
rect 3031 2396 3035 2400
rect 3151 2396 3155 2400
rect 3943 2399 3947 2403
rect 111 2384 115 2388
rect 535 2383 539 2387
rect 671 2383 675 2387
rect 815 2383 819 2387
rect 959 2383 963 2387
rect 1103 2383 1107 2387
rect 1247 2383 1251 2387
rect 1391 2383 1395 2387
rect 1527 2383 1531 2387
rect 1655 2383 1659 2387
rect 1791 2383 1795 2387
rect 1903 2383 1907 2387
rect 2007 2384 2011 2388
rect 111 2367 115 2371
rect 535 2364 539 2368
rect 671 2364 675 2368
rect 815 2364 819 2368
rect 959 2364 963 2368
rect 1103 2364 1107 2368
rect 1247 2364 1251 2368
rect 1391 2364 1395 2368
rect 1527 2364 1531 2368
rect 1655 2364 1659 2368
rect 1791 2364 1795 2368
rect 1903 2364 1907 2368
rect 2007 2367 2011 2371
rect 2047 2329 2051 2333
rect 2167 2332 2171 2336
rect 2359 2332 2363 2336
rect 2535 2332 2539 2336
rect 2703 2332 2707 2336
rect 2871 2332 2875 2336
rect 3031 2332 3035 2336
rect 3199 2332 3203 2336
rect 3943 2329 3947 2333
rect 2047 2312 2051 2316
rect 2167 2313 2171 2317
rect 2359 2313 2363 2317
rect 2535 2313 2539 2317
rect 2703 2313 2707 2317
rect 2871 2313 2875 2317
rect 3031 2313 3035 2317
rect 3199 2313 3203 2317
rect 3943 2312 3947 2316
rect 111 2297 115 2301
rect 535 2300 539 2304
rect 647 2300 651 2304
rect 767 2300 771 2304
rect 895 2300 899 2304
rect 1031 2300 1035 2304
rect 1167 2300 1171 2304
rect 1295 2300 1299 2304
rect 1423 2300 1427 2304
rect 1551 2300 1555 2304
rect 1671 2300 1675 2304
rect 1799 2300 1803 2304
rect 1903 2300 1907 2304
rect 2007 2297 2011 2301
rect 111 2280 115 2284
rect 535 2281 539 2285
rect 647 2281 651 2285
rect 767 2281 771 2285
rect 895 2281 899 2285
rect 1031 2281 1035 2285
rect 1167 2281 1171 2285
rect 1295 2281 1299 2285
rect 1423 2281 1427 2285
rect 1551 2281 1555 2285
rect 1671 2281 1675 2285
rect 1799 2281 1803 2285
rect 1903 2281 1907 2285
rect 2007 2280 2011 2284
rect 2047 2260 2051 2264
rect 2071 2259 2075 2263
rect 2167 2259 2171 2263
rect 2287 2259 2291 2263
rect 2423 2259 2427 2263
rect 2559 2259 2563 2263
rect 2703 2259 2707 2263
rect 2839 2259 2843 2263
rect 2983 2259 2987 2263
rect 3127 2259 3131 2263
rect 3271 2259 3275 2263
rect 3943 2260 3947 2264
rect 2047 2243 2051 2247
rect 2071 2240 2075 2244
rect 2167 2240 2171 2244
rect 2287 2240 2291 2244
rect 2423 2240 2427 2244
rect 2559 2240 2563 2244
rect 2703 2240 2707 2244
rect 2839 2240 2843 2244
rect 2983 2240 2987 2244
rect 3127 2240 3131 2244
rect 3271 2240 3275 2244
rect 3943 2243 3947 2247
rect 111 2224 115 2228
rect 415 2223 419 2227
rect 535 2223 539 2227
rect 671 2223 675 2227
rect 823 2223 827 2227
rect 991 2223 995 2227
rect 1175 2223 1179 2227
rect 1367 2223 1371 2227
rect 1567 2223 1571 2227
rect 1767 2223 1771 2227
rect 2007 2224 2011 2228
rect 111 2207 115 2211
rect 415 2204 419 2208
rect 535 2204 539 2208
rect 671 2204 675 2208
rect 823 2204 827 2208
rect 991 2204 995 2208
rect 1175 2204 1179 2208
rect 1367 2204 1371 2208
rect 1567 2204 1571 2208
rect 1767 2204 1771 2208
rect 2007 2207 2011 2211
rect 2047 2177 2051 2181
rect 2071 2180 2075 2184
rect 2295 2180 2299 2184
rect 2503 2180 2507 2184
rect 2687 2180 2691 2184
rect 2863 2180 2867 2184
rect 3023 2180 3027 2184
rect 3175 2180 3179 2184
rect 3319 2180 3323 2184
rect 3471 2180 3475 2184
rect 3943 2177 3947 2181
rect 2047 2160 2051 2164
rect 2071 2161 2075 2165
rect 2295 2161 2299 2165
rect 2503 2161 2507 2165
rect 2687 2161 2691 2165
rect 2863 2161 2867 2165
rect 3023 2161 3027 2165
rect 3175 2161 3179 2165
rect 3319 2161 3323 2165
rect 3471 2161 3475 2165
rect 3943 2160 3947 2164
rect 111 2133 115 2137
rect 135 2136 139 2140
rect 247 2136 251 2140
rect 391 2136 395 2140
rect 551 2136 555 2140
rect 711 2136 715 2140
rect 871 2136 875 2140
rect 1031 2136 1035 2140
rect 1191 2136 1195 2140
rect 1351 2136 1355 2140
rect 1511 2136 1515 2140
rect 1679 2136 1683 2140
rect 2007 2133 2011 2137
rect 111 2116 115 2120
rect 135 2117 139 2121
rect 247 2117 251 2121
rect 391 2117 395 2121
rect 551 2117 555 2121
rect 711 2117 715 2121
rect 871 2117 875 2121
rect 1031 2117 1035 2121
rect 1191 2117 1195 2121
rect 1351 2117 1355 2121
rect 1511 2117 1515 2121
rect 1679 2117 1683 2121
rect 2007 2116 2011 2120
rect 2047 2084 2051 2088
rect 2399 2083 2403 2087
rect 2495 2083 2499 2087
rect 2591 2083 2595 2087
rect 2687 2083 2691 2087
rect 2783 2083 2787 2087
rect 2879 2083 2883 2087
rect 2975 2083 2979 2087
rect 3071 2083 3075 2087
rect 3167 2083 3171 2087
rect 3263 2083 3267 2087
rect 3359 2083 3363 2087
rect 3455 2083 3459 2087
rect 3551 2083 3555 2087
rect 3647 2083 3651 2087
rect 3743 2083 3747 2087
rect 3839 2083 3843 2087
rect 3943 2084 3947 2088
rect 2047 2067 2051 2071
rect 2399 2064 2403 2068
rect 2495 2064 2499 2068
rect 2591 2064 2595 2068
rect 2687 2064 2691 2068
rect 2783 2064 2787 2068
rect 2879 2064 2883 2068
rect 2975 2064 2979 2068
rect 3071 2064 3075 2068
rect 3167 2064 3171 2068
rect 3263 2064 3267 2068
rect 3359 2064 3363 2068
rect 3455 2064 3459 2068
rect 3551 2064 3555 2068
rect 3647 2064 3651 2068
rect 3743 2064 3747 2068
rect 3839 2064 3843 2068
rect 3943 2067 3947 2071
rect 111 2056 115 2060
rect 135 2055 139 2059
rect 247 2055 251 2059
rect 399 2055 403 2059
rect 551 2055 555 2059
rect 703 2055 707 2059
rect 847 2055 851 2059
rect 991 2055 995 2059
rect 1127 2055 1131 2059
rect 1255 2055 1259 2059
rect 1383 2055 1387 2059
rect 1519 2055 1523 2059
rect 2007 2056 2011 2060
rect 111 2039 115 2043
rect 135 2036 139 2040
rect 247 2036 251 2040
rect 399 2036 403 2040
rect 551 2036 555 2040
rect 703 2036 707 2040
rect 847 2036 851 2040
rect 991 2036 995 2040
rect 1127 2036 1131 2040
rect 1255 2036 1259 2040
rect 1383 2036 1387 2040
rect 1519 2036 1523 2040
rect 2007 2039 2011 2043
rect 2047 2001 2051 2005
rect 2191 2004 2195 2008
rect 2399 2004 2403 2008
rect 2647 2004 2651 2008
rect 2919 2004 2923 2008
rect 3215 2004 3219 2008
rect 3527 2004 3531 2008
rect 3839 2004 3843 2008
rect 3943 2001 3947 2005
rect 2047 1984 2051 1988
rect 2191 1985 2195 1989
rect 2399 1985 2403 1989
rect 2647 1985 2651 1989
rect 2919 1985 2923 1989
rect 3215 1985 3219 1989
rect 3527 1985 3531 1989
rect 3839 1985 3843 1989
rect 3943 1984 3947 1988
rect 111 1957 115 1961
rect 231 1960 235 1964
rect 391 1960 395 1964
rect 567 1960 571 1964
rect 751 1960 755 1964
rect 943 1960 947 1964
rect 1135 1960 1139 1964
rect 1335 1960 1339 1964
rect 1543 1960 1547 1964
rect 2007 1957 2011 1961
rect 111 1940 115 1944
rect 231 1941 235 1945
rect 391 1941 395 1945
rect 567 1941 571 1945
rect 751 1941 755 1945
rect 943 1941 947 1945
rect 1135 1941 1139 1945
rect 1335 1941 1339 1945
rect 1543 1941 1547 1945
rect 2007 1940 2011 1944
rect 2047 1920 2051 1924
rect 2071 1919 2075 1923
rect 2239 1919 2243 1923
rect 2447 1919 2451 1923
rect 2671 1919 2675 1923
rect 2895 1919 2899 1923
rect 3127 1919 3131 1923
rect 3359 1919 3363 1923
rect 3591 1919 3595 1923
rect 3831 1919 3835 1923
rect 3943 1920 3947 1924
rect 2047 1903 2051 1907
rect 2071 1900 2075 1904
rect 2239 1900 2243 1904
rect 2447 1900 2451 1904
rect 2671 1900 2675 1904
rect 2895 1900 2899 1904
rect 3127 1900 3131 1904
rect 3359 1900 3363 1904
rect 3591 1900 3595 1904
rect 3831 1900 3835 1904
rect 3943 1903 3947 1907
rect 111 1888 115 1892
rect 511 1887 515 1891
rect 623 1887 627 1891
rect 743 1887 747 1891
rect 863 1887 867 1891
rect 983 1887 987 1891
rect 1103 1887 1107 1891
rect 1223 1887 1227 1891
rect 1335 1887 1339 1891
rect 1455 1887 1459 1891
rect 1575 1887 1579 1891
rect 1695 1887 1699 1891
rect 2007 1888 2011 1892
rect 111 1871 115 1875
rect 511 1868 515 1872
rect 623 1868 627 1872
rect 743 1868 747 1872
rect 863 1868 867 1872
rect 983 1868 987 1872
rect 1103 1868 1107 1872
rect 1223 1868 1227 1872
rect 1335 1868 1339 1872
rect 1455 1868 1459 1872
rect 1575 1868 1579 1872
rect 1695 1868 1699 1872
rect 2007 1871 2011 1875
rect 2047 1837 2051 1841
rect 2071 1840 2075 1844
rect 2199 1840 2203 1844
rect 2367 1840 2371 1844
rect 2543 1840 2547 1844
rect 2719 1840 2723 1844
rect 2887 1840 2891 1844
rect 3039 1840 3043 1844
rect 3183 1840 3187 1844
rect 3319 1840 3323 1844
rect 3455 1840 3459 1844
rect 3583 1840 3587 1844
rect 3711 1840 3715 1844
rect 3839 1840 3843 1844
rect 3943 1837 3947 1841
rect 2047 1820 2051 1824
rect 2071 1821 2075 1825
rect 2199 1821 2203 1825
rect 2367 1821 2371 1825
rect 2543 1821 2547 1825
rect 2719 1821 2723 1825
rect 2887 1821 2891 1825
rect 3039 1821 3043 1825
rect 3183 1821 3187 1825
rect 3319 1821 3323 1825
rect 3455 1821 3459 1825
rect 3583 1821 3587 1825
rect 3711 1821 3715 1825
rect 3839 1821 3843 1825
rect 3943 1820 3947 1824
rect 111 1797 115 1801
rect 615 1800 619 1804
rect 711 1800 715 1804
rect 815 1800 819 1804
rect 927 1800 931 1804
rect 1039 1800 1043 1804
rect 1159 1800 1163 1804
rect 1279 1800 1283 1804
rect 1399 1800 1403 1804
rect 1519 1800 1523 1804
rect 1639 1800 1643 1804
rect 2007 1797 2011 1801
rect 111 1780 115 1784
rect 615 1781 619 1785
rect 711 1781 715 1785
rect 815 1781 819 1785
rect 927 1781 931 1785
rect 1039 1781 1043 1785
rect 1159 1781 1163 1785
rect 1279 1781 1283 1785
rect 1399 1781 1403 1785
rect 1519 1781 1523 1785
rect 1639 1781 1643 1785
rect 2007 1780 2011 1784
rect 2047 1764 2051 1768
rect 2071 1763 2075 1767
rect 2183 1763 2187 1767
rect 2327 1763 2331 1767
rect 2487 1763 2491 1767
rect 2655 1763 2659 1767
rect 2831 1763 2835 1767
rect 3023 1763 3027 1767
rect 3223 1763 3227 1767
rect 3431 1763 3435 1767
rect 3647 1763 3651 1767
rect 3839 1763 3843 1767
rect 3943 1764 3947 1768
rect 2047 1747 2051 1751
rect 2071 1744 2075 1748
rect 2183 1744 2187 1748
rect 2327 1744 2331 1748
rect 2487 1744 2491 1748
rect 2655 1744 2659 1748
rect 2831 1744 2835 1748
rect 3023 1744 3027 1748
rect 3223 1744 3227 1748
rect 3431 1744 3435 1748
rect 3647 1744 3651 1748
rect 3839 1744 3843 1748
rect 3943 1747 3947 1751
rect 111 1728 115 1732
rect 367 1727 371 1731
rect 495 1727 499 1731
rect 639 1727 643 1731
rect 799 1727 803 1731
rect 967 1727 971 1731
rect 1143 1727 1147 1731
rect 1327 1727 1331 1731
rect 1511 1727 1515 1731
rect 1703 1727 1707 1731
rect 2007 1728 2011 1732
rect 111 1711 115 1715
rect 367 1708 371 1712
rect 495 1708 499 1712
rect 639 1708 643 1712
rect 799 1708 803 1712
rect 967 1708 971 1712
rect 1143 1708 1147 1712
rect 1327 1708 1331 1712
rect 1511 1708 1515 1712
rect 1703 1708 1707 1712
rect 2007 1711 2011 1715
rect 2047 1673 2051 1677
rect 2223 1676 2227 1680
rect 2327 1676 2331 1680
rect 2439 1676 2443 1680
rect 2559 1676 2563 1680
rect 2687 1676 2691 1680
rect 2823 1676 2827 1680
rect 2967 1676 2971 1680
rect 3127 1676 3131 1680
rect 3303 1676 3307 1680
rect 3487 1676 3491 1680
rect 3671 1676 3675 1680
rect 3839 1676 3843 1680
rect 3943 1673 3947 1677
rect 2047 1656 2051 1660
rect 2223 1657 2227 1661
rect 2327 1657 2331 1661
rect 2439 1657 2443 1661
rect 2559 1657 2563 1661
rect 2687 1657 2691 1661
rect 2823 1657 2827 1661
rect 2967 1657 2971 1661
rect 3127 1657 3131 1661
rect 3303 1657 3307 1661
rect 3487 1657 3491 1661
rect 3671 1657 3675 1661
rect 3839 1657 3843 1661
rect 3943 1656 3947 1660
rect 111 1641 115 1645
rect 135 1644 139 1648
rect 247 1644 251 1648
rect 399 1644 403 1648
rect 567 1644 571 1648
rect 743 1644 747 1648
rect 935 1644 939 1648
rect 1135 1644 1139 1648
rect 1343 1644 1347 1648
rect 1551 1644 1555 1648
rect 1767 1644 1771 1648
rect 2007 1641 2011 1645
rect 111 1624 115 1628
rect 135 1625 139 1629
rect 247 1625 251 1629
rect 399 1625 403 1629
rect 567 1625 571 1629
rect 743 1625 747 1629
rect 935 1625 939 1629
rect 1135 1625 1139 1629
rect 1343 1625 1347 1629
rect 1551 1625 1555 1629
rect 1767 1625 1771 1629
rect 2007 1624 2011 1628
rect 2047 1600 2051 1604
rect 2391 1599 2395 1603
rect 2503 1599 2507 1603
rect 2615 1599 2619 1603
rect 2735 1599 2739 1603
rect 2855 1599 2859 1603
rect 2975 1599 2979 1603
rect 3095 1599 3099 1603
rect 3215 1599 3219 1603
rect 3335 1599 3339 1603
rect 3455 1599 3459 1603
rect 3943 1600 3947 1604
rect 2047 1583 2051 1587
rect 2391 1580 2395 1584
rect 2503 1580 2507 1584
rect 2615 1580 2619 1584
rect 2735 1580 2739 1584
rect 2855 1580 2859 1584
rect 2975 1580 2979 1584
rect 3095 1580 3099 1584
rect 3215 1580 3219 1584
rect 3335 1580 3339 1584
rect 3455 1580 3459 1584
rect 3943 1583 3947 1587
rect 111 1568 115 1572
rect 135 1567 139 1571
rect 255 1567 259 1571
rect 423 1567 427 1571
rect 615 1567 619 1571
rect 831 1567 835 1571
rect 1063 1567 1067 1571
rect 1311 1567 1315 1571
rect 1567 1567 1571 1571
rect 1831 1567 1835 1571
rect 2007 1568 2011 1572
rect 111 1551 115 1555
rect 135 1548 139 1552
rect 255 1548 259 1552
rect 423 1548 427 1552
rect 615 1548 619 1552
rect 831 1548 835 1552
rect 1063 1548 1067 1552
rect 1311 1548 1315 1552
rect 1567 1548 1571 1552
rect 1831 1548 1835 1552
rect 2007 1551 2011 1555
rect 2047 1517 2051 1521
rect 2543 1520 2547 1524
rect 2671 1520 2675 1524
rect 2799 1520 2803 1524
rect 2935 1520 2939 1524
rect 3071 1520 3075 1524
rect 3207 1520 3211 1524
rect 3335 1520 3339 1524
rect 3463 1520 3467 1524
rect 3591 1520 3595 1524
rect 3727 1520 3731 1524
rect 3839 1520 3843 1524
rect 3943 1517 3947 1521
rect 2047 1500 2051 1504
rect 2543 1501 2547 1505
rect 2671 1501 2675 1505
rect 2799 1501 2803 1505
rect 2935 1501 2939 1505
rect 3071 1501 3075 1505
rect 3207 1501 3211 1505
rect 3335 1501 3339 1505
rect 3463 1501 3467 1505
rect 3591 1501 3595 1505
rect 3727 1501 3731 1505
rect 3839 1501 3843 1505
rect 3943 1500 3947 1504
rect 111 1481 115 1485
rect 239 1484 243 1488
rect 407 1484 411 1488
rect 583 1484 587 1488
rect 775 1484 779 1488
rect 967 1484 971 1488
rect 1159 1484 1163 1488
rect 1351 1484 1355 1488
rect 1543 1484 1547 1488
rect 1735 1484 1739 1488
rect 1903 1484 1907 1488
rect 2007 1481 2011 1485
rect 111 1464 115 1468
rect 239 1465 243 1469
rect 407 1465 411 1469
rect 583 1465 587 1469
rect 775 1465 779 1469
rect 967 1465 971 1469
rect 1159 1465 1163 1469
rect 1351 1465 1355 1469
rect 1543 1465 1547 1469
rect 1735 1465 1739 1469
rect 1903 1465 1907 1469
rect 2007 1464 2011 1468
rect 2047 1436 2051 1440
rect 2519 1435 2523 1439
rect 2631 1435 2635 1439
rect 2759 1435 2763 1439
rect 2895 1435 2899 1439
rect 3031 1435 3035 1439
rect 3175 1435 3179 1439
rect 3311 1435 3315 1439
rect 3447 1435 3451 1439
rect 3583 1435 3587 1439
rect 3719 1435 3723 1439
rect 3839 1435 3843 1439
rect 3943 1436 3947 1440
rect 2047 1419 2051 1423
rect 2519 1416 2523 1420
rect 2631 1416 2635 1420
rect 2759 1416 2763 1420
rect 2895 1416 2899 1420
rect 3031 1416 3035 1420
rect 3175 1416 3179 1420
rect 3311 1416 3315 1420
rect 3447 1416 3451 1420
rect 3583 1416 3587 1420
rect 3719 1416 3723 1420
rect 3839 1416 3843 1420
rect 3943 1419 3947 1423
rect 111 1404 115 1408
rect 463 1403 467 1407
rect 583 1403 587 1407
rect 711 1403 715 1407
rect 855 1403 859 1407
rect 1007 1403 1011 1407
rect 1167 1403 1171 1407
rect 1335 1403 1339 1407
rect 1511 1403 1515 1407
rect 1687 1403 1691 1407
rect 1871 1403 1875 1407
rect 2007 1404 2011 1408
rect 111 1387 115 1391
rect 463 1384 467 1388
rect 583 1384 587 1388
rect 711 1384 715 1388
rect 855 1384 859 1388
rect 1007 1384 1011 1388
rect 1167 1384 1171 1388
rect 1335 1384 1339 1388
rect 1511 1384 1515 1388
rect 1687 1384 1691 1388
rect 1871 1384 1875 1388
rect 2007 1387 2011 1391
rect 2047 1353 2051 1357
rect 2399 1356 2403 1360
rect 2535 1356 2539 1360
rect 2679 1356 2683 1360
rect 2823 1356 2827 1360
rect 2967 1356 2971 1360
rect 3111 1356 3115 1360
rect 3255 1356 3259 1360
rect 3407 1356 3411 1360
rect 3559 1356 3563 1360
rect 3711 1356 3715 1360
rect 3839 1356 3843 1360
rect 3943 1353 3947 1357
rect 2047 1336 2051 1340
rect 2399 1337 2403 1341
rect 2535 1337 2539 1341
rect 2679 1337 2683 1341
rect 2823 1337 2827 1341
rect 2967 1337 2971 1341
rect 3111 1337 3115 1341
rect 3255 1337 3259 1341
rect 3407 1337 3411 1341
rect 3559 1337 3563 1341
rect 3711 1337 3715 1341
rect 3839 1337 3843 1341
rect 3943 1336 3947 1340
rect 111 1321 115 1325
rect 655 1324 659 1328
rect 767 1324 771 1328
rect 887 1324 891 1328
rect 1015 1324 1019 1328
rect 1143 1324 1147 1328
rect 1279 1324 1283 1328
rect 1415 1324 1419 1328
rect 1559 1324 1563 1328
rect 1703 1324 1707 1328
rect 1847 1324 1851 1328
rect 2007 1321 2011 1325
rect 111 1304 115 1308
rect 655 1305 659 1309
rect 767 1305 771 1309
rect 887 1305 891 1309
rect 1015 1305 1019 1309
rect 1143 1305 1147 1309
rect 1279 1305 1283 1309
rect 1415 1305 1419 1309
rect 1559 1305 1563 1309
rect 1703 1305 1707 1309
rect 1847 1305 1851 1309
rect 2007 1304 2011 1308
rect 2047 1280 2051 1284
rect 2247 1279 2251 1283
rect 2375 1279 2379 1283
rect 2511 1279 2515 1283
rect 2647 1279 2651 1283
rect 2791 1279 2795 1283
rect 2943 1279 2947 1283
rect 3111 1279 3115 1283
rect 3287 1279 3291 1283
rect 3471 1279 3475 1283
rect 3663 1279 3667 1283
rect 3839 1279 3843 1283
rect 3943 1280 3947 1284
rect 2047 1263 2051 1267
rect 2247 1260 2251 1264
rect 2375 1260 2379 1264
rect 2511 1260 2515 1264
rect 2647 1260 2651 1264
rect 2791 1260 2795 1264
rect 2943 1260 2947 1264
rect 3111 1260 3115 1264
rect 3287 1260 3291 1264
rect 3471 1260 3475 1264
rect 3663 1260 3667 1264
rect 3839 1260 3843 1264
rect 3943 1263 3947 1267
rect 111 1248 115 1252
rect 439 1247 443 1251
rect 551 1247 555 1251
rect 671 1247 675 1251
rect 799 1247 803 1251
rect 935 1247 939 1251
rect 1079 1247 1083 1251
rect 1231 1247 1235 1251
rect 1391 1247 1395 1251
rect 1551 1247 1555 1251
rect 1719 1247 1723 1251
rect 2007 1248 2011 1252
rect 111 1231 115 1235
rect 439 1228 443 1232
rect 551 1228 555 1232
rect 671 1228 675 1232
rect 799 1228 803 1232
rect 935 1228 939 1232
rect 1079 1228 1083 1232
rect 1231 1228 1235 1232
rect 1391 1228 1395 1232
rect 1551 1228 1555 1232
rect 1719 1228 1723 1232
rect 2007 1231 2011 1235
rect 2047 1193 2051 1197
rect 2071 1196 2075 1200
rect 2183 1196 2187 1200
rect 2303 1196 2307 1200
rect 2431 1196 2435 1200
rect 2559 1196 2563 1200
rect 2711 1196 2715 1200
rect 2887 1196 2891 1200
rect 3087 1196 3091 1200
rect 3311 1196 3315 1200
rect 3543 1196 3547 1200
rect 3783 1196 3787 1200
rect 3943 1193 3947 1197
rect 2047 1176 2051 1180
rect 2071 1177 2075 1181
rect 2183 1177 2187 1181
rect 2303 1177 2307 1181
rect 2431 1177 2435 1181
rect 2559 1177 2563 1181
rect 2711 1177 2715 1181
rect 2887 1177 2891 1181
rect 3087 1177 3091 1181
rect 3311 1177 3315 1181
rect 3543 1177 3547 1181
rect 3783 1177 3787 1181
rect 3943 1176 3947 1180
rect 111 1165 115 1169
rect 167 1168 171 1172
rect 303 1168 307 1172
rect 463 1168 467 1172
rect 631 1168 635 1172
rect 807 1168 811 1172
rect 983 1168 987 1172
rect 1159 1168 1163 1172
rect 1335 1168 1339 1172
rect 1511 1168 1515 1172
rect 1695 1168 1699 1172
rect 2007 1165 2011 1169
rect 111 1148 115 1152
rect 167 1149 171 1153
rect 303 1149 307 1153
rect 463 1149 467 1153
rect 631 1149 635 1153
rect 807 1149 811 1153
rect 983 1149 987 1153
rect 1159 1149 1163 1153
rect 1335 1149 1339 1153
rect 1511 1149 1515 1153
rect 1695 1149 1699 1153
rect 2007 1148 2011 1152
rect 2047 1120 2051 1124
rect 2071 1119 2075 1123
rect 2199 1119 2203 1123
rect 2351 1119 2355 1123
rect 2511 1119 2515 1123
rect 2679 1119 2683 1123
rect 2871 1119 2875 1123
rect 3087 1119 3091 1123
rect 3319 1119 3323 1123
rect 3559 1119 3563 1123
rect 3807 1119 3811 1123
rect 3943 1120 3947 1124
rect 2047 1103 2051 1107
rect 2071 1100 2075 1104
rect 2199 1100 2203 1104
rect 2351 1100 2355 1104
rect 2511 1100 2515 1104
rect 2679 1100 2683 1104
rect 2871 1100 2875 1104
rect 3087 1100 3091 1104
rect 3319 1100 3323 1104
rect 3559 1100 3563 1104
rect 3807 1100 3811 1104
rect 3943 1103 3947 1107
rect 111 1092 115 1096
rect 135 1091 139 1095
rect 239 1091 243 1095
rect 375 1091 379 1095
rect 527 1091 531 1095
rect 695 1091 699 1095
rect 863 1091 867 1095
rect 1039 1091 1043 1095
rect 1215 1091 1219 1095
rect 1391 1091 1395 1095
rect 1567 1091 1571 1095
rect 1743 1091 1747 1095
rect 1903 1091 1907 1095
rect 2007 1092 2011 1096
rect 111 1075 115 1079
rect 135 1072 139 1076
rect 239 1072 243 1076
rect 375 1072 379 1076
rect 527 1072 531 1076
rect 695 1072 699 1076
rect 863 1072 867 1076
rect 1039 1072 1043 1076
rect 1215 1072 1219 1076
rect 1391 1072 1395 1076
rect 1567 1072 1571 1076
rect 1743 1072 1747 1076
rect 1903 1072 1907 1076
rect 2007 1075 2011 1079
rect 2047 1025 2051 1029
rect 2071 1028 2075 1032
rect 2263 1028 2267 1032
rect 2487 1028 2491 1032
rect 2703 1028 2707 1032
rect 2919 1028 2923 1032
rect 3119 1028 3123 1032
rect 3311 1028 3315 1032
rect 3495 1028 3499 1032
rect 3679 1028 3683 1032
rect 3839 1028 3843 1032
rect 3943 1025 3947 1029
rect 111 1009 115 1013
rect 135 1012 139 1016
rect 287 1012 291 1016
rect 471 1012 475 1016
rect 655 1012 659 1016
rect 839 1012 843 1016
rect 1015 1012 1019 1016
rect 1199 1012 1203 1016
rect 1383 1012 1387 1016
rect 1567 1012 1571 1016
rect 2007 1009 2011 1013
rect 2047 1008 2051 1012
rect 2071 1009 2075 1013
rect 2263 1009 2267 1013
rect 2487 1009 2491 1013
rect 2703 1009 2707 1013
rect 2919 1009 2923 1013
rect 3119 1009 3123 1013
rect 3311 1009 3315 1013
rect 3495 1009 3499 1013
rect 3679 1009 3683 1013
rect 3839 1009 3843 1013
rect 3943 1008 3947 1012
rect 111 992 115 996
rect 135 993 139 997
rect 287 993 291 997
rect 471 993 475 997
rect 655 993 659 997
rect 839 993 843 997
rect 1015 993 1019 997
rect 1199 993 1203 997
rect 1383 993 1387 997
rect 1567 993 1571 997
rect 2007 992 2011 996
rect 2047 952 2051 956
rect 2303 951 2307 955
rect 2455 951 2459 955
rect 2615 951 2619 955
rect 2783 951 2787 955
rect 2951 951 2955 955
rect 3111 951 3115 955
rect 3263 951 3267 955
rect 3415 951 3419 955
rect 3559 951 3563 955
rect 3711 951 3715 955
rect 3839 951 3843 955
rect 3943 952 3947 956
rect 111 936 115 940
rect 135 935 139 939
rect 295 935 299 939
rect 471 935 475 939
rect 639 935 643 939
rect 799 935 803 939
rect 951 935 955 939
rect 1087 935 1091 939
rect 1223 935 1227 939
rect 1359 935 1363 939
rect 1495 935 1499 939
rect 2007 936 2011 940
rect 2047 935 2051 939
rect 2303 932 2307 936
rect 2455 932 2459 936
rect 2615 932 2619 936
rect 2783 932 2787 936
rect 2951 932 2955 936
rect 3111 932 3115 936
rect 3263 932 3267 936
rect 3415 932 3419 936
rect 3559 932 3563 936
rect 3711 932 3715 936
rect 3839 932 3843 936
rect 3943 935 3947 939
rect 111 919 115 923
rect 135 916 139 920
rect 295 916 299 920
rect 471 916 475 920
rect 639 916 643 920
rect 799 916 803 920
rect 951 916 955 920
rect 1087 916 1091 920
rect 1223 916 1227 920
rect 1359 916 1363 920
rect 1495 916 1499 920
rect 2007 919 2011 923
rect 2047 865 2051 869
rect 2559 868 2563 872
rect 2679 868 2683 872
rect 2807 868 2811 872
rect 2943 868 2947 872
rect 3079 868 3083 872
rect 3207 868 3211 872
rect 3335 868 3339 872
rect 3463 868 3467 872
rect 3591 868 3595 872
rect 3727 868 3731 872
rect 3839 868 3843 872
rect 3943 865 3947 869
rect 111 853 115 857
rect 159 856 163 860
rect 319 856 323 860
rect 471 856 475 860
rect 615 856 619 860
rect 751 856 755 860
rect 879 856 883 860
rect 999 856 1003 860
rect 1111 856 1115 860
rect 1231 856 1235 860
rect 1351 856 1355 860
rect 2007 853 2011 857
rect 2047 848 2051 852
rect 2559 849 2563 853
rect 2679 849 2683 853
rect 2807 849 2811 853
rect 2943 849 2947 853
rect 3079 849 3083 853
rect 3207 849 3211 853
rect 3335 849 3339 853
rect 3463 849 3467 853
rect 3591 849 3595 853
rect 3727 849 3731 853
rect 3839 849 3843 853
rect 3943 848 3947 852
rect 111 836 115 840
rect 159 837 163 841
rect 319 837 323 841
rect 471 837 475 841
rect 615 837 619 841
rect 751 837 755 841
rect 879 837 883 841
rect 999 837 1003 841
rect 1111 837 1115 841
rect 1231 837 1235 841
rect 1351 837 1355 841
rect 2007 836 2011 840
rect 2047 792 2051 796
rect 2335 791 2339 795
rect 2471 791 2475 795
rect 2615 791 2619 795
rect 2767 791 2771 795
rect 2919 791 2923 795
rect 3079 791 3083 795
rect 3239 791 3243 795
rect 3391 791 3395 795
rect 3543 791 3547 795
rect 3703 791 3707 795
rect 3839 791 3843 795
rect 3943 792 3947 796
rect 111 784 115 788
rect 223 783 227 787
rect 383 783 387 787
rect 535 783 539 787
rect 679 783 683 787
rect 815 783 819 787
rect 951 783 955 787
rect 1079 783 1083 787
rect 1199 783 1203 787
rect 1327 783 1331 787
rect 1455 783 1459 787
rect 2007 784 2011 788
rect 2047 775 2051 779
rect 2335 772 2339 776
rect 111 767 115 771
rect 2471 772 2475 776
rect 2615 772 2619 776
rect 2767 772 2771 776
rect 2919 772 2923 776
rect 3079 772 3083 776
rect 3239 772 3243 776
rect 3391 772 3395 776
rect 3543 772 3547 776
rect 3703 772 3707 776
rect 3839 772 3843 776
rect 3943 775 3947 779
rect 223 764 227 768
rect 383 764 387 768
rect 535 764 539 768
rect 679 764 683 768
rect 815 764 819 768
rect 951 764 955 768
rect 1079 764 1083 768
rect 1199 764 1203 768
rect 1327 764 1331 768
rect 1455 764 1459 768
rect 2007 767 2011 771
rect 2047 705 2051 709
rect 2071 708 2075 712
rect 2183 708 2187 712
rect 2335 708 2339 712
rect 2487 708 2491 712
rect 2639 708 2643 712
rect 2807 708 2811 712
rect 2983 708 2987 712
rect 3167 708 3171 712
rect 3367 708 3371 712
rect 3575 708 3579 712
rect 3783 708 3787 712
rect 111 697 115 701
rect 311 700 315 704
rect 471 700 475 704
rect 639 700 643 704
rect 807 700 811 704
rect 975 700 979 704
rect 1135 700 1139 704
rect 1295 700 1299 704
rect 1455 700 1459 704
rect 1607 700 1611 704
rect 1767 700 1771 704
rect 3943 705 3947 709
rect 1903 700 1907 704
rect 2007 697 2011 701
rect 2047 688 2051 692
rect 2071 689 2075 693
rect 2183 689 2187 693
rect 2335 689 2339 693
rect 2487 689 2491 693
rect 2639 689 2643 693
rect 2807 689 2811 693
rect 2983 689 2987 693
rect 3167 689 3171 693
rect 3367 689 3371 693
rect 3575 689 3579 693
rect 3783 689 3787 693
rect 3943 688 3947 692
rect 111 680 115 684
rect 311 681 315 685
rect 471 681 475 685
rect 639 681 643 685
rect 807 681 811 685
rect 975 681 979 685
rect 1135 681 1139 685
rect 1295 681 1299 685
rect 1455 681 1459 685
rect 1607 681 1611 685
rect 1767 681 1771 685
rect 1903 681 1907 685
rect 2007 680 2011 684
rect 111 628 115 632
rect 295 627 299 631
rect 447 627 451 631
rect 615 627 619 631
rect 783 627 787 631
rect 951 627 955 631
rect 1111 627 1115 631
rect 1263 627 1267 631
rect 1399 627 1403 631
rect 1535 627 1539 631
rect 1663 627 1667 631
rect 1791 627 1795 631
rect 1903 627 1907 631
rect 2007 628 2011 632
rect 2047 624 2051 628
rect 2071 623 2075 627
rect 2239 623 2243 627
rect 2423 623 2427 627
rect 2623 623 2627 627
rect 2839 623 2843 627
rect 3071 623 3075 627
rect 3319 623 3323 627
rect 3575 623 3579 627
rect 3839 623 3843 627
rect 3943 624 3947 628
rect 111 611 115 615
rect 295 608 299 612
rect 447 608 451 612
rect 615 608 619 612
rect 783 608 787 612
rect 951 608 955 612
rect 1111 608 1115 612
rect 1263 608 1267 612
rect 1399 608 1403 612
rect 1535 608 1539 612
rect 1663 608 1667 612
rect 1791 608 1795 612
rect 1903 608 1907 612
rect 2007 611 2011 615
rect 2047 607 2051 611
rect 2071 604 2075 608
rect 2239 604 2243 608
rect 2423 604 2427 608
rect 2623 604 2627 608
rect 2839 604 2843 608
rect 3071 604 3075 608
rect 3319 604 3323 608
rect 3575 604 3579 608
rect 3839 604 3843 608
rect 3943 607 3947 611
rect 111 541 115 545
rect 239 544 243 548
rect 415 544 419 548
rect 607 544 611 548
rect 799 544 803 548
rect 991 544 995 548
rect 1175 544 1179 548
rect 1351 544 1355 548
rect 1519 544 1523 548
rect 1687 544 1691 548
rect 1863 544 1867 548
rect 2007 541 2011 545
rect 2047 541 2051 545
rect 2191 544 2195 548
rect 2287 544 2291 548
rect 2383 544 2387 548
rect 2479 544 2483 548
rect 2583 544 2587 548
rect 2711 544 2715 548
rect 2871 544 2875 548
rect 3071 544 3075 548
rect 3303 544 3307 548
rect 3551 544 3555 548
rect 3807 544 3811 548
rect 3943 541 3947 545
rect 111 524 115 528
rect 239 525 243 529
rect 415 525 419 529
rect 607 525 611 529
rect 799 525 803 529
rect 991 525 995 529
rect 1175 525 1179 529
rect 1351 525 1355 529
rect 1519 525 1523 529
rect 1687 525 1691 529
rect 1863 525 1867 529
rect 2007 524 2011 528
rect 2047 524 2051 528
rect 2191 525 2195 529
rect 2287 525 2291 529
rect 2383 525 2387 529
rect 2479 525 2483 529
rect 2583 525 2587 529
rect 2711 525 2715 529
rect 2871 525 2875 529
rect 3071 525 3075 529
rect 3303 525 3307 529
rect 3551 525 3555 529
rect 3807 525 3811 529
rect 3943 524 3947 528
rect 111 472 115 476
rect 135 471 139 475
rect 287 471 291 475
rect 463 471 467 475
rect 639 471 643 475
rect 807 471 811 475
rect 967 471 971 475
rect 1119 471 1123 475
rect 1271 471 1275 475
rect 1415 471 1419 475
rect 1567 471 1571 475
rect 2007 472 2011 476
rect 2047 472 2051 476
rect 2431 471 2435 475
rect 2527 471 2531 475
rect 2623 471 2627 475
rect 2727 471 2731 475
rect 2847 471 2851 475
rect 2999 471 3003 475
rect 3175 471 3179 475
rect 3375 471 3379 475
rect 3591 471 3595 475
rect 3807 471 3811 475
rect 3943 472 3947 476
rect 111 455 115 459
rect 135 452 139 456
rect 287 452 291 456
rect 463 452 467 456
rect 639 452 643 456
rect 807 452 811 456
rect 967 452 971 456
rect 1119 452 1123 456
rect 1271 452 1275 456
rect 1415 452 1419 456
rect 1567 452 1571 456
rect 2007 455 2011 459
rect 2047 455 2051 459
rect 2431 452 2435 456
rect 2527 452 2531 456
rect 2623 452 2627 456
rect 2727 452 2731 456
rect 2847 452 2851 456
rect 2999 452 3003 456
rect 3175 452 3179 456
rect 3375 452 3379 456
rect 3591 452 3595 456
rect 3807 452 3811 456
rect 3943 455 3947 459
rect 111 385 115 389
rect 135 388 139 392
rect 279 388 283 392
rect 439 388 443 392
rect 583 388 587 392
rect 719 388 723 392
rect 847 388 851 392
rect 967 388 971 392
rect 1087 388 1091 392
rect 1207 388 1211 392
rect 1327 388 1331 392
rect 2007 385 2011 389
rect 2047 389 2051 393
rect 2431 392 2435 396
rect 2527 392 2531 396
rect 2623 392 2627 396
rect 2719 392 2723 396
rect 2815 392 2819 396
rect 2927 392 2931 396
rect 3063 392 3067 396
rect 3223 392 3227 396
rect 3399 392 3403 396
rect 3591 392 3595 396
rect 3783 392 3787 396
rect 3943 389 3947 393
rect 111 368 115 372
rect 135 369 139 373
rect 279 369 283 373
rect 439 369 443 373
rect 583 369 587 373
rect 719 369 723 373
rect 847 369 851 373
rect 967 369 971 373
rect 1087 369 1091 373
rect 1207 369 1211 373
rect 1327 369 1331 373
rect 2007 368 2011 372
rect 2047 372 2051 376
rect 2431 373 2435 377
rect 2527 373 2531 377
rect 2623 373 2627 377
rect 2719 373 2723 377
rect 2815 373 2819 377
rect 2927 373 2931 377
rect 3063 373 3067 377
rect 3223 373 3227 377
rect 3399 373 3403 377
rect 3591 373 3595 377
rect 3783 373 3787 377
rect 3943 372 3947 376
rect 111 316 115 320
rect 143 315 147 319
rect 319 315 323 319
rect 479 315 483 319
rect 631 315 635 319
rect 775 315 779 319
rect 903 315 907 319
rect 1031 315 1035 319
rect 1151 315 1155 319
rect 1271 315 1275 319
rect 1391 315 1395 319
rect 2007 316 2011 320
rect 2047 316 2051 320
rect 2191 315 2195 319
rect 2327 315 2331 319
rect 2471 315 2475 319
rect 2623 315 2627 319
rect 2783 315 2787 319
rect 2951 315 2955 319
rect 3119 315 3123 319
rect 3295 315 3299 319
rect 3471 315 3475 319
rect 3655 315 3659 319
rect 3839 315 3843 319
rect 3943 316 3947 320
rect 111 299 115 303
rect 143 296 147 300
rect 319 296 323 300
rect 479 296 483 300
rect 631 296 635 300
rect 775 296 779 300
rect 903 296 907 300
rect 1031 296 1035 300
rect 1151 296 1155 300
rect 1271 296 1275 300
rect 1391 296 1395 300
rect 2007 299 2011 303
rect 2047 299 2051 303
rect 2191 296 2195 300
rect 2327 296 2331 300
rect 2471 296 2475 300
rect 2623 296 2627 300
rect 2783 296 2787 300
rect 2951 296 2955 300
rect 3119 296 3123 300
rect 3295 296 3299 300
rect 3471 296 3475 300
rect 3655 296 3659 300
rect 3839 296 3843 300
rect 3943 299 3947 303
rect 111 229 115 233
rect 223 232 227 236
rect 391 232 395 236
rect 559 232 563 236
rect 735 232 739 236
rect 903 232 907 236
rect 1063 232 1067 236
rect 1215 232 1219 236
rect 1359 232 1363 236
rect 1511 232 1515 236
rect 1663 232 1667 236
rect 2007 229 2011 233
rect 2047 233 2051 237
rect 2071 236 2075 240
rect 2215 236 2219 240
rect 2399 236 2403 240
rect 2591 236 2595 240
rect 2791 236 2795 240
rect 2983 236 2987 240
rect 3167 236 3171 240
rect 3343 236 3347 240
rect 3511 236 3515 240
rect 3687 236 3691 240
rect 3839 236 3843 240
rect 3943 233 3947 237
rect 111 212 115 216
rect 223 213 227 217
rect 391 213 395 217
rect 559 213 563 217
rect 735 213 739 217
rect 903 213 907 217
rect 1063 213 1067 217
rect 1215 213 1219 217
rect 1359 213 1363 217
rect 1511 213 1515 217
rect 1663 213 1667 217
rect 2007 212 2011 216
rect 2047 216 2051 220
rect 2071 217 2075 221
rect 2215 217 2219 221
rect 2399 217 2403 221
rect 2591 217 2595 221
rect 2791 217 2795 221
rect 2983 217 2987 221
rect 3167 217 3171 221
rect 3343 217 3347 221
rect 3511 217 3515 221
rect 3687 217 3691 221
rect 3839 217 3843 221
rect 3943 216 3947 220
rect 2047 140 2051 144
rect 2071 139 2075 143
rect 2191 139 2195 143
rect 2343 139 2347 143
rect 2495 139 2499 143
rect 2647 139 2651 143
rect 2799 139 2803 143
rect 2943 139 2947 143
rect 3071 139 3075 143
rect 3191 139 3195 143
rect 3311 139 3315 143
rect 3423 139 3427 143
rect 3527 139 3531 143
rect 3639 139 3643 143
rect 3743 139 3747 143
rect 3839 139 3843 143
rect 3943 140 3947 144
rect 111 128 115 132
rect 151 127 155 131
rect 247 127 251 131
rect 343 127 347 131
rect 439 127 443 131
rect 535 127 539 131
rect 631 127 635 131
rect 727 127 731 131
rect 823 127 827 131
rect 919 127 923 131
rect 1015 127 1019 131
rect 1111 127 1115 131
rect 1207 127 1211 131
rect 1303 127 1307 131
rect 1407 127 1411 131
rect 1511 127 1515 131
rect 1615 127 1619 131
rect 1711 127 1715 131
rect 1807 127 1811 131
rect 1903 127 1907 131
rect 2007 128 2011 132
rect 2047 123 2051 127
rect 2071 120 2075 124
rect 2191 120 2195 124
rect 2343 120 2347 124
rect 2495 120 2499 124
rect 2647 120 2651 124
rect 2799 120 2803 124
rect 2943 120 2947 124
rect 3071 120 3075 124
rect 3191 120 3195 124
rect 3311 120 3315 124
rect 3423 120 3427 124
rect 3527 120 3531 124
rect 3639 120 3643 124
rect 3743 120 3747 124
rect 3839 120 3843 124
rect 3943 123 3947 127
rect 111 111 115 115
rect 151 108 155 112
rect 247 108 251 112
rect 343 108 347 112
rect 439 108 443 112
rect 535 108 539 112
rect 631 108 635 112
rect 727 108 731 112
rect 823 108 827 112
rect 919 108 923 112
rect 1015 108 1019 112
rect 1111 108 1115 112
rect 1207 108 1211 112
rect 1303 108 1307 112
rect 1407 108 1411 112
rect 1511 108 1515 112
rect 1615 108 1619 112
rect 1711 108 1715 112
rect 1807 108 1811 112
rect 1903 108 1907 112
rect 2007 111 2011 115
<< m3 >>
rect 2047 4022 2051 4023
rect 2047 4017 2051 4018
rect 2071 4022 2075 4023
rect 2071 4017 2075 4018
rect 2327 4022 2331 4023
rect 2327 4017 2331 4018
rect 2591 4022 2595 4023
rect 2591 4017 2595 4018
rect 2839 4022 2843 4023
rect 2839 4017 2843 4018
rect 3087 4022 3091 4023
rect 3087 4017 3091 4018
rect 3343 4022 3347 4023
rect 3343 4017 3347 4018
rect 3943 4022 3947 4023
rect 3943 4017 3947 4018
rect 111 4002 115 4003
rect 111 3997 115 3998
rect 311 4002 315 4003
rect 311 3997 315 3998
rect 511 4002 515 4003
rect 511 3997 515 3998
rect 703 4002 707 4003
rect 703 3997 707 3998
rect 887 4002 891 4003
rect 887 3997 891 3998
rect 1063 4002 1067 4003
rect 1063 3997 1067 3998
rect 1231 4002 1235 4003
rect 1231 3997 1235 3998
rect 1383 4002 1387 4003
rect 1383 3997 1387 3998
rect 1519 4002 1523 4003
rect 1519 3997 1523 3998
rect 1655 4002 1659 4003
rect 1655 3997 1659 3998
rect 1791 4002 1795 4003
rect 1791 3997 1795 3998
rect 1903 4002 1907 4003
rect 1903 3997 1907 3998
rect 2007 4002 2011 4003
rect 2007 3997 2011 3998
rect 112 3970 114 3997
rect 312 3973 314 3997
rect 512 3973 514 3997
rect 704 3973 706 3997
rect 888 3973 890 3997
rect 1064 3973 1066 3997
rect 1232 3973 1234 3997
rect 1384 3973 1386 3997
rect 1520 3973 1522 3997
rect 1656 3973 1658 3997
rect 1792 3973 1794 3997
rect 1904 3973 1906 3997
rect 310 3972 316 3973
rect 110 3969 116 3970
rect 110 3965 111 3969
rect 115 3965 116 3969
rect 310 3968 311 3972
rect 315 3968 316 3972
rect 310 3967 316 3968
rect 510 3972 516 3973
rect 510 3968 511 3972
rect 515 3968 516 3972
rect 510 3967 516 3968
rect 702 3972 708 3973
rect 702 3968 703 3972
rect 707 3968 708 3972
rect 702 3967 708 3968
rect 886 3972 892 3973
rect 886 3968 887 3972
rect 891 3968 892 3972
rect 886 3967 892 3968
rect 1062 3972 1068 3973
rect 1062 3968 1063 3972
rect 1067 3968 1068 3972
rect 1062 3967 1068 3968
rect 1230 3972 1236 3973
rect 1230 3968 1231 3972
rect 1235 3968 1236 3972
rect 1230 3967 1236 3968
rect 1382 3972 1388 3973
rect 1382 3968 1383 3972
rect 1387 3968 1388 3972
rect 1382 3967 1388 3968
rect 1518 3972 1524 3973
rect 1518 3968 1519 3972
rect 1523 3968 1524 3972
rect 1518 3967 1524 3968
rect 1654 3972 1660 3973
rect 1654 3968 1655 3972
rect 1659 3968 1660 3972
rect 1654 3967 1660 3968
rect 1790 3972 1796 3973
rect 1790 3968 1791 3972
rect 1795 3968 1796 3972
rect 1790 3967 1796 3968
rect 1902 3972 1908 3973
rect 1902 3968 1903 3972
rect 1907 3968 1908 3972
rect 2008 3970 2010 3997
rect 2048 3990 2050 4017
rect 2072 3993 2074 4017
rect 2328 3993 2330 4017
rect 2592 3993 2594 4017
rect 2840 3993 2842 4017
rect 3088 3993 3090 4017
rect 3344 3993 3346 4017
rect 2070 3992 2076 3993
rect 2046 3989 2052 3990
rect 2046 3985 2047 3989
rect 2051 3985 2052 3989
rect 2070 3988 2071 3992
rect 2075 3988 2076 3992
rect 2070 3987 2076 3988
rect 2326 3992 2332 3993
rect 2326 3988 2327 3992
rect 2331 3988 2332 3992
rect 2326 3987 2332 3988
rect 2590 3992 2596 3993
rect 2590 3988 2591 3992
rect 2595 3988 2596 3992
rect 2590 3987 2596 3988
rect 2838 3992 2844 3993
rect 2838 3988 2839 3992
rect 2843 3988 2844 3992
rect 2838 3987 2844 3988
rect 3086 3992 3092 3993
rect 3086 3988 3087 3992
rect 3091 3988 3092 3992
rect 3086 3987 3092 3988
rect 3342 3992 3348 3993
rect 3342 3988 3343 3992
rect 3347 3988 3348 3992
rect 3944 3990 3946 4017
rect 3342 3987 3348 3988
rect 3942 3989 3948 3990
rect 2046 3984 2052 3985
rect 3942 3985 3943 3989
rect 3947 3985 3948 3989
rect 3942 3984 3948 3985
rect 2070 3973 2076 3974
rect 2046 3972 2052 3973
rect 1902 3967 1908 3968
rect 2006 3969 2012 3970
rect 110 3964 116 3965
rect 2006 3965 2007 3969
rect 2011 3965 2012 3969
rect 2046 3968 2047 3972
rect 2051 3968 2052 3972
rect 2070 3969 2071 3973
rect 2075 3969 2076 3973
rect 2070 3968 2076 3969
rect 2326 3973 2332 3974
rect 2326 3969 2327 3973
rect 2331 3969 2332 3973
rect 2326 3968 2332 3969
rect 2590 3973 2596 3974
rect 2590 3969 2591 3973
rect 2595 3969 2596 3973
rect 2590 3968 2596 3969
rect 2838 3973 2844 3974
rect 2838 3969 2839 3973
rect 2843 3969 2844 3973
rect 2838 3968 2844 3969
rect 3086 3973 3092 3974
rect 3086 3969 3087 3973
rect 3091 3969 3092 3973
rect 3086 3968 3092 3969
rect 3342 3973 3348 3974
rect 3342 3969 3343 3973
rect 3347 3969 3348 3973
rect 3342 3968 3348 3969
rect 3942 3972 3948 3973
rect 3942 3968 3943 3972
rect 3947 3968 3948 3972
rect 2046 3967 2052 3968
rect 2006 3964 2012 3965
rect 310 3953 316 3954
rect 110 3952 116 3953
rect 110 3948 111 3952
rect 115 3948 116 3952
rect 310 3949 311 3953
rect 315 3949 316 3953
rect 310 3948 316 3949
rect 510 3953 516 3954
rect 510 3949 511 3953
rect 515 3949 516 3953
rect 510 3948 516 3949
rect 702 3953 708 3954
rect 702 3949 703 3953
rect 707 3949 708 3953
rect 702 3948 708 3949
rect 886 3953 892 3954
rect 886 3949 887 3953
rect 891 3949 892 3953
rect 886 3948 892 3949
rect 1062 3953 1068 3954
rect 1062 3949 1063 3953
rect 1067 3949 1068 3953
rect 1062 3948 1068 3949
rect 1230 3953 1236 3954
rect 1230 3949 1231 3953
rect 1235 3949 1236 3953
rect 1230 3948 1236 3949
rect 1382 3953 1388 3954
rect 1382 3949 1383 3953
rect 1387 3949 1388 3953
rect 1382 3948 1388 3949
rect 1518 3953 1524 3954
rect 1518 3949 1519 3953
rect 1523 3949 1524 3953
rect 1518 3948 1524 3949
rect 1654 3953 1660 3954
rect 1654 3949 1655 3953
rect 1659 3949 1660 3953
rect 1654 3948 1660 3949
rect 1790 3953 1796 3954
rect 1790 3949 1791 3953
rect 1795 3949 1796 3953
rect 1790 3948 1796 3949
rect 1902 3953 1908 3954
rect 1902 3949 1903 3953
rect 1907 3949 1908 3953
rect 1902 3948 1908 3949
rect 2006 3952 2012 3953
rect 2006 3948 2007 3952
rect 2011 3948 2012 3952
rect 110 3947 116 3948
rect 112 3927 114 3947
rect 312 3927 314 3948
rect 512 3927 514 3948
rect 704 3927 706 3948
rect 888 3927 890 3948
rect 1064 3927 1066 3948
rect 1232 3927 1234 3948
rect 1384 3927 1386 3948
rect 1520 3927 1522 3948
rect 1656 3927 1658 3948
rect 1792 3927 1794 3948
rect 1904 3927 1906 3948
rect 2006 3947 2012 3948
rect 2048 3947 2050 3967
rect 2072 3947 2074 3968
rect 2328 3947 2330 3968
rect 2592 3947 2594 3968
rect 2840 3947 2842 3968
rect 3088 3947 3090 3968
rect 3344 3947 3346 3968
rect 3942 3967 3948 3968
rect 3944 3947 3946 3967
rect 2008 3927 2010 3947
rect 2047 3946 2051 3947
rect 2047 3941 2051 3942
rect 2071 3946 2075 3947
rect 2071 3941 2075 3942
rect 2127 3946 2131 3947
rect 2127 3941 2131 3942
rect 2271 3946 2275 3947
rect 2271 3941 2275 3942
rect 2327 3946 2331 3947
rect 2327 3941 2331 3942
rect 2439 3946 2443 3947
rect 2439 3941 2443 3942
rect 2591 3946 2595 3947
rect 2591 3941 2595 3942
rect 2615 3946 2619 3947
rect 2615 3941 2619 3942
rect 2799 3946 2803 3947
rect 2799 3941 2803 3942
rect 2839 3946 2843 3947
rect 2839 3941 2843 3942
rect 2983 3946 2987 3947
rect 2983 3941 2987 3942
rect 3087 3946 3091 3947
rect 3087 3941 3091 3942
rect 3175 3946 3179 3947
rect 3175 3941 3179 3942
rect 3343 3946 3347 3947
rect 3343 3941 3347 3942
rect 3367 3946 3371 3947
rect 3367 3941 3371 3942
rect 3559 3946 3563 3947
rect 3559 3941 3563 3942
rect 3943 3946 3947 3947
rect 3943 3941 3947 3942
rect 111 3926 115 3927
rect 111 3921 115 3922
rect 279 3926 283 3927
rect 279 3921 283 3922
rect 311 3926 315 3927
rect 311 3921 315 3922
rect 415 3926 419 3927
rect 415 3921 419 3922
rect 511 3926 515 3927
rect 511 3921 515 3922
rect 567 3926 571 3927
rect 567 3921 571 3922
rect 703 3926 707 3927
rect 703 3921 707 3922
rect 735 3926 739 3927
rect 735 3921 739 3922
rect 887 3926 891 3927
rect 887 3921 891 3922
rect 911 3926 915 3927
rect 911 3921 915 3922
rect 1063 3926 1067 3927
rect 1063 3921 1067 3922
rect 1095 3926 1099 3927
rect 1095 3921 1099 3922
rect 1231 3926 1235 3927
rect 1231 3921 1235 3922
rect 1287 3926 1291 3927
rect 1287 3921 1291 3922
rect 1383 3926 1387 3927
rect 1383 3921 1387 3922
rect 1479 3926 1483 3927
rect 1479 3921 1483 3922
rect 1519 3926 1523 3927
rect 1519 3921 1523 3922
rect 1655 3926 1659 3927
rect 1655 3921 1659 3922
rect 1679 3926 1683 3927
rect 1679 3921 1683 3922
rect 1791 3926 1795 3927
rect 1791 3921 1795 3922
rect 1903 3926 1907 3927
rect 1903 3921 1907 3922
rect 2007 3926 2011 3927
rect 2007 3921 2011 3922
rect 2048 3921 2050 3941
rect 112 3901 114 3921
rect 110 3900 116 3901
rect 280 3900 282 3921
rect 416 3900 418 3921
rect 568 3900 570 3921
rect 736 3900 738 3921
rect 912 3900 914 3921
rect 1096 3900 1098 3921
rect 1288 3900 1290 3921
rect 1480 3900 1482 3921
rect 1680 3900 1682 3921
rect 2008 3901 2010 3921
rect 2046 3920 2052 3921
rect 2128 3920 2130 3941
rect 2272 3920 2274 3941
rect 2440 3920 2442 3941
rect 2616 3920 2618 3941
rect 2800 3920 2802 3941
rect 2984 3920 2986 3941
rect 3176 3920 3178 3941
rect 3368 3920 3370 3941
rect 3560 3920 3562 3941
rect 3944 3921 3946 3941
rect 3942 3920 3948 3921
rect 2046 3916 2047 3920
rect 2051 3916 2052 3920
rect 2046 3915 2052 3916
rect 2126 3919 2132 3920
rect 2126 3915 2127 3919
rect 2131 3915 2132 3919
rect 2126 3914 2132 3915
rect 2270 3919 2276 3920
rect 2270 3915 2271 3919
rect 2275 3915 2276 3919
rect 2270 3914 2276 3915
rect 2438 3919 2444 3920
rect 2438 3915 2439 3919
rect 2443 3915 2444 3919
rect 2438 3914 2444 3915
rect 2614 3919 2620 3920
rect 2614 3915 2615 3919
rect 2619 3915 2620 3919
rect 2614 3914 2620 3915
rect 2798 3919 2804 3920
rect 2798 3915 2799 3919
rect 2803 3915 2804 3919
rect 2798 3914 2804 3915
rect 2982 3919 2988 3920
rect 2982 3915 2983 3919
rect 2987 3915 2988 3919
rect 2982 3914 2988 3915
rect 3174 3919 3180 3920
rect 3174 3915 3175 3919
rect 3179 3915 3180 3919
rect 3174 3914 3180 3915
rect 3366 3919 3372 3920
rect 3366 3915 3367 3919
rect 3371 3915 3372 3919
rect 3366 3914 3372 3915
rect 3558 3919 3564 3920
rect 3558 3915 3559 3919
rect 3563 3915 3564 3919
rect 3942 3916 3943 3920
rect 3947 3916 3948 3920
rect 3942 3915 3948 3916
rect 3558 3914 3564 3915
rect 2046 3903 2052 3904
rect 2006 3900 2012 3901
rect 110 3896 111 3900
rect 115 3896 116 3900
rect 110 3895 116 3896
rect 278 3899 284 3900
rect 278 3895 279 3899
rect 283 3895 284 3899
rect 278 3894 284 3895
rect 414 3899 420 3900
rect 414 3895 415 3899
rect 419 3895 420 3899
rect 414 3894 420 3895
rect 566 3899 572 3900
rect 566 3895 567 3899
rect 571 3895 572 3899
rect 566 3894 572 3895
rect 734 3899 740 3900
rect 734 3895 735 3899
rect 739 3895 740 3899
rect 734 3894 740 3895
rect 910 3899 916 3900
rect 910 3895 911 3899
rect 915 3895 916 3899
rect 910 3894 916 3895
rect 1094 3899 1100 3900
rect 1094 3895 1095 3899
rect 1099 3895 1100 3899
rect 1094 3894 1100 3895
rect 1286 3899 1292 3900
rect 1286 3895 1287 3899
rect 1291 3895 1292 3899
rect 1286 3894 1292 3895
rect 1478 3899 1484 3900
rect 1478 3895 1479 3899
rect 1483 3895 1484 3899
rect 1478 3894 1484 3895
rect 1678 3899 1684 3900
rect 1678 3895 1679 3899
rect 1683 3895 1684 3899
rect 2006 3896 2007 3900
rect 2011 3896 2012 3900
rect 2046 3899 2047 3903
rect 2051 3899 2052 3903
rect 3942 3903 3948 3904
rect 2046 3898 2052 3899
rect 2126 3900 2132 3901
rect 2006 3895 2012 3896
rect 1678 3894 1684 3895
rect 110 3883 116 3884
rect 110 3879 111 3883
rect 115 3879 116 3883
rect 2006 3883 2012 3884
rect 110 3878 116 3879
rect 278 3880 284 3881
rect 112 3843 114 3878
rect 278 3876 279 3880
rect 283 3876 284 3880
rect 278 3875 284 3876
rect 414 3880 420 3881
rect 414 3876 415 3880
rect 419 3876 420 3880
rect 414 3875 420 3876
rect 566 3880 572 3881
rect 566 3876 567 3880
rect 571 3876 572 3880
rect 566 3875 572 3876
rect 734 3880 740 3881
rect 734 3876 735 3880
rect 739 3876 740 3880
rect 734 3875 740 3876
rect 910 3880 916 3881
rect 910 3876 911 3880
rect 915 3876 916 3880
rect 910 3875 916 3876
rect 1094 3880 1100 3881
rect 1094 3876 1095 3880
rect 1099 3876 1100 3880
rect 1094 3875 1100 3876
rect 1286 3880 1292 3881
rect 1286 3876 1287 3880
rect 1291 3876 1292 3880
rect 1286 3875 1292 3876
rect 1478 3880 1484 3881
rect 1478 3876 1479 3880
rect 1483 3876 1484 3880
rect 1478 3875 1484 3876
rect 1678 3880 1684 3881
rect 1678 3876 1679 3880
rect 1683 3876 1684 3880
rect 2006 3879 2007 3883
rect 2011 3879 2012 3883
rect 2006 3878 2012 3879
rect 1678 3875 1684 3876
rect 280 3843 282 3875
rect 416 3843 418 3875
rect 568 3843 570 3875
rect 736 3843 738 3875
rect 912 3843 914 3875
rect 1096 3843 1098 3875
rect 1288 3843 1290 3875
rect 1480 3843 1482 3875
rect 1680 3843 1682 3875
rect 2008 3843 2010 3878
rect 2048 3871 2050 3898
rect 2126 3896 2127 3900
rect 2131 3896 2132 3900
rect 2126 3895 2132 3896
rect 2270 3900 2276 3901
rect 2270 3896 2271 3900
rect 2275 3896 2276 3900
rect 2270 3895 2276 3896
rect 2438 3900 2444 3901
rect 2438 3896 2439 3900
rect 2443 3896 2444 3900
rect 2438 3895 2444 3896
rect 2614 3900 2620 3901
rect 2614 3896 2615 3900
rect 2619 3896 2620 3900
rect 2614 3895 2620 3896
rect 2798 3900 2804 3901
rect 2798 3896 2799 3900
rect 2803 3896 2804 3900
rect 2798 3895 2804 3896
rect 2982 3900 2988 3901
rect 2982 3896 2983 3900
rect 2987 3896 2988 3900
rect 2982 3895 2988 3896
rect 3174 3900 3180 3901
rect 3174 3896 3175 3900
rect 3179 3896 3180 3900
rect 3174 3895 3180 3896
rect 3366 3900 3372 3901
rect 3366 3896 3367 3900
rect 3371 3896 3372 3900
rect 3366 3895 3372 3896
rect 3558 3900 3564 3901
rect 3558 3896 3559 3900
rect 3563 3896 3564 3900
rect 3942 3899 3943 3903
rect 3947 3899 3948 3903
rect 3942 3898 3948 3899
rect 3558 3895 3564 3896
rect 2128 3871 2130 3895
rect 2272 3871 2274 3895
rect 2440 3871 2442 3895
rect 2616 3871 2618 3895
rect 2800 3871 2802 3895
rect 2984 3871 2986 3895
rect 3176 3871 3178 3895
rect 3368 3871 3370 3895
rect 3560 3871 3562 3895
rect 3944 3871 3946 3898
rect 2047 3870 2051 3871
rect 2047 3865 2051 3866
rect 2127 3870 2131 3871
rect 2127 3865 2131 3866
rect 2263 3870 2267 3871
rect 2263 3865 2267 3866
rect 2271 3870 2275 3871
rect 2271 3865 2275 3866
rect 2375 3870 2379 3871
rect 2375 3865 2379 3866
rect 2439 3870 2443 3871
rect 2439 3865 2443 3866
rect 2495 3870 2499 3871
rect 2495 3865 2499 3866
rect 2615 3870 2619 3871
rect 2615 3865 2619 3866
rect 2631 3870 2635 3871
rect 2631 3865 2635 3866
rect 2775 3870 2779 3871
rect 2775 3865 2779 3866
rect 2799 3870 2803 3871
rect 2799 3865 2803 3866
rect 2919 3870 2923 3871
rect 2919 3865 2923 3866
rect 2983 3870 2987 3871
rect 2983 3865 2987 3866
rect 3063 3870 3067 3871
rect 3063 3865 3067 3866
rect 3175 3870 3179 3871
rect 3175 3865 3179 3866
rect 3207 3870 3211 3871
rect 3207 3865 3211 3866
rect 3343 3870 3347 3871
rect 3343 3865 3347 3866
rect 3367 3870 3371 3871
rect 3367 3865 3371 3866
rect 3471 3870 3475 3871
rect 3471 3865 3475 3866
rect 3559 3870 3563 3871
rect 3559 3865 3563 3866
rect 3599 3870 3603 3871
rect 3599 3865 3603 3866
rect 3727 3870 3731 3871
rect 3727 3865 3731 3866
rect 3839 3870 3843 3871
rect 3839 3865 3843 3866
rect 3943 3870 3947 3871
rect 3943 3865 3947 3866
rect 111 3842 115 3843
rect 111 3837 115 3838
rect 231 3842 235 3843
rect 231 3837 235 3838
rect 279 3842 283 3843
rect 279 3837 283 3838
rect 335 3842 339 3843
rect 335 3837 339 3838
rect 415 3842 419 3843
rect 415 3837 419 3838
rect 439 3842 443 3843
rect 439 3837 443 3838
rect 535 3842 539 3843
rect 535 3837 539 3838
rect 567 3842 571 3843
rect 567 3837 571 3838
rect 631 3842 635 3843
rect 631 3837 635 3838
rect 727 3842 731 3843
rect 727 3837 731 3838
rect 735 3842 739 3843
rect 735 3837 739 3838
rect 831 3842 835 3843
rect 831 3837 835 3838
rect 911 3842 915 3843
rect 911 3837 915 3838
rect 935 3842 939 3843
rect 935 3837 939 3838
rect 1039 3842 1043 3843
rect 1039 3837 1043 3838
rect 1095 3842 1099 3843
rect 1095 3837 1099 3838
rect 1151 3842 1155 3843
rect 1151 3837 1155 3838
rect 1263 3842 1267 3843
rect 1263 3837 1267 3838
rect 1287 3842 1291 3843
rect 1287 3837 1291 3838
rect 1383 3842 1387 3843
rect 1383 3837 1387 3838
rect 1479 3842 1483 3843
rect 1479 3837 1483 3838
rect 1503 3842 1507 3843
rect 1503 3837 1507 3838
rect 1631 3842 1635 3843
rect 1631 3837 1635 3838
rect 1679 3842 1683 3843
rect 1679 3837 1683 3838
rect 2007 3842 2011 3843
rect 2048 3838 2050 3865
rect 2264 3841 2266 3865
rect 2376 3841 2378 3865
rect 2496 3841 2498 3865
rect 2632 3841 2634 3865
rect 2776 3841 2778 3865
rect 2920 3841 2922 3865
rect 3064 3841 3066 3865
rect 3208 3841 3210 3865
rect 3344 3841 3346 3865
rect 3472 3841 3474 3865
rect 3600 3841 3602 3865
rect 3728 3841 3730 3865
rect 3840 3841 3842 3865
rect 2262 3840 2268 3841
rect 2007 3837 2011 3838
rect 2046 3837 2052 3838
rect 112 3810 114 3837
rect 232 3813 234 3837
rect 336 3813 338 3837
rect 440 3813 442 3837
rect 536 3813 538 3837
rect 632 3813 634 3837
rect 728 3813 730 3837
rect 832 3813 834 3837
rect 936 3813 938 3837
rect 1040 3813 1042 3837
rect 1152 3813 1154 3837
rect 1264 3813 1266 3837
rect 1384 3813 1386 3837
rect 1504 3813 1506 3837
rect 1632 3813 1634 3837
rect 230 3812 236 3813
rect 110 3809 116 3810
rect 110 3805 111 3809
rect 115 3805 116 3809
rect 230 3808 231 3812
rect 235 3808 236 3812
rect 230 3807 236 3808
rect 334 3812 340 3813
rect 334 3808 335 3812
rect 339 3808 340 3812
rect 334 3807 340 3808
rect 438 3812 444 3813
rect 438 3808 439 3812
rect 443 3808 444 3812
rect 438 3807 444 3808
rect 534 3812 540 3813
rect 534 3808 535 3812
rect 539 3808 540 3812
rect 534 3807 540 3808
rect 630 3812 636 3813
rect 630 3808 631 3812
rect 635 3808 636 3812
rect 630 3807 636 3808
rect 726 3812 732 3813
rect 726 3808 727 3812
rect 731 3808 732 3812
rect 726 3807 732 3808
rect 830 3812 836 3813
rect 830 3808 831 3812
rect 835 3808 836 3812
rect 830 3807 836 3808
rect 934 3812 940 3813
rect 934 3808 935 3812
rect 939 3808 940 3812
rect 934 3807 940 3808
rect 1038 3812 1044 3813
rect 1038 3808 1039 3812
rect 1043 3808 1044 3812
rect 1038 3807 1044 3808
rect 1150 3812 1156 3813
rect 1150 3808 1151 3812
rect 1155 3808 1156 3812
rect 1150 3807 1156 3808
rect 1262 3812 1268 3813
rect 1262 3808 1263 3812
rect 1267 3808 1268 3812
rect 1262 3807 1268 3808
rect 1382 3812 1388 3813
rect 1382 3808 1383 3812
rect 1387 3808 1388 3812
rect 1382 3807 1388 3808
rect 1502 3812 1508 3813
rect 1502 3808 1503 3812
rect 1507 3808 1508 3812
rect 1502 3807 1508 3808
rect 1630 3812 1636 3813
rect 1630 3808 1631 3812
rect 1635 3808 1636 3812
rect 2008 3810 2010 3837
rect 2046 3833 2047 3837
rect 2051 3833 2052 3837
rect 2262 3836 2263 3840
rect 2267 3836 2268 3840
rect 2262 3835 2268 3836
rect 2374 3840 2380 3841
rect 2374 3836 2375 3840
rect 2379 3836 2380 3840
rect 2374 3835 2380 3836
rect 2494 3840 2500 3841
rect 2494 3836 2495 3840
rect 2499 3836 2500 3840
rect 2494 3835 2500 3836
rect 2630 3840 2636 3841
rect 2630 3836 2631 3840
rect 2635 3836 2636 3840
rect 2630 3835 2636 3836
rect 2774 3840 2780 3841
rect 2774 3836 2775 3840
rect 2779 3836 2780 3840
rect 2774 3835 2780 3836
rect 2918 3840 2924 3841
rect 2918 3836 2919 3840
rect 2923 3836 2924 3840
rect 2918 3835 2924 3836
rect 3062 3840 3068 3841
rect 3062 3836 3063 3840
rect 3067 3836 3068 3840
rect 3062 3835 3068 3836
rect 3206 3840 3212 3841
rect 3206 3836 3207 3840
rect 3211 3836 3212 3840
rect 3206 3835 3212 3836
rect 3342 3840 3348 3841
rect 3342 3836 3343 3840
rect 3347 3836 3348 3840
rect 3342 3835 3348 3836
rect 3470 3840 3476 3841
rect 3470 3836 3471 3840
rect 3475 3836 3476 3840
rect 3470 3835 3476 3836
rect 3598 3840 3604 3841
rect 3598 3836 3599 3840
rect 3603 3836 3604 3840
rect 3598 3835 3604 3836
rect 3726 3840 3732 3841
rect 3726 3836 3727 3840
rect 3731 3836 3732 3840
rect 3726 3835 3732 3836
rect 3838 3840 3844 3841
rect 3838 3836 3839 3840
rect 3843 3836 3844 3840
rect 3944 3838 3946 3865
rect 3838 3835 3844 3836
rect 3942 3837 3948 3838
rect 2046 3832 2052 3833
rect 3942 3833 3943 3837
rect 3947 3833 3948 3837
rect 3942 3832 3948 3833
rect 2262 3821 2268 3822
rect 2046 3820 2052 3821
rect 2046 3816 2047 3820
rect 2051 3816 2052 3820
rect 2262 3817 2263 3821
rect 2267 3817 2268 3821
rect 2262 3816 2268 3817
rect 2374 3821 2380 3822
rect 2374 3817 2375 3821
rect 2379 3817 2380 3821
rect 2374 3816 2380 3817
rect 2494 3821 2500 3822
rect 2494 3817 2495 3821
rect 2499 3817 2500 3821
rect 2494 3816 2500 3817
rect 2630 3821 2636 3822
rect 2630 3817 2631 3821
rect 2635 3817 2636 3821
rect 2630 3816 2636 3817
rect 2774 3821 2780 3822
rect 2774 3817 2775 3821
rect 2779 3817 2780 3821
rect 2774 3816 2780 3817
rect 2918 3821 2924 3822
rect 2918 3817 2919 3821
rect 2923 3817 2924 3821
rect 2918 3816 2924 3817
rect 3062 3821 3068 3822
rect 3062 3817 3063 3821
rect 3067 3817 3068 3821
rect 3062 3816 3068 3817
rect 3206 3821 3212 3822
rect 3206 3817 3207 3821
rect 3211 3817 3212 3821
rect 3206 3816 3212 3817
rect 3342 3821 3348 3822
rect 3342 3817 3343 3821
rect 3347 3817 3348 3821
rect 3342 3816 3348 3817
rect 3470 3821 3476 3822
rect 3470 3817 3471 3821
rect 3475 3817 3476 3821
rect 3470 3816 3476 3817
rect 3598 3821 3604 3822
rect 3598 3817 3599 3821
rect 3603 3817 3604 3821
rect 3598 3816 3604 3817
rect 3726 3821 3732 3822
rect 3726 3817 3727 3821
rect 3731 3817 3732 3821
rect 3726 3816 3732 3817
rect 3838 3821 3844 3822
rect 3838 3817 3839 3821
rect 3843 3817 3844 3821
rect 3838 3816 3844 3817
rect 3942 3820 3948 3821
rect 3942 3816 3943 3820
rect 3947 3816 3948 3820
rect 2046 3815 2052 3816
rect 1630 3807 1636 3808
rect 2006 3809 2012 3810
rect 110 3804 116 3805
rect 2006 3805 2007 3809
rect 2011 3805 2012 3809
rect 2006 3804 2012 3805
rect 230 3793 236 3794
rect 110 3792 116 3793
rect 110 3788 111 3792
rect 115 3788 116 3792
rect 230 3789 231 3793
rect 235 3789 236 3793
rect 230 3788 236 3789
rect 334 3793 340 3794
rect 334 3789 335 3793
rect 339 3789 340 3793
rect 334 3788 340 3789
rect 438 3793 444 3794
rect 438 3789 439 3793
rect 443 3789 444 3793
rect 438 3788 444 3789
rect 534 3793 540 3794
rect 534 3789 535 3793
rect 539 3789 540 3793
rect 534 3788 540 3789
rect 630 3793 636 3794
rect 630 3789 631 3793
rect 635 3789 636 3793
rect 630 3788 636 3789
rect 726 3793 732 3794
rect 726 3789 727 3793
rect 731 3789 732 3793
rect 726 3788 732 3789
rect 830 3793 836 3794
rect 830 3789 831 3793
rect 835 3789 836 3793
rect 830 3788 836 3789
rect 934 3793 940 3794
rect 934 3789 935 3793
rect 939 3789 940 3793
rect 934 3788 940 3789
rect 1038 3793 1044 3794
rect 1038 3789 1039 3793
rect 1043 3789 1044 3793
rect 1038 3788 1044 3789
rect 1150 3793 1156 3794
rect 1150 3789 1151 3793
rect 1155 3789 1156 3793
rect 1150 3788 1156 3789
rect 1262 3793 1268 3794
rect 1262 3789 1263 3793
rect 1267 3789 1268 3793
rect 1262 3788 1268 3789
rect 1382 3793 1388 3794
rect 1382 3789 1383 3793
rect 1387 3789 1388 3793
rect 1382 3788 1388 3789
rect 1502 3793 1508 3794
rect 1502 3789 1503 3793
rect 1507 3789 1508 3793
rect 1502 3788 1508 3789
rect 1630 3793 1636 3794
rect 1630 3789 1631 3793
rect 1635 3789 1636 3793
rect 1630 3788 1636 3789
rect 2006 3792 2012 3793
rect 2006 3788 2007 3792
rect 2011 3788 2012 3792
rect 110 3787 116 3788
rect 112 3767 114 3787
rect 232 3767 234 3788
rect 336 3767 338 3788
rect 440 3767 442 3788
rect 536 3767 538 3788
rect 632 3767 634 3788
rect 728 3767 730 3788
rect 832 3767 834 3788
rect 936 3767 938 3788
rect 1040 3767 1042 3788
rect 1152 3767 1154 3788
rect 1264 3767 1266 3788
rect 1384 3767 1386 3788
rect 1504 3767 1506 3788
rect 1632 3767 1634 3788
rect 2006 3787 2012 3788
rect 2008 3767 2010 3787
rect 2048 3779 2050 3815
rect 2264 3779 2266 3816
rect 2376 3779 2378 3816
rect 2496 3779 2498 3816
rect 2632 3779 2634 3816
rect 2776 3779 2778 3816
rect 2920 3779 2922 3816
rect 3064 3779 3066 3816
rect 3208 3779 3210 3816
rect 3344 3779 3346 3816
rect 3472 3779 3474 3816
rect 3600 3779 3602 3816
rect 3728 3779 3730 3816
rect 3840 3779 3842 3816
rect 3942 3815 3948 3816
rect 3944 3779 3946 3815
rect 2047 3778 2051 3779
rect 2047 3773 2051 3774
rect 2071 3778 2075 3779
rect 2071 3773 2075 3774
rect 2183 3778 2187 3779
rect 2183 3773 2187 3774
rect 2263 3778 2267 3779
rect 2263 3773 2267 3774
rect 2327 3778 2331 3779
rect 2327 3773 2331 3774
rect 2375 3778 2379 3779
rect 2375 3773 2379 3774
rect 2479 3778 2483 3779
rect 2479 3773 2483 3774
rect 2495 3778 2499 3779
rect 2495 3773 2499 3774
rect 2631 3778 2635 3779
rect 2631 3773 2635 3774
rect 2639 3778 2643 3779
rect 2639 3773 2643 3774
rect 2775 3778 2779 3779
rect 2775 3773 2779 3774
rect 2807 3778 2811 3779
rect 2807 3773 2811 3774
rect 2919 3778 2923 3779
rect 2919 3773 2923 3774
rect 2983 3778 2987 3779
rect 2983 3773 2987 3774
rect 3063 3778 3067 3779
rect 3063 3773 3067 3774
rect 3159 3778 3163 3779
rect 3159 3773 3163 3774
rect 3207 3778 3211 3779
rect 3207 3773 3211 3774
rect 3335 3778 3339 3779
rect 3335 3773 3339 3774
rect 3343 3778 3347 3779
rect 3343 3773 3347 3774
rect 3471 3778 3475 3779
rect 3471 3773 3475 3774
rect 3511 3778 3515 3779
rect 3511 3773 3515 3774
rect 3599 3778 3603 3779
rect 3599 3773 3603 3774
rect 3687 3778 3691 3779
rect 3687 3773 3691 3774
rect 3727 3778 3731 3779
rect 3727 3773 3731 3774
rect 3839 3778 3843 3779
rect 3839 3773 3843 3774
rect 3943 3778 3947 3779
rect 3943 3773 3947 3774
rect 111 3766 115 3767
rect 111 3761 115 3762
rect 159 3766 163 3767
rect 159 3761 163 3762
rect 231 3766 235 3767
rect 231 3761 235 3762
rect 335 3766 339 3767
rect 335 3761 339 3762
rect 351 3766 355 3767
rect 351 3761 355 3762
rect 439 3766 443 3767
rect 439 3761 443 3762
rect 535 3766 539 3767
rect 535 3761 539 3762
rect 551 3766 555 3767
rect 551 3761 555 3762
rect 631 3766 635 3767
rect 631 3761 635 3762
rect 727 3766 731 3767
rect 727 3761 731 3762
rect 751 3766 755 3767
rect 751 3761 755 3762
rect 831 3766 835 3767
rect 831 3761 835 3762
rect 935 3766 939 3767
rect 935 3761 939 3762
rect 959 3766 963 3767
rect 959 3761 963 3762
rect 1039 3766 1043 3767
rect 1039 3761 1043 3762
rect 1151 3766 1155 3767
rect 1151 3761 1155 3762
rect 1167 3766 1171 3767
rect 1167 3761 1171 3762
rect 1263 3766 1267 3767
rect 1263 3761 1267 3762
rect 1383 3766 1387 3767
rect 1383 3761 1387 3762
rect 1503 3766 1507 3767
rect 1503 3761 1507 3762
rect 1607 3766 1611 3767
rect 1607 3761 1611 3762
rect 1631 3766 1635 3767
rect 1631 3761 1635 3762
rect 2007 3766 2011 3767
rect 2007 3761 2011 3762
rect 112 3741 114 3761
rect 110 3740 116 3741
rect 160 3740 162 3761
rect 352 3740 354 3761
rect 552 3740 554 3761
rect 752 3740 754 3761
rect 960 3740 962 3761
rect 1168 3740 1170 3761
rect 1384 3740 1386 3761
rect 1608 3740 1610 3761
rect 2008 3741 2010 3761
rect 2048 3753 2050 3773
rect 2046 3752 2052 3753
rect 2072 3752 2074 3773
rect 2184 3752 2186 3773
rect 2328 3752 2330 3773
rect 2480 3752 2482 3773
rect 2640 3752 2642 3773
rect 2808 3752 2810 3773
rect 2984 3752 2986 3773
rect 3160 3752 3162 3773
rect 3336 3752 3338 3773
rect 3512 3752 3514 3773
rect 3688 3752 3690 3773
rect 3840 3752 3842 3773
rect 3944 3753 3946 3773
rect 3942 3752 3948 3753
rect 2046 3748 2047 3752
rect 2051 3748 2052 3752
rect 2046 3747 2052 3748
rect 2070 3751 2076 3752
rect 2070 3747 2071 3751
rect 2075 3747 2076 3751
rect 2070 3746 2076 3747
rect 2182 3751 2188 3752
rect 2182 3747 2183 3751
rect 2187 3747 2188 3751
rect 2182 3746 2188 3747
rect 2326 3751 2332 3752
rect 2326 3747 2327 3751
rect 2331 3747 2332 3751
rect 2326 3746 2332 3747
rect 2478 3751 2484 3752
rect 2478 3747 2479 3751
rect 2483 3747 2484 3751
rect 2478 3746 2484 3747
rect 2638 3751 2644 3752
rect 2638 3747 2639 3751
rect 2643 3747 2644 3751
rect 2638 3746 2644 3747
rect 2806 3751 2812 3752
rect 2806 3747 2807 3751
rect 2811 3747 2812 3751
rect 2806 3746 2812 3747
rect 2982 3751 2988 3752
rect 2982 3747 2983 3751
rect 2987 3747 2988 3751
rect 2982 3746 2988 3747
rect 3158 3751 3164 3752
rect 3158 3747 3159 3751
rect 3163 3747 3164 3751
rect 3158 3746 3164 3747
rect 3334 3751 3340 3752
rect 3334 3747 3335 3751
rect 3339 3747 3340 3751
rect 3334 3746 3340 3747
rect 3510 3751 3516 3752
rect 3510 3747 3511 3751
rect 3515 3747 3516 3751
rect 3510 3746 3516 3747
rect 3686 3751 3692 3752
rect 3686 3747 3687 3751
rect 3691 3747 3692 3751
rect 3686 3746 3692 3747
rect 3838 3751 3844 3752
rect 3838 3747 3839 3751
rect 3843 3747 3844 3751
rect 3942 3748 3943 3752
rect 3947 3748 3948 3752
rect 3942 3747 3948 3748
rect 3838 3746 3844 3747
rect 2006 3740 2012 3741
rect 110 3736 111 3740
rect 115 3736 116 3740
rect 110 3735 116 3736
rect 158 3739 164 3740
rect 158 3735 159 3739
rect 163 3735 164 3739
rect 158 3734 164 3735
rect 350 3739 356 3740
rect 350 3735 351 3739
rect 355 3735 356 3739
rect 350 3734 356 3735
rect 550 3739 556 3740
rect 550 3735 551 3739
rect 555 3735 556 3739
rect 550 3734 556 3735
rect 750 3739 756 3740
rect 750 3735 751 3739
rect 755 3735 756 3739
rect 750 3734 756 3735
rect 958 3739 964 3740
rect 958 3735 959 3739
rect 963 3735 964 3739
rect 958 3734 964 3735
rect 1166 3739 1172 3740
rect 1166 3735 1167 3739
rect 1171 3735 1172 3739
rect 1166 3734 1172 3735
rect 1382 3739 1388 3740
rect 1382 3735 1383 3739
rect 1387 3735 1388 3739
rect 1382 3734 1388 3735
rect 1606 3739 1612 3740
rect 1606 3735 1607 3739
rect 1611 3735 1612 3739
rect 2006 3736 2007 3740
rect 2011 3736 2012 3740
rect 2006 3735 2012 3736
rect 2046 3735 2052 3736
rect 1606 3734 1612 3735
rect 2046 3731 2047 3735
rect 2051 3731 2052 3735
rect 3942 3735 3948 3736
rect 2046 3730 2052 3731
rect 2070 3732 2076 3733
rect 110 3723 116 3724
rect 110 3719 111 3723
rect 115 3719 116 3723
rect 2006 3723 2012 3724
rect 110 3718 116 3719
rect 158 3720 164 3721
rect 112 3683 114 3718
rect 158 3716 159 3720
rect 163 3716 164 3720
rect 158 3715 164 3716
rect 350 3720 356 3721
rect 350 3716 351 3720
rect 355 3716 356 3720
rect 350 3715 356 3716
rect 550 3720 556 3721
rect 550 3716 551 3720
rect 555 3716 556 3720
rect 550 3715 556 3716
rect 750 3720 756 3721
rect 750 3716 751 3720
rect 755 3716 756 3720
rect 750 3715 756 3716
rect 958 3720 964 3721
rect 958 3716 959 3720
rect 963 3716 964 3720
rect 958 3715 964 3716
rect 1166 3720 1172 3721
rect 1166 3716 1167 3720
rect 1171 3716 1172 3720
rect 1166 3715 1172 3716
rect 1382 3720 1388 3721
rect 1382 3716 1383 3720
rect 1387 3716 1388 3720
rect 1382 3715 1388 3716
rect 1606 3720 1612 3721
rect 1606 3716 1607 3720
rect 1611 3716 1612 3720
rect 2006 3719 2007 3723
rect 2011 3719 2012 3723
rect 2006 3718 2012 3719
rect 1606 3715 1612 3716
rect 160 3683 162 3715
rect 352 3683 354 3715
rect 552 3683 554 3715
rect 752 3683 754 3715
rect 960 3683 962 3715
rect 1168 3683 1170 3715
rect 1384 3683 1386 3715
rect 1608 3683 1610 3715
rect 2008 3683 2010 3718
rect 2048 3691 2050 3730
rect 2070 3728 2071 3732
rect 2075 3728 2076 3732
rect 2070 3727 2076 3728
rect 2182 3732 2188 3733
rect 2182 3728 2183 3732
rect 2187 3728 2188 3732
rect 2182 3727 2188 3728
rect 2326 3732 2332 3733
rect 2326 3728 2327 3732
rect 2331 3728 2332 3732
rect 2326 3727 2332 3728
rect 2478 3732 2484 3733
rect 2478 3728 2479 3732
rect 2483 3728 2484 3732
rect 2478 3727 2484 3728
rect 2638 3732 2644 3733
rect 2638 3728 2639 3732
rect 2643 3728 2644 3732
rect 2638 3727 2644 3728
rect 2806 3732 2812 3733
rect 2806 3728 2807 3732
rect 2811 3728 2812 3732
rect 2806 3727 2812 3728
rect 2982 3732 2988 3733
rect 2982 3728 2983 3732
rect 2987 3728 2988 3732
rect 2982 3727 2988 3728
rect 3158 3732 3164 3733
rect 3158 3728 3159 3732
rect 3163 3728 3164 3732
rect 3158 3727 3164 3728
rect 3334 3732 3340 3733
rect 3334 3728 3335 3732
rect 3339 3728 3340 3732
rect 3334 3727 3340 3728
rect 3510 3732 3516 3733
rect 3510 3728 3511 3732
rect 3515 3728 3516 3732
rect 3510 3727 3516 3728
rect 3686 3732 3692 3733
rect 3686 3728 3687 3732
rect 3691 3728 3692 3732
rect 3686 3727 3692 3728
rect 3838 3732 3844 3733
rect 3838 3728 3839 3732
rect 3843 3728 3844 3732
rect 3942 3731 3943 3735
rect 3947 3731 3948 3735
rect 3942 3730 3948 3731
rect 3838 3727 3844 3728
rect 2072 3691 2074 3727
rect 2184 3691 2186 3727
rect 2328 3691 2330 3727
rect 2480 3691 2482 3727
rect 2640 3691 2642 3727
rect 2808 3691 2810 3727
rect 2984 3691 2986 3727
rect 3160 3691 3162 3727
rect 3336 3691 3338 3727
rect 3512 3691 3514 3727
rect 3688 3691 3690 3727
rect 3840 3691 3842 3727
rect 3944 3691 3946 3730
rect 2047 3690 2051 3691
rect 2047 3685 2051 3686
rect 2071 3690 2075 3691
rect 2071 3685 2075 3686
rect 2183 3690 2187 3691
rect 2183 3685 2187 3686
rect 2199 3690 2203 3691
rect 2199 3685 2203 3686
rect 2327 3690 2331 3691
rect 2327 3685 2331 3686
rect 2367 3690 2371 3691
rect 2367 3685 2371 3686
rect 2479 3690 2483 3691
rect 2479 3685 2483 3686
rect 2551 3690 2555 3691
rect 2551 3685 2555 3686
rect 2639 3690 2643 3691
rect 2639 3685 2643 3686
rect 2735 3690 2739 3691
rect 2735 3685 2739 3686
rect 2807 3690 2811 3691
rect 2807 3685 2811 3686
rect 2927 3690 2931 3691
rect 2927 3685 2931 3686
rect 2983 3690 2987 3691
rect 2983 3685 2987 3686
rect 3111 3690 3115 3691
rect 3111 3685 3115 3686
rect 3159 3690 3163 3691
rect 3159 3685 3163 3686
rect 3295 3690 3299 3691
rect 3295 3685 3299 3686
rect 3335 3690 3339 3691
rect 3335 3685 3339 3686
rect 3479 3690 3483 3691
rect 3479 3685 3483 3686
rect 3511 3690 3515 3691
rect 3511 3685 3515 3686
rect 3671 3690 3675 3691
rect 3671 3685 3675 3686
rect 3687 3690 3691 3691
rect 3687 3685 3691 3686
rect 3839 3690 3843 3691
rect 3839 3685 3843 3686
rect 3943 3690 3947 3691
rect 3943 3685 3947 3686
rect 111 3682 115 3683
rect 111 3677 115 3678
rect 151 3682 155 3683
rect 151 3677 155 3678
rect 159 3682 163 3683
rect 159 3677 163 3678
rect 351 3682 355 3683
rect 351 3677 355 3678
rect 383 3682 387 3683
rect 383 3677 387 3678
rect 551 3682 555 3683
rect 551 3677 555 3678
rect 615 3682 619 3683
rect 615 3677 619 3678
rect 751 3682 755 3683
rect 751 3677 755 3678
rect 839 3682 843 3683
rect 839 3677 843 3678
rect 959 3682 963 3683
rect 959 3677 963 3678
rect 1055 3682 1059 3683
rect 1055 3677 1059 3678
rect 1167 3682 1171 3683
rect 1167 3677 1171 3678
rect 1263 3682 1267 3683
rect 1263 3677 1267 3678
rect 1383 3682 1387 3683
rect 1383 3677 1387 3678
rect 1479 3682 1483 3683
rect 1479 3677 1483 3678
rect 1607 3682 1611 3683
rect 1607 3677 1611 3678
rect 1695 3682 1699 3683
rect 1695 3677 1699 3678
rect 2007 3682 2011 3683
rect 2007 3677 2011 3678
rect 112 3650 114 3677
rect 152 3653 154 3677
rect 384 3653 386 3677
rect 616 3653 618 3677
rect 840 3653 842 3677
rect 1056 3653 1058 3677
rect 1264 3653 1266 3677
rect 1480 3653 1482 3677
rect 1696 3653 1698 3677
rect 150 3652 156 3653
rect 110 3649 116 3650
rect 110 3645 111 3649
rect 115 3645 116 3649
rect 150 3648 151 3652
rect 155 3648 156 3652
rect 150 3647 156 3648
rect 382 3652 388 3653
rect 382 3648 383 3652
rect 387 3648 388 3652
rect 382 3647 388 3648
rect 614 3652 620 3653
rect 614 3648 615 3652
rect 619 3648 620 3652
rect 614 3647 620 3648
rect 838 3652 844 3653
rect 838 3648 839 3652
rect 843 3648 844 3652
rect 838 3647 844 3648
rect 1054 3652 1060 3653
rect 1054 3648 1055 3652
rect 1059 3648 1060 3652
rect 1054 3647 1060 3648
rect 1262 3652 1268 3653
rect 1262 3648 1263 3652
rect 1267 3648 1268 3652
rect 1262 3647 1268 3648
rect 1478 3652 1484 3653
rect 1478 3648 1479 3652
rect 1483 3648 1484 3652
rect 1478 3647 1484 3648
rect 1694 3652 1700 3653
rect 1694 3648 1695 3652
rect 1699 3648 1700 3652
rect 2008 3650 2010 3677
rect 2048 3658 2050 3685
rect 2072 3661 2074 3685
rect 2200 3661 2202 3685
rect 2368 3661 2370 3685
rect 2552 3661 2554 3685
rect 2736 3661 2738 3685
rect 2928 3661 2930 3685
rect 3112 3661 3114 3685
rect 3296 3661 3298 3685
rect 3480 3661 3482 3685
rect 3672 3661 3674 3685
rect 3840 3661 3842 3685
rect 2070 3660 2076 3661
rect 2046 3657 2052 3658
rect 2046 3653 2047 3657
rect 2051 3653 2052 3657
rect 2070 3656 2071 3660
rect 2075 3656 2076 3660
rect 2070 3655 2076 3656
rect 2198 3660 2204 3661
rect 2198 3656 2199 3660
rect 2203 3656 2204 3660
rect 2198 3655 2204 3656
rect 2366 3660 2372 3661
rect 2366 3656 2367 3660
rect 2371 3656 2372 3660
rect 2366 3655 2372 3656
rect 2550 3660 2556 3661
rect 2550 3656 2551 3660
rect 2555 3656 2556 3660
rect 2550 3655 2556 3656
rect 2734 3660 2740 3661
rect 2734 3656 2735 3660
rect 2739 3656 2740 3660
rect 2734 3655 2740 3656
rect 2926 3660 2932 3661
rect 2926 3656 2927 3660
rect 2931 3656 2932 3660
rect 2926 3655 2932 3656
rect 3110 3660 3116 3661
rect 3110 3656 3111 3660
rect 3115 3656 3116 3660
rect 3110 3655 3116 3656
rect 3294 3660 3300 3661
rect 3294 3656 3295 3660
rect 3299 3656 3300 3660
rect 3294 3655 3300 3656
rect 3478 3660 3484 3661
rect 3478 3656 3479 3660
rect 3483 3656 3484 3660
rect 3478 3655 3484 3656
rect 3670 3660 3676 3661
rect 3670 3656 3671 3660
rect 3675 3656 3676 3660
rect 3670 3655 3676 3656
rect 3838 3660 3844 3661
rect 3838 3656 3839 3660
rect 3843 3656 3844 3660
rect 3944 3658 3946 3685
rect 3838 3655 3844 3656
rect 3942 3657 3948 3658
rect 2046 3652 2052 3653
rect 3942 3653 3943 3657
rect 3947 3653 3948 3657
rect 3942 3652 3948 3653
rect 1694 3647 1700 3648
rect 2006 3649 2012 3650
rect 110 3644 116 3645
rect 2006 3645 2007 3649
rect 2011 3645 2012 3649
rect 2006 3644 2012 3645
rect 2070 3641 2076 3642
rect 2046 3640 2052 3641
rect 2046 3636 2047 3640
rect 2051 3636 2052 3640
rect 2070 3637 2071 3641
rect 2075 3637 2076 3641
rect 2070 3636 2076 3637
rect 2198 3641 2204 3642
rect 2198 3637 2199 3641
rect 2203 3637 2204 3641
rect 2198 3636 2204 3637
rect 2366 3641 2372 3642
rect 2366 3637 2367 3641
rect 2371 3637 2372 3641
rect 2366 3636 2372 3637
rect 2550 3641 2556 3642
rect 2550 3637 2551 3641
rect 2555 3637 2556 3641
rect 2550 3636 2556 3637
rect 2734 3641 2740 3642
rect 2734 3637 2735 3641
rect 2739 3637 2740 3641
rect 2734 3636 2740 3637
rect 2926 3641 2932 3642
rect 2926 3637 2927 3641
rect 2931 3637 2932 3641
rect 2926 3636 2932 3637
rect 3110 3641 3116 3642
rect 3110 3637 3111 3641
rect 3115 3637 3116 3641
rect 3110 3636 3116 3637
rect 3294 3641 3300 3642
rect 3294 3637 3295 3641
rect 3299 3637 3300 3641
rect 3294 3636 3300 3637
rect 3478 3641 3484 3642
rect 3478 3637 3479 3641
rect 3483 3637 3484 3641
rect 3478 3636 3484 3637
rect 3670 3641 3676 3642
rect 3670 3637 3671 3641
rect 3675 3637 3676 3641
rect 3670 3636 3676 3637
rect 3838 3641 3844 3642
rect 3838 3637 3839 3641
rect 3843 3637 3844 3641
rect 3838 3636 3844 3637
rect 3942 3640 3948 3641
rect 3942 3636 3943 3640
rect 3947 3636 3948 3640
rect 2046 3635 2052 3636
rect 150 3633 156 3634
rect 110 3632 116 3633
rect 110 3628 111 3632
rect 115 3628 116 3632
rect 150 3629 151 3633
rect 155 3629 156 3633
rect 150 3628 156 3629
rect 382 3633 388 3634
rect 382 3629 383 3633
rect 387 3629 388 3633
rect 382 3628 388 3629
rect 614 3633 620 3634
rect 614 3629 615 3633
rect 619 3629 620 3633
rect 614 3628 620 3629
rect 838 3633 844 3634
rect 838 3629 839 3633
rect 843 3629 844 3633
rect 838 3628 844 3629
rect 1054 3633 1060 3634
rect 1054 3629 1055 3633
rect 1059 3629 1060 3633
rect 1054 3628 1060 3629
rect 1262 3633 1268 3634
rect 1262 3629 1263 3633
rect 1267 3629 1268 3633
rect 1262 3628 1268 3629
rect 1478 3633 1484 3634
rect 1478 3629 1479 3633
rect 1483 3629 1484 3633
rect 1478 3628 1484 3629
rect 1694 3633 1700 3634
rect 1694 3629 1695 3633
rect 1699 3629 1700 3633
rect 1694 3628 1700 3629
rect 2006 3632 2012 3633
rect 2006 3628 2007 3632
rect 2011 3628 2012 3632
rect 110 3627 116 3628
rect 112 3603 114 3627
rect 152 3603 154 3628
rect 384 3603 386 3628
rect 616 3603 618 3628
rect 840 3603 842 3628
rect 1056 3603 1058 3628
rect 1264 3603 1266 3628
rect 1480 3603 1482 3628
rect 1696 3603 1698 3628
rect 2006 3627 2012 3628
rect 2008 3603 2010 3627
rect 2048 3611 2050 3635
rect 2072 3611 2074 3636
rect 2200 3611 2202 3636
rect 2368 3611 2370 3636
rect 2552 3611 2554 3636
rect 2736 3611 2738 3636
rect 2928 3611 2930 3636
rect 3112 3611 3114 3636
rect 3296 3611 3298 3636
rect 3480 3611 3482 3636
rect 3672 3611 3674 3636
rect 3840 3611 3842 3636
rect 3942 3635 3948 3636
rect 3944 3611 3946 3635
rect 2047 3610 2051 3611
rect 2047 3605 2051 3606
rect 2071 3610 2075 3611
rect 2071 3605 2075 3606
rect 2103 3610 2107 3611
rect 2103 3605 2107 3606
rect 2199 3610 2203 3611
rect 2199 3605 2203 3606
rect 2279 3610 2283 3611
rect 2279 3605 2283 3606
rect 2367 3610 2371 3611
rect 2367 3605 2371 3606
rect 2471 3610 2475 3611
rect 2471 3605 2475 3606
rect 2551 3610 2555 3611
rect 2551 3605 2555 3606
rect 2671 3610 2675 3611
rect 2671 3605 2675 3606
rect 2735 3610 2739 3611
rect 2735 3605 2739 3606
rect 2871 3610 2875 3611
rect 2871 3605 2875 3606
rect 2927 3610 2931 3611
rect 2927 3605 2931 3606
rect 3063 3610 3067 3611
rect 3063 3605 3067 3606
rect 3111 3610 3115 3611
rect 3111 3605 3115 3606
rect 3255 3610 3259 3611
rect 3255 3605 3259 3606
rect 3295 3610 3299 3611
rect 3295 3605 3299 3606
rect 3447 3610 3451 3611
rect 3447 3605 3451 3606
rect 3479 3610 3483 3611
rect 3479 3605 3483 3606
rect 3639 3610 3643 3611
rect 3639 3605 3643 3606
rect 3671 3610 3675 3611
rect 3671 3605 3675 3606
rect 3839 3610 3843 3611
rect 3839 3605 3843 3606
rect 3943 3610 3947 3611
rect 3943 3605 3947 3606
rect 111 3602 115 3603
rect 111 3597 115 3598
rect 151 3602 155 3603
rect 151 3597 155 3598
rect 167 3602 171 3603
rect 167 3597 171 3598
rect 359 3602 363 3603
rect 359 3597 363 3598
rect 383 3602 387 3603
rect 383 3597 387 3598
rect 559 3602 563 3603
rect 559 3597 563 3598
rect 615 3602 619 3603
rect 615 3597 619 3598
rect 775 3602 779 3603
rect 775 3597 779 3598
rect 839 3602 843 3603
rect 839 3597 843 3598
rect 991 3602 995 3603
rect 991 3597 995 3598
rect 1055 3602 1059 3603
rect 1055 3597 1059 3598
rect 1215 3602 1219 3603
rect 1215 3597 1219 3598
rect 1263 3602 1267 3603
rect 1263 3597 1267 3598
rect 1447 3602 1451 3603
rect 1447 3597 1451 3598
rect 1479 3602 1483 3603
rect 1479 3597 1483 3598
rect 1687 3602 1691 3603
rect 1687 3597 1691 3598
rect 1695 3602 1699 3603
rect 1695 3597 1699 3598
rect 2007 3602 2011 3603
rect 2007 3597 2011 3598
rect 112 3577 114 3597
rect 110 3576 116 3577
rect 168 3576 170 3597
rect 360 3576 362 3597
rect 560 3576 562 3597
rect 776 3576 778 3597
rect 992 3576 994 3597
rect 1216 3576 1218 3597
rect 1448 3576 1450 3597
rect 1688 3576 1690 3597
rect 2008 3577 2010 3597
rect 2048 3585 2050 3605
rect 2046 3584 2052 3585
rect 2104 3584 2106 3605
rect 2280 3584 2282 3605
rect 2472 3584 2474 3605
rect 2672 3584 2674 3605
rect 2872 3584 2874 3605
rect 3064 3584 3066 3605
rect 3256 3584 3258 3605
rect 3448 3584 3450 3605
rect 3640 3584 3642 3605
rect 3840 3584 3842 3605
rect 3944 3585 3946 3605
rect 3942 3584 3948 3585
rect 2046 3580 2047 3584
rect 2051 3580 2052 3584
rect 2046 3579 2052 3580
rect 2102 3583 2108 3584
rect 2102 3579 2103 3583
rect 2107 3579 2108 3583
rect 2102 3578 2108 3579
rect 2278 3583 2284 3584
rect 2278 3579 2279 3583
rect 2283 3579 2284 3583
rect 2278 3578 2284 3579
rect 2470 3583 2476 3584
rect 2470 3579 2471 3583
rect 2475 3579 2476 3583
rect 2470 3578 2476 3579
rect 2670 3583 2676 3584
rect 2670 3579 2671 3583
rect 2675 3579 2676 3583
rect 2670 3578 2676 3579
rect 2870 3583 2876 3584
rect 2870 3579 2871 3583
rect 2875 3579 2876 3583
rect 2870 3578 2876 3579
rect 3062 3583 3068 3584
rect 3062 3579 3063 3583
rect 3067 3579 3068 3583
rect 3062 3578 3068 3579
rect 3254 3583 3260 3584
rect 3254 3579 3255 3583
rect 3259 3579 3260 3583
rect 3254 3578 3260 3579
rect 3446 3583 3452 3584
rect 3446 3579 3447 3583
rect 3451 3579 3452 3583
rect 3446 3578 3452 3579
rect 3638 3583 3644 3584
rect 3638 3579 3639 3583
rect 3643 3579 3644 3583
rect 3638 3578 3644 3579
rect 3838 3583 3844 3584
rect 3838 3579 3839 3583
rect 3843 3579 3844 3583
rect 3942 3580 3943 3584
rect 3947 3580 3948 3584
rect 3942 3579 3948 3580
rect 3838 3578 3844 3579
rect 2006 3576 2012 3577
rect 110 3572 111 3576
rect 115 3572 116 3576
rect 110 3571 116 3572
rect 166 3575 172 3576
rect 166 3571 167 3575
rect 171 3571 172 3575
rect 166 3570 172 3571
rect 358 3575 364 3576
rect 358 3571 359 3575
rect 363 3571 364 3575
rect 358 3570 364 3571
rect 558 3575 564 3576
rect 558 3571 559 3575
rect 563 3571 564 3575
rect 558 3570 564 3571
rect 774 3575 780 3576
rect 774 3571 775 3575
rect 779 3571 780 3575
rect 774 3570 780 3571
rect 990 3575 996 3576
rect 990 3571 991 3575
rect 995 3571 996 3575
rect 990 3570 996 3571
rect 1214 3575 1220 3576
rect 1214 3571 1215 3575
rect 1219 3571 1220 3575
rect 1214 3570 1220 3571
rect 1446 3575 1452 3576
rect 1446 3571 1447 3575
rect 1451 3571 1452 3575
rect 1446 3570 1452 3571
rect 1686 3575 1692 3576
rect 1686 3571 1687 3575
rect 1691 3571 1692 3575
rect 2006 3572 2007 3576
rect 2011 3572 2012 3576
rect 2006 3571 2012 3572
rect 1686 3570 1692 3571
rect 2046 3567 2052 3568
rect 2046 3563 2047 3567
rect 2051 3563 2052 3567
rect 3942 3567 3948 3568
rect 2046 3562 2052 3563
rect 2102 3564 2108 3565
rect 110 3559 116 3560
rect 110 3555 111 3559
rect 115 3555 116 3559
rect 2006 3559 2012 3560
rect 110 3554 116 3555
rect 166 3556 172 3557
rect 112 3519 114 3554
rect 166 3552 167 3556
rect 171 3552 172 3556
rect 166 3551 172 3552
rect 358 3556 364 3557
rect 358 3552 359 3556
rect 363 3552 364 3556
rect 358 3551 364 3552
rect 558 3556 564 3557
rect 558 3552 559 3556
rect 563 3552 564 3556
rect 558 3551 564 3552
rect 774 3556 780 3557
rect 774 3552 775 3556
rect 779 3552 780 3556
rect 774 3551 780 3552
rect 990 3556 996 3557
rect 990 3552 991 3556
rect 995 3552 996 3556
rect 990 3551 996 3552
rect 1214 3556 1220 3557
rect 1214 3552 1215 3556
rect 1219 3552 1220 3556
rect 1214 3551 1220 3552
rect 1446 3556 1452 3557
rect 1446 3552 1447 3556
rect 1451 3552 1452 3556
rect 1446 3551 1452 3552
rect 1686 3556 1692 3557
rect 1686 3552 1687 3556
rect 1691 3552 1692 3556
rect 2006 3555 2007 3559
rect 2011 3555 2012 3559
rect 2006 3554 2012 3555
rect 1686 3551 1692 3552
rect 168 3519 170 3551
rect 360 3519 362 3551
rect 560 3519 562 3551
rect 776 3519 778 3551
rect 992 3519 994 3551
rect 1216 3519 1218 3551
rect 1448 3519 1450 3551
rect 1688 3519 1690 3551
rect 2008 3519 2010 3554
rect 2048 3531 2050 3562
rect 2102 3560 2103 3564
rect 2107 3560 2108 3564
rect 2102 3559 2108 3560
rect 2278 3564 2284 3565
rect 2278 3560 2279 3564
rect 2283 3560 2284 3564
rect 2278 3559 2284 3560
rect 2470 3564 2476 3565
rect 2470 3560 2471 3564
rect 2475 3560 2476 3564
rect 2470 3559 2476 3560
rect 2670 3564 2676 3565
rect 2670 3560 2671 3564
rect 2675 3560 2676 3564
rect 2670 3559 2676 3560
rect 2870 3564 2876 3565
rect 2870 3560 2871 3564
rect 2875 3560 2876 3564
rect 2870 3559 2876 3560
rect 3062 3564 3068 3565
rect 3062 3560 3063 3564
rect 3067 3560 3068 3564
rect 3062 3559 3068 3560
rect 3254 3564 3260 3565
rect 3254 3560 3255 3564
rect 3259 3560 3260 3564
rect 3254 3559 3260 3560
rect 3446 3564 3452 3565
rect 3446 3560 3447 3564
rect 3451 3560 3452 3564
rect 3446 3559 3452 3560
rect 3638 3564 3644 3565
rect 3638 3560 3639 3564
rect 3643 3560 3644 3564
rect 3638 3559 3644 3560
rect 3838 3564 3844 3565
rect 3838 3560 3839 3564
rect 3843 3560 3844 3564
rect 3942 3563 3943 3567
rect 3947 3563 3948 3567
rect 3942 3562 3948 3563
rect 3838 3559 3844 3560
rect 2104 3531 2106 3559
rect 2280 3531 2282 3559
rect 2472 3531 2474 3559
rect 2672 3531 2674 3559
rect 2872 3531 2874 3559
rect 3064 3531 3066 3559
rect 3256 3531 3258 3559
rect 3448 3531 3450 3559
rect 3640 3531 3642 3559
rect 3840 3531 3842 3559
rect 3944 3531 3946 3562
rect 2047 3530 2051 3531
rect 2047 3525 2051 3526
rect 2103 3530 2107 3531
rect 2103 3525 2107 3526
rect 2279 3530 2283 3531
rect 2279 3525 2283 3526
rect 2327 3530 2331 3531
rect 2327 3525 2331 3526
rect 2447 3530 2451 3531
rect 2447 3525 2451 3526
rect 2471 3530 2475 3531
rect 2471 3525 2475 3526
rect 2583 3530 2587 3531
rect 2583 3525 2587 3526
rect 2671 3530 2675 3531
rect 2671 3525 2675 3526
rect 2735 3530 2739 3531
rect 2735 3525 2739 3526
rect 2871 3530 2875 3531
rect 2871 3525 2875 3526
rect 2911 3530 2915 3531
rect 2911 3525 2915 3526
rect 3063 3530 3067 3531
rect 3063 3525 3067 3526
rect 3111 3530 3115 3531
rect 3111 3525 3115 3526
rect 3255 3530 3259 3531
rect 3255 3525 3259 3526
rect 3335 3530 3339 3531
rect 3335 3525 3339 3526
rect 3447 3530 3451 3531
rect 3447 3525 3451 3526
rect 3567 3530 3571 3531
rect 3567 3525 3571 3526
rect 3639 3530 3643 3531
rect 3639 3525 3643 3526
rect 3807 3530 3811 3531
rect 3807 3525 3811 3526
rect 3839 3530 3843 3531
rect 3839 3525 3843 3526
rect 3943 3530 3947 3531
rect 3943 3525 3947 3526
rect 111 3518 115 3519
rect 111 3513 115 3514
rect 167 3518 171 3519
rect 167 3513 171 3514
rect 295 3518 299 3519
rect 295 3513 299 3514
rect 359 3518 363 3519
rect 359 3513 363 3514
rect 431 3518 435 3519
rect 431 3513 435 3514
rect 559 3518 563 3519
rect 559 3513 563 3514
rect 583 3518 587 3519
rect 583 3513 587 3514
rect 743 3518 747 3519
rect 743 3513 747 3514
rect 775 3518 779 3519
rect 775 3513 779 3514
rect 911 3518 915 3519
rect 911 3513 915 3514
rect 991 3518 995 3519
rect 991 3513 995 3514
rect 1079 3518 1083 3519
rect 1079 3513 1083 3514
rect 1215 3518 1219 3519
rect 1215 3513 1219 3514
rect 1247 3518 1251 3519
rect 1247 3513 1251 3514
rect 1423 3518 1427 3519
rect 1423 3513 1427 3514
rect 1447 3518 1451 3519
rect 1447 3513 1451 3514
rect 1599 3518 1603 3519
rect 1599 3513 1603 3514
rect 1687 3518 1691 3519
rect 1687 3513 1691 3514
rect 1775 3518 1779 3519
rect 1775 3513 1779 3514
rect 2007 3518 2011 3519
rect 2007 3513 2011 3514
rect 112 3486 114 3513
rect 296 3489 298 3513
rect 432 3489 434 3513
rect 584 3489 586 3513
rect 744 3489 746 3513
rect 912 3489 914 3513
rect 1080 3489 1082 3513
rect 1248 3489 1250 3513
rect 1424 3489 1426 3513
rect 1600 3489 1602 3513
rect 1776 3489 1778 3513
rect 294 3488 300 3489
rect 110 3485 116 3486
rect 110 3481 111 3485
rect 115 3481 116 3485
rect 294 3484 295 3488
rect 299 3484 300 3488
rect 294 3483 300 3484
rect 430 3488 436 3489
rect 430 3484 431 3488
rect 435 3484 436 3488
rect 430 3483 436 3484
rect 582 3488 588 3489
rect 582 3484 583 3488
rect 587 3484 588 3488
rect 582 3483 588 3484
rect 742 3488 748 3489
rect 742 3484 743 3488
rect 747 3484 748 3488
rect 742 3483 748 3484
rect 910 3488 916 3489
rect 910 3484 911 3488
rect 915 3484 916 3488
rect 910 3483 916 3484
rect 1078 3488 1084 3489
rect 1078 3484 1079 3488
rect 1083 3484 1084 3488
rect 1078 3483 1084 3484
rect 1246 3488 1252 3489
rect 1246 3484 1247 3488
rect 1251 3484 1252 3488
rect 1246 3483 1252 3484
rect 1422 3488 1428 3489
rect 1422 3484 1423 3488
rect 1427 3484 1428 3488
rect 1422 3483 1428 3484
rect 1598 3488 1604 3489
rect 1598 3484 1599 3488
rect 1603 3484 1604 3488
rect 1598 3483 1604 3484
rect 1774 3488 1780 3489
rect 1774 3484 1775 3488
rect 1779 3484 1780 3488
rect 2008 3486 2010 3513
rect 2048 3498 2050 3525
rect 2328 3501 2330 3525
rect 2448 3501 2450 3525
rect 2584 3501 2586 3525
rect 2736 3501 2738 3525
rect 2912 3501 2914 3525
rect 3112 3501 3114 3525
rect 3336 3501 3338 3525
rect 3568 3501 3570 3525
rect 3808 3501 3810 3525
rect 2326 3500 2332 3501
rect 2046 3497 2052 3498
rect 2046 3493 2047 3497
rect 2051 3493 2052 3497
rect 2326 3496 2327 3500
rect 2331 3496 2332 3500
rect 2326 3495 2332 3496
rect 2446 3500 2452 3501
rect 2446 3496 2447 3500
rect 2451 3496 2452 3500
rect 2446 3495 2452 3496
rect 2582 3500 2588 3501
rect 2582 3496 2583 3500
rect 2587 3496 2588 3500
rect 2582 3495 2588 3496
rect 2734 3500 2740 3501
rect 2734 3496 2735 3500
rect 2739 3496 2740 3500
rect 2734 3495 2740 3496
rect 2910 3500 2916 3501
rect 2910 3496 2911 3500
rect 2915 3496 2916 3500
rect 2910 3495 2916 3496
rect 3110 3500 3116 3501
rect 3110 3496 3111 3500
rect 3115 3496 3116 3500
rect 3110 3495 3116 3496
rect 3334 3500 3340 3501
rect 3334 3496 3335 3500
rect 3339 3496 3340 3500
rect 3334 3495 3340 3496
rect 3566 3500 3572 3501
rect 3566 3496 3567 3500
rect 3571 3496 3572 3500
rect 3566 3495 3572 3496
rect 3806 3500 3812 3501
rect 3806 3496 3807 3500
rect 3811 3496 3812 3500
rect 3944 3498 3946 3525
rect 3806 3495 3812 3496
rect 3942 3497 3948 3498
rect 2046 3492 2052 3493
rect 3942 3493 3943 3497
rect 3947 3493 3948 3497
rect 3942 3492 3948 3493
rect 1774 3483 1780 3484
rect 2006 3485 2012 3486
rect 110 3480 116 3481
rect 2006 3481 2007 3485
rect 2011 3481 2012 3485
rect 2326 3481 2332 3482
rect 2006 3480 2012 3481
rect 2046 3480 2052 3481
rect 2046 3476 2047 3480
rect 2051 3476 2052 3480
rect 2326 3477 2327 3481
rect 2331 3477 2332 3481
rect 2326 3476 2332 3477
rect 2446 3481 2452 3482
rect 2446 3477 2447 3481
rect 2451 3477 2452 3481
rect 2446 3476 2452 3477
rect 2582 3481 2588 3482
rect 2582 3477 2583 3481
rect 2587 3477 2588 3481
rect 2582 3476 2588 3477
rect 2734 3481 2740 3482
rect 2734 3477 2735 3481
rect 2739 3477 2740 3481
rect 2734 3476 2740 3477
rect 2910 3481 2916 3482
rect 2910 3477 2911 3481
rect 2915 3477 2916 3481
rect 2910 3476 2916 3477
rect 3110 3481 3116 3482
rect 3110 3477 3111 3481
rect 3115 3477 3116 3481
rect 3110 3476 3116 3477
rect 3334 3481 3340 3482
rect 3334 3477 3335 3481
rect 3339 3477 3340 3481
rect 3334 3476 3340 3477
rect 3566 3481 3572 3482
rect 3566 3477 3567 3481
rect 3571 3477 3572 3481
rect 3566 3476 3572 3477
rect 3806 3481 3812 3482
rect 3806 3477 3807 3481
rect 3811 3477 3812 3481
rect 3806 3476 3812 3477
rect 3942 3480 3948 3481
rect 3942 3476 3943 3480
rect 3947 3476 3948 3480
rect 2046 3475 2052 3476
rect 294 3469 300 3470
rect 110 3468 116 3469
rect 110 3464 111 3468
rect 115 3464 116 3468
rect 294 3465 295 3469
rect 299 3465 300 3469
rect 294 3464 300 3465
rect 430 3469 436 3470
rect 430 3465 431 3469
rect 435 3465 436 3469
rect 430 3464 436 3465
rect 582 3469 588 3470
rect 582 3465 583 3469
rect 587 3465 588 3469
rect 582 3464 588 3465
rect 742 3469 748 3470
rect 742 3465 743 3469
rect 747 3465 748 3469
rect 742 3464 748 3465
rect 910 3469 916 3470
rect 910 3465 911 3469
rect 915 3465 916 3469
rect 910 3464 916 3465
rect 1078 3469 1084 3470
rect 1078 3465 1079 3469
rect 1083 3465 1084 3469
rect 1078 3464 1084 3465
rect 1246 3469 1252 3470
rect 1246 3465 1247 3469
rect 1251 3465 1252 3469
rect 1246 3464 1252 3465
rect 1422 3469 1428 3470
rect 1422 3465 1423 3469
rect 1427 3465 1428 3469
rect 1422 3464 1428 3465
rect 1598 3469 1604 3470
rect 1598 3465 1599 3469
rect 1603 3465 1604 3469
rect 1598 3464 1604 3465
rect 1774 3469 1780 3470
rect 1774 3465 1775 3469
rect 1779 3465 1780 3469
rect 1774 3464 1780 3465
rect 2006 3468 2012 3469
rect 2006 3464 2007 3468
rect 2011 3464 2012 3468
rect 110 3463 116 3464
rect 112 3423 114 3463
rect 296 3423 298 3464
rect 432 3423 434 3464
rect 584 3423 586 3464
rect 744 3423 746 3464
rect 912 3423 914 3464
rect 1080 3423 1082 3464
rect 1248 3423 1250 3464
rect 1424 3423 1426 3464
rect 1600 3423 1602 3464
rect 1776 3423 1778 3464
rect 2006 3463 2012 3464
rect 2008 3423 2010 3463
rect 2048 3455 2050 3475
rect 2328 3455 2330 3476
rect 2448 3455 2450 3476
rect 2584 3455 2586 3476
rect 2736 3455 2738 3476
rect 2912 3455 2914 3476
rect 3112 3455 3114 3476
rect 3336 3455 3338 3476
rect 3568 3455 3570 3476
rect 3808 3455 3810 3476
rect 3942 3475 3948 3476
rect 3944 3455 3946 3475
rect 2047 3454 2051 3455
rect 2047 3449 2051 3450
rect 2327 3454 2331 3455
rect 2327 3449 2331 3450
rect 2447 3454 2451 3455
rect 2447 3449 2451 3450
rect 2551 3454 2555 3455
rect 2551 3449 2555 3450
rect 2583 3454 2587 3455
rect 2583 3449 2587 3450
rect 2663 3454 2667 3455
rect 2663 3449 2667 3450
rect 2735 3454 2739 3455
rect 2735 3449 2739 3450
rect 2775 3454 2779 3455
rect 2775 3449 2779 3450
rect 2903 3454 2907 3455
rect 2903 3449 2907 3450
rect 2911 3454 2915 3455
rect 2911 3449 2915 3450
rect 3047 3454 3051 3455
rect 3047 3449 3051 3450
rect 3111 3454 3115 3455
rect 3111 3449 3115 3450
rect 3207 3454 3211 3455
rect 3207 3449 3211 3450
rect 3335 3454 3339 3455
rect 3335 3449 3339 3450
rect 3383 3454 3387 3455
rect 3383 3449 3387 3450
rect 3567 3454 3571 3455
rect 3567 3449 3571 3450
rect 3751 3454 3755 3455
rect 3751 3449 3755 3450
rect 3807 3454 3811 3455
rect 3807 3449 3811 3450
rect 3943 3454 3947 3455
rect 3943 3449 3947 3450
rect 2048 3429 2050 3449
rect 2046 3428 2052 3429
rect 2448 3428 2450 3449
rect 2552 3428 2554 3449
rect 2664 3428 2666 3449
rect 2776 3428 2778 3449
rect 2904 3428 2906 3449
rect 3048 3428 3050 3449
rect 3208 3428 3210 3449
rect 3384 3428 3386 3449
rect 3568 3428 3570 3449
rect 3752 3428 3754 3449
rect 3944 3429 3946 3449
rect 3942 3428 3948 3429
rect 2046 3424 2047 3428
rect 2051 3424 2052 3428
rect 2046 3423 2052 3424
rect 2446 3427 2452 3428
rect 2446 3423 2447 3427
rect 2451 3423 2452 3427
rect 111 3422 115 3423
rect 111 3417 115 3418
rect 295 3422 299 3423
rect 295 3417 299 3418
rect 431 3422 435 3423
rect 431 3417 435 3418
rect 495 3422 499 3423
rect 495 3417 499 3418
rect 583 3422 587 3423
rect 583 3417 587 3418
rect 647 3422 651 3423
rect 647 3417 651 3418
rect 743 3422 747 3423
rect 743 3417 747 3418
rect 799 3422 803 3423
rect 799 3417 803 3418
rect 911 3422 915 3423
rect 911 3417 915 3418
rect 959 3422 963 3423
rect 959 3417 963 3418
rect 1079 3422 1083 3423
rect 1079 3417 1083 3418
rect 1127 3422 1131 3423
rect 1127 3417 1131 3418
rect 1247 3422 1251 3423
rect 1247 3417 1251 3418
rect 1295 3422 1299 3423
rect 1295 3417 1299 3418
rect 1423 3422 1427 3423
rect 1423 3417 1427 3418
rect 1463 3422 1467 3423
rect 1463 3417 1467 3418
rect 1599 3422 1603 3423
rect 1599 3417 1603 3418
rect 1639 3422 1643 3423
rect 1639 3417 1643 3418
rect 1775 3422 1779 3423
rect 1775 3417 1779 3418
rect 1815 3422 1819 3423
rect 1815 3417 1819 3418
rect 2007 3422 2011 3423
rect 2446 3422 2452 3423
rect 2550 3427 2556 3428
rect 2550 3423 2551 3427
rect 2555 3423 2556 3427
rect 2550 3422 2556 3423
rect 2662 3427 2668 3428
rect 2662 3423 2663 3427
rect 2667 3423 2668 3427
rect 2662 3422 2668 3423
rect 2774 3427 2780 3428
rect 2774 3423 2775 3427
rect 2779 3423 2780 3427
rect 2774 3422 2780 3423
rect 2902 3427 2908 3428
rect 2902 3423 2903 3427
rect 2907 3423 2908 3427
rect 2902 3422 2908 3423
rect 3046 3427 3052 3428
rect 3046 3423 3047 3427
rect 3051 3423 3052 3427
rect 3046 3422 3052 3423
rect 3206 3427 3212 3428
rect 3206 3423 3207 3427
rect 3211 3423 3212 3427
rect 3206 3422 3212 3423
rect 3382 3427 3388 3428
rect 3382 3423 3383 3427
rect 3387 3423 3388 3427
rect 3382 3422 3388 3423
rect 3566 3427 3572 3428
rect 3566 3423 3567 3427
rect 3571 3423 3572 3427
rect 3566 3422 3572 3423
rect 3750 3427 3756 3428
rect 3750 3423 3751 3427
rect 3755 3423 3756 3427
rect 3942 3424 3943 3428
rect 3947 3424 3948 3428
rect 3942 3423 3948 3424
rect 3750 3422 3756 3423
rect 2007 3417 2011 3418
rect 112 3397 114 3417
rect 110 3396 116 3397
rect 496 3396 498 3417
rect 648 3396 650 3417
rect 800 3396 802 3417
rect 960 3396 962 3417
rect 1128 3396 1130 3417
rect 1296 3396 1298 3417
rect 1464 3396 1466 3417
rect 1640 3396 1642 3417
rect 1816 3396 1818 3417
rect 2008 3397 2010 3417
rect 2046 3411 2052 3412
rect 2046 3407 2047 3411
rect 2051 3407 2052 3411
rect 3942 3411 3948 3412
rect 2046 3406 2052 3407
rect 2446 3408 2452 3409
rect 2006 3396 2012 3397
rect 110 3392 111 3396
rect 115 3392 116 3396
rect 110 3391 116 3392
rect 494 3395 500 3396
rect 494 3391 495 3395
rect 499 3391 500 3395
rect 494 3390 500 3391
rect 646 3395 652 3396
rect 646 3391 647 3395
rect 651 3391 652 3395
rect 646 3390 652 3391
rect 798 3395 804 3396
rect 798 3391 799 3395
rect 803 3391 804 3395
rect 798 3390 804 3391
rect 958 3395 964 3396
rect 958 3391 959 3395
rect 963 3391 964 3395
rect 958 3390 964 3391
rect 1126 3395 1132 3396
rect 1126 3391 1127 3395
rect 1131 3391 1132 3395
rect 1126 3390 1132 3391
rect 1294 3395 1300 3396
rect 1294 3391 1295 3395
rect 1299 3391 1300 3395
rect 1294 3390 1300 3391
rect 1462 3395 1468 3396
rect 1462 3391 1463 3395
rect 1467 3391 1468 3395
rect 1462 3390 1468 3391
rect 1638 3395 1644 3396
rect 1638 3391 1639 3395
rect 1643 3391 1644 3395
rect 1638 3390 1644 3391
rect 1814 3395 1820 3396
rect 1814 3391 1815 3395
rect 1819 3391 1820 3395
rect 2006 3392 2007 3396
rect 2011 3392 2012 3396
rect 2006 3391 2012 3392
rect 1814 3390 1820 3391
rect 110 3379 116 3380
rect 110 3375 111 3379
rect 115 3375 116 3379
rect 2006 3379 2012 3380
rect 110 3374 116 3375
rect 494 3376 500 3377
rect 112 3335 114 3374
rect 494 3372 495 3376
rect 499 3372 500 3376
rect 494 3371 500 3372
rect 646 3376 652 3377
rect 646 3372 647 3376
rect 651 3372 652 3376
rect 646 3371 652 3372
rect 798 3376 804 3377
rect 798 3372 799 3376
rect 803 3372 804 3376
rect 798 3371 804 3372
rect 958 3376 964 3377
rect 958 3372 959 3376
rect 963 3372 964 3376
rect 958 3371 964 3372
rect 1126 3376 1132 3377
rect 1126 3372 1127 3376
rect 1131 3372 1132 3376
rect 1126 3371 1132 3372
rect 1294 3376 1300 3377
rect 1294 3372 1295 3376
rect 1299 3372 1300 3376
rect 1294 3371 1300 3372
rect 1462 3376 1468 3377
rect 1462 3372 1463 3376
rect 1467 3372 1468 3376
rect 1462 3371 1468 3372
rect 1638 3376 1644 3377
rect 1638 3372 1639 3376
rect 1643 3372 1644 3376
rect 1638 3371 1644 3372
rect 1814 3376 1820 3377
rect 1814 3372 1815 3376
rect 1819 3372 1820 3376
rect 2006 3375 2007 3379
rect 2011 3375 2012 3379
rect 2006 3374 2012 3375
rect 1814 3371 1820 3372
rect 496 3335 498 3371
rect 648 3335 650 3371
rect 800 3335 802 3371
rect 960 3335 962 3371
rect 1128 3335 1130 3371
rect 1296 3335 1298 3371
rect 1464 3335 1466 3371
rect 1640 3335 1642 3371
rect 1816 3335 1818 3371
rect 2008 3335 2010 3374
rect 2048 3367 2050 3406
rect 2446 3404 2447 3408
rect 2451 3404 2452 3408
rect 2446 3403 2452 3404
rect 2550 3408 2556 3409
rect 2550 3404 2551 3408
rect 2555 3404 2556 3408
rect 2550 3403 2556 3404
rect 2662 3408 2668 3409
rect 2662 3404 2663 3408
rect 2667 3404 2668 3408
rect 2662 3403 2668 3404
rect 2774 3408 2780 3409
rect 2774 3404 2775 3408
rect 2779 3404 2780 3408
rect 2774 3403 2780 3404
rect 2902 3408 2908 3409
rect 2902 3404 2903 3408
rect 2907 3404 2908 3408
rect 2902 3403 2908 3404
rect 3046 3408 3052 3409
rect 3046 3404 3047 3408
rect 3051 3404 3052 3408
rect 3046 3403 3052 3404
rect 3206 3408 3212 3409
rect 3206 3404 3207 3408
rect 3211 3404 3212 3408
rect 3206 3403 3212 3404
rect 3382 3408 3388 3409
rect 3382 3404 3383 3408
rect 3387 3404 3388 3408
rect 3382 3403 3388 3404
rect 3566 3408 3572 3409
rect 3566 3404 3567 3408
rect 3571 3404 3572 3408
rect 3566 3403 3572 3404
rect 3750 3408 3756 3409
rect 3750 3404 3751 3408
rect 3755 3404 3756 3408
rect 3942 3407 3943 3411
rect 3947 3407 3948 3411
rect 3942 3406 3948 3407
rect 3750 3403 3756 3404
rect 2448 3367 2450 3403
rect 2552 3367 2554 3403
rect 2664 3367 2666 3403
rect 2776 3367 2778 3403
rect 2904 3367 2906 3403
rect 3048 3367 3050 3403
rect 3208 3367 3210 3403
rect 3384 3367 3386 3403
rect 3568 3367 3570 3403
rect 3752 3367 3754 3403
rect 3944 3367 3946 3406
rect 2047 3366 2051 3367
rect 2047 3361 2051 3362
rect 2447 3366 2451 3367
rect 2447 3361 2451 3362
rect 2551 3366 2555 3367
rect 2551 3361 2555 3362
rect 2567 3366 2571 3367
rect 2567 3361 2571 3362
rect 2663 3366 2667 3367
rect 2663 3361 2667 3362
rect 2719 3366 2723 3367
rect 2719 3361 2723 3362
rect 2775 3366 2779 3367
rect 2775 3361 2779 3362
rect 2871 3366 2875 3367
rect 2871 3361 2875 3362
rect 2903 3366 2907 3367
rect 2903 3361 2907 3362
rect 3023 3366 3027 3367
rect 3023 3361 3027 3362
rect 3047 3366 3051 3367
rect 3047 3361 3051 3362
rect 3175 3366 3179 3367
rect 3175 3361 3179 3362
rect 3207 3366 3211 3367
rect 3207 3361 3211 3362
rect 3327 3366 3331 3367
rect 3327 3361 3331 3362
rect 3383 3366 3387 3367
rect 3383 3361 3387 3362
rect 3479 3366 3483 3367
rect 3479 3361 3483 3362
rect 3567 3366 3571 3367
rect 3567 3361 3571 3362
rect 3631 3366 3635 3367
rect 3631 3361 3635 3362
rect 3751 3366 3755 3367
rect 3751 3361 3755 3362
rect 3783 3366 3787 3367
rect 3783 3361 3787 3362
rect 3943 3366 3947 3367
rect 3943 3361 3947 3362
rect 111 3334 115 3335
rect 111 3329 115 3330
rect 135 3334 139 3335
rect 135 3329 139 3330
rect 295 3334 299 3335
rect 295 3329 299 3330
rect 479 3334 483 3335
rect 479 3329 483 3330
rect 495 3334 499 3335
rect 495 3329 499 3330
rect 647 3334 651 3335
rect 647 3329 651 3330
rect 671 3334 675 3335
rect 671 3329 675 3330
rect 799 3334 803 3335
rect 799 3329 803 3330
rect 863 3334 867 3335
rect 863 3329 867 3330
rect 959 3334 963 3335
rect 959 3329 963 3330
rect 1055 3334 1059 3335
rect 1055 3329 1059 3330
rect 1127 3334 1131 3335
rect 1127 3329 1131 3330
rect 1247 3334 1251 3335
rect 1247 3329 1251 3330
rect 1295 3334 1299 3335
rect 1295 3329 1299 3330
rect 1439 3334 1443 3335
rect 1439 3329 1443 3330
rect 1463 3334 1467 3335
rect 1463 3329 1467 3330
rect 1631 3334 1635 3335
rect 1631 3329 1635 3330
rect 1639 3334 1643 3335
rect 1639 3329 1643 3330
rect 1815 3334 1819 3335
rect 1815 3329 1819 3330
rect 1823 3334 1827 3335
rect 1823 3329 1827 3330
rect 2007 3334 2011 3335
rect 2048 3334 2050 3361
rect 2568 3337 2570 3361
rect 2720 3337 2722 3361
rect 2872 3337 2874 3361
rect 3024 3337 3026 3361
rect 3176 3337 3178 3361
rect 3328 3337 3330 3361
rect 3480 3337 3482 3361
rect 3632 3337 3634 3361
rect 3784 3337 3786 3361
rect 2566 3336 2572 3337
rect 2007 3329 2011 3330
rect 2046 3333 2052 3334
rect 2046 3329 2047 3333
rect 2051 3329 2052 3333
rect 2566 3332 2567 3336
rect 2571 3332 2572 3336
rect 2566 3331 2572 3332
rect 2718 3336 2724 3337
rect 2718 3332 2719 3336
rect 2723 3332 2724 3336
rect 2718 3331 2724 3332
rect 2870 3336 2876 3337
rect 2870 3332 2871 3336
rect 2875 3332 2876 3336
rect 2870 3331 2876 3332
rect 3022 3336 3028 3337
rect 3022 3332 3023 3336
rect 3027 3332 3028 3336
rect 3022 3331 3028 3332
rect 3174 3336 3180 3337
rect 3174 3332 3175 3336
rect 3179 3332 3180 3336
rect 3174 3331 3180 3332
rect 3326 3336 3332 3337
rect 3326 3332 3327 3336
rect 3331 3332 3332 3336
rect 3326 3331 3332 3332
rect 3478 3336 3484 3337
rect 3478 3332 3479 3336
rect 3483 3332 3484 3336
rect 3478 3331 3484 3332
rect 3630 3336 3636 3337
rect 3630 3332 3631 3336
rect 3635 3332 3636 3336
rect 3630 3331 3636 3332
rect 3782 3336 3788 3337
rect 3782 3332 3783 3336
rect 3787 3332 3788 3336
rect 3944 3334 3946 3361
rect 3782 3331 3788 3332
rect 3942 3333 3948 3334
rect 112 3302 114 3329
rect 136 3305 138 3329
rect 296 3305 298 3329
rect 480 3305 482 3329
rect 672 3305 674 3329
rect 864 3305 866 3329
rect 1056 3305 1058 3329
rect 1248 3305 1250 3329
rect 1440 3305 1442 3329
rect 1632 3305 1634 3329
rect 1824 3305 1826 3329
rect 134 3304 140 3305
rect 110 3301 116 3302
rect 110 3297 111 3301
rect 115 3297 116 3301
rect 134 3300 135 3304
rect 139 3300 140 3304
rect 134 3299 140 3300
rect 294 3304 300 3305
rect 294 3300 295 3304
rect 299 3300 300 3304
rect 294 3299 300 3300
rect 478 3304 484 3305
rect 478 3300 479 3304
rect 483 3300 484 3304
rect 478 3299 484 3300
rect 670 3304 676 3305
rect 670 3300 671 3304
rect 675 3300 676 3304
rect 670 3299 676 3300
rect 862 3304 868 3305
rect 862 3300 863 3304
rect 867 3300 868 3304
rect 862 3299 868 3300
rect 1054 3304 1060 3305
rect 1054 3300 1055 3304
rect 1059 3300 1060 3304
rect 1054 3299 1060 3300
rect 1246 3304 1252 3305
rect 1246 3300 1247 3304
rect 1251 3300 1252 3304
rect 1246 3299 1252 3300
rect 1438 3304 1444 3305
rect 1438 3300 1439 3304
rect 1443 3300 1444 3304
rect 1438 3299 1444 3300
rect 1630 3304 1636 3305
rect 1630 3300 1631 3304
rect 1635 3300 1636 3304
rect 1630 3299 1636 3300
rect 1822 3304 1828 3305
rect 1822 3300 1823 3304
rect 1827 3300 1828 3304
rect 2008 3302 2010 3329
rect 2046 3328 2052 3329
rect 3942 3329 3943 3333
rect 3947 3329 3948 3333
rect 3942 3328 3948 3329
rect 2566 3317 2572 3318
rect 2046 3316 2052 3317
rect 2046 3312 2047 3316
rect 2051 3312 2052 3316
rect 2566 3313 2567 3317
rect 2571 3313 2572 3317
rect 2566 3312 2572 3313
rect 2718 3317 2724 3318
rect 2718 3313 2719 3317
rect 2723 3313 2724 3317
rect 2718 3312 2724 3313
rect 2870 3317 2876 3318
rect 2870 3313 2871 3317
rect 2875 3313 2876 3317
rect 2870 3312 2876 3313
rect 3022 3317 3028 3318
rect 3022 3313 3023 3317
rect 3027 3313 3028 3317
rect 3022 3312 3028 3313
rect 3174 3317 3180 3318
rect 3174 3313 3175 3317
rect 3179 3313 3180 3317
rect 3174 3312 3180 3313
rect 3326 3317 3332 3318
rect 3326 3313 3327 3317
rect 3331 3313 3332 3317
rect 3326 3312 3332 3313
rect 3478 3317 3484 3318
rect 3478 3313 3479 3317
rect 3483 3313 3484 3317
rect 3478 3312 3484 3313
rect 3630 3317 3636 3318
rect 3630 3313 3631 3317
rect 3635 3313 3636 3317
rect 3630 3312 3636 3313
rect 3782 3317 3788 3318
rect 3782 3313 3783 3317
rect 3787 3313 3788 3317
rect 3782 3312 3788 3313
rect 3942 3316 3948 3317
rect 3942 3312 3943 3316
rect 3947 3312 3948 3316
rect 2046 3311 2052 3312
rect 1822 3299 1828 3300
rect 2006 3301 2012 3302
rect 110 3296 116 3297
rect 2006 3297 2007 3301
rect 2011 3297 2012 3301
rect 2006 3296 2012 3297
rect 2048 3287 2050 3311
rect 2568 3287 2570 3312
rect 2720 3287 2722 3312
rect 2872 3287 2874 3312
rect 3024 3287 3026 3312
rect 3176 3287 3178 3312
rect 3328 3287 3330 3312
rect 3480 3287 3482 3312
rect 3632 3287 3634 3312
rect 3784 3287 3786 3312
rect 3942 3311 3948 3312
rect 3944 3287 3946 3311
rect 2047 3286 2051 3287
rect 134 3285 140 3286
rect 110 3284 116 3285
rect 110 3280 111 3284
rect 115 3280 116 3284
rect 134 3281 135 3285
rect 139 3281 140 3285
rect 134 3280 140 3281
rect 294 3285 300 3286
rect 294 3281 295 3285
rect 299 3281 300 3285
rect 294 3280 300 3281
rect 478 3285 484 3286
rect 478 3281 479 3285
rect 483 3281 484 3285
rect 478 3280 484 3281
rect 670 3285 676 3286
rect 670 3281 671 3285
rect 675 3281 676 3285
rect 670 3280 676 3281
rect 862 3285 868 3286
rect 862 3281 863 3285
rect 867 3281 868 3285
rect 862 3280 868 3281
rect 1054 3285 1060 3286
rect 1054 3281 1055 3285
rect 1059 3281 1060 3285
rect 1054 3280 1060 3281
rect 1246 3285 1252 3286
rect 1246 3281 1247 3285
rect 1251 3281 1252 3285
rect 1246 3280 1252 3281
rect 1438 3285 1444 3286
rect 1438 3281 1439 3285
rect 1443 3281 1444 3285
rect 1438 3280 1444 3281
rect 1630 3285 1636 3286
rect 1630 3281 1631 3285
rect 1635 3281 1636 3285
rect 1630 3280 1636 3281
rect 1822 3285 1828 3286
rect 1822 3281 1823 3285
rect 1827 3281 1828 3285
rect 1822 3280 1828 3281
rect 2006 3284 2012 3285
rect 2006 3280 2007 3284
rect 2011 3280 2012 3284
rect 2047 3281 2051 3282
rect 2415 3286 2419 3287
rect 2415 3281 2419 3282
rect 2551 3286 2555 3287
rect 2551 3281 2555 3282
rect 2567 3286 2571 3287
rect 2567 3281 2571 3282
rect 2687 3286 2691 3287
rect 2687 3281 2691 3282
rect 2719 3286 2723 3287
rect 2719 3281 2723 3282
rect 2831 3286 2835 3287
rect 2831 3281 2835 3282
rect 2871 3286 2875 3287
rect 2871 3281 2875 3282
rect 2975 3286 2979 3287
rect 2975 3281 2979 3282
rect 3023 3286 3027 3287
rect 3023 3281 3027 3282
rect 3119 3286 3123 3287
rect 3119 3281 3123 3282
rect 3175 3286 3179 3287
rect 3175 3281 3179 3282
rect 3255 3286 3259 3287
rect 3255 3281 3259 3282
rect 3327 3286 3331 3287
rect 3327 3281 3331 3282
rect 3383 3286 3387 3287
rect 3383 3281 3387 3282
rect 3479 3286 3483 3287
rect 3479 3281 3483 3282
rect 3503 3286 3507 3287
rect 3503 3281 3507 3282
rect 3623 3286 3627 3287
rect 3623 3281 3627 3282
rect 3631 3286 3635 3287
rect 3631 3281 3635 3282
rect 3743 3286 3747 3287
rect 3743 3281 3747 3282
rect 3783 3286 3787 3287
rect 3783 3281 3787 3282
rect 3839 3286 3843 3287
rect 3839 3281 3843 3282
rect 3943 3286 3947 3287
rect 3943 3281 3947 3282
rect 110 3279 116 3280
rect 112 3255 114 3279
rect 136 3255 138 3280
rect 296 3255 298 3280
rect 480 3255 482 3280
rect 672 3255 674 3280
rect 864 3255 866 3280
rect 1056 3255 1058 3280
rect 1248 3255 1250 3280
rect 1440 3255 1442 3280
rect 1632 3255 1634 3280
rect 1824 3255 1826 3280
rect 2006 3279 2012 3280
rect 2008 3255 2010 3279
rect 2048 3261 2050 3281
rect 2046 3260 2052 3261
rect 2416 3260 2418 3281
rect 2552 3260 2554 3281
rect 2688 3260 2690 3281
rect 2832 3260 2834 3281
rect 2976 3260 2978 3281
rect 3120 3260 3122 3281
rect 3256 3260 3258 3281
rect 3384 3260 3386 3281
rect 3504 3260 3506 3281
rect 3624 3260 3626 3281
rect 3744 3260 3746 3281
rect 3840 3260 3842 3281
rect 3944 3261 3946 3281
rect 3942 3260 3948 3261
rect 2046 3256 2047 3260
rect 2051 3256 2052 3260
rect 2046 3255 2052 3256
rect 2414 3259 2420 3260
rect 2414 3255 2415 3259
rect 2419 3255 2420 3259
rect 111 3254 115 3255
rect 111 3249 115 3250
rect 135 3254 139 3255
rect 135 3249 139 3250
rect 295 3254 299 3255
rect 295 3249 299 3250
rect 319 3254 323 3255
rect 319 3249 323 3250
rect 479 3254 483 3255
rect 479 3249 483 3250
rect 519 3254 523 3255
rect 519 3249 523 3250
rect 671 3254 675 3255
rect 671 3249 675 3250
rect 719 3254 723 3255
rect 719 3249 723 3250
rect 863 3254 867 3255
rect 863 3249 867 3250
rect 911 3254 915 3255
rect 911 3249 915 3250
rect 1055 3254 1059 3255
rect 1055 3249 1059 3250
rect 1095 3254 1099 3255
rect 1095 3249 1099 3250
rect 1247 3254 1251 3255
rect 1247 3249 1251 3250
rect 1271 3254 1275 3255
rect 1271 3249 1275 3250
rect 1439 3254 1443 3255
rect 1439 3249 1443 3250
rect 1447 3254 1451 3255
rect 1447 3249 1451 3250
rect 1623 3254 1627 3255
rect 1623 3249 1627 3250
rect 1631 3254 1635 3255
rect 1631 3249 1635 3250
rect 1799 3254 1803 3255
rect 1799 3249 1803 3250
rect 1823 3254 1827 3255
rect 1823 3249 1827 3250
rect 2007 3254 2011 3255
rect 2414 3254 2420 3255
rect 2550 3259 2556 3260
rect 2550 3255 2551 3259
rect 2555 3255 2556 3259
rect 2550 3254 2556 3255
rect 2686 3259 2692 3260
rect 2686 3255 2687 3259
rect 2691 3255 2692 3259
rect 2686 3254 2692 3255
rect 2830 3259 2836 3260
rect 2830 3255 2831 3259
rect 2835 3255 2836 3259
rect 2830 3254 2836 3255
rect 2974 3259 2980 3260
rect 2974 3255 2975 3259
rect 2979 3255 2980 3259
rect 2974 3254 2980 3255
rect 3118 3259 3124 3260
rect 3118 3255 3119 3259
rect 3123 3255 3124 3259
rect 3118 3254 3124 3255
rect 3254 3259 3260 3260
rect 3254 3255 3255 3259
rect 3259 3255 3260 3259
rect 3254 3254 3260 3255
rect 3382 3259 3388 3260
rect 3382 3255 3383 3259
rect 3387 3255 3388 3259
rect 3382 3254 3388 3255
rect 3502 3259 3508 3260
rect 3502 3255 3503 3259
rect 3507 3255 3508 3259
rect 3502 3254 3508 3255
rect 3622 3259 3628 3260
rect 3622 3255 3623 3259
rect 3627 3255 3628 3259
rect 3622 3254 3628 3255
rect 3742 3259 3748 3260
rect 3742 3255 3743 3259
rect 3747 3255 3748 3259
rect 3742 3254 3748 3255
rect 3838 3259 3844 3260
rect 3838 3255 3839 3259
rect 3843 3255 3844 3259
rect 3942 3256 3943 3260
rect 3947 3256 3948 3260
rect 3942 3255 3948 3256
rect 3838 3254 3844 3255
rect 2007 3249 2011 3250
rect 112 3229 114 3249
rect 110 3228 116 3229
rect 136 3228 138 3249
rect 320 3228 322 3249
rect 520 3228 522 3249
rect 720 3228 722 3249
rect 912 3228 914 3249
rect 1096 3228 1098 3249
rect 1272 3228 1274 3249
rect 1448 3228 1450 3249
rect 1624 3228 1626 3249
rect 1800 3228 1802 3249
rect 2008 3229 2010 3249
rect 2046 3243 2052 3244
rect 2046 3239 2047 3243
rect 2051 3239 2052 3243
rect 3942 3243 3948 3244
rect 2046 3238 2052 3239
rect 2414 3240 2420 3241
rect 2006 3228 2012 3229
rect 110 3224 111 3228
rect 115 3224 116 3228
rect 110 3223 116 3224
rect 134 3227 140 3228
rect 134 3223 135 3227
rect 139 3223 140 3227
rect 134 3222 140 3223
rect 318 3227 324 3228
rect 318 3223 319 3227
rect 323 3223 324 3227
rect 318 3222 324 3223
rect 518 3227 524 3228
rect 518 3223 519 3227
rect 523 3223 524 3227
rect 518 3222 524 3223
rect 718 3227 724 3228
rect 718 3223 719 3227
rect 723 3223 724 3227
rect 718 3222 724 3223
rect 910 3227 916 3228
rect 910 3223 911 3227
rect 915 3223 916 3227
rect 910 3222 916 3223
rect 1094 3227 1100 3228
rect 1094 3223 1095 3227
rect 1099 3223 1100 3227
rect 1094 3222 1100 3223
rect 1270 3227 1276 3228
rect 1270 3223 1271 3227
rect 1275 3223 1276 3227
rect 1270 3222 1276 3223
rect 1446 3227 1452 3228
rect 1446 3223 1447 3227
rect 1451 3223 1452 3227
rect 1446 3222 1452 3223
rect 1622 3227 1628 3228
rect 1622 3223 1623 3227
rect 1627 3223 1628 3227
rect 1622 3222 1628 3223
rect 1798 3227 1804 3228
rect 1798 3223 1799 3227
rect 1803 3223 1804 3227
rect 2006 3224 2007 3228
rect 2011 3224 2012 3228
rect 2006 3223 2012 3224
rect 1798 3222 1804 3223
rect 110 3211 116 3212
rect 110 3207 111 3211
rect 115 3207 116 3211
rect 2006 3211 2012 3212
rect 110 3206 116 3207
rect 134 3208 140 3209
rect 112 3171 114 3206
rect 134 3204 135 3208
rect 139 3204 140 3208
rect 134 3203 140 3204
rect 318 3208 324 3209
rect 318 3204 319 3208
rect 323 3204 324 3208
rect 318 3203 324 3204
rect 518 3208 524 3209
rect 518 3204 519 3208
rect 523 3204 524 3208
rect 518 3203 524 3204
rect 718 3208 724 3209
rect 718 3204 719 3208
rect 723 3204 724 3208
rect 718 3203 724 3204
rect 910 3208 916 3209
rect 910 3204 911 3208
rect 915 3204 916 3208
rect 910 3203 916 3204
rect 1094 3208 1100 3209
rect 1094 3204 1095 3208
rect 1099 3204 1100 3208
rect 1094 3203 1100 3204
rect 1270 3208 1276 3209
rect 1270 3204 1271 3208
rect 1275 3204 1276 3208
rect 1270 3203 1276 3204
rect 1446 3208 1452 3209
rect 1446 3204 1447 3208
rect 1451 3204 1452 3208
rect 1446 3203 1452 3204
rect 1622 3208 1628 3209
rect 1622 3204 1623 3208
rect 1627 3204 1628 3208
rect 1622 3203 1628 3204
rect 1798 3208 1804 3209
rect 1798 3204 1799 3208
rect 1803 3204 1804 3208
rect 2006 3207 2007 3211
rect 2011 3207 2012 3211
rect 2006 3206 2012 3207
rect 1798 3203 1804 3204
rect 136 3171 138 3203
rect 320 3171 322 3203
rect 520 3171 522 3203
rect 720 3171 722 3203
rect 912 3171 914 3203
rect 1096 3171 1098 3203
rect 1272 3171 1274 3203
rect 1448 3171 1450 3203
rect 1624 3171 1626 3203
rect 1800 3171 1802 3203
rect 2008 3171 2010 3206
rect 2048 3199 2050 3238
rect 2414 3236 2415 3240
rect 2419 3236 2420 3240
rect 2414 3235 2420 3236
rect 2550 3240 2556 3241
rect 2550 3236 2551 3240
rect 2555 3236 2556 3240
rect 2550 3235 2556 3236
rect 2686 3240 2692 3241
rect 2686 3236 2687 3240
rect 2691 3236 2692 3240
rect 2686 3235 2692 3236
rect 2830 3240 2836 3241
rect 2830 3236 2831 3240
rect 2835 3236 2836 3240
rect 2830 3235 2836 3236
rect 2974 3240 2980 3241
rect 2974 3236 2975 3240
rect 2979 3236 2980 3240
rect 2974 3235 2980 3236
rect 3118 3240 3124 3241
rect 3118 3236 3119 3240
rect 3123 3236 3124 3240
rect 3118 3235 3124 3236
rect 3254 3240 3260 3241
rect 3254 3236 3255 3240
rect 3259 3236 3260 3240
rect 3254 3235 3260 3236
rect 3382 3240 3388 3241
rect 3382 3236 3383 3240
rect 3387 3236 3388 3240
rect 3382 3235 3388 3236
rect 3502 3240 3508 3241
rect 3502 3236 3503 3240
rect 3507 3236 3508 3240
rect 3502 3235 3508 3236
rect 3622 3240 3628 3241
rect 3622 3236 3623 3240
rect 3627 3236 3628 3240
rect 3622 3235 3628 3236
rect 3742 3240 3748 3241
rect 3742 3236 3743 3240
rect 3747 3236 3748 3240
rect 3742 3235 3748 3236
rect 3838 3240 3844 3241
rect 3838 3236 3839 3240
rect 3843 3236 3844 3240
rect 3942 3239 3943 3243
rect 3947 3239 3948 3243
rect 3942 3238 3948 3239
rect 3838 3235 3844 3236
rect 2416 3199 2418 3235
rect 2552 3199 2554 3235
rect 2688 3199 2690 3235
rect 2832 3199 2834 3235
rect 2976 3199 2978 3235
rect 3120 3199 3122 3235
rect 3256 3199 3258 3235
rect 3384 3199 3386 3235
rect 3504 3199 3506 3235
rect 3624 3199 3626 3235
rect 3744 3199 3746 3235
rect 3840 3199 3842 3235
rect 3944 3199 3946 3238
rect 2047 3198 2051 3199
rect 2047 3193 2051 3194
rect 2247 3198 2251 3199
rect 2247 3193 2251 3194
rect 2399 3198 2403 3199
rect 2399 3193 2403 3194
rect 2415 3198 2419 3199
rect 2415 3193 2419 3194
rect 2551 3198 2555 3199
rect 2551 3193 2555 3194
rect 2559 3198 2563 3199
rect 2559 3193 2563 3194
rect 2687 3198 2691 3199
rect 2687 3193 2691 3194
rect 2727 3198 2731 3199
rect 2727 3193 2731 3194
rect 2831 3198 2835 3199
rect 2831 3193 2835 3194
rect 2903 3198 2907 3199
rect 2903 3193 2907 3194
rect 2975 3198 2979 3199
rect 2975 3193 2979 3194
rect 3079 3198 3083 3199
rect 3079 3193 3083 3194
rect 3119 3198 3123 3199
rect 3119 3193 3123 3194
rect 3255 3198 3259 3199
rect 3255 3193 3259 3194
rect 3263 3198 3267 3199
rect 3263 3193 3267 3194
rect 3383 3198 3387 3199
rect 3383 3193 3387 3194
rect 3447 3198 3451 3199
rect 3447 3193 3451 3194
rect 3503 3198 3507 3199
rect 3503 3193 3507 3194
rect 3623 3198 3627 3199
rect 3623 3193 3627 3194
rect 3631 3198 3635 3199
rect 3631 3193 3635 3194
rect 3743 3198 3747 3199
rect 3743 3193 3747 3194
rect 3815 3198 3819 3199
rect 3815 3193 3819 3194
rect 3839 3198 3843 3199
rect 3839 3193 3843 3194
rect 3943 3198 3947 3199
rect 3943 3193 3947 3194
rect 111 3170 115 3171
rect 111 3165 115 3166
rect 135 3170 139 3171
rect 135 3165 139 3166
rect 143 3170 147 3171
rect 143 3165 147 3166
rect 319 3170 323 3171
rect 319 3165 323 3166
rect 343 3170 347 3171
rect 343 3165 347 3166
rect 519 3170 523 3171
rect 519 3165 523 3166
rect 543 3170 547 3171
rect 543 3165 547 3166
rect 719 3170 723 3171
rect 719 3165 723 3166
rect 743 3170 747 3171
rect 743 3165 747 3166
rect 911 3170 915 3171
rect 911 3165 915 3166
rect 927 3170 931 3171
rect 927 3165 931 3166
rect 1095 3170 1099 3171
rect 1095 3165 1099 3166
rect 1103 3170 1107 3171
rect 1103 3165 1107 3166
rect 1263 3170 1267 3171
rect 1263 3165 1267 3166
rect 1271 3170 1275 3171
rect 1271 3165 1275 3166
rect 1423 3170 1427 3171
rect 1423 3165 1427 3166
rect 1447 3170 1451 3171
rect 1447 3165 1451 3166
rect 1575 3170 1579 3171
rect 1575 3165 1579 3166
rect 1623 3170 1627 3171
rect 1623 3165 1627 3166
rect 1735 3170 1739 3171
rect 1735 3165 1739 3166
rect 1799 3170 1803 3171
rect 1799 3165 1803 3166
rect 2007 3170 2011 3171
rect 2048 3166 2050 3193
rect 2248 3169 2250 3193
rect 2400 3169 2402 3193
rect 2560 3169 2562 3193
rect 2728 3169 2730 3193
rect 2904 3169 2906 3193
rect 3080 3169 3082 3193
rect 3264 3169 3266 3193
rect 3448 3169 3450 3193
rect 3632 3169 3634 3193
rect 3816 3169 3818 3193
rect 2246 3168 2252 3169
rect 2007 3165 2011 3166
rect 2046 3165 2052 3166
rect 112 3138 114 3165
rect 144 3141 146 3165
rect 344 3141 346 3165
rect 544 3141 546 3165
rect 744 3141 746 3165
rect 928 3141 930 3165
rect 1104 3141 1106 3165
rect 1264 3141 1266 3165
rect 1424 3141 1426 3165
rect 1576 3141 1578 3165
rect 1736 3141 1738 3165
rect 142 3140 148 3141
rect 110 3137 116 3138
rect 110 3133 111 3137
rect 115 3133 116 3137
rect 142 3136 143 3140
rect 147 3136 148 3140
rect 142 3135 148 3136
rect 342 3140 348 3141
rect 342 3136 343 3140
rect 347 3136 348 3140
rect 342 3135 348 3136
rect 542 3140 548 3141
rect 542 3136 543 3140
rect 547 3136 548 3140
rect 542 3135 548 3136
rect 742 3140 748 3141
rect 742 3136 743 3140
rect 747 3136 748 3140
rect 742 3135 748 3136
rect 926 3140 932 3141
rect 926 3136 927 3140
rect 931 3136 932 3140
rect 926 3135 932 3136
rect 1102 3140 1108 3141
rect 1102 3136 1103 3140
rect 1107 3136 1108 3140
rect 1102 3135 1108 3136
rect 1262 3140 1268 3141
rect 1262 3136 1263 3140
rect 1267 3136 1268 3140
rect 1262 3135 1268 3136
rect 1422 3140 1428 3141
rect 1422 3136 1423 3140
rect 1427 3136 1428 3140
rect 1422 3135 1428 3136
rect 1574 3140 1580 3141
rect 1574 3136 1575 3140
rect 1579 3136 1580 3140
rect 1574 3135 1580 3136
rect 1734 3140 1740 3141
rect 1734 3136 1735 3140
rect 1739 3136 1740 3140
rect 2008 3138 2010 3165
rect 2046 3161 2047 3165
rect 2051 3161 2052 3165
rect 2246 3164 2247 3168
rect 2251 3164 2252 3168
rect 2246 3163 2252 3164
rect 2398 3168 2404 3169
rect 2398 3164 2399 3168
rect 2403 3164 2404 3168
rect 2398 3163 2404 3164
rect 2558 3168 2564 3169
rect 2558 3164 2559 3168
rect 2563 3164 2564 3168
rect 2558 3163 2564 3164
rect 2726 3168 2732 3169
rect 2726 3164 2727 3168
rect 2731 3164 2732 3168
rect 2726 3163 2732 3164
rect 2902 3168 2908 3169
rect 2902 3164 2903 3168
rect 2907 3164 2908 3168
rect 2902 3163 2908 3164
rect 3078 3168 3084 3169
rect 3078 3164 3079 3168
rect 3083 3164 3084 3168
rect 3078 3163 3084 3164
rect 3262 3168 3268 3169
rect 3262 3164 3263 3168
rect 3267 3164 3268 3168
rect 3262 3163 3268 3164
rect 3446 3168 3452 3169
rect 3446 3164 3447 3168
rect 3451 3164 3452 3168
rect 3446 3163 3452 3164
rect 3630 3168 3636 3169
rect 3630 3164 3631 3168
rect 3635 3164 3636 3168
rect 3630 3163 3636 3164
rect 3814 3168 3820 3169
rect 3814 3164 3815 3168
rect 3819 3164 3820 3168
rect 3944 3166 3946 3193
rect 3814 3163 3820 3164
rect 3942 3165 3948 3166
rect 2046 3160 2052 3161
rect 3942 3161 3943 3165
rect 3947 3161 3948 3165
rect 3942 3160 3948 3161
rect 2246 3149 2252 3150
rect 2046 3148 2052 3149
rect 2046 3144 2047 3148
rect 2051 3144 2052 3148
rect 2246 3145 2247 3149
rect 2251 3145 2252 3149
rect 2246 3144 2252 3145
rect 2398 3149 2404 3150
rect 2398 3145 2399 3149
rect 2403 3145 2404 3149
rect 2398 3144 2404 3145
rect 2558 3149 2564 3150
rect 2558 3145 2559 3149
rect 2563 3145 2564 3149
rect 2558 3144 2564 3145
rect 2726 3149 2732 3150
rect 2726 3145 2727 3149
rect 2731 3145 2732 3149
rect 2726 3144 2732 3145
rect 2902 3149 2908 3150
rect 2902 3145 2903 3149
rect 2907 3145 2908 3149
rect 2902 3144 2908 3145
rect 3078 3149 3084 3150
rect 3078 3145 3079 3149
rect 3083 3145 3084 3149
rect 3078 3144 3084 3145
rect 3262 3149 3268 3150
rect 3262 3145 3263 3149
rect 3267 3145 3268 3149
rect 3262 3144 3268 3145
rect 3446 3149 3452 3150
rect 3446 3145 3447 3149
rect 3451 3145 3452 3149
rect 3446 3144 3452 3145
rect 3630 3149 3636 3150
rect 3630 3145 3631 3149
rect 3635 3145 3636 3149
rect 3630 3144 3636 3145
rect 3814 3149 3820 3150
rect 3814 3145 3815 3149
rect 3819 3145 3820 3149
rect 3814 3144 3820 3145
rect 3942 3148 3948 3149
rect 3942 3144 3943 3148
rect 3947 3144 3948 3148
rect 2046 3143 2052 3144
rect 1734 3135 1740 3136
rect 2006 3137 2012 3138
rect 110 3132 116 3133
rect 2006 3133 2007 3137
rect 2011 3133 2012 3137
rect 2006 3132 2012 3133
rect 142 3121 148 3122
rect 110 3120 116 3121
rect 110 3116 111 3120
rect 115 3116 116 3120
rect 142 3117 143 3121
rect 147 3117 148 3121
rect 142 3116 148 3117
rect 342 3121 348 3122
rect 342 3117 343 3121
rect 347 3117 348 3121
rect 342 3116 348 3117
rect 542 3121 548 3122
rect 542 3117 543 3121
rect 547 3117 548 3121
rect 542 3116 548 3117
rect 742 3121 748 3122
rect 742 3117 743 3121
rect 747 3117 748 3121
rect 742 3116 748 3117
rect 926 3121 932 3122
rect 926 3117 927 3121
rect 931 3117 932 3121
rect 926 3116 932 3117
rect 1102 3121 1108 3122
rect 1102 3117 1103 3121
rect 1107 3117 1108 3121
rect 1102 3116 1108 3117
rect 1262 3121 1268 3122
rect 1262 3117 1263 3121
rect 1267 3117 1268 3121
rect 1262 3116 1268 3117
rect 1422 3121 1428 3122
rect 1422 3117 1423 3121
rect 1427 3117 1428 3121
rect 1422 3116 1428 3117
rect 1574 3121 1580 3122
rect 1574 3117 1575 3121
rect 1579 3117 1580 3121
rect 1574 3116 1580 3117
rect 1734 3121 1740 3122
rect 1734 3117 1735 3121
rect 1739 3117 1740 3121
rect 1734 3116 1740 3117
rect 2006 3120 2012 3121
rect 2006 3116 2007 3120
rect 2011 3116 2012 3120
rect 2048 3119 2050 3143
rect 2248 3119 2250 3144
rect 2400 3119 2402 3144
rect 2560 3119 2562 3144
rect 2728 3119 2730 3144
rect 2904 3119 2906 3144
rect 3080 3119 3082 3144
rect 3264 3119 3266 3144
rect 3448 3119 3450 3144
rect 3632 3119 3634 3144
rect 3816 3119 3818 3144
rect 3942 3143 3948 3144
rect 3944 3119 3946 3143
rect 110 3115 116 3116
rect 112 3095 114 3115
rect 144 3095 146 3116
rect 344 3095 346 3116
rect 544 3095 546 3116
rect 744 3095 746 3116
rect 928 3095 930 3116
rect 1104 3095 1106 3116
rect 1264 3095 1266 3116
rect 1424 3095 1426 3116
rect 1576 3095 1578 3116
rect 1736 3095 1738 3116
rect 2006 3115 2012 3116
rect 2047 3118 2051 3119
rect 2008 3095 2010 3115
rect 2047 3113 2051 3114
rect 2079 3118 2083 3119
rect 2079 3113 2083 3114
rect 2223 3118 2227 3119
rect 2223 3113 2227 3114
rect 2247 3118 2251 3119
rect 2247 3113 2251 3114
rect 2375 3118 2379 3119
rect 2375 3113 2379 3114
rect 2399 3118 2403 3119
rect 2399 3113 2403 3114
rect 2527 3118 2531 3119
rect 2527 3113 2531 3114
rect 2559 3118 2563 3119
rect 2559 3113 2563 3114
rect 2687 3118 2691 3119
rect 2687 3113 2691 3114
rect 2727 3118 2731 3119
rect 2727 3113 2731 3114
rect 2855 3118 2859 3119
rect 2855 3113 2859 3114
rect 2903 3118 2907 3119
rect 2903 3113 2907 3114
rect 3039 3118 3043 3119
rect 3039 3113 3043 3114
rect 3079 3118 3083 3119
rect 3079 3113 3083 3114
rect 3231 3118 3235 3119
rect 3231 3113 3235 3114
rect 3263 3118 3267 3119
rect 3263 3113 3267 3114
rect 3431 3118 3435 3119
rect 3431 3113 3435 3114
rect 3447 3118 3451 3119
rect 3447 3113 3451 3114
rect 3631 3118 3635 3119
rect 3631 3113 3635 3114
rect 3639 3118 3643 3119
rect 3639 3113 3643 3114
rect 3815 3118 3819 3119
rect 3815 3113 3819 3114
rect 3839 3118 3843 3119
rect 3839 3113 3843 3114
rect 3943 3118 3947 3119
rect 3943 3113 3947 3114
rect 111 3094 115 3095
rect 111 3089 115 3090
rect 143 3094 147 3095
rect 143 3089 147 3090
rect 263 3094 267 3095
rect 263 3089 267 3090
rect 343 3094 347 3095
rect 343 3089 347 3090
rect 439 3094 443 3095
rect 439 3089 443 3090
rect 543 3094 547 3095
rect 543 3089 547 3090
rect 615 3094 619 3095
rect 615 3089 619 3090
rect 743 3094 747 3095
rect 743 3089 747 3090
rect 799 3094 803 3095
rect 799 3089 803 3090
rect 927 3094 931 3095
rect 927 3089 931 3090
rect 975 3094 979 3095
rect 975 3089 979 3090
rect 1103 3094 1107 3095
rect 1103 3089 1107 3090
rect 1143 3094 1147 3095
rect 1143 3089 1147 3090
rect 1263 3094 1267 3095
rect 1263 3089 1267 3090
rect 1303 3094 1307 3095
rect 1303 3089 1307 3090
rect 1423 3094 1427 3095
rect 1423 3089 1427 3090
rect 1455 3094 1459 3095
rect 1455 3089 1459 3090
rect 1575 3094 1579 3095
rect 1575 3089 1579 3090
rect 1607 3094 1611 3095
rect 1607 3089 1611 3090
rect 1735 3094 1739 3095
rect 1735 3089 1739 3090
rect 1767 3094 1771 3095
rect 1767 3089 1771 3090
rect 2007 3094 2011 3095
rect 2048 3093 2050 3113
rect 2007 3089 2011 3090
rect 2046 3092 2052 3093
rect 2080 3092 2082 3113
rect 2224 3092 2226 3113
rect 2376 3092 2378 3113
rect 2528 3092 2530 3113
rect 2688 3092 2690 3113
rect 2856 3092 2858 3113
rect 3040 3092 3042 3113
rect 3232 3092 3234 3113
rect 3432 3092 3434 3113
rect 3640 3092 3642 3113
rect 3840 3092 3842 3113
rect 3944 3093 3946 3113
rect 3942 3092 3948 3093
rect 112 3069 114 3089
rect 110 3068 116 3069
rect 264 3068 266 3089
rect 440 3068 442 3089
rect 616 3068 618 3089
rect 800 3068 802 3089
rect 976 3068 978 3089
rect 1144 3068 1146 3089
rect 1304 3068 1306 3089
rect 1456 3068 1458 3089
rect 1608 3068 1610 3089
rect 1768 3068 1770 3089
rect 2008 3069 2010 3089
rect 2046 3088 2047 3092
rect 2051 3088 2052 3092
rect 2046 3087 2052 3088
rect 2078 3091 2084 3092
rect 2078 3087 2079 3091
rect 2083 3087 2084 3091
rect 2078 3086 2084 3087
rect 2222 3091 2228 3092
rect 2222 3087 2223 3091
rect 2227 3087 2228 3091
rect 2222 3086 2228 3087
rect 2374 3091 2380 3092
rect 2374 3087 2375 3091
rect 2379 3087 2380 3091
rect 2374 3086 2380 3087
rect 2526 3091 2532 3092
rect 2526 3087 2527 3091
rect 2531 3087 2532 3091
rect 2526 3086 2532 3087
rect 2686 3091 2692 3092
rect 2686 3087 2687 3091
rect 2691 3087 2692 3091
rect 2686 3086 2692 3087
rect 2854 3091 2860 3092
rect 2854 3087 2855 3091
rect 2859 3087 2860 3091
rect 2854 3086 2860 3087
rect 3038 3091 3044 3092
rect 3038 3087 3039 3091
rect 3043 3087 3044 3091
rect 3038 3086 3044 3087
rect 3230 3091 3236 3092
rect 3230 3087 3231 3091
rect 3235 3087 3236 3091
rect 3230 3086 3236 3087
rect 3430 3091 3436 3092
rect 3430 3087 3431 3091
rect 3435 3087 3436 3091
rect 3430 3086 3436 3087
rect 3638 3091 3644 3092
rect 3638 3087 3639 3091
rect 3643 3087 3644 3091
rect 3638 3086 3644 3087
rect 3838 3091 3844 3092
rect 3838 3087 3839 3091
rect 3843 3087 3844 3091
rect 3942 3088 3943 3092
rect 3947 3088 3948 3092
rect 3942 3087 3948 3088
rect 3838 3086 3844 3087
rect 2046 3075 2052 3076
rect 2046 3071 2047 3075
rect 2051 3071 2052 3075
rect 3942 3075 3948 3076
rect 2046 3070 2052 3071
rect 2078 3072 2084 3073
rect 2006 3068 2012 3069
rect 110 3064 111 3068
rect 115 3064 116 3068
rect 110 3063 116 3064
rect 262 3067 268 3068
rect 262 3063 263 3067
rect 267 3063 268 3067
rect 262 3062 268 3063
rect 438 3067 444 3068
rect 438 3063 439 3067
rect 443 3063 444 3067
rect 438 3062 444 3063
rect 614 3067 620 3068
rect 614 3063 615 3067
rect 619 3063 620 3067
rect 614 3062 620 3063
rect 798 3067 804 3068
rect 798 3063 799 3067
rect 803 3063 804 3067
rect 798 3062 804 3063
rect 974 3067 980 3068
rect 974 3063 975 3067
rect 979 3063 980 3067
rect 974 3062 980 3063
rect 1142 3067 1148 3068
rect 1142 3063 1143 3067
rect 1147 3063 1148 3067
rect 1142 3062 1148 3063
rect 1302 3067 1308 3068
rect 1302 3063 1303 3067
rect 1307 3063 1308 3067
rect 1302 3062 1308 3063
rect 1454 3067 1460 3068
rect 1454 3063 1455 3067
rect 1459 3063 1460 3067
rect 1454 3062 1460 3063
rect 1606 3067 1612 3068
rect 1606 3063 1607 3067
rect 1611 3063 1612 3067
rect 1606 3062 1612 3063
rect 1766 3067 1772 3068
rect 1766 3063 1767 3067
rect 1771 3063 1772 3067
rect 2006 3064 2007 3068
rect 2011 3064 2012 3068
rect 2006 3063 2012 3064
rect 1766 3062 1772 3063
rect 110 3051 116 3052
rect 110 3047 111 3051
rect 115 3047 116 3051
rect 2006 3051 2012 3052
rect 110 3046 116 3047
rect 262 3048 268 3049
rect 112 2995 114 3046
rect 262 3044 263 3048
rect 267 3044 268 3048
rect 262 3043 268 3044
rect 438 3048 444 3049
rect 438 3044 439 3048
rect 443 3044 444 3048
rect 438 3043 444 3044
rect 614 3048 620 3049
rect 614 3044 615 3048
rect 619 3044 620 3048
rect 614 3043 620 3044
rect 798 3048 804 3049
rect 798 3044 799 3048
rect 803 3044 804 3048
rect 798 3043 804 3044
rect 974 3048 980 3049
rect 974 3044 975 3048
rect 979 3044 980 3048
rect 974 3043 980 3044
rect 1142 3048 1148 3049
rect 1142 3044 1143 3048
rect 1147 3044 1148 3048
rect 1142 3043 1148 3044
rect 1302 3048 1308 3049
rect 1302 3044 1303 3048
rect 1307 3044 1308 3048
rect 1302 3043 1308 3044
rect 1454 3048 1460 3049
rect 1454 3044 1455 3048
rect 1459 3044 1460 3048
rect 1454 3043 1460 3044
rect 1606 3048 1612 3049
rect 1606 3044 1607 3048
rect 1611 3044 1612 3048
rect 1606 3043 1612 3044
rect 1766 3048 1772 3049
rect 1766 3044 1767 3048
rect 1771 3044 1772 3048
rect 2006 3047 2007 3051
rect 2011 3047 2012 3051
rect 2006 3046 2012 3047
rect 1766 3043 1772 3044
rect 264 2995 266 3043
rect 440 2995 442 3043
rect 616 2995 618 3043
rect 800 2995 802 3043
rect 976 2995 978 3043
rect 1144 2995 1146 3043
rect 1304 2995 1306 3043
rect 1456 2995 1458 3043
rect 1608 2995 1610 3043
rect 1768 2995 1770 3043
rect 2008 2995 2010 3046
rect 2048 3035 2050 3070
rect 2078 3068 2079 3072
rect 2083 3068 2084 3072
rect 2078 3067 2084 3068
rect 2222 3072 2228 3073
rect 2222 3068 2223 3072
rect 2227 3068 2228 3072
rect 2222 3067 2228 3068
rect 2374 3072 2380 3073
rect 2374 3068 2375 3072
rect 2379 3068 2380 3072
rect 2374 3067 2380 3068
rect 2526 3072 2532 3073
rect 2526 3068 2527 3072
rect 2531 3068 2532 3072
rect 2526 3067 2532 3068
rect 2686 3072 2692 3073
rect 2686 3068 2687 3072
rect 2691 3068 2692 3072
rect 2686 3067 2692 3068
rect 2854 3072 2860 3073
rect 2854 3068 2855 3072
rect 2859 3068 2860 3072
rect 2854 3067 2860 3068
rect 3038 3072 3044 3073
rect 3038 3068 3039 3072
rect 3043 3068 3044 3072
rect 3038 3067 3044 3068
rect 3230 3072 3236 3073
rect 3230 3068 3231 3072
rect 3235 3068 3236 3072
rect 3230 3067 3236 3068
rect 3430 3072 3436 3073
rect 3430 3068 3431 3072
rect 3435 3068 3436 3072
rect 3430 3067 3436 3068
rect 3638 3072 3644 3073
rect 3638 3068 3639 3072
rect 3643 3068 3644 3072
rect 3638 3067 3644 3068
rect 3838 3072 3844 3073
rect 3838 3068 3839 3072
rect 3843 3068 3844 3072
rect 3942 3071 3943 3075
rect 3947 3071 3948 3075
rect 3942 3070 3948 3071
rect 3838 3067 3844 3068
rect 2080 3035 2082 3067
rect 2224 3035 2226 3067
rect 2376 3035 2378 3067
rect 2528 3035 2530 3067
rect 2688 3035 2690 3067
rect 2856 3035 2858 3067
rect 3040 3035 3042 3067
rect 3232 3035 3234 3067
rect 3432 3035 3434 3067
rect 3640 3035 3642 3067
rect 3840 3035 3842 3067
rect 3944 3035 3946 3070
rect 2047 3034 2051 3035
rect 2047 3029 2051 3030
rect 2071 3034 2075 3035
rect 2071 3029 2075 3030
rect 2079 3034 2083 3035
rect 2079 3029 2083 3030
rect 2183 3034 2187 3035
rect 2183 3029 2187 3030
rect 2223 3034 2227 3035
rect 2223 3029 2227 3030
rect 2327 3034 2331 3035
rect 2327 3029 2331 3030
rect 2375 3034 2379 3035
rect 2375 3029 2379 3030
rect 2479 3034 2483 3035
rect 2479 3029 2483 3030
rect 2527 3034 2531 3035
rect 2527 3029 2531 3030
rect 2655 3034 2659 3035
rect 2655 3029 2659 3030
rect 2687 3034 2691 3035
rect 2687 3029 2691 3030
rect 2855 3034 2859 3035
rect 2855 3029 2859 3030
rect 3039 3034 3043 3035
rect 3039 3029 3043 3030
rect 3087 3034 3091 3035
rect 3087 3029 3091 3030
rect 3231 3034 3235 3035
rect 3231 3029 3235 3030
rect 3335 3034 3339 3035
rect 3335 3029 3339 3030
rect 3431 3034 3435 3035
rect 3431 3029 3435 3030
rect 3599 3034 3603 3035
rect 3599 3029 3603 3030
rect 3639 3034 3643 3035
rect 3639 3029 3643 3030
rect 3839 3034 3843 3035
rect 3839 3029 3843 3030
rect 3943 3034 3947 3035
rect 3943 3029 3947 3030
rect 2048 3002 2050 3029
rect 2072 3005 2074 3029
rect 2184 3005 2186 3029
rect 2328 3005 2330 3029
rect 2480 3005 2482 3029
rect 2656 3005 2658 3029
rect 2856 3005 2858 3029
rect 3088 3005 3090 3029
rect 3336 3005 3338 3029
rect 3600 3005 3602 3029
rect 3840 3005 3842 3029
rect 2070 3004 2076 3005
rect 2046 3001 2052 3002
rect 2046 2997 2047 3001
rect 2051 2997 2052 3001
rect 2070 3000 2071 3004
rect 2075 3000 2076 3004
rect 2070 2999 2076 3000
rect 2182 3004 2188 3005
rect 2182 3000 2183 3004
rect 2187 3000 2188 3004
rect 2182 2999 2188 3000
rect 2326 3004 2332 3005
rect 2326 3000 2327 3004
rect 2331 3000 2332 3004
rect 2326 2999 2332 3000
rect 2478 3004 2484 3005
rect 2478 3000 2479 3004
rect 2483 3000 2484 3004
rect 2478 2999 2484 3000
rect 2654 3004 2660 3005
rect 2654 3000 2655 3004
rect 2659 3000 2660 3004
rect 2654 2999 2660 3000
rect 2854 3004 2860 3005
rect 2854 3000 2855 3004
rect 2859 3000 2860 3004
rect 2854 2999 2860 3000
rect 3086 3004 3092 3005
rect 3086 3000 3087 3004
rect 3091 3000 3092 3004
rect 3086 2999 3092 3000
rect 3334 3004 3340 3005
rect 3334 3000 3335 3004
rect 3339 3000 3340 3004
rect 3334 2999 3340 3000
rect 3598 3004 3604 3005
rect 3598 3000 3599 3004
rect 3603 3000 3604 3004
rect 3598 2999 3604 3000
rect 3838 3004 3844 3005
rect 3838 3000 3839 3004
rect 3843 3000 3844 3004
rect 3944 3002 3946 3029
rect 3838 2999 3844 3000
rect 3942 3001 3948 3002
rect 2046 2996 2052 2997
rect 3942 2997 3943 3001
rect 3947 2997 3948 3001
rect 3942 2996 3948 2997
rect 111 2994 115 2995
rect 111 2989 115 2990
rect 263 2994 267 2995
rect 263 2989 267 2990
rect 343 2994 347 2995
rect 343 2989 347 2990
rect 439 2994 443 2995
rect 439 2989 443 2990
rect 543 2994 547 2995
rect 543 2989 547 2990
rect 615 2994 619 2995
rect 615 2989 619 2990
rect 655 2994 659 2995
rect 655 2989 659 2990
rect 783 2994 787 2995
rect 783 2989 787 2990
rect 799 2994 803 2995
rect 799 2989 803 2990
rect 935 2994 939 2995
rect 935 2989 939 2990
rect 975 2994 979 2995
rect 975 2989 979 2990
rect 1103 2994 1107 2995
rect 1103 2989 1107 2990
rect 1143 2994 1147 2995
rect 1143 2989 1147 2990
rect 1295 2994 1299 2995
rect 1295 2989 1299 2990
rect 1303 2994 1307 2995
rect 1303 2989 1307 2990
rect 1455 2994 1459 2995
rect 1455 2989 1459 2990
rect 1495 2994 1499 2995
rect 1495 2989 1499 2990
rect 1607 2994 1611 2995
rect 1607 2989 1611 2990
rect 1711 2994 1715 2995
rect 1711 2989 1715 2990
rect 1767 2994 1771 2995
rect 1767 2989 1771 2990
rect 1903 2994 1907 2995
rect 1903 2989 1907 2990
rect 2007 2994 2011 2995
rect 2007 2989 2011 2990
rect 112 2962 114 2989
rect 344 2965 346 2989
rect 440 2965 442 2989
rect 544 2965 546 2989
rect 656 2965 658 2989
rect 784 2965 786 2989
rect 936 2965 938 2989
rect 1104 2965 1106 2989
rect 1296 2965 1298 2989
rect 1496 2965 1498 2989
rect 1712 2965 1714 2989
rect 1904 2965 1906 2989
rect 342 2964 348 2965
rect 110 2961 116 2962
rect 110 2957 111 2961
rect 115 2957 116 2961
rect 342 2960 343 2964
rect 347 2960 348 2964
rect 342 2959 348 2960
rect 438 2964 444 2965
rect 438 2960 439 2964
rect 443 2960 444 2964
rect 438 2959 444 2960
rect 542 2964 548 2965
rect 542 2960 543 2964
rect 547 2960 548 2964
rect 542 2959 548 2960
rect 654 2964 660 2965
rect 654 2960 655 2964
rect 659 2960 660 2964
rect 654 2959 660 2960
rect 782 2964 788 2965
rect 782 2960 783 2964
rect 787 2960 788 2964
rect 782 2959 788 2960
rect 934 2964 940 2965
rect 934 2960 935 2964
rect 939 2960 940 2964
rect 934 2959 940 2960
rect 1102 2964 1108 2965
rect 1102 2960 1103 2964
rect 1107 2960 1108 2964
rect 1102 2959 1108 2960
rect 1294 2964 1300 2965
rect 1294 2960 1295 2964
rect 1299 2960 1300 2964
rect 1294 2959 1300 2960
rect 1494 2964 1500 2965
rect 1494 2960 1495 2964
rect 1499 2960 1500 2964
rect 1494 2959 1500 2960
rect 1710 2964 1716 2965
rect 1710 2960 1711 2964
rect 1715 2960 1716 2964
rect 1710 2959 1716 2960
rect 1902 2964 1908 2965
rect 1902 2960 1903 2964
rect 1907 2960 1908 2964
rect 2008 2962 2010 2989
rect 2070 2985 2076 2986
rect 2046 2984 2052 2985
rect 2046 2980 2047 2984
rect 2051 2980 2052 2984
rect 2070 2981 2071 2985
rect 2075 2981 2076 2985
rect 2070 2980 2076 2981
rect 2182 2985 2188 2986
rect 2182 2981 2183 2985
rect 2187 2981 2188 2985
rect 2182 2980 2188 2981
rect 2326 2985 2332 2986
rect 2326 2981 2327 2985
rect 2331 2981 2332 2985
rect 2326 2980 2332 2981
rect 2478 2985 2484 2986
rect 2478 2981 2479 2985
rect 2483 2981 2484 2985
rect 2478 2980 2484 2981
rect 2654 2985 2660 2986
rect 2654 2981 2655 2985
rect 2659 2981 2660 2985
rect 2654 2980 2660 2981
rect 2854 2985 2860 2986
rect 2854 2981 2855 2985
rect 2859 2981 2860 2985
rect 2854 2980 2860 2981
rect 3086 2985 3092 2986
rect 3086 2981 3087 2985
rect 3091 2981 3092 2985
rect 3086 2980 3092 2981
rect 3334 2985 3340 2986
rect 3334 2981 3335 2985
rect 3339 2981 3340 2985
rect 3334 2980 3340 2981
rect 3598 2985 3604 2986
rect 3598 2981 3599 2985
rect 3603 2981 3604 2985
rect 3598 2980 3604 2981
rect 3838 2985 3844 2986
rect 3838 2981 3839 2985
rect 3843 2981 3844 2985
rect 3838 2980 3844 2981
rect 3942 2984 3948 2985
rect 3942 2980 3943 2984
rect 3947 2980 3948 2984
rect 2046 2979 2052 2980
rect 1902 2959 1908 2960
rect 2006 2961 2012 2962
rect 110 2956 116 2957
rect 2006 2957 2007 2961
rect 2011 2957 2012 2961
rect 2006 2956 2012 2957
rect 2048 2955 2050 2979
rect 2072 2955 2074 2980
rect 2184 2955 2186 2980
rect 2328 2955 2330 2980
rect 2480 2955 2482 2980
rect 2656 2955 2658 2980
rect 2856 2955 2858 2980
rect 3088 2955 3090 2980
rect 3336 2955 3338 2980
rect 3600 2955 3602 2980
rect 3840 2955 3842 2980
rect 3942 2979 3948 2980
rect 3944 2955 3946 2979
rect 2047 2954 2051 2955
rect 2047 2949 2051 2950
rect 2071 2954 2075 2955
rect 2071 2949 2075 2950
rect 2183 2954 2187 2955
rect 2183 2949 2187 2950
rect 2263 2954 2267 2955
rect 2263 2949 2267 2950
rect 2327 2954 2331 2955
rect 2327 2949 2331 2950
rect 2479 2954 2483 2955
rect 2479 2949 2483 2950
rect 2487 2954 2491 2955
rect 2487 2949 2491 2950
rect 2655 2954 2659 2955
rect 2655 2949 2659 2950
rect 2735 2954 2739 2955
rect 2735 2949 2739 2950
rect 2855 2954 2859 2955
rect 2855 2949 2859 2950
rect 2999 2954 3003 2955
rect 2999 2949 3003 2950
rect 3087 2954 3091 2955
rect 3087 2949 3091 2950
rect 3279 2954 3283 2955
rect 3279 2949 3283 2950
rect 3335 2954 3339 2955
rect 3335 2949 3339 2950
rect 3567 2954 3571 2955
rect 3567 2949 3571 2950
rect 3599 2954 3603 2955
rect 3599 2949 3603 2950
rect 3839 2954 3843 2955
rect 3839 2949 3843 2950
rect 3943 2954 3947 2955
rect 3943 2949 3947 2950
rect 342 2945 348 2946
rect 110 2944 116 2945
rect 110 2940 111 2944
rect 115 2940 116 2944
rect 342 2941 343 2945
rect 347 2941 348 2945
rect 342 2940 348 2941
rect 438 2945 444 2946
rect 438 2941 439 2945
rect 443 2941 444 2945
rect 438 2940 444 2941
rect 542 2945 548 2946
rect 542 2941 543 2945
rect 547 2941 548 2945
rect 542 2940 548 2941
rect 654 2945 660 2946
rect 654 2941 655 2945
rect 659 2941 660 2945
rect 654 2940 660 2941
rect 782 2945 788 2946
rect 782 2941 783 2945
rect 787 2941 788 2945
rect 782 2940 788 2941
rect 934 2945 940 2946
rect 934 2941 935 2945
rect 939 2941 940 2945
rect 934 2940 940 2941
rect 1102 2945 1108 2946
rect 1102 2941 1103 2945
rect 1107 2941 1108 2945
rect 1102 2940 1108 2941
rect 1294 2945 1300 2946
rect 1294 2941 1295 2945
rect 1299 2941 1300 2945
rect 1294 2940 1300 2941
rect 1494 2945 1500 2946
rect 1494 2941 1495 2945
rect 1499 2941 1500 2945
rect 1494 2940 1500 2941
rect 1710 2945 1716 2946
rect 1710 2941 1711 2945
rect 1715 2941 1716 2945
rect 1710 2940 1716 2941
rect 1902 2945 1908 2946
rect 1902 2941 1903 2945
rect 1907 2941 1908 2945
rect 1902 2940 1908 2941
rect 2006 2944 2012 2945
rect 2006 2940 2007 2944
rect 2011 2940 2012 2944
rect 110 2939 116 2940
rect 112 2919 114 2939
rect 344 2919 346 2940
rect 440 2919 442 2940
rect 544 2919 546 2940
rect 656 2919 658 2940
rect 784 2919 786 2940
rect 936 2919 938 2940
rect 1104 2919 1106 2940
rect 1296 2919 1298 2940
rect 1496 2919 1498 2940
rect 1712 2919 1714 2940
rect 1904 2919 1906 2940
rect 2006 2939 2012 2940
rect 2008 2919 2010 2939
rect 2048 2929 2050 2949
rect 2046 2928 2052 2929
rect 2072 2928 2074 2949
rect 2264 2928 2266 2949
rect 2488 2928 2490 2949
rect 2736 2928 2738 2949
rect 3000 2928 3002 2949
rect 3280 2928 3282 2949
rect 3568 2928 3570 2949
rect 3840 2928 3842 2949
rect 3944 2929 3946 2949
rect 3942 2928 3948 2929
rect 2046 2924 2047 2928
rect 2051 2924 2052 2928
rect 2046 2923 2052 2924
rect 2070 2927 2076 2928
rect 2070 2923 2071 2927
rect 2075 2923 2076 2927
rect 2070 2922 2076 2923
rect 2262 2927 2268 2928
rect 2262 2923 2263 2927
rect 2267 2923 2268 2927
rect 2262 2922 2268 2923
rect 2486 2927 2492 2928
rect 2486 2923 2487 2927
rect 2491 2923 2492 2927
rect 2486 2922 2492 2923
rect 2734 2927 2740 2928
rect 2734 2923 2735 2927
rect 2739 2923 2740 2927
rect 2734 2922 2740 2923
rect 2998 2927 3004 2928
rect 2998 2923 2999 2927
rect 3003 2923 3004 2927
rect 2998 2922 3004 2923
rect 3278 2927 3284 2928
rect 3278 2923 3279 2927
rect 3283 2923 3284 2927
rect 3278 2922 3284 2923
rect 3566 2927 3572 2928
rect 3566 2923 3567 2927
rect 3571 2923 3572 2927
rect 3566 2922 3572 2923
rect 3838 2927 3844 2928
rect 3838 2923 3839 2927
rect 3843 2923 3844 2927
rect 3942 2924 3943 2928
rect 3947 2924 3948 2928
rect 3942 2923 3948 2924
rect 3838 2922 3844 2923
rect 111 2918 115 2919
rect 111 2913 115 2914
rect 207 2918 211 2919
rect 207 2913 211 2914
rect 327 2918 331 2919
rect 327 2913 331 2914
rect 343 2918 347 2919
rect 343 2913 347 2914
rect 439 2918 443 2919
rect 439 2913 443 2914
rect 447 2918 451 2919
rect 447 2913 451 2914
rect 543 2918 547 2919
rect 543 2913 547 2914
rect 575 2918 579 2919
rect 575 2913 579 2914
rect 655 2918 659 2919
rect 655 2913 659 2914
rect 703 2918 707 2919
rect 703 2913 707 2914
rect 783 2918 787 2919
rect 783 2913 787 2914
rect 847 2918 851 2919
rect 847 2913 851 2914
rect 935 2918 939 2919
rect 935 2913 939 2914
rect 999 2918 1003 2919
rect 999 2913 1003 2914
rect 1103 2918 1107 2919
rect 1103 2913 1107 2914
rect 1167 2918 1171 2919
rect 1167 2913 1171 2914
rect 1295 2918 1299 2919
rect 1295 2913 1299 2914
rect 1351 2918 1355 2919
rect 1351 2913 1355 2914
rect 1495 2918 1499 2919
rect 1495 2913 1499 2914
rect 1535 2918 1539 2919
rect 1535 2913 1539 2914
rect 1711 2918 1715 2919
rect 1711 2913 1715 2914
rect 1727 2918 1731 2919
rect 1727 2913 1731 2914
rect 1903 2918 1907 2919
rect 1903 2913 1907 2914
rect 2007 2918 2011 2919
rect 2007 2913 2011 2914
rect 112 2893 114 2913
rect 110 2892 116 2893
rect 208 2892 210 2913
rect 328 2892 330 2913
rect 448 2892 450 2913
rect 576 2892 578 2913
rect 704 2892 706 2913
rect 848 2892 850 2913
rect 1000 2892 1002 2913
rect 1168 2892 1170 2913
rect 1352 2892 1354 2913
rect 1536 2892 1538 2913
rect 1728 2892 1730 2913
rect 1904 2892 1906 2913
rect 2008 2893 2010 2913
rect 2046 2911 2052 2912
rect 2046 2907 2047 2911
rect 2051 2907 2052 2911
rect 3942 2911 3948 2912
rect 2046 2906 2052 2907
rect 2070 2908 2076 2909
rect 2006 2892 2012 2893
rect 110 2888 111 2892
rect 115 2888 116 2892
rect 110 2887 116 2888
rect 206 2891 212 2892
rect 206 2887 207 2891
rect 211 2887 212 2891
rect 206 2886 212 2887
rect 326 2891 332 2892
rect 326 2887 327 2891
rect 331 2887 332 2891
rect 326 2886 332 2887
rect 446 2891 452 2892
rect 446 2887 447 2891
rect 451 2887 452 2891
rect 446 2886 452 2887
rect 574 2891 580 2892
rect 574 2887 575 2891
rect 579 2887 580 2891
rect 574 2886 580 2887
rect 702 2891 708 2892
rect 702 2887 703 2891
rect 707 2887 708 2891
rect 702 2886 708 2887
rect 846 2891 852 2892
rect 846 2887 847 2891
rect 851 2887 852 2891
rect 846 2886 852 2887
rect 998 2891 1004 2892
rect 998 2887 999 2891
rect 1003 2887 1004 2891
rect 998 2886 1004 2887
rect 1166 2891 1172 2892
rect 1166 2887 1167 2891
rect 1171 2887 1172 2891
rect 1166 2886 1172 2887
rect 1350 2891 1356 2892
rect 1350 2887 1351 2891
rect 1355 2887 1356 2891
rect 1350 2886 1356 2887
rect 1534 2891 1540 2892
rect 1534 2887 1535 2891
rect 1539 2887 1540 2891
rect 1534 2886 1540 2887
rect 1726 2891 1732 2892
rect 1726 2887 1727 2891
rect 1731 2887 1732 2891
rect 1726 2886 1732 2887
rect 1902 2891 1908 2892
rect 1902 2887 1903 2891
rect 1907 2887 1908 2891
rect 2006 2888 2007 2892
rect 2011 2888 2012 2892
rect 2006 2887 2012 2888
rect 1902 2886 1908 2887
rect 110 2875 116 2876
rect 110 2871 111 2875
rect 115 2871 116 2875
rect 2006 2875 2012 2876
rect 110 2870 116 2871
rect 206 2872 212 2873
rect 112 2839 114 2870
rect 206 2868 207 2872
rect 211 2868 212 2872
rect 206 2867 212 2868
rect 326 2872 332 2873
rect 326 2868 327 2872
rect 331 2868 332 2872
rect 326 2867 332 2868
rect 446 2872 452 2873
rect 446 2868 447 2872
rect 451 2868 452 2872
rect 446 2867 452 2868
rect 574 2872 580 2873
rect 574 2868 575 2872
rect 579 2868 580 2872
rect 574 2867 580 2868
rect 702 2872 708 2873
rect 702 2868 703 2872
rect 707 2868 708 2872
rect 702 2867 708 2868
rect 846 2872 852 2873
rect 846 2868 847 2872
rect 851 2868 852 2872
rect 846 2867 852 2868
rect 998 2872 1004 2873
rect 998 2868 999 2872
rect 1003 2868 1004 2872
rect 998 2867 1004 2868
rect 1166 2872 1172 2873
rect 1166 2868 1167 2872
rect 1171 2868 1172 2872
rect 1166 2867 1172 2868
rect 1350 2872 1356 2873
rect 1350 2868 1351 2872
rect 1355 2868 1356 2872
rect 1350 2867 1356 2868
rect 1534 2872 1540 2873
rect 1534 2868 1535 2872
rect 1539 2868 1540 2872
rect 1534 2867 1540 2868
rect 1726 2872 1732 2873
rect 1726 2868 1727 2872
rect 1731 2868 1732 2872
rect 1726 2867 1732 2868
rect 1902 2872 1908 2873
rect 1902 2868 1903 2872
rect 1907 2868 1908 2872
rect 2006 2871 2007 2875
rect 2011 2871 2012 2875
rect 2048 2871 2050 2906
rect 2070 2904 2071 2908
rect 2075 2904 2076 2908
rect 2070 2903 2076 2904
rect 2262 2908 2268 2909
rect 2262 2904 2263 2908
rect 2267 2904 2268 2908
rect 2262 2903 2268 2904
rect 2486 2908 2492 2909
rect 2486 2904 2487 2908
rect 2491 2904 2492 2908
rect 2486 2903 2492 2904
rect 2734 2908 2740 2909
rect 2734 2904 2735 2908
rect 2739 2904 2740 2908
rect 2734 2903 2740 2904
rect 2998 2908 3004 2909
rect 2998 2904 2999 2908
rect 3003 2904 3004 2908
rect 2998 2903 3004 2904
rect 3278 2908 3284 2909
rect 3278 2904 3279 2908
rect 3283 2904 3284 2908
rect 3278 2903 3284 2904
rect 3566 2908 3572 2909
rect 3566 2904 3567 2908
rect 3571 2904 3572 2908
rect 3566 2903 3572 2904
rect 3838 2908 3844 2909
rect 3838 2904 3839 2908
rect 3843 2904 3844 2908
rect 3942 2907 3943 2911
rect 3947 2907 3948 2911
rect 3942 2906 3948 2907
rect 3838 2903 3844 2904
rect 2072 2871 2074 2903
rect 2264 2871 2266 2903
rect 2488 2871 2490 2903
rect 2736 2871 2738 2903
rect 3000 2871 3002 2903
rect 3280 2871 3282 2903
rect 3568 2871 3570 2903
rect 3840 2871 3842 2903
rect 3944 2871 3946 2906
rect 2006 2870 2012 2871
rect 2047 2870 2051 2871
rect 1902 2867 1908 2868
rect 208 2839 210 2867
rect 328 2839 330 2867
rect 448 2839 450 2867
rect 576 2839 578 2867
rect 704 2839 706 2867
rect 848 2839 850 2867
rect 1000 2839 1002 2867
rect 1168 2839 1170 2867
rect 1352 2839 1354 2867
rect 1536 2839 1538 2867
rect 1728 2839 1730 2867
rect 1904 2839 1906 2867
rect 2008 2839 2010 2870
rect 2047 2865 2051 2866
rect 2071 2870 2075 2871
rect 2071 2865 2075 2866
rect 2263 2870 2267 2871
rect 2263 2865 2267 2866
rect 2487 2870 2491 2871
rect 2487 2865 2491 2866
rect 2671 2870 2675 2871
rect 2671 2865 2675 2866
rect 2735 2870 2739 2871
rect 2735 2865 2739 2866
rect 2887 2870 2891 2871
rect 2887 2865 2891 2866
rect 2999 2870 3003 2871
rect 2999 2865 3003 2866
rect 3095 2870 3099 2871
rect 3095 2865 3099 2866
rect 3279 2870 3283 2871
rect 3279 2865 3283 2866
rect 3287 2870 3291 2871
rect 3287 2865 3291 2866
rect 3479 2870 3483 2871
rect 3479 2865 3483 2866
rect 3567 2870 3571 2871
rect 3567 2865 3571 2866
rect 3671 2870 3675 2871
rect 3671 2865 3675 2866
rect 3839 2870 3843 2871
rect 3839 2865 3843 2866
rect 3943 2870 3947 2871
rect 3943 2865 3947 2866
rect 111 2838 115 2839
rect 111 2833 115 2834
rect 135 2838 139 2839
rect 135 2833 139 2834
rect 207 2838 211 2839
rect 207 2833 211 2834
rect 247 2838 251 2839
rect 247 2833 251 2834
rect 327 2838 331 2839
rect 327 2833 331 2834
rect 399 2838 403 2839
rect 399 2833 403 2834
rect 447 2838 451 2839
rect 447 2833 451 2834
rect 551 2838 555 2839
rect 551 2833 555 2834
rect 575 2838 579 2839
rect 575 2833 579 2834
rect 703 2838 707 2839
rect 703 2833 707 2834
rect 711 2838 715 2839
rect 711 2833 715 2834
rect 847 2838 851 2839
rect 847 2833 851 2834
rect 879 2838 883 2839
rect 879 2833 883 2834
rect 999 2838 1003 2839
rect 999 2833 1003 2834
rect 1047 2838 1051 2839
rect 1047 2833 1051 2834
rect 1167 2838 1171 2839
rect 1167 2833 1171 2834
rect 1223 2838 1227 2839
rect 1223 2833 1227 2834
rect 1351 2838 1355 2839
rect 1351 2833 1355 2834
rect 1399 2838 1403 2839
rect 1399 2833 1403 2834
rect 1535 2838 1539 2839
rect 1535 2833 1539 2834
rect 1575 2838 1579 2839
rect 1575 2833 1579 2834
rect 1727 2838 1731 2839
rect 1727 2833 1731 2834
rect 1751 2838 1755 2839
rect 1751 2833 1755 2834
rect 1903 2838 1907 2839
rect 1903 2833 1907 2834
rect 2007 2838 2011 2839
rect 2048 2838 2050 2865
rect 2672 2841 2674 2865
rect 2888 2841 2890 2865
rect 3096 2841 3098 2865
rect 3288 2841 3290 2865
rect 3480 2841 3482 2865
rect 3672 2841 3674 2865
rect 3840 2841 3842 2865
rect 2670 2840 2676 2841
rect 2007 2833 2011 2834
rect 2046 2837 2052 2838
rect 2046 2833 2047 2837
rect 2051 2833 2052 2837
rect 2670 2836 2671 2840
rect 2675 2836 2676 2840
rect 2670 2835 2676 2836
rect 2886 2840 2892 2841
rect 2886 2836 2887 2840
rect 2891 2836 2892 2840
rect 2886 2835 2892 2836
rect 3094 2840 3100 2841
rect 3094 2836 3095 2840
rect 3099 2836 3100 2840
rect 3094 2835 3100 2836
rect 3286 2840 3292 2841
rect 3286 2836 3287 2840
rect 3291 2836 3292 2840
rect 3286 2835 3292 2836
rect 3478 2840 3484 2841
rect 3478 2836 3479 2840
rect 3483 2836 3484 2840
rect 3478 2835 3484 2836
rect 3670 2840 3676 2841
rect 3670 2836 3671 2840
rect 3675 2836 3676 2840
rect 3670 2835 3676 2836
rect 3838 2840 3844 2841
rect 3838 2836 3839 2840
rect 3843 2836 3844 2840
rect 3944 2838 3946 2865
rect 3838 2835 3844 2836
rect 3942 2837 3948 2838
rect 112 2806 114 2833
rect 136 2809 138 2833
rect 248 2809 250 2833
rect 400 2809 402 2833
rect 552 2809 554 2833
rect 712 2809 714 2833
rect 880 2809 882 2833
rect 1048 2809 1050 2833
rect 1224 2809 1226 2833
rect 1400 2809 1402 2833
rect 1576 2809 1578 2833
rect 1752 2809 1754 2833
rect 1904 2809 1906 2833
rect 134 2808 140 2809
rect 110 2805 116 2806
rect 110 2801 111 2805
rect 115 2801 116 2805
rect 134 2804 135 2808
rect 139 2804 140 2808
rect 134 2803 140 2804
rect 246 2808 252 2809
rect 246 2804 247 2808
rect 251 2804 252 2808
rect 246 2803 252 2804
rect 398 2808 404 2809
rect 398 2804 399 2808
rect 403 2804 404 2808
rect 398 2803 404 2804
rect 550 2808 556 2809
rect 550 2804 551 2808
rect 555 2804 556 2808
rect 550 2803 556 2804
rect 710 2808 716 2809
rect 710 2804 711 2808
rect 715 2804 716 2808
rect 710 2803 716 2804
rect 878 2808 884 2809
rect 878 2804 879 2808
rect 883 2804 884 2808
rect 878 2803 884 2804
rect 1046 2808 1052 2809
rect 1046 2804 1047 2808
rect 1051 2804 1052 2808
rect 1046 2803 1052 2804
rect 1222 2808 1228 2809
rect 1222 2804 1223 2808
rect 1227 2804 1228 2808
rect 1222 2803 1228 2804
rect 1398 2808 1404 2809
rect 1398 2804 1399 2808
rect 1403 2804 1404 2808
rect 1398 2803 1404 2804
rect 1574 2808 1580 2809
rect 1574 2804 1575 2808
rect 1579 2804 1580 2808
rect 1574 2803 1580 2804
rect 1750 2808 1756 2809
rect 1750 2804 1751 2808
rect 1755 2804 1756 2808
rect 1750 2803 1756 2804
rect 1902 2808 1908 2809
rect 1902 2804 1903 2808
rect 1907 2804 1908 2808
rect 2008 2806 2010 2833
rect 2046 2832 2052 2833
rect 3942 2833 3943 2837
rect 3947 2833 3948 2837
rect 3942 2832 3948 2833
rect 2670 2821 2676 2822
rect 2046 2820 2052 2821
rect 2046 2816 2047 2820
rect 2051 2816 2052 2820
rect 2670 2817 2671 2821
rect 2675 2817 2676 2821
rect 2670 2816 2676 2817
rect 2886 2821 2892 2822
rect 2886 2817 2887 2821
rect 2891 2817 2892 2821
rect 2886 2816 2892 2817
rect 3094 2821 3100 2822
rect 3094 2817 3095 2821
rect 3099 2817 3100 2821
rect 3094 2816 3100 2817
rect 3286 2821 3292 2822
rect 3286 2817 3287 2821
rect 3291 2817 3292 2821
rect 3286 2816 3292 2817
rect 3478 2821 3484 2822
rect 3478 2817 3479 2821
rect 3483 2817 3484 2821
rect 3478 2816 3484 2817
rect 3670 2821 3676 2822
rect 3670 2817 3671 2821
rect 3675 2817 3676 2821
rect 3670 2816 3676 2817
rect 3838 2821 3844 2822
rect 3838 2817 3839 2821
rect 3843 2817 3844 2821
rect 3838 2816 3844 2817
rect 3942 2820 3948 2821
rect 3942 2816 3943 2820
rect 3947 2816 3948 2820
rect 2046 2815 2052 2816
rect 1902 2803 1908 2804
rect 2006 2805 2012 2806
rect 110 2800 116 2801
rect 2006 2801 2007 2805
rect 2011 2801 2012 2805
rect 2006 2800 2012 2801
rect 2048 2795 2050 2815
rect 2672 2795 2674 2816
rect 2888 2795 2890 2816
rect 3096 2795 3098 2816
rect 3288 2795 3290 2816
rect 3480 2795 3482 2816
rect 3672 2795 3674 2816
rect 3840 2795 3842 2816
rect 3942 2815 3948 2816
rect 3944 2795 3946 2815
rect 2047 2794 2051 2795
rect 134 2789 140 2790
rect 110 2788 116 2789
rect 110 2784 111 2788
rect 115 2784 116 2788
rect 134 2785 135 2789
rect 139 2785 140 2789
rect 134 2784 140 2785
rect 246 2789 252 2790
rect 246 2785 247 2789
rect 251 2785 252 2789
rect 246 2784 252 2785
rect 398 2789 404 2790
rect 398 2785 399 2789
rect 403 2785 404 2789
rect 398 2784 404 2785
rect 550 2789 556 2790
rect 550 2785 551 2789
rect 555 2785 556 2789
rect 550 2784 556 2785
rect 710 2789 716 2790
rect 710 2785 711 2789
rect 715 2785 716 2789
rect 710 2784 716 2785
rect 878 2789 884 2790
rect 878 2785 879 2789
rect 883 2785 884 2789
rect 878 2784 884 2785
rect 1046 2789 1052 2790
rect 1046 2785 1047 2789
rect 1051 2785 1052 2789
rect 1046 2784 1052 2785
rect 1222 2789 1228 2790
rect 1222 2785 1223 2789
rect 1227 2785 1228 2789
rect 1222 2784 1228 2785
rect 1398 2789 1404 2790
rect 1398 2785 1399 2789
rect 1403 2785 1404 2789
rect 1398 2784 1404 2785
rect 1574 2789 1580 2790
rect 1574 2785 1575 2789
rect 1579 2785 1580 2789
rect 1574 2784 1580 2785
rect 1750 2789 1756 2790
rect 1750 2785 1751 2789
rect 1755 2785 1756 2789
rect 1750 2784 1756 2785
rect 1902 2789 1908 2790
rect 2047 2789 2051 2790
rect 2071 2794 2075 2795
rect 2071 2789 2075 2790
rect 2199 2794 2203 2795
rect 2199 2789 2203 2790
rect 2343 2794 2347 2795
rect 2343 2789 2347 2790
rect 2479 2794 2483 2795
rect 2479 2789 2483 2790
rect 2607 2794 2611 2795
rect 2607 2789 2611 2790
rect 2671 2794 2675 2795
rect 2671 2789 2675 2790
rect 2727 2794 2731 2795
rect 2727 2789 2731 2790
rect 2839 2794 2843 2795
rect 2839 2789 2843 2790
rect 2887 2794 2891 2795
rect 2887 2789 2891 2790
rect 2943 2794 2947 2795
rect 2943 2789 2947 2790
rect 3047 2794 3051 2795
rect 3047 2789 3051 2790
rect 3095 2794 3099 2795
rect 3095 2789 3099 2790
rect 3143 2794 3147 2795
rect 3143 2789 3147 2790
rect 3239 2794 3243 2795
rect 3239 2789 3243 2790
rect 3287 2794 3291 2795
rect 3287 2789 3291 2790
rect 3343 2794 3347 2795
rect 3343 2789 3347 2790
rect 3447 2794 3451 2795
rect 3447 2789 3451 2790
rect 3479 2794 3483 2795
rect 3479 2789 3483 2790
rect 3551 2794 3555 2795
rect 3551 2789 3555 2790
rect 3647 2794 3651 2795
rect 3647 2789 3651 2790
rect 3671 2794 3675 2795
rect 3671 2789 3675 2790
rect 3743 2794 3747 2795
rect 3743 2789 3747 2790
rect 3839 2794 3843 2795
rect 3839 2789 3843 2790
rect 3943 2794 3947 2795
rect 3943 2789 3947 2790
rect 1902 2785 1903 2789
rect 1907 2785 1908 2789
rect 1902 2784 1908 2785
rect 2006 2788 2012 2789
rect 2006 2784 2007 2788
rect 2011 2784 2012 2788
rect 110 2783 116 2784
rect 112 2755 114 2783
rect 136 2755 138 2784
rect 248 2755 250 2784
rect 400 2755 402 2784
rect 552 2755 554 2784
rect 712 2755 714 2784
rect 880 2755 882 2784
rect 1048 2755 1050 2784
rect 1224 2755 1226 2784
rect 1400 2755 1402 2784
rect 1576 2755 1578 2784
rect 1752 2755 1754 2784
rect 1904 2755 1906 2784
rect 2006 2783 2012 2784
rect 2008 2755 2010 2783
rect 2048 2769 2050 2789
rect 2046 2768 2052 2769
rect 2072 2768 2074 2789
rect 2200 2768 2202 2789
rect 2344 2768 2346 2789
rect 2480 2768 2482 2789
rect 2608 2768 2610 2789
rect 2728 2768 2730 2789
rect 2840 2768 2842 2789
rect 2944 2768 2946 2789
rect 3048 2768 3050 2789
rect 3144 2768 3146 2789
rect 3240 2768 3242 2789
rect 3344 2768 3346 2789
rect 3448 2768 3450 2789
rect 3552 2768 3554 2789
rect 3648 2768 3650 2789
rect 3744 2768 3746 2789
rect 3840 2768 3842 2789
rect 3944 2769 3946 2789
rect 3942 2768 3948 2769
rect 2046 2764 2047 2768
rect 2051 2764 2052 2768
rect 2046 2763 2052 2764
rect 2070 2767 2076 2768
rect 2070 2763 2071 2767
rect 2075 2763 2076 2767
rect 2070 2762 2076 2763
rect 2198 2767 2204 2768
rect 2198 2763 2199 2767
rect 2203 2763 2204 2767
rect 2198 2762 2204 2763
rect 2342 2767 2348 2768
rect 2342 2763 2343 2767
rect 2347 2763 2348 2767
rect 2342 2762 2348 2763
rect 2478 2767 2484 2768
rect 2478 2763 2479 2767
rect 2483 2763 2484 2767
rect 2478 2762 2484 2763
rect 2606 2767 2612 2768
rect 2606 2763 2607 2767
rect 2611 2763 2612 2767
rect 2606 2762 2612 2763
rect 2726 2767 2732 2768
rect 2726 2763 2727 2767
rect 2731 2763 2732 2767
rect 2726 2762 2732 2763
rect 2838 2767 2844 2768
rect 2838 2763 2839 2767
rect 2843 2763 2844 2767
rect 2838 2762 2844 2763
rect 2942 2767 2948 2768
rect 2942 2763 2943 2767
rect 2947 2763 2948 2767
rect 2942 2762 2948 2763
rect 3046 2767 3052 2768
rect 3046 2763 3047 2767
rect 3051 2763 3052 2767
rect 3046 2762 3052 2763
rect 3142 2767 3148 2768
rect 3142 2763 3143 2767
rect 3147 2763 3148 2767
rect 3142 2762 3148 2763
rect 3238 2767 3244 2768
rect 3238 2763 3239 2767
rect 3243 2763 3244 2767
rect 3238 2762 3244 2763
rect 3342 2767 3348 2768
rect 3342 2763 3343 2767
rect 3347 2763 3348 2767
rect 3342 2762 3348 2763
rect 3446 2767 3452 2768
rect 3446 2763 3447 2767
rect 3451 2763 3452 2767
rect 3446 2762 3452 2763
rect 3550 2767 3556 2768
rect 3550 2763 3551 2767
rect 3555 2763 3556 2767
rect 3550 2762 3556 2763
rect 3646 2767 3652 2768
rect 3646 2763 3647 2767
rect 3651 2763 3652 2767
rect 3646 2762 3652 2763
rect 3742 2767 3748 2768
rect 3742 2763 3743 2767
rect 3747 2763 3748 2767
rect 3742 2762 3748 2763
rect 3838 2767 3844 2768
rect 3838 2763 3839 2767
rect 3843 2763 3844 2767
rect 3942 2764 3943 2768
rect 3947 2764 3948 2768
rect 3942 2763 3948 2764
rect 3838 2762 3844 2763
rect 111 2754 115 2755
rect 111 2749 115 2750
rect 135 2754 139 2755
rect 135 2749 139 2750
rect 247 2754 251 2755
rect 247 2749 251 2750
rect 255 2754 259 2755
rect 255 2749 259 2750
rect 399 2754 403 2755
rect 399 2749 403 2750
rect 407 2754 411 2755
rect 407 2749 411 2750
rect 551 2754 555 2755
rect 551 2749 555 2750
rect 575 2754 579 2755
rect 575 2749 579 2750
rect 711 2754 715 2755
rect 711 2749 715 2750
rect 743 2754 747 2755
rect 743 2749 747 2750
rect 879 2754 883 2755
rect 879 2749 883 2750
rect 919 2754 923 2755
rect 919 2749 923 2750
rect 1047 2754 1051 2755
rect 1047 2749 1051 2750
rect 1087 2754 1091 2755
rect 1087 2749 1091 2750
rect 1223 2754 1227 2755
rect 1223 2749 1227 2750
rect 1255 2754 1259 2755
rect 1255 2749 1259 2750
rect 1399 2754 1403 2755
rect 1399 2749 1403 2750
rect 1423 2754 1427 2755
rect 1423 2749 1427 2750
rect 1575 2754 1579 2755
rect 1575 2749 1579 2750
rect 1599 2754 1603 2755
rect 1599 2749 1603 2750
rect 1751 2754 1755 2755
rect 1751 2749 1755 2750
rect 1903 2754 1907 2755
rect 1903 2749 1907 2750
rect 2007 2754 2011 2755
rect 2007 2749 2011 2750
rect 2046 2751 2052 2752
rect 112 2729 114 2749
rect 110 2728 116 2729
rect 136 2728 138 2749
rect 256 2728 258 2749
rect 408 2728 410 2749
rect 576 2728 578 2749
rect 744 2728 746 2749
rect 920 2728 922 2749
rect 1088 2728 1090 2749
rect 1256 2728 1258 2749
rect 1424 2728 1426 2749
rect 1600 2728 1602 2749
rect 2008 2729 2010 2749
rect 2046 2747 2047 2751
rect 2051 2747 2052 2751
rect 3942 2751 3948 2752
rect 2046 2746 2052 2747
rect 2070 2748 2076 2749
rect 2006 2728 2012 2729
rect 110 2724 111 2728
rect 115 2724 116 2728
rect 110 2723 116 2724
rect 134 2727 140 2728
rect 134 2723 135 2727
rect 139 2723 140 2727
rect 134 2722 140 2723
rect 254 2727 260 2728
rect 254 2723 255 2727
rect 259 2723 260 2727
rect 254 2722 260 2723
rect 406 2727 412 2728
rect 406 2723 407 2727
rect 411 2723 412 2727
rect 406 2722 412 2723
rect 574 2727 580 2728
rect 574 2723 575 2727
rect 579 2723 580 2727
rect 574 2722 580 2723
rect 742 2727 748 2728
rect 742 2723 743 2727
rect 747 2723 748 2727
rect 742 2722 748 2723
rect 918 2727 924 2728
rect 918 2723 919 2727
rect 923 2723 924 2727
rect 918 2722 924 2723
rect 1086 2727 1092 2728
rect 1086 2723 1087 2727
rect 1091 2723 1092 2727
rect 1086 2722 1092 2723
rect 1254 2727 1260 2728
rect 1254 2723 1255 2727
rect 1259 2723 1260 2727
rect 1254 2722 1260 2723
rect 1422 2727 1428 2728
rect 1422 2723 1423 2727
rect 1427 2723 1428 2727
rect 1422 2722 1428 2723
rect 1598 2727 1604 2728
rect 1598 2723 1599 2727
rect 1603 2723 1604 2727
rect 2006 2724 2007 2728
rect 2011 2724 2012 2728
rect 2006 2723 2012 2724
rect 1598 2722 1604 2723
rect 110 2711 116 2712
rect 110 2707 111 2711
rect 115 2707 116 2711
rect 2006 2711 2012 2712
rect 110 2706 116 2707
rect 134 2708 140 2709
rect 112 2679 114 2706
rect 134 2704 135 2708
rect 139 2704 140 2708
rect 134 2703 140 2704
rect 254 2708 260 2709
rect 254 2704 255 2708
rect 259 2704 260 2708
rect 254 2703 260 2704
rect 406 2708 412 2709
rect 406 2704 407 2708
rect 411 2704 412 2708
rect 406 2703 412 2704
rect 574 2708 580 2709
rect 574 2704 575 2708
rect 579 2704 580 2708
rect 574 2703 580 2704
rect 742 2708 748 2709
rect 742 2704 743 2708
rect 747 2704 748 2708
rect 742 2703 748 2704
rect 918 2708 924 2709
rect 918 2704 919 2708
rect 923 2704 924 2708
rect 918 2703 924 2704
rect 1086 2708 1092 2709
rect 1086 2704 1087 2708
rect 1091 2704 1092 2708
rect 1086 2703 1092 2704
rect 1254 2708 1260 2709
rect 1254 2704 1255 2708
rect 1259 2704 1260 2708
rect 1254 2703 1260 2704
rect 1422 2708 1428 2709
rect 1422 2704 1423 2708
rect 1427 2704 1428 2708
rect 1422 2703 1428 2704
rect 1598 2708 1604 2709
rect 1598 2704 1599 2708
rect 1603 2704 1604 2708
rect 2006 2707 2007 2711
rect 2011 2707 2012 2711
rect 2006 2706 2012 2707
rect 1598 2703 1604 2704
rect 136 2679 138 2703
rect 256 2679 258 2703
rect 408 2679 410 2703
rect 576 2679 578 2703
rect 744 2679 746 2703
rect 920 2679 922 2703
rect 1088 2679 1090 2703
rect 1256 2679 1258 2703
rect 1424 2679 1426 2703
rect 1600 2679 1602 2703
rect 2008 2679 2010 2706
rect 2048 2699 2050 2746
rect 2070 2744 2071 2748
rect 2075 2744 2076 2748
rect 2070 2743 2076 2744
rect 2198 2748 2204 2749
rect 2198 2744 2199 2748
rect 2203 2744 2204 2748
rect 2198 2743 2204 2744
rect 2342 2748 2348 2749
rect 2342 2744 2343 2748
rect 2347 2744 2348 2748
rect 2342 2743 2348 2744
rect 2478 2748 2484 2749
rect 2478 2744 2479 2748
rect 2483 2744 2484 2748
rect 2478 2743 2484 2744
rect 2606 2748 2612 2749
rect 2606 2744 2607 2748
rect 2611 2744 2612 2748
rect 2606 2743 2612 2744
rect 2726 2748 2732 2749
rect 2726 2744 2727 2748
rect 2731 2744 2732 2748
rect 2726 2743 2732 2744
rect 2838 2748 2844 2749
rect 2838 2744 2839 2748
rect 2843 2744 2844 2748
rect 2838 2743 2844 2744
rect 2942 2748 2948 2749
rect 2942 2744 2943 2748
rect 2947 2744 2948 2748
rect 2942 2743 2948 2744
rect 3046 2748 3052 2749
rect 3046 2744 3047 2748
rect 3051 2744 3052 2748
rect 3046 2743 3052 2744
rect 3142 2748 3148 2749
rect 3142 2744 3143 2748
rect 3147 2744 3148 2748
rect 3142 2743 3148 2744
rect 3238 2748 3244 2749
rect 3238 2744 3239 2748
rect 3243 2744 3244 2748
rect 3238 2743 3244 2744
rect 3342 2748 3348 2749
rect 3342 2744 3343 2748
rect 3347 2744 3348 2748
rect 3342 2743 3348 2744
rect 3446 2748 3452 2749
rect 3446 2744 3447 2748
rect 3451 2744 3452 2748
rect 3446 2743 3452 2744
rect 3550 2748 3556 2749
rect 3550 2744 3551 2748
rect 3555 2744 3556 2748
rect 3550 2743 3556 2744
rect 3646 2748 3652 2749
rect 3646 2744 3647 2748
rect 3651 2744 3652 2748
rect 3646 2743 3652 2744
rect 3742 2748 3748 2749
rect 3742 2744 3743 2748
rect 3747 2744 3748 2748
rect 3742 2743 3748 2744
rect 3838 2748 3844 2749
rect 3838 2744 3839 2748
rect 3843 2744 3844 2748
rect 3942 2747 3943 2751
rect 3947 2747 3948 2751
rect 3942 2746 3948 2747
rect 3838 2743 3844 2744
rect 2072 2699 2074 2743
rect 2200 2699 2202 2743
rect 2344 2699 2346 2743
rect 2480 2699 2482 2743
rect 2608 2699 2610 2743
rect 2728 2699 2730 2743
rect 2840 2699 2842 2743
rect 2944 2699 2946 2743
rect 3048 2699 3050 2743
rect 3144 2699 3146 2743
rect 3240 2699 3242 2743
rect 3344 2699 3346 2743
rect 3448 2699 3450 2743
rect 3552 2699 3554 2743
rect 3648 2699 3650 2743
rect 3744 2699 3746 2743
rect 3840 2699 3842 2743
rect 3944 2699 3946 2746
rect 2047 2698 2051 2699
rect 2047 2693 2051 2694
rect 2071 2698 2075 2699
rect 2071 2693 2075 2694
rect 2095 2698 2099 2699
rect 2095 2693 2099 2694
rect 2199 2698 2203 2699
rect 2199 2693 2203 2694
rect 2263 2698 2267 2699
rect 2263 2693 2267 2694
rect 2343 2698 2347 2699
rect 2343 2693 2347 2694
rect 2439 2698 2443 2699
rect 2439 2693 2443 2694
rect 2479 2698 2483 2699
rect 2479 2693 2483 2694
rect 2607 2698 2611 2699
rect 2607 2693 2611 2694
rect 2615 2698 2619 2699
rect 2615 2693 2619 2694
rect 2727 2698 2731 2699
rect 2727 2693 2731 2694
rect 2783 2698 2787 2699
rect 2783 2693 2787 2694
rect 2839 2698 2843 2699
rect 2839 2693 2843 2694
rect 2943 2698 2947 2699
rect 2943 2693 2947 2694
rect 3047 2698 3051 2699
rect 3047 2693 3051 2694
rect 3095 2698 3099 2699
rect 3095 2693 3099 2694
rect 3143 2698 3147 2699
rect 3143 2693 3147 2694
rect 3239 2698 3243 2699
rect 3239 2693 3243 2694
rect 3343 2698 3347 2699
rect 3343 2693 3347 2694
rect 3383 2698 3387 2699
rect 3383 2693 3387 2694
rect 3447 2698 3451 2699
rect 3447 2693 3451 2694
rect 3535 2698 3539 2699
rect 3535 2693 3539 2694
rect 3551 2698 3555 2699
rect 3551 2693 3555 2694
rect 3647 2698 3651 2699
rect 3647 2693 3651 2694
rect 3743 2698 3747 2699
rect 3743 2693 3747 2694
rect 3839 2698 3843 2699
rect 3839 2693 3843 2694
rect 3943 2698 3947 2699
rect 3943 2693 3947 2694
rect 111 2678 115 2679
rect 111 2673 115 2674
rect 135 2678 139 2679
rect 135 2673 139 2674
rect 167 2678 171 2679
rect 167 2673 171 2674
rect 255 2678 259 2679
rect 255 2673 259 2674
rect 359 2678 363 2679
rect 359 2673 363 2674
rect 407 2678 411 2679
rect 407 2673 411 2674
rect 559 2678 563 2679
rect 559 2673 563 2674
rect 575 2678 579 2679
rect 575 2673 579 2674
rect 743 2678 747 2679
rect 743 2673 747 2674
rect 759 2678 763 2679
rect 759 2673 763 2674
rect 919 2678 923 2679
rect 919 2673 923 2674
rect 951 2678 955 2679
rect 951 2673 955 2674
rect 1087 2678 1091 2679
rect 1087 2673 1091 2674
rect 1143 2678 1147 2679
rect 1143 2673 1147 2674
rect 1255 2678 1259 2679
rect 1255 2673 1259 2674
rect 1327 2678 1331 2679
rect 1327 2673 1331 2674
rect 1423 2678 1427 2679
rect 1423 2673 1427 2674
rect 1511 2678 1515 2679
rect 1511 2673 1515 2674
rect 1599 2678 1603 2679
rect 1599 2673 1603 2674
rect 1703 2678 1707 2679
rect 1703 2673 1707 2674
rect 2007 2678 2011 2679
rect 2007 2673 2011 2674
rect 112 2646 114 2673
rect 168 2649 170 2673
rect 360 2649 362 2673
rect 560 2649 562 2673
rect 760 2649 762 2673
rect 952 2649 954 2673
rect 1144 2649 1146 2673
rect 1328 2649 1330 2673
rect 1512 2649 1514 2673
rect 1704 2649 1706 2673
rect 166 2648 172 2649
rect 110 2645 116 2646
rect 110 2641 111 2645
rect 115 2641 116 2645
rect 166 2644 167 2648
rect 171 2644 172 2648
rect 166 2643 172 2644
rect 358 2648 364 2649
rect 358 2644 359 2648
rect 363 2644 364 2648
rect 358 2643 364 2644
rect 558 2648 564 2649
rect 558 2644 559 2648
rect 563 2644 564 2648
rect 558 2643 564 2644
rect 758 2648 764 2649
rect 758 2644 759 2648
rect 763 2644 764 2648
rect 758 2643 764 2644
rect 950 2648 956 2649
rect 950 2644 951 2648
rect 955 2644 956 2648
rect 950 2643 956 2644
rect 1142 2648 1148 2649
rect 1142 2644 1143 2648
rect 1147 2644 1148 2648
rect 1142 2643 1148 2644
rect 1326 2648 1332 2649
rect 1326 2644 1327 2648
rect 1331 2644 1332 2648
rect 1326 2643 1332 2644
rect 1510 2648 1516 2649
rect 1510 2644 1511 2648
rect 1515 2644 1516 2648
rect 1510 2643 1516 2644
rect 1702 2648 1708 2649
rect 1702 2644 1703 2648
rect 1707 2644 1708 2648
rect 2008 2646 2010 2673
rect 2048 2666 2050 2693
rect 2096 2669 2098 2693
rect 2264 2669 2266 2693
rect 2440 2669 2442 2693
rect 2616 2669 2618 2693
rect 2784 2669 2786 2693
rect 2944 2669 2946 2693
rect 3096 2669 3098 2693
rect 3240 2669 3242 2693
rect 3384 2669 3386 2693
rect 3536 2669 3538 2693
rect 2094 2668 2100 2669
rect 2046 2665 2052 2666
rect 2046 2661 2047 2665
rect 2051 2661 2052 2665
rect 2094 2664 2095 2668
rect 2099 2664 2100 2668
rect 2094 2663 2100 2664
rect 2262 2668 2268 2669
rect 2262 2664 2263 2668
rect 2267 2664 2268 2668
rect 2262 2663 2268 2664
rect 2438 2668 2444 2669
rect 2438 2664 2439 2668
rect 2443 2664 2444 2668
rect 2438 2663 2444 2664
rect 2614 2668 2620 2669
rect 2614 2664 2615 2668
rect 2619 2664 2620 2668
rect 2614 2663 2620 2664
rect 2782 2668 2788 2669
rect 2782 2664 2783 2668
rect 2787 2664 2788 2668
rect 2782 2663 2788 2664
rect 2942 2668 2948 2669
rect 2942 2664 2943 2668
rect 2947 2664 2948 2668
rect 2942 2663 2948 2664
rect 3094 2668 3100 2669
rect 3094 2664 3095 2668
rect 3099 2664 3100 2668
rect 3094 2663 3100 2664
rect 3238 2668 3244 2669
rect 3238 2664 3239 2668
rect 3243 2664 3244 2668
rect 3238 2663 3244 2664
rect 3382 2668 3388 2669
rect 3382 2664 3383 2668
rect 3387 2664 3388 2668
rect 3382 2663 3388 2664
rect 3534 2668 3540 2669
rect 3534 2664 3535 2668
rect 3539 2664 3540 2668
rect 3944 2666 3946 2693
rect 3534 2663 3540 2664
rect 3942 2665 3948 2666
rect 2046 2660 2052 2661
rect 3942 2661 3943 2665
rect 3947 2661 3948 2665
rect 3942 2660 3948 2661
rect 2094 2649 2100 2650
rect 2046 2648 2052 2649
rect 1702 2643 1708 2644
rect 2006 2645 2012 2646
rect 110 2640 116 2641
rect 2006 2641 2007 2645
rect 2011 2641 2012 2645
rect 2046 2644 2047 2648
rect 2051 2644 2052 2648
rect 2094 2645 2095 2649
rect 2099 2645 2100 2649
rect 2094 2644 2100 2645
rect 2262 2649 2268 2650
rect 2262 2645 2263 2649
rect 2267 2645 2268 2649
rect 2262 2644 2268 2645
rect 2438 2649 2444 2650
rect 2438 2645 2439 2649
rect 2443 2645 2444 2649
rect 2438 2644 2444 2645
rect 2614 2649 2620 2650
rect 2614 2645 2615 2649
rect 2619 2645 2620 2649
rect 2614 2644 2620 2645
rect 2782 2649 2788 2650
rect 2782 2645 2783 2649
rect 2787 2645 2788 2649
rect 2782 2644 2788 2645
rect 2942 2649 2948 2650
rect 2942 2645 2943 2649
rect 2947 2645 2948 2649
rect 2942 2644 2948 2645
rect 3094 2649 3100 2650
rect 3094 2645 3095 2649
rect 3099 2645 3100 2649
rect 3094 2644 3100 2645
rect 3238 2649 3244 2650
rect 3238 2645 3239 2649
rect 3243 2645 3244 2649
rect 3238 2644 3244 2645
rect 3382 2649 3388 2650
rect 3382 2645 3383 2649
rect 3387 2645 3388 2649
rect 3382 2644 3388 2645
rect 3534 2649 3540 2650
rect 3534 2645 3535 2649
rect 3539 2645 3540 2649
rect 3534 2644 3540 2645
rect 3942 2648 3948 2649
rect 3942 2644 3943 2648
rect 3947 2644 3948 2648
rect 2046 2643 2052 2644
rect 2006 2640 2012 2641
rect 166 2629 172 2630
rect 110 2628 116 2629
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 166 2625 167 2629
rect 171 2625 172 2629
rect 166 2624 172 2625
rect 358 2629 364 2630
rect 358 2625 359 2629
rect 363 2625 364 2629
rect 358 2624 364 2625
rect 558 2629 564 2630
rect 558 2625 559 2629
rect 563 2625 564 2629
rect 558 2624 564 2625
rect 758 2629 764 2630
rect 758 2625 759 2629
rect 763 2625 764 2629
rect 758 2624 764 2625
rect 950 2629 956 2630
rect 950 2625 951 2629
rect 955 2625 956 2629
rect 950 2624 956 2625
rect 1142 2629 1148 2630
rect 1142 2625 1143 2629
rect 1147 2625 1148 2629
rect 1142 2624 1148 2625
rect 1326 2629 1332 2630
rect 1326 2625 1327 2629
rect 1331 2625 1332 2629
rect 1326 2624 1332 2625
rect 1510 2629 1516 2630
rect 1510 2625 1511 2629
rect 1515 2625 1516 2629
rect 1510 2624 1516 2625
rect 1702 2629 1708 2630
rect 1702 2625 1703 2629
rect 1707 2625 1708 2629
rect 1702 2624 1708 2625
rect 2006 2628 2012 2629
rect 2006 2624 2007 2628
rect 2011 2624 2012 2628
rect 110 2623 116 2624
rect 112 2587 114 2623
rect 168 2587 170 2624
rect 360 2587 362 2624
rect 560 2587 562 2624
rect 760 2587 762 2624
rect 952 2587 954 2624
rect 1144 2587 1146 2624
rect 1328 2587 1330 2624
rect 1512 2587 1514 2624
rect 1704 2587 1706 2624
rect 2006 2623 2012 2624
rect 2008 2587 2010 2623
rect 2048 2615 2050 2643
rect 2096 2615 2098 2644
rect 2264 2615 2266 2644
rect 2440 2615 2442 2644
rect 2616 2615 2618 2644
rect 2784 2615 2786 2644
rect 2944 2615 2946 2644
rect 3096 2615 3098 2644
rect 3240 2615 3242 2644
rect 3384 2615 3386 2644
rect 3536 2615 3538 2644
rect 3942 2643 3948 2644
rect 3944 2615 3946 2643
rect 2047 2614 2051 2615
rect 2047 2609 2051 2610
rect 2095 2614 2099 2615
rect 2095 2609 2099 2610
rect 2215 2614 2219 2615
rect 2215 2609 2219 2610
rect 2263 2614 2267 2615
rect 2263 2609 2267 2610
rect 2367 2614 2371 2615
rect 2367 2609 2371 2610
rect 2439 2614 2443 2615
rect 2439 2609 2443 2610
rect 2519 2614 2523 2615
rect 2519 2609 2523 2610
rect 2615 2614 2619 2615
rect 2615 2609 2619 2610
rect 2671 2614 2675 2615
rect 2671 2609 2675 2610
rect 2783 2614 2787 2615
rect 2783 2609 2787 2610
rect 2815 2614 2819 2615
rect 2815 2609 2819 2610
rect 2943 2614 2947 2615
rect 2943 2609 2947 2610
rect 2951 2614 2955 2615
rect 2951 2609 2955 2610
rect 3087 2614 3091 2615
rect 3087 2609 3091 2610
rect 3095 2614 3099 2615
rect 3095 2609 3099 2610
rect 3223 2614 3227 2615
rect 3223 2609 3227 2610
rect 3239 2614 3243 2615
rect 3239 2609 3243 2610
rect 3367 2614 3371 2615
rect 3367 2609 3371 2610
rect 3383 2614 3387 2615
rect 3383 2609 3387 2610
rect 3535 2614 3539 2615
rect 3535 2609 3539 2610
rect 3943 2614 3947 2615
rect 3943 2609 3947 2610
rect 2048 2589 2050 2609
rect 2046 2588 2052 2589
rect 2216 2588 2218 2609
rect 2368 2588 2370 2609
rect 2520 2588 2522 2609
rect 2672 2588 2674 2609
rect 2816 2588 2818 2609
rect 2952 2588 2954 2609
rect 3088 2588 3090 2609
rect 3224 2588 3226 2609
rect 3368 2588 3370 2609
rect 3944 2589 3946 2609
rect 3942 2588 3948 2589
rect 111 2586 115 2587
rect 111 2581 115 2582
rect 167 2586 171 2587
rect 167 2581 171 2582
rect 359 2586 363 2587
rect 359 2581 363 2582
rect 559 2586 563 2587
rect 559 2581 563 2582
rect 575 2586 579 2587
rect 575 2581 579 2582
rect 687 2586 691 2587
rect 687 2581 691 2582
rect 759 2586 763 2587
rect 759 2581 763 2582
rect 807 2586 811 2587
rect 807 2581 811 2582
rect 935 2586 939 2587
rect 935 2581 939 2582
rect 951 2586 955 2587
rect 951 2581 955 2582
rect 1071 2586 1075 2587
rect 1071 2581 1075 2582
rect 1143 2586 1147 2587
rect 1143 2581 1147 2582
rect 1207 2586 1211 2587
rect 1207 2581 1211 2582
rect 1327 2586 1331 2587
rect 1327 2581 1331 2582
rect 1351 2586 1355 2587
rect 1351 2581 1355 2582
rect 1495 2586 1499 2587
rect 1495 2581 1499 2582
rect 1511 2586 1515 2587
rect 1511 2581 1515 2582
rect 1647 2586 1651 2587
rect 1647 2581 1651 2582
rect 1703 2586 1707 2587
rect 1703 2581 1707 2582
rect 1799 2586 1803 2587
rect 1799 2581 1803 2582
rect 2007 2586 2011 2587
rect 2046 2584 2047 2588
rect 2051 2584 2052 2588
rect 2046 2583 2052 2584
rect 2214 2587 2220 2588
rect 2214 2583 2215 2587
rect 2219 2583 2220 2587
rect 2214 2582 2220 2583
rect 2366 2587 2372 2588
rect 2366 2583 2367 2587
rect 2371 2583 2372 2587
rect 2366 2582 2372 2583
rect 2518 2587 2524 2588
rect 2518 2583 2519 2587
rect 2523 2583 2524 2587
rect 2518 2582 2524 2583
rect 2670 2587 2676 2588
rect 2670 2583 2671 2587
rect 2675 2583 2676 2587
rect 2670 2582 2676 2583
rect 2814 2587 2820 2588
rect 2814 2583 2815 2587
rect 2819 2583 2820 2587
rect 2814 2582 2820 2583
rect 2950 2587 2956 2588
rect 2950 2583 2951 2587
rect 2955 2583 2956 2587
rect 2950 2582 2956 2583
rect 3086 2587 3092 2588
rect 3086 2583 3087 2587
rect 3091 2583 3092 2587
rect 3086 2582 3092 2583
rect 3222 2587 3228 2588
rect 3222 2583 3223 2587
rect 3227 2583 3228 2587
rect 3222 2582 3228 2583
rect 3366 2587 3372 2588
rect 3366 2583 3367 2587
rect 3371 2583 3372 2587
rect 3942 2584 3943 2588
rect 3947 2584 3948 2588
rect 3942 2583 3948 2584
rect 3366 2582 3372 2583
rect 2007 2581 2011 2582
rect 112 2561 114 2581
rect 110 2560 116 2561
rect 576 2560 578 2581
rect 688 2560 690 2581
rect 808 2560 810 2581
rect 936 2560 938 2581
rect 1072 2560 1074 2581
rect 1208 2560 1210 2581
rect 1352 2560 1354 2581
rect 1496 2560 1498 2581
rect 1648 2560 1650 2581
rect 1800 2560 1802 2581
rect 2008 2561 2010 2581
rect 2046 2571 2052 2572
rect 2046 2567 2047 2571
rect 2051 2567 2052 2571
rect 3942 2571 3948 2572
rect 2046 2566 2052 2567
rect 2214 2568 2220 2569
rect 2006 2560 2012 2561
rect 110 2556 111 2560
rect 115 2556 116 2560
rect 110 2555 116 2556
rect 574 2559 580 2560
rect 574 2555 575 2559
rect 579 2555 580 2559
rect 574 2554 580 2555
rect 686 2559 692 2560
rect 686 2555 687 2559
rect 691 2555 692 2559
rect 686 2554 692 2555
rect 806 2559 812 2560
rect 806 2555 807 2559
rect 811 2555 812 2559
rect 806 2554 812 2555
rect 934 2559 940 2560
rect 934 2555 935 2559
rect 939 2555 940 2559
rect 934 2554 940 2555
rect 1070 2559 1076 2560
rect 1070 2555 1071 2559
rect 1075 2555 1076 2559
rect 1070 2554 1076 2555
rect 1206 2559 1212 2560
rect 1206 2555 1207 2559
rect 1211 2555 1212 2559
rect 1206 2554 1212 2555
rect 1350 2559 1356 2560
rect 1350 2555 1351 2559
rect 1355 2555 1356 2559
rect 1350 2554 1356 2555
rect 1494 2559 1500 2560
rect 1494 2555 1495 2559
rect 1499 2555 1500 2559
rect 1494 2554 1500 2555
rect 1646 2559 1652 2560
rect 1646 2555 1647 2559
rect 1651 2555 1652 2559
rect 1646 2554 1652 2555
rect 1798 2559 1804 2560
rect 1798 2555 1799 2559
rect 1803 2555 1804 2559
rect 2006 2556 2007 2560
rect 2011 2556 2012 2560
rect 2006 2555 2012 2556
rect 1798 2554 1804 2555
rect 110 2543 116 2544
rect 110 2539 111 2543
rect 115 2539 116 2543
rect 2006 2543 2012 2544
rect 110 2538 116 2539
rect 574 2540 580 2541
rect 112 2507 114 2538
rect 574 2536 575 2540
rect 579 2536 580 2540
rect 574 2535 580 2536
rect 686 2540 692 2541
rect 686 2536 687 2540
rect 691 2536 692 2540
rect 686 2535 692 2536
rect 806 2540 812 2541
rect 806 2536 807 2540
rect 811 2536 812 2540
rect 806 2535 812 2536
rect 934 2540 940 2541
rect 934 2536 935 2540
rect 939 2536 940 2540
rect 934 2535 940 2536
rect 1070 2540 1076 2541
rect 1070 2536 1071 2540
rect 1075 2536 1076 2540
rect 1070 2535 1076 2536
rect 1206 2540 1212 2541
rect 1206 2536 1207 2540
rect 1211 2536 1212 2540
rect 1206 2535 1212 2536
rect 1350 2540 1356 2541
rect 1350 2536 1351 2540
rect 1355 2536 1356 2540
rect 1350 2535 1356 2536
rect 1494 2540 1500 2541
rect 1494 2536 1495 2540
rect 1499 2536 1500 2540
rect 1494 2535 1500 2536
rect 1646 2540 1652 2541
rect 1646 2536 1647 2540
rect 1651 2536 1652 2540
rect 1646 2535 1652 2536
rect 1798 2540 1804 2541
rect 1798 2536 1799 2540
rect 1803 2536 1804 2540
rect 2006 2539 2007 2543
rect 2011 2539 2012 2543
rect 2006 2538 2012 2539
rect 1798 2535 1804 2536
rect 576 2507 578 2535
rect 688 2507 690 2535
rect 808 2507 810 2535
rect 936 2507 938 2535
rect 1072 2507 1074 2535
rect 1208 2507 1210 2535
rect 1352 2507 1354 2535
rect 1496 2507 1498 2535
rect 1648 2507 1650 2535
rect 1800 2507 1802 2535
rect 2008 2507 2010 2538
rect 2048 2535 2050 2566
rect 2214 2564 2215 2568
rect 2219 2564 2220 2568
rect 2214 2563 2220 2564
rect 2366 2568 2372 2569
rect 2366 2564 2367 2568
rect 2371 2564 2372 2568
rect 2366 2563 2372 2564
rect 2518 2568 2524 2569
rect 2518 2564 2519 2568
rect 2523 2564 2524 2568
rect 2518 2563 2524 2564
rect 2670 2568 2676 2569
rect 2670 2564 2671 2568
rect 2675 2564 2676 2568
rect 2670 2563 2676 2564
rect 2814 2568 2820 2569
rect 2814 2564 2815 2568
rect 2819 2564 2820 2568
rect 2814 2563 2820 2564
rect 2950 2568 2956 2569
rect 2950 2564 2951 2568
rect 2955 2564 2956 2568
rect 2950 2563 2956 2564
rect 3086 2568 3092 2569
rect 3086 2564 3087 2568
rect 3091 2564 3092 2568
rect 3086 2563 3092 2564
rect 3222 2568 3228 2569
rect 3222 2564 3223 2568
rect 3227 2564 3228 2568
rect 3222 2563 3228 2564
rect 3366 2568 3372 2569
rect 3366 2564 3367 2568
rect 3371 2564 3372 2568
rect 3942 2567 3943 2571
rect 3947 2567 3948 2571
rect 3942 2566 3948 2567
rect 3366 2563 3372 2564
rect 2216 2535 2218 2563
rect 2368 2535 2370 2563
rect 2520 2535 2522 2563
rect 2672 2535 2674 2563
rect 2816 2535 2818 2563
rect 2952 2535 2954 2563
rect 3088 2535 3090 2563
rect 3224 2535 3226 2563
rect 3368 2535 3370 2563
rect 3944 2535 3946 2566
rect 2047 2534 2051 2535
rect 2047 2529 2051 2530
rect 2095 2534 2099 2535
rect 2095 2529 2099 2530
rect 2215 2534 2219 2535
rect 2215 2529 2219 2530
rect 2343 2534 2347 2535
rect 2343 2529 2347 2530
rect 2367 2534 2371 2535
rect 2367 2529 2371 2530
rect 2471 2534 2475 2535
rect 2471 2529 2475 2530
rect 2519 2534 2523 2535
rect 2519 2529 2523 2530
rect 2599 2534 2603 2535
rect 2599 2529 2603 2530
rect 2671 2534 2675 2535
rect 2671 2529 2675 2530
rect 2719 2534 2723 2535
rect 2719 2529 2723 2530
rect 2815 2534 2819 2535
rect 2815 2529 2819 2530
rect 2839 2534 2843 2535
rect 2839 2529 2843 2530
rect 2951 2534 2955 2535
rect 2951 2529 2955 2530
rect 2967 2534 2971 2535
rect 2967 2529 2971 2530
rect 3087 2534 3091 2535
rect 3087 2529 3091 2530
rect 3095 2534 3099 2535
rect 3095 2529 3099 2530
rect 3223 2534 3227 2535
rect 3223 2529 3227 2530
rect 3367 2534 3371 2535
rect 3367 2529 3371 2530
rect 3943 2534 3947 2535
rect 3943 2529 3947 2530
rect 111 2506 115 2507
rect 111 2501 115 2502
rect 503 2506 507 2507
rect 503 2501 507 2502
rect 575 2506 579 2507
rect 575 2501 579 2502
rect 607 2506 611 2507
rect 607 2501 611 2502
rect 687 2506 691 2507
rect 687 2501 691 2502
rect 719 2506 723 2507
rect 719 2501 723 2502
rect 807 2506 811 2507
rect 807 2501 811 2502
rect 847 2506 851 2507
rect 847 2501 851 2502
rect 935 2506 939 2507
rect 935 2501 939 2502
rect 983 2506 987 2507
rect 983 2501 987 2502
rect 1071 2506 1075 2507
rect 1071 2501 1075 2502
rect 1127 2506 1131 2507
rect 1127 2501 1131 2502
rect 1207 2506 1211 2507
rect 1207 2501 1211 2502
rect 1279 2506 1283 2507
rect 1279 2501 1283 2502
rect 1351 2506 1355 2507
rect 1351 2501 1355 2502
rect 1431 2506 1435 2507
rect 1431 2501 1435 2502
rect 1495 2506 1499 2507
rect 1495 2501 1499 2502
rect 1583 2506 1587 2507
rect 1583 2501 1587 2502
rect 1647 2506 1651 2507
rect 1647 2501 1651 2502
rect 1743 2506 1747 2507
rect 1743 2501 1747 2502
rect 1799 2506 1803 2507
rect 1799 2501 1803 2502
rect 1903 2506 1907 2507
rect 1903 2501 1907 2502
rect 2007 2506 2011 2507
rect 2048 2502 2050 2529
rect 2096 2505 2098 2529
rect 2216 2505 2218 2529
rect 2344 2505 2346 2529
rect 2472 2505 2474 2529
rect 2600 2505 2602 2529
rect 2720 2505 2722 2529
rect 2840 2505 2842 2529
rect 2968 2505 2970 2529
rect 3096 2505 3098 2529
rect 3224 2505 3226 2529
rect 2094 2504 2100 2505
rect 2007 2501 2011 2502
rect 2046 2501 2052 2502
rect 112 2474 114 2501
rect 504 2477 506 2501
rect 608 2477 610 2501
rect 720 2477 722 2501
rect 848 2477 850 2501
rect 984 2477 986 2501
rect 1128 2477 1130 2501
rect 1280 2477 1282 2501
rect 1432 2477 1434 2501
rect 1584 2477 1586 2501
rect 1744 2477 1746 2501
rect 1904 2477 1906 2501
rect 502 2476 508 2477
rect 110 2473 116 2474
rect 110 2469 111 2473
rect 115 2469 116 2473
rect 502 2472 503 2476
rect 507 2472 508 2476
rect 502 2471 508 2472
rect 606 2476 612 2477
rect 606 2472 607 2476
rect 611 2472 612 2476
rect 606 2471 612 2472
rect 718 2476 724 2477
rect 718 2472 719 2476
rect 723 2472 724 2476
rect 718 2471 724 2472
rect 846 2476 852 2477
rect 846 2472 847 2476
rect 851 2472 852 2476
rect 846 2471 852 2472
rect 982 2476 988 2477
rect 982 2472 983 2476
rect 987 2472 988 2476
rect 982 2471 988 2472
rect 1126 2476 1132 2477
rect 1126 2472 1127 2476
rect 1131 2472 1132 2476
rect 1126 2471 1132 2472
rect 1278 2476 1284 2477
rect 1278 2472 1279 2476
rect 1283 2472 1284 2476
rect 1278 2471 1284 2472
rect 1430 2476 1436 2477
rect 1430 2472 1431 2476
rect 1435 2472 1436 2476
rect 1430 2471 1436 2472
rect 1582 2476 1588 2477
rect 1582 2472 1583 2476
rect 1587 2472 1588 2476
rect 1582 2471 1588 2472
rect 1742 2476 1748 2477
rect 1742 2472 1743 2476
rect 1747 2472 1748 2476
rect 1742 2471 1748 2472
rect 1902 2476 1908 2477
rect 1902 2472 1903 2476
rect 1907 2472 1908 2476
rect 2008 2474 2010 2501
rect 2046 2497 2047 2501
rect 2051 2497 2052 2501
rect 2094 2500 2095 2504
rect 2099 2500 2100 2504
rect 2094 2499 2100 2500
rect 2214 2504 2220 2505
rect 2214 2500 2215 2504
rect 2219 2500 2220 2504
rect 2214 2499 2220 2500
rect 2342 2504 2348 2505
rect 2342 2500 2343 2504
rect 2347 2500 2348 2504
rect 2342 2499 2348 2500
rect 2470 2504 2476 2505
rect 2470 2500 2471 2504
rect 2475 2500 2476 2504
rect 2470 2499 2476 2500
rect 2598 2504 2604 2505
rect 2598 2500 2599 2504
rect 2603 2500 2604 2504
rect 2598 2499 2604 2500
rect 2718 2504 2724 2505
rect 2718 2500 2719 2504
rect 2723 2500 2724 2504
rect 2718 2499 2724 2500
rect 2838 2504 2844 2505
rect 2838 2500 2839 2504
rect 2843 2500 2844 2504
rect 2838 2499 2844 2500
rect 2966 2504 2972 2505
rect 2966 2500 2967 2504
rect 2971 2500 2972 2504
rect 2966 2499 2972 2500
rect 3094 2504 3100 2505
rect 3094 2500 3095 2504
rect 3099 2500 3100 2504
rect 3094 2499 3100 2500
rect 3222 2504 3228 2505
rect 3222 2500 3223 2504
rect 3227 2500 3228 2504
rect 3944 2502 3946 2529
rect 3222 2499 3228 2500
rect 3942 2501 3948 2502
rect 2046 2496 2052 2497
rect 3942 2497 3943 2501
rect 3947 2497 3948 2501
rect 3942 2496 3948 2497
rect 2094 2485 2100 2486
rect 2046 2484 2052 2485
rect 2046 2480 2047 2484
rect 2051 2480 2052 2484
rect 2094 2481 2095 2485
rect 2099 2481 2100 2485
rect 2094 2480 2100 2481
rect 2214 2485 2220 2486
rect 2214 2481 2215 2485
rect 2219 2481 2220 2485
rect 2214 2480 2220 2481
rect 2342 2485 2348 2486
rect 2342 2481 2343 2485
rect 2347 2481 2348 2485
rect 2342 2480 2348 2481
rect 2470 2485 2476 2486
rect 2470 2481 2471 2485
rect 2475 2481 2476 2485
rect 2470 2480 2476 2481
rect 2598 2485 2604 2486
rect 2598 2481 2599 2485
rect 2603 2481 2604 2485
rect 2598 2480 2604 2481
rect 2718 2485 2724 2486
rect 2718 2481 2719 2485
rect 2723 2481 2724 2485
rect 2718 2480 2724 2481
rect 2838 2485 2844 2486
rect 2838 2481 2839 2485
rect 2843 2481 2844 2485
rect 2838 2480 2844 2481
rect 2966 2485 2972 2486
rect 2966 2481 2967 2485
rect 2971 2481 2972 2485
rect 2966 2480 2972 2481
rect 3094 2485 3100 2486
rect 3094 2481 3095 2485
rect 3099 2481 3100 2485
rect 3094 2480 3100 2481
rect 3222 2485 3228 2486
rect 3222 2481 3223 2485
rect 3227 2481 3228 2485
rect 3222 2480 3228 2481
rect 3942 2484 3948 2485
rect 3942 2480 3943 2484
rect 3947 2480 3948 2484
rect 2046 2479 2052 2480
rect 1902 2471 1908 2472
rect 2006 2473 2012 2474
rect 110 2468 116 2469
rect 2006 2469 2007 2473
rect 2011 2469 2012 2473
rect 2006 2468 2012 2469
rect 502 2457 508 2458
rect 110 2456 116 2457
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 502 2453 503 2457
rect 507 2453 508 2457
rect 502 2452 508 2453
rect 606 2457 612 2458
rect 606 2453 607 2457
rect 611 2453 612 2457
rect 606 2452 612 2453
rect 718 2457 724 2458
rect 718 2453 719 2457
rect 723 2453 724 2457
rect 718 2452 724 2453
rect 846 2457 852 2458
rect 846 2453 847 2457
rect 851 2453 852 2457
rect 846 2452 852 2453
rect 982 2457 988 2458
rect 982 2453 983 2457
rect 987 2453 988 2457
rect 982 2452 988 2453
rect 1126 2457 1132 2458
rect 1126 2453 1127 2457
rect 1131 2453 1132 2457
rect 1126 2452 1132 2453
rect 1278 2457 1284 2458
rect 1278 2453 1279 2457
rect 1283 2453 1284 2457
rect 1278 2452 1284 2453
rect 1430 2457 1436 2458
rect 1430 2453 1431 2457
rect 1435 2453 1436 2457
rect 1430 2452 1436 2453
rect 1582 2457 1588 2458
rect 1582 2453 1583 2457
rect 1587 2453 1588 2457
rect 1582 2452 1588 2453
rect 1742 2457 1748 2458
rect 1742 2453 1743 2457
rect 1747 2453 1748 2457
rect 1742 2452 1748 2453
rect 1902 2457 1908 2458
rect 1902 2453 1903 2457
rect 1907 2453 1908 2457
rect 1902 2452 1908 2453
rect 2006 2456 2012 2457
rect 2006 2452 2007 2456
rect 2011 2452 2012 2456
rect 110 2451 116 2452
rect 112 2415 114 2451
rect 504 2415 506 2452
rect 608 2415 610 2452
rect 720 2415 722 2452
rect 848 2415 850 2452
rect 984 2415 986 2452
rect 1128 2415 1130 2452
rect 1280 2415 1282 2452
rect 1432 2415 1434 2452
rect 1584 2415 1586 2452
rect 1744 2415 1746 2452
rect 1904 2415 1906 2452
rect 2006 2451 2012 2452
rect 2008 2415 2010 2451
rect 2048 2447 2050 2479
rect 2096 2447 2098 2480
rect 2216 2447 2218 2480
rect 2344 2447 2346 2480
rect 2472 2447 2474 2480
rect 2600 2447 2602 2480
rect 2720 2447 2722 2480
rect 2840 2447 2842 2480
rect 2968 2447 2970 2480
rect 3096 2447 3098 2480
rect 3224 2447 3226 2480
rect 3942 2479 3948 2480
rect 3944 2447 3946 2479
rect 2047 2446 2051 2447
rect 2047 2441 2051 2442
rect 2071 2446 2075 2447
rect 2071 2441 2075 2442
rect 2095 2446 2099 2447
rect 2095 2441 2099 2442
rect 2191 2446 2195 2447
rect 2191 2441 2195 2442
rect 2215 2446 2219 2447
rect 2215 2441 2219 2442
rect 2319 2446 2323 2447
rect 2319 2441 2323 2442
rect 2343 2446 2347 2447
rect 2343 2441 2347 2442
rect 2439 2446 2443 2447
rect 2439 2441 2443 2442
rect 2471 2446 2475 2447
rect 2471 2441 2475 2442
rect 2559 2446 2563 2447
rect 2559 2441 2563 2442
rect 2599 2446 2603 2447
rect 2599 2441 2603 2442
rect 2679 2446 2683 2447
rect 2679 2441 2683 2442
rect 2719 2446 2723 2447
rect 2719 2441 2723 2442
rect 2791 2446 2795 2447
rect 2791 2441 2795 2442
rect 2839 2446 2843 2447
rect 2839 2441 2843 2442
rect 2911 2446 2915 2447
rect 2911 2441 2915 2442
rect 2967 2446 2971 2447
rect 2967 2441 2971 2442
rect 3031 2446 3035 2447
rect 3031 2441 3035 2442
rect 3095 2446 3099 2447
rect 3095 2441 3099 2442
rect 3151 2446 3155 2447
rect 3151 2441 3155 2442
rect 3223 2446 3227 2447
rect 3223 2441 3227 2442
rect 3943 2446 3947 2447
rect 3943 2441 3947 2442
rect 2048 2421 2050 2441
rect 2046 2420 2052 2421
rect 2072 2420 2074 2441
rect 2192 2420 2194 2441
rect 2320 2420 2322 2441
rect 2440 2420 2442 2441
rect 2560 2420 2562 2441
rect 2680 2420 2682 2441
rect 2792 2420 2794 2441
rect 2912 2420 2914 2441
rect 3032 2420 3034 2441
rect 3152 2420 3154 2441
rect 3944 2421 3946 2441
rect 3942 2420 3948 2421
rect 2046 2416 2047 2420
rect 2051 2416 2052 2420
rect 2046 2415 2052 2416
rect 2070 2419 2076 2420
rect 2070 2415 2071 2419
rect 2075 2415 2076 2419
rect 111 2414 115 2415
rect 111 2409 115 2410
rect 503 2414 507 2415
rect 503 2409 507 2410
rect 535 2414 539 2415
rect 535 2409 539 2410
rect 607 2414 611 2415
rect 607 2409 611 2410
rect 671 2414 675 2415
rect 671 2409 675 2410
rect 719 2414 723 2415
rect 719 2409 723 2410
rect 815 2414 819 2415
rect 815 2409 819 2410
rect 847 2414 851 2415
rect 847 2409 851 2410
rect 959 2414 963 2415
rect 959 2409 963 2410
rect 983 2414 987 2415
rect 983 2409 987 2410
rect 1103 2414 1107 2415
rect 1103 2409 1107 2410
rect 1127 2414 1131 2415
rect 1127 2409 1131 2410
rect 1247 2414 1251 2415
rect 1247 2409 1251 2410
rect 1279 2414 1283 2415
rect 1279 2409 1283 2410
rect 1391 2414 1395 2415
rect 1391 2409 1395 2410
rect 1431 2414 1435 2415
rect 1431 2409 1435 2410
rect 1527 2414 1531 2415
rect 1527 2409 1531 2410
rect 1583 2414 1587 2415
rect 1583 2409 1587 2410
rect 1655 2414 1659 2415
rect 1655 2409 1659 2410
rect 1743 2414 1747 2415
rect 1743 2409 1747 2410
rect 1791 2414 1795 2415
rect 1791 2409 1795 2410
rect 1903 2414 1907 2415
rect 1903 2409 1907 2410
rect 2007 2414 2011 2415
rect 2070 2414 2076 2415
rect 2190 2419 2196 2420
rect 2190 2415 2191 2419
rect 2195 2415 2196 2419
rect 2190 2414 2196 2415
rect 2318 2419 2324 2420
rect 2318 2415 2319 2419
rect 2323 2415 2324 2419
rect 2318 2414 2324 2415
rect 2438 2419 2444 2420
rect 2438 2415 2439 2419
rect 2443 2415 2444 2419
rect 2438 2414 2444 2415
rect 2558 2419 2564 2420
rect 2558 2415 2559 2419
rect 2563 2415 2564 2419
rect 2558 2414 2564 2415
rect 2678 2419 2684 2420
rect 2678 2415 2679 2419
rect 2683 2415 2684 2419
rect 2678 2414 2684 2415
rect 2790 2419 2796 2420
rect 2790 2415 2791 2419
rect 2795 2415 2796 2419
rect 2790 2414 2796 2415
rect 2910 2419 2916 2420
rect 2910 2415 2911 2419
rect 2915 2415 2916 2419
rect 2910 2414 2916 2415
rect 3030 2419 3036 2420
rect 3030 2415 3031 2419
rect 3035 2415 3036 2419
rect 3030 2414 3036 2415
rect 3150 2419 3156 2420
rect 3150 2415 3151 2419
rect 3155 2415 3156 2419
rect 3942 2416 3943 2420
rect 3947 2416 3948 2420
rect 3942 2415 3948 2416
rect 3150 2414 3156 2415
rect 2007 2409 2011 2410
rect 112 2389 114 2409
rect 110 2388 116 2389
rect 536 2388 538 2409
rect 672 2388 674 2409
rect 816 2388 818 2409
rect 960 2388 962 2409
rect 1104 2388 1106 2409
rect 1248 2388 1250 2409
rect 1392 2388 1394 2409
rect 1528 2388 1530 2409
rect 1656 2388 1658 2409
rect 1792 2388 1794 2409
rect 1904 2388 1906 2409
rect 2008 2389 2010 2409
rect 2046 2403 2052 2404
rect 2046 2399 2047 2403
rect 2051 2399 2052 2403
rect 3942 2403 3948 2404
rect 2046 2398 2052 2399
rect 2070 2400 2076 2401
rect 2006 2388 2012 2389
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 110 2383 116 2384
rect 534 2387 540 2388
rect 534 2383 535 2387
rect 539 2383 540 2387
rect 534 2382 540 2383
rect 670 2387 676 2388
rect 670 2383 671 2387
rect 675 2383 676 2387
rect 670 2382 676 2383
rect 814 2387 820 2388
rect 814 2383 815 2387
rect 819 2383 820 2387
rect 814 2382 820 2383
rect 958 2387 964 2388
rect 958 2383 959 2387
rect 963 2383 964 2387
rect 958 2382 964 2383
rect 1102 2387 1108 2388
rect 1102 2383 1103 2387
rect 1107 2383 1108 2387
rect 1102 2382 1108 2383
rect 1246 2387 1252 2388
rect 1246 2383 1247 2387
rect 1251 2383 1252 2387
rect 1246 2382 1252 2383
rect 1390 2387 1396 2388
rect 1390 2383 1391 2387
rect 1395 2383 1396 2387
rect 1390 2382 1396 2383
rect 1526 2387 1532 2388
rect 1526 2383 1527 2387
rect 1531 2383 1532 2387
rect 1526 2382 1532 2383
rect 1654 2387 1660 2388
rect 1654 2383 1655 2387
rect 1659 2383 1660 2387
rect 1654 2382 1660 2383
rect 1790 2387 1796 2388
rect 1790 2383 1791 2387
rect 1795 2383 1796 2387
rect 1790 2382 1796 2383
rect 1902 2387 1908 2388
rect 1902 2383 1903 2387
rect 1907 2383 1908 2387
rect 2006 2384 2007 2388
rect 2011 2384 2012 2388
rect 2006 2383 2012 2384
rect 1902 2382 1908 2383
rect 110 2371 116 2372
rect 110 2367 111 2371
rect 115 2367 116 2371
rect 2006 2371 2012 2372
rect 110 2366 116 2367
rect 534 2368 540 2369
rect 112 2335 114 2366
rect 534 2364 535 2368
rect 539 2364 540 2368
rect 534 2363 540 2364
rect 670 2368 676 2369
rect 670 2364 671 2368
rect 675 2364 676 2368
rect 670 2363 676 2364
rect 814 2368 820 2369
rect 814 2364 815 2368
rect 819 2364 820 2368
rect 814 2363 820 2364
rect 958 2368 964 2369
rect 958 2364 959 2368
rect 963 2364 964 2368
rect 958 2363 964 2364
rect 1102 2368 1108 2369
rect 1102 2364 1103 2368
rect 1107 2364 1108 2368
rect 1102 2363 1108 2364
rect 1246 2368 1252 2369
rect 1246 2364 1247 2368
rect 1251 2364 1252 2368
rect 1246 2363 1252 2364
rect 1390 2368 1396 2369
rect 1390 2364 1391 2368
rect 1395 2364 1396 2368
rect 1390 2363 1396 2364
rect 1526 2368 1532 2369
rect 1526 2364 1527 2368
rect 1531 2364 1532 2368
rect 1526 2363 1532 2364
rect 1654 2368 1660 2369
rect 1654 2364 1655 2368
rect 1659 2364 1660 2368
rect 1654 2363 1660 2364
rect 1790 2368 1796 2369
rect 1790 2364 1791 2368
rect 1795 2364 1796 2368
rect 1790 2363 1796 2364
rect 1902 2368 1908 2369
rect 1902 2364 1903 2368
rect 1907 2364 1908 2368
rect 2006 2367 2007 2371
rect 2011 2367 2012 2371
rect 2048 2367 2050 2398
rect 2070 2396 2071 2400
rect 2075 2396 2076 2400
rect 2070 2395 2076 2396
rect 2190 2400 2196 2401
rect 2190 2396 2191 2400
rect 2195 2396 2196 2400
rect 2190 2395 2196 2396
rect 2318 2400 2324 2401
rect 2318 2396 2319 2400
rect 2323 2396 2324 2400
rect 2318 2395 2324 2396
rect 2438 2400 2444 2401
rect 2438 2396 2439 2400
rect 2443 2396 2444 2400
rect 2438 2395 2444 2396
rect 2558 2400 2564 2401
rect 2558 2396 2559 2400
rect 2563 2396 2564 2400
rect 2558 2395 2564 2396
rect 2678 2400 2684 2401
rect 2678 2396 2679 2400
rect 2683 2396 2684 2400
rect 2678 2395 2684 2396
rect 2790 2400 2796 2401
rect 2790 2396 2791 2400
rect 2795 2396 2796 2400
rect 2790 2395 2796 2396
rect 2910 2400 2916 2401
rect 2910 2396 2911 2400
rect 2915 2396 2916 2400
rect 2910 2395 2916 2396
rect 3030 2400 3036 2401
rect 3030 2396 3031 2400
rect 3035 2396 3036 2400
rect 3030 2395 3036 2396
rect 3150 2400 3156 2401
rect 3150 2396 3151 2400
rect 3155 2396 3156 2400
rect 3942 2399 3943 2403
rect 3947 2399 3948 2403
rect 3942 2398 3948 2399
rect 3150 2395 3156 2396
rect 2072 2367 2074 2395
rect 2192 2367 2194 2395
rect 2320 2367 2322 2395
rect 2440 2367 2442 2395
rect 2560 2367 2562 2395
rect 2680 2367 2682 2395
rect 2792 2367 2794 2395
rect 2912 2367 2914 2395
rect 3032 2367 3034 2395
rect 3152 2367 3154 2395
rect 3944 2367 3946 2398
rect 2006 2366 2012 2367
rect 2047 2366 2051 2367
rect 1902 2363 1908 2364
rect 536 2335 538 2363
rect 672 2335 674 2363
rect 816 2335 818 2363
rect 960 2335 962 2363
rect 1104 2335 1106 2363
rect 1248 2335 1250 2363
rect 1392 2335 1394 2363
rect 1528 2335 1530 2363
rect 1656 2335 1658 2363
rect 1792 2335 1794 2363
rect 1904 2335 1906 2363
rect 2008 2335 2010 2366
rect 2047 2361 2051 2362
rect 2071 2366 2075 2367
rect 2071 2361 2075 2362
rect 2167 2366 2171 2367
rect 2167 2361 2171 2362
rect 2191 2366 2195 2367
rect 2191 2361 2195 2362
rect 2319 2366 2323 2367
rect 2319 2361 2323 2362
rect 2359 2366 2363 2367
rect 2359 2361 2363 2362
rect 2439 2366 2443 2367
rect 2439 2361 2443 2362
rect 2535 2366 2539 2367
rect 2535 2361 2539 2362
rect 2559 2366 2563 2367
rect 2559 2361 2563 2362
rect 2679 2366 2683 2367
rect 2679 2361 2683 2362
rect 2703 2366 2707 2367
rect 2703 2361 2707 2362
rect 2791 2366 2795 2367
rect 2791 2361 2795 2362
rect 2871 2366 2875 2367
rect 2871 2361 2875 2362
rect 2911 2366 2915 2367
rect 2911 2361 2915 2362
rect 3031 2366 3035 2367
rect 3031 2361 3035 2362
rect 3151 2366 3155 2367
rect 3151 2361 3155 2362
rect 3199 2366 3203 2367
rect 3199 2361 3203 2362
rect 3943 2366 3947 2367
rect 3943 2361 3947 2362
rect 111 2334 115 2335
rect 111 2329 115 2330
rect 535 2334 539 2335
rect 535 2329 539 2330
rect 647 2334 651 2335
rect 647 2329 651 2330
rect 671 2334 675 2335
rect 671 2329 675 2330
rect 767 2334 771 2335
rect 767 2329 771 2330
rect 815 2334 819 2335
rect 815 2329 819 2330
rect 895 2334 899 2335
rect 895 2329 899 2330
rect 959 2334 963 2335
rect 959 2329 963 2330
rect 1031 2334 1035 2335
rect 1031 2329 1035 2330
rect 1103 2334 1107 2335
rect 1103 2329 1107 2330
rect 1167 2334 1171 2335
rect 1167 2329 1171 2330
rect 1247 2334 1251 2335
rect 1247 2329 1251 2330
rect 1295 2334 1299 2335
rect 1295 2329 1299 2330
rect 1391 2334 1395 2335
rect 1391 2329 1395 2330
rect 1423 2334 1427 2335
rect 1423 2329 1427 2330
rect 1527 2334 1531 2335
rect 1527 2329 1531 2330
rect 1551 2334 1555 2335
rect 1551 2329 1555 2330
rect 1655 2334 1659 2335
rect 1655 2329 1659 2330
rect 1671 2334 1675 2335
rect 1671 2329 1675 2330
rect 1791 2334 1795 2335
rect 1791 2329 1795 2330
rect 1799 2334 1803 2335
rect 1799 2329 1803 2330
rect 1903 2334 1907 2335
rect 1903 2329 1907 2330
rect 2007 2334 2011 2335
rect 2048 2334 2050 2361
rect 2168 2337 2170 2361
rect 2360 2337 2362 2361
rect 2536 2337 2538 2361
rect 2704 2337 2706 2361
rect 2872 2337 2874 2361
rect 3032 2337 3034 2361
rect 3200 2337 3202 2361
rect 2166 2336 2172 2337
rect 2007 2329 2011 2330
rect 2046 2333 2052 2334
rect 2046 2329 2047 2333
rect 2051 2329 2052 2333
rect 2166 2332 2167 2336
rect 2171 2332 2172 2336
rect 2166 2331 2172 2332
rect 2358 2336 2364 2337
rect 2358 2332 2359 2336
rect 2363 2332 2364 2336
rect 2358 2331 2364 2332
rect 2534 2336 2540 2337
rect 2534 2332 2535 2336
rect 2539 2332 2540 2336
rect 2534 2331 2540 2332
rect 2702 2336 2708 2337
rect 2702 2332 2703 2336
rect 2707 2332 2708 2336
rect 2702 2331 2708 2332
rect 2870 2336 2876 2337
rect 2870 2332 2871 2336
rect 2875 2332 2876 2336
rect 2870 2331 2876 2332
rect 3030 2336 3036 2337
rect 3030 2332 3031 2336
rect 3035 2332 3036 2336
rect 3030 2331 3036 2332
rect 3198 2336 3204 2337
rect 3198 2332 3199 2336
rect 3203 2332 3204 2336
rect 3944 2334 3946 2361
rect 3198 2331 3204 2332
rect 3942 2333 3948 2334
rect 112 2302 114 2329
rect 536 2305 538 2329
rect 648 2305 650 2329
rect 768 2305 770 2329
rect 896 2305 898 2329
rect 1032 2305 1034 2329
rect 1168 2305 1170 2329
rect 1296 2305 1298 2329
rect 1424 2305 1426 2329
rect 1552 2305 1554 2329
rect 1672 2305 1674 2329
rect 1800 2305 1802 2329
rect 1904 2305 1906 2329
rect 534 2304 540 2305
rect 110 2301 116 2302
rect 110 2297 111 2301
rect 115 2297 116 2301
rect 534 2300 535 2304
rect 539 2300 540 2304
rect 534 2299 540 2300
rect 646 2304 652 2305
rect 646 2300 647 2304
rect 651 2300 652 2304
rect 646 2299 652 2300
rect 766 2304 772 2305
rect 766 2300 767 2304
rect 771 2300 772 2304
rect 766 2299 772 2300
rect 894 2304 900 2305
rect 894 2300 895 2304
rect 899 2300 900 2304
rect 894 2299 900 2300
rect 1030 2304 1036 2305
rect 1030 2300 1031 2304
rect 1035 2300 1036 2304
rect 1030 2299 1036 2300
rect 1166 2304 1172 2305
rect 1166 2300 1167 2304
rect 1171 2300 1172 2304
rect 1166 2299 1172 2300
rect 1294 2304 1300 2305
rect 1294 2300 1295 2304
rect 1299 2300 1300 2304
rect 1294 2299 1300 2300
rect 1422 2304 1428 2305
rect 1422 2300 1423 2304
rect 1427 2300 1428 2304
rect 1422 2299 1428 2300
rect 1550 2304 1556 2305
rect 1550 2300 1551 2304
rect 1555 2300 1556 2304
rect 1550 2299 1556 2300
rect 1670 2304 1676 2305
rect 1670 2300 1671 2304
rect 1675 2300 1676 2304
rect 1670 2299 1676 2300
rect 1798 2304 1804 2305
rect 1798 2300 1799 2304
rect 1803 2300 1804 2304
rect 1798 2299 1804 2300
rect 1902 2304 1908 2305
rect 1902 2300 1903 2304
rect 1907 2300 1908 2304
rect 2008 2302 2010 2329
rect 2046 2328 2052 2329
rect 3942 2329 3943 2333
rect 3947 2329 3948 2333
rect 3942 2328 3948 2329
rect 2166 2317 2172 2318
rect 2046 2316 2052 2317
rect 2046 2312 2047 2316
rect 2051 2312 2052 2316
rect 2166 2313 2167 2317
rect 2171 2313 2172 2317
rect 2166 2312 2172 2313
rect 2358 2317 2364 2318
rect 2358 2313 2359 2317
rect 2363 2313 2364 2317
rect 2358 2312 2364 2313
rect 2534 2317 2540 2318
rect 2534 2313 2535 2317
rect 2539 2313 2540 2317
rect 2534 2312 2540 2313
rect 2702 2317 2708 2318
rect 2702 2313 2703 2317
rect 2707 2313 2708 2317
rect 2702 2312 2708 2313
rect 2870 2317 2876 2318
rect 2870 2313 2871 2317
rect 2875 2313 2876 2317
rect 2870 2312 2876 2313
rect 3030 2317 3036 2318
rect 3030 2313 3031 2317
rect 3035 2313 3036 2317
rect 3030 2312 3036 2313
rect 3198 2317 3204 2318
rect 3198 2313 3199 2317
rect 3203 2313 3204 2317
rect 3198 2312 3204 2313
rect 3942 2316 3948 2317
rect 3942 2312 3943 2316
rect 3947 2312 3948 2316
rect 2046 2311 2052 2312
rect 1902 2299 1908 2300
rect 2006 2301 2012 2302
rect 110 2296 116 2297
rect 2006 2297 2007 2301
rect 2011 2297 2012 2301
rect 2006 2296 2012 2297
rect 2048 2291 2050 2311
rect 2168 2291 2170 2312
rect 2360 2291 2362 2312
rect 2536 2291 2538 2312
rect 2704 2291 2706 2312
rect 2872 2291 2874 2312
rect 3032 2291 3034 2312
rect 3200 2291 3202 2312
rect 3942 2311 3948 2312
rect 3944 2291 3946 2311
rect 2047 2290 2051 2291
rect 534 2285 540 2286
rect 110 2284 116 2285
rect 110 2280 111 2284
rect 115 2280 116 2284
rect 534 2281 535 2285
rect 539 2281 540 2285
rect 534 2280 540 2281
rect 646 2285 652 2286
rect 646 2281 647 2285
rect 651 2281 652 2285
rect 646 2280 652 2281
rect 766 2285 772 2286
rect 766 2281 767 2285
rect 771 2281 772 2285
rect 766 2280 772 2281
rect 894 2285 900 2286
rect 894 2281 895 2285
rect 899 2281 900 2285
rect 894 2280 900 2281
rect 1030 2285 1036 2286
rect 1030 2281 1031 2285
rect 1035 2281 1036 2285
rect 1030 2280 1036 2281
rect 1166 2285 1172 2286
rect 1166 2281 1167 2285
rect 1171 2281 1172 2285
rect 1166 2280 1172 2281
rect 1294 2285 1300 2286
rect 1294 2281 1295 2285
rect 1299 2281 1300 2285
rect 1294 2280 1300 2281
rect 1422 2285 1428 2286
rect 1422 2281 1423 2285
rect 1427 2281 1428 2285
rect 1422 2280 1428 2281
rect 1550 2285 1556 2286
rect 1550 2281 1551 2285
rect 1555 2281 1556 2285
rect 1550 2280 1556 2281
rect 1670 2285 1676 2286
rect 1670 2281 1671 2285
rect 1675 2281 1676 2285
rect 1670 2280 1676 2281
rect 1798 2285 1804 2286
rect 1798 2281 1799 2285
rect 1803 2281 1804 2285
rect 1798 2280 1804 2281
rect 1902 2285 1908 2286
rect 2047 2285 2051 2286
rect 2071 2290 2075 2291
rect 2071 2285 2075 2286
rect 2167 2290 2171 2291
rect 2167 2285 2171 2286
rect 2287 2290 2291 2291
rect 2287 2285 2291 2286
rect 2359 2290 2363 2291
rect 2359 2285 2363 2286
rect 2423 2290 2427 2291
rect 2423 2285 2427 2286
rect 2535 2290 2539 2291
rect 2535 2285 2539 2286
rect 2559 2290 2563 2291
rect 2559 2285 2563 2286
rect 2703 2290 2707 2291
rect 2703 2285 2707 2286
rect 2839 2290 2843 2291
rect 2839 2285 2843 2286
rect 2871 2290 2875 2291
rect 2871 2285 2875 2286
rect 2983 2290 2987 2291
rect 2983 2285 2987 2286
rect 3031 2290 3035 2291
rect 3031 2285 3035 2286
rect 3127 2290 3131 2291
rect 3127 2285 3131 2286
rect 3199 2290 3203 2291
rect 3199 2285 3203 2286
rect 3271 2290 3275 2291
rect 3271 2285 3275 2286
rect 3943 2290 3947 2291
rect 3943 2285 3947 2286
rect 1902 2281 1903 2285
rect 1907 2281 1908 2285
rect 1902 2280 1908 2281
rect 2006 2284 2012 2285
rect 2006 2280 2007 2284
rect 2011 2280 2012 2284
rect 110 2279 116 2280
rect 112 2255 114 2279
rect 536 2255 538 2280
rect 648 2255 650 2280
rect 768 2255 770 2280
rect 896 2255 898 2280
rect 1032 2255 1034 2280
rect 1168 2255 1170 2280
rect 1296 2255 1298 2280
rect 1424 2255 1426 2280
rect 1552 2255 1554 2280
rect 1672 2255 1674 2280
rect 1800 2255 1802 2280
rect 1904 2255 1906 2280
rect 2006 2279 2012 2280
rect 2008 2255 2010 2279
rect 2048 2265 2050 2285
rect 2046 2264 2052 2265
rect 2072 2264 2074 2285
rect 2168 2264 2170 2285
rect 2288 2264 2290 2285
rect 2424 2264 2426 2285
rect 2560 2264 2562 2285
rect 2704 2264 2706 2285
rect 2840 2264 2842 2285
rect 2984 2264 2986 2285
rect 3128 2264 3130 2285
rect 3272 2264 3274 2285
rect 3944 2265 3946 2285
rect 3942 2264 3948 2265
rect 2046 2260 2047 2264
rect 2051 2260 2052 2264
rect 2046 2259 2052 2260
rect 2070 2263 2076 2264
rect 2070 2259 2071 2263
rect 2075 2259 2076 2263
rect 2070 2258 2076 2259
rect 2166 2263 2172 2264
rect 2166 2259 2167 2263
rect 2171 2259 2172 2263
rect 2166 2258 2172 2259
rect 2286 2263 2292 2264
rect 2286 2259 2287 2263
rect 2291 2259 2292 2263
rect 2286 2258 2292 2259
rect 2422 2263 2428 2264
rect 2422 2259 2423 2263
rect 2427 2259 2428 2263
rect 2422 2258 2428 2259
rect 2558 2263 2564 2264
rect 2558 2259 2559 2263
rect 2563 2259 2564 2263
rect 2558 2258 2564 2259
rect 2702 2263 2708 2264
rect 2702 2259 2703 2263
rect 2707 2259 2708 2263
rect 2702 2258 2708 2259
rect 2838 2263 2844 2264
rect 2838 2259 2839 2263
rect 2843 2259 2844 2263
rect 2838 2258 2844 2259
rect 2982 2263 2988 2264
rect 2982 2259 2983 2263
rect 2987 2259 2988 2263
rect 2982 2258 2988 2259
rect 3126 2263 3132 2264
rect 3126 2259 3127 2263
rect 3131 2259 3132 2263
rect 3126 2258 3132 2259
rect 3270 2263 3276 2264
rect 3270 2259 3271 2263
rect 3275 2259 3276 2263
rect 3942 2260 3943 2264
rect 3947 2260 3948 2264
rect 3942 2259 3948 2260
rect 3270 2258 3276 2259
rect 111 2254 115 2255
rect 111 2249 115 2250
rect 415 2254 419 2255
rect 415 2249 419 2250
rect 535 2254 539 2255
rect 535 2249 539 2250
rect 647 2254 651 2255
rect 647 2249 651 2250
rect 671 2254 675 2255
rect 671 2249 675 2250
rect 767 2254 771 2255
rect 767 2249 771 2250
rect 823 2254 827 2255
rect 823 2249 827 2250
rect 895 2254 899 2255
rect 895 2249 899 2250
rect 991 2254 995 2255
rect 991 2249 995 2250
rect 1031 2254 1035 2255
rect 1031 2249 1035 2250
rect 1167 2254 1171 2255
rect 1167 2249 1171 2250
rect 1175 2254 1179 2255
rect 1175 2249 1179 2250
rect 1295 2254 1299 2255
rect 1295 2249 1299 2250
rect 1367 2254 1371 2255
rect 1367 2249 1371 2250
rect 1423 2254 1427 2255
rect 1423 2249 1427 2250
rect 1551 2254 1555 2255
rect 1551 2249 1555 2250
rect 1567 2254 1571 2255
rect 1567 2249 1571 2250
rect 1671 2254 1675 2255
rect 1671 2249 1675 2250
rect 1767 2254 1771 2255
rect 1767 2249 1771 2250
rect 1799 2254 1803 2255
rect 1799 2249 1803 2250
rect 1903 2254 1907 2255
rect 1903 2249 1907 2250
rect 2007 2254 2011 2255
rect 2007 2249 2011 2250
rect 112 2229 114 2249
rect 110 2228 116 2229
rect 416 2228 418 2249
rect 536 2228 538 2249
rect 672 2228 674 2249
rect 824 2228 826 2249
rect 992 2228 994 2249
rect 1176 2228 1178 2249
rect 1368 2228 1370 2249
rect 1568 2228 1570 2249
rect 1768 2228 1770 2249
rect 2008 2229 2010 2249
rect 2046 2247 2052 2248
rect 2046 2243 2047 2247
rect 2051 2243 2052 2247
rect 3942 2247 3948 2248
rect 2046 2242 2052 2243
rect 2070 2244 2076 2245
rect 2006 2228 2012 2229
rect 110 2224 111 2228
rect 115 2224 116 2228
rect 110 2223 116 2224
rect 414 2227 420 2228
rect 414 2223 415 2227
rect 419 2223 420 2227
rect 414 2222 420 2223
rect 534 2227 540 2228
rect 534 2223 535 2227
rect 539 2223 540 2227
rect 534 2222 540 2223
rect 670 2227 676 2228
rect 670 2223 671 2227
rect 675 2223 676 2227
rect 670 2222 676 2223
rect 822 2227 828 2228
rect 822 2223 823 2227
rect 827 2223 828 2227
rect 822 2222 828 2223
rect 990 2227 996 2228
rect 990 2223 991 2227
rect 995 2223 996 2227
rect 990 2222 996 2223
rect 1174 2227 1180 2228
rect 1174 2223 1175 2227
rect 1179 2223 1180 2227
rect 1174 2222 1180 2223
rect 1366 2227 1372 2228
rect 1366 2223 1367 2227
rect 1371 2223 1372 2227
rect 1366 2222 1372 2223
rect 1566 2227 1572 2228
rect 1566 2223 1567 2227
rect 1571 2223 1572 2227
rect 1566 2222 1572 2223
rect 1766 2227 1772 2228
rect 1766 2223 1767 2227
rect 1771 2223 1772 2227
rect 2006 2224 2007 2228
rect 2011 2224 2012 2228
rect 2006 2223 2012 2224
rect 1766 2222 1772 2223
rect 2048 2215 2050 2242
rect 2070 2240 2071 2244
rect 2075 2240 2076 2244
rect 2070 2239 2076 2240
rect 2166 2244 2172 2245
rect 2166 2240 2167 2244
rect 2171 2240 2172 2244
rect 2166 2239 2172 2240
rect 2286 2244 2292 2245
rect 2286 2240 2287 2244
rect 2291 2240 2292 2244
rect 2286 2239 2292 2240
rect 2422 2244 2428 2245
rect 2422 2240 2423 2244
rect 2427 2240 2428 2244
rect 2422 2239 2428 2240
rect 2558 2244 2564 2245
rect 2558 2240 2559 2244
rect 2563 2240 2564 2244
rect 2558 2239 2564 2240
rect 2702 2244 2708 2245
rect 2702 2240 2703 2244
rect 2707 2240 2708 2244
rect 2702 2239 2708 2240
rect 2838 2244 2844 2245
rect 2838 2240 2839 2244
rect 2843 2240 2844 2244
rect 2838 2239 2844 2240
rect 2982 2244 2988 2245
rect 2982 2240 2983 2244
rect 2987 2240 2988 2244
rect 2982 2239 2988 2240
rect 3126 2244 3132 2245
rect 3126 2240 3127 2244
rect 3131 2240 3132 2244
rect 3126 2239 3132 2240
rect 3270 2244 3276 2245
rect 3270 2240 3271 2244
rect 3275 2240 3276 2244
rect 3942 2243 3943 2247
rect 3947 2243 3948 2247
rect 3942 2242 3948 2243
rect 3270 2239 3276 2240
rect 2072 2215 2074 2239
rect 2168 2215 2170 2239
rect 2288 2215 2290 2239
rect 2424 2215 2426 2239
rect 2560 2215 2562 2239
rect 2704 2215 2706 2239
rect 2840 2215 2842 2239
rect 2984 2215 2986 2239
rect 3128 2215 3130 2239
rect 3272 2215 3274 2239
rect 3944 2215 3946 2242
rect 2047 2214 2051 2215
rect 110 2211 116 2212
rect 110 2207 111 2211
rect 115 2207 116 2211
rect 2006 2211 2012 2212
rect 110 2206 116 2207
rect 414 2208 420 2209
rect 112 2171 114 2206
rect 414 2204 415 2208
rect 419 2204 420 2208
rect 414 2203 420 2204
rect 534 2208 540 2209
rect 534 2204 535 2208
rect 539 2204 540 2208
rect 534 2203 540 2204
rect 670 2208 676 2209
rect 670 2204 671 2208
rect 675 2204 676 2208
rect 670 2203 676 2204
rect 822 2208 828 2209
rect 822 2204 823 2208
rect 827 2204 828 2208
rect 822 2203 828 2204
rect 990 2208 996 2209
rect 990 2204 991 2208
rect 995 2204 996 2208
rect 990 2203 996 2204
rect 1174 2208 1180 2209
rect 1174 2204 1175 2208
rect 1179 2204 1180 2208
rect 1174 2203 1180 2204
rect 1366 2208 1372 2209
rect 1366 2204 1367 2208
rect 1371 2204 1372 2208
rect 1366 2203 1372 2204
rect 1566 2208 1572 2209
rect 1566 2204 1567 2208
rect 1571 2204 1572 2208
rect 1566 2203 1572 2204
rect 1766 2208 1772 2209
rect 1766 2204 1767 2208
rect 1771 2204 1772 2208
rect 2006 2207 2007 2211
rect 2011 2207 2012 2211
rect 2047 2209 2051 2210
rect 2071 2214 2075 2215
rect 2071 2209 2075 2210
rect 2167 2214 2171 2215
rect 2167 2209 2171 2210
rect 2287 2214 2291 2215
rect 2287 2209 2291 2210
rect 2295 2214 2299 2215
rect 2295 2209 2299 2210
rect 2423 2214 2427 2215
rect 2423 2209 2427 2210
rect 2503 2214 2507 2215
rect 2503 2209 2507 2210
rect 2559 2214 2563 2215
rect 2559 2209 2563 2210
rect 2687 2214 2691 2215
rect 2687 2209 2691 2210
rect 2703 2214 2707 2215
rect 2703 2209 2707 2210
rect 2839 2214 2843 2215
rect 2839 2209 2843 2210
rect 2863 2214 2867 2215
rect 2863 2209 2867 2210
rect 2983 2214 2987 2215
rect 2983 2209 2987 2210
rect 3023 2214 3027 2215
rect 3023 2209 3027 2210
rect 3127 2214 3131 2215
rect 3127 2209 3131 2210
rect 3175 2214 3179 2215
rect 3175 2209 3179 2210
rect 3271 2214 3275 2215
rect 3271 2209 3275 2210
rect 3319 2214 3323 2215
rect 3319 2209 3323 2210
rect 3471 2214 3475 2215
rect 3471 2209 3475 2210
rect 3943 2214 3947 2215
rect 3943 2209 3947 2210
rect 2006 2206 2012 2207
rect 1766 2203 1772 2204
rect 416 2171 418 2203
rect 536 2171 538 2203
rect 672 2171 674 2203
rect 824 2171 826 2203
rect 992 2171 994 2203
rect 1176 2171 1178 2203
rect 1368 2171 1370 2203
rect 1568 2171 1570 2203
rect 1768 2171 1770 2203
rect 2008 2171 2010 2206
rect 2048 2182 2050 2209
rect 2072 2185 2074 2209
rect 2296 2185 2298 2209
rect 2504 2185 2506 2209
rect 2688 2185 2690 2209
rect 2864 2185 2866 2209
rect 3024 2185 3026 2209
rect 3176 2185 3178 2209
rect 3320 2185 3322 2209
rect 3472 2185 3474 2209
rect 2070 2184 2076 2185
rect 2046 2181 2052 2182
rect 2046 2177 2047 2181
rect 2051 2177 2052 2181
rect 2070 2180 2071 2184
rect 2075 2180 2076 2184
rect 2070 2179 2076 2180
rect 2294 2184 2300 2185
rect 2294 2180 2295 2184
rect 2299 2180 2300 2184
rect 2294 2179 2300 2180
rect 2502 2184 2508 2185
rect 2502 2180 2503 2184
rect 2507 2180 2508 2184
rect 2502 2179 2508 2180
rect 2686 2184 2692 2185
rect 2686 2180 2687 2184
rect 2691 2180 2692 2184
rect 2686 2179 2692 2180
rect 2862 2184 2868 2185
rect 2862 2180 2863 2184
rect 2867 2180 2868 2184
rect 2862 2179 2868 2180
rect 3022 2184 3028 2185
rect 3022 2180 3023 2184
rect 3027 2180 3028 2184
rect 3022 2179 3028 2180
rect 3174 2184 3180 2185
rect 3174 2180 3175 2184
rect 3179 2180 3180 2184
rect 3174 2179 3180 2180
rect 3318 2184 3324 2185
rect 3318 2180 3319 2184
rect 3323 2180 3324 2184
rect 3318 2179 3324 2180
rect 3470 2184 3476 2185
rect 3470 2180 3471 2184
rect 3475 2180 3476 2184
rect 3944 2182 3946 2209
rect 3470 2179 3476 2180
rect 3942 2181 3948 2182
rect 2046 2176 2052 2177
rect 3942 2177 3943 2181
rect 3947 2177 3948 2181
rect 3942 2176 3948 2177
rect 111 2170 115 2171
rect 111 2165 115 2166
rect 135 2170 139 2171
rect 135 2165 139 2166
rect 247 2170 251 2171
rect 247 2165 251 2166
rect 391 2170 395 2171
rect 391 2165 395 2166
rect 415 2170 419 2171
rect 415 2165 419 2166
rect 535 2170 539 2171
rect 535 2165 539 2166
rect 551 2170 555 2171
rect 551 2165 555 2166
rect 671 2170 675 2171
rect 671 2165 675 2166
rect 711 2170 715 2171
rect 711 2165 715 2166
rect 823 2170 827 2171
rect 823 2165 827 2166
rect 871 2170 875 2171
rect 871 2165 875 2166
rect 991 2170 995 2171
rect 991 2165 995 2166
rect 1031 2170 1035 2171
rect 1031 2165 1035 2166
rect 1175 2170 1179 2171
rect 1175 2165 1179 2166
rect 1191 2170 1195 2171
rect 1191 2165 1195 2166
rect 1351 2170 1355 2171
rect 1351 2165 1355 2166
rect 1367 2170 1371 2171
rect 1367 2165 1371 2166
rect 1511 2170 1515 2171
rect 1511 2165 1515 2166
rect 1567 2170 1571 2171
rect 1567 2165 1571 2166
rect 1679 2170 1683 2171
rect 1679 2165 1683 2166
rect 1767 2170 1771 2171
rect 1767 2165 1771 2166
rect 2007 2170 2011 2171
rect 2007 2165 2011 2166
rect 2070 2165 2076 2166
rect 112 2138 114 2165
rect 136 2141 138 2165
rect 248 2141 250 2165
rect 392 2141 394 2165
rect 552 2141 554 2165
rect 712 2141 714 2165
rect 872 2141 874 2165
rect 1032 2141 1034 2165
rect 1192 2141 1194 2165
rect 1352 2141 1354 2165
rect 1512 2141 1514 2165
rect 1680 2141 1682 2165
rect 134 2140 140 2141
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 134 2136 135 2140
rect 139 2136 140 2140
rect 134 2135 140 2136
rect 246 2140 252 2141
rect 246 2136 247 2140
rect 251 2136 252 2140
rect 246 2135 252 2136
rect 390 2140 396 2141
rect 390 2136 391 2140
rect 395 2136 396 2140
rect 390 2135 396 2136
rect 550 2140 556 2141
rect 550 2136 551 2140
rect 555 2136 556 2140
rect 550 2135 556 2136
rect 710 2140 716 2141
rect 710 2136 711 2140
rect 715 2136 716 2140
rect 710 2135 716 2136
rect 870 2140 876 2141
rect 870 2136 871 2140
rect 875 2136 876 2140
rect 870 2135 876 2136
rect 1030 2140 1036 2141
rect 1030 2136 1031 2140
rect 1035 2136 1036 2140
rect 1030 2135 1036 2136
rect 1190 2140 1196 2141
rect 1190 2136 1191 2140
rect 1195 2136 1196 2140
rect 1190 2135 1196 2136
rect 1350 2140 1356 2141
rect 1350 2136 1351 2140
rect 1355 2136 1356 2140
rect 1350 2135 1356 2136
rect 1510 2140 1516 2141
rect 1510 2136 1511 2140
rect 1515 2136 1516 2140
rect 1510 2135 1516 2136
rect 1678 2140 1684 2141
rect 1678 2136 1679 2140
rect 1683 2136 1684 2140
rect 2008 2138 2010 2165
rect 2046 2164 2052 2165
rect 2046 2160 2047 2164
rect 2051 2160 2052 2164
rect 2070 2161 2071 2165
rect 2075 2161 2076 2165
rect 2070 2160 2076 2161
rect 2294 2165 2300 2166
rect 2294 2161 2295 2165
rect 2299 2161 2300 2165
rect 2294 2160 2300 2161
rect 2502 2165 2508 2166
rect 2502 2161 2503 2165
rect 2507 2161 2508 2165
rect 2502 2160 2508 2161
rect 2686 2165 2692 2166
rect 2686 2161 2687 2165
rect 2691 2161 2692 2165
rect 2686 2160 2692 2161
rect 2862 2165 2868 2166
rect 2862 2161 2863 2165
rect 2867 2161 2868 2165
rect 2862 2160 2868 2161
rect 3022 2165 3028 2166
rect 3022 2161 3023 2165
rect 3027 2161 3028 2165
rect 3022 2160 3028 2161
rect 3174 2165 3180 2166
rect 3174 2161 3175 2165
rect 3179 2161 3180 2165
rect 3174 2160 3180 2161
rect 3318 2165 3324 2166
rect 3318 2161 3319 2165
rect 3323 2161 3324 2165
rect 3318 2160 3324 2161
rect 3470 2165 3476 2166
rect 3470 2161 3471 2165
rect 3475 2161 3476 2165
rect 3470 2160 3476 2161
rect 3942 2164 3948 2165
rect 3942 2160 3943 2164
rect 3947 2160 3948 2164
rect 2046 2159 2052 2160
rect 1678 2135 1684 2136
rect 2006 2137 2012 2138
rect 110 2132 116 2133
rect 2006 2133 2007 2137
rect 2011 2133 2012 2137
rect 2006 2132 2012 2133
rect 134 2121 140 2122
rect 110 2120 116 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 134 2117 135 2121
rect 139 2117 140 2121
rect 134 2116 140 2117
rect 246 2121 252 2122
rect 246 2117 247 2121
rect 251 2117 252 2121
rect 246 2116 252 2117
rect 390 2121 396 2122
rect 390 2117 391 2121
rect 395 2117 396 2121
rect 390 2116 396 2117
rect 550 2121 556 2122
rect 550 2117 551 2121
rect 555 2117 556 2121
rect 550 2116 556 2117
rect 710 2121 716 2122
rect 710 2117 711 2121
rect 715 2117 716 2121
rect 710 2116 716 2117
rect 870 2121 876 2122
rect 870 2117 871 2121
rect 875 2117 876 2121
rect 870 2116 876 2117
rect 1030 2121 1036 2122
rect 1030 2117 1031 2121
rect 1035 2117 1036 2121
rect 1030 2116 1036 2117
rect 1190 2121 1196 2122
rect 1190 2117 1191 2121
rect 1195 2117 1196 2121
rect 1190 2116 1196 2117
rect 1350 2121 1356 2122
rect 1350 2117 1351 2121
rect 1355 2117 1356 2121
rect 1350 2116 1356 2117
rect 1510 2121 1516 2122
rect 1510 2117 1511 2121
rect 1515 2117 1516 2121
rect 1510 2116 1516 2117
rect 1678 2121 1684 2122
rect 1678 2117 1679 2121
rect 1683 2117 1684 2121
rect 1678 2116 1684 2117
rect 2006 2120 2012 2121
rect 2006 2116 2007 2120
rect 2011 2116 2012 2120
rect 110 2115 116 2116
rect 112 2087 114 2115
rect 136 2087 138 2116
rect 248 2087 250 2116
rect 392 2087 394 2116
rect 552 2087 554 2116
rect 712 2087 714 2116
rect 872 2087 874 2116
rect 1032 2087 1034 2116
rect 1192 2087 1194 2116
rect 1352 2087 1354 2116
rect 1512 2087 1514 2116
rect 1680 2087 1682 2116
rect 2006 2115 2012 2116
rect 2048 2115 2050 2159
rect 2072 2115 2074 2160
rect 2296 2115 2298 2160
rect 2504 2115 2506 2160
rect 2688 2115 2690 2160
rect 2864 2115 2866 2160
rect 3024 2115 3026 2160
rect 3176 2115 3178 2160
rect 3320 2115 3322 2160
rect 3472 2115 3474 2160
rect 3942 2159 3948 2160
rect 3944 2115 3946 2159
rect 2008 2087 2010 2115
rect 2047 2114 2051 2115
rect 2047 2109 2051 2110
rect 2071 2114 2075 2115
rect 2071 2109 2075 2110
rect 2295 2114 2299 2115
rect 2295 2109 2299 2110
rect 2399 2114 2403 2115
rect 2399 2109 2403 2110
rect 2495 2114 2499 2115
rect 2495 2109 2499 2110
rect 2503 2114 2507 2115
rect 2503 2109 2507 2110
rect 2591 2114 2595 2115
rect 2591 2109 2595 2110
rect 2687 2114 2691 2115
rect 2687 2109 2691 2110
rect 2783 2114 2787 2115
rect 2783 2109 2787 2110
rect 2863 2114 2867 2115
rect 2863 2109 2867 2110
rect 2879 2114 2883 2115
rect 2879 2109 2883 2110
rect 2975 2114 2979 2115
rect 2975 2109 2979 2110
rect 3023 2114 3027 2115
rect 3023 2109 3027 2110
rect 3071 2114 3075 2115
rect 3071 2109 3075 2110
rect 3167 2114 3171 2115
rect 3167 2109 3171 2110
rect 3175 2114 3179 2115
rect 3175 2109 3179 2110
rect 3263 2114 3267 2115
rect 3263 2109 3267 2110
rect 3319 2114 3323 2115
rect 3319 2109 3323 2110
rect 3359 2114 3363 2115
rect 3359 2109 3363 2110
rect 3455 2114 3459 2115
rect 3455 2109 3459 2110
rect 3471 2114 3475 2115
rect 3471 2109 3475 2110
rect 3551 2114 3555 2115
rect 3551 2109 3555 2110
rect 3647 2114 3651 2115
rect 3647 2109 3651 2110
rect 3743 2114 3747 2115
rect 3743 2109 3747 2110
rect 3839 2114 3843 2115
rect 3839 2109 3843 2110
rect 3943 2114 3947 2115
rect 3943 2109 3947 2110
rect 2048 2089 2050 2109
rect 2046 2088 2052 2089
rect 2400 2088 2402 2109
rect 2496 2088 2498 2109
rect 2592 2088 2594 2109
rect 2688 2088 2690 2109
rect 2784 2088 2786 2109
rect 2880 2088 2882 2109
rect 2976 2088 2978 2109
rect 3072 2088 3074 2109
rect 3168 2088 3170 2109
rect 3264 2088 3266 2109
rect 3360 2088 3362 2109
rect 3456 2088 3458 2109
rect 3552 2088 3554 2109
rect 3648 2088 3650 2109
rect 3744 2088 3746 2109
rect 3840 2088 3842 2109
rect 3944 2089 3946 2109
rect 3942 2088 3948 2089
rect 111 2086 115 2087
rect 111 2081 115 2082
rect 135 2086 139 2087
rect 135 2081 139 2082
rect 247 2086 251 2087
rect 247 2081 251 2082
rect 391 2086 395 2087
rect 391 2081 395 2082
rect 399 2086 403 2087
rect 399 2081 403 2082
rect 551 2086 555 2087
rect 551 2081 555 2082
rect 703 2086 707 2087
rect 703 2081 707 2082
rect 711 2086 715 2087
rect 711 2081 715 2082
rect 847 2086 851 2087
rect 847 2081 851 2082
rect 871 2086 875 2087
rect 871 2081 875 2082
rect 991 2086 995 2087
rect 991 2081 995 2082
rect 1031 2086 1035 2087
rect 1031 2081 1035 2082
rect 1127 2086 1131 2087
rect 1127 2081 1131 2082
rect 1191 2086 1195 2087
rect 1191 2081 1195 2082
rect 1255 2086 1259 2087
rect 1255 2081 1259 2082
rect 1351 2086 1355 2087
rect 1351 2081 1355 2082
rect 1383 2086 1387 2087
rect 1383 2081 1387 2082
rect 1511 2086 1515 2087
rect 1511 2081 1515 2082
rect 1519 2086 1523 2087
rect 1519 2081 1523 2082
rect 1679 2086 1683 2087
rect 1679 2081 1683 2082
rect 2007 2086 2011 2087
rect 2046 2084 2047 2088
rect 2051 2084 2052 2088
rect 2046 2083 2052 2084
rect 2398 2087 2404 2088
rect 2398 2083 2399 2087
rect 2403 2083 2404 2087
rect 2398 2082 2404 2083
rect 2494 2087 2500 2088
rect 2494 2083 2495 2087
rect 2499 2083 2500 2087
rect 2494 2082 2500 2083
rect 2590 2087 2596 2088
rect 2590 2083 2591 2087
rect 2595 2083 2596 2087
rect 2590 2082 2596 2083
rect 2686 2087 2692 2088
rect 2686 2083 2687 2087
rect 2691 2083 2692 2087
rect 2686 2082 2692 2083
rect 2782 2087 2788 2088
rect 2782 2083 2783 2087
rect 2787 2083 2788 2087
rect 2782 2082 2788 2083
rect 2878 2087 2884 2088
rect 2878 2083 2879 2087
rect 2883 2083 2884 2087
rect 2878 2082 2884 2083
rect 2974 2087 2980 2088
rect 2974 2083 2975 2087
rect 2979 2083 2980 2087
rect 2974 2082 2980 2083
rect 3070 2087 3076 2088
rect 3070 2083 3071 2087
rect 3075 2083 3076 2087
rect 3070 2082 3076 2083
rect 3166 2087 3172 2088
rect 3166 2083 3167 2087
rect 3171 2083 3172 2087
rect 3166 2082 3172 2083
rect 3262 2087 3268 2088
rect 3262 2083 3263 2087
rect 3267 2083 3268 2087
rect 3262 2082 3268 2083
rect 3358 2087 3364 2088
rect 3358 2083 3359 2087
rect 3363 2083 3364 2087
rect 3358 2082 3364 2083
rect 3454 2087 3460 2088
rect 3454 2083 3455 2087
rect 3459 2083 3460 2087
rect 3454 2082 3460 2083
rect 3550 2087 3556 2088
rect 3550 2083 3551 2087
rect 3555 2083 3556 2087
rect 3550 2082 3556 2083
rect 3646 2087 3652 2088
rect 3646 2083 3647 2087
rect 3651 2083 3652 2087
rect 3646 2082 3652 2083
rect 3742 2087 3748 2088
rect 3742 2083 3743 2087
rect 3747 2083 3748 2087
rect 3742 2082 3748 2083
rect 3838 2087 3844 2088
rect 3838 2083 3839 2087
rect 3843 2083 3844 2087
rect 3942 2084 3943 2088
rect 3947 2084 3948 2088
rect 3942 2083 3948 2084
rect 3838 2082 3844 2083
rect 2007 2081 2011 2082
rect 112 2061 114 2081
rect 110 2060 116 2061
rect 136 2060 138 2081
rect 248 2060 250 2081
rect 400 2060 402 2081
rect 552 2060 554 2081
rect 704 2060 706 2081
rect 848 2060 850 2081
rect 992 2060 994 2081
rect 1128 2060 1130 2081
rect 1256 2060 1258 2081
rect 1384 2060 1386 2081
rect 1520 2060 1522 2081
rect 2008 2061 2010 2081
rect 2046 2071 2052 2072
rect 2046 2067 2047 2071
rect 2051 2067 2052 2071
rect 3942 2071 3948 2072
rect 2046 2066 2052 2067
rect 2398 2068 2404 2069
rect 2006 2060 2012 2061
rect 110 2056 111 2060
rect 115 2056 116 2060
rect 110 2055 116 2056
rect 134 2059 140 2060
rect 134 2055 135 2059
rect 139 2055 140 2059
rect 134 2054 140 2055
rect 246 2059 252 2060
rect 246 2055 247 2059
rect 251 2055 252 2059
rect 246 2054 252 2055
rect 398 2059 404 2060
rect 398 2055 399 2059
rect 403 2055 404 2059
rect 398 2054 404 2055
rect 550 2059 556 2060
rect 550 2055 551 2059
rect 555 2055 556 2059
rect 550 2054 556 2055
rect 702 2059 708 2060
rect 702 2055 703 2059
rect 707 2055 708 2059
rect 702 2054 708 2055
rect 846 2059 852 2060
rect 846 2055 847 2059
rect 851 2055 852 2059
rect 846 2054 852 2055
rect 990 2059 996 2060
rect 990 2055 991 2059
rect 995 2055 996 2059
rect 990 2054 996 2055
rect 1126 2059 1132 2060
rect 1126 2055 1127 2059
rect 1131 2055 1132 2059
rect 1126 2054 1132 2055
rect 1254 2059 1260 2060
rect 1254 2055 1255 2059
rect 1259 2055 1260 2059
rect 1254 2054 1260 2055
rect 1382 2059 1388 2060
rect 1382 2055 1383 2059
rect 1387 2055 1388 2059
rect 1382 2054 1388 2055
rect 1518 2059 1524 2060
rect 1518 2055 1519 2059
rect 1523 2055 1524 2059
rect 2006 2056 2007 2060
rect 2011 2056 2012 2060
rect 2006 2055 2012 2056
rect 1518 2054 1524 2055
rect 110 2043 116 2044
rect 110 2039 111 2043
rect 115 2039 116 2043
rect 2006 2043 2012 2044
rect 110 2038 116 2039
rect 134 2040 140 2041
rect 112 1995 114 2038
rect 134 2036 135 2040
rect 139 2036 140 2040
rect 134 2035 140 2036
rect 246 2040 252 2041
rect 246 2036 247 2040
rect 251 2036 252 2040
rect 246 2035 252 2036
rect 398 2040 404 2041
rect 398 2036 399 2040
rect 403 2036 404 2040
rect 398 2035 404 2036
rect 550 2040 556 2041
rect 550 2036 551 2040
rect 555 2036 556 2040
rect 550 2035 556 2036
rect 702 2040 708 2041
rect 702 2036 703 2040
rect 707 2036 708 2040
rect 702 2035 708 2036
rect 846 2040 852 2041
rect 846 2036 847 2040
rect 851 2036 852 2040
rect 846 2035 852 2036
rect 990 2040 996 2041
rect 990 2036 991 2040
rect 995 2036 996 2040
rect 990 2035 996 2036
rect 1126 2040 1132 2041
rect 1126 2036 1127 2040
rect 1131 2036 1132 2040
rect 1126 2035 1132 2036
rect 1254 2040 1260 2041
rect 1254 2036 1255 2040
rect 1259 2036 1260 2040
rect 1254 2035 1260 2036
rect 1382 2040 1388 2041
rect 1382 2036 1383 2040
rect 1387 2036 1388 2040
rect 1382 2035 1388 2036
rect 1518 2040 1524 2041
rect 1518 2036 1519 2040
rect 1523 2036 1524 2040
rect 2006 2039 2007 2043
rect 2011 2039 2012 2043
rect 2048 2039 2050 2066
rect 2398 2064 2399 2068
rect 2403 2064 2404 2068
rect 2398 2063 2404 2064
rect 2494 2068 2500 2069
rect 2494 2064 2495 2068
rect 2499 2064 2500 2068
rect 2494 2063 2500 2064
rect 2590 2068 2596 2069
rect 2590 2064 2591 2068
rect 2595 2064 2596 2068
rect 2590 2063 2596 2064
rect 2686 2068 2692 2069
rect 2686 2064 2687 2068
rect 2691 2064 2692 2068
rect 2686 2063 2692 2064
rect 2782 2068 2788 2069
rect 2782 2064 2783 2068
rect 2787 2064 2788 2068
rect 2782 2063 2788 2064
rect 2878 2068 2884 2069
rect 2878 2064 2879 2068
rect 2883 2064 2884 2068
rect 2878 2063 2884 2064
rect 2974 2068 2980 2069
rect 2974 2064 2975 2068
rect 2979 2064 2980 2068
rect 2974 2063 2980 2064
rect 3070 2068 3076 2069
rect 3070 2064 3071 2068
rect 3075 2064 3076 2068
rect 3070 2063 3076 2064
rect 3166 2068 3172 2069
rect 3166 2064 3167 2068
rect 3171 2064 3172 2068
rect 3166 2063 3172 2064
rect 3262 2068 3268 2069
rect 3262 2064 3263 2068
rect 3267 2064 3268 2068
rect 3262 2063 3268 2064
rect 3358 2068 3364 2069
rect 3358 2064 3359 2068
rect 3363 2064 3364 2068
rect 3358 2063 3364 2064
rect 3454 2068 3460 2069
rect 3454 2064 3455 2068
rect 3459 2064 3460 2068
rect 3454 2063 3460 2064
rect 3550 2068 3556 2069
rect 3550 2064 3551 2068
rect 3555 2064 3556 2068
rect 3550 2063 3556 2064
rect 3646 2068 3652 2069
rect 3646 2064 3647 2068
rect 3651 2064 3652 2068
rect 3646 2063 3652 2064
rect 3742 2068 3748 2069
rect 3742 2064 3743 2068
rect 3747 2064 3748 2068
rect 3742 2063 3748 2064
rect 3838 2068 3844 2069
rect 3838 2064 3839 2068
rect 3843 2064 3844 2068
rect 3942 2067 3943 2071
rect 3947 2067 3948 2071
rect 3942 2066 3948 2067
rect 3838 2063 3844 2064
rect 2400 2039 2402 2063
rect 2496 2039 2498 2063
rect 2592 2039 2594 2063
rect 2688 2039 2690 2063
rect 2784 2039 2786 2063
rect 2880 2039 2882 2063
rect 2976 2039 2978 2063
rect 3072 2039 3074 2063
rect 3168 2039 3170 2063
rect 3264 2039 3266 2063
rect 3360 2039 3362 2063
rect 3456 2039 3458 2063
rect 3552 2039 3554 2063
rect 3648 2039 3650 2063
rect 3744 2039 3746 2063
rect 3840 2039 3842 2063
rect 3944 2039 3946 2066
rect 2006 2038 2012 2039
rect 2047 2038 2051 2039
rect 1518 2035 1524 2036
rect 136 1995 138 2035
rect 248 1995 250 2035
rect 400 1995 402 2035
rect 552 1995 554 2035
rect 704 1995 706 2035
rect 848 1995 850 2035
rect 992 1995 994 2035
rect 1128 1995 1130 2035
rect 1256 1995 1258 2035
rect 1384 1995 1386 2035
rect 1520 1995 1522 2035
rect 2008 1995 2010 2038
rect 2047 2033 2051 2034
rect 2191 2038 2195 2039
rect 2191 2033 2195 2034
rect 2399 2038 2403 2039
rect 2399 2033 2403 2034
rect 2495 2038 2499 2039
rect 2495 2033 2499 2034
rect 2591 2038 2595 2039
rect 2591 2033 2595 2034
rect 2647 2038 2651 2039
rect 2647 2033 2651 2034
rect 2687 2038 2691 2039
rect 2687 2033 2691 2034
rect 2783 2038 2787 2039
rect 2783 2033 2787 2034
rect 2879 2038 2883 2039
rect 2879 2033 2883 2034
rect 2919 2038 2923 2039
rect 2919 2033 2923 2034
rect 2975 2038 2979 2039
rect 2975 2033 2979 2034
rect 3071 2038 3075 2039
rect 3071 2033 3075 2034
rect 3167 2038 3171 2039
rect 3167 2033 3171 2034
rect 3215 2038 3219 2039
rect 3215 2033 3219 2034
rect 3263 2038 3267 2039
rect 3263 2033 3267 2034
rect 3359 2038 3363 2039
rect 3359 2033 3363 2034
rect 3455 2038 3459 2039
rect 3455 2033 3459 2034
rect 3527 2038 3531 2039
rect 3527 2033 3531 2034
rect 3551 2038 3555 2039
rect 3551 2033 3555 2034
rect 3647 2038 3651 2039
rect 3647 2033 3651 2034
rect 3743 2038 3747 2039
rect 3743 2033 3747 2034
rect 3839 2038 3843 2039
rect 3839 2033 3843 2034
rect 3943 2038 3947 2039
rect 3943 2033 3947 2034
rect 2048 2006 2050 2033
rect 2192 2009 2194 2033
rect 2400 2009 2402 2033
rect 2648 2009 2650 2033
rect 2920 2009 2922 2033
rect 3216 2009 3218 2033
rect 3528 2009 3530 2033
rect 3840 2009 3842 2033
rect 2190 2008 2196 2009
rect 2046 2005 2052 2006
rect 2046 2001 2047 2005
rect 2051 2001 2052 2005
rect 2190 2004 2191 2008
rect 2195 2004 2196 2008
rect 2190 2003 2196 2004
rect 2398 2008 2404 2009
rect 2398 2004 2399 2008
rect 2403 2004 2404 2008
rect 2398 2003 2404 2004
rect 2646 2008 2652 2009
rect 2646 2004 2647 2008
rect 2651 2004 2652 2008
rect 2646 2003 2652 2004
rect 2918 2008 2924 2009
rect 2918 2004 2919 2008
rect 2923 2004 2924 2008
rect 2918 2003 2924 2004
rect 3214 2008 3220 2009
rect 3214 2004 3215 2008
rect 3219 2004 3220 2008
rect 3214 2003 3220 2004
rect 3526 2008 3532 2009
rect 3526 2004 3527 2008
rect 3531 2004 3532 2008
rect 3526 2003 3532 2004
rect 3838 2008 3844 2009
rect 3838 2004 3839 2008
rect 3843 2004 3844 2008
rect 3944 2006 3946 2033
rect 3838 2003 3844 2004
rect 3942 2005 3948 2006
rect 2046 2000 2052 2001
rect 3942 2001 3943 2005
rect 3947 2001 3948 2005
rect 3942 2000 3948 2001
rect 111 1994 115 1995
rect 111 1989 115 1990
rect 135 1994 139 1995
rect 135 1989 139 1990
rect 231 1994 235 1995
rect 231 1989 235 1990
rect 247 1994 251 1995
rect 247 1989 251 1990
rect 391 1994 395 1995
rect 391 1989 395 1990
rect 399 1994 403 1995
rect 399 1989 403 1990
rect 551 1994 555 1995
rect 551 1989 555 1990
rect 567 1994 571 1995
rect 567 1989 571 1990
rect 703 1994 707 1995
rect 703 1989 707 1990
rect 751 1994 755 1995
rect 751 1989 755 1990
rect 847 1994 851 1995
rect 847 1989 851 1990
rect 943 1994 947 1995
rect 943 1989 947 1990
rect 991 1994 995 1995
rect 991 1989 995 1990
rect 1127 1994 1131 1995
rect 1127 1989 1131 1990
rect 1135 1994 1139 1995
rect 1135 1989 1139 1990
rect 1255 1994 1259 1995
rect 1255 1989 1259 1990
rect 1335 1994 1339 1995
rect 1335 1989 1339 1990
rect 1383 1994 1387 1995
rect 1383 1989 1387 1990
rect 1519 1994 1523 1995
rect 1519 1989 1523 1990
rect 1543 1994 1547 1995
rect 1543 1989 1547 1990
rect 2007 1994 2011 1995
rect 2007 1989 2011 1990
rect 2190 1989 2196 1990
rect 112 1962 114 1989
rect 232 1965 234 1989
rect 392 1965 394 1989
rect 568 1965 570 1989
rect 752 1965 754 1989
rect 944 1965 946 1989
rect 1136 1965 1138 1989
rect 1336 1965 1338 1989
rect 1544 1965 1546 1989
rect 230 1964 236 1965
rect 110 1961 116 1962
rect 110 1957 111 1961
rect 115 1957 116 1961
rect 230 1960 231 1964
rect 235 1960 236 1964
rect 230 1959 236 1960
rect 390 1964 396 1965
rect 390 1960 391 1964
rect 395 1960 396 1964
rect 390 1959 396 1960
rect 566 1964 572 1965
rect 566 1960 567 1964
rect 571 1960 572 1964
rect 566 1959 572 1960
rect 750 1964 756 1965
rect 750 1960 751 1964
rect 755 1960 756 1964
rect 750 1959 756 1960
rect 942 1964 948 1965
rect 942 1960 943 1964
rect 947 1960 948 1964
rect 942 1959 948 1960
rect 1134 1964 1140 1965
rect 1134 1960 1135 1964
rect 1139 1960 1140 1964
rect 1134 1959 1140 1960
rect 1334 1964 1340 1965
rect 1334 1960 1335 1964
rect 1339 1960 1340 1964
rect 1334 1959 1340 1960
rect 1542 1964 1548 1965
rect 1542 1960 1543 1964
rect 1547 1960 1548 1964
rect 2008 1962 2010 1989
rect 2046 1988 2052 1989
rect 2046 1984 2047 1988
rect 2051 1984 2052 1988
rect 2190 1985 2191 1989
rect 2195 1985 2196 1989
rect 2190 1984 2196 1985
rect 2398 1989 2404 1990
rect 2398 1985 2399 1989
rect 2403 1985 2404 1989
rect 2398 1984 2404 1985
rect 2646 1989 2652 1990
rect 2646 1985 2647 1989
rect 2651 1985 2652 1989
rect 2646 1984 2652 1985
rect 2918 1989 2924 1990
rect 2918 1985 2919 1989
rect 2923 1985 2924 1989
rect 2918 1984 2924 1985
rect 3214 1989 3220 1990
rect 3214 1985 3215 1989
rect 3219 1985 3220 1989
rect 3214 1984 3220 1985
rect 3526 1989 3532 1990
rect 3526 1985 3527 1989
rect 3531 1985 3532 1989
rect 3526 1984 3532 1985
rect 3838 1989 3844 1990
rect 3838 1985 3839 1989
rect 3843 1985 3844 1989
rect 3838 1984 3844 1985
rect 3942 1988 3948 1989
rect 3942 1984 3943 1988
rect 3947 1984 3948 1988
rect 2046 1983 2052 1984
rect 1542 1959 1548 1960
rect 2006 1961 2012 1962
rect 110 1956 116 1957
rect 2006 1957 2007 1961
rect 2011 1957 2012 1961
rect 2006 1956 2012 1957
rect 2048 1951 2050 1983
rect 2192 1951 2194 1984
rect 2400 1951 2402 1984
rect 2648 1951 2650 1984
rect 2920 1951 2922 1984
rect 3216 1951 3218 1984
rect 3528 1951 3530 1984
rect 3840 1951 3842 1984
rect 3942 1983 3948 1984
rect 3944 1951 3946 1983
rect 2047 1950 2051 1951
rect 230 1945 236 1946
rect 110 1944 116 1945
rect 110 1940 111 1944
rect 115 1940 116 1944
rect 230 1941 231 1945
rect 235 1941 236 1945
rect 230 1940 236 1941
rect 390 1945 396 1946
rect 390 1941 391 1945
rect 395 1941 396 1945
rect 390 1940 396 1941
rect 566 1945 572 1946
rect 566 1941 567 1945
rect 571 1941 572 1945
rect 566 1940 572 1941
rect 750 1945 756 1946
rect 750 1941 751 1945
rect 755 1941 756 1945
rect 750 1940 756 1941
rect 942 1945 948 1946
rect 942 1941 943 1945
rect 947 1941 948 1945
rect 942 1940 948 1941
rect 1134 1945 1140 1946
rect 1134 1941 1135 1945
rect 1139 1941 1140 1945
rect 1134 1940 1140 1941
rect 1334 1945 1340 1946
rect 1334 1941 1335 1945
rect 1339 1941 1340 1945
rect 1334 1940 1340 1941
rect 1542 1945 1548 1946
rect 2047 1945 2051 1946
rect 2071 1950 2075 1951
rect 2071 1945 2075 1946
rect 2191 1950 2195 1951
rect 2191 1945 2195 1946
rect 2239 1950 2243 1951
rect 2239 1945 2243 1946
rect 2399 1950 2403 1951
rect 2399 1945 2403 1946
rect 2447 1950 2451 1951
rect 2447 1945 2451 1946
rect 2647 1950 2651 1951
rect 2647 1945 2651 1946
rect 2671 1950 2675 1951
rect 2671 1945 2675 1946
rect 2895 1950 2899 1951
rect 2895 1945 2899 1946
rect 2919 1950 2923 1951
rect 2919 1945 2923 1946
rect 3127 1950 3131 1951
rect 3127 1945 3131 1946
rect 3215 1950 3219 1951
rect 3215 1945 3219 1946
rect 3359 1950 3363 1951
rect 3359 1945 3363 1946
rect 3527 1950 3531 1951
rect 3527 1945 3531 1946
rect 3591 1950 3595 1951
rect 3591 1945 3595 1946
rect 3831 1950 3835 1951
rect 3831 1945 3835 1946
rect 3839 1950 3843 1951
rect 3839 1945 3843 1946
rect 3943 1950 3947 1951
rect 3943 1945 3947 1946
rect 1542 1941 1543 1945
rect 1547 1941 1548 1945
rect 1542 1940 1548 1941
rect 2006 1944 2012 1945
rect 2006 1940 2007 1944
rect 2011 1940 2012 1944
rect 110 1939 116 1940
rect 112 1919 114 1939
rect 232 1919 234 1940
rect 392 1919 394 1940
rect 568 1919 570 1940
rect 752 1919 754 1940
rect 944 1919 946 1940
rect 1136 1919 1138 1940
rect 1336 1919 1338 1940
rect 1544 1919 1546 1940
rect 2006 1939 2012 1940
rect 2008 1919 2010 1939
rect 2048 1925 2050 1945
rect 2046 1924 2052 1925
rect 2072 1924 2074 1945
rect 2240 1924 2242 1945
rect 2448 1924 2450 1945
rect 2672 1924 2674 1945
rect 2896 1924 2898 1945
rect 3128 1924 3130 1945
rect 3360 1924 3362 1945
rect 3592 1924 3594 1945
rect 3832 1924 3834 1945
rect 3944 1925 3946 1945
rect 3942 1924 3948 1925
rect 2046 1920 2047 1924
rect 2051 1920 2052 1924
rect 2046 1919 2052 1920
rect 2070 1923 2076 1924
rect 2070 1919 2071 1923
rect 2075 1919 2076 1923
rect 111 1918 115 1919
rect 111 1913 115 1914
rect 231 1918 235 1919
rect 231 1913 235 1914
rect 391 1918 395 1919
rect 391 1913 395 1914
rect 511 1918 515 1919
rect 511 1913 515 1914
rect 567 1918 571 1919
rect 567 1913 571 1914
rect 623 1918 627 1919
rect 623 1913 627 1914
rect 743 1918 747 1919
rect 743 1913 747 1914
rect 751 1918 755 1919
rect 751 1913 755 1914
rect 863 1918 867 1919
rect 863 1913 867 1914
rect 943 1918 947 1919
rect 943 1913 947 1914
rect 983 1918 987 1919
rect 983 1913 987 1914
rect 1103 1918 1107 1919
rect 1103 1913 1107 1914
rect 1135 1918 1139 1919
rect 1135 1913 1139 1914
rect 1223 1918 1227 1919
rect 1223 1913 1227 1914
rect 1335 1918 1339 1919
rect 1335 1913 1339 1914
rect 1455 1918 1459 1919
rect 1455 1913 1459 1914
rect 1543 1918 1547 1919
rect 1543 1913 1547 1914
rect 1575 1918 1579 1919
rect 1575 1913 1579 1914
rect 1695 1918 1699 1919
rect 1695 1913 1699 1914
rect 2007 1918 2011 1919
rect 2070 1918 2076 1919
rect 2238 1923 2244 1924
rect 2238 1919 2239 1923
rect 2243 1919 2244 1923
rect 2238 1918 2244 1919
rect 2446 1923 2452 1924
rect 2446 1919 2447 1923
rect 2451 1919 2452 1923
rect 2446 1918 2452 1919
rect 2670 1923 2676 1924
rect 2670 1919 2671 1923
rect 2675 1919 2676 1923
rect 2670 1918 2676 1919
rect 2894 1923 2900 1924
rect 2894 1919 2895 1923
rect 2899 1919 2900 1923
rect 2894 1918 2900 1919
rect 3126 1923 3132 1924
rect 3126 1919 3127 1923
rect 3131 1919 3132 1923
rect 3126 1918 3132 1919
rect 3358 1923 3364 1924
rect 3358 1919 3359 1923
rect 3363 1919 3364 1923
rect 3358 1918 3364 1919
rect 3590 1923 3596 1924
rect 3590 1919 3591 1923
rect 3595 1919 3596 1923
rect 3590 1918 3596 1919
rect 3830 1923 3836 1924
rect 3830 1919 3831 1923
rect 3835 1919 3836 1923
rect 3942 1920 3943 1924
rect 3947 1920 3948 1924
rect 3942 1919 3948 1920
rect 3830 1918 3836 1919
rect 2007 1913 2011 1914
rect 112 1893 114 1913
rect 110 1892 116 1893
rect 512 1892 514 1913
rect 624 1892 626 1913
rect 744 1892 746 1913
rect 864 1892 866 1913
rect 984 1892 986 1913
rect 1104 1892 1106 1913
rect 1224 1892 1226 1913
rect 1336 1892 1338 1913
rect 1456 1892 1458 1913
rect 1576 1892 1578 1913
rect 1696 1892 1698 1913
rect 2008 1893 2010 1913
rect 2046 1907 2052 1908
rect 2046 1903 2047 1907
rect 2051 1903 2052 1907
rect 3942 1907 3948 1908
rect 2046 1902 2052 1903
rect 2070 1904 2076 1905
rect 2006 1892 2012 1893
rect 110 1888 111 1892
rect 115 1888 116 1892
rect 110 1887 116 1888
rect 510 1891 516 1892
rect 510 1887 511 1891
rect 515 1887 516 1891
rect 510 1886 516 1887
rect 622 1891 628 1892
rect 622 1887 623 1891
rect 627 1887 628 1891
rect 622 1886 628 1887
rect 742 1891 748 1892
rect 742 1887 743 1891
rect 747 1887 748 1891
rect 742 1886 748 1887
rect 862 1891 868 1892
rect 862 1887 863 1891
rect 867 1887 868 1891
rect 862 1886 868 1887
rect 982 1891 988 1892
rect 982 1887 983 1891
rect 987 1887 988 1891
rect 982 1886 988 1887
rect 1102 1891 1108 1892
rect 1102 1887 1103 1891
rect 1107 1887 1108 1891
rect 1102 1886 1108 1887
rect 1222 1891 1228 1892
rect 1222 1887 1223 1891
rect 1227 1887 1228 1891
rect 1222 1886 1228 1887
rect 1334 1891 1340 1892
rect 1334 1887 1335 1891
rect 1339 1887 1340 1891
rect 1334 1886 1340 1887
rect 1454 1891 1460 1892
rect 1454 1887 1455 1891
rect 1459 1887 1460 1891
rect 1454 1886 1460 1887
rect 1574 1891 1580 1892
rect 1574 1887 1575 1891
rect 1579 1887 1580 1891
rect 1574 1886 1580 1887
rect 1694 1891 1700 1892
rect 1694 1887 1695 1891
rect 1699 1887 1700 1891
rect 2006 1888 2007 1892
rect 2011 1888 2012 1892
rect 2006 1887 2012 1888
rect 1694 1886 1700 1887
rect 110 1875 116 1876
rect 110 1871 111 1875
rect 115 1871 116 1875
rect 2006 1875 2012 1876
rect 2048 1875 2050 1902
rect 2070 1900 2071 1904
rect 2075 1900 2076 1904
rect 2070 1899 2076 1900
rect 2238 1904 2244 1905
rect 2238 1900 2239 1904
rect 2243 1900 2244 1904
rect 2238 1899 2244 1900
rect 2446 1904 2452 1905
rect 2446 1900 2447 1904
rect 2451 1900 2452 1904
rect 2446 1899 2452 1900
rect 2670 1904 2676 1905
rect 2670 1900 2671 1904
rect 2675 1900 2676 1904
rect 2670 1899 2676 1900
rect 2894 1904 2900 1905
rect 2894 1900 2895 1904
rect 2899 1900 2900 1904
rect 2894 1899 2900 1900
rect 3126 1904 3132 1905
rect 3126 1900 3127 1904
rect 3131 1900 3132 1904
rect 3126 1899 3132 1900
rect 3358 1904 3364 1905
rect 3358 1900 3359 1904
rect 3363 1900 3364 1904
rect 3358 1899 3364 1900
rect 3590 1904 3596 1905
rect 3590 1900 3591 1904
rect 3595 1900 3596 1904
rect 3590 1899 3596 1900
rect 3830 1904 3836 1905
rect 3830 1900 3831 1904
rect 3835 1900 3836 1904
rect 3942 1903 3943 1907
rect 3947 1903 3948 1907
rect 3942 1902 3948 1903
rect 3830 1899 3836 1900
rect 2072 1875 2074 1899
rect 2240 1875 2242 1899
rect 2448 1875 2450 1899
rect 2672 1875 2674 1899
rect 2896 1875 2898 1899
rect 3128 1875 3130 1899
rect 3360 1875 3362 1899
rect 3592 1875 3594 1899
rect 3832 1875 3834 1899
rect 3944 1875 3946 1902
rect 110 1870 116 1871
rect 510 1872 516 1873
rect 112 1835 114 1870
rect 510 1868 511 1872
rect 515 1868 516 1872
rect 510 1867 516 1868
rect 622 1872 628 1873
rect 622 1868 623 1872
rect 627 1868 628 1872
rect 622 1867 628 1868
rect 742 1872 748 1873
rect 742 1868 743 1872
rect 747 1868 748 1872
rect 742 1867 748 1868
rect 862 1872 868 1873
rect 862 1868 863 1872
rect 867 1868 868 1872
rect 862 1867 868 1868
rect 982 1872 988 1873
rect 982 1868 983 1872
rect 987 1868 988 1872
rect 982 1867 988 1868
rect 1102 1872 1108 1873
rect 1102 1868 1103 1872
rect 1107 1868 1108 1872
rect 1102 1867 1108 1868
rect 1222 1872 1228 1873
rect 1222 1868 1223 1872
rect 1227 1868 1228 1872
rect 1222 1867 1228 1868
rect 1334 1872 1340 1873
rect 1334 1868 1335 1872
rect 1339 1868 1340 1872
rect 1334 1867 1340 1868
rect 1454 1872 1460 1873
rect 1454 1868 1455 1872
rect 1459 1868 1460 1872
rect 1454 1867 1460 1868
rect 1574 1872 1580 1873
rect 1574 1868 1575 1872
rect 1579 1868 1580 1872
rect 1574 1867 1580 1868
rect 1694 1872 1700 1873
rect 1694 1868 1695 1872
rect 1699 1868 1700 1872
rect 2006 1871 2007 1875
rect 2011 1871 2012 1875
rect 2006 1870 2012 1871
rect 2047 1874 2051 1875
rect 1694 1867 1700 1868
rect 512 1835 514 1867
rect 624 1835 626 1867
rect 744 1835 746 1867
rect 864 1835 866 1867
rect 984 1835 986 1867
rect 1104 1835 1106 1867
rect 1224 1835 1226 1867
rect 1336 1835 1338 1867
rect 1456 1835 1458 1867
rect 1576 1835 1578 1867
rect 1696 1835 1698 1867
rect 2008 1835 2010 1870
rect 2047 1869 2051 1870
rect 2071 1874 2075 1875
rect 2071 1869 2075 1870
rect 2199 1874 2203 1875
rect 2199 1869 2203 1870
rect 2239 1874 2243 1875
rect 2239 1869 2243 1870
rect 2367 1874 2371 1875
rect 2367 1869 2371 1870
rect 2447 1874 2451 1875
rect 2447 1869 2451 1870
rect 2543 1874 2547 1875
rect 2543 1869 2547 1870
rect 2671 1874 2675 1875
rect 2671 1869 2675 1870
rect 2719 1874 2723 1875
rect 2719 1869 2723 1870
rect 2887 1874 2891 1875
rect 2887 1869 2891 1870
rect 2895 1874 2899 1875
rect 2895 1869 2899 1870
rect 3039 1874 3043 1875
rect 3039 1869 3043 1870
rect 3127 1874 3131 1875
rect 3127 1869 3131 1870
rect 3183 1874 3187 1875
rect 3183 1869 3187 1870
rect 3319 1874 3323 1875
rect 3319 1869 3323 1870
rect 3359 1874 3363 1875
rect 3359 1869 3363 1870
rect 3455 1874 3459 1875
rect 3455 1869 3459 1870
rect 3583 1874 3587 1875
rect 3583 1869 3587 1870
rect 3591 1874 3595 1875
rect 3591 1869 3595 1870
rect 3711 1874 3715 1875
rect 3711 1869 3715 1870
rect 3831 1874 3835 1875
rect 3831 1869 3835 1870
rect 3839 1874 3843 1875
rect 3839 1869 3843 1870
rect 3943 1874 3947 1875
rect 3943 1869 3947 1870
rect 2048 1842 2050 1869
rect 2072 1845 2074 1869
rect 2200 1845 2202 1869
rect 2368 1845 2370 1869
rect 2544 1845 2546 1869
rect 2720 1845 2722 1869
rect 2888 1845 2890 1869
rect 3040 1845 3042 1869
rect 3184 1845 3186 1869
rect 3320 1845 3322 1869
rect 3456 1845 3458 1869
rect 3584 1845 3586 1869
rect 3712 1845 3714 1869
rect 3840 1845 3842 1869
rect 2070 1844 2076 1845
rect 2046 1841 2052 1842
rect 2046 1837 2047 1841
rect 2051 1837 2052 1841
rect 2070 1840 2071 1844
rect 2075 1840 2076 1844
rect 2070 1839 2076 1840
rect 2198 1844 2204 1845
rect 2198 1840 2199 1844
rect 2203 1840 2204 1844
rect 2198 1839 2204 1840
rect 2366 1844 2372 1845
rect 2366 1840 2367 1844
rect 2371 1840 2372 1844
rect 2366 1839 2372 1840
rect 2542 1844 2548 1845
rect 2542 1840 2543 1844
rect 2547 1840 2548 1844
rect 2542 1839 2548 1840
rect 2718 1844 2724 1845
rect 2718 1840 2719 1844
rect 2723 1840 2724 1844
rect 2718 1839 2724 1840
rect 2886 1844 2892 1845
rect 2886 1840 2887 1844
rect 2891 1840 2892 1844
rect 2886 1839 2892 1840
rect 3038 1844 3044 1845
rect 3038 1840 3039 1844
rect 3043 1840 3044 1844
rect 3038 1839 3044 1840
rect 3182 1844 3188 1845
rect 3182 1840 3183 1844
rect 3187 1840 3188 1844
rect 3182 1839 3188 1840
rect 3318 1844 3324 1845
rect 3318 1840 3319 1844
rect 3323 1840 3324 1844
rect 3318 1839 3324 1840
rect 3454 1844 3460 1845
rect 3454 1840 3455 1844
rect 3459 1840 3460 1844
rect 3454 1839 3460 1840
rect 3582 1844 3588 1845
rect 3582 1840 3583 1844
rect 3587 1840 3588 1844
rect 3582 1839 3588 1840
rect 3710 1844 3716 1845
rect 3710 1840 3711 1844
rect 3715 1840 3716 1844
rect 3710 1839 3716 1840
rect 3838 1844 3844 1845
rect 3838 1840 3839 1844
rect 3843 1840 3844 1844
rect 3944 1842 3946 1869
rect 3838 1839 3844 1840
rect 3942 1841 3948 1842
rect 2046 1836 2052 1837
rect 3942 1837 3943 1841
rect 3947 1837 3948 1841
rect 3942 1836 3948 1837
rect 111 1834 115 1835
rect 111 1829 115 1830
rect 511 1834 515 1835
rect 511 1829 515 1830
rect 615 1834 619 1835
rect 615 1829 619 1830
rect 623 1834 627 1835
rect 623 1829 627 1830
rect 711 1834 715 1835
rect 711 1829 715 1830
rect 743 1834 747 1835
rect 743 1829 747 1830
rect 815 1834 819 1835
rect 815 1829 819 1830
rect 863 1834 867 1835
rect 863 1829 867 1830
rect 927 1834 931 1835
rect 927 1829 931 1830
rect 983 1834 987 1835
rect 983 1829 987 1830
rect 1039 1834 1043 1835
rect 1039 1829 1043 1830
rect 1103 1834 1107 1835
rect 1103 1829 1107 1830
rect 1159 1834 1163 1835
rect 1159 1829 1163 1830
rect 1223 1834 1227 1835
rect 1223 1829 1227 1830
rect 1279 1834 1283 1835
rect 1279 1829 1283 1830
rect 1335 1834 1339 1835
rect 1335 1829 1339 1830
rect 1399 1834 1403 1835
rect 1399 1829 1403 1830
rect 1455 1834 1459 1835
rect 1455 1829 1459 1830
rect 1519 1834 1523 1835
rect 1519 1829 1523 1830
rect 1575 1834 1579 1835
rect 1575 1829 1579 1830
rect 1639 1834 1643 1835
rect 1639 1829 1643 1830
rect 1695 1834 1699 1835
rect 1695 1829 1699 1830
rect 2007 1834 2011 1835
rect 2007 1829 2011 1830
rect 112 1802 114 1829
rect 616 1805 618 1829
rect 712 1805 714 1829
rect 816 1805 818 1829
rect 928 1805 930 1829
rect 1040 1805 1042 1829
rect 1160 1805 1162 1829
rect 1280 1805 1282 1829
rect 1400 1805 1402 1829
rect 1520 1805 1522 1829
rect 1640 1805 1642 1829
rect 614 1804 620 1805
rect 110 1801 116 1802
rect 110 1797 111 1801
rect 115 1797 116 1801
rect 614 1800 615 1804
rect 619 1800 620 1804
rect 614 1799 620 1800
rect 710 1804 716 1805
rect 710 1800 711 1804
rect 715 1800 716 1804
rect 710 1799 716 1800
rect 814 1804 820 1805
rect 814 1800 815 1804
rect 819 1800 820 1804
rect 814 1799 820 1800
rect 926 1804 932 1805
rect 926 1800 927 1804
rect 931 1800 932 1804
rect 926 1799 932 1800
rect 1038 1804 1044 1805
rect 1038 1800 1039 1804
rect 1043 1800 1044 1804
rect 1038 1799 1044 1800
rect 1158 1804 1164 1805
rect 1158 1800 1159 1804
rect 1163 1800 1164 1804
rect 1158 1799 1164 1800
rect 1278 1804 1284 1805
rect 1278 1800 1279 1804
rect 1283 1800 1284 1804
rect 1278 1799 1284 1800
rect 1398 1804 1404 1805
rect 1398 1800 1399 1804
rect 1403 1800 1404 1804
rect 1398 1799 1404 1800
rect 1518 1804 1524 1805
rect 1518 1800 1519 1804
rect 1523 1800 1524 1804
rect 1518 1799 1524 1800
rect 1638 1804 1644 1805
rect 1638 1800 1639 1804
rect 1643 1800 1644 1804
rect 2008 1802 2010 1829
rect 2070 1825 2076 1826
rect 2046 1824 2052 1825
rect 2046 1820 2047 1824
rect 2051 1820 2052 1824
rect 2070 1821 2071 1825
rect 2075 1821 2076 1825
rect 2070 1820 2076 1821
rect 2198 1825 2204 1826
rect 2198 1821 2199 1825
rect 2203 1821 2204 1825
rect 2198 1820 2204 1821
rect 2366 1825 2372 1826
rect 2366 1821 2367 1825
rect 2371 1821 2372 1825
rect 2366 1820 2372 1821
rect 2542 1825 2548 1826
rect 2542 1821 2543 1825
rect 2547 1821 2548 1825
rect 2542 1820 2548 1821
rect 2718 1825 2724 1826
rect 2718 1821 2719 1825
rect 2723 1821 2724 1825
rect 2718 1820 2724 1821
rect 2886 1825 2892 1826
rect 2886 1821 2887 1825
rect 2891 1821 2892 1825
rect 2886 1820 2892 1821
rect 3038 1825 3044 1826
rect 3038 1821 3039 1825
rect 3043 1821 3044 1825
rect 3038 1820 3044 1821
rect 3182 1825 3188 1826
rect 3182 1821 3183 1825
rect 3187 1821 3188 1825
rect 3182 1820 3188 1821
rect 3318 1825 3324 1826
rect 3318 1821 3319 1825
rect 3323 1821 3324 1825
rect 3318 1820 3324 1821
rect 3454 1825 3460 1826
rect 3454 1821 3455 1825
rect 3459 1821 3460 1825
rect 3454 1820 3460 1821
rect 3582 1825 3588 1826
rect 3582 1821 3583 1825
rect 3587 1821 3588 1825
rect 3582 1820 3588 1821
rect 3710 1825 3716 1826
rect 3710 1821 3711 1825
rect 3715 1821 3716 1825
rect 3710 1820 3716 1821
rect 3838 1825 3844 1826
rect 3838 1821 3839 1825
rect 3843 1821 3844 1825
rect 3838 1820 3844 1821
rect 3942 1824 3948 1825
rect 3942 1820 3943 1824
rect 3947 1820 3948 1824
rect 2046 1819 2052 1820
rect 1638 1799 1644 1800
rect 2006 1801 2012 1802
rect 110 1796 116 1797
rect 2006 1797 2007 1801
rect 2011 1797 2012 1801
rect 2006 1796 2012 1797
rect 2048 1795 2050 1819
rect 2072 1795 2074 1820
rect 2200 1795 2202 1820
rect 2368 1795 2370 1820
rect 2544 1795 2546 1820
rect 2720 1795 2722 1820
rect 2888 1795 2890 1820
rect 3040 1795 3042 1820
rect 3184 1795 3186 1820
rect 3320 1795 3322 1820
rect 3456 1795 3458 1820
rect 3584 1795 3586 1820
rect 3712 1795 3714 1820
rect 3840 1795 3842 1820
rect 3942 1819 3948 1820
rect 3944 1795 3946 1819
rect 2047 1794 2051 1795
rect 2047 1789 2051 1790
rect 2071 1794 2075 1795
rect 2071 1789 2075 1790
rect 2183 1794 2187 1795
rect 2183 1789 2187 1790
rect 2199 1794 2203 1795
rect 2199 1789 2203 1790
rect 2327 1794 2331 1795
rect 2327 1789 2331 1790
rect 2367 1794 2371 1795
rect 2367 1789 2371 1790
rect 2487 1794 2491 1795
rect 2487 1789 2491 1790
rect 2543 1794 2547 1795
rect 2543 1789 2547 1790
rect 2655 1794 2659 1795
rect 2655 1789 2659 1790
rect 2719 1794 2723 1795
rect 2719 1789 2723 1790
rect 2831 1794 2835 1795
rect 2831 1789 2835 1790
rect 2887 1794 2891 1795
rect 2887 1789 2891 1790
rect 3023 1794 3027 1795
rect 3023 1789 3027 1790
rect 3039 1794 3043 1795
rect 3039 1789 3043 1790
rect 3183 1794 3187 1795
rect 3183 1789 3187 1790
rect 3223 1794 3227 1795
rect 3223 1789 3227 1790
rect 3319 1794 3323 1795
rect 3319 1789 3323 1790
rect 3431 1794 3435 1795
rect 3431 1789 3435 1790
rect 3455 1794 3459 1795
rect 3455 1789 3459 1790
rect 3583 1794 3587 1795
rect 3583 1789 3587 1790
rect 3647 1794 3651 1795
rect 3647 1789 3651 1790
rect 3711 1794 3715 1795
rect 3711 1789 3715 1790
rect 3839 1794 3843 1795
rect 3839 1789 3843 1790
rect 3943 1794 3947 1795
rect 3943 1789 3947 1790
rect 614 1785 620 1786
rect 110 1784 116 1785
rect 110 1780 111 1784
rect 115 1780 116 1784
rect 614 1781 615 1785
rect 619 1781 620 1785
rect 614 1780 620 1781
rect 710 1785 716 1786
rect 710 1781 711 1785
rect 715 1781 716 1785
rect 710 1780 716 1781
rect 814 1785 820 1786
rect 814 1781 815 1785
rect 819 1781 820 1785
rect 814 1780 820 1781
rect 926 1785 932 1786
rect 926 1781 927 1785
rect 931 1781 932 1785
rect 926 1780 932 1781
rect 1038 1785 1044 1786
rect 1038 1781 1039 1785
rect 1043 1781 1044 1785
rect 1038 1780 1044 1781
rect 1158 1785 1164 1786
rect 1158 1781 1159 1785
rect 1163 1781 1164 1785
rect 1158 1780 1164 1781
rect 1278 1785 1284 1786
rect 1278 1781 1279 1785
rect 1283 1781 1284 1785
rect 1278 1780 1284 1781
rect 1398 1785 1404 1786
rect 1398 1781 1399 1785
rect 1403 1781 1404 1785
rect 1398 1780 1404 1781
rect 1518 1785 1524 1786
rect 1518 1781 1519 1785
rect 1523 1781 1524 1785
rect 1518 1780 1524 1781
rect 1638 1785 1644 1786
rect 1638 1781 1639 1785
rect 1643 1781 1644 1785
rect 1638 1780 1644 1781
rect 2006 1784 2012 1785
rect 2006 1780 2007 1784
rect 2011 1780 2012 1784
rect 110 1779 116 1780
rect 112 1759 114 1779
rect 616 1759 618 1780
rect 712 1759 714 1780
rect 816 1759 818 1780
rect 928 1759 930 1780
rect 1040 1759 1042 1780
rect 1160 1759 1162 1780
rect 1280 1759 1282 1780
rect 1400 1759 1402 1780
rect 1520 1759 1522 1780
rect 1640 1759 1642 1780
rect 2006 1779 2012 1780
rect 2008 1759 2010 1779
rect 2048 1769 2050 1789
rect 2046 1768 2052 1769
rect 2072 1768 2074 1789
rect 2184 1768 2186 1789
rect 2328 1768 2330 1789
rect 2488 1768 2490 1789
rect 2656 1768 2658 1789
rect 2832 1768 2834 1789
rect 3024 1768 3026 1789
rect 3224 1768 3226 1789
rect 3432 1768 3434 1789
rect 3648 1768 3650 1789
rect 3840 1768 3842 1789
rect 3944 1769 3946 1789
rect 3942 1768 3948 1769
rect 2046 1764 2047 1768
rect 2051 1764 2052 1768
rect 2046 1763 2052 1764
rect 2070 1767 2076 1768
rect 2070 1763 2071 1767
rect 2075 1763 2076 1767
rect 2070 1762 2076 1763
rect 2182 1767 2188 1768
rect 2182 1763 2183 1767
rect 2187 1763 2188 1767
rect 2182 1762 2188 1763
rect 2326 1767 2332 1768
rect 2326 1763 2327 1767
rect 2331 1763 2332 1767
rect 2326 1762 2332 1763
rect 2486 1767 2492 1768
rect 2486 1763 2487 1767
rect 2491 1763 2492 1767
rect 2486 1762 2492 1763
rect 2654 1767 2660 1768
rect 2654 1763 2655 1767
rect 2659 1763 2660 1767
rect 2654 1762 2660 1763
rect 2830 1767 2836 1768
rect 2830 1763 2831 1767
rect 2835 1763 2836 1767
rect 2830 1762 2836 1763
rect 3022 1767 3028 1768
rect 3022 1763 3023 1767
rect 3027 1763 3028 1767
rect 3022 1762 3028 1763
rect 3222 1767 3228 1768
rect 3222 1763 3223 1767
rect 3227 1763 3228 1767
rect 3222 1762 3228 1763
rect 3430 1767 3436 1768
rect 3430 1763 3431 1767
rect 3435 1763 3436 1767
rect 3430 1762 3436 1763
rect 3646 1767 3652 1768
rect 3646 1763 3647 1767
rect 3651 1763 3652 1767
rect 3646 1762 3652 1763
rect 3838 1767 3844 1768
rect 3838 1763 3839 1767
rect 3843 1763 3844 1767
rect 3942 1764 3943 1768
rect 3947 1764 3948 1768
rect 3942 1763 3948 1764
rect 3838 1762 3844 1763
rect 111 1758 115 1759
rect 111 1753 115 1754
rect 367 1758 371 1759
rect 367 1753 371 1754
rect 495 1758 499 1759
rect 495 1753 499 1754
rect 615 1758 619 1759
rect 615 1753 619 1754
rect 639 1758 643 1759
rect 639 1753 643 1754
rect 711 1758 715 1759
rect 711 1753 715 1754
rect 799 1758 803 1759
rect 799 1753 803 1754
rect 815 1758 819 1759
rect 815 1753 819 1754
rect 927 1758 931 1759
rect 927 1753 931 1754
rect 967 1758 971 1759
rect 967 1753 971 1754
rect 1039 1758 1043 1759
rect 1039 1753 1043 1754
rect 1143 1758 1147 1759
rect 1143 1753 1147 1754
rect 1159 1758 1163 1759
rect 1159 1753 1163 1754
rect 1279 1758 1283 1759
rect 1279 1753 1283 1754
rect 1327 1758 1331 1759
rect 1327 1753 1331 1754
rect 1399 1758 1403 1759
rect 1399 1753 1403 1754
rect 1511 1758 1515 1759
rect 1511 1753 1515 1754
rect 1519 1758 1523 1759
rect 1519 1753 1523 1754
rect 1639 1758 1643 1759
rect 1639 1753 1643 1754
rect 1703 1758 1707 1759
rect 1703 1753 1707 1754
rect 2007 1758 2011 1759
rect 2007 1753 2011 1754
rect 112 1733 114 1753
rect 110 1732 116 1733
rect 368 1732 370 1753
rect 496 1732 498 1753
rect 640 1732 642 1753
rect 800 1732 802 1753
rect 968 1732 970 1753
rect 1144 1732 1146 1753
rect 1328 1732 1330 1753
rect 1512 1732 1514 1753
rect 1704 1732 1706 1753
rect 2008 1733 2010 1753
rect 2046 1751 2052 1752
rect 2046 1747 2047 1751
rect 2051 1747 2052 1751
rect 3942 1751 3948 1752
rect 2046 1746 2052 1747
rect 2070 1748 2076 1749
rect 2006 1732 2012 1733
rect 110 1728 111 1732
rect 115 1728 116 1732
rect 110 1727 116 1728
rect 366 1731 372 1732
rect 366 1727 367 1731
rect 371 1727 372 1731
rect 366 1726 372 1727
rect 494 1731 500 1732
rect 494 1727 495 1731
rect 499 1727 500 1731
rect 494 1726 500 1727
rect 638 1731 644 1732
rect 638 1727 639 1731
rect 643 1727 644 1731
rect 638 1726 644 1727
rect 798 1731 804 1732
rect 798 1727 799 1731
rect 803 1727 804 1731
rect 798 1726 804 1727
rect 966 1731 972 1732
rect 966 1727 967 1731
rect 971 1727 972 1731
rect 966 1726 972 1727
rect 1142 1731 1148 1732
rect 1142 1727 1143 1731
rect 1147 1727 1148 1731
rect 1142 1726 1148 1727
rect 1326 1731 1332 1732
rect 1326 1727 1327 1731
rect 1331 1727 1332 1731
rect 1326 1726 1332 1727
rect 1510 1731 1516 1732
rect 1510 1727 1511 1731
rect 1515 1727 1516 1731
rect 1510 1726 1516 1727
rect 1702 1731 1708 1732
rect 1702 1727 1703 1731
rect 1707 1727 1708 1731
rect 2006 1728 2007 1732
rect 2011 1728 2012 1732
rect 2006 1727 2012 1728
rect 1702 1726 1708 1727
rect 110 1715 116 1716
rect 110 1711 111 1715
rect 115 1711 116 1715
rect 2006 1715 2012 1716
rect 110 1710 116 1711
rect 366 1712 372 1713
rect 112 1679 114 1710
rect 366 1708 367 1712
rect 371 1708 372 1712
rect 366 1707 372 1708
rect 494 1712 500 1713
rect 494 1708 495 1712
rect 499 1708 500 1712
rect 494 1707 500 1708
rect 638 1712 644 1713
rect 638 1708 639 1712
rect 643 1708 644 1712
rect 638 1707 644 1708
rect 798 1712 804 1713
rect 798 1708 799 1712
rect 803 1708 804 1712
rect 798 1707 804 1708
rect 966 1712 972 1713
rect 966 1708 967 1712
rect 971 1708 972 1712
rect 966 1707 972 1708
rect 1142 1712 1148 1713
rect 1142 1708 1143 1712
rect 1147 1708 1148 1712
rect 1142 1707 1148 1708
rect 1326 1712 1332 1713
rect 1326 1708 1327 1712
rect 1331 1708 1332 1712
rect 1326 1707 1332 1708
rect 1510 1712 1516 1713
rect 1510 1708 1511 1712
rect 1515 1708 1516 1712
rect 1510 1707 1516 1708
rect 1702 1712 1708 1713
rect 1702 1708 1703 1712
rect 1707 1708 1708 1712
rect 2006 1711 2007 1715
rect 2011 1711 2012 1715
rect 2048 1711 2050 1746
rect 2070 1744 2071 1748
rect 2075 1744 2076 1748
rect 2070 1743 2076 1744
rect 2182 1748 2188 1749
rect 2182 1744 2183 1748
rect 2187 1744 2188 1748
rect 2182 1743 2188 1744
rect 2326 1748 2332 1749
rect 2326 1744 2327 1748
rect 2331 1744 2332 1748
rect 2326 1743 2332 1744
rect 2486 1748 2492 1749
rect 2486 1744 2487 1748
rect 2491 1744 2492 1748
rect 2486 1743 2492 1744
rect 2654 1748 2660 1749
rect 2654 1744 2655 1748
rect 2659 1744 2660 1748
rect 2654 1743 2660 1744
rect 2830 1748 2836 1749
rect 2830 1744 2831 1748
rect 2835 1744 2836 1748
rect 2830 1743 2836 1744
rect 3022 1748 3028 1749
rect 3022 1744 3023 1748
rect 3027 1744 3028 1748
rect 3022 1743 3028 1744
rect 3222 1748 3228 1749
rect 3222 1744 3223 1748
rect 3227 1744 3228 1748
rect 3222 1743 3228 1744
rect 3430 1748 3436 1749
rect 3430 1744 3431 1748
rect 3435 1744 3436 1748
rect 3430 1743 3436 1744
rect 3646 1748 3652 1749
rect 3646 1744 3647 1748
rect 3651 1744 3652 1748
rect 3646 1743 3652 1744
rect 3838 1748 3844 1749
rect 3838 1744 3839 1748
rect 3843 1744 3844 1748
rect 3942 1747 3943 1751
rect 3947 1747 3948 1751
rect 3942 1746 3948 1747
rect 3838 1743 3844 1744
rect 2072 1711 2074 1743
rect 2184 1711 2186 1743
rect 2328 1711 2330 1743
rect 2488 1711 2490 1743
rect 2656 1711 2658 1743
rect 2832 1711 2834 1743
rect 3024 1711 3026 1743
rect 3224 1711 3226 1743
rect 3432 1711 3434 1743
rect 3648 1711 3650 1743
rect 3840 1711 3842 1743
rect 3944 1711 3946 1746
rect 2006 1710 2012 1711
rect 2047 1710 2051 1711
rect 1702 1707 1708 1708
rect 368 1679 370 1707
rect 496 1679 498 1707
rect 640 1679 642 1707
rect 800 1679 802 1707
rect 968 1679 970 1707
rect 1144 1679 1146 1707
rect 1328 1679 1330 1707
rect 1512 1679 1514 1707
rect 1704 1679 1706 1707
rect 2008 1679 2010 1710
rect 2047 1705 2051 1706
rect 2071 1710 2075 1711
rect 2071 1705 2075 1706
rect 2183 1710 2187 1711
rect 2183 1705 2187 1706
rect 2223 1710 2227 1711
rect 2223 1705 2227 1706
rect 2327 1710 2331 1711
rect 2327 1705 2331 1706
rect 2439 1710 2443 1711
rect 2439 1705 2443 1706
rect 2487 1710 2491 1711
rect 2487 1705 2491 1706
rect 2559 1710 2563 1711
rect 2559 1705 2563 1706
rect 2655 1710 2659 1711
rect 2655 1705 2659 1706
rect 2687 1710 2691 1711
rect 2687 1705 2691 1706
rect 2823 1710 2827 1711
rect 2823 1705 2827 1706
rect 2831 1710 2835 1711
rect 2831 1705 2835 1706
rect 2967 1710 2971 1711
rect 2967 1705 2971 1706
rect 3023 1710 3027 1711
rect 3023 1705 3027 1706
rect 3127 1710 3131 1711
rect 3127 1705 3131 1706
rect 3223 1710 3227 1711
rect 3223 1705 3227 1706
rect 3303 1710 3307 1711
rect 3303 1705 3307 1706
rect 3431 1710 3435 1711
rect 3431 1705 3435 1706
rect 3487 1710 3491 1711
rect 3487 1705 3491 1706
rect 3647 1710 3651 1711
rect 3647 1705 3651 1706
rect 3671 1710 3675 1711
rect 3671 1705 3675 1706
rect 3839 1710 3843 1711
rect 3839 1705 3843 1706
rect 3943 1710 3947 1711
rect 3943 1705 3947 1706
rect 111 1678 115 1679
rect 111 1673 115 1674
rect 135 1678 139 1679
rect 135 1673 139 1674
rect 247 1678 251 1679
rect 247 1673 251 1674
rect 367 1678 371 1679
rect 367 1673 371 1674
rect 399 1678 403 1679
rect 399 1673 403 1674
rect 495 1678 499 1679
rect 495 1673 499 1674
rect 567 1678 571 1679
rect 567 1673 571 1674
rect 639 1678 643 1679
rect 639 1673 643 1674
rect 743 1678 747 1679
rect 743 1673 747 1674
rect 799 1678 803 1679
rect 799 1673 803 1674
rect 935 1678 939 1679
rect 935 1673 939 1674
rect 967 1678 971 1679
rect 967 1673 971 1674
rect 1135 1678 1139 1679
rect 1135 1673 1139 1674
rect 1143 1678 1147 1679
rect 1143 1673 1147 1674
rect 1327 1678 1331 1679
rect 1327 1673 1331 1674
rect 1343 1678 1347 1679
rect 1343 1673 1347 1674
rect 1511 1678 1515 1679
rect 1511 1673 1515 1674
rect 1551 1678 1555 1679
rect 1551 1673 1555 1674
rect 1703 1678 1707 1679
rect 1703 1673 1707 1674
rect 1767 1678 1771 1679
rect 1767 1673 1771 1674
rect 2007 1678 2011 1679
rect 2048 1678 2050 1705
rect 2224 1681 2226 1705
rect 2328 1681 2330 1705
rect 2440 1681 2442 1705
rect 2560 1681 2562 1705
rect 2688 1681 2690 1705
rect 2824 1681 2826 1705
rect 2968 1681 2970 1705
rect 3128 1681 3130 1705
rect 3304 1681 3306 1705
rect 3488 1681 3490 1705
rect 3672 1681 3674 1705
rect 3840 1681 3842 1705
rect 2222 1680 2228 1681
rect 2007 1673 2011 1674
rect 2046 1677 2052 1678
rect 2046 1673 2047 1677
rect 2051 1673 2052 1677
rect 2222 1676 2223 1680
rect 2227 1676 2228 1680
rect 2222 1675 2228 1676
rect 2326 1680 2332 1681
rect 2326 1676 2327 1680
rect 2331 1676 2332 1680
rect 2326 1675 2332 1676
rect 2438 1680 2444 1681
rect 2438 1676 2439 1680
rect 2443 1676 2444 1680
rect 2438 1675 2444 1676
rect 2558 1680 2564 1681
rect 2558 1676 2559 1680
rect 2563 1676 2564 1680
rect 2558 1675 2564 1676
rect 2686 1680 2692 1681
rect 2686 1676 2687 1680
rect 2691 1676 2692 1680
rect 2686 1675 2692 1676
rect 2822 1680 2828 1681
rect 2822 1676 2823 1680
rect 2827 1676 2828 1680
rect 2822 1675 2828 1676
rect 2966 1680 2972 1681
rect 2966 1676 2967 1680
rect 2971 1676 2972 1680
rect 2966 1675 2972 1676
rect 3126 1680 3132 1681
rect 3126 1676 3127 1680
rect 3131 1676 3132 1680
rect 3126 1675 3132 1676
rect 3302 1680 3308 1681
rect 3302 1676 3303 1680
rect 3307 1676 3308 1680
rect 3302 1675 3308 1676
rect 3486 1680 3492 1681
rect 3486 1676 3487 1680
rect 3491 1676 3492 1680
rect 3486 1675 3492 1676
rect 3670 1680 3676 1681
rect 3670 1676 3671 1680
rect 3675 1676 3676 1680
rect 3670 1675 3676 1676
rect 3838 1680 3844 1681
rect 3838 1676 3839 1680
rect 3843 1676 3844 1680
rect 3944 1678 3946 1705
rect 3838 1675 3844 1676
rect 3942 1677 3948 1678
rect 112 1646 114 1673
rect 136 1649 138 1673
rect 248 1649 250 1673
rect 400 1649 402 1673
rect 568 1649 570 1673
rect 744 1649 746 1673
rect 936 1649 938 1673
rect 1136 1649 1138 1673
rect 1344 1649 1346 1673
rect 1552 1649 1554 1673
rect 1768 1649 1770 1673
rect 134 1648 140 1649
rect 110 1645 116 1646
rect 110 1641 111 1645
rect 115 1641 116 1645
rect 134 1644 135 1648
rect 139 1644 140 1648
rect 134 1643 140 1644
rect 246 1648 252 1649
rect 246 1644 247 1648
rect 251 1644 252 1648
rect 246 1643 252 1644
rect 398 1648 404 1649
rect 398 1644 399 1648
rect 403 1644 404 1648
rect 398 1643 404 1644
rect 566 1648 572 1649
rect 566 1644 567 1648
rect 571 1644 572 1648
rect 566 1643 572 1644
rect 742 1648 748 1649
rect 742 1644 743 1648
rect 747 1644 748 1648
rect 742 1643 748 1644
rect 934 1648 940 1649
rect 934 1644 935 1648
rect 939 1644 940 1648
rect 934 1643 940 1644
rect 1134 1648 1140 1649
rect 1134 1644 1135 1648
rect 1139 1644 1140 1648
rect 1134 1643 1140 1644
rect 1342 1648 1348 1649
rect 1342 1644 1343 1648
rect 1347 1644 1348 1648
rect 1342 1643 1348 1644
rect 1550 1648 1556 1649
rect 1550 1644 1551 1648
rect 1555 1644 1556 1648
rect 1550 1643 1556 1644
rect 1766 1648 1772 1649
rect 1766 1644 1767 1648
rect 1771 1644 1772 1648
rect 2008 1646 2010 1673
rect 2046 1672 2052 1673
rect 3942 1673 3943 1677
rect 3947 1673 3948 1677
rect 3942 1672 3948 1673
rect 2222 1661 2228 1662
rect 2046 1660 2052 1661
rect 2046 1656 2047 1660
rect 2051 1656 2052 1660
rect 2222 1657 2223 1661
rect 2227 1657 2228 1661
rect 2222 1656 2228 1657
rect 2326 1661 2332 1662
rect 2326 1657 2327 1661
rect 2331 1657 2332 1661
rect 2326 1656 2332 1657
rect 2438 1661 2444 1662
rect 2438 1657 2439 1661
rect 2443 1657 2444 1661
rect 2438 1656 2444 1657
rect 2558 1661 2564 1662
rect 2558 1657 2559 1661
rect 2563 1657 2564 1661
rect 2558 1656 2564 1657
rect 2686 1661 2692 1662
rect 2686 1657 2687 1661
rect 2691 1657 2692 1661
rect 2686 1656 2692 1657
rect 2822 1661 2828 1662
rect 2822 1657 2823 1661
rect 2827 1657 2828 1661
rect 2822 1656 2828 1657
rect 2966 1661 2972 1662
rect 2966 1657 2967 1661
rect 2971 1657 2972 1661
rect 2966 1656 2972 1657
rect 3126 1661 3132 1662
rect 3126 1657 3127 1661
rect 3131 1657 3132 1661
rect 3126 1656 3132 1657
rect 3302 1661 3308 1662
rect 3302 1657 3303 1661
rect 3307 1657 3308 1661
rect 3302 1656 3308 1657
rect 3486 1661 3492 1662
rect 3486 1657 3487 1661
rect 3491 1657 3492 1661
rect 3486 1656 3492 1657
rect 3670 1661 3676 1662
rect 3670 1657 3671 1661
rect 3675 1657 3676 1661
rect 3670 1656 3676 1657
rect 3838 1661 3844 1662
rect 3838 1657 3839 1661
rect 3843 1657 3844 1661
rect 3838 1656 3844 1657
rect 3942 1660 3948 1661
rect 3942 1656 3943 1660
rect 3947 1656 3948 1660
rect 2046 1655 2052 1656
rect 1766 1643 1772 1644
rect 2006 1645 2012 1646
rect 110 1640 116 1641
rect 2006 1641 2007 1645
rect 2011 1641 2012 1645
rect 2006 1640 2012 1641
rect 2048 1631 2050 1655
rect 2224 1631 2226 1656
rect 2328 1631 2330 1656
rect 2440 1631 2442 1656
rect 2560 1631 2562 1656
rect 2688 1631 2690 1656
rect 2824 1631 2826 1656
rect 2968 1631 2970 1656
rect 3128 1631 3130 1656
rect 3304 1631 3306 1656
rect 3488 1631 3490 1656
rect 3672 1631 3674 1656
rect 3840 1631 3842 1656
rect 3942 1655 3948 1656
rect 3944 1631 3946 1655
rect 2047 1630 2051 1631
rect 134 1629 140 1630
rect 110 1628 116 1629
rect 110 1624 111 1628
rect 115 1624 116 1628
rect 134 1625 135 1629
rect 139 1625 140 1629
rect 134 1624 140 1625
rect 246 1629 252 1630
rect 246 1625 247 1629
rect 251 1625 252 1629
rect 246 1624 252 1625
rect 398 1629 404 1630
rect 398 1625 399 1629
rect 403 1625 404 1629
rect 398 1624 404 1625
rect 566 1629 572 1630
rect 566 1625 567 1629
rect 571 1625 572 1629
rect 566 1624 572 1625
rect 742 1629 748 1630
rect 742 1625 743 1629
rect 747 1625 748 1629
rect 742 1624 748 1625
rect 934 1629 940 1630
rect 934 1625 935 1629
rect 939 1625 940 1629
rect 934 1624 940 1625
rect 1134 1629 1140 1630
rect 1134 1625 1135 1629
rect 1139 1625 1140 1629
rect 1134 1624 1140 1625
rect 1342 1629 1348 1630
rect 1342 1625 1343 1629
rect 1347 1625 1348 1629
rect 1342 1624 1348 1625
rect 1550 1629 1556 1630
rect 1550 1625 1551 1629
rect 1555 1625 1556 1629
rect 1550 1624 1556 1625
rect 1766 1629 1772 1630
rect 1766 1625 1767 1629
rect 1771 1625 1772 1629
rect 1766 1624 1772 1625
rect 2006 1628 2012 1629
rect 2006 1624 2007 1628
rect 2011 1624 2012 1628
rect 2047 1625 2051 1626
rect 2223 1630 2227 1631
rect 2223 1625 2227 1626
rect 2327 1630 2331 1631
rect 2327 1625 2331 1626
rect 2391 1630 2395 1631
rect 2391 1625 2395 1626
rect 2439 1630 2443 1631
rect 2439 1625 2443 1626
rect 2503 1630 2507 1631
rect 2503 1625 2507 1626
rect 2559 1630 2563 1631
rect 2559 1625 2563 1626
rect 2615 1630 2619 1631
rect 2615 1625 2619 1626
rect 2687 1630 2691 1631
rect 2687 1625 2691 1626
rect 2735 1630 2739 1631
rect 2735 1625 2739 1626
rect 2823 1630 2827 1631
rect 2823 1625 2827 1626
rect 2855 1630 2859 1631
rect 2855 1625 2859 1626
rect 2967 1630 2971 1631
rect 2967 1625 2971 1626
rect 2975 1630 2979 1631
rect 2975 1625 2979 1626
rect 3095 1630 3099 1631
rect 3095 1625 3099 1626
rect 3127 1630 3131 1631
rect 3127 1625 3131 1626
rect 3215 1630 3219 1631
rect 3215 1625 3219 1626
rect 3303 1630 3307 1631
rect 3303 1625 3307 1626
rect 3335 1630 3339 1631
rect 3335 1625 3339 1626
rect 3455 1630 3459 1631
rect 3455 1625 3459 1626
rect 3487 1630 3491 1631
rect 3487 1625 3491 1626
rect 3671 1630 3675 1631
rect 3671 1625 3675 1626
rect 3839 1630 3843 1631
rect 3839 1625 3843 1626
rect 3943 1630 3947 1631
rect 3943 1625 3947 1626
rect 110 1623 116 1624
rect 112 1599 114 1623
rect 136 1599 138 1624
rect 248 1599 250 1624
rect 400 1599 402 1624
rect 568 1599 570 1624
rect 744 1599 746 1624
rect 936 1599 938 1624
rect 1136 1599 1138 1624
rect 1344 1599 1346 1624
rect 1552 1599 1554 1624
rect 1768 1599 1770 1624
rect 2006 1623 2012 1624
rect 2008 1599 2010 1623
rect 2048 1605 2050 1625
rect 2046 1604 2052 1605
rect 2392 1604 2394 1625
rect 2504 1604 2506 1625
rect 2616 1604 2618 1625
rect 2736 1604 2738 1625
rect 2856 1604 2858 1625
rect 2976 1604 2978 1625
rect 3096 1604 3098 1625
rect 3216 1604 3218 1625
rect 3336 1604 3338 1625
rect 3456 1604 3458 1625
rect 3944 1605 3946 1625
rect 3942 1604 3948 1605
rect 2046 1600 2047 1604
rect 2051 1600 2052 1604
rect 2046 1599 2052 1600
rect 2390 1603 2396 1604
rect 2390 1599 2391 1603
rect 2395 1599 2396 1603
rect 111 1598 115 1599
rect 111 1593 115 1594
rect 135 1598 139 1599
rect 135 1593 139 1594
rect 247 1598 251 1599
rect 247 1593 251 1594
rect 255 1598 259 1599
rect 255 1593 259 1594
rect 399 1598 403 1599
rect 399 1593 403 1594
rect 423 1598 427 1599
rect 423 1593 427 1594
rect 567 1598 571 1599
rect 567 1593 571 1594
rect 615 1598 619 1599
rect 615 1593 619 1594
rect 743 1598 747 1599
rect 743 1593 747 1594
rect 831 1598 835 1599
rect 831 1593 835 1594
rect 935 1598 939 1599
rect 935 1593 939 1594
rect 1063 1598 1067 1599
rect 1063 1593 1067 1594
rect 1135 1598 1139 1599
rect 1135 1593 1139 1594
rect 1311 1598 1315 1599
rect 1311 1593 1315 1594
rect 1343 1598 1347 1599
rect 1343 1593 1347 1594
rect 1551 1598 1555 1599
rect 1551 1593 1555 1594
rect 1567 1598 1571 1599
rect 1567 1593 1571 1594
rect 1767 1598 1771 1599
rect 1767 1593 1771 1594
rect 1831 1598 1835 1599
rect 1831 1593 1835 1594
rect 2007 1598 2011 1599
rect 2390 1598 2396 1599
rect 2502 1603 2508 1604
rect 2502 1599 2503 1603
rect 2507 1599 2508 1603
rect 2502 1598 2508 1599
rect 2614 1603 2620 1604
rect 2614 1599 2615 1603
rect 2619 1599 2620 1603
rect 2614 1598 2620 1599
rect 2734 1603 2740 1604
rect 2734 1599 2735 1603
rect 2739 1599 2740 1603
rect 2734 1598 2740 1599
rect 2854 1603 2860 1604
rect 2854 1599 2855 1603
rect 2859 1599 2860 1603
rect 2854 1598 2860 1599
rect 2974 1603 2980 1604
rect 2974 1599 2975 1603
rect 2979 1599 2980 1603
rect 2974 1598 2980 1599
rect 3094 1603 3100 1604
rect 3094 1599 3095 1603
rect 3099 1599 3100 1603
rect 3094 1598 3100 1599
rect 3214 1603 3220 1604
rect 3214 1599 3215 1603
rect 3219 1599 3220 1603
rect 3214 1598 3220 1599
rect 3334 1603 3340 1604
rect 3334 1599 3335 1603
rect 3339 1599 3340 1603
rect 3334 1598 3340 1599
rect 3454 1603 3460 1604
rect 3454 1599 3455 1603
rect 3459 1599 3460 1603
rect 3942 1600 3943 1604
rect 3947 1600 3948 1604
rect 3942 1599 3948 1600
rect 3454 1598 3460 1599
rect 2007 1593 2011 1594
rect 112 1573 114 1593
rect 110 1572 116 1573
rect 136 1572 138 1593
rect 256 1572 258 1593
rect 424 1572 426 1593
rect 616 1572 618 1593
rect 832 1572 834 1593
rect 1064 1572 1066 1593
rect 1312 1572 1314 1593
rect 1568 1572 1570 1593
rect 1832 1572 1834 1593
rect 2008 1573 2010 1593
rect 2046 1587 2052 1588
rect 2046 1583 2047 1587
rect 2051 1583 2052 1587
rect 3942 1587 3948 1588
rect 2046 1582 2052 1583
rect 2390 1584 2396 1585
rect 2006 1572 2012 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 110 1567 116 1568
rect 134 1571 140 1572
rect 134 1567 135 1571
rect 139 1567 140 1571
rect 134 1566 140 1567
rect 254 1571 260 1572
rect 254 1567 255 1571
rect 259 1567 260 1571
rect 254 1566 260 1567
rect 422 1571 428 1572
rect 422 1567 423 1571
rect 427 1567 428 1571
rect 422 1566 428 1567
rect 614 1571 620 1572
rect 614 1567 615 1571
rect 619 1567 620 1571
rect 614 1566 620 1567
rect 830 1571 836 1572
rect 830 1567 831 1571
rect 835 1567 836 1571
rect 830 1566 836 1567
rect 1062 1571 1068 1572
rect 1062 1567 1063 1571
rect 1067 1567 1068 1571
rect 1062 1566 1068 1567
rect 1310 1571 1316 1572
rect 1310 1567 1311 1571
rect 1315 1567 1316 1571
rect 1310 1566 1316 1567
rect 1566 1571 1572 1572
rect 1566 1567 1567 1571
rect 1571 1567 1572 1571
rect 1566 1566 1572 1567
rect 1830 1571 1836 1572
rect 1830 1567 1831 1571
rect 1835 1567 1836 1571
rect 2006 1568 2007 1572
rect 2011 1568 2012 1572
rect 2006 1567 2012 1568
rect 1830 1566 1836 1567
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 2006 1555 2012 1556
rect 2048 1555 2050 1582
rect 2390 1580 2391 1584
rect 2395 1580 2396 1584
rect 2390 1579 2396 1580
rect 2502 1584 2508 1585
rect 2502 1580 2503 1584
rect 2507 1580 2508 1584
rect 2502 1579 2508 1580
rect 2614 1584 2620 1585
rect 2614 1580 2615 1584
rect 2619 1580 2620 1584
rect 2614 1579 2620 1580
rect 2734 1584 2740 1585
rect 2734 1580 2735 1584
rect 2739 1580 2740 1584
rect 2734 1579 2740 1580
rect 2854 1584 2860 1585
rect 2854 1580 2855 1584
rect 2859 1580 2860 1584
rect 2854 1579 2860 1580
rect 2974 1584 2980 1585
rect 2974 1580 2975 1584
rect 2979 1580 2980 1584
rect 2974 1579 2980 1580
rect 3094 1584 3100 1585
rect 3094 1580 3095 1584
rect 3099 1580 3100 1584
rect 3094 1579 3100 1580
rect 3214 1584 3220 1585
rect 3214 1580 3215 1584
rect 3219 1580 3220 1584
rect 3214 1579 3220 1580
rect 3334 1584 3340 1585
rect 3334 1580 3335 1584
rect 3339 1580 3340 1584
rect 3334 1579 3340 1580
rect 3454 1584 3460 1585
rect 3454 1580 3455 1584
rect 3459 1580 3460 1584
rect 3942 1583 3943 1587
rect 3947 1583 3948 1587
rect 3942 1582 3948 1583
rect 3454 1579 3460 1580
rect 2392 1555 2394 1579
rect 2504 1555 2506 1579
rect 2616 1555 2618 1579
rect 2736 1555 2738 1579
rect 2856 1555 2858 1579
rect 2976 1555 2978 1579
rect 3096 1555 3098 1579
rect 3216 1555 3218 1579
rect 3336 1555 3338 1579
rect 3456 1555 3458 1579
rect 3944 1555 3946 1582
rect 110 1550 116 1551
rect 134 1552 140 1553
rect 112 1519 114 1550
rect 134 1548 135 1552
rect 139 1548 140 1552
rect 134 1547 140 1548
rect 254 1552 260 1553
rect 254 1548 255 1552
rect 259 1548 260 1552
rect 254 1547 260 1548
rect 422 1552 428 1553
rect 422 1548 423 1552
rect 427 1548 428 1552
rect 422 1547 428 1548
rect 614 1552 620 1553
rect 614 1548 615 1552
rect 619 1548 620 1552
rect 614 1547 620 1548
rect 830 1552 836 1553
rect 830 1548 831 1552
rect 835 1548 836 1552
rect 830 1547 836 1548
rect 1062 1552 1068 1553
rect 1062 1548 1063 1552
rect 1067 1548 1068 1552
rect 1062 1547 1068 1548
rect 1310 1552 1316 1553
rect 1310 1548 1311 1552
rect 1315 1548 1316 1552
rect 1310 1547 1316 1548
rect 1566 1552 1572 1553
rect 1566 1548 1567 1552
rect 1571 1548 1572 1552
rect 1566 1547 1572 1548
rect 1830 1552 1836 1553
rect 1830 1548 1831 1552
rect 1835 1548 1836 1552
rect 2006 1551 2007 1555
rect 2011 1551 2012 1555
rect 2006 1550 2012 1551
rect 2047 1554 2051 1555
rect 1830 1547 1836 1548
rect 136 1519 138 1547
rect 256 1519 258 1547
rect 424 1519 426 1547
rect 616 1519 618 1547
rect 832 1519 834 1547
rect 1064 1519 1066 1547
rect 1312 1519 1314 1547
rect 1568 1519 1570 1547
rect 1832 1519 1834 1547
rect 2008 1519 2010 1550
rect 2047 1549 2051 1550
rect 2391 1554 2395 1555
rect 2391 1549 2395 1550
rect 2503 1554 2507 1555
rect 2503 1549 2507 1550
rect 2543 1554 2547 1555
rect 2543 1549 2547 1550
rect 2615 1554 2619 1555
rect 2615 1549 2619 1550
rect 2671 1554 2675 1555
rect 2671 1549 2675 1550
rect 2735 1554 2739 1555
rect 2735 1549 2739 1550
rect 2799 1554 2803 1555
rect 2799 1549 2803 1550
rect 2855 1554 2859 1555
rect 2855 1549 2859 1550
rect 2935 1554 2939 1555
rect 2935 1549 2939 1550
rect 2975 1554 2979 1555
rect 2975 1549 2979 1550
rect 3071 1554 3075 1555
rect 3071 1549 3075 1550
rect 3095 1554 3099 1555
rect 3095 1549 3099 1550
rect 3207 1554 3211 1555
rect 3207 1549 3211 1550
rect 3215 1554 3219 1555
rect 3215 1549 3219 1550
rect 3335 1554 3339 1555
rect 3335 1549 3339 1550
rect 3455 1554 3459 1555
rect 3455 1549 3459 1550
rect 3463 1554 3467 1555
rect 3463 1549 3467 1550
rect 3591 1554 3595 1555
rect 3591 1549 3595 1550
rect 3727 1554 3731 1555
rect 3727 1549 3731 1550
rect 3839 1554 3843 1555
rect 3839 1549 3843 1550
rect 3943 1554 3947 1555
rect 3943 1549 3947 1550
rect 2048 1522 2050 1549
rect 2544 1525 2546 1549
rect 2672 1525 2674 1549
rect 2800 1525 2802 1549
rect 2936 1525 2938 1549
rect 3072 1525 3074 1549
rect 3208 1525 3210 1549
rect 3336 1525 3338 1549
rect 3464 1525 3466 1549
rect 3592 1525 3594 1549
rect 3728 1525 3730 1549
rect 3840 1525 3842 1549
rect 2542 1524 2548 1525
rect 2046 1521 2052 1522
rect 111 1518 115 1519
rect 111 1513 115 1514
rect 135 1518 139 1519
rect 135 1513 139 1514
rect 239 1518 243 1519
rect 239 1513 243 1514
rect 255 1518 259 1519
rect 255 1513 259 1514
rect 407 1518 411 1519
rect 407 1513 411 1514
rect 423 1518 427 1519
rect 423 1513 427 1514
rect 583 1518 587 1519
rect 583 1513 587 1514
rect 615 1518 619 1519
rect 615 1513 619 1514
rect 775 1518 779 1519
rect 775 1513 779 1514
rect 831 1518 835 1519
rect 831 1513 835 1514
rect 967 1518 971 1519
rect 967 1513 971 1514
rect 1063 1518 1067 1519
rect 1063 1513 1067 1514
rect 1159 1518 1163 1519
rect 1159 1513 1163 1514
rect 1311 1518 1315 1519
rect 1311 1513 1315 1514
rect 1351 1518 1355 1519
rect 1351 1513 1355 1514
rect 1543 1518 1547 1519
rect 1543 1513 1547 1514
rect 1567 1518 1571 1519
rect 1567 1513 1571 1514
rect 1735 1518 1739 1519
rect 1735 1513 1739 1514
rect 1831 1518 1835 1519
rect 1831 1513 1835 1514
rect 1903 1518 1907 1519
rect 1903 1513 1907 1514
rect 2007 1518 2011 1519
rect 2046 1517 2047 1521
rect 2051 1517 2052 1521
rect 2542 1520 2543 1524
rect 2547 1520 2548 1524
rect 2542 1519 2548 1520
rect 2670 1524 2676 1525
rect 2670 1520 2671 1524
rect 2675 1520 2676 1524
rect 2670 1519 2676 1520
rect 2798 1524 2804 1525
rect 2798 1520 2799 1524
rect 2803 1520 2804 1524
rect 2798 1519 2804 1520
rect 2934 1524 2940 1525
rect 2934 1520 2935 1524
rect 2939 1520 2940 1524
rect 2934 1519 2940 1520
rect 3070 1524 3076 1525
rect 3070 1520 3071 1524
rect 3075 1520 3076 1524
rect 3070 1519 3076 1520
rect 3206 1524 3212 1525
rect 3206 1520 3207 1524
rect 3211 1520 3212 1524
rect 3206 1519 3212 1520
rect 3334 1524 3340 1525
rect 3334 1520 3335 1524
rect 3339 1520 3340 1524
rect 3334 1519 3340 1520
rect 3462 1524 3468 1525
rect 3462 1520 3463 1524
rect 3467 1520 3468 1524
rect 3462 1519 3468 1520
rect 3590 1524 3596 1525
rect 3590 1520 3591 1524
rect 3595 1520 3596 1524
rect 3590 1519 3596 1520
rect 3726 1524 3732 1525
rect 3726 1520 3727 1524
rect 3731 1520 3732 1524
rect 3726 1519 3732 1520
rect 3838 1524 3844 1525
rect 3838 1520 3839 1524
rect 3843 1520 3844 1524
rect 3944 1522 3946 1549
rect 3838 1519 3844 1520
rect 3942 1521 3948 1522
rect 2046 1516 2052 1517
rect 3942 1517 3943 1521
rect 3947 1517 3948 1521
rect 3942 1516 3948 1517
rect 2007 1513 2011 1514
rect 112 1486 114 1513
rect 240 1489 242 1513
rect 408 1489 410 1513
rect 584 1489 586 1513
rect 776 1489 778 1513
rect 968 1489 970 1513
rect 1160 1489 1162 1513
rect 1352 1489 1354 1513
rect 1544 1489 1546 1513
rect 1736 1489 1738 1513
rect 1904 1489 1906 1513
rect 238 1488 244 1489
rect 110 1485 116 1486
rect 110 1481 111 1485
rect 115 1481 116 1485
rect 238 1484 239 1488
rect 243 1484 244 1488
rect 238 1483 244 1484
rect 406 1488 412 1489
rect 406 1484 407 1488
rect 411 1484 412 1488
rect 406 1483 412 1484
rect 582 1488 588 1489
rect 582 1484 583 1488
rect 587 1484 588 1488
rect 582 1483 588 1484
rect 774 1488 780 1489
rect 774 1484 775 1488
rect 779 1484 780 1488
rect 774 1483 780 1484
rect 966 1488 972 1489
rect 966 1484 967 1488
rect 971 1484 972 1488
rect 966 1483 972 1484
rect 1158 1488 1164 1489
rect 1158 1484 1159 1488
rect 1163 1484 1164 1488
rect 1158 1483 1164 1484
rect 1350 1488 1356 1489
rect 1350 1484 1351 1488
rect 1355 1484 1356 1488
rect 1350 1483 1356 1484
rect 1542 1488 1548 1489
rect 1542 1484 1543 1488
rect 1547 1484 1548 1488
rect 1542 1483 1548 1484
rect 1734 1488 1740 1489
rect 1734 1484 1735 1488
rect 1739 1484 1740 1488
rect 1734 1483 1740 1484
rect 1902 1488 1908 1489
rect 1902 1484 1903 1488
rect 1907 1484 1908 1488
rect 2008 1486 2010 1513
rect 2542 1505 2548 1506
rect 2046 1504 2052 1505
rect 2046 1500 2047 1504
rect 2051 1500 2052 1504
rect 2542 1501 2543 1505
rect 2547 1501 2548 1505
rect 2542 1500 2548 1501
rect 2670 1505 2676 1506
rect 2670 1501 2671 1505
rect 2675 1501 2676 1505
rect 2670 1500 2676 1501
rect 2798 1505 2804 1506
rect 2798 1501 2799 1505
rect 2803 1501 2804 1505
rect 2798 1500 2804 1501
rect 2934 1505 2940 1506
rect 2934 1501 2935 1505
rect 2939 1501 2940 1505
rect 2934 1500 2940 1501
rect 3070 1505 3076 1506
rect 3070 1501 3071 1505
rect 3075 1501 3076 1505
rect 3070 1500 3076 1501
rect 3206 1505 3212 1506
rect 3206 1501 3207 1505
rect 3211 1501 3212 1505
rect 3206 1500 3212 1501
rect 3334 1505 3340 1506
rect 3334 1501 3335 1505
rect 3339 1501 3340 1505
rect 3334 1500 3340 1501
rect 3462 1505 3468 1506
rect 3462 1501 3463 1505
rect 3467 1501 3468 1505
rect 3462 1500 3468 1501
rect 3590 1505 3596 1506
rect 3590 1501 3591 1505
rect 3595 1501 3596 1505
rect 3590 1500 3596 1501
rect 3726 1505 3732 1506
rect 3726 1501 3727 1505
rect 3731 1501 3732 1505
rect 3726 1500 3732 1501
rect 3838 1505 3844 1506
rect 3838 1501 3839 1505
rect 3843 1501 3844 1505
rect 3838 1500 3844 1501
rect 3942 1504 3948 1505
rect 3942 1500 3943 1504
rect 3947 1500 3948 1504
rect 2046 1499 2052 1500
rect 1902 1483 1908 1484
rect 2006 1485 2012 1486
rect 110 1480 116 1481
rect 2006 1481 2007 1485
rect 2011 1481 2012 1485
rect 2006 1480 2012 1481
rect 238 1469 244 1470
rect 110 1468 116 1469
rect 110 1464 111 1468
rect 115 1464 116 1468
rect 238 1465 239 1469
rect 243 1465 244 1469
rect 238 1464 244 1465
rect 406 1469 412 1470
rect 406 1465 407 1469
rect 411 1465 412 1469
rect 406 1464 412 1465
rect 582 1469 588 1470
rect 582 1465 583 1469
rect 587 1465 588 1469
rect 582 1464 588 1465
rect 774 1469 780 1470
rect 774 1465 775 1469
rect 779 1465 780 1469
rect 774 1464 780 1465
rect 966 1469 972 1470
rect 966 1465 967 1469
rect 971 1465 972 1469
rect 966 1464 972 1465
rect 1158 1469 1164 1470
rect 1158 1465 1159 1469
rect 1163 1465 1164 1469
rect 1158 1464 1164 1465
rect 1350 1469 1356 1470
rect 1350 1465 1351 1469
rect 1355 1465 1356 1469
rect 1350 1464 1356 1465
rect 1542 1469 1548 1470
rect 1542 1465 1543 1469
rect 1547 1465 1548 1469
rect 1542 1464 1548 1465
rect 1734 1469 1740 1470
rect 1734 1465 1735 1469
rect 1739 1465 1740 1469
rect 1734 1464 1740 1465
rect 1902 1469 1908 1470
rect 1902 1465 1903 1469
rect 1907 1465 1908 1469
rect 1902 1464 1908 1465
rect 2006 1468 2012 1469
rect 2006 1464 2007 1468
rect 2011 1464 2012 1468
rect 2048 1467 2050 1499
rect 2544 1467 2546 1500
rect 2672 1467 2674 1500
rect 2800 1467 2802 1500
rect 2936 1467 2938 1500
rect 3072 1467 3074 1500
rect 3208 1467 3210 1500
rect 3336 1467 3338 1500
rect 3464 1467 3466 1500
rect 3592 1467 3594 1500
rect 3728 1467 3730 1500
rect 3840 1467 3842 1500
rect 3942 1499 3948 1500
rect 3944 1467 3946 1499
rect 110 1463 116 1464
rect 112 1435 114 1463
rect 240 1435 242 1464
rect 408 1435 410 1464
rect 584 1435 586 1464
rect 776 1435 778 1464
rect 968 1435 970 1464
rect 1160 1435 1162 1464
rect 1352 1435 1354 1464
rect 1544 1435 1546 1464
rect 1736 1435 1738 1464
rect 1904 1435 1906 1464
rect 2006 1463 2012 1464
rect 2047 1466 2051 1467
rect 2008 1435 2010 1463
rect 2047 1461 2051 1462
rect 2519 1466 2523 1467
rect 2519 1461 2523 1462
rect 2543 1466 2547 1467
rect 2543 1461 2547 1462
rect 2631 1466 2635 1467
rect 2631 1461 2635 1462
rect 2671 1466 2675 1467
rect 2671 1461 2675 1462
rect 2759 1466 2763 1467
rect 2759 1461 2763 1462
rect 2799 1466 2803 1467
rect 2799 1461 2803 1462
rect 2895 1466 2899 1467
rect 2895 1461 2899 1462
rect 2935 1466 2939 1467
rect 2935 1461 2939 1462
rect 3031 1466 3035 1467
rect 3031 1461 3035 1462
rect 3071 1466 3075 1467
rect 3071 1461 3075 1462
rect 3175 1466 3179 1467
rect 3175 1461 3179 1462
rect 3207 1466 3211 1467
rect 3207 1461 3211 1462
rect 3311 1466 3315 1467
rect 3311 1461 3315 1462
rect 3335 1466 3339 1467
rect 3335 1461 3339 1462
rect 3447 1466 3451 1467
rect 3447 1461 3451 1462
rect 3463 1466 3467 1467
rect 3463 1461 3467 1462
rect 3583 1466 3587 1467
rect 3583 1461 3587 1462
rect 3591 1466 3595 1467
rect 3591 1461 3595 1462
rect 3719 1466 3723 1467
rect 3719 1461 3723 1462
rect 3727 1466 3731 1467
rect 3727 1461 3731 1462
rect 3839 1466 3843 1467
rect 3839 1461 3843 1462
rect 3943 1466 3947 1467
rect 3943 1461 3947 1462
rect 2048 1441 2050 1461
rect 2046 1440 2052 1441
rect 2520 1440 2522 1461
rect 2632 1440 2634 1461
rect 2760 1440 2762 1461
rect 2896 1440 2898 1461
rect 3032 1440 3034 1461
rect 3176 1440 3178 1461
rect 3312 1440 3314 1461
rect 3448 1440 3450 1461
rect 3584 1440 3586 1461
rect 3720 1440 3722 1461
rect 3840 1440 3842 1461
rect 3944 1441 3946 1461
rect 3942 1440 3948 1441
rect 2046 1436 2047 1440
rect 2051 1436 2052 1440
rect 2046 1435 2052 1436
rect 2518 1439 2524 1440
rect 2518 1435 2519 1439
rect 2523 1435 2524 1439
rect 111 1434 115 1435
rect 111 1429 115 1430
rect 239 1434 243 1435
rect 239 1429 243 1430
rect 407 1434 411 1435
rect 407 1429 411 1430
rect 463 1434 467 1435
rect 463 1429 467 1430
rect 583 1434 587 1435
rect 583 1429 587 1430
rect 711 1434 715 1435
rect 711 1429 715 1430
rect 775 1434 779 1435
rect 775 1429 779 1430
rect 855 1434 859 1435
rect 855 1429 859 1430
rect 967 1434 971 1435
rect 967 1429 971 1430
rect 1007 1434 1011 1435
rect 1007 1429 1011 1430
rect 1159 1434 1163 1435
rect 1159 1429 1163 1430
rect 1167 1434 1171 1435
rect 1167 1429 1171 1430
rect 1335 1434 1339 1435
rect 1335 1429 1339 1430
rect 1351 1434 1355 1435
rect 1351 1429 1355 1430
rect 1511 1434 1515 1435
rect 1511 1429 1515 1430
rect 1543 1434 1547 1435
rect 1543 1429 1547 1430
rect 1687 1434 1691 1435
rect 1687 1429 1691 1430
rect 1735 1434 1739 1435
rect 1735 1429 1739 1430
rect 1871 1434 1875 1435
rect 1871 1429 1875 1430
rect 1903 1434 1907 1435
rect 1903 1429 1907 1430
rect 2007 1434 2011 1435
rect 2518 1434 2524 1435
rect 2630 1439 2636 1440
rect 2630 1435 2631 1439
rect 2635 1435 2636 1439
rect 2630 1434 2636 1435
rect 2758 1439 2764 1440
rect 2758 1435 2759 1439
rect 2763 1435 2764 1439
rect 2758 1434 2764 1435
rect 2894 1439 2900 1440
rect 2894 1435 2895 1439
rect 2899 1435 2900 1439
rect 2894 1434 2900 1435
rect 3030 1439 3036 1440
rect 3030 1435 3031 1439
rect 3035 1435 3036 1439
rect 3030 1434 3036 1435
rect 3174 1439 3180 1440
rect 3174 1435 3175 1439
rect 3179 1435 3180 1439
rect 3174 1434 3180 1435
rect 3310 1439 3316 1440
rect 3310 1435 3311 1439
rect 3315 1435 3316 1439
rect 3310 1434 3316 1435
rect 3446 1439 3452 1440
rect 3446 1435 3447 1439
rect 3451 1435 3452 1439
rect 3446 1434 3452 1435
rect 3582 1439 3588 1440
rect 3582 1435 3583 1439
rect 3587 1435 3588 1439
rect 3582 1434 3588 1435
rect 3718 1439 3724 1440
rect 3718 1435 3719 1439
rect 3723 1435 3724 1439
rect 3718 1434 3724 1435
rect 3838 1439 3844 1440
rect 3838 1435 3839 1439
rect 3843 1435 3844 1439
rect 3942 1436 3943 1440
rect 3947 1436 3948 1440
rect 3942 1435 3948 1436
rect 3838 1434 3844 1435
rect 2007 1429 2011 1430
rect 112 1409 114 1429
rect 110 1408 116 1409
rect 464 1408 466 1429
rect 584 1408 586 1429
rect 712 1408 714 1429
rect 856 1408 858 1429
rect 1008 1408 1010 1429
rect 1168 1408 1170 1429
rect 1336 1408 1338 1429
rect 1512 1408 1514 1429
rect 1688 1408 1690 1429
rect 1872 1408 1874 1429
rect 2008 1409 2010 1429
rect 2046 1423 2052 1424
rect 2046 1419 2047 1423
rect 2051 1419 2052 1423
rect 3942 1423 3948 1424
rect 2046 1418 2052 1419
rect 2518 1420 2524 1421
rect 2006 1408 2012 1409
rect 110 1404 111 1408
rect 115 1404 116 1408
rect 110 1403 116 1404
rect 462 1407 468 1408
rect 462 1403 463 1407
rect 467 1403 468 1407
rect 462 1402 468 1403
rect 582 1407 588 1408
rect 582 1403 583 1407
rect 587 1403 588 1407
rect 582 1402 588 1403
rect 710 1407 716 1408
rect 710 1403 711 1407
rect 715 1403 716 1407
rect 710 1402 716 1403
rect 854 1407 860 1408
rect 854 1403 855 1407
rect 859 1403 860 1407
rect 854 1402 860 1403
rect 1006 1407 1012 1408
rect 1006 1403 1007 1407
rect 1011 1403 1012 1407
rect 1006 1402 1012 1403
rect 1166 1407 1172 1408
rect 1166 1403 1167 1407
rect 1171 1403 1172 1407
rect 1166 1402 1172 1403
rect 1334 1407 1340 1408
rect 1334 1403 1335 1407
rect 1339 1403 1340 1407
rect 1334 1402 1340 1403
rect 1510 1407 1516 1408
rect 1510 1403 1511 1407
rect 1515 1403 1516 1407
rect 1510 1402 1516 1403
rect 1686 1407 1692 1408
rect 1686 1403 1687 1407
rect 1691 1403 1692 1407
rect 1686 1402 1692 1403
rect 1870 1407 1876 1408
rect 1870 1403 1871 1407
rect 1875 1403 1876 1407
rect 2006 1404 2007 1408
rect 2011 1404 2012 1408
rect 2006 1403 2012 1404
rect 1870 1402 1876 1403
rect 110 1391 116 1392
rect 110 1387 111 1391
rect 115 1387 116 1391
rect 2006 1391 2012 1392
rect 2048 1391 2050 1418
rect 2518 1416 2519 1420
rect 2523 1416 2524 1420
rect 2518 1415 2524 1416
rect 2630 1420 2636 1421
rect 2630 1416 2631 1420
rect 2635 1416 2636 1420
rect 2630 1415 2636 1416
rect 2758 1420 2764 1421
rect 2758 1416 2759 1420
rect 2763 1416 2764 1420
rect 2758 1415 2764 1416
rect 2894 1420 2900 1421
rect 2894 1416 2895 1420
rect 2899 1416 2900 1420
rect 2894 1415 2900 1416
rect 3030 1420 3036 1421
rect 3030 1416 3031 1420
rect 3035 1416 3036 1420
rect 3030 1415 3036 1416
rect 3174 1420 3180 1421
rect 3174 1416 3175 1420
rect 3179 1416 3180 1420
rect 3174 1415 3180 1416
rect 3310 1420 3316 1421
rect 3310 1416 3311 1420
rect 3315 1416 3316 1420
rect 3310 1415 3316 1416
rect 3446 1420 3452 1421
rect 3446 1416 3447 1420
rect 3451 1416 3452 1420
rect 3446 1415 3452 1416
rect 3582 1420 3588 1421
rect 3582 1416 3583 1420
rect 3587 1416 3588 1420
rect 3582 1415 3588 1416
rect 3718 1420 3724 1421
rect 3718 1416 3719 1420
rect 3723 1416 3724 1420
rect 3718 1415 3724 1416
rect 3838 1420 3844 1421
rect 3838 1416 3839 1420
rect 3843 1416 3844 1420
rect 3942 1419 3943 1423
rect 3947 1419 3948 1423
rect 3942 1418 3948 1419
rect 3838 1415 3844 1416
rect 2520 1391 2522 1415
rect 2632 1391 2634 1415
rect 2760 1391 2762 1415
rect 2896 1391 2898 1415
rect 3032 1391 3034 1415
rect 3176 1391 3178 1415
rect 3312 1391 3314 1415
rect 3448 1391 3450 1415
rect 3584 1391 3586 1415
rect 3720 1391 3722 1415
rect 3840 1391 3842 1415
rect 3944 1391 3946 1418
rect 110 1386 116 1387
rect 462 1388 468 1389
rect 112 1359 114 1386
rect 462 1384 463 1388
rect 467 1384 468 1388
rect 462 1383 468 1384
rect 582 1388 588 1389
rect 582 1384 583 1388
rect 587 1384 588 1388
rect 582 1383 588 1384
rect 710 1388 716 1389
rect 710 1384 711 1388
rect 715 1384 716 1388
rect 710 1383 716 1384
rect 854 1388 860 1389
rect 854 1384 855 1388
rect 859 1384 860 1388
rect 854 1383 860 1384
rect 1006 1388 1012 1389
rect 1006 1384 1007 1388
rect 1011 1384 1012 1388
rect 1006 1383 1012 1384
rect 1166 1388 1172 1389
rect 1166 1384 1167 1388
rect 1171 1384 1172 1388
rect 1166 1383 1172 1384
rect 1334 1388 1340 1389
rect 1334 1384 1335 1388
rect 1339 1384 1340 1388
rect 1334 1383 1340 1384
rect 1510 1388 1516 1389
rect 1510 1384 1511 1388
rect 1515 1384 1516 1388
rect 1510 1383 1516 1384
rect 1686 1388 1692 1389
rect 1686 1384 1687 1388
rect 1691 1384 1692 1388
rect 1686 1383 1692 1384
rect 1870 1388 1876 1389
rect 1870 1384 1871 1388
rect 1875 1384 1876 1388
rect 2006 1387 2007 1391
rect 2011 1387 2012 1391
rect 2006 1386 2012 1387
rect 2047 1390 2051 1391
rect 1870 1383 1876 1384
rect 464 1359 466 1383
rect 584 1359 586 1383
rect 712 1359 714 1383
rect 856 1359 858 1383
rect 1008 1359 1010 1383
rect 1168 1359 1170 1383
rect 1336 1359 1338 1383
rect 1512 1359 1514 1383
rect 1688 1359 1690 1383
rect 1872 1359 1874 1383
rect 2008 1359 2010 1386
rect 2047 1385 2051 1386
rect 2399 1390 2403 1391
rect 2399 1385 2403 1386
rect 2519 1390 2523 1391
rect 2519 1385 2523 1386
rect 2535 1390 2539 1391
rect 2535 1385 2539 1386
rect 2631 1390 2635 1391
rect 2631 1385 2635 1386
rect 2679 1390 2683 1391
rect 2679 1385 2683 1386
rect 2759 1390 2763 1391
rect 2759 1385 2763 1386
rect 2823 1390 2827 1391
rect 2823 1385 2827 1386
rect 2895 1390 2899 1391
rect 2895 1385 2899 1386
rect 2967 1390 2971 1391
rect 2967 1385 2971 1386
rect 3031 1390 3035 1391
rect 3031 1385 3035 1386
rect 3111 1390 3115 1391
rect 3111 1385 3115 1386
rect 3175 1390 3179 1391
rect 3175 1385 3179 1386
rect 3255 1390 3259 1391
rect 3255 1385 3259 1386
rect 3311 1390 3315 1391
rect 3311 1385 3315 1386
rect 3407 1390 3411 1391
rect 3407 1385 3411 1386
rect 3447 1390 3451 1391
rect 3447 1385 3451 1386
rect 3559 1390 3563 1391
rect 3559 1385 3563 1386
rect 3583 1390 3587 1391
rect 3583 1385 3587 1386
rect 3711 1390 3715 1391
rect 3711 1385 3715 1386
rect 3719 1390 3723 1391
rect 3719 1385 3723 1386
rect 3839 1390 3843 1391
rect 3839 1385 3843 1386
rect 3943 1390 3947 1391
rect 3943 1385 3947 1386
rect 111 1358 115 1359
rect 111 1353 115 1354
rect 463 1358 467 1359
rect 463 1353 467 1354
rect 583 1358 587 1359
rect 583 1353 587 1354
rect 655 1358 659 1359
rect 655 1353 659 1354
rect 711 1358 715 1359
rect 711 1353 715 1354
rect 767 1358 771 1359
rect 767 1353 771 1354
rect 855 1358 859 1359
rect 855 1353 859 1354
rect 887 1358 891 1359
rect 887 1353 891 1354
rect 1007 1358 1011 1359
rect 1007 1353 1011 1354
rect 1015 1358 1019 1359
rect 1015 1353 1019 1354
rect 1143 1358 1147 1359
rect 1143 1353 1147 1354
rect 1167 1358 1171 1359
rect 1167 1353 1171 1354
rect 1279 1358 1283 1359
rect 1279 1353 1283 1354
rect 1335 1358 1339 1359
rect 1335 1353 1339 1354
rect 1415 1358 1419 1359
rect 1415 1353 1419 1354
rect 1511 1358 1515 1359
rect 1511 1353 1515 1354
rect 1559 1358 1563 1359
rect 1559 1353 1563 1354
rect 1687 1358 1691 1359
rect 1687 1353 1691 1354
rect 1703 1358 1707 1359
rect 1703 1353 1707 1354
rect 1847 1358 1851 1359
rect 1847 1353 1851 1354
rect 1871 1358 1875 1359
rect 1871 1353 1875 1354
rect 2007 1358 2011 1359
rect 2048 1358 2050 1385
rect 2400 1361 2402 1385
rect 2536 1361 2538 1385
rect 2680 1361 2682 1385
rect 2824 1361 2826 1385
rect 2968 1361 2970 1385
rect 3112 1361 3114 1385
rect 3256 1361 3258 1385
rect 3408 1361 3410 1385
rect 3560 1361 3562 1385
rect 3712 1361 3714 1385
rect 3840 1361 3842 1385
rect 2398 1360 2404 1361
rect 2007 1353 2011 1354
rect 2046 1357 2052 1358
rect 2046 1353 2047 1357
rect 2051 1353 2052 1357
rect 2398 1356 2399 1360
rect 2403 1356 2404 1360
rect 2398 1355 2404 1356
rect 2534 1360 2540 1361
rect 2534 1356 2535 1360
rect 2539 1356 2540 1360
rect 2534 1355 2540 1356
rect 2678 1360 2684 1361
rect 2678 1356 2679 1360
rect 2683 1356 2684 1360
rect 2678 1355 2684 1356
rect 2822 1360 2828 1361
rect 2822 1356 2823 1360
rect 2827 1356 2828 1360
rect 2822 1355 2828 1356
rect 2966 1360 2972 1361
rect 2966 1356 2967 1360
rect 2971 1356 2972 1360
rect 2966 1355 2972 1356
rect 3110 1360 3116 1361
rect 3110 1356 3111 1360
rect 3115 1356 3116 1360
rect 3110 1355 3116 1356
rect 3254 1360 3260 1361
rect 3254 1356 3255 1360
rect 3259 1356 3260 1360
rect 3254 1355 3260 1356
rect 3406 1360 3412 1361
rect 3406 1356 3407 1360
rect 3411 1356 3412 1360
rect 3406 1355 3412 1356
rect 3558 1360 3564 1361
rect 3558 1356 3559 1360
rect 3563 1356 3564 1360
rect 3558 1355 3564 1356
rect 3710 1360 3716 1361
rect 3710 1356 3711 1360
rect 3715 1356 3716 1360
rect 3710 1355 3716 1356
rect 3838 1360 3844 1361
rect 3838 1356 3839 1360
rect 3843 1356 3844 1360
rect 3944 1358 3946 1385
rect 3838 1355 3844 1356
rect 3942 1357 3948 1358
rect 112 1326 114 1353
rect 656 1329 658 1353
rect 768 1329 770 1353
rect 888 1329 890 1353
rect 1016 1329 1018 1353
rect 1144 1329 1146 1353
rect 1280 1329 1282 1353
rect 1416 1329 1418 1353
rect 1560 1329 1562 1353
rect 1704 1329 1706 1353
rect 1848 1329 1850 1353
rect 654 1328 660 1329
rect 110 1325 116 1326
rect 110 1321 111 1325
rect 115 1321 116 1325
rect 654 1324 655 1328
rect 659 1324 660 1328
rect 654 1323 660 1324
rect 766 1328 772 1329
rect 766 1324 767 1328
rect 771 1324 772 1328
rect 766 1323 772 1324
rect 886 1328 892 1329
rect 886 1324 887 1328
rect 891 1324 892 1328
rect 886 1323 892 1324
rect 1014 1328 1020 1329
rect 1014 1324 1015 1328
rect 1019 1324 1020 1328
rect 1014 1323 1020 1324
rect 1142 1328 1148 1329
rect 1142 1324 1143 1328
rect 1147 1324 1148 1328
rect 1142 1323 1148 1324
rect 1278 1328 1284 1329
rect 1278 1324 1279 1328
rect 1283 1324 1284 1328
rect 1278 1323 1284 1324
rect 1414 1328 1420 1329
rect 1414 1324 1415 1328
rect 1419 1324 1420 1328
rect 1414 1323 1420 1324
rect 1558 1328 1564 1329
rect 1558 1324 1559 1328
rect 1563 1324 1564 1328
rect 1558 1323 1564 1324
rect 1702 1328 1708 1329
rect 1702 1324 1703 1328
rect 1707 1324 1708 1328
rect 1702 1323 1708 1324
rect 1846 1328 1852 1329
rect 1846 1324 1847 1328
rect 1851 1324 1852 1328
rect 2008 1326 2010 1353
rect 2046 1352 2052 1353
rect 3942 1353 3943 1357
rect 3947 1353 3948 1357
rect 3942 1352 3948 1353
rect 2398 1341 2404 1342
rect 2046 1340 2052 1341
rect 2046 1336 2047 1340
rect 2051 1336 2052 1340
rect 2398 1337 2399 1341
rect 2403 1337 2404 1341
rect 2398 1336 2404 1337
rect 2534 1341 2540 1342
rect 2534 1337 2535 1341
rect 2539 1337 2540 1341
rect 2534 1336 2540 1337
rect 2678 1341 2684 1342
rect 2678 1337 2679 1341
rect 2683 1337 2684 1341
rect 2678 1336 2684 1337
rect 2822 1341 2828 1342
rect 2822 1337 2823 1341
rect 2827 1337 2828 1341
rect 2822 1336 2828 1337
rect 2966 1341 2972 1342
rect 2966 1337 2967 1341
rect 2971 1337 2972 1341
rect 2966 1336 2972 1337
rect 3110 1341 3116 1342
rect 3110 1337 3111 1341
rect 3115 1337 3116 1341
rect 3110 1336 3116 1337
rect 3254 1341 3260 1342
rect 3254 1337 3255 1341
rect 3259 1337 3260 1341
rect 3254 1336 3260 1337
rect 3406 1341 3412 1342
rect 3406 1337 3407 1341
rect 3411 1337 3412 1341
rect 3406 1336 3412 1337
rect 3558 1341 3564 1342
rect 3558 1337 3559 1341
rect 3563 1337 3564 1341
rect 3558 1336 3564 1337
rect 3710 1341 3716 1342
rect 3710 1337 3711 1341
rect 3715 1337 3716 1341
rect 3710 1336 3716 1337
rect 3838 1341 3844 1342
rect 3838 1337 3839 1341
rect 3843 1337 3844 1341
rect 3838 1336 3844 1337
rect 3942 1340 3948 1341
rect 3942 1336 3943 1340
rect 3947 1336 3948 1340
rect 2046 1335 2052 1336
rect 1846 1323 1852 1324
rect 2006 1325 2012 1326
rect 110 1320 116 1321
rect 2006 1321 2007 1325
rect 2011 1321 2012 1325
rect 2006 1320 2012 1321
rect 2048 1311 2050 1335
rect 2400 1311 2402 1336
rect 2536 1311 2538 1336
rect 2680 1311 2682 1336
rect 2824 1311 2826 1336
rect 2968 1311 2970 1336
rect 3112 1311 3114 1336
rect 3256 1311 3258 1336
rect 3408 1311 3410 1336
rect 3560 1311 3562 1336
rect 3712 1311 3714 1336
rect 3840 1311 3842 1336
rect 3942 1335 3948 1336
rect 3944 1311 3946 1335
rect 2047 1310 2051 1311
rect 654 1309 660 1310
rect 110 1308 116 1309
rect 110 1304 111 1308
rect 115 1304 116 1308
rect 654 1305 655 1309
rect 659 1305 660 1309
rect 654 1304 660 1305
rect 766 1309 772 1310
rect 766 1305 767 1309
rect 771 1305 772 1309
rect 766 1304 772 1305
rect 886 1309 892 1310
rect 886 1305 887 1309
rect 891 1305 892 1309
rect 886 1304 892 1305
rect 1014 1309 1020 1310
rect 1014 1305 1015 1309
rect 1019 1305 1020 1309
rect 1014 1304 1020 1305
rect 1142 1309 1148 1310
rect 1142 1305 1143 1309
rect 1147 1305 1148 1309
rect 1142 1304 1148 1305
rect 1278 1309 1284 1310
rect 1278 1305 1279 1309
rect 1283 1305 1284 1309
rect 1278 1304 1284 1305
rect 1414 1309 1420 1310
rect 1414 1305 1415 1309
rect 1419 1305 1420 1309
rect 1414 1304 1420 1305
rect 1558 1309 1564 1310
rect 1558 1305 1559 1309
rect 1563 1305 1564 1309
rect 1558 1304 1564 1305
rect 1702 1309 1708 1310
rect 1702 1305 1703 1309
rect 1707 1305 1708 1309
rect 1702 1304 1708 1305
rect 1846 1309 1852 1310
rect 1846 1305 1847 1309
rect 1851 1305 1852 1309
rect 1846 1304 1852 1305
rect 2006 1308 2012 1309
rect 2006 1304 2007 1308
rect 2011 1304 2012 1308
rect 2047 1305 2051 1306
rect 2247 1310 2251 1311
rect 2247 1305 2251 1306
rect 2375 1310 2379 1311
rect 2375 1305 2379 1306
rect 2399 1310 2403 1311
rect 2399 1305 2403 1306
rect 2511 1310 2515 1311
rect 2511 1305 2515 1306
rect 2535 1310 2539 1311
rect 2535 1305 2539 1306
rect 2647 1310 2651 1311
rect 2647 1305 2651 1306
rect 2679 1310 2683 1311
rect 2679 1305 2683 1306
rect 2791 1310 2795 1311
rect 2791 1305 2795 1306
rect 2823 1310 2827 1311
rect 2823 1305 2827 1306
rect 2943 1310 2947 1311
rect 2943 1305 2947 1306
rect 2967 1310 2971 1311
rect 2967 1305 2971 1306
rect 3111 1310 3115 1311
rect 3111 1305 3115 1306
rect 3255 1310 3259 1311
rect 3255 1305 3259 1306
rect 3287 1310 3291 1311
rect 3287 1305 3291 1306
rect 3407 1310 3411 1311
rect 3407 1305 3411 1306
rect 3471 1310 3475 1311
rect 3471 1305 3475 1306
rect 3559 1310 3563 1311
rect 3559 1305 3563 1306
rect 3663 1310 3667 1311
rect 3663 1305 3667 1306
rect 3711 1310 3715 1311
rect 3711 1305 3715 1306
rect 3839 1310 3843 1311
rect 3839 1305 3843 1306
rect 3943 1310 3947 1311
rect 3943 1305 3947 1306
rect 110 1303 116 1304
rect 112 1279 114 1303
rect 656 1279 658 1304
rect 768 1279 770 1304
rect 888 1279 890 1304
rect 1016 1279 1018 1304
rect 1144 1279 1146 1304
rect 1280 1279 1282 1304
rect 1416 1279 1418 1304
rect 1560 1279 1562 1304
rect 1704 1279 1706 1304
rect 1848 1279 1850 1304
rect 2006 1303 2012 1304
rect 2008 1279 2010 1303
rect 2048 1285 2050 1305
rect 2046 1284 2052 1285
rect 2248 1284 2250 1305
rect 2376 1284 2378 1305
rect 2512 1284 2514 1305
rect 2648 1284 2650 1305
rect 2792 1284 2794 1305
rect 2944 1284 2946 1305
rect 3112 1284 3114 1305
rect 3288 1284 3290 1305
rect 3472 1284 3474 1305
rect 3664 1284 3666 1305
rect 3840 1284 3842 1305
rect 3944 1285 3946 1305
rect 3942 1284 3948 1285
rect 2046 1280 2047 1284
rect 2051 1280 2052 1284
rect 2046 1279 2052 1280
rect 2246 1283 2252 1284
rect 2246 1279 2247 1283
rect 2251 1279 2252 1283
rect 111 1278 115 1279
rect 111 1273 115 1274
rect 439 1278 443 1279
rect 439 1273 443 1274
rect 551 1278 555 1279
rect 551 1273 555 1274
rect 655 1278 659 1279
rect 655 1273 659 1274
rect 671 1278 675 1279
rect 671 1273 675 1274
rect 767 1278 771 1279
rect 767 1273 771 1274
rect 799 1278 803 1279
rect 799 1273 803 1274
rect 887 1278 891 1279
rect 887 1273 891 1274
rect 935 1278 939 1279
rect 935 1273 939 1274
rect 1015 1278 1019 1279
rect 1015 1273 1019 1274
rect 1079 1278 1083 1279
rect 1079 1273 1083 1274
rect 1143 1278 1147 1279
rect 1143 1273 1147 1274
rect 1231 1278 1235 1279
rect 1231 1273 1235 1274
rect 1279 1278 1283 1279
rect 1279 1273 1283 1274
rect 1391 1278 1395 1279
rect 1391 1273 1395 1274
rect 1415 1278 1419 1279
rect 1415 1273 1419 1274
rect 1551 1278 1555 1279
rect 1551 1273 1555 1274
rect 1559 1278 1563 1279
rect 1559 1273 1563 1274
rect 1703 1278 1707 1279
rect 1703 1273 1707 1274
rect 1719 1278 1723 1279
rect 1719 1273 1723 1274
rect 1847 1278 1851 1279
rect 1847 1273 1851 1274
rect 2007 1278 2011 1279
rect 2246 1278 2252 1279
rect 2374 1283 2380 1284
rect 2374 1279 2375 1283
rect 2379 1279 2380 1283
rect 2374 1278 2380 1279
rect 2510 1283 2516 1284
rect 2510 1279 2511 1283
rect 2515 1279 2516 1283
rect 2510 1278 2516 1279
rect 2646 1283 2652 1284
rect 2646 1279 2647 1283
rect 2651 1279 2652 1283
rect 2646 1278 2652 1279
rect 2790 1283 2796 1284
rect 2790 1279 2791 1283
rect 2795 1279 2796 1283
rect 2790 1278 2796 1279
rect 2942 1283 2948 1284
rect 2942 1279 2943 1283
rect 2947 1279 2948 1283
rect 2942 1278 2948 1279
rect 3110 1283 3116 1284
rect 3110 1279 3111 1283
rect 3115 1279 3116 1283
rect 3110 1278 3116 1279
rect 3286 1283 3292 1284
rect 3286 1279 3287 1283
rect 3291 1279 3292 1283
rect 3286 1278 3292 1279
rect 3470 1283 3476 1284
rect 3470 1279 3471 1283
rect 3475 1279 3476 1283
rect 3470 1278 3476 1279
rect 3662 1283 3668 1284
rect 3662 1279 3663 1283
rect 3667 1279 3668 1283
rect 3662 1278 3668 1279
rect 3838 1283 3844 1284
rect 3838 1279 3839 1283
rect 3843 1279 3844 1283
rect 3942 1280 3943 1284
rect 3947 1280 3948 1284
rect 3942 1279 3948 1280
rect 3838 1278 3844 1279
rect 2007 1273 2011 1274
rect 112 1253 114 1273
rect 110 1252 116 1253
rect 440 1252 442 1273
rect 552 1252 554 1273
rect 672 1252 674 1273
rect 800 1252 802 1273
rect 936 1252 938 1273
rect 1080 1252 1082 1273
rect 1232 1252 1234 1273
rect 1392 1252 1394 1273
rect 1552 1252 1554 1273
rect 1720 1252 1722 1273
rect 2008 1253 2010 1273
rect 2046 1267 2052 1268
rect 2046 1263 2047 1267
rect 2051 1263 2052 1267
rect 3942 1267 3948 1268
rect 2046 1262 2052 1263
rect 2246 1264 2252 1265
rect 2006 1252 2012 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 438 1251 444 1252
rect 438 1247 439 1251
rect 443 1247 444 1251
rect 438 1246 444 1247
rect 550 1251 556 1252
rect 550 1247 551 1251
rect 555 1247 556 1251
rect 550 1246 556 1247
rect 670 1251 676 1252
rect 670 1247 671 1251
rect 675 1247 676 1251
rect 670 1246 676 1247
rect 798 1251 804 1252
rect 798 1247 799 1251
rect 803 1247 804 1251
rect 798 1246 804 1247
rect 934 1251 940 1252
rect 934 1247 935 1251
rect 939 1247 940 1251
rect 934 1246 940 1247
rect 1078 1251 1084 1252
rect 1078 1247 1079 1251
rect 1083 1247 1084 1251
rect 1078 1246 1084 1247
rect 1230 1251 1236 1252
rect 1230 1247 1231 1251
rect 1235 1247 1236 1251
rect 1230 1246 1236 1247
rect 1390 1251 1396 1252
rect 1390 1247 1391 1251
rect 1395 1247 1396 1251
rect 1390 1246 1396 1247
rect 1550 1251 1556 1252
rect 1550 1247 1551 1251
rect 1555 1247 1556 1251
rect 1550 1246 1556 1247
rect 1718 1251 1724 1252
rect 1718 1247 1719 1251
rect 1723 1247 1724 1251
rect 2006 1248 2007 1252
rect 2011 1248 2012 1252
rect 2006 1247 2012 1248
rect 1718 1246 1724 1247
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 2006 1235 2012 1236
rect 110 1230 116 1231
rect 438 1232 444 1233
rect 112 1203 114 1230
rect 438 1228 439 1232
rect 443 1228 444 1232
rect 438 1227 444 1228
rect 550 1232 556 1233
rect 550 1228 551 1232
rect 555 1228 556 1232
rect 550 1227 556 1228
rect 670 1232 676 1233
rect 670 1228 671 1232
rect 675 1228 676 1232
rect 670 1227 676 1228
rect 798 1232 804 1233
rect 798 1228 799 1232
rect 803 1228 804 1232
rect 798 1227 804 1228
rect 934 1232 940 1233
rect 934 1228 935 1232
rect 939 1228 940 1232
rect 934 1227 940 1228
rect 1078 1232 1084 1233
rect 1078 1228 1079 1232
rect 1083 1228 1084 1232
rect 1078 1227 1084 1228
rect 1230 1232 1236 1233
rect 1230 1228 1231 1232
rect 1235 1228 1236 1232
rect 1230 1227 1236 1228
rect 1390 1232 1396 1233
rect 1390 1228 1391 1232
rect 1395 1228 1396 1232
rect 1390 1227 1396 1228
rect 1550 1232 1556 1233
rect 1550 1228 1551 1232
rect 1555 1228 1556 1232
rect 1550 1227 1556 1228
rect 1718 1232 1724 1233
rect 1718 1228 1719 1232
rect 1723 1228 1724 1232
rect 2006 1231 2007 1235
rect 2011 1231 2012 1235
rect 2048 1231 2050 1262
rect 2246 1260 2247 1264
rect 2251 1260 2252 1264
rect 2246 1259 2252 1260
rect 2374 1264 2380 1265
rect 2374 1260 2375 1264
rect 2379 1260 2380 1264
rect 2374 1259 2380 1260
rect 2510 1264 2516 1265
rect 2510 1260 2511 1264
rect 2515 1260 2516 1264
rect 2510 1259 2516 1260
rect 2646 1264 2652 1265
rect 2646 1260 2647 1264
rect 2651 1260 2652 1264
rect 2646 1259 2652 1260
rect 2790 1264 2796 1265
rect 2790 1260 2791 1264
rect 2795 1260 2796 1264
rect 2790 1259 2796 1260
rect 2942 1264 2948 1265
rect 2942 1260 2943 1264
rect 2947 1260 2948 1264
rect 2942 1259 2948 1260
rect 3110 1264 3116 1265
rect 3110 1260 3111 1264
rect 3115 1260 3116 1264
rect 3110 1259 3116 1260
rect 3286 1264 3292 1265
rect 3286 1260 3287 1264
rect 3291 1260 3292 1264
rect 3286 1259 3292 1260
rect 3470 1264 3476 1265
rect 3470 1260 3471 1264
rect 3475 1260 3476 1264
rect 3470 1259 3476 1260
rect 3662 1264 3668 1265
rect 3662 1260 3663 1264
rect 3667 1260 3668 1264
rect 3662 1259 3668 1260
rect 3838 1264 3844 1265
rect 3838 1260 3839 1264
rect 3843 1260 3844 1264
rect 3942 1263 3943 1267
rect 3947 1263 3948 1267
rect 3942 1262 3948 1263
rect 3838 1259 3844 1260
rect 2248 1231 2250 1259
rect 2376 1231 2378 1259
rect 2512 1231 2514 1259
rect 2648 1231 2650 1259
rect 2792 1231 2794 1259
rect 2944 1231 2946 1259
rect 3112 1231 3114 1259
rect 3288 1231 3290 1259
rect 3472 1231 3474 1259
rect 3664 1231 3666 1259
rect 3840 1231 3842 1259
rect 3944 1231 3946 1262
rect 2006 1230 2012 1231
rect 2047 1230 2051 1231
rect 1718 1227 1724 1228
rect 440 1203 442 1227
rect 552 1203 554 1227
rect 672 1203 674 1227
rect 800 1203 802 1227
rect 936 1203 938 1227
rect 1080 1203 1082 1227
rect 1232 1203 1234 1227
rect 1392 1203 1394 1227
rect 1552 1203 1554 1227
rect 1720 1203 1722 1227
rect 2008 1203 2010 1230
rect 2047 1225 2051 1226
rect 2071 1230 2075 1231
rect 2071 1225 2075 1226
rect 2183 1230 2187 1231
rect 2183 1225 2187 1226
rect 2247 1230 2251 1231
rect 2247 1225 2251 1226
rect 2303 1230 2307 1231
rect 2303 1225 2307 1226
rect 2375 1230 2379 1231
rect 2375 1225 2379 1226
rect 2431 1230 2435 1231
rect 2431 1225 2435 1226
rect 2511 1230 2515 1231
rect 2511 1225 2515 1226
rect 2559 1230 2563 1231
rect 2559 1225 2563 1226
rect 2647 1230 2651 1231
rect 2647 1225 2651 1226
rect 2711 1230 2715 1231
rect 2711 1225 2715 1226
rect 2791 1230 2795 1231
rect 2791 1225 2795 1226
rect 2887 1230 2891 1231
rect 2887 1225 2891 1226
rect 2943 1230 2947 1231
rect 2943 1225 2947 1226
rect 3087 1230 3091 1231
rect 3087 1225 3091 1226
rect 3111 1230 3115 1231
rect 3111 1225 3115 1226
rect 3287 1230 3291 1231
rect 3287 1225 3291 1226
rect 3311 1230 3315 1231
rect 3311 1225 3315 1226
rect 3471 1230 3475 1231
rect 3471 1225 3475 1226
rect 3543 1230 3547 1231
rect 3543 1225 3547 1226
rect 3663 1230 3667 1231
rect 3663 1225 3667 1226
rect 3783 1230 3787 1231
rect 3783 1225 3787 1226
rect 3839 1230 3843 1231
rect 3839 1225 3843 1226
rect 3943 1230 3947 1231
rect 3943 1225 3947 1226
rect 111 1202 115 1203
rect 111 1197 115 1198
rect 167 1202 171 1203
rect 167 1197 171 1198
rect 303 1202 307 1203
rect 303 1197 307 1198
rect 439 1202 443 1203
rect 439 1197 443 1198
rect 463 1202 467 1203
rect 463 1197 467 1198
rect 551 1202 555 1203
rect 551 1197 555 1198
rect 631 1202 635 1203
rect 631 1197 635 1198
rect 671 1202 675 1203
rect 671 1197 675 1198
rect 799 1202 803 1203
rect 799 1197 803 1198
rect 807 1202 811 1203
rect 807 1197 811 1198
rect 935 1202 939 1203
rect 935 1197 939 1198
rect 983 1202 987 1203
rect 983 1197 987 1198
rect 1079 1202 1083 1203
rect 1079 1197 1083 1198
rect 1159 1202 1163 1203
rect 1159 1197 1163 1198
rect 1231 1202 1235 1203
rect 1231 1197 1235 1198
rect 1335 1202 1339 1203
rect 1335 1197 1339 1198
rect 1391 1202 1395 1203
rect 1391 1197 1395 1198
rect 1511 1202 1515 1203
rect 1511 1197 1515 1198
rect 1551 1202 1555 1203
rect 1551 1197 1555 1198
rect 1695 1202 1699 1203
rect 1695 1197 1699 1198
rect 1719 1202 1723 1203
rect 1719 1197 1723 1198
rect 2007 1202 2011 1203
rect 2048 1198 2050 1225
rect 2072 1201 2074 1225
rect 2184 1201 2186 1225
rect 2304 1201 2306 1225
rect 2432 1201 2434 1225
rect 2560 1201 2562 1225
rect 2712 1201 2714 1225
rect 2888 1201 2890 1225
rect 3088 1201 3090 1225
rect 3312 1201 3314 1225
rect 3544 1201 3546 1225
rect 3784 1201 3786 1225
rect 2070 1200 2076 1201
rect 2007 1197 2011 1198
rect 2046 1197 2052 1198
rect 112 1170 114 1197
rect 168 1173 170 1197
rect 304 1173 306 1197
rect 464 1173 466 1197
rect 632 1173 634 1197
rect 808 1173 810 1197
rect 984 1173 986 1197
rect 1160 1173 1162 1197
rect 1336 1173 1338 1197
rect 1512 1173 1514 1197
rect 1696 1173 1698 1197
rect 166 1172 172 1173
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 166 1168 167 1172
rect 171 1168 172 1172
rect 166 1167 172 1168
rect 302 1172 308 1173
rect 302 1168 303 1172
rect 307 1168 308 1172
rect 302 1167 308 1168
rect 462 1172 468 1173
rect 462 1168 463 1172
rect 467 1168 468 1172
rect 462 1167 468 1168
rect 630 1172 636 1173
rect 630 1168 631 1172
rect 635 1168 636 1172
rect 630 1167 636 1168
rect 806 1172 812 1173
rect 806 1168 807 1172
rect 811 1168 812 1172
rect 806 1167 812 1168
rect 982 1172 988 1173
rect 982 1168 983 1172
rect 987 1168 988 1172
rect 982 1167 988 1168
rect 1158 1172 1164 1173
rect 1158 1168 1159 1172
rect 1163 1168 1164 1172
rect 1158 1167 1164 1168
rect 1334 1172 1340 1173
rect 1334 1168 1335 1172
rect 1339 1168 1340 1172
rect 1334 1167 1340 1168
rect 1510 1172 1516 1173
rect 1510 1168 1511 1172
rect 1515 1168 1516 1172
rect 1510 1167 1516 1168
rect 1694 1172 1700 1173
rect 1694 1168 1695 1172
rect 1699 1168 1700 1172
rect 2008 1170 2010 1197
rect 2046 1193 2047 1197
rect 2051 1193 2052 1197
rect 2070 1196 2071 1200
rect 2075 1196 2076 1200
rect 2070 1195 2076 1196
rect 2182 1200 2188 1201
rect 2182 1196 2183 1200
rect 2187 1196 2188 1200
rect 2182 1195 2188 1196
rect 2302 1200 2308 1201
rect 2302 1196 2303 1200
rect 2307 1196 2308 1200
rect 2302 1195 2308 1196
rect 2430 1200 2436 1201
rect 2430 1196 2431 1200
rect 2435 1196 2436 1200
rect 2430 1195 2436 1196
rect 2558 1200 2564 1201
rect 2558 1196 2559 1200
rect 2563 1196 2564 1200
rect 2558 1195 2564 1196
rect 2710 1200 2716 1201
rect 2710 1196 2711 1200
rect 2715 1196 2716 1200
rect 2710 1195 2716 1196
rect 2886 1200 2892 1201
rect 2886 1196 2887 1200
rect 2891 1196 2892 1200
rect 2886 1195 2892 1196
rect 3086 1200 3092 1201
rect 3086 1196 3087 1200
rect 3091 1196 3092 1200
rect 3086 1195 3092 1196
rect 3310 1200 3316 1201
rect 3310 1196 3311 1200
rect 3315 1196 3316 1200
rect 3310 1195 3316 1196
rect 3542 1200 3548 1201
rect 3542 1196 3543 1200
rect 3547 1196 3548 1200
rect 3542 1195 3548 1196
rect 3782 1200 3788 1201
rect 3782 1196 3783 1200
rect 3787 1196 3788 1200
rect 3944 1198 3946 1225
rect 3782 1195 3788 1196
rect 3942 1197 3948 1198
rect 2046 1192 2052 1193
rect 3942 1193 3943 1197
rect 3947 1193 3948 1197
rect 3942 1192 3948 1193
rect 2070 1181 2076 1182
rect 2046 1180 2052 1181
rect 2046 1176 2047 1180
rect 2051 1176 2052 1180
rect 2070 1177 2071 1181
rect 2075 1177 2076 1181
rect 2070 1176 2076 1177
rect 2182 1181 2188 1182
rect 2182 1177 2183 1181
rect 2187 1177 2188 1181
rect 2182 1176 2188 1177
rect 2302 1181 2308 1182
rect 2302 1177 2303 1181
rect 2307 1177 2308 1181
rect 2302 1176 2308 1177
rect 2430 1181 2436 1182
rect 2430 1177 2431 1181
rect 2435 1177 2436 1181
rect 2430 1176 2436 1177
rect 2558 1181 2564 1182
rect 2558 1177 2559 1181
rect 2563 1177 2564 1181
rect 2558 1176 2564 1177
rect 2710 1181 2716 1182
rect 2710 1177 2711 1181
rect 2715 1177 2716 1181
rect 2710 1176 2716 1177
rect 2886 1181 2892 1182
rect 2886 1177 2887 1181
rect 2891 1177 2892 1181
rect 2886 1176 2892 1177
rect 3086 1181 3092 1182
rect 3086 1177 3087 1181
rect 3091 1177 3092 1181
rect 3086 1176 3092 1177
rect 3310 1181 3316 1182
rect 3310 1177 3311 1181
rect 3315 1177 3316 1181
rect 3310 1176 3316 1177
rect 3542 1181 3548 1182
rect 3542 1177 3543 1181
rect 3547 1177 3548 1181
rect 3542 1176 3548 1177
rect 3782 1181 3788 1182
rect 3782 1177 3783 1181
rect 3787 1177 3788 1181
rect 3782 1176 3788 1177
rect 3942 1180 3948 1181
rect 3942 1176 3943 1180
rect 3947 1176 3948 1180
rect 2046 1175 2052 1176
rect 1694 1167 1700 1168
rect 2006 1169 2012 1170
rect 110 1164 116 1165
rect 2006 1165 2007 1169
rect 2011 1165 2012 1169
rect 2006 1164 2012 1165
rect 166 1153 172 1154
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 166 1149 167 1153
rect 171 1149 172 1153
rect 166 1148 172 1149
rect 302 1153 308 1154
rect 302 1149 303 1153
rect 307 1149 308 1153
rect 302 1148 308 1149
rect 462 1153 468 1154
rect 462 1149 463 1153
rect 467 1149 468 1153
rect 462 1148 468 1149
rect 630 1153 636 1154
rect 630 1149 631 1153
rect 635 1149 636 1153
rect 630 1148 636 1149
rect 806 1153 812 1154
rect 806 1149 807 1153
rect 811 1149 812 1153
rect 806 1148 812 1149
rect 982 1153 988 1154
rect 982 1149 983 1153
rect 987 1149 988 1153
rect 982 1148 988 1149
rect 1158 1153 1164 1154
rect 1158 1149 1159 1153
rect 1163 1149 1164 1153
rect 1158 1148 1164 1149
rect 1334 1153 1340 1154
rect 1334 1149 1335 1153
rect 1339 1149 1340 1153
rect 1334 1148 1340 1149
rect 1510 1153 1516 1154
rect 1510 1149 1511 1153
rect 1515 1149 1516 1153
rect 1510 1148 1516 1149
rect 1694 1153 1700 1154
rect 1694 1149 1695 1153
rect 1699 1149 1700 1153
rect 1694 1148 1700 1149
rect 2006 1152 2012 1153
rect 2006 1148 2007 1152
rect 2011 1148 2012 1152
rect 2048 1151 2050 1175
rect 2072 1151 2074 1176
rect 2184 1151 2186 1176
rect 2304 1151 2306 1176
rect 2432 1151 2434 1176
rect 2560 1151 2562 1176
rect 2712 1151 2714 1176
rect 2888 1151 2890 1176
rect 3088 1151 3090 1176
rect 3312 1151 3314 1176
rect 3544 1151 3546 1176
rect 3784 1151 3786 1176
rect 3942 1175 3948 1176
rect 3944 1151 3946 1175
rect 110 1147 116 1148
rect 112 1123 114 1147
rect 168 1123 170 1148
rect 304 1123 306 1148
rect 464 1123 466 1148
rect 632 1123 634 1148
rect 808 1123 810 1148
rect 984 1123 986 1148
rect 1160 1123 1162 1148
rect 1336 1123 1338 1148
rect 1512 1123 1514 1148
rect 1696 1123 1698 1148
rect 2006 1147 2012 1148
rect 2047 1150 2051 1151
rect 2008 1123 2010 1147
rect 2047 1145 2051 1146
rect 2071 1150 2075 1151
rect 2071 1145 2075 1146
rect 2183 1150 2187 1151
rect 2183 1145 2187 1146
rect 2199 1150 2203 1151
rect 2199 1145 2203 1146
rect 2303 1150 2307 1151
rect 2303 1145 2307 1146
rect 2351 1150 2355 1151
rect 2351 1145 2355 1146
rect 2431 1150 2435 1151
rect 2431 1145 2435 1146
rect 2511 1150 2515 1151
rect 2511 1145 2515 1146
rect 2559 1150 2563 1151
rect 2559 1145 2563 1146
rect 2679 1150 2683 1151
rect 2679 1145 2683 1146
rect 2711 1150 2715 1151
rect 2711 1145 2715 1146
rect 2871 1150 2875 1151
rect 2871 1145 2875 1146
rect 2887 1150 2891 1151
rect 2887 1145 2891 1146
rect 3087 1150 3091 1151
rect 3087 1145 3091 1146
rect 3311 1150 3315 1151
rect 3311 1145 3315 1146
rect 3319 1150 3323 1151
rect 3319 1145 3323 1146
rect 3543 1150 3547 1151
rect 3543 1145 3547 1146
rect 3559 1150 3563 1151
rect 3559 1145 3563 1146
rect 3783 1150 3787 1151
rect 3783 1145 3787 1146
rect 3807 1150 3811 1151
rect 3807 1145 3811 1146
rect 3943 1150 3947 1151
rect 3943 1145 3947 1146
rect 2048 1125 2050 1145
rect 2046 1124 2052 1125
rect 2072 1124 2074 1145
rect 2200 1124 2202 1145
rect 2352 1124 2354 1145
rect 2512 1124 2514 1145
rect 2680 1124 2682 1145
rect 2872 1124 2874 1145
rect 3088 1124 3090 1145
rect 3320 1124 3322 1145
rect 3560 1124 3562 1145
rect 3808 1124 3810 1145
rect 3944 1125 3946 1145
rect 3942 1124 3948 1125
rect 111 1122 115 1123
rect 111 1117 115 1118
rect 135 1122 139 1123
rect 135 1117 139 1118
rect 167 1122 171 1123
rect 167 1117 171 1118
rect 239 1122 243 1123
rect 239 1117 243 1118
rect 303 1122 307 1123
rect 303 1117 307 1118
rect 375 1122 379 1123
rect 375 1117 379 1118
rect 463 1122 467 1123
rect 463 1117 467 1118
rect 527 1122 531 1123
rect 527 1117 531 1118
rect 631 1122 635 1123
rect 631 1117 635 1118
rect 695 1122 699 1123
rect 695 1117 699 1118
rect 807 1122 811 1123
rect 807 1117 811 1118
rect 863 1122 867 1123
rect 863 1117 867 1118
rect 983 1122 987 1123
rect 983 1117 987 1118
rect 1039 1122 1043 1123
rect 1039 1117 1043 1118
rect 1159 1122 1163 1123
rect 1159 1117 1163 1118
rect 1215 1122 1219 1123
rect 1215 1117 1219 1118
rect 1335 1122 1339 1123
rect 1335 1117 1339 1118
rect 1391 1122 1395 1123
rect 1391 1117 1395 1118
rect 1511 1122 1515 1123
rect 1511 1117 1515 1118
rect 1567 1122 1571 1123
rect 1567 1117 1571 1118
rect 1695 1122 1699 1123
rect 1695 1117 1699 1118
rect 1743 1122 1747 1123
rect 1743 1117 1747 1118
rect 1903 1122 1907 1123
rect 1903 1117 1907 1118
rect 2007 1122 2011 1123
rect 2046 1120 2047 1124
rect 2051 1120 2052 1124
rect 2046 1119 2052 1120
rect 2070 1123 2076 1124
rect 2070 1119 2071 1123
rect 2075 1119 2076 1123
rect 2070 1118 2076 1119
rect 2198 1123 2204 1124
rect 2198 1119 2199 1123
rect 2203 1119 2204 1123
rect 2198 1118 2204 1119
rect 2350 1123 2356 1124
rect 2350 1119 2351 1123
rect 2355 1119 2356 1123
rect 2350 1118 2356 1119
rect 2510 1123 2516 1124
rect 2510 1119 2511 1123
rect 2515 1119 2516 1123
rect 2510 1118 2516 1119
rect 2678 1123 2684 1124
rect 2678 1119 2679 1123
rect 2683 1119 2684 1123
rect 2678 1118 2684 1119
rect 2870 1123 2876 1124
rect 2870 1119 2871 1123
rect 2875 1119 2876 1123
rect 2870 1118 2876 1119
rect 3086 1123 3092 1124
rect 3086 1119 3087 1123
rect 3091 1119 3092 1123
rect 3086 1118 3092 1119
rect 3318 1123 3324 1124
rect 3318 1119 3319 1123
rect 3323 1119 3324 1123
rect 3318 1118 3324 1119
rect 3558 1123 3564 1124
rect 3558 1119 3559 1123
rect 3563 1119 3564 1123
rect 3558 1118 3564 1119
rect 3806 1123 3812 1124
rect 3806 1119 3807 1123
rect 3811 1119 3812 1123
rect 3942 1120 3943 1124
rect 3947 1120 3948 1124
rect 3942 1119 3948 1120
rect 3806 1118 3812 1119
rect 2007 1117 2011 1118
rect 112 1097 114 1117
rect 110 1096 116 1097
rect 136 1096 138 1117
rect 240 1096 242 1117
rect 376 1096 378 1117
rect 528 1096 530 1117
rect 696 1096 698 1117
rect 864 1096 866 1117
rect 1040 1096 1042 1117
rect 1216 1096 1218 1117
rect 1392 1096 1394 1117
rect 1568 1096 1570 1117
rect 1744 1096 1746 1117
rect 1904 1096 1906 1117
rect 2008 1097 2010 1117
rect 2046 1107 2052 1108
rect 2046 1103 2047 1107
rect 2051 1103 2052 1107
rect 3942 1107 3948 1108
rect 2046 1102 2052 1103
rect 2070 1104 2076 1105
rect 2006 1096 2012 1097
rect 110 1092 111 1096
rect 115 1092 116 1096
rect 110 1091 116 1092
rect 134 1095 140 1096
rect 134 1091 135 1095
rect 139 1091 140 1095
rect 134 1090 140 1091
rect 238 1095 244 1096
rect 238 1091 239 1095
rect 243 1091 244 1095
rect 238 1090 244 1091
rect 374 1095 380 1096
rect 374 1091 375 1095
rect 379 1091 380 1095
rect 374 1090 380 1091
rect 526 1095 532 1096
rect 526 1091 527 1095
rect 531 1091 532 1095
rect 526 1090 532 1091
rect 694 1095 700 1096
rect 694 1091 695 1095
rect 699 1091 700 1095
rect 694 1090 700 1091
rect 862 1095 868 1096
rect 862 1091 863 1095
rect 867 1091 868 1095
rect 862 1090 868 1091
rect 1038 1095 1044 1096
rect 1038 1091 1039 1095
rect 1043 1091 1044 1095
rect 1038 1090 1044 1091
rect 1214 1095 1220 1096
rect 1214 1091 1215 1095
rect 1219 1091 1220 1095
rect 1214 1090 1220 1091
rect 1390 1095 1396 1096
rect 1390 1091 1391 1095
rect 1395 1091 1396 1095
rect 1390 1090 1396 1091
rect 1566 1095 1572 1096
rect 1566 1091 1567 1095
rect 1571 1091 1572 1095
rect 1566 1090 1572 1091
rect 1742 1095 1748 1096
rect 1742 1091 1743 1095
rect 1747 1091 1748 1095
rect 1742 1090 1748 1091
rect 1902 1095 1908 1096
rect 1902 1091 1903 1095
rect 1907 1091 1908 1095
rect 2006 1092 2007 1096
rect 2011 1092 2012 1096
rect 2006 1091 2012 1092
rect 1902 1090 1908 1091
rect 110 1079 116 1080
rect 110 1075 111 1079
rect 115 1075 116 1079
rect 2006 1079 2012 1080
rect 110 1074 116 1075
rect 134 1076 140 1077
rect 112 1047 114 1074
rect 134 1072 135 1076
rect 139 1072 140 1076
rect 134 1071 140 1072
rect 238 1076 244 1077
rect 238 1072 239 1076
rect 243 1072 244 1076
rect 238 1071 244 1072
rect 374 1076 380 1077
rect 374 1072 375 1076
rect 379 1072 380 1076
rect 374 1071 380 1072
rect 526 1076 532 1077
rect 526 1072 527 1076
rect 531 1072 532 1076
rect 526 1071 532 1072
rect 694 1076 700 1077
rect 694 1072 695 1076
rect 699 1072 700 1076
rect 694 1071 700 1072
rect 862 1076 868 1077
rect 862 1072 863 1076
rect 867 1072 868 1076
rect 862 1071 868 1072
rect 1038 1076 1044 1077
rect 1038 1072 1039 1076
rect 1043 1072 1044 1076
rect 1038 1071 1044 1072
rect 1214 1076 1220 1077
rect 1214 1072 1215 1076
rect 1219 1072 1220 1076
rect 1214 1071 1220 1072
rect 1390 1076 1396 1077
rect 1390 1072 1391 1076
rect 1395 1072 1396 1076
rect 1390 1071 1396 1072
rect 1566 1076 1572 1077
rect 1566 1072 1567 1076
rect 1571 1072 1572 1076
rect 1566 1071 1572 1072
rect 1742 1076 1748 1077
rect 1742 1072 1743 1076
rect 1747 1072 1748 1076
rect 1742 1071 1748 1072
rect 1902 1076 1908 1077
rect 1902 1072 1903 1076
rect 1907 1072 1908 1076
rect 2006 1075 2007 1079
rect 2011 1075 2012 1079
rect 2006 1074 2012 1075
rect 1902 1071 1908 1072
rect 136 1047 138 1071
rect 240 1047 242 1071
rect 376 1047 378 1071
rect 528 1047 530 1071
rect 696 1047 698 1071
rect 864 1047 866 1071
rect 1040 1047 1042 1071
rect 1216 1047 1218 1071
rect 1392 1047 1394 1071
rect 1568 1047 1570 1071
rect 1744 1047 1746 1071
rect 1904 1047 1906 1071
rect 2008 1047 2010 1074
rect 2048 1063 2050 1102
rect 2070 1100 2071 1104
rect 2075 1100 2076 1104
rect 2070 1099 2076 1100
rect 2198 1104 2204 1105
rect 2198 1100 2199 1104
rect 2203 1100 2204 1104
rect 2198 1099 2204 1100
rect 2350 1104 2356 1105
rect 2350 1100 2351 1104
rect 2355 1100 2356 1104
rect 2350 1099 2356 1100
rect 2510 1104 2516 1105
rect 2510 1100 2511 1104
rect 2515 1100 2516 1104
rect 2510 1099 2516 1100
rect 2678 1104 2684 1105
rect 2678 1100 2679 1104
rect 2683 1100 2684 1104
rect 2678 1099 2684 1100
rect 2870 1104 2876 1105
rect 2870 1100 2871 1104
rect 2875 1100 2876 1104
rect 2870 1099 2876 1100
rect 3086 1104 3092 1105
rect 3086 1100 3087 1104
rect 3091 1100 3092 1104
rect 3086 1099 3092 1100
rect 3318 1104 3324 1105
rect 3318 1100 3319 1104
rect 3323 1100 3324 1104
rect 3318 1099 3324 1100
rect 3558 1104 3564 1105
rect 3558 1100 3559 1104
rect 3563 1100 3564 1104
rect 3558 1099 3564 1100
rect 3806 1104 3812 1105
rect 3806 1100 3807 1104
rect 3811 1100 3812 1104
rect 3942 1103 3943 1107
rect 3947 1103 3948 1107
rect 3942 1102 3948 1103
rect 3806 1099 3812 1100
rect 2072 1063 2074 1099
rect 2200 1063 2202 1099
rect 2352 1063 2354 1099
rect 2512 1063 2514 1099
rect 2680 1063 2682 1099
rect 2872 1063 2874 1099
rect 3088 1063 3090 1099
rect 3320 1063 3322 1099
rect 3560 1063 3562 1099
rect 3808 1063 3810 1099
rect 3944 1063 3946 1102
rect 2047 1062 2051 1063
rect 2047 1057 2051 1058
rect 2071 1062 2075 1063
rect 2071 1057 2075 1058
rect 2199 1062 2203 1063
rect 2199 1057 2203 1058
rect 2263 1062 2267 1063
rect 2263 1057 2267 1058
rect 2351 1062 2355 1063
rect 2351 1057 2355 1058
rect 2487 1062 2491 1063
rect 2487 1057 2491 1058
rect 2511 1062 2515 1063
rect 2511 1057 2515 1058
rect 2679 1062 2683 1063
rect 2679 1057 2683 1058
rect 2703 1062 2707 1063
rect 2703 1057 2707 1058
rect 2871 1062 2875 1063
rect 2871 1057 2875 1058
rect 2919 1062 2923 1063
rect 2919 1057 2923 1058
rect 3087 1062 3091 1063
rect 3087 1057 3091 1058
rect 3119 1062 3123 1063
rect 3119 1057 3123 1058
rect 3311 1062 3315 1063
rect 3311 1057 3315 1058
rect 3319 1062 3323 1063
rect 3319 1057 3323 1058
rect 3495 1062 3499 1063
rect 3495 1057 3499 1058
rect 3559 1062 3563 1063
rect 3559 1057 3563 1058
rect 3679 1062 3683 1063
rect 3679 1057 3683 1058
rect 3807 1062 3811 1063
rect 3807 1057 3811 1058
rect 3839 1062 3843 1063
rect 3839 1057 3843 1058
rect 3943 1062 3947 1063
rect 3943 1057 3947 1058
rect 111 1046 115 1047
rect 111 1041 115 1042
rect 135 1046 139 1047
rect 135 1041 139 1042
rect 239 1046 243 1047
rect 239 1041 243 1042
rect 287 1046 291 1047
rect 287 1041 291 1042
rect 375 1046 379 1047
rect 375 1041 379 1042
rect 471 1046 475 1047
rect 471 1041 475 1042
rect 527 1046 531 1047
rect 527 1041 531 1042
rect 655 1046 659 1047
rect 655 1041 659 1042
rect 695 1046 699 1047
rect 695 1041 699 1042
rect 839 1046 843 1047
rect 839 1041 843 1042
rect 863 1046 867 1047
rect 863 1041 867 1042
rect 1015 1046 1019 1047
rect 1015 1041 1019 1042
rect 1039 1046 1043 1047
rect 1039 1041 1043 1042
rect 1199 1046 1203 1047
rect 1199 1041 1203 1042
rect 1215 1046 1219 1047
rect 1215 1041 1219 1042
rect 1383 1046 1387 1047
rect 1383 1041 1387 1042
rect 1391 1046 1395 1047
rect 1391 1041 1395 1042
rect 1567 1046 1571 1047
rect 1567 1041 1571 1042
rect 1743 1046 1747 1047
rect 1743 1041 1747 1042
rect 1903 1046 1907 1047
rect 1903 1041 1907 1042
rect 2007 1046 2011 1047
rect 2007 1041 2011 1042
rect 112 1014 114 1041
rect 136 1017 138 1041
rect 288 1017 290 1041
rect 472 1017 474 1041
rect 656 1017 658 1041
rect 840 1017 842 1041
rect 1016 1017 1018 1041
rect 1200 1017 1202 1041
rect 1384 1017 1386 1041
rect 1568 1017 1570 1041
rect 134 1016 140 1017
rect 110 1013 116 1014
rect 110 1009 111 1013
rect 115 1009 116 1013
rect 134 1012 135 1016
rect 139 1012 140 1016
rect 134 1011 140 1012
rect 286 1016 292 1017
rect 286 1012 287 1016
rect 291 1012 292 1016
rect 286 1011 292 1012
rect 470 1016 476 1017
rect 470 1012 471 1016
rect 475 1012 476 1016
rect 470 1011 476 1012
rect 654 1016 660 1017
rect 654 1012 655 1016
rect 659 1012 660 1016
rect 654 1011 660 1012
rect 838 1016 844 1017
rect 838 1012 839 1016
rect 843 1012 844 1016
rect 838 1011 844 1012
rect 1014 1016 1020 1017
rect 1014 1012 1015 1016
rect 1019 1012 1020 1016
rect 1014 1011 1020 1012
rect 1198 1016 1204 1017
rect 1198 1012 1199 1016
rect 1203 1012 1204 1016
rect 1198 1011 1204 1012
rect 1382 1016 1388 1017
rect 1382 1012 1383 1016
rect 1387 1012 1388 1016
rect 1382 1011 1388 1012
rect 1566 1016 1572 1017
rect 1566 1012 1567 1016
rect 1571 1012 1572 1016
rect 2008 1014 2010 1041
rect 2048 1030 2050 1057
rect 2072 1033 2074 1057
rect 2264 1033 2266 1057
rect 2488 1033 2490 1057
rect 2704 1033 2706 1057
rect 2920 1033 2922 1057
rect 3120 1033 3122 1057
rect 3312 1033 3314 1057
rect 3496 1033 3498 1057
rect 3680 1033 3682 1057
rect 3840 1033 3842 1057
rect 2070 1032 2076 1033
rect 2046 1029 2052 1030
rect 2046 1025 2047 1029
rect 2051 1025 2052 1029
rect 2070 1028 2071 1032
rect 2075 1028 2076 1032
rect 2070 1027 2076 1028
rect 2262 1032 2268 1033
rect 2262 1028 2263 1032
rect 2267 1028 2268 1032
rect 2262 1027 2268 1028
rect 2486 1032 2492 1033
rect 2486 1028 2487 1032
rect 2491 1028 2492 1032
rect 2486 1027 2492 1028
rect 2702 1032 2708 1033
rect 2702 1028 2703 1032
rect 2707 1028 2708 1032
rect 2702 1027 2708 1028
rect 2918 1032 2924 1033
rect 2918 1028 2919 1032
rect 2923 1028 2924 1032
rect 2918 1027 2924 1028
rect 3118 1032 3124 1033
rect 3118 1028 3119 1032
rect 3123 1028 3124 1032
rect 3118 1027 3124 1028
rect 3310 1032 3316 1033
rect 3310 1028 3311 1032
rect 3315 1028 3316 1032
rect 3310 1027 3316 1028
rect 3494 1032 3500 1033
rect 3494 1028 3495 1032
rect 3499 1028 3500 1032
rect 3494 1027 3500 1028
rect 3678 1032 3684 1033
rect 3678 1028 3679 1032
rect 3683 1028 3684 1032
rect 3678 1027 3684 1028
rect 3838 1032 3844 1033
rect 3838 1028 3839 1032
rect 3843 1028 3844 1032
rect 3944 1030 3946 1057
rect 3838 1027 3844 1028
rect 3942 1029 3948 1030
rect 2046 1024 2052 1025
rect 3942 1025 3943 1029
rect 3947 1025 3948 1029
rect 3942 1024 3948 1025
rect 1566 1011 1572 1012
rect 2006 1013 2012 1014
rect 2070 1013 2076 1014
rect 110 1008 116 1009
rect 2006 1009 2007 1013
rect 2011 1009 2012 1013
rect 2006 1008 2012 1009
rect 2046 1012 2052 1013
rect 2046 1008 2047 1012
rect 2051 1008 2052 1012
rect 2070 1009 2071 1013
rect 2075 1009 2076 1013
rect 2070 1008 2076 1009
rect 2262 1013 2268 1014
rect 2262 1009 2263 1013
rect 2267 1009 2268 1013
rect 2262 1008 2268 1009
rect 2486 1013 2492 1014
rect 2486 1009 2487 1013
rect 2491 1009 2492 1013
rect 2486 1008 2492 1009
rect 2702 1013 2708 1014
rect 2702 1009 2703 1013
rect 2707 1009 2708 1013
rect 2702 1008 2708 1009
rect 2918 1013 2924 1014
rect 2918 1009 2919 1013
rect 2923 1009 2924 1013
rect 2918 1008 2924 1009
rect 3118 1013 3124 1014
rect 3118 1009 3119 1013
rect 3123 1009 3124 1013
rect 3118 1008 3124 1009
rect 3310 1013 3316 1014
rect 3310 1009 3311 1013
rect 3315 1009 3316 1013
rect 3310 1008 3316 1009
rect 3494 1013 3500 1014
rect 3494 1009 3495 1013
rect 3499 1009 3500 1013
rect 3494 1008 3500 1009
rect 3678 1013 3684 1014
rect 3678 1009 3679 1013
rect 3683 1009 3684 1013
rect 3678 1008 3684 1009
rect 3838 1013 3844 1014
rect 3838 1009 3839 1013
rect 3843 1009 3844 1013
rect 3838 1008 3844 1009
rect 3942 1012 3948 1013
rect 3942 1008 3943 1012
rect 3947 1008 3948 1012
rect 2046 1007 2052 1008
rect 134 997 140 998
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 134 993 135 997
rect 139 993 140 997
rect 134 992 140 993
rect 286 997 292 998
rect 286 993 287 997
rect 291 993 292 997
rect 286 992 292 993
rect 470 997 476 998
rect 470 993 471 997
rect 475 993 476 997
rect 470 992 476 993
rect 654 997 660 998
rect 654 993 655 997
rect 659 993 660 997
rect 654 992 660 993
rect 838 997 844 998
rect 838 993 839 997
rect 843 993 844 997
rect 838 992 844 993
rect 1014 997 1020 998
rect 1014 993 1015 997
rect 1019 993 1020 997
rect 1014 992 1020 993
rect 1198 997 1204 998
rect 1198 993 1199 997
rect 1203 993 1204 997
rect 1198 992 1204 993
rect 1382 997 1388 998
rect 1382 993 1383 997
rect 1387 993 1388 997
rect 1382 992 1388 993
rect 1566 997 1572 998
rect 1566 993 1567 997
rect 1571 993 1572 997
rect 1566 992 1572 993
rect 2006 996 2012 997
rect 2006 992 2007 996
rect 2011 992 2012 996
rect 110 991 116 992
rect 112 967 114 991
rect 136 967 138 992
rect 288 967 290 992
rect 472 967 474 992
rect 656 967 658 992
rect 840 967 842 992
rect 1016 967 1018 992
rect 1200 967 1202 992
rect 1384 967 1386 992
rect 1568 967 1570 992
rect 2006 991 2012 992
rect 2008 967 2010 991
rect 2048 983 2050 1007
rect 2072 983 2074 1008
rect 2264 983 2266 1008
rect 2488 983 2490 1008
rect 2704 983 2706 1008
rect 2920 983 2922 1008
rect 3120 983 3122 1008
rect 3312 983 3314 1008
rect 3496 983 3498 1008
rect 3680 983 3682 1008
rect 3840 983 3842 1008
rect 3942 1007 3948 1008
rect 3944 983 3946 1007
rect 2047 982 2051 983
rect 2047 977 2051 978
rect 2071 982 2075 983
rect 2071 977 2075 978
rect 2263 982 2267 983
rect 2263 977 2267 978
rect 2303 982 2307 983
rect 2303 977 2307 978
rect 2455 982 2459 983
rect 2455 977 2459 978
rect 2487 982 2491 983
rect 2487 977 2491 978
rect 2615 982 2619 983
rect 2615 977 2619 978
rect 2703 982 2707 983
rect 2703 977 2707 978
rect 2783 982 2787 983
rect 2783 977 2787 978
rect 2919 982 2923 983
rect 2919 977 2923 978
rect 2951 982 2955 983
rect 2951 977 2955 978
rect 3111 982 3115 983
rect 3111 977 3115 978
rect 3119 982 3123 983
rect 3119 977 3123 978
rect 3263 982 3267 983
rect 3263 977 3267 978
rect 3311 982 3315 983
rect 3311 977 3315 978
rect 3415 982 3419 983
rect 3415 977 3419 978
rect 3495 982 3499 983
rect 3495 977 3499 978
rect 3559 982 3563 983
rect 3559 977 3563 978
rect 3679 982 3683 983
rect 3679 977 3683 978
rect 3711 982 3715 983
rect 3711 977 3715 978
rect 3839 982 3843 983
rect 3839 977 3843 978
rect 3943 982 3947 983
rect 3943 977 3947 978
rect 111 966 115 967
rect 111 961 115 962
rect 135 966 139 967
rect 135 961 139 962
rect 287 966 291 967
rect 287 961 291 962
rect 295 966 299 967
rect 295 961 299 962
rect 471 966 475 967
rect 471 961 475 962
rect 639 966 643 967
rect 639 961 643 962
rect 655 966 659 967
rect 655 961 659 962
rect 799 966 803 967
rect 799 961 803 962
rect 839 966 843 967
rect 839 961 843 962
rect 951 966 955 967
rect 951 961 955 962
rect 1015 966 1019 967
rect 1015 961 1019 962
rect 1087 966 1091 967
rect 1087 961 1091 962
rect 1199 966 1203 967
rect 1199 961 1203 962
rect 1223 966 1227 967
rect 1223 961 1227 962
rect 1359 966 1363 967
rect 1359 961 1363 962
rect 1383 966 1387 967
rect 1383 961 1387 962
rect 1495 966 1499 967
rect 1495 961 1499 962
rect 1567 966 1571 967
rect 1567 961 1571 962
rect 2007 966 2011 967
rect 2007 961 2011 962
rect 112 941 114 961
rect 110 940 116 941
rect 136 940 138 961
rect 296 940 298 961
rect 472 940 474 961
rect 640 940 642 961
rect 800 940 802 961
rect 952 940 954 961
rect 1088 940 1090 961
rect 1224 940 1226 961
rect 1360 940 1362 961
rect 1496 940 1498 961
rect 2008 941 2010 961
rect 2048 957 2050 977
rect 2046 956 2052 957
rect 2304 956 2306 977
rect 2456 956 2458 977
rect 2616 956 2618 977
rect 2784 956 2786 977
rect 2952 956 2954 977
rect 3112 956 3114 977
rect 3264 956 3266 977
rect 3416 956 3418 977
rect 3560 956 3562 977
rect 3712 956 3714 977
rect 3840 956 3842 977
rect 3944 957 3946 977
rect 3942 956 3948 957
rect 2046 952 2047 956
rect 2051 952 2052 956
rect 2046 951 2052 952
rect 2302 955 2308 956
rect 2302 951 2303 955
rect 2307 951 2308 955
rect 2302 950 2308 951
rect 2454 955 2460 956
rect 2454 951 2455 955
rect 2459 951 2460 955
rect 2454 950 2460 951
rect 2614 955 2620 956
rect 2614 951 2615 955
rect 2619 951 2620 955
rect 2614 950 2620 951
rect 2782 955 2788 956
rect 2782 951 2783 955
rect 2787 951 2788 955
rect 2782 950 2788 951
rect 2950 955 2956 956
rect 2950 951 2951 955
rect 2955 951 2956 955
rect 2950 950 2956 951
rect 3110 955 3116 956
rect 3110 951 3111 955
rect 3115 951 3116 955
rect 3110 950 3116 951
rect 3262 955 3268 956
rect 3262 951 3263 955
rect 3267 951 3268 955
rect 3262 950 3268 951
rect 3414 955 3420 956
rect 3414 951 3415 955
rect 3419 951 3420 955
rect 3414 950 3420 951
rect 3558 955 3564 956
rect 3558 951 3559 955
rect 3563 951 3564 955
rect 3558 950 3564 951
rect 3710 955 3716 956
rect 3710 951 3711 955
rect 3715 951 3716 955
rect 3710 950 3716 951
rect 3838 955 3844 956
rect 3838 951 3839 955
rect 3843 951 3844 955
rect 3942 952 3943 956
rect 3947 952 3948 956
rect 3942 951 3948 952
rect 3838 950 3844 951
rect 2006 940 2012 941
rect 110 936 111 940
rect 115 936 116 940
rect 110 935 116 936
rect 134 939 140 940
rect 134 935 135 939
rect 139 935 140 939
rect 134 934 140 935
rect 294 939 300 940
rect 294 935 295 939
rect 299 935 300 939
rect 294 934 300 935
rect 470 939 476 940
rect 470 935 471 939
rect 475 935 476 939
rect 470 934 476 935
rect 638 939 644 940
rect 638 935 639 939
rect 643 935 644 939
rect 638 934 644 935
rect 798 939 804 940
rect 798 935 799 939
rect 803 935 804 939
rect 798 934 804 935
rect 950 939 956 940
rect 950 935 951 939
rect 955 935 956 939
rect 950 934 956 935
rect 1086 939 1092 940
rect 1086 935 1087 939
rect 1091 935 1092 939
rect 1086 934 1092 935
rect 1222 939 1228 940
rect 1222 935 1223 939
rect 1227 935 1228 939
rect 1222 934 1228 935
rect 1358 939 1364 940
rect 1358 935 1359 939
rect 1363 935 1364 939
rect 1358 934 1364 935
rect 1494 939 1500 940
rect 1494 935 1495 939
rect 1499 935 1500 939
rect 2006 936 2007 940
rect 2011 936 2012 940
rect 2006 935 2012 936
rect 2046 939 2052 940
rect 2046 935 2047 939
rect 2051 935 2052 939
rect 3942 939 3948 940
rect 1494 934 1500 935
rect 2046 934 2052 935
rect 2302 936 2308 937
rect 110 923 116 924
rect 110 919 111 923
rect 115 919 116 923
rect 2006 923 2012 924
rect 110 918 116 919
rect 134 920 140 921
rect 112 891 114 918
rect 134 916 135 920
rect 139 916 140 920
rect 134 915 140 916
rect 294 920 300 921
rect 294 916 295 920
rect 299 916 300 920
rect 294 915 300 916
rect 470 920 476 921
rect 470 916 471 920
rect 475 916 476 920
rect 470 915 476 916
rect 638 920 644 921
rect 638 916 639 920
rect 643 916 644 920
rect 638 915 644 916
rect 798 920 804 921
rect 798 916 799 920
rect 803 916 804 920
rect 798 915 804 916
rect 950 920 956 921
rect 950 916 951 920
rect 955 916 956 920
rect 950 915 956 916
rect 1086 920 1092 921
rect 1086 916 1087 920
rect 1091 916 1092 920
rect 1086 915 1092 916
rect 1222 920 1228 921
rect 1222 916 1223 920
rect 1227 916 1228 920
rect 1222 915 1228 916
rect 1358 920 1364 921
rect 1358 916 1359 920
rect 1363 916 1364 920
rect 1358 915 1364 916
rect 1494 920 1500 921
rect 1494 916 1495 920
rect 1499 916 1500 920
rect 2006 919 2007 923
rect 2011 919 2012 923
rect 2006 918 2012 919
rect 1494 915 1500 916
rect 136 891 138 915
rect 296 891 298 915
rect 472 891 474 915
rect 640 891 642 915
rect 800 891 802 915
rect 952 891 954 915
rect 1088 891 1090 915
rect 1224 891 1226 915
rect 1360 891 1362 915
rect 1496 891 1498 915
rect 2008 891 2010 918
rect 2048 903 2050 934
rect 2302 932 2303 936
rect 2307 932 2308 936
rect 2302 931 2308 932
rect 2454 936 2460 937
rect 2454 932 2455 936
rect 2459 932 2460 936
rect 2454 931 2460 932
rect 2614 936 2620 937
rect 2614 932 2615 936
rect 2619 932 2620 936
rect 2614 931 2620 932
rect 2782 936 2788 937
rect 2782 932 2783 936
rect 2787 932 2788 936
rect 2782 931 2788 932
rect 2950 936 2956 937
rect 2950 932 2951 936
rect 2955 932 2956 936
rect 2950 931 2956 932
rect 3110 936 3116 937
rect 3110 932 3111 936
rect 3115 932 3116 936
rect 3110 931 3116 932
rect 3262 936 3268 937
rect 3262 932 3263 936
rect 3267 932 3268 936
rect 3262 931 3268 932
rect 3414 936 3420 937
rect 3414 932 3415 936
rect 3419 932 3420 936
rect 3414 931 3420 932
rect 3558 936 3564 937
rect 3558 932 3559 936
rect 3563 932 3564 936
rect 3558 931 3564 932
rect 3710 936 3716 937
rect 3710 932 3711 936
rect 3715 932 3716 936
rect 3710 931 3716 932
rect 3838 936 3844 937
rect 3838 932 3839 936
rect 3843 932 3844 936
rect 3942 935 3943 939
rect 3947 935 3948 939
rect 3942 934 3948 935
rect 3838 931 3844 932
rect 2304 903 2306 931
rect 2456 903 2458 931
rect 2616 903 2618 931
rect 2784 903 2786 931
rect 2952 903 2954 931
rect 3112 903 3114 931
rect 3264 903 3266 931
rect 3416 903 3418 931
rect 3560 903 3562 931
rect 3712 903 3714 931
rect 3840 903 3842 931
rect 3944 903 3946 934
rect 2047 902 2051 903
rect 2047 897 2051 898
rect 2303 902 2307 903
rect 2303 897 2307 898
rect 2455 902 2459 903
rect 2455 897 2459 898
rect 2559 902 2563 903
rect 2559 897 2563 898
rect 2615 902 2619 903
rect 2615 897 2619 898
rect 2679 902 2683 903
rect 2679 897 2683 898
rect 2783 902 2787 903
rect 2783 897 2787 898
rect 2807 902 2811 903
rect 2807 897 2811 898
rect 2943 902 2947 903
rect 2943 897 2947 898
rect 2951 902 2955 903
rect 2951 897 2955 898
rect 3079 902 3083 903
rect 3079 897 3083 898
rect 3111 902 3115 903
rect 3111 897 3115 898
rect 3207 902 3211 903
rect 3207 897 3211 898
rect 3263 902 3267 903
rect 3263 897 3267 898
rect 3335 902 3339 903
rect 3335 897 3339 898
rect 3415 902 3419 903
rect 3415 897 3419 898
rect 3463 902 3467 903
rect 3463 897 3467 898
rect 3559 902 3563 903
rect 3559 897 3563 898
rect 3591 902 3595 903
rect 3591 897 3595 898
rect 3711 902 3715 903
rect 3711 897 3715 898
rect 3727 902 3731 903
rect 3727 897 3731 898
rect 3839 902 3843 903
rect 3839 897 3843 898
rect 3943 902 3947 903
rect 3943 897 3947 898
rect 111 890 115 891
rect 111 885 115 886
rect 135 890 139 891
rect 135 885 139 886
rect 159 890 163 891
rect 159 885 163 886
rect 295 890 299 891
rect 295 885 299 886
rect 319 890 323 891
rect 319 885 323 886
rect 471 890 475 891
rect 471 885 475 886
rect 615 890 619 891
rect 615 885 619 886
rect 639 890 643 891
rect 639 885 643 886
rect 751 890 755 891
rect 751 885 755 886
rect 799 890 803 891
rect 799 885 803 886
rect 879 890 883 891
rect 879 885 883 886
rect 951 890 955 891
rect 951 885 955 886
rect 999 890 1003 891
rect 999 885 1003 886
rect 1087 890 1091 891
rect 1087 885 1091 886
rect 1111 890 1115 891
rect 1111 885 1115 886
rect 1223 890 1227 891
rect 1223 885 1227 886
rect 1231 890 1235 891
rect 1231 885 1235 886
rect 1351 890 1355 891
rect 1351 885 1355 886
rect 1359 890 1363 891
rect 1359 885 1363 886
rect 1495 890 1499 891
rect 1495 885 1499 886
rect 2007 890 2011 891
rect 2007 885 2011 886
rect 112 858 114 885
rect 160 861 162 885
rect 320 861 322 885
rect 472 861 474 885
rect 616 861 618 885
rect 752 861 754 885
rect 880 861 882 885
rect 1000 861 1002 885
rect 1112 861 1114 885
rect 1232 861 1234 885
rect 1352 861 1354 885
rect 158 860 164 861
rect 110 857 116 858
rect 110 853 111 857
rect 115 853 116 857
rect 158 856 159 860
rect 163 856 164 860
rect 158 855 164 856
rect 318 860 324 861
rect 318 856 319 860
rect 323 856 324 860
rect 318 855 324 856
rect 470 860 476 861
rect 470 856 471 860
rect 475 856 476 860
rect 470 855 476 856
rect 614 860 620 861
rect 614 856 615 860
rect 619 856 620 860
rect 614 855 620 856
rect 750 860 756 861
rect 750 856 751 860
rect 755 856 756 860
rect 750 855 756 856
rect 878 860 884 861
rect 878 856 879 860
rect 883 856 884 860
rect 878 855 884 856
rect 998 860 1004 861
rect 998 856 999 860
rect 1003 856 1004 860
rect 998 855 1004 856
rect 1110 860 1116 861
rect 1110 856 1111 860
rect 1115 856 1116 860
rect 1110 855 1116 856
rect 1230 860 1236 861
rect 1230 856 1231 860
rect 1235 856 1236 860
rect 1230 855 1236 856
rect 1350 860 1356 861
rect 1350 856 1351 860
rect 1355 856 1356 860
rect 2008 858 2010 885
rect 2048 870 2050 897
rect 2560 873 2562 897
rect 2680 873 2682 897
rect 2808 873 2810 897
rect 2944 873 2946 897
rect 3080 873 3082 897
rect 3208 873 3210 897
rect 3336 873 3338 897
rect 3464 873 3466 897
rect 3592 873 3594 897
rect 3728 873 3730 897
rect 3840 873 3842 897
rect 2558 872 2564 873
rect 2046 869 2052 870
rect 2046 865 2047 869
rect 2051 865 2052 869
rect 2558 868 2559 872
rect 2563 868 2564 872
rect 2558 867 2564 868
rect 2678 872 2684 873
rect 2678 868 2679 872
rect 2683 868 2684 872
rect 2678 867 2684 868
rect 2806 872 2812 873
rect 2806 868 2807 872
rect 2811 868 2812 872
rect 2806 867 2812 868
rect 2942 872 2948 873
rect 2942 868 2943 872
rect 2947 868 2948 872
rect 2942 867 2948 868
rect 3078 872 3084 873
rect 3078 868 3079 872
rect 3083 868 3084 872
rect 3078 867 3084 868
rect 3206 872 3212 873
rect 3206 868 3207 872
rect 3211 868 3212 872
rect 3206 867 3212 868
rect 3334 872 3340 873
rect 3334 868 3335 872
rect 3339 868 3340 872
rect 3334 867 3340 868
rect 3462 872 3468 873
rect 3462 868 3463 872
rect 3467 868 3468 872
rect 3462 867 3468 868
rect 3590 872 3596 873
rect 3590 868 3591 872
rect 3595 868 3596 872
rect 3590 867 3596 868
rect 3726 872 3732 873
rect 3726 868 3727 872
rect 3731 868 3732 872
rect 3726 867 3732 868
rect 3838 872 3844 873
rect 3838 868 3839 872
rect 3843 868 3844 872
rect 3944 870 3946 897
rect 3838 867 3844 868
rect 3942 869 3948 870
rect 2046 864 2052 865
rect 3942 865 3943 869
rect 3947 865 3948 869
rect 3942 864 3948 865
rect 1350 855 1356 856
rect 2006 857 2012 858
rect 110 852 116 853
rect 2006 853 2007 857
rect 2011 853 2012 857
rect 2558 853 2564 854
rect 2006 852 2012 853
rect 2046 852 2052 853
rect 2046 848 2047 852
rect 2051 848 2052 852
rect 2558 849 2559 853
rect 2563 849 2564 853
rect 2558 848 2564 849
rect 2678 853 2684 854
rect 2678 849 2679 853
rect 2683 849 2684 853
rect 2678 848 2684 849
rect 2806 853 2812 854
rect 2806 849 2807 853
rect 2811 849 2812 853
rect 2806 848 2812 849
rect 2942 853 2948 854
rect 2942 849 2943 853
rect 2947 849 2948 853
rect 2942 848 2948 849
rect 3078 853 3084 854
rect 3078 849 3079 853
rect 3083 849 3084 853
rect 3078 848 3084 849
rect 3206 853 3212 854
rect 3206 849 3207 853
rect 3211 849 3212 853
rect 3206 848 3212 849
rect 3334 853 3340 854
rect 3334 849 3335 853
rect 3339 849 3340 853
rect 3334 848 3340 849
rect 3462 853 3468 854
rect 3462 849 3463 853
rect 3467 849 3468 853
rect 3462 848 3468 849
rect 3590 853 3596 854
rect 3590 849 3591 853
rect 3595 849 3596 853
rect 3590 848 3596 849
rect 3726 853 3732 854
rect 3726 849 3727 853
rect 3731 849 3732 853
rect 3726 848 3732 849
rect 3838 853 3844 854
rect 3838 849 3839 853
rect 3843 849 3844 853
rect 3838 848 3844 849
rect 3942 852 3948 853
rect 3942 848 3943 852
rect 3947 848 3948 852
rect 2046 847 2052 848
rect 158 841 164 842
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 158 837 159 841
rect 163 837 164 841
rect 158 836 164 837
rect 318 841 324 842
rect 318 837 319 841
rect 323 837 324 841
rect 318 836 324 837
rect 470 841 476 842
rect 470 837 471 841
rect 475 837 476 841
rect 470 836 476 837
rect 614 841 620 842
rect 614 837 615 841
rect 619 837 620 841
rect 614 836 620 837
rect 750 841 756 842
rect 750 837 751 841
rect 755 837 756 841
rect 750 836 756 837
rect 878 841 884 842
rect 878 837 879 841
rect 883 837 884 841
rect 878 836 884 837
rect 998 841 1004 842
rect 998 837 999 841
rect 1003 837 1004 841
rect 998 836 1004 837
rect 1110 841 1116 842
rect 1110 837 1111 841
rect 1115 837 1116 841
rect 1110 836 1116 837
rect 1230 841 1236 842
rect 1230 837 1231 841
rect 1235 837 1236 841
rect 1230 836 1236 837
rect 1350 841 1356 842
rect 1350 837 1351 841
rect 1355 837 1356 841
rect 1350 836 1356 837
rect 2006 840 2012 841
rect 2006 836 2007 840
rect 2011 836 2012 840
rect 110 835 116 836
rect 112 815 114 835
rect 160 815 162 836
rect 320 815 322 836
rect 472 815 474 836
rect 616 815 618 836
rect 752 815 754 836
rect 880 815 882 836
rect 1000 815 1002 836
rect 1112 815 1114 836
rect 1232 815 1234 836
rect 1352 815 1354 836
rect 2006 835 2012 836
rect 2008 815 2010 835
rect 2048 823 2050 847
rect 2560 823 2562 848
rect 2680 823 2682 848
rect 2808 823 2810 848
rect 2944 823 2946 848
rect 3080 823 3082 848
rect 3208 823 3210 848
rect 3336 823 3338 848
rect 3464 823 3466 848
rect 3592 823 3594 848
rect 3728 823 3730 848
rect 3840 823 3842 848
rect 3942 847 3948 848
rect 3944 823 3946 847
rect 2047 822 2051 823
rect 2047 817 2051 818
rect 2335 822 2339 823
rect 2335 817 2339 818
rect 2471 822 2475 823
rect 2471 817 2475 818
rect 2559 822 2563 823
rect 2559 817 2563 818
rect 2615 822 2619 823
rect 2615 817 2619 818
rect 2679 822 2683 823
rect 2679 817 2683 818
rect 2767 822 2771 823
rect 2767 817 2771 818
rect 2807 822 2811 823
rect 2807 817 2811 818
rect 2919 822 2923 823
rect 2919 817 2923 818
rect 2943 822 2947 823
rect 2943 817 2947 818
rect 3079 822 3083 823
rect 3079 817 3083 818
rect 3207 822 3211 823
rect 3207 817 3211 818
rect 3239 822 3243 823
rect 3239 817 3243 818
rect 3335 822 3339 823
rect 3335 817 3339 818
rect 3391 822 3395 823
rect 3391 817 3395 818
rect 3463 822 3467 823
rect 3463 817 3467 818
rect 3543 822 3547 823
rect 3543 817 3547 818
rect 3591 822 3595 823
rect 3591 817 3595 818
rect 3703 822 3707 823
rect 3703 817 3707 818
rect 3727 822 3731 823
rect 3727 817 3731 818
rect 3839 822 3843 823
rect 3839 817 3843 818
rect 3943 822 3947 823
rect 3943 817 3947 818
rect 111 814 115 815
rect 111 809 115 810
rect 159 814 163 815
rect 159 809 163 810
rect 223 814 227 815
rect 223 809 227 810
rect 319 814 323 815
rect 319 809 323 810
rect 383 814 387 815
rect 383 809 387 810
rect 471 814 475 815
rect 471 809 475 810
rect 535 814 539 815
rect 535 809 539 810
rect 615 814 619 815
rect 615 809 619 810
rect 679 814 683 815
rect 679 809 683 810
rect 751 814 755 815
rect 751 809 755 810
rect 815 814 819 815
rect 815 809 819 810
rect 879 814 883 815
rect 879 809 883 810
rect 951 814 955 815
rect 951 809 955 810
rect 999 814 1003 815
rect 999 809 1003 810
rect 1079 814 1083 815
rect 1079 809 1083 810
rect 1111 814 1115 815
rect 1111 809 1115 810
rect 1199 814 1203 815
rect 1199 809 1203 810
rect 1231 814 1235 815
rect 1231 809 1235 810
rect 1327 814 1331 815
rect 1327 809 1331 810
rect 1351 814 1355 815
rect 1351 809 1355 810
rect 1455 814 1459 815
rect 1455 809 1459 810
rect 2007 814 2011 815
rect 2007 809 2011 810
rect 112 789 114 809
rect 110 788 116 789
rect 224 788 226 809
rect 384 788 386 809
rect 536 788 538 809
rect 680 788 682 809
rect 816 788 818 809
rect 952 788 954 809
rect 1080 788 1082 809
rect 1200 788 1202 809
rect 1328 788 1330 809
rect 1456 788 1458 809
rect 2008 789 2010 809
rect 2048 797 2050 817
rect 2046 796 2052 797
rect 2336 796 2338 817
rect 2472 796 2474 817
rect 2616 796 2618 817
rect 2768 796 2770 817
rect 2920 796 2922 817
rect 3080 796 3082 817
rect 3240 796 3242 817
rect 3392 796 3394 817
rect 3544 796 3546 817
rect 3704 796 3706 817
rect 3840 796 3842 817
rect 3944 797 3946 817
rect 3942 796 3948 797
rect 2046 792 2047 796
rect 2051 792 2052 796
rect 2046 791 2052 792
rect 2334 795 2340 796
rect 2334 791 2335 795
rect 2339 791 2340 795
rect 2334 790 2340 791
rect 2470 795 2476 796
rect 2470 791 2471 795
rect 2475 791 2476 795
rect 2470 790 2476 791
rect 2614 795 2620 796
rect 2614 791 2615 795
rect 2619 791 2620 795
rect 2614 790 2620 791
rect 2766 795 2772 796
rect 2766 791 2767 795
rect 2771 791 2772 795
rect 2766 790 2772 791
rect 2918 795 2924 796
rect 2918 791 2919 795
rect 2923 791 2924 795
rect 2918 790 2924 791
rect 3078 795 3084 796
rect 3078 791 3079 795
rect 3083 791 3084 795
rect 3078 790 3084 791
rect 3238 795 3244 796
rect 3238 791 3239 795
rect 3243 791 3244 795
rect 3238 790 3244 791
rect 3390 795 3396 796
rect 3390 791 3391 795
rect 3395 791 3396 795
rect 3390 790 3396 791
rect 3542 795 3548 796
rect 3542 791 3543 795
rect 3547 791 3548 795
rect 3542 790 3548 791
rect 3702 795 3708 796
rect 3702 791 3703 795
rect 3707 791 3708 795
rect 3702 790 3708 791
rect 3838 795 3844 796
rect 3838 791 3839 795
rect 3843 791 3844 795
rect 3942 792 3943 796
rect 3947 792 3948 796
rect 3942 791 3948 792
rect 3838 790 3844 791
rect 2006 788 2012 789
rect 110 784 111 788
rect 115 784 116 788
rect 110 783 116 784
rect 222 787 228 788
rect 222 783 223 787
rect 227 783 228 787
rect 222 782 228 783
rect 382 787 388 788
rect 382 783 383 787
rect 387 783 388 787
rect 382 782 388 783
rect 534 787 540 788
rect 534 783 535 787
rect 539 783 540 787
rect 534 782 540 783
rect 678 787 684 788
rect 678 783 679 787
rect 683 783 684 787
rect 678 782 684 783
rect 814 787 820 788
rect 814 783 815 787
rect 819 783 820 787
rect 814 782 820 783
rect 950 787 956 788
rect 950 783 951 787
rect 955 783 956 787
rect 950 782 956 783
rect 1078 787 1084 788
rect 1078 783 1079 787
rect 1083 783 1084 787
rect 1078 782 1084 783
rect 1198 787 1204 788
rect 1198 783 1199 787
rect 1203 783 1204 787
rect 1198 782 1204 783
rect 1326 787 1332 788
rect 1326 783 1327 787
rect 1331 783 1332 787
rect 1326 782 1332 783
rect 1454 787 1460 788
rect 1454 783 1455 787
rect 1459 783 1460 787
rect 2006 784 2007 788
rect 2011 784 2012 788
rect 2006 783 2012 784
rect 1454 782 1460 783
rect 2046 779 2052 780
rect 2046 775 2047 779
rect 2051 775 2052 779
rect 3942 779 3948 780
rect 2046 774 2052 775
rect 2334 776 2340 777
rect 110 771 116 772
rect 110 767 111 771
rect 115 767 116 771
rect 2006 771 2012 772
rect 110 766 116 767
rect 222 768 228 769
rect 112 735 114 766
rect 222 764 223 768
rect 227 764 228 768
rect 222 763 228 764
rect 382 768 388 769
rect 382 764 383 768
rect 387 764 388 768
rect 382 763 388 764
rect 534 768 540 769
rect 534 764 535 768
rect 539 764 540 768
rect 534 763 540 764
rect 678 768 684 769
rect 678 764 679 768
rect 683 764 684 768
rect 678 763 684 764
rect 814 768 820 769
rect 814 764 815 768
rect 819 764 820 768
rect 814 763 820 764
rect 950 768 956 769
rect 950 764 951 768
rect 955 764 956 768
rect 950 763 956 764
rect 1078 768 1084 769
rect 1078 764 1079 768
rect 1083 764 1084 768
rect 1078 763 1084 764
rect 1198 768 1204 769
rect 1198 764 1199 768
rect 1203 764 1204 768
rect 1198 763 1204 764
rect 1326 768 1332 769
rect 1326 764 1327 768
rect 1331 764 1332 768
rect 1326 763 1332 764
rect 1454 768 1460 769
rect 1454 764 1455 768
rect 1459 764 1460 768
rect 2006 767 2007 771
rect 2011 767 2012 771
rect 2006 766 2012 767
rect 1454 763 1460 764
rect 224 735 226 763
rect 384 735 386 763
rect 536 735 538 763
rect 680 735 682 763
rect 816 735 818 763
rect 952 735 954 763
rect 1080 735 1082 763
rect 1200 735 1202 763
rect 1328 735 1330 763
rect 1456 735 1458 763
rect 2008 735 2010 766
rect 2048 743 2050 774
rect 2334 772 2335 776
rect 2339 772 2340 776
rect 2334 771 2340 772
rect 2470 776 2476 777
rect 2470 772 2471 776
rect 2475 772 2476 776
rect 2470 771 2476 772
rect 2614 776 2620 777
rect 2614 772 2615 776
rect 2619 772 2620 776
rect 2614 771 2620 772
rect 2766 776 2772 777
rect 2766 772 2767 776
rect 2771 772 2772 776
rect 2766 771 2772 772
rect 2918 776 2924 777
rect 2918 772 2919 776
rect 2923 772 2924 776
rect 2918 771 2924 772
rect 3078 776 3084 777
rect 3078 772 3079 776
rect 3083 772 3084 776
rect 3078 771 3084 772
rect 3238 776 3244 777
rect 3238 772 3239 776
rect 3243 772 3244 776
rect 3238 771 3244 772
rect 3390 776 3396 777
rect 3390 772 3391 776
rect 3395 772 3396 776
rect 3390 771 3396 772
rect 3542 776 3548 777
rect 3542 772 3543 776
rect 3547 772 3548 776
rect 3542 771 3548 772
rect 3702 776 3708 777
rect 3702 772 3703 776
rect 3707 772 3708 776
rect 3702 771 3708 772
rect 3838 776 3844 777
rect 3838 772 3839 776
rect 3843 772 3844 776
rect 3942 775 3943 779
rect 3947 775 3948 779
rect 3942 774 3948 775
rect 3838 771 3844 772
rect 2336 743 2338 771
rect 2472 743 2474 771
rect 2616 743 2618 771
rect 2768 743 2770 771
rect 2920 743 2922 771
rect 3080 743 3082 771
rect 3240 743 3242 771
rect 3392 743 3394 771
rect 3544 743 3546 771
rect 3704 743 3706 771
rect 3840 743 3842 771
rect 3944 743 3946 774
rect 2047 742 2051 743
rect 2047 737 2051 738
rect 2071 742 2075 743
rect 2071 737 2075 738
rect 2183 742 2187 743
rect 2183 737 2187 738
rect 2335 742 2339 743
rect 2335 737 2339 738
rect 2471 742 2475 743
rect 2471 737 2475 738
rect 2487 742 2491 743
rect 2487 737 2491 738
rect 2615 742 2619 743
rect 2615 737 2619 738
rect 2639 742 2643 743
rect 2639 737 2643 738
rect 2767 742 2771 743
rect 2767 737 2771 738
rect 2807 742 2811 743
rect 2807 737 2811 738
rect 2919 742 2923 743
rect 2919 737 2923 738
rect 2983 742 2987 743
rect 2983 737 2987 738
rect 3079 742 3083 743
rect 3079 737 3083 738
rect 3167 742 3171 743
rect 3167 737 3171 738
rect 3239 742 3243 743
rect 3239 737 3243 738
rect 3367 742 3371 743
rect 3367 737 3371 738
rect 3391 742 3395 743
rect 3391 737 3395 738
rect 3543 742 3547 743
rect 3543 737 3547 738
rect 3575 742 3579 743
rect 3575 737 3579 738
rect 3703 742 3707 743
rect 3703 737 3707 738
rect 3783 742 3787 743
rect 3783 737 3787 738
rect 3839 742 3843 743
rect 3839 737 3843 738
rect 3943 742 3947 743
rect 3943 737 3947 738
rect 111 734 115 735
rect 111 729 115 730
rect 223 734 227 735
rect 223 729 227 730
rect 311 734 315 735
rect 311 729 315 730
rect 383 734 387 735
rect 383 729 387 730
rect 471 734 475 735
rect 471 729 475 730
rect 535 734 539 735
rect 535 729 539 730
rect 639 734 643 735
rect 639 729 643 730
rect 679 734 683 735
rect 679 729 683 730
rect 807 734 811 735
rect 807 729 811 730
rect 815 734 819 735
rect 815 729 819 730
rect 951 734 955 735
rect 951 729 955 730
rect 975 734 979 735
rect 975 729 979 730
rect 1079 734 1083 735
rect 1079 729 1083 730
rect 1135 734 1139 735
rect 1135 729 1139 730
rect 1199 734 1203 735
rect 1199 729 1203 730
rect 1295 734 1299 735
rect 1295 729 1299 730
rect 1327 734 1331 735
rect 1327 729 1331 730
rect 1455 734 1459 735
rect 1455 729 1459 730
rect 1607 734 1611 735
rect 1607 729 1611 730
rect 1767 734 1771 735
rect 1767 729 1771 730
rect 1903 734 1907 735
rect 1903 729 1907 730
rect 2007 734 2011 735
rect 2007 729 2011 730
rect 112 702 114 729
rect 312 705 314 729
rect 472 705 474 729
rect 640 705 642 729
rect 808 705 810 729
rect 976 705 978 729
rect 1136 705 1138 729
rect 1296 705 1298 729
rect 1456 705 1458 729
rect 1608 705 1610 729
rect 1768 705 1770 729
rect 1904 705 1906 729
rect 310 704 316 705
rect 110 701 116 702
rect 110 697 111 701
rect 115 697 116 701
rect 310 700 311 704
rect 315 700 316 704
rect 310 699 316 700
rect 470 704 476 705
rect 470 700 471 704
rect 475 700 476 704
rect 470 699 476 700
rect 638 704 644 705
rect 638 700 639 704
rect 643 700 644 704
rect 638 699 644 700
rect 806 704 812 705
rect 806 700 807 704
rect 811 700 812 704
rect 806 699 812 700
rect 974 704 980 705
rect 974 700 975 704
rect 979 700 980 704
rect 974 699 980 700
rect 1134 704 1140 705
rect 1134 700 1135 704
rect 1139 700 1140 704
rect 1134 699 1140 700
rect 1294 704 1300 705
rect 1294 700 1295 704
rect 1299 700 1300 704
rect 1294 699 1300 700
rect 1454 704 1460 705
rect 1454 700 1455 704
rect 1459 700 1460 704
rect 1454 699 1460 700
rect 1606 704 1612 705
rect 1606 700 1607 704
rect 1611 700 1612 704
rect 1606 699 1612 700
rect 1766 704 1772 705
rect 1766 700 1767 704
rect 1771 700 1772 704
rect 1766 699 1772 700
rect 1902 704 1908 705
rect 1902 700 1903 704
rect 1907 700 1908 704
rect 2008 702 2010 729
rect 2048 710 2050 737
rect 2072 713 2074 737
rect 2184 713 2186 737
rect 2336 713 2338 737
rect 2488 713 2490 737
rect 2640 713 2642 737
rect 2808 713 2810 737
rect 2984 713 2986 737
rect 3168 713 3170 737
rect 3368 713 3370 737
rect 3576 713 3578 737
rect 3784 713 3786 737
rect 2070 712 2076 713
rect 2046 709 2052 710
rect 2046 705 2047 709
rect 2051 705 2052 709
rect 2070 708 2071 712
rect 2075 708 2076 712
rect 2070 707 2076 708
rect 2182 712 2188 713
rect 2182 708 2183 712
rect 2187 708 2188 712
rect 2182 707 2188 708
rect 2334 712 2340 713
rect 2334 708 2335 712
rect 2339 708 2340 712
rect 2334 707 2340 708
rect 2486 712 2492 713
rect 2486 708 2487 712
rect 2491 708 2492 712
rect 2486 707 2492 708
rect 2638 712 2644 713
rect 2638 708 2639 712
rect 2643 708 2644 712
rect 2638 707 2644 708
rect 2806 712 2812 713
rect 2806 708 2807 712
rect 2811 708 2812 712
rect 2806 707 2812 708
rect 2982 712 2988 713
rect 2982 708 2983 712
rect 2987 708 2988 712
rect 2982 707 2988 708
rect 3166 712 3172 713
rect 3166 708 3167 712
rect 3171 708 3172 712
rect 3166 707 3172 708
rect 3366 712 3372 713
rect 3366 708 3367 712
rect 3371 708 3372 712
rect 3366 707 3372 708
rect 3574 712 3580 713
rect 3574 708 3575 712
rect 3579 708 3580 712
rect 3574 707 3580 708
rect 3782 712 3788 713
rect 3782 708 3783 712
rect 3787 708 3788 712
rect 3944 710 3946 737
rect 3782 707 3788 708
rect 3942 709 3948 710
rect 2046 704 2052 705
rect 3942 705 3943 709
rect 3947 705 3948 709
rect 3942 704 3948 705
rect 1902 699 1908 700
rect 2006 701 2012 702
rect 110 696 116 697
rect 2006 697 2007 701
rect 2011 697 2012 701
rect 2006 696 2012 697
rect 2070 693 2076 694
rect 2046 692 2052 693
rect 2046 688 2047 692
rect 2051 688 2052 692
rect 2070 689 2071 693
rect 2075 689 2076 693
rect 2070 688 2076 689
rect 2182 693 2188 694
rect 2182 689 2183 693
rect 2187 689 2188 693
rect 2182 688 2188 689
rect 2334 693 2340 694
rect 2334 689 2335 693
rect 2339 689 2340 693
rect 2334 688 2340 689
rect 2486 693 2492 694
rect 2486 689 2487 693
rect 2491 689 2492 693
rect 2486 688 2492 689
rect 2638 693 2644 694
rect 2638 689 2639 693
rect 2643 689 2644 693
rect 2638 688 2644 689
rect 2806 693 2812 694
rect 2806 689 2807 693
rect 2811 689 2812 693
rect 2806 688 2812 689
rect 2982 693 2988 694
rect 2982 689 2983 693
rect 2987 689 2988 693
rect 2982 688 2988 689
rect 3166 693 3172 694
rect 3166 689 3167 693
rect 3171 689 3172 693
rect 3166 688 3172 689
rect 3366 693 3372 694
rect 3366 689 3367 693
rect 3371 689 3372 693
rect 3366 688 3372 689
rect 3574 693 3580 694
rect 3574 689 3575 693
rect 3579 689 3580 693
rect 3574 688 3580 689
rect 3782 693 3788 694
rect 3782 689 3783 693
rect 3787 689 3788 693
rect 3782 688 3788 689
rect 3942 692 3948 693
rect 3942 688 3943 692
rect 3947 688 3948 692
rect 2046 687 2052 688
rect 310 685 316 686
rect 110 684 116 685
rect 110 680 111 684
rect 115 680 116 684
rect 310 681 311 685
rect 315 681 316 685
rect 310 680 316 681
rect 470 685 476 686
rect 470 681 471 685
rect 475 681 476 685
rect 470 680 476 681
rect 638 685 644 686
rect 638 681 639 685
rect 643 681 644 685
rect 638 680 644 681
rect 806 685 812 686
rect 806 681 807 685
rect 811 681 812 685
rect 806 680 812 681
rect 974 685 980 686
rect 974 681 975 685
rect 979 681 980 685
rect 974 680 980 681
rect 1134 685 1140 686
rect 1134 681 1135 685
rect 1139 681 1140 685
rect 1134 680 1140 681
rect 1294 685 1300 686
rect 1294 681 1295 685
rect 1299 681 1300 685
rect 1294 680 1300 681
rect 1454 685 1460 686
rect 1454 681 1455 685
rect 1459 681 1460 685
rect 1454 680 1460 681
rect 1606 685 1612 686
rect 1606 681 1607 685
rect 1611 681 1612 685
rect 1606 680 1612 681
rect 1766 685 1772 686
rect 1766 681 1767 685
rect 1771 681 1772 685
rect 1766 680 1772 681
rect 1902 685 1908 686
rect 1902 681 1903 685
rect 1907 681 1908 685
rect 1902 680 1908 681
rect 2006 684 2012 685
rect 2006 680 2007 684
rect 2011 680 2012 684
rect 110 679 116 680
rect 112 659 114 679
rect 312 659 314 680
rect 472 659 474 680
rect 640 659 642 680
rect 808 659 810 680
rect 976 659 978 680
rect 1136 659 1138 680
rect 1296 659 1298 680
rect 1456 659 1458 680
rect 1608 659 1610 680
rect 1768 659 1770 680
rect 1904 659 1906 680
rect 2006 679 2012 680
rect 2008 659 2010 679
rect 111 658 115 659
rect 111 653 115 654
rect 295 658 299 659
rect 295 653 299 654
rect 311 658 315 659
rect 311 653 315 654
rect 447 658 451 659
rect 447 653 451 654
rect 471 658 475 659
rect 471 653 475 654
rect 615 658 619 659
rect 615 653 619 654
rect 639 658 643 659
rect 639 653 643 654
rect 783 658 787 659
rect 783 653 787 654
rect 807 658 811 659
rect 807 653 811 654
rect 951 658 955 659
rect 951 653 955 654
rect 975 658 979 659
rect 975 653 979 654
rect 1111 658 1115 659
rect 1111 653 1115 654
rect 1135 658 1139 659
rect 1135 653 1139 654
rect 1263 658 1267 659
rect 1263 653 1267 654
rect 1295 658 1299 659
rect 1295 653 1299 654
rect 1399 658 1403 659
rect 1399 653 1403 654
rect 1455 658 1459 659
rect 1455 653 1459 654
rect 1535 658 1539 659
rect 1535 653 1539 654
rect 1607 658 1611 659
rect 1607 653 1611 654
rect 1663 658 1667 659
rect 1663 653 1667 654
rect 1767 658 1771 659
rect 1767 653 1771 654
rect 1791 658 1795 659
rect 1791 653 1795 654
rect 1903 658 1907 659
rect 1903 653 1907 654
rect 2007 658 2011 659
rect 2048 655 2050 687
rect 2072 655 2074 688
rect 2184 655 2186 688
rect 2336 655 2338 688
rect 2488 655 2490 688
rect 2640 655 2642 688
rect 2808 655 2810 688
rect 2984 655 2986 688
rect 3168 655 3170 688
rect 3368 655 3370 688
rect 3576 655 3578 688
rect 3784 655 3786 688
rect 3942 687 3948 688
rect 3944 655 3946 687
rect 2007 653 2011 654
rect 2047 654 2051 655
rect 112 633 114 653
rect 110 632 116 633
rect 296 632 298 653
rect 448 632 450 653
rect 616 632 618 653
rect 784 632 786 653
rect 952 632 954 653
rect 1112 632 1114 653
rect 1264 632 1266 653
rect 1400 632 1402 653
rect 1536 632 1538 653
rect 1664 632 1666 653
rect 1792 632 1794 653
rect 1904 632 1906 653
rect 2008 633 2010 653
rect 2047 649 2051 650
rect 2071 654 2075 655
rect 2071 649 2075 650
rect 2183 654 2187 655
rect 2183 649 2187 650
rect 2239 654 2243 655
rect 2239 649 2243 650
rect 2335 654 2339 655
rect 2335 649 2339 650
rect 2423 654 2427 655
rect 2423 649 2427 650
rect 2487 654 2491 655
rect 2487 649 2491 650
rect 2623 654 2627 655
rect 2623 649 2627 650
rect 2639 654 2643 655
rect 2639 649 2643 650
rect 2807 654 2811 655
rect 2807 649 2811 650
rect 2839 654 2843 655
rect 2839 649 2843 650
rect 2983 654 2987 655
rect 2983 649 2987 650
rect 3071 654 3075 655
rect 3071 649 3075 650
rect 3167 654 3171 655
rect 3167 649 3171 650
rect 3319 654 3323 655
rect 3319 649 3323 650
rect 3367 654 3371 655
rect 3367 649 3371 650
rect 3575 654 3579 655
rect 3575 649 3579 650
rect 3783 654 3787 655
rect 3783 649 3787 650
rect 3839 654 3843 655
rect 3839 649 3843 650
rect 3943 654 3947 655
rect 3943 649 3947 650
rect 2006 632 2012 633
rect 110 628 111 632
rect 115 628 116 632
rect 110 627 116 628
rect 294 631 300 632
rect 294 627 295 631
rect 299 627 300 631
rect 294 626 300 627
rect 446 631 452 632
rect 446 627 447 631
rect 451 627 452 631
rect 446 626 452 627
rect 614 631 620 632
rect 614 627 615 631
rect 619 627 620 631
rect 614 626 620 627
rect 782 631 788 632
rect 782 627 783 631
rect 787 627 788 631
rect 782 626 788 627
rect 950 631 956 632
rect 950 627 951 631
rect 955 627 956 631
rect 950 626 956 627
rect 1110 631 1116 632
rect 1110 627 1111 631
rect 1115 627 1116 631
rect 1110 626 1116 627
rect 1262 631 1268 632
rect 1262 627 1263 631
rect 1267 627 1268 631
rect 1262 626 1268 627
rect 1398 631 1404 632
rect 1398 627 1399 631
rect 1403 627 1404 631
rect 1398 626 1404 627
rect 1534 631 1540 632
rect 1534 627 1535 631
rect 1539 627 1540 631
rect 1534 626 1540 627
rect 1662 631 1668 632
rect 1662 627 1663 631
rect 1667 627 1668 631
rect 1662 626 1668 627
rect 1790 631 1796 632
rect 1790 627 1791 631
rect 1795 627 1796 631
rect 1790 626 1796 627
rect 1902 631 1908 632
rect 1902 627 1903 631
rect 1907 627 1908 631
rect 2006 628 2007 632
rect 2011 628 2012 632
rect 2048 629 2050 649
rect 2006 627 2012 628
rect 2046 628 2052 629
rect 2072 628 2074 649
rect 2240 628 2242 649
rect 2424 628 2426 649
rect 2624 628 2626 649
rect 2840 628 2842 649
rect 3072 628 3074 649
rect 3320 628 3322 649
rect 3576 628 3578 649
rect 3840 628 3842 649
rect 3944 629 3946 649
rect 3942 628 3948 629
rect 1902 626 1908 627
rect 2046 624 2047 628
rect 2051 624 2052 628
rect 2046 623 2052 624
rect 2070 627 2076 628
rect 2070 623 2071 627
rect 2075 623 2076 627
rect 2070 622 2076 623
rect 2238 627 2244 628
rect 2238 623 2239 627
rect 2243 623 2244 627
rect 2238 622 2244 623
rect 2422 627 2428 628
rect 2422 623 2423 627
rect 2427 623 2428 627
rect 2422 622 2428 623
rect 2622 627 2628 628
rect 2622 623 2623 627
rect 2627 623 2628 627
rect 2622 622 2628 623
rect 2838 627 2844 628
rect 2838 623 2839 627
rect 2843 623 2844 627
rect 2838 622 2844 623
rect 3070 627 3076 628
rect 3070 623 3071 627
rect 3075 623 3076 627
rect 3070 622 3076 623
rect 3318 627 3324 628
rect 3318 623 3319 627
rect 3323 623 3324 627
rect 3318 622 3324 623
rect 3574 627 3580 628
rect 3574 623 3575 627
rect 3579 623 3580 627
rect 3574 622 3580 623
rect 3838 627 3844 628
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3942 624 3943 628
rect 3947 624 3948 628
rect 3942 623 3948 624
rect 3838 622 3844 623
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 2006 615 2012 616
rect 110 610 116 611
rect 294 612 300 613
rect 112 579 114 610
rect 294 608 295 612
rect 299 608 300 612
rect 294 607 300 608
rect 446 612 452 613
rect 446 608 447 612
rect 451 608 452 612
rect 446 607 452 608
rect 614 612 620 613
rect 614 608 615 612
rect 619 608 620 612
rect 614 607 620 608
rect 782 612 788 613
rect 782 608 783 612
rect 787 608 788 612
rect 782 607 788 608
rect 950 612 956 613
rect 950 608 951 612
rect 955 608 956 612
rect 950 607 956 608
rect 1110 612 1116 613
rect 1110 608 1111 612
rect 1115 608 1116 612
rect 1110 607 1116 608
rect 1262 612 1268 613
rect 1262 608 1263 612
rect 1267 608 1268 612
rect 1262 607 1268 608
rect 1398 612 1404 613
rect 1398 608 1399 612
rect 1403 608 1404 612
rect 1398 607 1404 608
rect 1534 612 1540 613
rect 1534 608 1535 612
rect 1539 608 1540 612
rect 1534 607 1540 608
rect 1662 612 1668 613
rect 1662 608 1663 612
rect 1667 608 1668 612
rect 1662 607 1668 608
rect 1790 612 1796 613
rect 1790 608 1791 612
rect 1795 608 1796 612
rect 1790 607 1796 608
rect 1902 612 1908 613
rect 1902 608 1903 612
rect 1907 608 1908 612
rect 2006 611 2007 615
rect 2011 611 2012 615
rect 2006 610 2012 611
rect 2046 611 2052 612
rect 1902 607 1908 608
rect 296 579 298 607
rect 448 579 450 607
rect 616 579 618 607
rect 784 579 786 607
rect 952 579 954 607
rect 1112 579 1114 607
rect 1264 579 1266 607
rect 1400 579 1402 607
rect 1536 579 1538 607
rect 1664 579 1666 607
rect 1792 579 1794 607
rect 1904 579 1906 607
rect 2008 579 2010 610
rect 2046 607 2047 611
rect 2051 607 2052 611
rect 3942 611 3948 612
rect 2046 606 2052 607
rect 2070 608 2076 609
rect 2048 579 2050 606
rect 2070 604 2071 608
rect 2075 604 2076 608
rect 2070 603 2076 604
rect 2238 608 2244 609
rect 2238 604 2239 608
rect 2243 604 2244 608
rect 2238 603 2244 604
rect 2422 608 2428 609
rect 2422 604 2423 608
rect 2427 604 2428 608
rect 2422 603 2428 604
rect 2622 608 2628 609
rect 2622 604 2623 608
rect 2627 604 2628 608
rect 2622 603 2628 604
rect 2838 608 2844 609
rect 2838 604 2839 608
rect 2843 604 2844 608
rect 2838 603 2844 604
rect 3070 608 3076 609
rect 3070 604 3071 608
rect 3075 604 3076 608
rect 3070 603 3076 604
rect 3318 608 3324 609
rect 3318 604 3319 608
rect 3323 604 3324 608
rect 3318 603 3324 604
rect 3574 608 3580 609
rect 3574 604 3575 608
rect 3579 604 3580 608
rect 3574 603 3580 604
rect 3838 608 3844 609
rect 3838 604 3839 608
rect 3843 604 3844 608
rect 3942 607 3943 611
rect 3947 607 3948 611
rect 3942 606 3948 607
rect 3838 603 3844 604
rect 2072 579 2074 603
rect 2240 579 2242 603
rect 2424 579 2426 603
rect 2624 579 2626 603
rect 2840 579 2842 603
rect 3072 579 3074 603
rect 3320 579 3322 603
rect 3576 579 3578 603
rect 3840 579 3842 603
rect 3944 579 3946 606
rect 111 578 115 579
rect 111 573 115 574
rect 239 578 243 579
rect 239 573 243 574
rect 295 578 299 579
rect 295 573 299 574
rect 415 578 419 579
rect 415 573 419 574
rect 447 578 451 579
rect 447 573 451 574
rect 607 578 611 579
rect 607 573 611 574
rect 615 578 619 579
rect 615 573 619 574
rect 783 578 787 579
rect 783 573 787 574
rect 799 578 803 579
rect 799 573 803 574
rect 951 578 955 579
rect 951 573 955 574
rect 991 578 995 579
rect 991 573 995 574
rect 1111 578 1115 579
rect 1111 573 1115 574
rect 1175 578 1179 579
rect 1175 573 1179 574
rect 1263 578 1267 579
rect 1263 573 1267 574
rect 1351 578 1355 579
rect 1351 573 1355 574
rect 1399 578 1403 579
rect 1399 573 1403 574
rect 1519 578 1523 579
rect 1519 573 1523 574
rect 1535 578 1539 579
rect 1535 573 1539 574
rect 1663 578 1667 579
rect 1663 573 1667 574
rect 1687 578 1691 579
rect 1687 573 1691 574
rect 1791 578 1795 579
rect 1791 573 1795 574
rect 1863 578 1867 579
rect 1863 573 1867 574
rect 1903 578 1907 579
rect 1903 573 1907 574
rect 2007 578 2011 579
rect 2007 573 2011 574
rect 2047 578 2051 579
rect 2047 573 2051 574
rect 2071 578 2075 579
rect 2071 573 2075 574
rect 2191 578 2195 579
rect 2191 573 2195 574
rect 2239 578 2243 579
rect 2239 573 2243 574
rect 2287 578 2291 579
rect 2287 573 2291 574
rect 2383 578 2387 579
rect 2383 573 2387 574
rect 2423 578 2427 579
rect 2423 573 2427 574
rect 2479 578 2483 579
rect 2479 573 2483 574
rect 2583 578 2587 579
rect 2583 573 2587 574
rect 2623 578 2627 579
rect 2623 573 2627 574
rect 2711 578 2715 579
rect 2711 573 2715 574
rect 2839 578 2843 579
rect 2839 573 2843 574
rect 2871 578 2875 579
rect 2871 573 2875 574
rect 3071 578 3075 579
rect 3071 573 3075 574
rect 3303 578 3307 579
rect 3303 573 3307 574
rect 3319 578 3323 579
rect 3319 573 3323 574
rect 3551 578 3555 579
rect 3551 573 3555 574
rect 3575 578 3579 579
rect 3575 573 3579 574
rect 3807 578 3811 579
rect 3807 573 3811 574
rect 3839 578 3843 579
rect 3839 573 3843 574
rect 3943 578 3947 579
rect 3943 573 3947 574
rect 112 546 114 573
rect 240 549 242 573
rect 416 549 418 573
rect 608 549 610 573
rect 800 549 802 573
rect 992 549 994 573
rect 1176 549 1178 573
rect 1352 549 1354 573
rect 1520 549 1522 573
rect 1688 549 1690 573
rect 1864 549 1866 573
rect 238 548 244 549
rect 110 545 116 546
rect 110 541 111 545
rect 115 541 116 545
rect 238 544 239 548
rect 243 544 244 548
rect 238 543 244 544
rect 414 548 420 549
rect 414 544 415 548
rect 419 544 420 548
rect 414 543 420 544
rect 606 548 612 549
rect 606 544 607 548
rect 611 544 612 548
rect 606 543 612 544
rect 798 548 804 549
rect 798 544 799 548
rect 803 544 804 548
rect 798 543 804 544
rect 990 548 996 549
rect 990 544 991 548
rect 995 544 996 548
rect 990 543 996 544
rect 1174 548 1180 549
rect 1174 544 1175 548
rect 1179 544 1180 548
rect 1174 543 1180 544
rect 1350 548 1356 549
rect 1350 544 1351 548
rect 1355 544 1356 548
rect 1350 543 1356 544
rect 1518 548 1524 549
rect 1518 544 1519 548
rect 1523 544 1524 548
rect 1518 543 1524 544
rect 1686 548 1692 549
rect 1686 544 1687 548
rect 1691 544 1692 548
rect 1686 543 1692 544
rect 1862 548 1868 549
rect 1862 544 1863 548
rect 1867 544 1868 548
rect 2008 546 2010 573
rect 2048 546 2050 573
rect 2192 549 2194 573
rect 2288 549 2290 573
rect 2384 549 2386 573
rect 2480 549 2482 573
rect 2584 549 2586 573
rect 2712 549 2714 573
rect 2872 549 2874 573
rect 3072 549 3074 573
rect 3304 549 3306 573
rect 3552 549 3554 573
rect 3808 549 3810 573
rect 2190 548 2196 549
rect 1862 543 1868 544
rect 2006 545 2012 546
rect 110 540 116 541
rect 2006 541 2007 545
rect 2011 541 2012 545
rect 2006 540 2012 541
rect 2046 545 2052 546
rect 2046 541 2047 545
rect 2051 541 2052 545
rect 2190 544 2191 548
rect 2195 544 2196 548
rect 2190 543 2196 544
rect 2286 548 2292 549
rect 2286 544 2287 548
rect 2291 544 2292 548
rect 2286 543 2292 544
rect 2382 548 2388 549
rect 2382 544 2383 548
rect 2387 544 2388 548
rect 2382 543 2388 544
rect 2478 548 2484 549
rect 2478 544 2479 548
rect 2483 544 2484 548
rect 2478 543 2484 544
rect 2582 548 2588 549
rect 2582 544 2583 548
rect 2587 544 2588 548
rect 2582 543 2588 544
rect 2710 548 2716 549
rect 2710 544 2711 548
rect 2715 544 2716 548
rect 2710 543 2716 544
rect 2870 548 2876 549
rect 2870 544 2871 548
rect 2875 544 2876 548
rect 2870 543 2876 544
rect 3070 548 3076 549
rect 3070 544 3071 548
rect 3075 544 3076 548
rect 3070 543 3076 544
rect 3302 548 3308 549
rect 3302 544 3303 548
rect 3307 544 3308 548
rect 3302 543 3308 544
rect 3550 548 3556 549
rect 3550 544 3551 548
rect 3555 544 3556 548
rect 3550 543 3556 544
rect 3806 548 3812 549
rect 3806 544 3807 548
rect 3811 544 3812 548
rect 3944 546 3946 573
rect 3806 543 3812 544
rect 3942 545 3948 546
rect 2046 540 2052 541
rect 3942 541 3943 545
rect 3947 541 3948 545
rect 3942 540 3948 541
rect 238 529 244 530
rect 110 528 116 529
rect 110 524 111 528
rect 115 524 116 528
rect 238 525 239 529
rect 243 525 244 529
rect 238 524 244 525
rect 414 529 420 530
rect 414 525 415 529
rect 419 525 420 529
rect 414 524 420 525
rect 606 529 612 530
rect 606 525 607 529
rect 611 525 612 529
rect 606 524 612 525
rect 798 529 804 530
rect 798 525 799 529
rect 803 525 804 529
rect 798 524 804 525
rect 990 529 996 530
rect 990 525 991 529
rect 995 525 996 529
rect 990 524 996 525
rect 1174 529 1180 530
rect 1174 525 1175 529
rect 1179 525 1180 529
rect 1174 524 1180 525
rect 1350 529 1356 530
rect 1350 525 1351 529
rect 1355 525 1356 529
rect 1350 524 1356 525
rect 1518 529 1524 530
rect 1518 525 1519 529
rect 1523 525 1524 529
rect 1518 524 1524 525
rect 1686 529 1692 530
rect 1686 525 1687 529
rect 1691 525 1692 529
rect 1686 524 1692 525
rect 1862 529 1868 530
rect 2190 529 2196 530
rect 1862 525 1863 529
rect 1867 525 1868 529
rect 1862 524 1868 525
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 110 523 116 524
rect 112 503 114 523
rect 240 503 242 524
rect 416 503 418 524
rect 608 503 610 524
rect 800 503 802 524
rect 992 503 994 524
rect 1176 503 1178 524
rect 1352 503 1354 524
rect 1520 503 1522 524
rect 1688 503 1690 524
rect 1864 503 1866 524
rect 2006 523 2012 524
rect 2046 528 2052 529
rect 2046 524 2047 528
rect 2051 524 2052 528
rect 2190 525 2191 529
rect 2195 525 2196 529
rect 2190 524 2196 525
rect 2286 529 2292 530
rect 2286 525 2287 529
rect 2291 525 2292 529
rect 2286 524 2292 525
rect 2382 529 2388 530
rect 2382 525 2383 529
rect 2387 525 2388 529
rect 2382 524 2388 525
rect 2478 529 2484 530
rect 2478 525 2479 529
rect 2483 525 2484 529
rect 2478 524 2484 525
rect 2582 529 2588 530
rect 2582 525 2583 529
rect 2587 525 2588 529
rect 2582 524 2588 525
rect 2710 529 2716 530
rect 2710 525 2711 529
rect 2715 525 2716 529
rect 2710 524 2716 525
rect 2870 529 2876 530
rect 2870 525 2871 529
rect 2875 525 2876 529
rect 2870 524 2876 525
rect 3070 529 3076 530
rect 3070 525 3071 529
rect 3075 525 3076 529
rect 3070 524 3076 525
rect 3302 529 3308 530
rect 3302 525 3303 529
rect 3307 525 3308 529
rect 3302 524 3308 525
rect 3550 529 3556 530
rect 3550 525 3551 529
rect 3555 525 3556 529
rect 3550 524 3556 525
rect 3806 529 3812 530
rect 3806 525 3807 529
rect 3811 525 3812 529
rect 3806 524 3812 525
rect 3942 528 3948 529
rect 3942 524 3943 528
rect 3947 524 3948 528
rect 2046 523 2052 524
rect 2008 503 2010 523
rect 2048 503 2050 523
rect 2192 503 2194 524
rect 2288 503 2290 524
rect 2384 503 2386 524
rect 2480 503 2482 524
rect 2584 503 2586 524
rect 2712 503 2714 524
rect 2872 503 2874 524
rect 3072 503 3074 524
rect 3304 503 3306 524
rect 3552 503 3554 524
rect 3808 503 3810 524
rect 3942 523 3948 524
rect 3944 503 3946 523
rect 111 502 115 503
rect 111 497 115 498
rect 135 502 139 503
rect 135 497 139 498
rect 239 502 243 503
rect 239 497 243 498
rect 287 502 291 503
rect 287 497 291 498
rect 415 502 419 503
rect 415 497 419 498
rect 463 502 467 503
rect 463 497 467 498
rect 607 502 611 503
rect 607 497 611 498
rect 639 502 643 503
rect 639 497 643 498
rect 799 502 803 503
rect 799 497 803 498
rect 807 502 811 503
rect 807 497 811 498
rect 967 502 971 503
rect 967 497 971 498
rect 991 502 995 503
rect 991 497 995 498
rect 1119 502 1123 503
rect 1119 497 1123 498
rect 1175 502 1179 503
rect 1175 497 1179 498
rect 1271 502 1275 503
rect 1271 497 1275 498
rect 1351 502 1355 503
rect 1351 497 1355 498
rect 1415 502 1419 503
rect 1415 497 1419 498
rect 1519 502 1523 503
rect 1519 497 1523 498
rect 1567 502 1571 503
rect 1567 497 1571 498
rect 1687 502 1691 503
rect 1687 497 1691 498
rect 1863 502 1867 503
rect 1863 497 1867 498
rect 2007 502 2011 503
rect 2007 497 2011 498
rect 2047 502 2051 503
rect 2047 497 2051 498
rect 2191 502 2195 503
rect 2191 497 2195 498
rect 2287 502 2291 503
rect 2287 497 2291 498
rect 2383 502 2387 503
rect 2383 497 2387 498
rect 2431 502 2435 503
rect 2431 497 2435 498
rect 2479 502 2483 503
rect 2479 497 2483 498
rect 2527 502 2531 503
rect 2527 497 2531 498
rect 2583 502 2587 503
rect 2583 497 2587 498
rect 2623 502 2627 503
rect 2623 497 2627 498
rect 2711 502 2715 503
rect 2711 497 2715 498
rect 2727 502 2731 503
rect 2727 497 2731 498
rect 2847 502 2851 503
rect 2847 497 2851 498
rect 2871 502 2875 503
rect 2871 497 2875 498
rect 2999 502 3003 503
rect 2999 497 3003 498
rect 3071 502 3075 503
rect 3071 497 3075 498
rect 3175 502 3179 503
rect 3175 497 3179 498
rect 3303 502 3307 503
rect 3303 497 3307 498
rect 3375 502 3379 503
rect 3375 497 3379 498
rect 3551 502 3555 503
rect 3551 497 3555 498
rect 3591 502 3595 503
rect 3591 497 3595 498
rect 3807 502 3811 503
rect 3807 497 3811 498
rect 3943 502 3947 503
rect 3943 497 3947 498
rect 112 477 114 497
rect 110 476 116 477
rect 136 476 138 497
rect 288 476 290 497
rect 464 476 466 497
rect 640 476 642 497
rect 808 476 810 497
rect 968 476 970 497
rect 1120 476 1122 497
rect 1272 476 1274 497
rect 1416 476 1418 497
rect 1568 476 1570 497
rect 2008 477 2010 497
rect 2048 477 2050 497
rect 2006 476 2012 477
rect 110 472 111 476
rect 115 472 116 476
rect 110 471 116 472
rect 134 475 140 476
rect 134 471 135 475
rect 139 471 140 475
rect 134 470 140 471
rect 286 475 292 476
rect 286 471 287 475
rect 291 471 292 475
rect 286 470 292 471
rect 462 475 468 476
rect 462 471 463 475
rect 467 471 468 475
rect 462 470 468 471
rect 638 475 644 476
rect 638 471 639 475
rect 643 471 644 475
rect 638 470 644 471
rect 806 475 812 476
rect 806 471 807 475
rect 811 471 812 475
rect 806 470 812 471
rect 966 475 972 476
rect 966 471 967 475
rect 971 471 972 475
rect 966 470 972 471
rect 1118 475 1124 476
rect 1118 471 1119 475
rect 1123 471 1124 475
rect 1118 470 1124 471
rect 1270 475 1276 476
rect 1270 471 1271 475
rect 1275 471 1276 475
rect 1270 470 1276 471
rect 1414 475 1420 476
rect 1414 471 1415 475
rect 1419 471 1420 475
rect 1414 470 1420 471
rect 1566 475 1572 476
rect 1566 471 1567 475
rect 1571 471 1572 475
rect 2006 472 2007 476
rect 2011 472 2012 476
rect 2006 471 2012 472
rect 2046 476 2052 477
rect 2432 476 2434 497
rect 2528 476 2530 497
rect 2624 476 2626 497
rect 2728 476 2730 497
rect 2848 476 2850 497
rect 3000 476 3002 497
rect 3176 476 3178 497
rect 3376 476 3378 497
rect 3592 476 3594 497
rect 3808 476 3810 497
rect 3944 477 3946 497
rect 3942 476 3948 477
rect 2046 472 2047 476
rect 2051 472 2052 476
rect 2046 471 2052 472
rect 2430 475 2436 476
rect 2430 471 2431 475
rect 2435 471 2436 475
rect 1566 470 1572 471
rect 2430 470 2436 471
rect 2526 475 2532 476
rect 2526 471 2527 475
rect 2531 471 2532 475
rect 2526 470 2532 471
rect 2622 475 2628 476
rect 2622 471 2623 475
rect 2627 471 2628 475
rect 2622 470 2628 471
rect 2726 475 2732 476
rect 2726 471 2727 475
rect 2731 471 2732 475
rect 2726 470 2732 471
rect 2846 475 2852 476
rect 2846 471 2847 475
rect 2851 471 2852 475
rect 2846 470 2852 471
rect 2998 475 3004 476
rect 2998 471 2999 475
rect 3003 471 3004 475
rect 2998 470 3004 471
rect 3174 475 3180 476
rect 3174 471 3175 475
rect 3179 471 3180 475
rect 3174 470 3180 471
rect 3374 475 3380 476
rect 3374 471 3375 475
rect 3379 471 3380 475
rect 3374 470 3380 471
rect 3590 475 3596 476
rect 3590 471 3591 475
rect 3595 471 3596 475
rect 3590 470 3596 471
rect 3806 475 3812 476
rect 3806 471 3807 475
rect 3811 471 3812 475
rect 3942 472 3943 476
rect 3947 472 3948 476
rect 3942 471 3948 472
rect 3806 470 3812 471
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 2006 459 2012 460
rect 110 454 116 455
rect 134 456 140 457
rect 112 423 114 454
rect 134 452 135 456
rect 139 452 140 456
rect 134 451 140 452
rect 286 456 292 457
rect 286 452 287 456
rect 291 452 292 456
rect 286 451 292 452
rect 462 456 468 457
rect 462 452 463 456
rect 467 452 468 456
rect 462 451 468 452
rect 638 456 644 457
rect 638 452 639 456
rect 643 452 644 456
rect 638 451 644 452
rect 806 456 812 457
rect 806 452 807 456
rect 811 452 812 456
rect 806 451 812 452
rect 966 456 972 457
rect 966 452 967 456
rect 971 452 972 456
rect 966 451 972 452
rect 1118 456 1124 457
rect 1118 452 1119 456
rect 1123 452 1124 456
rect 1118 451 1124 452
rect 1270 456 1276 457
rect 1270 452 1271 456
rect 1275 452 1276 456
rect 1270 451 1276 452
rect 1414 456 1420 457
rect 1414 452 1415 456
rect 1419 452 1420 456
rect 1414 451 1420 452
rect 1566 456 1572 457
rect 1566 452 1567 456
rect 1571 452 1572 456
rect 2006 455 2007 459
rect 2011 455 2012 459
rect 2006 454 2012 455
rect 2046 459 2052 460
rect 2046 455 2047 459
rect 2051 455 2052 459
rect 3942 459 3948 460
rect 2046 454 2052 455
rect 2430 456 2436 457
rect 1566 451 1572 452
rect 136 423 138 451
rect 288 423 290 451
rect 464 423 466 451
rect 640 423 642 451
rect 808 423 810 451
rect 968 423 970 451
rect 1120 423 1122 451
rect 1272 423 1274 451
rect 1416 423 1418 451
rect 1568 423 1570 451
rect 2008 423 2010 454
rect 2048 427 2050 454
rect 2430 452 2431 456
rect 2435 452 2436 456
rect 2430 451 2436 452
rect 2526 456 2532 457
rect 2526 452 2527 456
rect 2531 452 2532 456
rect 2526 451 2532 452
rect 2622 456 2628 457
rect 2622 452 2623 456
rect 2627 452 2628 456
rect 2622 451 2628 452
rect 2726 456 2732 457
rect 2726 452 2727 456
rect 2731 452 2732 456
rect 2726 451 2732 452
rect 2846 456 2852 457
rect 2846 452 2847 456
rect 2851 452 2852 456
rect 2846 451 2852 452
rect 2998 456 3004 457
rect 2998 452 2999 456
rect 3003 452 3004 456
rect 2998 451 3004 452
rect 3174 456 3180 457
rect 3174 452 3175 456
rect 3179 452 3180 456
rect 3174 451 3180 452
rect 3374 456 3380 457
rect 3374 452 3375 456
rect 3379 452 3380 456
rect 3374 451 3380 452
rect 3590 456 3596 457
rect 3590 452 3591 456
rect 3595 452 3596 456
rect 3590 451 3596 452
rect 3806 456 3812 457
rect 3806 452 3807 456
rect 3811 452 3812 456
rect 3942 455 3943 459
rect 3947 455 3948 459
rect 3942 454 3948 455
rect 3806 451 3812 452
rect 2432 427 2434 451
rect 2528 427 2530 451
rect 2624 427 2626 451
rect 2728 427 2730 451
rect 2848 427 2850 451
rect 3000 427 3002 451
rect 3176 427 3178 451
rect 3376 427 3378 451
rect 3592 427 3594 451
rect 3808 427 3810 451
rect 3944 427 3946 454
rect 2047 426 2051 427
rect 111 422 115 423
rect 111 417 115 418
rect 135 422 139 423
rect 135 417 139 418
rect 279 422 283 423
rect 279 417 283 418
rect 287 422 291 423
rect 287 417 291 418
rect 439 422 443 423
rect 439 417 443 418
rect 463 422 467 423
rect 463 417 467 418
rect 583 422 587 423
rect 583 417 587 418
rect 639 422 643 423
rect 639 417 643 418
rect 719 422 723 423
rect 719 417 723 418
rect 807 422 811 423
rect 807 417 811 418
rect 847 422 851 423
rect 847 417 851 418
rect 967 422 971 423
rect 967 417 971 418
rect 1087 422 1091 423
rect 1087 417 1091 418
rect 1119 422 1123 423
rect 1119 417 1123 418
rect 1207 422 1211 423
rect 1207 417 1211 418
rect 1271 422 1275 423
rect 1271 417 1275 418
rect 1327 422 1331 423
rect 1327 417 1331 418
rect 1415 422 1419 423
rect 1415 417 1419 418
rect 1567 422 1571 423
rect 1567 417 1571 418
rect 2007 422 2011 423
rect 2047 421 2051 422
rect 2431 426 2435 427
rect 2431 421 2435 422
rect 2527 426 2531 427
rect 2527 421 2531 422
rect 2623 426 2627 427
rect 2623 421 2627 422
rect 2719 426 2723 427
rect 2719 421 2723 422
rect 2727 426 2731 427
rect 2727 421 2731 422
rect 2815 426 2819 427
rect 2815 421 2819 422
rect 2847 426 2851 427
rect 2847 421 2851 422
rect 2927 426 2931 427
rect 2927 421 2931 422
rect 2999 426 3003 427
rect 2999 421 3003 422
rect 3063 426 3067 427
rect 3063 421 3067 422
rect 3175 426 3179 427
rect 3175 421 3179 422
rect 3223 426 3227 427
rect 3223 421 3227 422
rect 3375 426 3379 427
rect 3375 421 3379 422
rect 3399 426 3403 427
rect 3399 421 3403 422
rect 3591 426 3595 427
rect 3591 421 3595 422
rect 3783 426 3787 427
rect 3783 421 3787 422
rect 3807 426 3811 427
rect 3807 421 3811 422
rect 3943 426 3947 427
rect 3943 421 3947 422
rect 2007 417 2011 418
rect 112 390 114 417
rect 136 393 138 417
rect 280 393 282 417
rect 440 393 442 417
rect 584 393 586 417
rect 720 393 722 417
rect 848 393 850 417
rect 968 393 970 417
rect 1088 393 1090 417
rect 1208 393 1210 417
rect 1328 393 1330 417
rect 134 392 140 393
rect 110 389 116 390
rect 110 385 111 389
rect 115 385 116 389
rect 134 388 135 392
rect 139 388 140 392
rect 134 387 140 388
rect 278 392 284 393
rect 278 388 279 392
rect 283 388 284 392
rect 278 387 284 388
rect 438 392 444 393
rect 438 388 439 392
rect 443 388 444 392
rect 438 387 444 388
rect 582 392 588 393
rect 582 388 583 392
rect 587 388 588 392
rect 582 387 588 388
rect 718 392 724 393
rect 718 388 719 392
rect 723 388 724 392
rect 718 387 724 388
rect 846 392 852 393
rect 846 388 847 392
rect 851 388 852 392
rect 846 387 852 388
rect 966 392 972 393
rect 966 388 967 392
rect 971 388 972 392
rect 966 387 972 388
rect 1086 392 1092 393
rect 1086 388 1087 392
rect 1091 388 1092 392
rect 1086 387 1092 388
rect 1206 392 1212 393
rect 1206 388 1207 392
rect 1211 388 1212 392
rect 1206 387 1212 388
rect 1326 392 1332 393
rect 1326 388 1327 392
rect 1331 388 1332 392
rect 2008 390 2010 417
rect 2048 394 2050 421
rect 2432 397 2434 421
rect 2528 397 2530 421
rect 2624 397 2626 421
rect 2720 397 2722 421
rect 2816 397 2818 421
rect 2928 397 2930 421
rect 3064 397 3066 421
rect 3224 397 3226 421
rect 3400 397 3402 421
rect 3592 397 3594 421
rect 3784 397 3786 421
rect 2430 396 2436 397
rect 2046 393 2052 394
rect 1326 387 1332 388
rect 2006 389 2012 390
rect 110 384 116 385
rect 2006 385 2007 389
rect 2011 385 2012 389
rect 2046 389 2047 393
rect 2051 389 2052 393
rect 2430 392 2431 396
rect 2435 392 2436 396
rect 2430 391 2436 392
rect 2526 396 2532 397
rect 2526 392 2527 396
rect 2531 392 2532 396
rect 2526 391 2532 392
rect 2622 396 2628 397
rect 2622 392 2623 396
rect 2627 392 2628 396
rect 2622 391 2628 392
rect 2718 396 2724 397
rect 2718 392 2719 396
rect 2723 392 2724 396
rect 2718 391 2724 392
rect 2814 396 2820 397
rect 2814 392 2815 396
rect 2819 392 2820 396
rect 2814 391 2820 392
rect 2926 396 2932 397
rect 2926 392 2927 396
rect 2931 392 2932 396
rect 2926 391 2932 392
rect 3062 396 3068 397
rect 3062 392 3063 396
rect 3067 392 3068 396
rect 3062 391 3068 392
rect 3222 396 3228 397
rect 3222 392 3223 396
rect 3227 392 3228 396
rect 3222 391 3228 392
rect 3398 396 3404 397
rect 3398 392 3399 396
rect 3403 392 3404 396
rect 3398 391 3404 392
rect 3590 396 3596 397
rect 3590 392 3591 396
rect 3595 392 3596 396
rect 3590 391 3596 392
rect 3782 396 3788 397
rect 3782 392 3783 396
rect 3787 392 3788 396
rect 3944 394 3946 421
rect 3782 391 3788 392
rect 3942 393 3948 394
rect 2046 388 2052 389
rect 3942 389 3943 393
rect 3947 389 3948 393
rect 3942 388 3948 389
rect 2006 384 2012 385
rect 2430 377 2436 378
rect 2046 376 2052 377
rect 134 373 140 374
rect 110 372 116 373
rect 110 368 111 372
rect 115 368 116 372
rect 134 369 135 373
rect 139 369 140 373
rect 134 368 140 369
rect 278 373 284 374
rect 278 369 279 373
rect 283 369 284 373
rect 278 368 284 369
rect 438 373 444 374
rect 438 369 439 373
rect 443 369 444 373
rect 438 368 444 369
rect 582 373 588 374
rect 582 369 583 373
rect 587 369 588 373
rect 582 368 588 369
rect 718 373 724 374
rect 718 369 719 373
rect 723 369 724 373
rect 718 368 724 369
rect 846 373 852 374
rect 846 369 847 373
rect 851 369 852 373
rect 846 368 852 369
rect 966 373 972 374
rect 966 369 967 373
rect 971 369 972 373
rect 966 368 972 369
rect 1086 373 1092 374
rect 1086 369 1087 373
rect 1091 369 1092 373
rect 1086 368 1092 369
rect 1206 373 1212 374
rect 1206 369 1207 373
rect 1211 369 1212 373
rect 1206 368 1212 369
rect 1326 373 1332 374
rect 1326 369 1327 373
rect 1331 369 1332 373
rect 1326 368 1332 369
rect 2006 372 2012 373
rect 2006 368 2007 372
rect 2011 368 2012 372
rect 2046 372 2047 376
rect 2051 372 2052 376
rect 2430 373 2431 377
rect 2435 373 2436 377
rect 2430 372 2436 373
rect 2526 377 2532 378
rect 2526 373 2527 377
rect 2531 373 2532 377
rect 2526 372 2532 373
rect 2622 377 2628 378
rect 2622 373 2623 377
rect 2627 373 2628 377
rect 2622 372 2628 373
rect 2718 377 2724 378
rect 2718 373 2719 377
rect 2723 373 2724 377
rect 2718 372 2724 373
rect 2814 377 2820 378
rect 2814 373 2815 377
rect 2819 373 2820 377
rect 2814 372 2820 373
rect 2926 377 2932 378
rect 2926 373 2927 377
rect 2931 373 2932 377
rect 2926 372 2932 373
rect 3062 377 3068 378
rect 3062 373 3063 377
rect 3067 373 3068 377
rect 3062 372 3068 373
rect 3222 377 3228 378
rect 3222 373 3223 377
rect 3227 373 3228 377
rect 3222 372 3228 373
rect 3398 377 3404 378
rect 3398 373 3399 377
rect 3403 373 3404 377
rect 3398 372 3404 373
rect 3590 377 3596 378
rect 3590 373 3591 377
rect 3595 373 3596 377
rect 3590 372 3596 373
rect 3782 377 3788 378
rect 3782 373 3783 377
rect 3787 373 3788 377
rect 3782 372 3788 373
rect 3942 376 3948 377
rect 3942 372 3943 376
rect 3947 372 3948 376
rect 2046 371 2052 372
rect 110 367 116 368
rect 112 347 114 367
rect 136 347 138 368
rect 280 347 282 368
rect 440 347 442 368
rect 584 347 586 368
rect 720 347 722 368
rect 848 347 850 368
rect 968 347 970 368
rect 1088 347 1090 368
rect 1208 347 1210 368
rect 1328 347 1330 368
rect 2006 367 2012 368
rect 2008 347 2010 367
rect 2048 347 2050 371
rect 2432 347 2434 372
rect 2528 347 2530 372
rect 2624 347 2626 372
rect 2720 347 2722 372
rect 2816 347 2818 372
rect 2928 347 2930 372
rect 3064 347 3066 372
rect 3224 347 3226 372
rect 3400 347 3402 372
rect 3592 347 3594 372
rect 3784 347 3786 372
rect 3942 371 3948 372
rect 3944 347 3946 371
rect 111 346 115 347
rect 111 341 115 342
rect 135 346 139 347
rect 135 341 139 342
rect 143 346 147 347
rect 143 341 147 342
rect 279 346 283 347
rect 279 341 283 342
rect 319 346 323 347
rect 319 341 323 342
rect 439 346 443 347
rect 439 341 443 342
rect 479 346 483 347
rect 479 341 483 342
rect 583 346 587 347
rect 583 341 587 342
rect 631 346 635 347
rect 631 341 635 342
rect 719 346 723 347
rect 719 341 723 342
rect 775 346 779 347
rect 775 341 779 342
rect 847 346 851 347
rect 847 341 851 342
rect 903 346 907 347
rect 903 341 907 342
rect 967 346 971 347
rect 967 341 971 342
rect 1031 346 1035 347
rect 1031 341 1035 342
rect 1087 346 1091 347
rect 1087 341 1091 342
rect 1151 346 1155 347
rect 1151 341 1155 342
rect 1207 346 1211 347
rect 1207 341 1211 342
rect 1271 346 1275 347
rect 1271 341 1275 342
rect 1327 346 1331 347
rect 1327 341 1331 342
rect 1391 346 1395 347
rect 1391 341 1395 342
rect 2007 346 2011 347
rect 2007 341 2011 342
rect 2047 346 2051 347
rect 2047 341 2051 342
rect 2191 346 2195 347
rect 2191 341 2195 342
rect 2327 346 2331 347
rect 2327 341 2331 342
rect 2431 346 2435 347
rect 2431 341 2435 342
rect 2471 346 2475 347
rect 2471 341 2475 342
rect 2527 346 2531 347
rect 2527 341 2531 342
rect 2623 346 2627 347
rect 2623 341 2627 342
rect 2719 346 2723 347
rect 2719 341 2723 342
rect 2783 346 2787 347
rect 2783 341 2787 342
rect 2815 346 2819 347
rect 2815 341 2819 342
rect 2927 346 2931 347
rect 2927 341 2931 342
rect 2951 346 2955 347
rect 2951 341 2955 342
rect 3063 346 3067 347
rect 3063 341 3067 342
rect 3119 346 3123 347
rect 3119 341 3123 342
rect 3223 346 3227 347
rect 3223 341 3227 342
rect 3295 346 3299 347
rect 3295 341 3299 342
rect 3399 346 3403 347
rect 3399 341 3403 342
rect 3471 346 3475 347
rect 3471 341 3475 342
rect 3591 346 3595 347
rect 3591 341 3595 342
rect 3655 346 3659 347
rect 3655 341 3659 342
rect 3783 346 3787 347
rect 3783 341 3787 342
rect 3839 346 3843 347
rect 3839 341 3843 342
rect 3943 346 3947 347
rect 3943 341 3947 342
rect 112 321 114 341
rect 110 320 116 321
rect 144 320 146 341
rect 320 320 322 341
rect 480 320 482 341
rect 632 320 634 341
rect 776 320 778 341
rect 904 320 906 341
rect 1032 320 1034 341
rect 1152 320 1154 341
rect 1272 320 1274 341
rect 1392 320 1394 341
rect 2008 321 2010 341
rect 2048 321 2050 341
rect 2006 320 2012 321
rect 110 316 111 320
rect 115 316 116 320
rect 110 315 116 316
rect 142 319 148 320
rect 142 315 143 319
rect 147 315 148 319
rect 142 314 148 315
rect 318 319 324 320
rect 318 315 319 319
rect 323 315 324 319
rect 318 314 324 315
rect 478 319 484 320
rect 478 315 479 319
rect 483 315 484 319
rect 478 314 484 315
rect 630 319 636 320
rect 630 315 631 319
rect 635 315 636 319
rect 630 314 636 315
rect 774 319 780 320
rect 774 315 775 319
rect 779 315 780 319
rect 774 314 780 315
rect 902 319 908 320
rect 902 315 903 319
rect 907 315 908 319
rect 902 314 908 315
rect 1030 319 1036 320
rect 1030 315 1031 319
rect 1035 315 1036 319
rect 1030 314 1036 315
rect 1150 319 1156 320
rect 1150 315 1151 319
rect 1155 315 1156 319
rect 1150 314 1156 315
rect 1270 319 1276 320
rect 1270 315 1271 319
rect 1275 315 1276 319
rect 1270 314 1276 315
rect 1390 319 1396 320
rect 1390 315 1391 319
rect 1395 315 1396 319
rect 2006 316 2007 320
rect 2011 316 2012 320
rect 2006 315 2012 316
rect 2046 320 2052 321
rect 2192 320 2194 341
rect 2328 320 2330 341
rect 2472 320 2474 341
rect 2624 320 2626 341
rect 2784 320 2786 341
rect 2952 320 2954 341
rect 3120 320 3122 341
rect 3296 320 3298 341
rect 3472 320 3474 341
rect 3656 320 3658 341
rect 3840 320 3842 341
rect 3944 321 3946 341
rect 3942 320 3948 321
rect 2046 316 2047 320
rect 2051 316 2052 320
rect 2046 315 2052 316
rect 2190 319 2196 320
rect 2190 315 2191 319
rect 2195 315 2196 319
rect 1390 314 1396 315
rect 2190 314 2196 315
rect 2326 319 2332 320
rect 2326 315 2327 319
rect 2331 315 2332 319
rect 2326 314 2332 315
rect 2470 319 2476 320
rect 2470 315 2471 319
rect 2475 315 2476 319
rect 2470 314 2476 315
rect 2622 319 2628 320
rect 2622 315 2623 319
rect 2627 315 2628 319
rect 2622 314 2628 315
rect 2782 319 2788 320
rect 2782 315 2783 319
rect 2787 315 2788 319
rect 2782 314 2788 315
rect 2950 319 2956 320
rect 2950 315 2951 319
rect 2955 315 2956 319
rect 2950 314 2956 315
rect 3118 319 3124 320
rect 3118 315 3119 319
rect 3123 315 3124 319
rect 3118 314 3124 315
rect 3294 319 3300 320
rect 3294 315 3295 319
rect 3299 315 3300 319
rect 3294 314 3300 315
rect 3470 319 3476 320
rect 3470 315 3471 319
rect 3475 315 3476 319
rect 3470 314 3476 315
rect 3654 319 3660 320
rect 3654 315 3655 319
rect 3659 315 3660 319
rect 3654 314 3660 315
rect 3838 319 3844 320
rect 3838 315 3839 319
rect 3843 315 3844 319
rect 3942 316 3943 320
rect 3947 316 3948 320
rect 3942 315 3948 316
rect 3838 314 3844 315
rect 110 303 116 304
rect 110 299 111 303
rect 115 299 116 303
rect 2006 303 2012 304
rect 110 298 116 299
rect 142 300 148 301
rect 112 267 114 298
rect 142 296 143 300
rect 147 296 148 300
rect 142 295 148 296
rect 318 300 324 301
rect 318 296 319 300
rect 323 296 324 300
rect 318 295 324 296
rect 478 300 484 301
rect 478 296 479 300
rect 483 296 484 300
rect 478 295 484 296
rect 630 300 636 301
rect 630 296 631 300
rect 635 296 636 300
rect 630 295 636 296
rect 774 300 780 301
rect 774 296 775 300
rect 779 296 780 300
rect 774 295 780 296
rect 902 300 908 301
rect 902 296 903 300
rect 907 296 908 300
rect 902 295 908 296
rect 1030 300 1036 301
rect 1030 296 1031 300
rect 1035 296 1036 300
rect 1030 295 1036 296
rect 1150 300 1156 301
rect 1150 296 1151 300
rect 1155 296 1156 300
rect 1150 295 1156 296
rect 1270 300 1276 301
rect 1270 296 1271 300
rect 1275 296 1276 300
rect 1270 295 1276 296
rect 1390 300 1396 301
rect 1390 296 1391 300
rect 1395 296 1396 300
rect 2006 299 2007 303
rect 2011 299 2012 303
rect 2006 298 2012 299
rect 2046 303 2052 304
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 3942 303 3948 304
rect 2046 298 2052 299
rect 2190 300 2196 301
rect 1390 295 1396 296
rect 144 267 146 295
rect 320 267 322 295
rect 480 267 482 295
rect 632 267 634 295
rect 776 267 778 295
rect 904 267 906 295
rect 1032 267 1034 295
rect 1152 267 1154 295
rect 1272 267 1274 295
rect 1392 267 1394 295
rect 2008 267 2010 298
rect 2048 271 2050 298
rect 2190 296 2191 300
rect 2195 296 2196 300
rect 2190 295 2196 296
rect 2326 300 2332 301
rect 2326 296 2327 300
rect 2331 296 2332 300
rect 2326 295 2332 296
rect 2470 300 2476 301
rect 2470 296 2471 300
rect 2475 296 2476 300
rect 2470 295 2476 296
rect 2622 300 2628 301
rect 2622 296 2623 300
rect 2627 296 2628 300
rect 2622 295 2628 296
rect 2782 300 2788 301
rect 2782 296 2783 300
rect 2787 296 2788 300
rect 2782 295 2788 296
rect 2950 300 2956 301
rect 2950 296 2951 300
rect 2955 296 2956 300
rect 2950 295 2956 296
rect 3118 300 3124 301
rect 3118 296 3119 300
rect 3123 296 3124 300
rect 3118 295 3124 296
rect 3294 300 3300 301
rect 3294 296 3295 300
rect 3299 296 3300 300
rect 3294 295 3300 296
rect 3470 300 3476 301
rect 3470 296 3471 300
rect 3475 296 3476 300
rect 3470 295 3476 296
rect 3654 300 3660 301
rect 3654 296 3655 300
rect 3659 296 3660 300
rect 3654 295 3660 296
rect 3838 300 3844 301
rect 3838 296 3839 300
rect 3843 296 3844 300
rect 3942 299 3943 303
rect 3947 299 3948 303
rect 3942 298 3948 299
rect 3838 295 3844 296
rect 2192 271 2194 295
rect 2328 271 2330 295
rect 2472 271 2474 295
rect 2624 271 2626 295
rect 2784 271 2786 295
rect 2952 271 2954 295
rect 3120 271 3122 295
rect 3296 271 3298 295
rect 3472 271 3474 295
rect 3656 271 3658 295
rect 3840 271 3842 295
rect 3944 271 3946 298
rect 2047 270 2051 271
rect 111 266 115 267
rect 111 261 115 262
rect 143 266 147 267
rect 143 261 147 262
rect 223 266 227 267
rect 223 261 227 262
rect 319 266 323 267
rect 319 261 323 262
rect 391 266 395 267
rect 391 261 395 262
rect 479 266 483 267
rect 479 261 483 262
rect 559 266 563 267
rect 559 261 563 262
rect 631 266 635 267
rect 631 261 635 262
rect 735 266 739 267
rect 735 261 739 262
rect 775 266 779 267
rect 775 261 779 262
rect 903 266 907 267
rect 903 261 907 262
rect 1031 266 1035 267
rect 1031 261 1035 262
rect 1063 266 1067 267
rect 1063 261 1067 262
rect 1151 266 1155 267
rect 1151 261 1155 262
rect 1215 266 1219 267
rect 1215 261 1219 262
rect 1271 266 1275 267
rect 1271 261 1275 262
rect 1359 266 1363 267
rect 1359 261 1363 262
rect 1391 266 1395 267
rect 1391 261 1395 262
rect 1511 266 1515 267
rect 1511 261 1515 262
rect 1663 266 1667 267
rect 1663 261 1667 262
rect 2007 266 2011 267
rect 2047 265 2051 266
rect 2071 270 2075 271
rect 2071 265 2075 266
rect 2191 270 2195 271
rect 2191 265 2195 266
rect 2215 270 2219 271
rect 2215 265 2219 266
rect 2327 270 2331 271
rect 2327 265 2331 266
rect 2399 270 2403 271
rect 2399 265 2403 266
rect 2471 270 2475 271
rect 2471 265 2475 266
rect 2591 270 2595 271
rect 2591 265 2595 266
rect 2623 270 2627 271
rect 2623 265 2627 266
rect 2783 270 2787 271
rect 2783 265 2787 266
rect 2791 270 2795 271
rect 2791 265 2795 266
rect 2951 270 2955 271
rect 2951 265 2955 266
rect 2983 270 2987 271
rect 2983 265 2987 266
rect 3119 270 3123 271
rect 3119 265 3123 266
rect 3167 270 3171 271
rect 3167 265 3171 266
rect 3295 270 3299 271
rect 3295 265 3299 266
rect 3343 270 3347 271
rect 3343 265 3347 266
rect 3471 270 3475 271
rect 3471 265 3475 266
rect 3511 270 3515 271
rect 3511 265 3515 266
rect 3655 270 3659 271
rect 3655 265 3659 266
rect 3687 270 3691 271
rect 3687 265 3691 266
rect 3839 270 3843 271
rect 3839 265 3843 266
rect 3943 270 3947 271
rect 3943 265 3947 266
rect 2007 261 2011 262
rect 112 234 114 261
rect 224 237 226 261
rect 392 237 394 261
rect 560 237 562 261
rect 736 237 738 261
rect 904 237 906 261
rect 1064 237 1066 261
rect 1216 237 1218 261
rect 1360 237 1362 261
rect 1512 237 1514 261
rect 1664 237 1666 261
rect 222 236 228 237
rect 110 233 116 234
rect 110 229 111 233
rect 115 229 116 233
rect 222 232 223 236
rect 227 232 228 236
rect 222 231 228 232
rect 390 236 396 237
rect 390 232 391 236
rect 395 232 396 236
rect 390 231 396 232
rect 558 236 564 237
rect 558 232 559 236
rect 563 232 564 236
rect 558 231 564 232
rect 734 236 740 237
rect 734 232 735 236
rect 739 232 740 236
rect 734 231 740 232
rect 902 236 908 237
rect 902 232 903 236
rect 907 232 908 236
rect 902 231 908 232
rect 1062 236 1068 237
rect 1062 232 1063 236
rect 1067 232 1068 236
rect 1062 231 1068 232
rect 1214 236 1220 237
rect 1214 232 1215 236
rect 1219 232 1220 236
rect 1214 231 1220 232
rect 1358 236 1364 237
rect 1358 232 1359 236
rect 1363 232 1364 236
rect 1358 231 1364 232
rect 1510 236 1516 237
rect 1510 232 1511 236
rect 1515 232 1516 236
rect 1510 231 1516 232
rect 1662 236 1668 237
rect 1662 232 1663 236
rect 1667 232 1668 236
rect 2008 234 2010 261
rect 2048 238 2050 265
rect 2072 241 2074 265
rect 2216 241 2218 265
rect 2400 241 2402 265
rect 2592 241 2594 265
rect 2792 241 2794 265
rect 2984 241 2986 265
rect 3168 241 3170 265
rect 3344 241 3346 265
rect 3512 241 3514 265
rect 3688 241 3690 265
rect 3840 241 3842 265
rect 2070 240 2076 241
rect 2046 237 2052 238
rect 1662 231 1668 232
rect 2006 233 2012 234
rect 110 228 116 229
rect 2006 229 2007 233
rect 2011 229 2012 233
rect 2046 233 2047 237
rect 2051 233 2052 237
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2214 240 2220 241
rect 2214 236 2215 240
rect 2219 236 2220 240
rect 2214 235 2220 236
rect 2398 240 2404 241
rect 2398 236 2399 240
rect 2403 236 2404 240
rect 2398 235 2404 236
rect 2590 240 2596 241
rect 2590 236 2591 240
rect 2595 236 2596 240
rect 2590 235 2596 236
rect 2790 240 2796 241
rect 2790 236 2791 240
rect 2795 236 2796 240
rect 2790 235 2796 236
rect 2982 240 2988 241
rect 2982 236 2983 240
rect 2987 236 2988 240
rect 2982 235 2988 236
rect 3166 240 3172 241
rect 3166 236 3167 240
rect 3171 236 3172 240
rect 3166 235 3172 236
rect 3342 240 3348 241
rect 3342 236 3343 240
rect 3347 236 3348 240
rect 3342 235 3348 236
rect 3510 240 3516 241
rect 3510 236 3511 240
rect 3515 236 3516 240
rect 3510 235 3516 236
rect 3686 240 3692 241
rect 3686 236 3687 240
rect 3691 236 3692 240
rect 3686 235 3692 236
rect 3838 240 3844 241
rect 3838 236 3839 240
rect 3843 236 3844 240
rect 3944 238 3946 265
rect 3838 235 3844 236
rect 3942 237 3948 238
rect 2046 232 2052 233
rect 3942 233 3943 237
rect 3947 233 3948 237
rect 3942 232 3948 233
rect 2006 228 2012 229
rect 2070 221 2076 222
rect 2046 220 2052 221
rect 222 217 228 218
rect 110 216 116 217
rect 110 212 111 216
rect 115 212 116 216
rect 222 213 223 217
rect 227 213 228 217
rect 222 212 228 213
rect 390 217 396 218
rect 390 213 391 217
rect 395 213 396 217
rect 390 212 396 213
rect 558 217 564 218
rect 558 213 559 217
rect 563 213 564 217
rect 558 212 564 213
rect 734 217 740 218
rect 734 213 735 217
rect 739 213 740 217
rect 734 212 740 213
rect 902 217 908 218
rect 902 213 903 217
rect 907 213 908 217
rect 902 212 908 213
rect 1062 217 1068 218
rect 1062 213 1063 217
rect 1067 213 1068 217
rect 1062 212 1068 213
rect 1214 217 1220 218
rect 1214 213 1215 217
rect 1219 213 1220 217
rect 1214 212 1220 213
rect 1358 217 1364 218
rect 1358 213 1359 217
rect 1363 213 1364 217
rect 1358 212 1364 213
rect 1510 217 1516 218
rect 1510 213 1511 217
rect 1515 213 1516 217
rect 1510 212 1516 213
rect 1662 217 1668 218
rect 1662 213 1663 217
rect 1667 213 1668 217
rect 1662 212 1668 213
rect 2006 216 2012 217
rect 2006 212 2007 216
rect 2011 212 2012 216
rect 2046 216 2047 220
rect 2051 216 2052 220
rect 2070 217 2071 221
rect 2075 217 2076 221
rect 2070 216 2076 217
rect 2214 221 2220 222
rect 2214 217 2215 221
rect 2219 217 2220 221
rect 2214 216 2220 217
rect 2398 221 2404 222
rect 2398 217 2399 221
rect 2403 217 2404 221
rect 2398 216 2404 217
rect 2590 221 2596 222
rect 2590 217 2591 221
rect 2595 217 2596 221
rect 2590 216 2596 217
rect 2790 221 2796 222
rect 2790 217 2791 221
rect 2795 217 2796 221
rect 2790 216 2796 217
rect 2982 221 2988 222
rect 2982 217 2983 221
rect 2987 217 2988 221
rect 2982 216 2988 217
rect 3166 221 3172 222
rect 3166 217 3167 221
rect 3171 217 3172 221
rect 3166 216 3172 217
rect 3342 221 3348 222
rect 3342 217 3343 221
rect 3347 217 3348 221
rect 3342 216 3348 217
rect 3510 221 3516 222
rect 3510 217 3511 221
rect 3515 217 3516 221
rect 3510 216 3516 217
rect 3686 221 3692 222
rect 3686 217 3687 221
rect 3691 217 3692 221
rect 3686 216 3692 217
rect 3838 221 3844 222
rect 3838 217 3839 221
rect 3843 217 3844 221
rect 3838 216 3844 217
rect 3942 220 3948 221
rect 3942 216 3943 220
rect 3947 216 3948 220
rect 2046 215 2052 216
rect 110 211 116 212
rect 112 159 114 211
rect 224 159 226 212
rect 392 159 394 212
rect 560 159 562 212
rect 736 159 738 212
rect 904 159 906 212
rect 1064 159 1066 212
rect 1216 159 1218 212
rect 1360 159 1362 212
rect 1512 159 1514 212
rect 1664 159 1666 212
rect 2006 211 2012 212
rect 2008 159 2010 211
rect 2048 171 2050 215
rect 2072 171 2074 216
rect 2216 171 2218 216
rect 2400 171 2402 216
rect 2592 171 2594 216
rect 2792 171 2794 216
rect 2984 171 2986 216
rect 3168 171 3170 216
rect 3344 171 3346 216
rect 3512 171 3514 216
rect 3688 171 3690 216
rect 3840 171 3842 216
rect 3942 215 3948 216
rect 3944 171 3946 215
rect 2047 170 2051 171
rect 2047 165 2051 166
rect 2071 170 2075 171
rect 2071 165 2075 166
rect 2191 170 2195 171
rect 2191 165 2195 166
rect 2215 170 2219 171
rect 2215 165 2219 166
rect 2343 170 2347 171
rect 2343 165 2347 166
rect 2399 170 2403 171
rect 2399 165 2403 166
rect 2495 170 2499 171
rect 2495 165 2499 166
rect 2591 170 2595 171
rect 2591 165 2595 166
rect 2647 170 2651 171
rect 2647 165 2651 166
rect 2791 170 2795 171
rect 2791 165 2795 166
rect 2799 170 2803 171
rect 2799 165 2803 166
rect 2943 170 2947 171
rect 2943 165 2947 166
rect 2983 170 2987 171
rect 2983 165 2987 166
rect 3071 170 3075 171
rect 3071 165 3075 166
rect 3167 170 3171 171
rect 3167 165 3171 166
rect 3191 170 3195 171
rect 3191 165 3195 166
rect 3311 170 3315 171
rect 3311 165 3315 166
rect 3343 170 3347 171
rect 3343 165 3347 166
rect 3423 170 3427 171
rect 3423 165 3427 166
rect 3511 170 3515 171
rect 3511 165 3515 166
rect 3527 170 3531 171
rect 3527 165 3531 166
rect 3639 170 3643 171
rect 3639 165 3643 166
rect 3687 170 3691 171
rect 3687 165 3691 166
rect 3743 170 3747 171
rect 3743 165 3747 166
rect 3839 170 3843 171
rect 3839 165 3843 166
rect 3943 170 3947 171
rect 3943 165 3947 166
rect 111 158 115 159
rect 111 153 115 154
rect 151 158 155 159
rect 151 153 155 154
rect 223 158 227 159
rect 223 153 227 154
rect 247 158 251 159
rect 247 153 251 154
rect 343 158 347 159
rect 343 153 347 154
rect 391 158 395 159
rect 391 153 395 154
rect 439 158 443 159
rect 439 153 443 154
rect 535 158 539 159
rect 535 153 539 154
rect 559 158 563 159
rect 559 153 563 154
rect 631 158 635 159
rect 631 153 635 154
rect 727 158 731 159
rect 727 153 731 154
rect 735 158 739 159
rect 735 153 739 154
rect 823 158 827 159
rect 823 153 827 154
rect 903 158 907 159
rect 903 153 907 154
rect 919 158 923 159
rect 919 153 923 154
rect 1015 158 1019 159
rect 1015 153 1019 154
rect 1063 158 1067 159
rect 1063 153 1067 154
rect 1111 158 1115 159
rect 1111 153 1115 154
rect 1207 158 1211 159
rect 1207 153 1211 154
rect 1215 158 1219 159
rect 1215 153 1219 154
rect 1303 158 1307 159
rect 1303 153 1307 154
rect 1359 158 1363 159
rect 1359 153 1363 154
rect 1407 158 1411 159
rect 1407 153 1411 154
rect 1511 158 1515 159
rect 1511 153 1515 154
rect 1615 158 1619 159
rect 1615 153 1619 154
rect 1663 158 1667 159
rect 1663 153 1667 154
rect 1711 158 1715 159
rect 1711 153 1715 154
rect 1807 158 1811 159
rect 1807 153 1811 154
rect 1903 158 1907 159
rect 1903 153 1907 154
rect 2007 158 2011 159
rect 2007 153 2011 154
rect 112 133 114 153
rect 110 132 116 133
rect 152 132 154 153
rect 248 132 250 153
rect 344 132 346 153
rect 440 132 442 153
rect 536 132 538 153
rect 632 132 634 153
rect 728 132 730 153
rect 824 132 826 153
rect 920 132 922 153
rect 1016 132 1018 153
rect 1112 132 1114 153
rect 1208 132 1210 153
rect 1304 132 1306 153
rect 1408 132 1410 153
rect 1512 132 1514 153
rect 1616 132 1618 153
rect 1712 132 1714 153
rect 1808 132 1810 153
rect 1904 132 1906 153
rect 2008 133 2010 153
rect 2048 145 2050 165
rect 2046 144 2052 145
rect 2072 144 2074 165
rect 2192 144 2194 165
rect 2344 144 2346 165
rect 2496 144 2498 165
rect 2648 144 2650 165
rect 2800 144 2802 165
rect 2944 144 2946 165
rect 3072 144 3074 165
rect 3192 144 3194 165
rect 3312 144 3314 165
rect 3424 144 3426 165
rect 3528 144 3530 165
rect 3640 144 3642 165
rect 3744 144 3746 165
rect 3840 144 3842 165
rect 3944 145 3946 165
rect 3942 144 3948 145
rect 2046 140 2047 144
rect 2051 140 2052 144
rect 2046 139 2052 140
rect 2070 143 2076 144
rect 2070 139 2071 143
rect 2075 139 2076 143
rect 2070 138 2076 139
rect 2190 143 2196 144
rect 2190 139 2191 143
rect 2195 139 2196 143
rect 2190 138 2196 139
rect 2342 143 2348 144
rect 2342 139 2343 143
rect 2347 139 2348 143
rect 2342 138 2348 139
rect 2494 143 2500 144
rect 2494 139 2495 143
rect 2499 139 2500 143
rect 2494 138 2500 139
rect 2646 143 2652 144
rect 2646 139 2647 143
rect 2651 139 2652 143
rect 2646 138 2652 139
rect 2798 143 2804 144
rect 2798 139 2799 143
rect 2803 139 2804 143
rect 2798 138 2804 139
rect 2942 143 2948 144
rect 2942 139 2943 143
rect 2947 139 2948 143
rect 2942 138 2948 139
rect 3070 143 3076 144
rect 3070 139 3071 143
rect 3075 139 3076 143
rect 3070 138 3076 139
rect 3190 143 3196 144
rect 3190 139 3191 143
rect 3195 139 3196 143
rect 3190 138 3196 139
rect 3310 143 3316 144
rect 3310 139 3311 143
rect 3315 139 3316 143
rect 3310 138 3316 139
rect 3422 143 3428 144
rect 3422 139 3423 143
rect 3427 139 3428 143
rect 3422 138 3428 139
rect 3526 143 3532 144
rect 3526 139 3527 143
rect 3531 139 3532 143
rect 3526 138 3532 139
rect 3638 143 3644 144
rect 3638 139 3639 143
rect 3643 139 3644 143
rect 3638 138 3644 139
rect 3742 143 3748 144
rect 3742 139 3743 143
rect 3747 139 3748 143
rect 3742 138 3748 139
rect 3838 143 3844 144
rect 3838 139 3839 143
rect 3843 139 3844 143
rect 3942 140 3943 144
rect 3947 140 3948 144
rect 3942 139 3948 140
rect 3838 138 3844 139
rect 2006 132 2012 133
rect 110 128 111 132
rect 115 128 116 132
rect 110 127 116 128
rect 150 131 156 132
rect 150 127 151 131
rect 155 127 156 131
rect 150 126 156 127
rect 246 131 252 132
rect 246 127 247 131
rect 251 127 252 131
rect 246 126 252 127
rect 342 131 348 132
rect 342 127 343 131
rect 347 127 348 131
rect 342 126 348 127
rect 438 131 444 132
rect 438 127 439 131
rect 443 127 444 131
rect 438 126 444 127
rect 534 131 540 132
rect 534 127 535 131
rect 539 127 540 131
rect 534 126 540 127
rect 630 131 636 132
rect 630 127 631 131
rect 635 127 636 131
rect 630 126 636 127
rect 726 131 732 132
rect 726 127 727 131
rect 731 127 732 131
rect 726 126 732 127
rect 822 131 828 132
rect 822 127 823 131
rect 827 127 828 131
rect 822 126 828 127
rect 918 131 924 132
rect 918 127 919 131
rect 923 127 924 131
rect 918 126 924 127
rect 1014 131 1020 132
rect 1014 127 1015 131
rect 1019 127 1020 131
rect 1014 126 1020 127
rect 1110 131 1116 132
rect 1110 127 1111 131
rect 1115 127 1116 131
rect 1110 126 1116 127
rect 1206 131 1212 132
rect 1206 127 1207 131
rect 1211 127 1212 131
rect 1206 126 1212 127
rect 1302 131 1308 132
rect 1302 127 1303 131
rect 1307 127 1308 131
rect 1302 126 1308 127
rect 1406 131 1412 132
rect 1406 127 1407 131
rect 1411 127 1412 131
rect 1406 126 1412 127
rect 1510 131 1516 132
rect 1510 127 1511 131
rect 1515 127 1516 131
rect 1510 126 1516 127
rect 1614 131 1620 132
rect 1614 127 1615 131
rect 1619 127 1620 131
rect 1614 126 1620 127
rect 1710 131 1716 132
rect 1710 127 1711 131
rect 1715 127 1716 131
rect 1710 126 1716 127
rect 1806 131 1812 132
rect 1806 127 1807 131
rect 1811 127 1812 131
rect 1806 126 1812 127
rect 1902 131 1908 132
rect 1902 127 1903 131
rect 1907 127 1908 131
rect 2006 128 2007 132
rect 2011 128 2012 132
rect 2006 127 2012 128
rect 2046 127 2052 128
rect 1902 126 1908 127
rect 2046 123 2047 127
rect 2051 123 2052 127
rect 3942 127 3948 128
rect 2046 122 2052 123
rect 2070 124 2076 125
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 2006 115 2012 116
rect 110 110 116 111
rect 150 112 156 113
rect 112 83 114 110
rect 150 108 151 112
rect 155 108 156 112
rect 150 107 156 108
rect 246 112 252 113
rect 246 108 247 112
rect 251 108 252 112
rect 246 107 252 108
rect 342 112 348 113
rect 342 108 343 112
rect 347 108 348 112
rect 342 107 348 108
rect 438 112 444 113
rect 438 108 439 112
rect 443 108 444 112
rect 438 107 444 108
rect 534 112 540 113
rect 534 108 535 112
rect 539 108 540 112
rect 534 107 540 108
rect 630 112 636 113
rect 630 108 631 112
rect 635 108 636 112
rect 630 107 636 108
rect 726 112 732 113
rect 726 108 727 112
rect 731 108 732 112
rect 726 107 732 108
rect 822 112 828 113
rect 822 108 823 112
rect 827 108 828 112
rect 822 107 828 108
rect 918 112 924 113
rect 918 108 919 112
rect 923 108 924 112
rect 918 107 924 108
rect 1014 112 1020 113
rect 1014 108 1015 112
rect 1019 108 1020 112
rect 1014 107 1020 108
rect 1110 112 1116 113
rect 1110 108 1111 112
rect 1115 108 1116 112
rect 1110 107 1116 108
rect 1206 112 1212 113
rect 1206 108 1207 112
rect 1211 108 1212 112
rect 1206 107 1212 108
rect 1302 112 1308 113
rect 1302 108 1303 112
rect 1307 108 1308 112
rect 1302 107 1308 108
rect 1406 112 1412 113
rect 1406 108 1407 112
rect 1411 108 1412 112
rect 1406 107 1412 108
rect 1510 112 1516 113
rect 1510 108 1511 112
rect 1515 108 1516 112
rect 1510 107 1516 108
rect 1614 112 1620 113
rect 1614 108 1615 112
rect 1619 108 1620 112
rect 1614 107 1620 108
rect 1710 112 1716 113
rect 1710 108 1711 112
rect 1715 108 1716 112
rect 1710 107 1716 108
rect 1806 112 1812 113
rect 1806 108 1807 112
rect 1811 108 1812 112
rect 1806 107 1812 108
rect 1902 112 1908 113
rect 1902 108 1903 112
rect 1907 108 1908 112
rect 2006 111 2007 115
rect 2011 111 2012 115
rect 2006 110 2012 111
rect 1902 107 1908 108
rect 152 83 154 107
rect 248 83 250 107
rect 344 83 346 107
rect 440 83 442 107
rect 536 83 538 107
rect 632 83 634 107
rect 728 83 730 107
rect 824 83 826 107
rect 920 83 922 107
rect 1016 83 1018 107
rect 1112 83 1114 107
rect 1208 83 1210 107
rect 1304 83 1306 107
rect 1408 83 1410 107
rect 1512 83 1514 107
rect 1616 83 1618 107
rect 1712 83 1714 107
rect 1808 83 1810 107
rect 1904 83 1906 107
rect 2008 83 2010 110
rect 2048 95 2050 122
rect 2070 120 2071 124
rect 2075 120 2076 124
rect 2070 119 2076 120
rect 2190 124 2196 125
rect 2190 120 2191 124
rect 2195 120 2196 124
rect 2190 119 2196 120
rect 2342 124 2348 125
rect 2342 120 2343 124
rect 2347 120 2348 124
rect 2342 119 2348 120
rect 2494 124 2500 125
rect 2494 120 2495 124
rect 2499 120 2500 124
rect 2494 119 2500 120
rect 2646 124 2652 125
rect 2646 120 2647 124
rect 2651 120 2652 124
rect 2646 119 2652 120
rect 2798 124 2804 125
rect 2798 120 2799 124
rect 2803 120 2804 124
rect 2798 119 2804 120
rect 2942 124 2948 125
rect 2942 120 2943 124
rect 2947 120 2948 124
rect 2942 119 2948 120
rect 3070 124 3076 125
rect 3070 120 3071 124
rect 3075 120 3076 124
rect 3070 119 3076 120
rect 3190 124 3196 125
rect 3190 120 3191 124
rect 3195 120 3196 124
rect 3190 119 3196 120
rect 3310 124 3316 125
rect 3310 120 3311 124
rect 3315 120 3316 124
rect 3310 119 3316 120
rect 3422 124 3428 125
rect 3422 120 3423 124
rect 3427 120 3428 124
rect 3422 119 3428 120
rect 3526 124 3532 125
rect 3526 120 3527 124
rect 3531 120 3532 124
rect 3526 119 3532 120
rect 3638 124 3644 125
rect 3638 120 3639 124
rect 3643 120 3644 124
rect 3638 119 3644 120
rect 3742 124 3748 125
rect 3742 120 3743 124
rect 3747 120 3748 124
rect 3742 119 3748 120
rect 3838 124 3844 125
rect 3838 120 3839 124
rect 3843 120 3844 124
rect 3942 123 3943 127
rect 3947 123 3948 127
rect 3942 122 3948 123
rect 3838 119 3844 120
rect 2072 95 2074 119
rect 2192 95 2194 119
rect 2344 95 2346 119
rect 2496 95 2498 119
rect 2648 95 2650 119
rect 2800 95 2802 119
rect 2944 95 2946 119
rect 3072 95 3074 119
rect 3192 95 3194 119
rect 3312 95 3314 119
rect 3424 95 3426 119
rect 3528 95 3530 119
rect 3640 95 3642 119
rect 3744 95 3746 119
rect 3840 95 3842 119
rect 3944 95 3946 122
rect 2047 94 2051 95
rect 2047 89 2051 90
rect 2071 94 2075 95
rect 2071 89 2075 90
rect 2191 94 2195 95
rect 2191 89 2195 90
rect 2343 94 2347 95
rect 2343 89 2347 90
rect 2495 94 2499 95
rect 2495 89 2499 90
rect 2647 94 2651 95
rect 2647 89 2651 90
rect 2799 94 2803 95
rect 2799 89 2803 90
rect 2943 94 2947 95
rect 2943 89 2947 90
rect 3071 94 3075 95
rect 3071 89 3075 90
rect 3191 94 3195 95
rect 3191 89 3195 90
rect 3311 94 3315 95
rect 3311 89 3315 90
rect 3423 94 3427 95
rect 3423 89 3427 90
rect 3527 94 3531 95
rect 3527 89 3531 90
rect 3639 94 3643 95
rect 3639 89 3643 90
rect 3743 94 3747 95
rect 3743 89 3747 90
rect 3839 94 3843 95
rect 3839 89 3843 90
rect 3943 94 3947 95
rect 3943 89 3947 90
rect 111 82 115 83
rect 111 77 115 78
rect 151 82 155 83
rect 151 77 155 78
rect 247 82 251 83
rect 247 77 251 78
rect 343 82 347 83
rect 343 77 347 78
rect 439 82 443 83
rect 439 77 443 78
rect 535 82 539 83
rect 535 77 539 78
rect 631 82 635 83
rect 631 77 635 78
rect 727 82 731 83
rect 727 77 731 78
rect 823 82 827 83
rect 823 77 827 78
rect 919 82 923 83
rect 919 77 923 78
rect 1015 82 1019 83
rect 1015 77 1019 78
rect 1111 82 1115 83
rect 1111 77 1115 78
rect 1207 82 1211 83
rect 1207 77 1211 78
rect 1303 82 1307 83
rect 1303 77 1307 78
rect 1407 82 1411 83
rect 1407 77 1411 78
rect 1511 82 1515 83
rect 1511 77 1515 78
rect 1615 82 1619 83
rect 1615 77 1619 78
rect 1711 82 1715 83
rect 1711 77 1715 78
rect 1807 82 1811 83
rect 1807 77 1811 78
rect 1903 82 1907 83
rect 1903 77 1907 78
rect 2007 82 2011 83
rect 2007 77 2011 78
<< m4c >>
rect 2047 4018 2051 4022
rect 2071 4018 2075 4022
rect 2327 4018 2331 4022
rect 2591 4018 2595 4022
rect 2839 4018 2843 4022
rect 3087 4018 3091 4022
rect 3343 4018 3347 4022
rect 3943 4018 3947 4022
rect 111 3998 115 4002
rect 311 3998 315 4002
rect 511 3998 515 4002
rect 703 3998 707 4002
rect 887 3998 891 4002
rect 1063 3998 1067 4002
rect 1231 3998 1235 4002
rect 1383 3998 1387 4002
rect 1519 3998 1523 4002
rect 1655 3998 1659 4002
rect 1791 3998 1795 4002
rect 1903 3998 1907 4002
rect 2007 3998 2011 4002
rect 2047 3942 2051 3946
rect 2071 3942 2075 3946
rect 2127 3942 2131 3946
rect 2271 3942 2275 3946
rect 2327 3942 2331 3946
rect 2439 3942 2443 3946
rect 2591 3942 2595 3946
rect 2615 3942 2619 3946
rect 2799 3942 2803 3946
rect 2839 3942 2843 3946
rect 2983 3942 2987 3946
rect 3087 3942 3091 3946
rect 3175 3942 3179 3946
rect 3343 3942 3347 3946
rect 3367 3942 3371 3946
rect 3559 3942 3563 3946
rect 3943 3942 3947 3946
rect 111 3922 115 3926
rect 279 3922 283 3926
rect 311 3922 315 3926
rect 415 3922 419 3926
rect 511 3922 515 3926
rect 567 3922 571 3926
rect 703 3922 707 3926
rect 735 3922 739 3926
rect 887 3922 891 3926
rect 911 3922 915 3926
rect 1063 3922 1067 3926
rect 1095 3922 1099 3926
rect 1231 3922 1235 3926
rect 1287 3922 1291 3926
rect 1383 3922 1387 3926
rect 1479 3922 1483 3926
rect 1519 3922 1523 3926
rect 1655 3922 1659 3926
rect 1679 3922 1683 3926
rect 1791 3922 1795 3926
rect 1903 3922 1907 3926
rect 2007 3922 2011 3926
rect 2047 3866 2051 3870
rect 2127 3866 2131 3870
rect 2263 3866 2267 3870
rect 2271 3866 2275 3870
rect 2375 3866 2379 3870
rect 2439 3866 2443 3870
rect 2495 3866 2499 3870
rect 2615 3866 2619 3870
rect 2631 3866 2635 3870
rect 2775 3866 2779 3870
rect 2799 3866 2803 3870
rect 2919 3866 2923 3870
rect 2983 3866 2987 3870
rect 3063 3866 3067 3870
rect 3175 3866 3179 3870
rect 3207 3866 3211 3870
rect 3343 3866 3347 3870
rect 3367 3866 3371 3870
rect 3471 3866 3475 3870
rect 3559 3866 3563 3870
rect 3599 3866 3603 3870
rect 3727 3866 3731 3870
rect 3839 3866 3843 3870
rect 3943 3866 3947 3870
rect 111 3838 115 3842
rect 231 3838 235 3842
rect 279 3838 283 3842
rect 335 3838 339 3842
rect 415 3838 419 3842
rect 439 3838 443 3842
rect 535 3838 539 3842
rect 567 3838 571 3842
rect 631 3838 635 3842
rect 727 3838 731 3842
rect 735 3838 739 3842
rect 831 3838 835 3842
rect 911 3838 915 3842
rect 935 3838 939 3842
rect 1039 3838 1043 3842
rect 1095 3838 1099 3842
rect 1151 3838 1155 3842
rect 1263 3838 1267 3842
rect 1287 3838 1291 3842
rect 1383 3838 1387 3842
rect 1479 3838 1483 3842
rect 1503 3838 1507 3842
rect 1631 3838 1635 3842
rect 1679 3838 1683 3842
rect 2007 3838 2011 3842
rect 2047 3774 2051 3778
rect 2071 3774 2075 3778
rect 2183 3774 2187 3778
rect 2263 3774 2267 3778
rect 2327 3774 2331 3778
rect 2375 3774 2379 3778
rect 2479 3774 2483 3778
rect 2495 3774 2499 3778
rect 2631 3774 2635 3778
rect 2639 3774 2643 3778
rect 2775 3774 2779 3778
rect 2807 3774 2811 3778
rect 2919 3774 2923 3778
rect 2983 3774 2987 3778
rect 3063 3774 3067 3778
rect 3159 3774 3163 3778
rect 3207 3774 3211 3778
rect 3335 3774 3339 3778
rect 3343 3774 3347 3778
rect 3471 3774 3475 3778
rect 3511 3774 3515 3778
rect 3599 3774 3603 3778
rect 3687 3774 3691 3778
rect 3727 3774 3731 3778
rect 3839 3774 3843 3778
rect 3943 3774 3947 3778
rect 111 3762 115 3766
rect 159 3762 163 3766
rect 231 3762 235 3766
rect 335 3762 339 3766
rect 351 3762 355 3766
rect 439 3762 443 3766
rect 535 3762 539 3766
rect 551 3762 555 3766
rect 631 3762 635 3766
rect 727 3762 731 3766
rect 751 3762 755 3766
rect 831 3762 835 3766
rect 935 3762 939 3766
rect 959 3762 963 3766
rect 1039 3762 1043 3766
rect 1151 3762 1155 3766
rect 1167 3762 1171 3766
rect 1263 3762 1267 3766
rect 1383 3762 1387 3766
rect 1503 3762 1507 3766
rect 1607 3762 1611 3766
rect 1631 3762 1635 3766
rect 2007 3762 2011 3766
rect 2047 3686 2051 3690
rect 2071 3686 2075 3690
rect 2183 3686 2187 3690
rect 2199 3686 2203 3690
rect 2327 3686 2331 3690
rect 2367 3686 2371 3690
rect 2479 3686 2483 3690
rect 2551 3686 2555 3690
rect 2639 3686 2643 3690
rect 2735 3686 2739 3690
rect 2807 3686 2811 3690
rect 2927 3686 2931 3690
rect 2983 3686 2987 3690
rect 3111 3686 3115 3690
rect 3159 3686 3163 3690
rect 3295 3686 3299 3690
rect 3335 3686 3339 3690
rect 3479 3686 3483 3690
rect 3511 3686 3515 3690
rect 3671 3686 3675 3690
rect 3687 3686 3691 3690
rect 3839 3686 3843 3690
rect 3943 3686 3947 3690
rect 111 3678 115 3682
rect 151 3678 155 3682
rect 159 3678 163 3682
rect 351 3678 355 3682
rect 383 3678 387 3682
rect 551 3678 555 3682
rect 615 3678 619 3682
rect 751 3678 755 3682
rect 839 3678 843 3682
rect 959 3678 963 3682
rect 1055 3678 1059 3682
rect 1167 3678 1171 3682
rect 1263 3678 1267 3682
rect 1383 3678 1387 3682
rect 1479 3678 1483 3682
rect 1607 3678 1611 3682
rect 1695 3678 1699 3682
rect 2007 3678 2011 3682
rect 2047 3606 2051 3610
rect 2071 3606 2075 3610
rect 2103 3606 2107 3610
rect 2199 3606 2203 3610
rect 2279 3606 2283 3610
rect 2367 3606 2371 3610
rect 2471 3606 2475 3610
rect 2551 3606 2555 3610
rect 2671 3606 2675 3610
rect 2735 3606 2739 3610
rect 2871 3606 2875 3610
rect 2927 3606 2931 3610
rect 3063 3606 3067 3610
rect 3111 3606 3115 3610
rect 3255 3606 3259 3610
rect 3295 3606 3299 3610
rect 3447 3606 3451 3610
rect 3479 3606 3483 3610
rect 3639 3606 3643 3610
rect 3671 3606 3675 3610
rect 3839 3606 3843 3610
rect 3943 3606 3947 3610
rect 111 3598 115 3602
rect 151 3598 155 3602
rect 167 3598 171 3602
rect 359 3598 363 3602
rect 383 3598 387 3602
rect 559 3598 563 3602
rect 615 3598 619 3602
rect 775 3598 779 3602
rect 839 3598 843 3602
rect 991 3598 995 3602
rect 1055 3598 1059 3602
rect 1215 3598 1219 3602
rect 1263 3598 1267 3602
rect 1447 3598 1451 3602
rect 1479 3598 1483 3602
rect 1687 3598 1691 3602
rect 1695 3598 1699 3602
rect 2007 3598 2011 3602
rect 2047 3526 2051 3530
rect 2103 3526 2107 3530
rect 2279 3526 2283 3530
rect 2327 3526 2331 3530
rect 2447 3526 2451 3530
rect 2471 3526 2475 3530
rect 2583 3526 2587 3530
rect 2671 3526 2675 3530
rect 2735 3526 2739 3530
rect 2871 3526 2875 3530
rect 2911 3526 2915 3530
rect 3063 3526 3067 3530
rect 3111 3526 3115 3530
rect 3255 3526 3259 3530
rect 3335 3526 3339 3530
rect 3447 3526 3451 3530
rect 3567 3526 3571 3530
rect 3639 3526 3643 3530
rect 3807 3526 3811 3530
rect 3839 3526 3843 3530
rect 3943 3526 3947 3530
rect 111 3514 115 3518
rect 167 3514 171 3518
rect 295 3514 299 3518
rect 359 3514 363 3518
rect 431 3514 435 3518
rect 559 3514 563 3518
rect 583 3514 587 3518
rect 743 3514 747 3518
rect 775 3514 779 3518
rect 911 3514 915 3518
rect 991 3514 995 3518
rect 1079 3514 1083 3518
rect 1215 3514 1219 3518
rect 1247 3514 1251 3518
rect 1423 3514 1427 3518
rect 1447 3514 1451 3518
rect 1599 3514 1603 3518
rect 1687 3514 1691 3518
rect 1775 3514 1779 3518
rect 2007 3514 2011 3518
rect 2047 3450 2051 3454
rect 2327 3450 2331 3454
rect 2447 3450 2451 3454
rect 2551 3450 2555 3454
rect 2583 3450 2587 3454
rect 2663 3450 2667 3454
rect 2735 3450 2739 3454
rect 2775 3450 2779 3454
rect 2903 3450 2907 3454
rect 2911 3450 2915 3454
rect 3047 3450 3051 3454
rect 3111 3450 3115 3454
rect 3207 3450 3211 3454
rect 3335 3450 3339 3454
rect 3383 3450 3387 3454
rect 3567 3450 3571 3454
rect 3751 3450 3755 3454
rect 3807 3450 3811 3454
rect 3943 3450 3947 3454
rect 111 3418 115 3422
rect 295 3418 299 3422
rect 431 3418 435 3422
rect 495 3418 499 3422
rect 583 3418 587 3422
rect 647 3418 651 3422
rect 743 3418 747 3422
rect 799 3418 803 3422
rect 911 3418 915 3422
rect 959 3418 963 3422
rect 1079 3418 1083 3422
rect 1127 3418 1131 3422
rect 1247 3418 1251 3422
rect 1295 3418 1299 3422
rect 1423 3418 1427 3422
rect 1463 3418 1467 3422
rect 1599 3418 1603 3422
rect 1639 3418 1643 3422
rect 1775 3418 1779 3422
rect 1815 3418 1819 3422
rect 2007 3418 2011 3422
rect 2047 3362 2051 3366
rect 2447 3362 2451 3366
rect 2551 3362 2555 3366
rect 2567 3362 2571 3366
rect 2663 3362 2667 3366
rect 2719 3362 2723 3366
rect 2775 3362 2779 3366
rect 2871 3362 2875 3366
rect 2903 3362 2907 3366
rect 3023 3362 3027 3366
rect 3047 3362 3051 3366
rect 3175 3362 3179 3366
rect 3207 3362 3211 3366
rect 3327 3362 3331 3366
rect 3383 3362 3387 3366
rect 3479 3362 3483 3366
rect 3567 3362 3571 3366
rect 3631 3362 3635 3366
rect 3751 3362 3755 3366
rect 3783 3362 3787 3366
rect 3943 3362 3947 3366
rect 111 3330 115 3334
rect 135 3330 139 3334
rect 295 3330 299 3334
rect 479 3330 483 3334
rect 495 3330 499 3334
rect 647 3330 651 3334
rect 671 3330 675 3334
rect 799 3330 803 3334
rect 863 3330 867 3334
rect 959 3330 963 3334
rect 1055 3330 1059 3334
rect 1127 3330 1131 3334
rect 1247 3330 1251 3334
rect 1295 3330 1299 3334
rect 1439 3330 1443 3334
rect 1463 3330 1467 3334
rect 1631 3330 1635 3334
rect 1639 3330 1643 3334
rect 1815 3330 1819 3334
rect 1823 3330 1827 3334
rect 2007 3330 2011 3334
rect 2047 3282 2051 3286
rect 2415 3282 2419 3286
rect 2551 3282 2555 3286
rect 2567 3282 2571 3286
rect 2687 3282 2691 3286
rect 2719 3282 2723 3286
rect 2831 3282 2835 3286
rect 2871 3282 2875 3286
rect 2975 3282 2979 3286
rect 3023 3282 3027 3286
rect 3119 3282 3123 3286
rect 3175 3282 3179 3286
rect 3255 3282 3259 3286
rect 3327 3282 3331 3286
rect 3383 3282 3387 3286
rect 3479 3282 3483 3286
rect 3503 3282 3507 3286
rect 3623 3282 3627 3286
rect 3631 3282 3635 3286
rect 3743 3282 3747 3286
rect 3783 3282 3787 3286
rect 3839 3282 3843 3286
rect 3943 3282 3947 3286
rect 111 3250 115 3254
rect 135 3250 139 3254
rect 295 3250 299 3254
rect 319 3250 323 3254
rect 479 3250 483 3254
rect 519 3250 523 3254
rect 671 3250 675 3254
rect 719 3250 723 3254
rect 863 3250 867 3254
rect 911 3250 915 3254
rect 1055 3250 1059 3254
rect 1095 3250 1099 3254
rect 1247 3250 1251 3254
rect 1271 3250 1275 3254
rect 1439 3250 1443 3254
rect 1447 3250 1451 3254
rect 1623 3250 1627 3254
rect 1631 3250 1635 3254
rect 1799 3250 1803 3254
rect 1823 3250 1827 3254
rect 2007 3250 2011 3254
rect 2047 3194 2051 3198
rect 2247 3194 2251 3198
rect 2399 3194 2403 3198
rect 2415 3194 2419 3198
rect 2551 3194 2555 3198
rect 2559 3194 2563 3198
rect 2687 3194 2691 3198
rect 2727 3194 2731 3198
rect 2831 3194 2835 3198
rect 2903 3194 2907 3198
rect 2975 3194 2979 3198
rect 3079 3194 3083 3198
rect 3119 3194 3123 3198
rect 3255 3194 3259 3198
rect 3263 3194 3267 3198
rect 3383 3194 3387 3198
rect 3447 3194 3451 3198
rect 3503 3194 3507 3198
rect 3623 3194 3627 3198
rect 3631 3194 3635 3198
rect 3743 3194 3747 3198
rect 3815 3194 3819 3198
rect 3839 3194 3843 3198
rect 3943 3194 3947 3198
rect 111 3166 115 3170
rect 135 3166 139 3170
rect 143 3166 147 3170
rect 319 3166 323 3170
rect 343 3166 347 3170
rect 519 3166 523 3170
rect 543 3166 547 3170
rect 719 3166 723 3170
rect 743 3166 747 3170
rect 911 3166 915 3170
rect 927 3166 931 3170
rect 1095 3166 1099 3170
rect 1103 3166 1107 3170
rect 1263 3166 1267 3170
rect 1271 3166 1275 3170
rect 1423 3166 1427 3170
rect 1447 3166 1451 3170
rect 1575 3166 1579 3170
rect 1623 3166 1627 3170
rect 1735 3166 1739 3170
rect 1799 3166 1803 3170
rect 2007 3166 2011 3170
rect 2047 3114 2051 3118
rect 2079 3114 2083 3118
rect 2223 3114 2227 3118
rect 2247 3114 2251 3118
rect 2375 3114 2379 3118
rect 2399 3114 2403 3118
rect 2527 3114 2531 3118
rect 2559 3114 2563 3118
rect 2687 3114 2691 3118
rect 2727 3114 2731 3118
rect 2855 3114 2859 3118
rect 2903 3114 2907 3118
rect 3039 3114 3043 3118
rect 3079 3114 3083 3118
rect 3231 3114 3235 3118
rect 3263 3114 3267 3118
rect 3431 3114 3435 3118
rect 3447 3114 3451 3118
rect 3631 3114 3635 3118
rect 3639 3114 3643 3118
rect 3815 3114 3819 3118
rect 3839 3114 3843 3118
rect 3943 3114 3947 3118
rect 111 3090 115 3094
rect 143 3090 147 3094
rect 263 3090 267 3094
rect 343 3090 347 3094
rect 439 3090 443 3094
rect 543 3090 547 3094
rect 615 3090 619 3094
rect 743 3090 747 3094
rect 799 3090 803 3094
rect 927 3090 931 3094
rect 975 3090 979 3094
rect 1103 3090 1107 3094
rect 1143 3090 1147 3094
rect 1263 3090 1267 3094
rect 1303 3090 1307 3094
rect 1423 3090 1427 3094
rect 1455 3090 1459 3094
rect 1575 3090 1579 3094
rect 1607 3090 1611 3094
rect 1735 3090 1739 3094
rect 1767 3090 1771 3094
rect 2007 3090 2011 3094
rect 2047 3030 2051 3034
rect 2071 3030 2075 3034
rect 2079 3030 2083 3034
rect 2183 3030 2187 3034
rect 2223 3030 2227 3034
rect 2327 3030 2331 3034
rect 2375 3030 2379 3034
rect 2479 3030 2483 3034
rect 2527 3030 2531 3034
rect 2655 3030 2659 3034
rect 2687 3030 2691 3034
rect 2855 3030 2859 3034
rect 3039 3030 3043 3034
rect 3087 3030 3091 3034
rect 3231 3030 3235 3034
rect 3335 3030 3339 3034
rect 3431 3030 3435 3034
rect 3599 3030 3603 3034
rect 3639 3030 3643 3034
rect 3839 3030 3843 3034
rect 3943 3030 3947 3034
rect 111 2990 115 2994
rect 263 2990 267 2994
rect 343 2990 347 2994
rect 439 2990 443 2994
rect 543 2990 547 2994
rect 615 2990 619 2994
rect 655 2990 659 2994
rect 783 2990 787 2994
rect 799 2990 803 2994
rect 935 2990 939 2994
rect 975 2990 979 2994
rect 1103 2990 1107 2994
rect 1143 2990 1147 2994
rect 1295 2990 1299 2994
rect 1303 2990 1307 2994
rect 1455 2990 1459 2994
rect 1495 2990 1499 2994
rect 1607 2990 1611 2994
rect 1711 2990 1715 2994
rect 1767 2990 1771 2994
rect 1903 2990 1907 2994
rect 2007 2990 2011 2994
rect 2047 2950 2051 2954
rect 2071 2950 2075 2954
rect 2183 2950 2187 2954
rect 2263 2950 2267 2954
rect 2327 2950 2331 2954
rect 2479 2950 2483 2954
rect 2487 2950 2491 2954
rect 2655 2950 2659 2954
rect 2735 2950 2739 2954
rect 2855 2950 2859 2954
rect 2999 2950 3003 2954
rect 3087 2950 3091 2954
rect 3279 2950 3283 2954
rect 3335 2950 3339 2954
rect 3567 2950 3571 2954
rect 3599 2950 3603 2954
rect 3839 2950 3843 2954
rect 3943 2950 3947 2954
rect 111 2914 115 2918
rect 207 2914 211 2918
rect 327 2914 331 2918
rect 343 2914 347 2918
rect 439 2914 443 2918
rect 447 2914 451 2918
rect 543 2914 547 2918
rect 575 2914 579 2918
rect 655 2914 659 2918
rect 703 2914 707 2918
rect 783 2914 787 2918
rect 847 2914 851 2918
rect 935 2914 939 2918
rect 999 2914 1003 2918
rect 1103 2914 1107 2918
rect 1167 2914 1171 2918
rect 1295 2914 1299 2918
rect 1351 2914 1355 2918
rect 1495 2914 1499 2918
rect 1535 2914 1539 2918
rect 1711 2914 1715 2918
rect 1727 2914 1731 2918
rect 1903 2914 1907 2918
rect 2007 2914 2011 2918
rect 2047 2866 2051 2870
rect 2071 2866 2075 2870
rect 2263 2866 2267 2870
rect 2487 2866 2491 2870
rect 2671 2866 2675 2870
rect 2735 2866 2739 2870
rect 2887 2866 2891 2870
rect 2999 2866 3003 2870
rect 3095 2866 3099 2870
rect 3279 2866 3283 2870
rect 3287 2866 3291 2870
rect 3479 2866 3483 2870
rect 3567 2866 3571 2870
rect 3671 2866 3675 2870
rect 3839 2866 3843 2870
rect 3943 2866 3947 2870
rect 111 2834 115 2838
rect 135 2834 139 2838
rect 207 2834 211 2838
rect 247 2834 251 2838
rect 327 2834 331 2838
rect 399 2834 403 2838
rect 447 2834 451 2838
rect 551 2834 555 2838
rect 575 2834 579 2838
rect 703 2834 707 2838
rect 711 2834 715 2838
rect 847 2834 851 2838
rect 879 2834 883 2838
rect 999 2834 1003 2838
rect 1047 2834 1051 2838
rect 1167 2834 1171 2838
rect 1223 2834 1227 2838
rect 1351 2834 1355 2838
rect 1399 2834 1403 2838
rect 1535 2834 1539 2838
rect 1575 2834 1579 2838
rect 1727 2834 1731 2838
rect 1751 2834 1755 2838
rect 1903 2834 1907 2838
rect 2007 2834 2011 2838
rect 2047 2790 2051 2794
rect 2071 2790 2075 2794
rect 2199 2790 2203 2794
rect 2343 2790 2347 2794
rect 2479 2790 2483 2794
rect 2607 2790 2611 2794
rect 2671 2790 2675 2794
rect 2727 2790 2731 2794
rect 2839 2790 2843 2794
rect 2887 2790 2891 2794
rect 2943 2790 2947 2794
rect 3047 2790 3051 2794
rect 3095 2790 3099 2794
rect 3143 2790 3147 2794
rect 3239 2790 3243 2794
rect 3287 2790 3291 2794
rect 3343 2790 3347 2794
rect 3447 2790 3451 2794
rect 3479 2790 3483 2794
rect 3551 2790 3555 2794
rect 3647 2790 3651 2794
rect 3671 2790 3675 2794
rect 3743 2790 3747 2794
rect 3839 2790 3843 2794
rect 3943 2790 3947 2794
rect 111 2750 115 2754
rect 135 2750 139 2754
rect 247 2750 251 2754
rect 255 2750 259 2754
rect 399 2750 403 2754
rect 407 2750 411 2754
rect 551 2750 555 2754
rect 575 2750 579 2754
rect 711 2750 715 2754
rect 743 2750 747 2754
rect 879 2750 883 2754
rect 919 2750 923 2754
rect 1047 2750 1051 2754
rect 1087 2750 1091 2754
rect 1223 2750 1227 2754
rect 1255 2750 1259 2754
rect 1399 2750 1403 2754
rect 1423 2750 1427 2754
rect 1575 2750 1579 2754
rect 1599 2750 1603 2754
rect 1751 2750 1755 2754
rect 1903 2750 1907 2754
rect 2007 2750 2011 2754
rect 2047 2694 2051 2698
rect 2071 2694 2075 2698
rect 2095 2694 2099 2698
rect 2199 2694 2203 2698
rect 2263 2694 2267 2698
rect 2343 2694 2347 2698
rect 2439 2694 2443 2698
rect 2479 2694 2483 2698
rect 2607 2694 2611 2698
rect 2615 2694 2619 2698
rect 2727 2694 2731 2698
rect 2783 2694 2787 2698
rect 2839 2694 2843 2698
rect 2943 2694 2947 2698
rect 3047 2694 3051 2698
rect 3095 2694 3099 2698
rect 3143 2694 3147 2698
rect 3239 2694 3243 2698
rect 3343 2694 3347 2698
rect 3383 2694 3387 2698
rect 3447 2694 3451 2698
rect 3535 2694 3539 2698
rect 3551 2694 3555 2698
rect 3647 2694 3651 2698
rect 3743 2694 3747 2698
rect 3839 2694 3843 2698
rect 3943 2694 3947 2698
rect 111 2674 115 2678
rect 135 2674 139 2678
rect 167 2674 171 2678
rect 255 2674 259 2678
rect 359 2674 363 2678
rect 407 2674 411 2678
rect 559 2674 563 2678
rect 575 2674 579 2678
rect 743 2674 747 2678
rect 759 2674 763 2678
rect 919 2674 923 2678
rect 951 2674 955 2678
rect 1087 2674 1091 2678
rect 1143 2674 1147 2678
rect 1255 2674 1259 2678
rect 1327 2674 1331 2678
rect 1423 2674 1427 2678
rect 1511 2674 1515 2678
rect 1599 2674 1603 2678
rect 1703 2674 1707 2678
rect 2007 2674 2011 2678
rect 2047 2610 2051 2614
rect 2095 2610 2099 2614
rect 2215 2610 2219 2614
rect 2263 2610 2267 2614
rect 2367 2610 2371 2614
rect 2439 2610 2443 2614
rect 2519 2610 2523 2614
rect 2615 2610 2619 2614
rect 2671 2610 2675 2614
rect 2783 2610 2787 2614
rect 2815 2610 2819 2614
rect 2943 2610 2947 2614
rect 2951 2610 2955 2614
rect 3087 2610 3091 2614
rect 3095 2610 3099 2614
rect 3223 2610 3227 2614
rect 3239 2610 3243 2614
rect 3367 2610 3371 2614
rect 3383 2610 3387 2614
rect 3535 2610 3539 2614
rect 3943 2610 3947 2614
rect 111 2582 115 2586
rect 167 2582 171 2586
rect 359 2582 363 2586
rect 559 2582 563 2586
rect 575 2582 579 2586
rect 687 2582 691 2586
rect 759 2582 763 2586
rect 807 2582 811 2586
rect 935 2582 939 2586
rect 951 2582 955 2586
rect 1071 2582 1075 2586
rect 1143 2582 1147 2586
rect 1207 2582 1211 2586
rect 1327 2582 1331 2586
rect 1351 2582 1355 2586
rect 1495 2582 1499 2586
rect 1511 2582 1515 2586
rect 1647 2582 1651 2586
rect 1703 2582 1707 2586
rect 1799 2582 1803 2586
rect 2007 2582 2011 2586
rect 2047 2530 2051 2534
rect 2095 2530 2099 2534
rect 2215 2530 2219 2534
rect 2343 2530 2347 2534
rect 2367 2530 2371 2534
rect 2471 2530 2475 2534
rect 2519 2530 2523 2534
rect 2599 2530 2603 2534
rect 2671 2530 2675 2534
rect 2719 2530 2723 2534
rect 2815 2530 2819 2534
rect 2839 2530 2843 2534
rect 2951 2530 2955 2534
rect 2967 2530 2971 2534
rect 3087 2530 3091 2534
rect 3095 2530 3099 2534
rect 3223 2530 3227 2534
rect 3367 2530 3371 2534
rect 3943 2530 3947 2534
rect 111 2502 115 2506
rect 503 2502 507 2506
rect 575 2502 579 2506
rect 607 2502 611 2506
rect 687 2502 691 2506
rect 719 2502 723 2506
rect 807 2502 811 2506
rect 847 2502 851 2506
rect 935 2502 939 2506
rect 983 2502 987 2506
rect 1071 2502 1075 2506
rect 1127 2502 1131 2506
rect 1207 2502 1211 2506
rect 1279 2502 1283 2506
rect 1351 2502 1355 2506
rect 1431 2502 1435 2506
rect 1495 2502 1499 2506
rect 1583 2502 1587 2506
rect 1647 2502 1651 2506
rect 1743 2502 1747 2506
rect 1799 2502 1803 2506
rect 1903 2502 1907 2506
rect 2007 2502 2011 2506
rect 2047 2442 2051 2446
rect 2071 2442 2075 2446
rect 2095 2442 2099 2446
rect 2191 2442 2195 2446
rect 2215 2442 2219 2446
rect 2319 2442 2323 2446
rect 2343 2442 2347 2446
rect 2439 2442 2443 2446
rect 2471 2442 2475 2446
rect 2559 2442 2563 2446
rect 2599 2442 2603 2446
rect 2679 2442 2683 2446
rect 2719 2442 2723 2446
rect 2791 2442 2795 2446
rect 2839 2442 2843 2446
rect 2911 2442 2915 2446
rect 2967 2442 2971 2446
rect 3031 2442 3035 2446
rect 3095 2442 3099 2446
rect 3151 2442 3155 2446
rect 3223 2442 3227 2446
rect 3943 2442 3947 2446
rect 111 2410 115 2414
rect 503 2410 507 2414
rect 535 2410 539 2414
rect 607 2410 611 2414
rect 671 2410 675 2414
rect 719 2410 723 2414
rect 815 2410 819 2414
rect 847 2410 851 2414
rect 959 2410 963 2414
rect 983 2410 987 2414
rect 1103 2410 1107 2414
rect 1127 2410 1131 2414
rect 1247 2410 1251 2414
rect 1279 2410 1283 2414
rect 1391 2410 1395 2414
rect 1431 2410 1435 2414
rect 1527 2410 1531 2414
rect 1583 2410 1587 2414
rect 1655 2410 1659 2414
rect 1743 2410 1747 2414
rect 1791 2410 1795 2414
rect 1903 2410 1907 2414
rect 2007 2410 2011 2414
rect 2047 2362 2051 2366
rect 2071 2362 2075 2366
rect 2167 2362 2171 2366
rect 2191 2362 2195 2366
rect 2319 2362 2323 2366
rect 2359 2362 2363 2366
rect 2439 2362 2443 2366
rect 2535 2362 2539 2366
rect 2559 2362 2563 2366
rect 2679 2362 2683 2366
rect 2703 2362 2707 2366
rect 2791 2362 2795 2366
rect 2871 2362 2875 2366
rect 2911 2362 2915 2366
rect 3031 2362 3035 2366
rect 3151 2362 3155 2366
rect 3199 2362 3203 2366
rect 3943 2362 3947 2366
rect 111 2330 115 2334
rect 535 2330 539 2334
rect 647 2330 651 2334
rect 671 2330 675 2334
rect 767 2330 771 2334
rect 815 2330 819 2334
rect 895 2330 899 2334
rect 959 2330 963 2334
rect 1031 2330 1035 2334
rect 1103 2330 1107 2334
rect 1167 2330 1171 2334
rect 1247 2330 1251 2334
rect 1295 2330 1299 2334
rect 1391 2330 1395 2334
rect 1423 2330 1427 2334
rect 1527 2330 1531 2334
rect 1551 2330 1555 2334
rect 1655 2330 1659 2334
rect 1671 2330 1675 2334
rect 1791 2330 1795 2334
rect 1799 2330 1803 2334
rect 1903 2330 1907 2334
rect 2007 2330 2011 2334
rect 2047 2286 2051 2290
rect 2071 2286 2075 2290
rect 2167 2286 2171 2290
rect 2287 2286 2291 2290
rect 2359 2286 2363 2290
rect 2423 2286 2427 2290
rect 2535 2286 2539 2290
rect 2559 2286 2563 2290
rect 2703 2286 2707 2290
rect 2839 2286 2843 2290
rect 2871 2286 2875 2290
rect 2983 2286 2987 2290
rect 3031 2286 3035 2290
rect 3127 2286 3131 2290
rect 3199 2286 3203 2290
rect 3271 2286 3275 2290
rect 3943 2286 3947 2290
rect 111 2250 115 2254
rect 415 2250 419 2254
rect 535 2250 539 2254
rect 647 2250 651 2254
rect 671 2250 675 2254
rect 767 2250 771 2254
rect 823 2250 827 2254
rect 895 2250 899 2254
rect 991 2250 995 2254
rect 1031 2250 1035 2254
rect 1167 2250 1171 2254
rect 1175 2250 1179 2254
rect 1295 2250 1299 2254
rect 1367 2250 1371 2254
rect 1423 2250 1427 2254
rect 1551 2250 1555 2254
rect 1567 2250 1571 2254
rect 1671 2250 1675 2254
rect 1767 2250 1771 2254
rect 1799 2250 1803 2254
rect 1903 2250 1907 2254
rect 2007 2250 2011 2254
rect 2047 2210 2051 2214
rect 2071 2210 2075 2214
rect 2167 2210 2171 2214
rect 2287 2210 2291 2214
rect 2295 2210 2299 2214
rect 2423 2210 2427 2214
rect 2503 2210 2507 2214
rect 2559 2210 2563 2214
rect 2687 2210 2691 2214
rect 2703 2210 2707 2214
rect 2839 2210 2843 2214
rect 2863 2210 2867 2214
rect 2983 2210 2987 2214
rect 3023 2210 3027 2214
rect 3127 2210 3131 2214
rect 3175 2210 3179 2214
rect 3271 2210 3275 2214
rect 3319 2210 3323 2214
rect 3471 2210 3475 2214
rect 3943 2210 3947 2214
rect 111 2166 115 2170
rect 135 2166 139 2170
rect 247 2166 251 2170
rect 391 2166 395 2170
rect 415 2166 419 2170
rect 535 2166 539 2170
rect 551 2166 555 2170
rect 671 2166 675 2170
rect 711 2166 715 2170
rect 823 2166 827 2170
rect 871 2166 875 2170
rect 991 2166 995 2170
rect 1031 2166 1035 2170
rect 1175 2166 1179 2170
rect 1191 2166 1195 2170
rect 1351 2166 1355 2170
rect 1367 2166 1371 2170
rect 1511 2166 1515 2170
rect 1567 2166 1571 2170
rect 1679 2166 1683 2170
rect 1767 2166 1771 2170
rect 2007 2166 2011 2170
rect 2047 2110 2051 2114
rect 2071 2110 2075 2114
rect 2295 2110 2299 2114
rect 2399 2110 2403 2114
rect 2495 2110 2499 2114
rect 2503 2110 2507 2114
rect 2591 2110 2595 2114
rect 2687 2110 2691 2114
rect 2783 2110 2787 2114
rect 2863 2110 2867 2114
rect 2879 2110 2883 2114
rect 2975 2110 2979 2114
rect 3023 2110 3027 2114
rect 3071 2110 3075 2114
rect 3167 2110 3171 2114
rect 3175 2110 3179 2114
rect 3263 2110 3267 2114
rect 3319 2110 3323 2114
rect 3359 2110 3363 2114
rect 3455 2110 3459 2114
rect 3471 2110 3475 2114
rect 3551 2110 3555 2114
rect 3647 2110 3651 2114
rect 3743 2110 3747 2114
rect 3839 2110 3843 2114
rect 3943 2110 3947 2114
rect 111 2082 115 2086
rect 135 2082 139 2086
rect 247 2082 251 2086
rect 391 2082 395 2086
rect 399 2082 403 2086
rect 551 2082 555 2086
rect 703 2082 707 2086
rect 711 2082 715 2086
rect 847 2082 851 2086
rect 871 2082 875 2086
rect 991 2082 995 2086
rect 1031 2082 1035 2086
rect 1127 2082 1131 2086
rect 1191 2082 1195 2086
rect 1255 2082 1259 2086
rect 1351 2082 1355 2086
rect 1383 2082 1387 2086
rect 1511 2082 1515 2086
rect 1519 2082 1523 2086
rect 1679 2082 1683 2086
rect 2007 2082 2011 2086
rect 2047 2034 2051 2038
rect 2191 2034 2195 2038
rect 2399 2034 2403 2038
rect 2495 2034 2499 2038
rect 2591 2034 2595 2038
rect 2647 2034 2651 2038
rect 2687 2034 2691 2038
rect 2783 2034 2787 2038
rect 2879 2034 2883 2038
rect 2919 2034 2923 2038
rect 2975 2034 2979 2038
rect 3071 2034 3075 2038
rect 3167 2034 3171 2038
rect 3215 2034 3219 2038
rect 3263 2034 3267 2038
rect 3359 2034 3363 2038
rect 3455 2034 3459 2038
rect 3527 2034 3531 2038
rect 3551 2034 3555 2038
rect 3647 2034 3651 2038
rect 3743 2034 3747 2038
rect 3839 2034 3843 2038
rect 3943 2034 3947 2038
rect 111 1990 115 1994
rect 135 1990 139 1994
rect 231 1990 235 1994
rect 247 1990 251 1994
rect 391 1990 395 1994
rect 399 1990 403 1994
rect 551 1990 555 1994
rect 567 1990 571 1994
rect 703 1990 707 1994
rect 751 1990 755 1994
rect 847 1990 851 1994
rect 943 1990 947 1994
rect 991 1990 995 1994
rect 1127 1990 1131 1994
rect 1135 1990 1139 1994
rect 1255 1990 1259 1994
rect 1335 1990 1339 1994
rect 1383 1990 1387 1994
rect 1519 1990 1523 1994
rect 1543 1990 1547 1994
rect 2007 1990 2011 1994
rect 2047 1946 2051 1950
rect 2071 1946 2075 1950
rect 2191 1946 2195 1950
rect 2239 1946 2243 1950
rect 2399 1946 2403 1950
rect 2447 1946 2451 1950
rect 2647 1946 2651 1950
rect 2671 1946 2675 1950
rect 2895 1946 2899 1950
rect 2919 1946 2923 1950
rect 3127 1946 3131 1950
rect 3215 1946 3219 1950
rect 3359 1946 3363 1950
rect 3527 1946 3531 1950
rect 3591 1946 3595 1950
rect 3831 1946 3835 1950
rect 3839 1946 3843 1950
rect 3943 1946 3947 1950
rect 111 1914 115 1918
rect 231 1914 235 1918
rect 391 1914 395 1918
rect 511 1914 515 1918
rect 567 1914 571 1918
rect 623 1914 627 1918
rect 743 1914 747 1918
rect 751 1914 755 1918
rect 863 1914 867 1918
rect 943 1914 947 1918
rect 983 1914 987 1918
rect 1103 1914 1107 1918
rect 1135 1914 1139 1918
rect 1223 1914 1227 1918
rect 1335 1914 1339 1918
rect 1455 1914 1459 1918
rect 1543 1914 1547 1918
rect 1575 1914 1579 1918
rect 1695 1914 1699 1918
rect 2007 1914 2011 1918
rect 2047 1870 2051 1874
rect 2071 1870 2075 1874
rect 2199 1870 2203 1874
rect 2239 1870 2243 1874
rect 2367 1870 2371 1874
rect 2447 1870 2451 1874
rect 2543 1870 2547 1874
rect 2671 1870 2675 1874
rect 2719 1870 2723 1874
rect 2887 1870 2891 1874
rect 2895 1870 2899 1874
rect 3039 1870 3043 1874
rect 3127 1870 3131 1874
rect 3183 1870 3187 1874
rect 3319 1870 3323 1874
rect 3359 1870 3363 1874
rect 3455 1870 3459 1874
rect 3583 1870 3587 1874
rect 3591 1870 3595 1874
rect 3711 1870 3715 1874
rect 3831 1870 3835 1874
rect 3839 1870 3843 1874
rect 3943 1870 3947 1874
rect 111 1830 115 1834
rect 511 1830 515 1834
rect 615 1830 619 1834
rect 623 1830 627 1834
rect 711 1830 715 1834
rect 743 1830 747 1834
rect 815 1830 819 1834
rect 863 1830 867 1834
rect 927 1830 931 1834
rect 983 1830 987 1834
rect 1039 1830 1043 1834
rect 1103 1830 1107 1834
rect 1159 1830 1163 1834
rect 1223 1830 1227 1834
rect 1279 1830 1283 1834
rect 1335 1830 1339 1834
rect 1399 1830 1403 1834
rect 1455 1830 1459 1834
rect 1519 1830 1523 1834
rect 1575 1830 1579 1834
rect 1639 1830 1643 1834
rect 1695 1830 1699 1834
rect 2007 1830 2011 1834
rect 2047 1790 2051 1794
rect 2071 1790 2075 1794
rect 2183 1790 2187 1794
rect 2199 1790 2203 1794
rect 2327 1790 2331 1794
rect 2367 1790 2371 1794
rect 2487 1790 2491 1794
rect 2543 1790 2547 1794
rect 2655 1790 2659 1794
rect 2719 1790 2723 1794
rect 2831 1790 2835 1794
rect 2887 1790 2891 1794
rect 3023 1790 3027 1794
rect 3039 1790 3043 1794
rect 3183 1790 3187 1794
rect 3223 1790 3227 1794
rect 3319 1790 3323 1794
rect 3431 1790 3435 1794
rect 3455 1790 3459 1794
rect 3583 1790 3587 1794
rect 3647 1790 3651 1794
rect 3711 1790 3715 1794
rect 3839 1790 3843 1794
rect 3943 1790 3947 1794
rect 111 1754 115 1758
rect 367 1754 371 1758
rect 495 1754 499 1758
rect 615 1754 619 1758
rect 639 1754 643 1758
rect 711 1754 715 1758
rect 799 1754 803 1758
rect 815 1754 819 1758
rect 927 1754 931 1758
rect 967 1754 971 1758
rect 1039 1754 1043 1758
rect 1143 1754 1147 1758
rect 1159 1754 1163 1758
rect 1279 1754 1283 1758
rect 1327 1754 1331 1758
rect 1399 1754 1403 1758
rect 1511 1754 1515 1758
rect 1519 1754 1523 1758
rect 1639 1754 1643 1758
rect 1703 1754 1707 1758
rect 2007 1754 2011 1758
rect 2047 1706 2051 1710
rect 2071 1706 2075 1710
rect 2183 1706 2187 1710
rect 2223 1706 2227 1710
rect 2327 1706 2331 1710
rect 2439 1706 2443 1710
rect 2487 1706 2491 1710
rect 2559 1706 2563 1710
rect 2655 1706 2659 1710
rect 2687 1706 2691 1710
rect 2823 1706 2827 1710
rect 2831 1706 2835 1710
rect 2967 1706 2971 1710
rect 3023 1706 3027 1710
rect 3127 1706 3131 1710
rect 3223 1706 3227 1710
rect 3303 1706 3307 1710
rect 3431 1706 3435 1710
rect 3487 1706 3491 1710
rect 3647 1706 3651 1710
rect 3671 1706 3675 1710
rect 3839 1706 3843 1710
rect 3943 1706 3947 1710
rect 111 1674 115 1678
rect 135 1674 139 1678
rect 247 1674 251 1678
rect 367 1674 371 1678
rect 399 1674 403 1678
rect 495 1674 499 1678
rect 567 1674 571 1678
rect 639 1674 643 1678
rect 743 1674 747 1678
rect 799 1674 803 1678
rect 935 1674 939 1678
rect 967 1674 971 1678
rect 1135 1674 1139 1678
rect 1143 1674 1147 1678
rect 1327 1674 1331 1678
rect 1343 1674 1347 1678
rect 1511 1674 1515 1678
rect 1551 1674 1555 1678
rect 1703 1674 1707 1678
rect 1767 1674 1771 1678
rect 2007 1674 2011 1678
rect 2047 1626 2051 1630
rect 2223 1626 2227 1630
rect 2327 1626 2331 1630
rect 2391 1626 2395 1630
rect 2439 1626 2443 1630
rect 2503 1626 2507 1630
rect 2559 1626 2563 1630
rect 2615 1626 2619 1630
rect 2687 1626 2691 1630
rect 2735 1626 2739 1630
rect 2823 1626 2827 1630
rect 2855 1626 2859 1630
rect 2967 1626 2971 1630
rect 2975 1626 2979 1630
rect 3095 1626 3099 1630
rect 3127 1626 3131 1630
rect 3215 1626 3219 1630
rect 3303 1626 3307 1630
rect 3335 1626 3339 1630
rect 3455 1626 3459 1630
rect 3487 1626 3491 1630
rect 3671 1626 3675 1630
rect 3839 1626 3843 1630
rect 3943 1626 3947 1630
rect 111 1594 115 1598
rect 135 1594 139 1598
rect 247 1594 251 1598
rect 255 1594 259 1598
rect 399 1594 403 1598
rect 423 1594 427 1598
rect 567 1594 571 1598
rect 615 1594 619 1598
rect 743 1594 747 1598
rect 831 1594 835 1598
rect 935 1594 939 1598
rect 1063 1594 1067 1598
rect 1135 1594 1139 1598
rect 1311 1594 1315 1598
rect 1343 1594 1347 1598
rect 1551 1594 1555 1598
rect 1567 1594 1571 1598
rect 1767 1594 1771 1598
rect 1831 1594 1835 1598
rect 2007 1594 2011 1598
rect 2047 1550 2051 1554
rect 2391 1550 2395 1554
rect 2503 1550 2507 1554
rect 2543 1550 2547 1554
rect 2615 1550 2619 1554
rect 2671 1550 2675 1554
rect 2735 1550 2739 1554
rect 2799 1550 2803 1554
rect 2855 1550 2859 1554
rect 2935 1550 2939 1554
rect 2975 1550 2979 1554
rect 3071 1550 3075 1554
rect 3095 1550 3099 1554
rect 3207 1550 3211 1554
rect 3215 1550 3219 1554
rect 3335 1550 3339 1554
rect 3455 1550 3459 1554
rect 3463 1550 3467 1554
rect 3591 1550 3595 1554
rect 3727 1550 3731 1554
rect 3839 1550 3843 1554
rect 3943 1550 3947 1554
rect 111 1514 115 1518
rect 135 1514 139 1518
rect 239 1514 243 1518
rect 255 1514 259 1518
rect 407 1514 411 1518
rect 423 1514 427 1518
rect 583 1514 587 1518
rect 615 1514 619 1518
rect 775 1514 779 1518
rect 831 1514 835 1518
rect 967 1514 971 1518
rect 1063 1514 1067 1518
rect 1159 1514 1163 1518
rect 1311 1514 1315 1518
rect 1351 1514 1355 1518
rect 1543 1514 1547 1518
rect 1567 1514 1571 1518
rect 1735 1514 1739 1518
rect 1831 1514 1835 1518
rect 1903 1514 1907 1518
rect 2007 1514 2011 1518
rect 2047 1462 2051 1466
rect 2519 1462 2523 1466
rect 2543 1462 2547 1466
rect 2631 1462 2635 1466
rect 2671 1462 2675 1466
rect 2759 1462 2763 1466
rect 2799 1462 2803 1466
rect 2895 1462 2899 1466
rect 2935 1462 2939 1466
rect 3031 1462 3035 1466
rect 3071 1462 3075 1466
rect 3175 1462 3179 1466
rect 3207 1462 3211 1466
rect 3311 1462 3315 1466
rect 3335 1462 3339 1466
rect 3447 1462 3451 1466
rect 3463 1462 3467 1466
rect 3583 1462 3587 1466
rect 3591 1462 3595 1466
rect 3719 1462 3723 1466
rect 3727 1462 3731 1466
rect 3839 1462 3843 1466
rect 3943 1462 3947 1466
rect 111 1430 115 1434
rect 239 1430 243 1434
rect 407 1430 411 1434
rect 463 1430 467 1434
rect 583 1430 587 1434
rect 711 1430 715 1434
rect 775 1430 779 1434
rect 855 1430 859 1434
rect 967 1430 971 1434
rect 1007 1430 1011 1434
rect 1159 1430 1163 1434
rect 1167 1430 1171 1434
rect 1335 1430 1339 1434
rect 1351 1430 1355 1434
rect 1511 1430 1515 1434
rect 1543 1430 1547 1434
rect 1687 1430 1691 1434
rect 1735 1430 1739 1434
rect 1871 1430 1875 1434
rect 1903 1430 1907 1434
rect 2007 1430 2011 1434
rect 2047 1386 2051 1390
rect 2399 1386 2403 1390
rect 2519 1386 2523 1390
rect 2535 1386 2539 1390
rect 2631 1386 2635 1390
rect 2679 1386 2683 1390
rect 2759 1386 2763 1390
rect 2823 1386 2827 1390
rect 2895 1386 2899 1390
rect 2967 1386 2971 1390
rect 3031 1386 3035 1390
rect 3111 1386 3115 1390
rect 3175 1386 3179 1390
rect 3255 1386 3259 1390
rect 3311 1386 3315 1390
rect 3407 1386 3411 1390
rect 3447 1386 3451 1390
rect 3559 1386 3563 1390
rect 3583 1386 3587 1390
rect 3711 1386 3715 1390
rect 3719 1386 3723 1390
rect 3839 1386 3843 1390
rect 3943 1386 3947 1390
rect 111 1354 115 1358
rect 463 1354 467 1358
rect 583 1354 587 1358
rect 655 1354 659 1358
rect 711 1354 715 1358
rect 767 1354 771 1358
rect 855 1354 859 1358
rect 887 1354 891 1358
rect 1007 1354 1011 1358
rect 1015 1354 1019 1358
rect 1143 1354 1147 1358
rect 1167 1354 1171 1358
rect 1279 1354 1283 1358
rect 1335 1354 1339 1358
rect 1415 1354 1419 1358
rect 1511 1354 1515 1358
rect 1559 1354 1563 1358
rect 1687 1354 1691 1358
rect 1703 1354 1707 1358
rect 1847 1354 1851 1358
rect 1871 1354 1875 1358
rect 2007 1354 2011 1358
rect 2047 1306 2051 1310
rect 2247 1306 2251 1310
rect 2375 1306 2379 1310
rect 2399 1306 2403 1310
rect 2511 1306 2515 1310
rect 2535 1306 2539 1310
rect 2647 1306 2651 1310
rect 2679 1306 2683 1310
rect 2791 1306 2795 1310
rect 2823 1306 2827 1310
rect 2943 1306 2947 1310
rect 2967 1306 2971 1310
rect 3111 1306 3115 1310
rect 3255 1306 3259 1310
rect 3287 1306 3291 1310
rect 3407 1306 3411 1310
rect 3471 1306 3475 1310
rect 3559 1306 3563 1310
rect 3663 1306 3667 1310
rect 3711 1306 3715 1310
rect 3839 1306 3843 1310
rect 3943 1306 3947 1310
rect 111 1274 115 1278
rect 439 1274 443 1278
rect 551 1274 555 1278
rect 655 1274 659 1278
rect 671 1274 675 1278
rect 767 1274 771 1278
rect 799 1274 803 1278
rect 887 1274 891 1278
rect 935 1274 939 1278
rect 1015 1274 1019 1278
rect 1079 1274 1083 1278
rect 1143 1274 1147 1278
rect 1231 1274 1235 1278
rect 1279 1274 1283 1278
rect 1391 1274 1395 1278
rect 1415 1274 1419 1278
rect 1551 1274 1555 1278
rect 1559 1274 1563 1278
rect 1703 1274 1707 1278
rect 1719 1274 1723 1278
rect 1847 1274 1851 1278
rect 2007 1274 2011 1278
rect 2047 1226 2051 1230
rect 2071 1226 2075 1230
rect 2183 1226 2187 1230
rect 2247 1226 2251 1230
rect 2303 1226 2307 1230
rect 2375 1226 2379 1230
rect 2431 1226 2435 1230
rect 2511 1226 2515 1230
rect 2559 1226 2563 1230
rect 2647 1226 2651 1230
rect 2711 1226 2715 1230
rect 2791 1226 2795 1230
rect 2887 1226 2891 1230
rect 2943 1226 2947 1230
rect 3087 1226 3091 1230
rect 3111 1226 3115 1230
rect 3287 1226 3291 1230
rect 3311 1226 3315 1230
rect 3471 1226 3475 1230
rect 3543 1226 3547 1230
rect 3663 1226 3667 1230
rect 3783 1226 3787 1230
rect 3839 1226 3843 1230
rect 3943 1226 3947 1230
rect 111 1198 115 1202
rect 167 1198 171 1202
rect 303 1198 307 1202
rect 439 1198 443 1202
rect 463 1198 467 1202
rect 551 1198 555 1202
rect 631 1198 635 1202
rect 671 1198 675 1202
rect 799 1198 803 1202
rect 807 1198 811 1202
rect 935 1198 939 1202
rect 983 1198 987 1202
rect 1079 1198 1083 1202
rect 1159 1198 1163 1202
rect 1231 1198 1235 1202
rect 1335 1198 1339 1202
rect 1391 1198 1395 1202
rect 1511 1198 1515 1202
rect 1551 1198 1555 1202
rect 1695 1198 1699 1202
rect 1719 1198 1723 1202
rect 2007 1198 2011 1202
rect 2047 1146 2051 1150
rect 2071 1146 2075 1150
rect 2183 1146 2187 1150
rect 2199 1146 2203 1150
rect 2303 1146 2307 1150
rect 2351 1146 2355 1150
rect 2431 1146 2435 1150
rect 2511 1146 2515 1150
rect 2559 1146 2563 1150
rect 2679 1146 2683 1150
rect 2711 1146 2715 1150
rect 2871 1146 2875 1150
rect 2887 1146 2891 1150
rect 3087 1146 3091 1150
rect 3311 1146 3315 1150
rect 3319 1146 3323 1150
rect 3543 1146 3547 1150
rect 3559 1146 3563 1150
rect 3783 1146 3787 1150
rect 3807 1146 3811 1150
rect 3943 1146 3947 1150
rect 111 1118 115 1122
rect 135 1118 139 1122
rect 167 1118 171 1122
rect 239 1118 243 1122
rect 303 1118 307 1122
rect 375 1118 379 1122
rect 463 1118 467 1122
rect 527 1118 531 1122
rect 631 1118 635 1122
rect 695 1118 699 1122
rect 807 1118 811 1122
rect 863 1118 867 1122
rect 983 1118 987 1122
rect 1039 1118 1043 1122
rect 1159 1118 1163 1122
rect 1215 1118 1219 1122
rect 1335 1118 1339 1122
rect 1391 1118 1395 1122
rect 1511 1118 1515 1122
rect 1567 1118 1571 1122
rect 1695 1118 1699 1122
rect 1743 1118 1747 1122
rect 1903 1118 1907 1122
rect 2007 1118 2011 1122
rect 2047 1058 2051 1062
rect 2071 1058 2075 1062
rect 2199 1058 2203 1062
rect 2263 1058 2267 1062
rect 2351 1058 2355 1062
rect 2487 1058 2491 1062
rect 2511 1058 2515 1062
rect 2679 1058 2683 1062
rect 2703 1058 2707 1062
rect 2871 1058 2875 1062
rect 2919 1058 2923 1062
rect 3087 1058 3091 1062
rect 3119 1058 3123 1062
rect 3311 1058 3315 1062
rect 3319 1058 3323 1062
rect 3495 1058 3499 1062
rect 3559 1058 3563 1062
rect 3679 1058 3683 1062
rect 3807 1058 3811 1062
rect 3839 1058 3843 1062
rect 3943 1058 3947 1062
rect 111 1042 115 1046
rect 135 1042 139 1046
rect 239 1042 243 1046
rect 287 1042 291 1046
rect 375 1042 379 1046
rect 471 1042 475 1046
rect 527 1042 531 1046
rect 655 1042 659 1046
rect 695 1042 699 1046
rect 839 1042 843 1046
rect 863 1042 867 1046
rect 1015 1042 1019 1046
rect 1039 1042 1043 1046
rect 1199 1042 1203 1046
rect 1215 1042 1219 1046
rect 1383 1042 1387 1046
rect 1391 1042 1395 1046
rect 1567 1042 1571 1046
rect 1743 1042 1747 1046
rect 1903 1042 1907 1046
rect 2007 1042 2011 1046
rect 2047 978 2051 982
rect 2071 978 2075 982
rect 2263 978 2267 982
rect 2303 978 2307 982
rect 2455 978 2459 982
rect 2487 978 2491 982
rect 2615 978 2619 982
rect 2703 978 2707 982
rect 2783 978 2787 982
rect 2919 978 2923 982
rect 2951 978 2955 982
rect 3111 978 3115 982
rect 3119 978 3123 982
rect 3263 978 3267 982
rect 3311 978 3315 982
rect 3415 978 3419 982
rect 3495 978 3499 982
rect 3559 978 3563 982
rect 3679 978 3683 982
rect 3711 978 3715 982
rect 3839 978 3843 982
rect 3943 978 3947 982
rect 111 962 115 966
rect 135 962 139 966
rect 287 962 291 966
rect 295 962 299 966
rect 471 962 475 966
rect 639 962 643 966
rect 655 962 659 966
rect 799 962 803 966
rect 839 962 843 966
rect 951 962 955 966
rect 1015 962 1019 966
rect 1087 962 1091 966
rect 1199 962 1203 966
rect 1223 962 1227 966
rect 1359 962 1363 966
rect 1383 962 1387 966
rect 1495 962 1499 966
rect 1567 962 1571 966
rect 2007 962 2011 966
rect 2047 898 2051 902
rect 2303 898 2307 902
rect 2455 898 2459 902
rect 2559 898 2563 902
rect 2615 898 2619 902
rect 2679 898 2683 902
rect 2783 898 2787 902
rect 2807 898 2811 902
rect 2943 898 2947 902
rect 2951 898 2955 902
rect 3079 898 3083 902
rect 3111 898 3115 902
rect 3207 898 3211 902
rect 3263 898 3267 902
rect 3335 898 3339 902
rect 3415 898 3419 902
rect 3463 898 3467 902
rect 3559 898 3563 902
rect 3591 898 3595 902
rect 3711 898 3715 902
rect 3727 898 3731 902
rect 3839 898 3843 902
rect 3943 898 3947 902
rect 111 886 115 890
rect 135 886 139 890
rect 159 886 163 890
rect 295 886 299 890
rect 319 886 323 890
rect 471 886 475 890
rect 615 886 619 890
rect 639 886 643 890
rect 751 886 755 890
rect 799 886 803 890
rect 879 886 883 890
rect 951 886 955 890
rect 999 886 1003 890
rect 1087 886 1091 890
rect 1111 886 1115 890
rect 1223 886 1227 890
rect 1231 886 1235 890
rect 1351 886 1355 890
rect 1359 886 1363 890
rect 1495 886 1499 890
rect 2007 886 2011 890
rect 2047 818 2051 822
rect 2335 818 2339 822
rect 2471 818 2475 822
rect 2559 818 2563 822
rect 2615 818 2619 822
rect 2679 818 2683 822
rect 2767 818 2771 822
rect 2807 818 2811 822
rect 2919 818 2923 822
rect 2943 818 2947 822
rect 3079 818 3083 822
rect 3207 818 3211 822
rect 3239 818 3243 822
rect 3335 818 3339 822
rect 3391 818 3395 822
rect 3463 818 3467 822
rect 3543 818 3547 822
rect 3591 818 3595 822
rect 3703 818 3707 822
rect 3727 818 3731 822
rect 3839 818 3843 822
rect 3943 818 3947 822
rect 111 810 115 814
rect 159 810 163 814
rect 223 810 227 814
rect 319 810 323 814
rect 383 810 387 814
rect 471 810 475 814
rect 535 810 539 814
rect 615 810 619 814
rect 679 810 683 814
rect 751 810 755 814
rect 815 810 819 814
rect 879 810 883 814
rect 951 810 955 814
rect 999 810 1003 814
rect 1079 810 1083 814
rect 1111 810 1115 814
rect 1199 810 1203 814
rect 1231 810 1235 814
rect 1327 810 1331 814
rect 1351 810 1355 814
rect 1455 810 1459 814
rect 2007 810 2011 814
rect 2047 738 2051 742
rect 2071 738 2075 742
rect 2183 738 2187 742
rect 2335 738 2339 742
rect 2471 738 2475 742
rect 2487 738 2491 742
rect 2615 738 2619 742
rect 2639 738 2643 742
rect 2767 738 2771 742
rect 2807 738 2811 742
rect 2919 738 2923 742
rect 2983 738 2987 742
rect 3079 738 3083 742
rect 3167 738 3171 742
rect 3239 738 3243 742
rect 3367 738 3371 742
rect 3391 738 3395 742
rect 3543 738 3547 742
rect 3575 738 3579 742
rect 3703 738 3707 742
rect 3783 738 3787 742
rect 3839 738 3843 742
rect 3943 738 3947 742
rect 111 730 115 734
rect 223 730 227 734
rect 311 730 315 734
rect 383 730 387 734
rect 471 730 475 734
rect 535 730 539 734
rect 639 730 643 734
rect 679 730 683 734
rect 807 730 811 734
rect 815 730 819 734
rect 951 730 955 734
rect 975 730 979 734
rect 1079 730 1083 734
rect 1135 730 1139 734
rect 1199 730 1203 734
rect 1295 730 1299 734
rect 1327 730 1331 734
rect 1455 730 1459 734
rect 1607 730 1611 734
rect 1767 730 1771 734
rect 1903 730 1907 734
rect 2007 730 2011 734
rect 111 654 115 658
rect 295 654 299 658
rect 311 654 315 658
rect 447 654 451 658
rect 471 654 475 658
rect 615 654 619 658
rect 639 654 643 658
rect 783 654 787 658
rect 807 654 811 658
rect 951 654 955 658
rect 975 654 979 658
rect 1111 654 1115 658
rect 1135 654 1139 658
rect 1263 654 1267 658
rect 1295 654 1299 658
rect 1399 654 1403 658
rect 1455 654 1459 658
rect 1535 654 1539 658
rect 1607 654 1611 658
rect 1663 654 1667 658
rect 1767 654 1771 658
rect 1791 654 1795 658
rect 1903 654 1907 658
rect 2007 654 2011 658
rect 2047 650 2051 654
rect 2071 650 2075 654
rect 2183 650 2187 654
rect 2239 650 2243 654
rect 2335 650 2339 654
rect 2423 650 2427 654
rect 2487 650 2491 654
rect 2623 650 2627 654
rect 2639 650 2643 654
rect 2807 650 2811 654
rect 2839 650 2843 654
rect 2983 650 2987 654
rect 3071 650 3075 654
rect 3167 650 3171 654
rect 3319 650 3323 654
rect 3367 650 3371 654
rect 3575 650 3579 654
rect 3783 650 3787 654
rect 3839 650 3843 654
rect 3943 650 3947 654
rect 111 574 115 578
rect 239 574 243 578
rect 295 574 299 578
rect 415 574 419 578
rect 447 574 451 578
rect 607 574 611 578
rect 615 574 619 578
rect 783 574 787 578
rect 799 574 803 578
rect 951 574 955 578
rect 991 574 995 578
rect 1111 574 1115 578
rect 1175 574 1179 578
rect 1263 574 1267 578
rect 1351 574 1355 578
rect 1399 574 1403 578
rect 1519 574 1523 578
rect 1535 574 1539 578
rect 1663 574 1667 578
rect 1687 574 1691 578
rect 1791 574 1795 578
rect 1863 574 1867 578
rect 1903 574 1907 578
rect 2007 574 2011 578
rect 2047 574 2051 578
rect 2071 574 2075 578
rect 2191 574 2195 578
rect 2239 574 2243 578
rect 2287 574 2291 578
rect 2383 574 2387 578
rect 2423 574 2427 578
rect 2479 574 2483 578
rect 2583 574 2587 578
rect 2623 574 2627 578
rect 2711 574 2715 578
rect 2839 574 2843 578
rect 2871 574 2875 578
rect 3071 574 3075 578
rect 3303 574 3307 578
rect 3319 574 3323 578
rect 3551 574 3555 578
rect 3575 574 3579 578
rect 3807 574 3811 578
rect 3839 574 3843 578
rect 3943 574 3947 578
rect 111 498 115 502
rect 135 498 139 502
rect 239 498 243 502
rect 287 498 291 502
rect 415 498 419 502
rect 463 498 467 502
rect 607 498 611 502
rect 639 498 643 502
rect 799 498 803 502
rect 807 498 811 502
rect 967 498 971 502
rect 991 498 995 502
rect 1119 498 1123 502
rect 1175 498 1179 502
rect 1271 498 1275 502
rect 1351 498 1355 502
rect 1415 498 1419 502
rect 1519 498 1523 502
rect 1567 498 1571 502
rect 1687 498 1691 502
rect 1863 498 1867 502
rect 2007 498 2011 502
rect 2047 498 2051 502
rect 2191 498 2195 502
rect 2287 498 2291 502
rect 2383 498 2387 502
rect 2431 498 2435 502
rect 2479 498 2483 502
rect 2527 498 2531 502
rect 2583 498 2587 502
rect 2623 498 2627 502
rect 2711 498 2715 502
rect 2727 498 2731 502
rect 2847 498 2851 502
rect 2871 498 2875 502
rect 2999 498 3003 502
rect 3071 498 3075 502
rect 3175 498 3179 502
rect 3303 498 3307 502
rect 3375 498 3379 502
rect 3551 498 3555 502
rect 3591 498 3595 502
rect 3807 498 3811 502
rect 3943 498 3947 502
rect 111 418 115 422
rect 135 418 139 422
rect 279 418 283 422
rect 287 418 291 422
rect 439 418 443 422
rect 463 418 467 422
rect 583 418 587 422
rect 639 418 643 422
rect 719 418 723 422
rect 807 418 811 422
rect 847 418 851 422
rect 967 418 971 422
rect 1087 418 1091 422
rect 1119 418 1123 422
rect 1207 418 1211 422
rect 1271 418 1275 422
rect 1327 418 1331 422
rect 1415 418 1419 422
rect 1567 418 1571 422
rect 2007 418 2011 422
rect 2047 422 2051 426
rect 2431 422 2435 426
rect 2527 422 2531 426
rect 2623 422 2627 426
rect 2719 422 2723 426
rect 2727 422 2731 426
rect 2815 422 2819 426
rect 2847 422 2851 426
rect 2927 422 2931 426
rect 2999 422 3003 426
rect 3063 422 3067 426
rect 3175 422 3179 426
rect 3223 422 3227 426
rect 3375 422 3379 426
rect 3399 422 3403 426
rect 3591 422 3595 426
rect 3783 422 3787 426
rect 3807 422 3811 426
rect 3943 422 3947 426
rect 111 342 115 346
rect 135 342 139 346
rect 143 342 147 346
rect 279 342 283 346
rect 319 342 323 346
rect 439 342 443 346
rect 479 342 483 346
rect 583 342 587 346
rect 631 342 635 346
rect 719 342 723 346
rect 775 342 779 346
rect 847 342 851 346
rect 903 342 907 346
rect 967 342 971 346
rect 1031 342 1035 346
rect 1087 342 1091 346
rect 1151 342 1155 346
rect 1207 342 1211 346
rect 1271 342 1275 346
rect 1327 342 1331 346
rect 1391 342 1395 346
rect 2007 342 2011 346
rect 2047 342 2051 346
rect 2191 342 2195 346
rect 2327 342 2331 346
rect 2431 342 2435 346
rect 2471 342 2475 346
rect 2527 342 2531 346
rect 2623 342 2627 346
rect 2719 342 2723 346
rect 2783 342 2787 346
rect 2815 342 2819 346
rect 2927 342 2931 346
rect 2951 342 2955 346
rect 3063 342 3067 346
rect 3119 342 3123 346
rect 3223 342 3227 346
rect 3295 342 3299 346
rect 3399 342 3403 346
rect 3471 342 3475 346
rect 3591 342 3595 346
rect 3655 342 3659 346
rect 3783 342 3787 346
rect 3839 342 3843 346
rect 3943 342 3947 346
rect 111 262 115 266
rect 143 262 147 266
rect 223 262 227 266
rect 319 262 323 266
rect 391 262 395 266
rect 479 262 483 266
rect 559 262 563 266
rect 631 262 635 266
rect 735 262 739 266
rect 775 262 779 266
rect 903 262 907 266
rect 1031 262 1035 266
rect 1063 262 1067 266
rect 1151 262 1155 266
rect 1215 262 1219 266
rect 1271 262 1275 266
rect 1359 262 1363 266
rect 1391 262 1395 266
rect 1511 262 1515 266
rect 1663 262 1667 266
rect 2007 262 2011 266
rect 2047 266 2051 270
rect 2071 266 2075 270
rect 2191 266 2195 270
rect 2215 266 2219 270
rect 2327 266 2331 270
rect 2399 266 2403 270
rect 2471 266 2475 270
rect 2591 266 2595 270
rect 2623 266 2627 270
rect 2783 266 2787 270
rect 2791 266 2795 270
rect 2951 266 2955 270
rect 2983 266 2987 270
rect 3119 266 3123 270
rect 3167 266 3171 270
rect 3295 266 3299 270
rect 3343 266 3347 270
rect 3471 266 3475 270
rect 3511 266 3515 270
rect 3655 266 3659 270
rect 3687 266 3691 270
rect 3839 266 3843 270
rect 3943 266 3947 270
rect 2047 166 2051 170
rect 2071 166 2075 170
rect 2191 166 2195 170
rect 2215 166 2219 170
rect 2343 166 2347 170
rect 2399 166 2403 170
rect 2495 166 2499 170
rect 2591 166 2595 170
rect 2647 166 2651 170
rect 2791 166 2795 170
rect 2799 166 2803 170
rect 2943 166 2947 170
rect 2983 166 2987 170
rect 3071 166 3075 170
rect 3167 166 3171 170
rect 3191 166 3195 170
rect 3311 166 3315 170
rect 3343 166 3347 170
rect 3423 166 3427 170
rect 3511 166 3515 170
rect 3527 166 3531 170
rect 3639 166 3643 170
rect 3687 166 3691 170
rect 3743 166 3747 170
rect 3839 166 3843 170
rect 3943 166 3947 170
rect 111 154 115 158
rect 151 154 155 158
rect 223 154 227 158
rect 247 154 251 158
rect 343 154 347 158
rect 391 154 395 158
rect 439 154 443 158
rect 535 154 539 158
rect 559 154 563 158
rect 631 154 635 158
rect 727 154 731 158
rect 735 154 739 158
rect 823 154 827 158
rect 903 154 907 158
rect 919 154 923 158
rect 1015 154 1019 158
rect 1063 154 1067 158
rect 1111 154 1115 158
rect 1207 154 1211 158
rect 1215 154 1219 158
rect 1303 154 1307 158
rect 1359 154 1363 158
rect 1407 154 1411 158
rect 1511 154 1515 158
rect 1615 154 1619 158
rect 1663 154 1667 158
rect 1711 154 1715 158
rect 1807 154 1811 158
rect 1903 154 1907 158
rect 2007 154 2011 158
rect 2047 90 2051 94
rect 2071 90 2075 94
rect 2191 90 2195 94
rect 2343 90 2347 94
rect 2495 90 2499 94
rect 2647 90 2651 94
rect 2799 90 2803 94
rect 2943 90 2947 94
rect 3071 90 3075 94
rect 3191 90 3195 94
rect 3311 90 3315 94
rect 3423 90 3427 94
rect 3527 90 3531 94
rect 3639 90 3643 94
rect 3743 90 3747 94
rect 3839 90 3843 94
rect 3943 90 3947 94
rect 111 78 115 82
rect 151 78 155 82
rect 247 78 251 82
rect 343 78 347 82
rect 439 78 443 82
rect 535 78 539 82
rect 631 78 635 82
rect 727 78 731 82
rect 823 78 827 82
rect 919 78 923 82
rect 1015 78 1019 82
rect 1111 78 1115 82
rect 1207 78 1211 82
rect 1303 78 1307 82
rect 1407 78 1411 82
rect 1511 78 1515 82
rect 1615 78 1619 82
rect 1711 78 1715 82
rect 1807 78 1811 82
rect 1903 78 1907 82
rect 2007 78 2011 82
<< m4 >>
rect 2018 4017 2019 4023
rect 2025 4022 3967 4023
rect 2025 4018 2047 4022
rect 2051 4018 2071 4022
rect 2075 4018 2327 4022
rect 2331 4018 2591 4022
rect 2595 4018 2839 4022
rect 2843 4018 3087 4022
rect 3091 4018 3343 4022
rect 3347 4018 3943 4022
rect 3947 4018 3967 4022
rect 2025 4017 3967 4018
rect 3973 4017 3974 4023
rect 84 3997 85 4003
rect 91 4002 2019 4003
rect 91 3998 111 4002
rect 115 3998 311 4002
rect 315 3998 511 4002
rect 515 3998 703 4002
rect 707 3998 887 4002
rect 891 3998 1063 4002
rect 1067 3998 1231 4002
rect 1235 3998 1383 4002
rect 1387 3998 1519 4002
rect 1523 3998 1655 4002
rect 1659 3998 1791 4002
rect 1795 3998 1903 4002
rect 1907 3998 2007 4002
rect 2011 3998 2019 4002
rect 91 3997 2019 3998
rect 2025 3997 2026 4003
rect 2030 3941 2031 3947
rect 2037 3946 3979 3947
rect 2037 3942 2047 3946
rect 2051 3942 2071 3946
rect 2075 3942 2127 3946
rect 2131 3942 2271 3946
rect 2275 3942 2327 3946
rect 2331 3942 2439 3946
rect 2443 3942 2591 3946
rect 2595 3942 2615 3946
rect 2619 3942 2799 3946
rect 2803 3942 2839 3946
rect 2843 3942 2983 3946
rect 2987 3942 3087 3946
rect 3091 3942 3175 3946
rect 3179 3942 3343 3946
rect 3347 3942 3367 3946
rect 3371 3942 3559 3946
rect 3563 3942 3943 3946
rect 3947 3942 3979 3946
rect 2037 3941 3979 3942
rect 3985 3941 3986 3947
rect 96 3921 97 3927
rect 103 3926 2031 3927
rect 103 3922 111 3926
rect 115 3922 279 3926
rect 283 3922 311 3926
rect 315 3922 415 3926
rect 419 3922 511 3926
rect 515 3922 567 3926
rect 571 3922 703 3926
rect 707 3922 735 3926
rect 739 3922 887 3926
rect 891 3922 911 3926
rect 915 3922 1063 3926
rect 1067 3922 1095 3926
rect 1099 3922 1231 3926
rect 1235 3922 1287 3926
rect 1291 3922 1383 3926
rect 1387 3922 1479 3926
rect 1483 3922 1519 3926
rect 1523 3922 1655 3926
rect 1659 3922 1679 3926
rect 1683 3922 1791 3926
rect 1795 3922 1903 3926
rect 1907 3922 2007 3926
rect 2011 3922 2031 3926
rect 103 3921 2031 3922
rect 2037 3921 2038 3927
rect 2018 3865 2019 3871
rect 2025 3870 3967 3871
rect 2025 3866 2047 3870
rect 2051 3866 2127 3870
rect 2131 3866 2263 3870
rect 2267 3866 2271 3870
rect 2275 3866 2375 3870
rect 2379 3866 2439 3870
rect 2443 3866 2495 3870
rect 2499 3866 2615 3870
rect 2619 3866 2631 3870
rect 2635 3866 2775 3870
rect 2779 3866 2799 3870
rect 2803 3866 2919 3870
rect 2923 3866 2983 3870
rect 2987 3866 3063 3870
rect 3067 3866 3175 3870
rect 3179 3866 3207 3870
rect 3211 3866 3343 3870
rect 3347 3866 3367 3870
rect 3371 3866 3471 3870
rect 3475 3866 3559 3870
rect 3563 3866 3599 3870
rect 3603 3866 3727 3870
rect 3731 3866 3839 3870
rect 3843 3866 3943 3870
rect 3947 3866 3967 3870
rect 2025 3865 3967 3866
rect 3973 3865 3974 3871
rect 84 3837 85 3843
rect 91 3842 2019 3843
rect 91 3838 111 3842
rect 115 3838 231 3842
rect 235 3838 279 3842
rect 283 3838 335 3842
rect 339 3838 415 3842
rect 419 3838 439 3842
rect 443 3838 535 3842
rect 539 3838 567 3842
rect 571 3838 631 3842
rect 635 3838 727 3842
rect 731 3838 735 3842
rect 739 3838 831 3842
rect 835 3838 911 3842
rect 915 3838 935 3842
rect 939 3838 1039 3842
rect 1043 3838 1095 3842
rect 1099 3838 1151 3842
rect 1155 3838 1263 3842
rect 1267 3838 1287 3842
rect 1291 3838 1383 3842
rect 1387 3838 1479 3842
rect 1483 3838 1503 3842
rect 1507 3838 1631 3842
rect 1635 3838 1679 3842
rect 1683 3838 2007 3842
rect 2011 3838 2019 3842
rect 91 3837 2019 3838
rect 2025 3837 2026 3843
rect 2030 3773 2031 3779
rect 2037 3778 3979 3779
rect 2037 3774 2047 3778
rect 2051 3774 2071 3778
rect 2075 3774 2183 3778
rect 2187 3774 2263 3778
rect 2267 3774 2327 3778
rect 2331 3774 2375 3778
rect 2379 3774 2479 3778
rect 2483 3774 2495 3778
rect 2499 3774 2631 3778
rect 2635 3774 2639 3778
rect 2643 3774 2775 3778
rect 2779 3774 2807 3778
rect 2811 3774 2919 3778
rect 2923 3774 2983 3778
rect 2987 3774 3063 3778
rect 3067 3774 3159 3778
rect 3163 3774 3207 3778
rect 3211 3774 3335 3778
rect 3339 3774 3343 3778
rect 3347 3774 3471 3778
rect 3475 3774 3511 3778
rect 3515 3774 3599 3778
rect 3603 3774 3687 3778
rect 3691 3774 3727 3778
rect 3731 3774 3839 3778
rect 3843 3774 3943 3778
rect 3947 3774 3979 3778
rect 2037 3773 3979 3774
rect 3985 3773 3986 3779
rect 96 3761 97 3767
rect 103 3766 2031 3767
rect 103 3762 111 3766
rect 115 3762 159 3766
rect 163 3762 231 3766
rect 235 3762 335 3766
rect 339 3762 351 3766
rect 355 3762 439 3766
rect 443 3762 535 3766
rect 539 3762 551 3766
rect 555 3762 631 3766
rect 635 3762 727 3766
rect 731 3762 751 3766
rect 755 3762 831 3766
rect 835 3762 935 3766
rect 939 3762 959 3766
rect 963 3762 1039 3766
rect 1043 3762 1151 3766
rect 1155 3762 1167 3766
rect 1171 3762 1263 3766
rect 1267 3762 1383 3766
rect 1387 3762 1503 3766
rect 1507 3762 1607 3766
rect 1611 3762 1631 3766
rect 1635 3762 2007 3766
rect 2011 3762 2031 3766
rect 103 3761 2031 3762
rect 2037 3761 2038 3767
rect 2018 3685 2019 3691
rect 2025 3690 3967 3691
rect 2025 3686 2047 3690
rect 2051 3686 2071 3690
rect 2075 3686 2183 3690
rect 2187 3686 2199 3690
rect 2203 3686 2327 3690
rect 2331 3686 2367 3690
rect 2371 3686 2479 3690
rect 2483 3686 2551 3690
rect 2555 3686 2639 3690
rect 2643 3686 2735 3690
rect 2739 3686 2807 3690
rect 2811 3686 2927 3690
rect 2931 3686 2983 3690
rect 2987 3686 3111 3690
rect 3115 3686 3159 3690
rect 3163 3686 3295 3690
rect 3299 3686 3335 3690
rect 3339 3686 3479 3690
rect 3483 3686 3511 3690
rect 3515 3686 3671 3690
rect 3675 3686 3687 3690
rect 3691 3686 3839 3690
rect 3843 3686 3943 3690
rect 3947 3686 3967 3690
rect 2025 3685 3967 3686
rect 3973 3685 3974 3691
rect 2018 3683 2026 3685
rect 84 3677 85 3683
rect 91 3682 2019 3683
rect 91 3678 111 3682
rect 115 3678 151 3682
rect 155 3678 159 3682
rect 163 3678 351 3682
rect 355 3678 383 3682
rect 387 3678 551 3682
rect 555 3678 615 3682
rect 619 3678 751 3682
rect 755 3678 839 3682
rect 843 3678 959 3682
rect 963 3678 1055 3682
rect 1059 3678 1167 3682
rect 1171 3678 1263 3682
rect 1267 3678 1383 3682
rect 1387 3678 1479 3682
rect 1483 3678 1607 3682
rect 1611 3678 1695 3682
rect 1699 3678 2007 3682
rect 2011 3678 2019 3682
rect 91 3677 2019 3678
rect 2025 3677 2026 3683
rect 2030 3605 2031 3611
rect 2037 3610 3979 3611
rect 2037 3606 2047 3610
rect 2051 3606 2071 3610
rect 2075 3606 2103 3610
rect 2107 3606 2199 3610
rect 2203 3606 2279 3610
rect 2283 3606 2367 3610
rect 2371 3606 2471 3610
rect 2475 3606 2551 3610
rect 2555 3606 2671 3610
rect 2675 3606 2735 3610
rect 2739 3606 2871 3610
rect 2875 3606 2927 3610
rect 2931 3606 3063 3610
rect 3067 3606 3111 3610
rect 3115 3606 3255 3610
rect 3259 3606 3295 3610
rect 3299 3606 3447 3610
rect 3451 3606 3479 3610
rect 3483 3606 3639 3610
rect 3643 3606 3671 3610
rect 3675 3606 3839 3610
rect 3843 3606 3943 3610
rect 3947 3606 3979 3610
rect 2037 3605 3979 3606
rect 3985 3605 3986 3611
rect 2030 3603 2038 3605
rect 96 3597 97 3603
rect 103 3602 2031 3603
rect 103 3598 111 3602
rect 115 3598 151 3602
rect 155 3598 167 3602
rect 171 3598 359 3602
rect 363 3598 383 3602
rect 387 3598 559 3602
rect 563 3598 615 3602
rect 619 3598 775 3602
rect 779 3598 839 3602
rect 843 3598 991 3602
rect 995 3598 1055 3602
rect 1059 3598 1215 3602
rect 1219 3598 1263 3602
rect 1267 3598 1447 3602
rect 1451 3598 1479 3602
rect 1483 3598 1687 3602
rect 1691 3598 1695 3602
rect 1699 3598 2007 3602
rect 2011 3598 2031 3602
rect 103 3597 2031 3598
rect 2037 3597 2038 3603
rect 2018 3525 2019 3531
rect 2025 3530 3967 3531
rect 2025 3526 2047 3530
rect 2051 3526 2103 3530
rect 2107 3526 2279 3530
rect 2283 3526 2327 3530
rect 2331 3526 2447 3530
rect 2451 3526 2471 3530
rect 2475 3526 2583 3530
rect 2587 3526 2671 3530
rect 2675 3526 2735 3530
rect 2739 3526 2871 3530
rect 2875 3526 2911 3530
rect 2915 3526 3063 3530
rect 3067 3526 3111 3530
rect 3115 3526 3255 3530
rect 3259 3526 3335 3530
rect 3339 3526 3447 3530
rect 3451 3526 3567 3530
rect 3571 3526 3639 3530
rect 3643 3526 3807 3530
rect 3811 3526 3839 3530
rect 3843 3526 3943 3530
rect 3947 3526 3967 3530
rect 2025 3525 3967 3526
rect 3973 3525 3974 3531
rect 84 3513 85 3519
rect 91 3518 2019 3519
rect 91 3514 111 3518
rect 115 3514 167 3518
rect 171 3514 295 3518
rect 299 3514 359 3518
rect 363 3514 431 3518
rect 435 3514 559 3518
rect 563 3514 583 3518
rect 587 3514 743 3518
rect 747 3514 775 3518
rect 779 3514 911 3518
rect 915 3514 991 3518
rect 995 3514 1079 3518
rect 1083 3514 1215 3518
rect 1219 3514 1247 3518
rect 1251 3514 1423 3518
rect 1427 3514 1447 3518
rect 1451 3514 1599 3518
rect 1603 3514 1687 3518
rect 1691 3514 1775 3518
rect 1779 3514 2007 3518
rect 2011 3514 2019 3518
rect 91 3513 2019 3514
rect 2025 3513 2026 3519
rect 2030 3449 2031 3455
rect 2037 3454 3979 3455
rect 2037 3450 2047 3454
rect 2051 3450 2327 3454
rect 2331 3450 2447 3454
rect 2451 3450 2551 3454
rect 2555 3450 2583 3454
rect 2587 3450 2663 3454
rect 2667 3450 2735 3454
rect 2739 3450 2775 3454
rect 2779 3450 2903 3454
rect 2907 3450 2911 3454
rect 2915 3450 3047 3454
rect 3051 3450 3111 3454
rect 3115 3450 3207 3454
rect 3211 3450 3335 3454
rect 3339 3450 3383 3454
rect 3387 3450 3567 3454
rect 3571 3450 3751 3454
rect 3755 3450 3807 3454
rect 3811 3450 3943 3454
rect 3947 3450 3979 3454
rect 2037 3449 3979 3450
rect 3985 3449 3986 3455
rect 96 3417 97 3423
rect 103 3422 2031 3423
rect 103 3418 111 3422
rect 115 3418 295 3422
rect 299 3418 431 3422
rect 435 3418 495 3422
rect 499 3418 583 3422
rect 587 3418 647 3422
rect 651 3418 743 3422
rect 747 3418 799 3422
rect 803 3418 911 3422
rect 915 3418 959 3422
rect 963 3418 1079 3422
rect 1083 3418 1127 3422
rect 1131 3418 1247 3422
rect 1251 3418 1295 3422
rect 1299 3418 1423 3422
rect 1427 3418 1463 3422
rect 1467 3418 1599 3422
rect 1603 3418 1639 3422
rect 1643 3418 1775 3422
rect 1779 3418 1815 3422
rect 1819 3418 2007 3422
rect 2011 3418 2031 3422
rect 103 3417 2031 3418
rect 2037 3417 2038 3423
rect 2018 3361 2019 3367
rect 2025 3366 3967 3367
rect 2025 3362 2047 3366
rect 2051 3362 2447 3366
rect 2451 3362 2551 3366
rect 2555 3362 2567 3366
rect 2571 3362 2663 3366
rect 2667 3362 2719 3366
rect 2723 3362 2775 3366
rect 2779 3362 2871 3366
rect 2875 3362 2903 3366
rect 2907 3362 3023 3366
rect 3027 3362 3047 3366
rect 3051 3362 3175 3366
rect 3179 3362 3207 3366
rect 3211 3362 3327 3366
rect 3331 3362 3383 3366
rect 3387 3362 3479 3366
rect 3483 3362 3567 3366
rect 3571 3362 3631 3366
rect 3635 3362 3751 3366
rect 3755 3362 3783 3366
rect 3787 3362 3943 3366
rect 3947 3362 3967 3366
rect 2025 3361 3967 3362
rect 3973 3361 3974 3367
rect 84 3329 85 3335
rect 91 3334 2019 3335
rect 91 3330 111 3334
rect 115 3330 135 3334
rect 139 3330 295 3334
rect 299 3330 479 3334
rect 483 3330 495 3334
rect 499 3330 647 3334
rect 651 3330 671 3334
rect 675 3330 799 3334
rect 803 3330 863 3334
rect 867 3330 959 3334
rect 963 3330 1055 3334
rect 1059 3330 1127 3334
rect 1131 3330 1247 3334
rect 1251 3330 1295 3334
rect 1299 3330 1439 3334
rect 1443 3330 1463 3334
rect 1467 3330 1631 3334
rect 1635 3330 1639 3334
rect 1643 3330 1815 3334
rect 1819 3330 1823 3334
rect 1827 3330 2007 3334
rect 2011 3330 2019 3334
rect 91 3329 2019 3330
rect 2025 3329 2026 3335
rect 2030 3281 2031 3287
rect 2037 3286 3979 3287
rect 2037 3282 2047 3286
rect 2051 3282 2415 3286
rect 2419 3282 2551 3286
rect 2555 3282 2567 3286
rect 2571 3282 2687 3286
rect 2691 3282 2719 3286
rect 2723 3282 2831 3286
rect 2835 3282 2871 3286
rect 2875 3282 2975 3286
rect 2979 3282 3023 3286
rect 3027 3282 3119 3286
rect 3123 3282 3175 3286
rect 3179 3282 3255 3286
rect 3259 3282 3327 3286
rect 3331 3282 3383 3286
rect 3387 3282 3479 3286
rect 3483 3282 3503 3286
rect 3507 3282 3623 3286
rect 3627 3282 3631 3286
rect 3635 3282 3743 3286
rect 3747 3282 3783 3286
rect 3787 3282 3839 3286
rect 3843 3282 3943 3286
rect 3947 3282 3979 3286
rect 2037 3281 3979 3282
rect 3985 3281 3986 3287
rect 96 3249 97 3255
rect 103 3254 2031 3255
rect 103 3250 111 3254
rect 115 3250 135 3254
rect 139 3250 295 3254
rect 299 3250 319 3254
rect 323 3250 479 3254
rect 483 3250 519 3254
rect 523 3250 671 3254
rect 675 3250 719 3254
rect 723 3250 863 3254
rect 867 3250 911 3254
rect 915 3250 1055 3254
rect 1059 3250 1095 3254
rect 1099 3250 1247 3254
rect 1251 3250 1271 3254
rect 1275 3250 1439 3254
rect 1443 3250 1447 3254
rect 1451 3250 1623 3254
rect 1627 3250 1631 3254
rect 1635 3250 1799 3254
rect 1803 3250 1823 3254
rect 1827 3250 2007 3254
rect 2011 3250 2031 3254
rect 103 3249 2031 3250
rect 2037 3249 2038 3255
rect 2018 3193 2019 3199
rect 2025 3198 3967 3199
rect 2025 3194 2047 3198
rect 2051 3194 2247 3198
rect 2251 3194 2399 3198
rect 2403 3194 2415 3198
rect 2419 3194 2551 3198
rect 2555 3194 2559 3198
rect 2563 3194 2687 3198
rect 2691 3194 2727 3198
rect 2731 3194 2831 3198
rect 2835 3194 2903 3198
rect 2907 3194 2975 3198
rect 2979 3194 3079 3198
rect 3083 3194 3119 3198
rect 3123 3194 3255 3198
rect 3259 3194 3263 3198
rect 3267 3194 3383 3198
rect 3387 3194 3447 3198
rect 3451 3194 3503 3198
rect 3507 3194 3623 3198
rect 3627 3194 3631 3198
rect 3635 3194 3743 3198
rect 3747 3194 3815 3198
rect 3819 3194 3839 3198
rect 3843 3194 3943 3198
rect 3947 3194 3967 3198
rect 2025 3193 3967 3194
rect 3973 3193 3974 3199
rect 84 3165 85 3171
rect 91 3170 2019 3171
rect 91 3166 111 3170
rect 115 3166 135 3170
rect 139 3166 143 3170
rect 147 3166 319 3170
rect 323 3166 343 3170
rect 347 3166 519 3170
rect 523 3166 543 3170
rect 547 3166 719 3170
rect 723 3166 743 3170
rect 747 3166 911 3170
rect 915 3166 927 3170
rect 931 3166 1095 3170
rect 1099 3166 1103 3170
rect 1107 3166 1263 3170
rect 1267 3166 1271 3170
rect 1275 3166 1423 3170
rect 1427 3166 1447 3170
rect 1451 3166 1575 3170
rect 1579 3166 1623 3170
rect 1627 3166 1735 3170
rect 1739 3166 1799 3170
rect 1803 3166 2007 3170
rect 2011 3166 2019 3170
rect 91 3165 2019 3166
rect 2025 3165 2026 3171
rect 2030 3113 2031 3119
rect 2037 3118 3979 3119
rect 2037 3114 2047 3118
rect 2051 3114 2079 3118
rect 2083 3114 2223 3118
rect 2227 3114 2247 3118
rect 2251 3114 2375 3118
rect 2379 3114 2399 3118
rect 2403 3114 2527 3118
rect 2531 3114 2559 3118
rect 2563 3114 2687 3118
rect 2691 3114 2727 3118
rect 2731 3114 2855 3118
rect 2859 3114 2903 3118
rect 2907 3114 3039 3118
rect 3043 3114 3079 3118
rect 3083 3114 3231 3118
rect 3235 3114 3263 3118
rect 3267 3114 3431 3118
rect 3435 3114 3447 3118
rect 3451 3114 3631 3118
rect 3635 3114 3639 3118
rect 3643 3114 3815 3118
rect 3819 3114 3839 3118
rect 3843 3114 3943 3118
rect 3947 3114 3979 3118
rect 2037 3113 3979 3114
rect 3985 3113 3986 3119
rect 96 3089 97 3095
rect 103 3094 2031 3095
rect 103 3090 111 3094
rect 115 3090 143 3094
rect 147 3090 263 3094
rect 267 3090 343 3094
rect 347 3090 439 3094
rect 443 3090 543 3094
rect 547 3090 615 3094
rect 619 3090 743 3094
rect 747 3090 799 3094
rect 803 3090 927 3094
rect 931 3090 975 3094
rect 979 3090 1103 3094
rect 1107 3090 1143 3094
rect 1147 3090 1263 3094
rect 1267 3090 1303 3094
rect 1307 3090 1423 3094
rect 1427 3090 1455 3094
rect 1459 3090 1575 3094
rect 1579 3090 1607 3094
rect 1611 3090 1735 3094
rect 1739 3090 1767 3094
rect 1771 3090 2007 3094
rect 2011 3090 2031 3094
rect 103 3089 2031 3090
rect 2037 3089 2038 3095
rect 2018 3029 2019 3035
rect 2025 3034 3967 3035
rect 2025 3030 2047 3034
rect 2051 3030 2071 3034
rect 2075 3030 2079 3034
rect 2083 3030 2183 3034
rect 2187 3030 2223 3034
rect 2227 3030 2327 3034
rect 2331 3030 2375 3034
rect 2379 3030 2479 3034
rect 2483 3030 2527 3034
rect 2531 3030 2655 3034
rect 2659 3030 2687 3034
rect 2691 3030 2855 3034
rect 2859 3030 3039 3034
rect 3043 3030 3087 3034
rect 3091 3030 3231 3034
rect 3235 3030 3335 3034
rect 3339 3030 3431 3034
rect 3435 3030 3599 3034
rect 3603 3030 3639 3034
rect 3643 3030 3839 3034
rect 3843 3030 3943 3034
rect 3947 3030 3967 3034
rect 2025 3029 3967 3030
rect 3973 3029 3974 3035
rect 84 2989 85 2995
rect 91 2994 2019 2995
rect 91 2990 111 2994
rect 115 2990 263 2994
rect 267 2990 343 2994
rect 347 2990 439 2994
rect 443 2990 543 2994
rect 547 2990 615 2994
rect 619 2990 655 2994
rect 659 2990 783 2994
rect 787 2990 799 2994
rect 803 2990 935 2994
rect 939 2990 975 2994
rect 979 2990 1103 2994
rect 1107 2990 1143 2994
rect 1147 2990 1295 2994
rect 1299 2990 1303 2994
rect 1307 2990 1455 2994
rect 1459 2990 1495 2994
rect 1499 2990 1607 2994
rect 1611 2990 1711 2994
rect 1715 2990 1767 2994
rect 1771 2990 1903 2994
rect 1907 2990 2007 2994
rect 2011 2990 2019 2994
rect 91 2989 2019 2990
rect 2025 2989 2026 2995
rect 2030 2949 2031 2955
rect 2037 2954 3979 2955
rect 2037 2950 2047 2954
rect 2051 2950 2071 2954
rect 2075 2950 2183 2954
rect 2187 2950 2263 2954
rect 2267 2950 2327 2954
rect 2331 2950 2479 2954
rect 2483 2950 2487 2954
rect 2491 2950 2655 2954
rect 2659 2950 2735 2954
rect 2739 2950 2855 2954
rect 2859 2950 2999 2954
rect 3003 2950 3087 2954
rect 3091 2950 3279 2954
rect 3283 2950 3335 2954
rect 3339 2950 3567 2954
rect 3571 2950 3599 2954
rect 3603 2950 3839 2954
rect 3843 2950 3943 2954
rect 3947 2950 3979 2954
rect 2037 2949 3979 2950
rect 3985 2949 3986 2955
rect 96 2913 97 2919
rect 103 2918 2031 2919
rect 103 2914 111 2918
rect 115 2914 207 2918
rect 211 2914 327 2918
rect 331 2914 343 2918
rect 347 2914 439 2918
rect 443 2914 447 2918
rect 451 2914 543 2918
rect 547 2914 575 2918
rect 579 2914 655 2918
rect 659 2914 703 2918
rect 707 2914 783 2918
rect 787 2914 847 2918
rect 851 2914 935 2918
rect 939 2914 999 2918
rect 1003 2914 1103 2918
rect 1107 2914 1167 2918
rect 1171 2914 1295 2918
rect 1299 2914 1351 2918
rect 1355 2914 1495 2918
rect 1499 2914 1535 2918
rect 1539 2914 1711 2918
rect 1715 2914 1727 2918
rect 1731 2914 1903 2918
rect 1907 2914 2007 2918
rect 2011 2914 2031 2918
rect 103 2913 2031 2914
rect 2037 2913 2038 2919
rect 2018 2865 2019 2871
rect 2025 2870 3967 2871
rect 2025 2866 2047 2870
rect 2051 2866 2071 2870
rect 2075 2866 2263 2870
rect 2267 2866 2487 2870
rect 2491 2866 2671 2870
rect 2675 2866 2735 2870
rect 2739 2866 2887 2870
rect 2891 2866 2999 2870
rect 3003 2866 3095 2870
rect 3099 2866 3279 2870
rect 3283 2866 3287 2870
rect 3291 2866 3479 2870
rect 3483 2866 3567 2870
rect 3571 2866 3671 2870
rect 3675 2866 3839 2870
rect 3843 2866 3943 2870
rect 3947 2866 3967 2870
rect 2025 2865 3967 2866
rect 3973 2865 3974 2871
rect 84 2833 85 2839
rect 91 2838 2019 2839
rect 91 2834 111 2838
rect 115 2834 135 2838
rect 139 2834 207 2838
rect 211 2834 247 2838
rect 251 2834 327 2838
rect 331 2834 399 2838
rect 403 2834 447 2838
rect 451 2834 551 2838
rect 555 2834 575 2838
rect 579 2834 703 2838
rect 707 2834 711 2838
rect 715 2834 847 2838
rect 851 2834 879 2838
rect 883 2834 999 2838
rect 1003 2834 1047 2838
rect 1051 2834 1167 2838
rect 1171 2834 1223 2838
rect 1227 2834 1351 2838
rect 1355 2834 1399 2838
rect 1403 2834 1535 2838
rect 1539 2834 1575 2838
rect 1579 2834 1727 2838
rect 1731 2834 1751 2838
rect 1755 2834 1903 2838
rect 1907 2834 2007 2838
rect 2011 2834 2019 2838
rect 91 2833 2019 2834
rect 2025 2833 2026 2839
rect 2030 2789 2031 2795
rect 2037 2794 3979 2795
rect 2037 2790 2047 2794
rect 2051 2790 2071 2794
rect 2075 2790 2199 2794
rect 2203 2790 2343 2794
rect 2347 2790 2479 2794
rect 2483 2790 2607 2794
rect 2611 2790 2671 2794
rect 2675 2790 2727 2794
rect 2731 2790 2839 2794
rect 2843 2790 2887 2794
rect 2891 2790 2943 2794
rect 2947 2790 3047 2794
rect 3051 2790 3095 2794
rect 3099 2790 3143 2794
rect 3147 2790 3239 2794
rect 3243 2790 3287 2794
rect 3291 2790 3343 2794
rect 3347 2790 3447 2794
rect 3451 2790 3479 2794
rect 3483 2790 3551 2794
rect 3555 2790 3647 2794
rect 3651 2790 3671 2794
rect 3675 2790 3743 2794
rect 3747 2790 3839 2794
rect 3843 2790 3943 2794
rect 3947 2790 3979 2794
rect 2037 2789 3979 2790
rect 3985 2789 3986 2795
rect 96 2749 97 2755
rect 103 2754 2031 2755
rect 103 2750 111 2754
rect 115 2750 135 2754
rect 139 2750 247 2754
rect 251 2750 255 2754
rect 259 2750 399 2754
rect 403 2750 407 2754
rect 411 2750 551 2754
rect 555 2750 575 2754
rect 579 2750 711 2754
rect 715 2750 743 2754
rect 747 2750 879 2754
rect 883 2750 919 2754
rect 923 2750 1047 2754
rect 1051 2750 1087 2754
rect 1091 2750 1223 2754
rect 1227 2750 1255 2754
rect 1259 2750 1399 2754
rect 1403 2750 1423 2754
rect 1427 2750 1575 2754
rect 1579 2750 1599 2754
rect 1603 2750 1751 2754
rect 1755 2750 1903 2754
rect 1907 2750 2007 2754
rect 2011 2750 2031 2754
rect 103 2749 2031 2750
rect 2037 2749 2038 2755
rect 2018 2693 2019 2699
rect 2025 2698 3967 2699
rect 2025 2694 2047 2698
rect 2051 2694 2071 2698
rect 2075 2694 2095 2698
rect 2099 2694 2199 2698
rect 2203 2694 2263 2698
rect 2267 2694 2343 2698
rect 2347 2694 2439 2698
rect 2443 2694 2479 2698
rect 2483 2694 2607 2698
rect 2611 2694 2615 2698
rect 2619 2694 2727 2698
rect 2731 2694 2783 2698
rect 2787 2694 2839 2698
rect 2843 2694 2943 2698
rect 2947 2694 3047 2698
rect 3051 2694 3095 2698
rect 3099 2694 3143 2698
rect 3147 2694 3239 2698
rect 3243 2694 3343 2698
rect 3347 2694 3383 2698
rect 3387 2694 3447 2698
rect 3451 2694 3535 2698
rect 3539 2694 3551 2698
rect 3555 2694 3647 2698
rect 3651 2694 3743 2698
rect 3747 2694 3839 2698
rect 3843 2694 3943 2698
rect 3947 2694 3967 2698
rect 2025 2693 3967 2694
rect 3973 2693 3974 2699
rect 84 2673 85 2679
rect 91 2678 2019 2679
rect 91 2674 111 2678
rect 115 2674 135 2678
rect 139 2674 167 2678
rect 171 2674 255 2678
rect 259 2674 359 2678
rect 363 2674 407 2678
rect 411 2674 559 2678
rect 563 2674 575 2678
rect 579 2674 743 2678
rect 747 2674 759 2678
rect 763 2674 919 2678
rect 923 2674 951 2678
rect 955 2674 1087 2678
rect 1091 2674 1143 2678
rect 1147 2674 1255 2678
rect 1259 2674 1327 2678
rect 1331 2674 1423 2678
rect 1427 2674 1511 2678
rect 1515 2674 1599 2678
rect 1603 2674 1703 2678
rect 1707 2674 2007 2678
rect 2011 2674 2019 2678
rect 91 2673 2019 2674
rect 2025 2673 2026 2679
rect 2030 2609 2031 2615
rect 2037 2614 3979 2615
rect 2037 2610 2047 2614
rect 2051 2610 2095 2614
rect 2099 2610 2215 2614
rect 2219 2610 2263 2614
rect 2267 2610 2367 2614
rect 2371 2610 2439 2614
rect 2443 2610 2519 2614
rect 2523 2610 2615 2614
rect 2619 2610 2671 2614
rect 2675 2610 2783 2614
rect 2787 2610 2815 2614
rect 2819 2610 2943 2614
rect 2947 2610 2951 2614
rect 2955 2610 3087 2614
rect 3091 2610 3095 2614
rect 3099 2610 3223 2614
rect 3227 2610 3239 2614
rect 3243 2610 3367 2614
rect 3371 2610 3383 2614
rect 3387 2610 3535 2614
rect 3539 2610 3943 2614
rect 3947 2610 3979 2614
rect 2037 2609 3979 2610
rect 3985 2609 3986 2615
rect 96 2581 97 2587
rect 103 2586 2031 2587
rect 103 2582 111 2586
rect 115 2582 167 2586
rect 171 2582 359 2586
rect 363 2582 559 2586
rect 563 2582 575 2586
rect 579 2582 687 2586
rect 691 2582 759 2586
rect 763 2582 807 2586
rect 811 2582 935 2586
rect 939 2582 951 2586
rect 955 2582 1071 2586
rect 1075 2582 1143 2586
rect 1147 2582 1207 2586
rect 1211 2582 1327 2586
rect 1331 2582 1351 2586
rect 1355 2582 1495 2586
rect 1499 2582 1511 2586
rect 1515 2582 1647 2586
rect 1651 2582 1703 2586
rect 1707 2582 1799 2586
rect 1803 2582 2007 2586
rect 2011 2582 2031 2586
rect 103 2581 2031 2582
rect 2037 2581 2038 2587
rect 2018 2529 2019 2535
rect 2025 2534 3967 2535
rect 2025 2530 2047 2534
rect 2051 2530 2095 2534
rect 2099 2530 2215 2534
rect 2219 2530 2343 2534
rect 2347 2530 2367 2534
rect 2371 2530 2471 2534
rect 2475 2530 2519 2534
rect 2523 2530 2599 2534
rect 2603 2530 2671 2534
rect 2675 2530 2719 2534
rect 2723 2530 2815 2534
rect 2819 2530 2839 2534
rect 2843 2530 2951 2534
rect 2955 2530 2967 2534
rect 2971 2530 3087 2534
rect 3091 2530 3095 2534
rect 3099 2530 3223 2534
rect 3227 2530 3367 2534
rect 3371 2530 3943 2534
rect 3947 2530 3967 2534
rect 2025 2529 3967 2530
rect 3973 2529 3974 2535
rect 84 2501 85 2507
rect 91 2506 2019 2507
rect 91 2502 111 2506
rect 115 2502 503 2506
rect 507 2502 575 2506
rect 579 2502 607 2506
rect 611 2502 687 2506
rect 691 2502 719 2506
rect 723 2502 807 2506
rect 811 2502 847 2506
rect 851 2502 935 2506
rect 939 2502 983 2506
rect 987 2502 1071 2506
rect 1075 2502 1127 2506
rect 1131 2502 1207 2506
rect 1211 2502 1279 2506
rect 1283 2502 1351 2506
rect 1355 2502 1431 2506
rect 1435 2502 1495 2506
rect 1499 2502 1583 2506
rect 1587 2502 1647 2506
rect 1651 2502 1743 2506
rect 1747 2502 1799 2506
rect 1803 2502 1903 2506
rect 1907 2502 2007 2506
rect 2011 2502 2019 2506
rect 91 2501 2019 2502
rect 2025 2501 2026 2507
rect 2030 2441 2031 2447
rect 2037 2446 3979 2447
rect 2037 2442 2047 2446
rect 2051 2442 2071 2446
rect 2075 2442 2095 2446
rect 2099 2442 2191 2446
rect 2195 2442 2215 2446
rect 2219 2442 2319 2446
rect 2323 2442 2343 2446
rect 2347 2442 2439 2446
rect 2443 2442 2471 2446
rect 2475 2442 2559 2446
rect 2563 2442 2599 2446
rect 2603 2442 2679 2446
rect 2683 2442 2719 2446
rect 2723 2442 2791 2446
rect 2795 2442 2839 2446
rect 2843 2442 2911 2446
rect 2915 2442 2967 2446
rect 2971 2442 3031 2446
rect 3035 2442 3095 2446
rect 3099 2442 3151 2446
rect 3155 2442 3223 2446
rect 3227 2442 3943 2446
rect 3947 2442 3979 2446
rect 2037 2441 3979 2442
rect 3985 2441 3986 2447
rect 96 2409 97 2415
rect 103 2414 2031 2415
rect 103 2410 111 2414
rect 115 2410 503 2414
rect 507 2410 535 2414
rect 539 2410 607 2414
rect 611 2410 671 2414
rect 675 2410 719 2414
rect 723 2410 815 2414
rect 819 2410 847 2414
rect 851 2410 959 2414
rect 963 2410 983 2414
rect 987 2410 1103 2414
rect 1107 2410 1127 2414
rect 1131 2410 1247 2414
rect 1251 2410 1279 2414
rect 1283 2410 1391 2414
rect 1395 2410 1431 2414
rect 1435 2410 1527 2414
rect 1531 2410 1583 2414
rect 1587 2410 1655 2414
rect 1659 2410 1743 2414
rect 1747 2410 1791 2414
rect 1795 2410 1903 2414
rect 1907 2410 2007 2414
rect 2011 2410 2031 2414
rect 103 2409 2031 2410
rect 2037 2409 2038 2415
rect 2018 2361 2019 2367
rect 2025 2366 3967 2367
rect 2025 2362 2047 2366
rect 2051 2362 2071 2366
rect 2075 2362 2167 2366
rect 2171 2362 2191 2366
rect 2195 2362 2319 2366
rect 2323 2362 2359 2366
rect 2363 2362 2439 2366
rect 2443 2362 2535 2366
rect 2539 2362 2559 2366
rect 2563 2362 2679 2366
rect 2683 2362 2703 2366
rect 2707 2362 2791 2366
rect 2795 2362 2871 2366
rect 2875 2362 2911 2366
rect 2915 2362 3031 2366
rect 3035 2362 3151 2366
rect 3155 2362 3199 2366
rect 3203 2362 3943 2366
rect 3947 2362 3967 2366
rect 2025 2361 3967 2362
rect 3973 2361 3974 2367
rect 84 2329 85 2335
rect 91 2334 2019 2335
rect 91 2330 111 2334
rect 115 2330 535 2334
rect 539 2330 647 2334
rect 651 2330 671 2334
rect 675 2330 767 2334
rect 771 2330 815 2334
rect 819 2330 895 2334
rect 899 2330 959 2334
rect 963 2330 1031 2334
rect 1035 2330 1103 2334
rect 1107 2330 1167 2334
rect 1171 2330 1247 2334
rect 1251 2330 1295 2334
rect 1299 2330 1391 2334
rect 1395 2330 1423 2334
rect 1427 2330 1527 2334
rect 1531 2330 1551 2334
rect 1555 2330 1655 2334
rect 1659 2330 1671 2334
rect 1675 2330 1791 2334
rect 1795 2330 1799 2334
rect 1803 2330 1903 2334
rect 1907 2330 2007 2334
rect 2011 2330 2019 2334
rect 91 2329 2019 2330
rect 2025 2329 2026 2335
rect 2030 2285 2031 2291
rect 2037 2290 3979 2291
rect 2037 2286 2047 2290
rect 2051 2286 2071 2290
rect 2075 2286 2167 2290
rect 2171 2286 2287 2290
rect 2291 2286 2359 2290
rect 2363 2286 2423 2290
rect 2427 2286 2535 2290
rect 2539 2286 2559 2290
rect 2563 2286 2703 2290
rect 2707 2286 2839 2290
rect 2843 2286 2871 2290
rect 2875 2286 2983 2290
rect 2987 2286 3031 2290
rect 3035 2286 3127 2290
rect 3131 2286 3199 2290
rect 3203 2286 3271 2290
rect 3275 2286 3943 2290
rect 3947 2286 3979 2290
rect 2037 2285 3979 2286
rect 3985 2285 3986 2291
rect 96 2249 97 2255
rect 103 2254 2031 2255
rect 103 2250 111 2254
rect 115 2250 415 2254
rect 419 2250 535 2254
rect 539 2250 647 2254
rect 651 2250 671 2254
rect 675 2250 767 2254
rect 771 2250 823 2254
rect 827 2250 895 2254
rect 899 2250 991 2254
rect 995 2250 1031 2254
rect 1035 2250 1167 2254
rect 1171 2250 1175 2254
rect 1179 2250 1295 2254
rect 1299 2250 1367 2254
rect 1371 2250 1423 2254
rect 1427 2250 1551 2254
rect 1555 2250 1567 2254
rect 1571 2250 1671 2254
rect 1675 2250 1767 2254
rect 1771 2250 1799 2254
rect 1803 2250 1903 2254
rect 1907 2250 2007 2254
rect 2011 2250 2031 2254
rect 103 2249 2031 2250
rect 2037 2249 2038 2255
rect 2018 2209 2019 2215
rect 2025 2214 3967 2215
rect 2025 2210 2047 2214
rect 2051 2210 2071 2214
rect 2075 2210 2167 2214
rect 2171 2210 2287 2214
rect 2291 2210 2295 2214
rect 2299 2210 2423 2214
rect 2427 2210 2503 2214
rect 2507 2210 2559 2214
rect 2563 2210 2687 2214
rect 2691 2210 2703 2214
rect 2707 2210 2839 2214
rect 2843 2210 2863 2214
rect 2867 2210 2983 2214
rect 2987 2210 3023 2214
rect 3027 2210 3127 2214
rect 3131 2210 3175 2214
rect 3179 2210 3271 2214
rect 3275 2210 3319 2214
rect 3323 2210 3471 2214
rect 3475 2210 3943 2214
rect 3947 2210 3967 2214
rect 2025 2209 3967 2210
rect 3973 2209 3974 2215
rect 84 2165 85 2171
rect 91 2170 2019 2171
rect 91 2166 111 2170
rect 115 2166 135 2170
rect 139 2166 247 2170
rect 251 2166 391 2170
rect 395 2166 415 2170
rect 419 2166 535 2170
rect 539 2166 551 2170
rect 555 2166 671 2170
rect 675 2166 711 2170
rect 715 2166 823 2170
rect 827 2166 871 2170
rect 875 2166 991 2170
rect 995 2166 1031 2170
rect 1035 2166 1175 2170
rect 1179 2166 1191 2170
rect 1195 2166 1351 2170
rect 1355 2166 1367 2170
rect 1371 2166 1511 2170
rect 1515 2166 1567 2170
rect 1571 2166 1679 2170
rect 1683 2166 1767 2170
rect 1771 2166 2007 2170
rect 2011 2166 2019 2170
rect 91 2165 2019 2166
rect 2025 2165 2026 2171
rect 2030 2109 2031 2115
rect 2037 2114 3979 2115
rect 2037 2110 2047 2114
rect 2051 2110 2071 2114
rect 2075 2110 2295 2114
rect 2299 2110 2399 2114
rect 2403 2110 2495 2114
rect 2499 2110 2503 2114
rect 2507 2110 2591 2114
rect 2595 2110 2687 2114
rect 2691 2110 2783 2114
rect 2787 2110 2863 2114
rect 2867 2110 2879 2114
rect 2883 2110 2975 2114
rect 2979 2110 3023 2114
rect 3027 2110 3071 2114
rect 3075 2110 3167 2114
rect 3171 2110 3175 2114
rect 3179 2110 3263 2114
rect 3267 2110 3319 2114
rect 3323 2110 3359 2114
rect 3363 2110 3455 2114
rect 3459 2110 3471 2114
rect 3475 2110 3551 2114
rect 3555 2110 3647 2114
rect 3651 2110 3743 2114
rect 3747 2110 3839 2114
rect 3843 2110 3943 2114
rect 3947 2110 3979 2114
rect 2037 2109 3979 2110
rect 3985 2109 3986 2115
rect 96 2081 97 2087
rect 103 2086 2031 2087
rect 103 2082 111 2086
rect 115 2082 135 2086
rect 139 2082 247 2086
rect 251 2082 391 2086
rect 395 2082 399 2086
rect 403 2082 551 2086
rect 555 2082 703 2086
rect 707 2082 711 2086
rect 715 2082 847 2086
rect 851 2082 871 2086
rect 875 2082 991 2086
rect 995 2082 1031 2086
rect 1035 2082 1127 2086
rect 1131 2082 1191 2086
rect 1195 2082 1255 2086
rect 1259 2082 1351 2086
rect 1355 2082 1383 2086
rect 1387 2082 1511 2086
rect 1515 2082 1519 2086
rect 1523 2082 1679 2086
rect 1683 2082 2007 2086
rect 2011 2082 2031 2086
rect 103 2081 2031 2082
rect 2037 2081 2038 2087
rect 2018 2033 2019 2039
rect 2025 2038 3967 2039
rect 2025 2034 2047 2038
rect 2051 2034 2191 2038
rect 2195 2034 2399 2038
rect 2403 2034 2495 2038
rect 2499 2034 2591 2038
rect 2595 2034 2647 2038
rect 2651 2034 2687 2038
rect 2691 2034 2783 2038
rect 2787 2034 2879 2038
rect 2883 2034 2919 2038
rect 2923 2034 2975 2038
rect 2979 2034 3071 2038
rect 3075 2034 3167 2038
rect 3171 2034 3215 2038
rect 3219 2034 3263 2038
rect 3267 2034 3359 2038
rect 3363 2034 3455 2038
rect 3459 2034 3527 2038
rect 3531 2034 3551 2038
rect 3555 2034 3647 2038
rect 3651 2034 3743 2038
rect 3747 2034 3839 2038
rect 3843 2034 3943 2038
rect 3947 2034 3967 2038
rect 2025 2033 3967 2034
rect 3973 2033 3974 2039
rect 84 1989 85 1995
rect 91 1994 2019 1995
rect 91 1990 111 1994
rect 115 1990 135 1994
rect 139 1990 231 1994
rect 235 1990 247 1994
rect 251 1990 391 1994
rect 395 1990 399 1994
rect 403 1990 551 1994
rect 555 1990 567 1994
rect 571 1990 703 1994
rect 707 1990 751 1994
rect 755 1990 847 1994
rect 851 1990 943 1994
rect 947 1990 991 1994
rect 995 1990 1127 1994
rect 1131 1990 1135 1994
rect 1139 1990 1255 1994
rect 1259 1990 1335 1994
rect 1339 1990 1383 1994
rect 1387 1990 1519 1994
rect 1523 1990 1543 1994
rect 1547 1990 2007 1994
rect 2011 1990 2019 1994
rect 91 1989 2019 1990
rect 2025 1989 2026 1995
rect 2030 1945 2031 1951
rect 2037 1950 3979 1951
rect 2037 1946 2047 1950
rect 2051 1946 2071 1950
rect 2075 1946 2191 1950
rect 2195 1946 2239 1950
rect 2243 1946 2399 1950
rect 2403 1946 2447 1950
rect 2451 1946 2647 1950
rect 2651 1946 2671 1950
rect 2675 1946 2895 1950
rect 2899 1946 2919 1950
rect 2923 1946 3127 1950
rect 3131 1946 3215 1950
rect 3219 1946 3359 1950
rect 3363 1946 3527 1950
rect 3531 1946 3591 1950
rect 3595 1946 3831 1950
rect 3835 1946 3839 1950
rect 3843 1946 3943 1950
rect 3947 1946 3979 1950
rect 2037 1945 3979 1946
rect 3985 1945 3986 1951
rect 96 1913 97 1919
rect 103 1918 2031 1919
rect 103 1914 111 1918
rect 115 1914 231 1918
rect 235 1914 391 1918
rect 395 1914 511 1918
rect 515 1914 567 1918
rect 571 1914 623 1918
rect 627 1914 743 1918
rect 747 1914 751 1918
rect 755 1914 863 1918
rect 867 1914 943 1918
rect 947 1914 983 1918
rect 987 1914 1103 1918
rect 1107 1914 1135 1918
rect 1139 1914 1223 1918
rect 1227 1914 1335 1918
rect 1339 1914 1455 1918
rect 1459 1914 1543 1918
rect 1547 1914 1575 1918
rect 1579 1914 1695 1918
rect 1699 1914 2007 1918
rect 2011 1914 2031 1918
rect 103 1913 2031 1914
rect 2037 1913 2038 1919
rect 2018 1869 2019 1875
rect 2025 1874 3967 1875
rect 2025 1870 2047 1874
rect 2051 1870 2071 1874
rect 2075 1870 2199 1874
rect 2203 1870 2239 1874
rect 2243 1870 2367 1874
rect 2371 1870 2447 1874
rect 2451 1870 2543 1874
rect 2547 1870 2671 1874
rect 2675 1870 2719 1874
rect 2723 1870 2887 1874
rect 2891 1870 2895 1874
rect 2899 1870 3039 1874
rect 3043 1870 3127 1874
rect 3131 1870 3183 1874
rect 3187 1870 3319 1874
rect 3323 1870 3359 1874
rect 3363 1870 3455 1874
rect 3459 1870 3583 1874
rect 3587 1870 3591 1874
rect 3595 1870 3711 1874
rect 3715 1870 3831 1874
rect 3835 1870 3839 1874
rect 3843 1870 3943 1874
rect 3947 1870 3967 1874
rect 2025 1869 3967 1870
rect 3973 1869 3974 1875
rect 84 1829 85 1835
rect 91 1834 2019 1835
rect 91 1830 111 1834
rect 115 1830 511 1834
rect 515 1830 615 1834
rect 619 1830 623 1834
rect 627 1830 711 1834
rect 715 1830 743 1834
rect 747 1830 815 1834
rect 819 1830 863 1834
rect 867 1830 927 1834
rect 931 1830 983 1834
rect 987 1830 1039 1834
rect 1043 1830 1103 1834
rect 1107 1830 1159 1834
rect 1163 1830 1223 1834
rect 1227 1830 1279 1834
rect 1283 1830 1335 1834
rect 1339 1830 1399 1834
rect 1403 1830 1455 1834
rect 1459 1830 1519 1834
rect 1523 1830 1575 1834
rect 1579 1830 1639 1834
rect 1643 1830 1695 1834
rect 1699 1830 2007 1834
rect 2011 1830 2019 1834
rect 91 1829 2019 1830
rect 2025 1829 2026 1835
rect 2030 1789 2031 1795
rect 2037 1794 3979 1795
rect 2037 1790 2047 1794
rect 2051 1790 2071 1794
rect 2075 1790 2183 1794
rect 2187 1790 2199 1794
rect 2203 1790 2327 1794
rect 2331 1790 2367 1794
rect 2371 1790 2487 1794
rect 2491 1790 2543 1794
rect 2547 1790 2655 1794
rect 2659 1790 2719 1794
rect 2723 1790 2831 1794
rect 2835 1790 2887 1794
rect 2891 1790 3023 1794
rect 3027 1790 3039 1794
rect 3043 1790 3183 1794
rect 3187 1790 3223 1794
rect 3227 1790 3319 1794
rect 3323 1790 3431 1794
rect 3435 1790 3455 1794
rect 3459 1790 3583 1794
rect 3587 1790 3647 1794
rect 3651 1790 3711 1794
rect 3715 1790 3839 1794
rect 3843 1790 3943 1794
rect 3947 1790 3979 1794
rect 2037 1789 3979 1790
rect 3985 1789 3986 1795
rect 96 1753 97 1759
rect 103 1758 2031 1759
rect 103 1754 111 1758
rect 115 1754 367 1758
rect 371 1754 495 1758
rect 499 1754 615 1758
rect 619 1754 639 1758
rect 643 1754 711 1758
rect 715 1754 799 1758
rect 803 1754 815 1758
rect 819 1754 927 1758
rect 931 1754 967 1758
rect 971 1754 1039 1758
rect 1043 1754 1143 1758
rect 1147 1754 1159 1758
rect 1163 1754 1279 1758
rect 1283 1754 1327 1758
rect 1331 1754 1399 1758
rect 1403 1754 1511 1758
rect 1515 1754 1519 1758
rect 1523 1754 1639 1758
rect 1643 1754 1703 1758
rect 1707 1754 2007 1758
rect 2011 1754 2031 1758
rect 103 1753 2031 1754
rect 2037 1753 2038 1759
rect 2018 1705 2019 1711
rect 2025 1710 3967 1711
rect 2025 1706 2047 1710
rect 2051 1706 2071 1710
rect 2075 1706 2183 1710
rect 2187 1706 2223 1710
rect 2227 1706 2327 1710
rect 2331 1706 2439 1710
rect 2443 1706 2487 1710
rect 2491 1706 2559 1710
rect 2563 1706 2655 1710
rect 2659 1706 2687 1710
rect 2691 1706 2823 1710
rect 2827 1706 2831 1710
rect 2835 1706 2967 1710
rect 2971 1706 3023 1710
rect 3027 1706 3127 1710
rect 3131 1706 3223 1710
rect 3227 1706 3303 1710
rect 3307 1706 3431 1710
rect 3435 1706 3487 1710
rect 3491 1706 3647 1710
rect 3651 1706 3671 1710
rect 3675 1706 3839 1710
rect 3843 1706 3943 1710
rect 3947 1706 3967 1710
rect 2025 1705 3967 1706
rect 3973 1705 3974 1711
rect 84 1673 85 1679
rect 91 1678 2019 1679
rect 91 1674 111 1678
rect 115 1674 135 1678
rect 139 1674 247 1678
rect 251 1674 367 1678
rect 371 1674 399 1678
rect 403 1674 495 1678
rect 499 1674 567 1678
rect 571 1674 639 1678
rect 643 1674 743 1678
rect 747 1674 799 1678
rect 803 1674 935 1678
rect 939 1674 967 1678
rect 971 1674 1135 1678
rect 1139 1674 1143 1678
rect 1147 1674 1327 1678
rect 1331 1674 1343 1678
rect 1347 1674 1511 1678
rect 1515 1674 1551 1678
rect 1555 1674 1703 1678
rect 1707 1674 1767 1678
rect 1771 1674 2007 1678
rect 2011 1674 2019 1678
rect 91 1673 2019 1674
rect 2025 1673 2026 1679
rect 2030 1625 2031 1631
rect 2037 1630 3979 1631
rect 2037 1626 2047 1630
rect 2051 1626 2223 1630
rect 2227 1626 2327 1630
rect 2331 1626 2391 1630
rect 2395 1626 2439 1630
rect 2443 1626 2503 1630
rect 2507 1626 2559 1630
rect 2563 1626 2615 1630
rect 2619 1626 2687 1630
rect 2691 1626 2735 1630
rect 2739 1626 2823 1630
rect 2827 1626 2855 1630
rect 2859 1626 2967 1630
rect 2971 1626 2975 1630
rect 2979 1626 3095 1630
rect 3099 1626 3127 1630
rect 3131 1626 3215 1630
rect 3219 1626 3303 1630
rect 3307 1626 3335 1630
rect 3339 1626 3455 1630
rect 3459 1626 3487 1630
rect 3491 1626 3671 1630
rect 3675 1626 3839 1630
rect 3843 1626 3943 1630
rect 3947 1626 3979 1630
rect 2037 1625 3979 1626
rect 3985 1625 3986 1631
rect 96 1593 97 1599
rect 103 1598 2031 1599
rect 103 1594 111 1598
rect 115 1594 135 1598
rect 139 1594 247 1598
rect 251 1594 255 1598
rect 259 1594 399 1598
rect 403 1594 423 1598
rect 427 1594 567 1598
rect 571 1594 615 1598
rect 619 1594 743 1598
rect 747 1594 831 1598
rect 835 1594 935 1598
rect 939 1594 1063 1598
rect 1067 1594 1135 1598
rect 1139 1594 1311 1598
rect 1315 1594 1343 1598
rect 1347 1594 1551 1598
rect 1555 1594 1567 1598
rect 1571 1594 1767 1598
rect 1771 1594 1831 1598
rect 1835 1594 2007 1598
rect 2011 1594 2031 1598
rect 103 1593 2031 1594
rect 2037 1593 2038 1599
rect 2018 1549 2019 1555
rect 2025 1554 3967 1555
rect 2025 1550 2047 1554
rect 2051 1550 2391 1554
rect 2395 1550 2503 1554
rect 2507 1550 2543 1554
rect 2547 1550 2615 1554
rect 2619 1550 2671 1554
rect 2675 1550 2735 1554
rect 2739 1550 2799 1554
rect 2803 1550 2855 1554
rect 2859 1550 2935 1554
rect 2939 1550 2975 1554
rect 2979 1550 3071 1554
rect 3075 1550 3095 1554
rect 3099 1550 3207 1554
rect 3211 1550 3215 1554
rect 3219 1550 3335 1554
rect 3339 1550 3455 1554
rect 3459 1550 3463 1554
rect 3467 1550 3591 1554
rect 3595 1550 3727 1554
rect 3731 1550 3839 1554
rect 3843 1550 3943 1554
rect 3947 1550 3967 1554
rect 2025 1549 3967 1550
rect 3973 1549 3974 1555
rect 84 1513 85 1519
rect 91 1518 2019 1519
rect 91 1514 111 1518
rect 115 1514 135 1518
rect 139 1514 239 1518
rect 243 1514 255 1518
rect 259 1514 407 1518
rect 411 1514 423 1518
rect 427 1514 583 1518
rect 587 1514 615 1518
rect 619 1514 775 1518
rect 779 1514 831 1518
rect 835 1514 967 1518
rect 971 1514 1063 1518
rect 1067 1514 1159 1518
rect 1163 1514 1311 1518
rect 1315 1514 1351 1518
rect 1355 1514 1543 1518
rect 1547 1514 1567 1518
rect 1571 1514 1735 1518
rect 1739 1514 1831 1518
rect 1835 1514 1903 1518
rect 1907 1514 2007 1518
rect 2011 1514 2019 1518
rect 91 1513 2019 1514
rect 2025 1513 2026 1519
rect 2030 1461 2031 1467
rect 2037 1466 3979 1467
rect 2037 1462 2047 1466
rect 2051 1462 2519 1466
rect 2523 1462 2543 1466
rect 2547 1462 2631 1466
rect 2635 1462 2671 1466
rect 2675 1462 2759 1466
rect 2763 1462 2799 1466
rect 2803 1462 2895 1466
rect 2899 1462 2935 1466
rect 2939 1462 3031 1466
rect 3035 1462 3071 1466
rect 3075 1462 3175 1466
rect 3179 1462 3207 1466
rect 3211 1462 3311 1466
rect 3315 1462 3335 1466
rect 3339 1462 3447 1466
rect 3451 1462 3463 1466
rect 3467 1462 3583 1466
rect 3587 1462 3591 1466
rect 3595 1462 3719 1466
rect 3723 1462 3727 1466
rect 3731 1462 3839 1466
rect 3843 1462 3943 1466
rect 3947 1462 3979 1466
rect 2037 1461 3979 1462
rect 3985 1461 3986 1467
rect 96 1429 97 1435
rect 103 1434 2031 1435
rect 103 1430 111 1434
rect 115 1430 239 1434
rect 243 1430 407 1434
rect 411 1430 463 1434
rect 467 1430 583 1434
rect 587 1430 711 1434
rect 715 1430 775 1434
rect 779 1430 855 1434
rect 859 1430 967 1434
rect 971 1430 1007 1434
rect 1011 1430 1159 1434
rect 1163 1430 1167 1434
rect 1171 1430 1335 1434
rect 1339 1430 1351 1434
rect 1355 1430 1511 1434
rect 1515 1430 1543 1434
rect 1547 1430 1687 1434
rect 1691 1430 1735 1434
rect 1739 1430 1871 1434
rect 1875 1430 1903 1434
rect 1907 1430 2007 1434
rect 2011 1430 2031 1434
rect 103 1429 2031 1430
rect 2037 1429 2038 1435
rect 2018 1385 2019 1391
rect 2025 1390 3967 1391
rect 2025 1386 2047 1390
rect 2051 1386 2399 1390
rect 2403 1386 2519 1390
rect 2523 1386 2535 1390
rect 2539 1386 2631 1390
rect 2635 1386 2679 1390
rect 2683 1386 2759 1390
rect 2763 1386 2823 1390
rect 2827 1386 2895 1390
rect 2899 1386 2967 1390
rect 2971 1386 3031 1390
rect 3035 1386 3111 1390
rect 3115 1386 3175 1390
rect 3179 1386 3255 1390
rect 3259 1386 3311 1390
rect 3315 1386 3407 1390
rect 3411 1386 3447 1390
rect 3451 1386 3559 1390
rect 3563 1386 3583 1390
rect 3587 1386 3711 1390
rect 3715 1386 3719 1390
rect 3723 1386 3839 1390
rect 3843 1386 3943 1390
rect 3947 1386 3967 1390
rect 2025 1385 3967 1386
rect 3973 1385 3974 1391
rect 84 1353 85 1359
rect 91 1358 2019 1359
rect 91 1354 111 1358
rect 115 1354 463 1358
rect 467 1354 583 1358
rect 587 1354 655 1358
rect 659 1354 711 1358
rect 715 1354 767 1358
rect 771 1354 855 1358
rect 859 1354 887 1358
rect 891 1354 1007 1358
rect 1011 1354 1015 1358
rect 1019 1354 1143 1358
rect 1147 1354 1167 1358
rect 1171 1354 1279 1358
rect 1283 1354 1335 1358
rect 1339 1354 1415 1358
rect 1419 1354 1511 1358
rect 1515 1354 1559 1358
rect 1563 1354 1687 1358
rect 1691 1354 1703 1358
rect 1707 1354 1847 1358
rect 1851 1354 1871 1358
rect 1875 1354 2007 1358
rect 2011 1354 2019 1358
rect 91 1353 2019 1354
rect 2025 1353 2026 1359
rect 2030 1305 2031 1311
rect 2037 1310 3979 1311
rect 2037 1306 2047 1310
rect 2051 1306 2247 1310
rect 2251 1306 2375 1310
rect 2379 1306 2399 1310
rect 2403 1306 2511 1310
rect 2515 1306 2535 1310
rect 2539 1306 2647 1310
rect 2651 1306 2679 1310
rect 2683 1306 2791 1310
rect 2795 1306 2823 1310
rect 2827 1306 2943 1310
rect 2947 1306 2967 1310
rect 2971 1306 3111 1310
rect 3115 1306 3255 1310
rect 3259 1306 3287 1310
rect 3291 1306 3407 1310
rect 3411 1306 3471 1310
rect 3475 1306 3559 1310
rect 3563 1306 3663 1310
rect 3667 1306 3711 1310
rect 3715 1306 3839 1310
rect 3843 1306 3943 1310
rect 3947 1306 3979 1310
rect 2037 1305 3979 1306
rect 3985 1305 3986 1311
rect 96 1273 97 1279
rect 103 1278 2031 1279
rect 103 1274 111 1278
rect 115 1274 439 1278
rect 443 1274 551 1278
rect 555 1274 655 1278
rect 659 1274 671 1278
rect 675 1274 767 1278
rect 771 1274 799 1278
rect 803 1274 887 1278
rect 891 1274 935 1278
rect 939 1274 1015 1278
rect 1019 1274 1079 1278
rect 1083 1274 1143 1278
rect 1147 1274 1231 1278
rect 1235 1274 1279 1278
rect 1283 1274 1391 1278
rect 1395 1274 1415 1278
rect 1419 1274 1551 1278
rect 1555 1274 1559 1278
rect 1563 1274 1703 1278
rect 1707 1274 1719 1278
rect 1723 1274 1847 1278
rect 1851 1274 2007 1278
rect 2011 1274 2031 1278
rect 103 1273 2031 1274
rect 2037 1273 2038 1279
rect 2018 1225 2019 1231
rect 2025 1230 3967 1231
rect 2025 1226 2047 1230
rect 2051 1226 2071 1230
rect 2075 1226 2183 1230
rect 2187 1226 2247 1230
rect 2251 1226 2303 1230
rect 2307 1226 2375 1230
rect 2379 1226 2431 1230
rect 2435 1226 2511 1230
rect 2515 1226 2559 1230
rect 2563 1226 2647 1230
rect 2651 1226 2711 1230
rect 2715 1226 2791 1230
rect 2795 1226 2887 1230
rect 2891 1226 2943 1230
rect 2947 1226 3087 1230
rect 3091 1226 3111 1230
rect 3115 1226 3287 1230
rect 3291 1226 3311 1230
rect 3315 1226 3471 1230
rect 3475 1226 3543 1230
rect 3547 1226 3663 1230
rect 3667 1226 3783 1230
rect 3787 1226 3839 1230
rect 3843 1226 3943 1230
rect 3947 1226 3967 1230
rect 2025 1225 3967 1226
rect 3973 1225 3974 1231
rect 84 1197 85 1203
rect 91 1202 2019 1203
rect 91 1198 111 1202
rect 115 1198 167 1202
rect 171 1198 303 1202
rect 307 1198 439 1202
rect 443 1198 463 1202
rect 467 1198 551 1202
rect 555 1198 631 1202
rect 635 1198 671 1202
rect 675 1198 799 1202
rect 803 1198 807 1202
rect 811 1198 935 1202
rect 939 1198 983 1202
rect 987 1198 1079 1202
rect 1083 1198 1159 1202
rect 1163 1198 1231 1202
rect 1235 1198 1335 1202
rect 1339 1198 1391 1202
rect 1395 1198 1511 1202
rect 1515 1198 1551 1202
rect 1555 1198 1695 1202
rect 1699 1198 1719 1202
rect 1723 1198 2007 1202
rect 2011 1198 2019 1202
rect 91 1197 2019 1198
rect 2025 1197 2026 1203
rect 2030 1145 2031 1151
rect 2037 1150 3979 1151
rect 2037 1146 2047 1150
rect 2051 1146 2071 1150
rect 2075 1146 2183 1150
rect 2187 1146 2199 1150
rect 2203 1146 2303 1150
rect 2307 1146 2351 1150
rect 2355 1146 2431 1150
rect 2435 1146 2511 1150
rect 2515 1146 2559 1150
rect 2563 1146 2679 1150
rect 2683 1146 2711 1150
rect 2715 1146 2871 1150
rect 2875 1146 2887 1150
rect 2891 1146 3087 1150
rect 3091 1146 3311 1150
rect 3315 1146 3319 1150
rect 3323 1146 3543 1150
rect 3547 1146 3559 1150
rect 3563 1146 3783 1150
rect 3787 1146 3807 1150
rect 3811 1146 3943 1150
rect 3947 1146 3979 1150
rect 2037 1145 3979 1146
rect 3985 1145 3986 1151
rect 96 1117 97 1123
rect 103 1122 2031 1123
rect 103 1118 111 1122
rect 115 1118 135 1122
rect 139 1118 167 1122
rect 171 1118 239 1122
rect 243 1118 303 1122
rect 307 1118 375 1122
rect 379 1118 463 1122
rect 467 1118 527 1122
rect 531 1118 631 1122
rect 635 1118 695 1122
rect 699 1118 807 1122
rect 811 1118 863 1122
rect 867 1118 983 1122
rect 987 1118 1039 1122
rect 1043 1118 1159 1122
rect 1163 1118 1215 1122
rect 1219 1118 1335 1122
rect 1339 1118 1391 1122
rect 1395 1118 1511 1122
rect 1515 1118 1567 1122
rect 1571 1118 1695 1122
rect 1699 1118 1743 1122
rect 1747 1118 1903 1122
rect 1907 1118 2007 1122
rect 2011 1118 2031 1122
rect 103 1117 2031 1118
rect 2037 1117 2038 1123
rect 2018 1057 2019 1063
rect 2025 1062 3967 1063
rect 2025 1058 2047 1062
rect 2051 1058 2071 1062
rect 2075 1058 2199 1062
rect 2203 1058 2263 1062
rect 2267 1058 2351 1062
rect 2355 1058 2487 1062
rect 2491 1058 2511 1062
rect 2515 1058 2679 1062
rect 2683 1058 2703 1062
rect 2707 1058 2871 1062
rect 2875 1058 2919 1062
rect 2923 1058 3087 1062
rect 3091 1058 3119 1062
rect 3123 1058 3311 1062
rect 3315 1058 3319 1062
rect 3323 1058 3495 1062
rect 3499 1058 3559 1062
rect 3563 1058 3679 1062
rect 3683 1058 3807 1062
rect 3811 1058 3839 1062
rect 3843 1058 3943 1062
rect 3947 1058 3967 1062
rect 2025 1057 3967 1058
rect 3973 1057 3974 1063
rect 84 1041 85 1047
rect 91 1046 2019 1047
rect 91 1042 111 1046
rect 115 1042 135 1046
rect 139 1042 239 1046
rect 243 1042 287 1046
rect 291 1042 375 1046
rect 379 1042 471 1046
rect 475 1042 527 1046
rect 531 1042 655 1046
rect 659 1042 695 1046
rect 699 1042 839 1046
rect 843 1042 863 1046
rect 867 1042 1015 1046
rect 1019 1042 1039 1046
rect 1043 1042 1199 1046
rect 1203 1042 1215 1046
rect 1219 1042 1383 1046
rect 1387 1042 1391 1046
rect 1395 1042 1567 1046
rect 1571 1042 1743 1046
rect 1747 1042 1903 1046
rect 1907 1042 2007 1046
rect 2011 1042 2019 1046
rect 91 1041 2019 1042
rect 2025 1041 2026 1047
rect 2030 977 2031 983
rect 2037 982 3979 983
rect 2037 978 2047 982
rect 2051 978 2071 982
rect 2075 978 2263 982
rect 2267 978 2303 982
rect 2307 978 2455 982
rect 2459 978 2487 982
rect 2491 978 2615 982
rect 2619 978 2703 982
rect 2707 978 2783 982
rect 2787 978 2919 982
rect 2923 978 2951 982
rect 2955 978 3111 982
rect 3115 978 3119 982
rect 3123 978 3263 982
rect 3267 978 3311 982
rect 3315 978 3415 982
rect 3419 978 3495 982
rect 3499 978 3559 982
rect 3563 978 3679 982
rect 3683 978 3711 982
rect 3715 978 3839 982
rect 3843 978 3943 982
rect 3947 978 3979 982
rect 2037 977 3979 978
rect 3985 977 3986 983
rect 96 961 97 967
rect 103 966 2031 967
rect 103 962 111 966
rect 115 962 135 966
rect 139 962 287 966
rect 291 962 295 966
rect 299 962 471 966
rect 475 962 639 966
rect 643 962 655 966
rect 659 962 799 966
rect 803 962 839 966
rect 843 962 951 966
rect 955 962 1015 966
rect 1019 962 1087 966
rect 1091 962 1199 966
rect 1203 962 1223 966
rect 1227 962 1359 966
rect 1363 962 1383 966
rect 1387 962 1495 966
rect 1499 962 1567 966
rect 1571 962 2007 966
rect 2011 962 2031 966
rect 103 961 2031 962
rect 2037 961 2038 967
rect 2018 897 2019 903
rect 2025 902 3967 903
rect 2025 898 2047 902
rect 2051 898 2303 902
rect 2307 898 2455 902
rect 2459 898 2559 902
rect 2563 898 2615 902
rect 2619 898 2679 902
rect 2683 898 2783 902
rect 2787 898 2807 902
rect 2811 898 2943 902
rect 2947 898 2951 902
rect 2955 898 3079 902
rect 3083 898 3111 902
rect 3115 898 3207 902
rect 3211 898 3263 902
rect 3267 898 3335 902
rect 3339 898 3415 902
rect 3419 898 3463 902
rect 3467 898 3559 902
rect 3563 898 3591 902
rect 3595 898 3711 902
rect 3715 898 3727 902
rect 3731 898 3839 902
rect 3843 898 3943 902
rect 3947 898 3967 902
rect 2025 897 3967 898
rect 3973 897 3974 903
rect 84 885 85 891
rect 91 890 2019 891
rect 91 886 111 890
rect 115 886 135 890
rect 139 886 159 890
rect 163 886 295 890
rect 299 886 319 890
rect 323 886 471 890
rect 475 886 615 890
rect 619 886 639 890
rect 643 886 751 890
rect 755 886 799 890
rect 803 886 879 890
rect 883 886 951 890
rect 955 886 999 890
rect 1003 886 1087 890
rect 1091 886 1111 890
rect 1115 886 1223 890
rect 1227 886 1231 890
rect 1235 886 1351 890
rect 1355 886 1359 890
rect 1363 886 1495 890
rect 1499 886 2007 890
rect 2011 886 2019 890
rect 91 885 2019 886
rect 2025 885 2026 891
rect 2030 817 2031 823
rect 2037 822 3979 823
rect 2037 818 2047 822
rect 2051 818 2335 822
rect 2339 818 2471 822
rect 2475 818 2559 822
rect 2563 818 2615 822
rect 2619 818 2679 822
rect 2683 818 2767 822
rect 2771 818 2807 822
rect 2811 818 2919 822
rect 2923 818 2943 822
rect 2947 818 3079 822
rect 3083 818 3207 822
rect 3211 818 3239 822
rect 3243 818 3335 822
rect 3339 818 3391 822
rect 3395 818 3463 822
rect 3467 818 3543 822
rect 3547 818 3591 822
rect 3595 818 3703 822
rect 3707 818 3727 822
rect 3731 818 3839 822
rect 3843 818 3943 822
rect 3947 818 3979 822
rect 2037 817 3979 818
rect 3985 817 3986 823
rect 2030 815 2038 817
rect 96 809 97 815
rect 103 814 2031 815
rect 103 810 111 814
rect 115 810 159 814
rect 163 810 223 814
rect 227 810 319 814
rect 323 810 383 814
rect 387 810 471 814
rect 475 810 535 814
rect 539 810 615 814
rect 619 810 679 814
rect 683 810 751 814
rect 755 810 815 814
rect 819 810 879 814
rect 883 810 951 814
rect 955 810 999 814
rect 1003 810 1079 814
rect 1083 810 1111 814
rect 1115 810 1199 814
rect 1203 810 1231 814
rect 1235 810 1327 814
rect 1331 810 1351 814
rect 1355 810 1455 814
rect 1459 810 2007 814
rect 2011 810 2031 814
rect 103 809 2031 810
rect 2037 809 2038 815
rect 2018 737 2019 743
rect 2025 742 3967 743
rect 2025 738 2047 742
rect 2051 738 2071 742
rect 2075 738 2183 742
rect 2187 738 2335 742
rect 2339 738 2471 742
rect 2475 738 2487 742
rect 2491 738 2615 742
rect 2619 738 2639 742
rect 2643 738 2767 742
rect 2771 738 2807 742
rect 2811 738 2919 742
rect 2923 738 2983 742
rect 2987 738 3079 742
rect 3083 738 3167 742
rect 3171 738 3239 742
rect 3243 738 3367 742
rect 3371 738 3391 742
rect 3395 738 3543 742
rect 3547 738 3575 742
rect 3579 738 3703 742
rect 3707 738 3783 742
rect 3787 738 3839 742
rect 3843 738 3943 742
rect 3947 738 3967 742
rect 2025 737 3967 738
rect 3973 737 3974 743
rect 2018 735 2026 737
rect 84 729 85 735
rect 91 734 2019 735
rect 91 730 111 734
rect 115 730 223 734
rect 227 730 311 734
rect 315 730 383 734
rect 387 730 471 734
rect 475 730 535 734
rect 539 730 639 734
rect 643 730 679 734
rect 683 730 807 734
rect 811 730 815 734
rect 819 730 951 734
rect 955 730 975 734
rect 979 730 1079 734
rect 1083 730 1135 734
rect 1139 730 1199 734
rect 1203 730 1295 734
rect 1299 730 1327 734
rect 1331 730 1455 734
rect 1459 730 1607 734
rect 1611 730 1767 734
rect 1771 730 1903 734
rect 1907 730 2007 734
rect 2011 730 2019 734
rect 91 729 2019 730
rect 2025 729 2026 735
rect 96 653 97 659
rect 103 658 2031 659
rect 103 654 111 658
rect 115 654 295 658
rect 299 654 311 658
rect 315 654 447 658
rect 451 654 471 658
rect 475 654 615 658
rect 619 654 639 658
rect 643 654 783 658
rect 787 654 807 658
rect 811 654 951 658
rect 955 654 975 658
rect 979 654 1111 658
rect 1115 654 1135 658
rect 1139 654 1263 658
rect 1267 654 1295 658
rect 1299 654 1399 658
rect 1403 654 1455 658
rect 1459 654 1535 658
rect 1539 654 1607 658
rect 1611 654 1663 658
rect 1667 654 1767 658
rect 1771 654 1791 658
rect 1795 654 1903 658
rect 1907 654 2007 658
rect 2011 654 2031 658
rect 103 653 2031 654
rect 2037 655 2038 659
rect 2037 654 3986 655
rect 2037 653 2047 654
rect 2030 650 2047 653
rect 2051 650 2071 654
rect 2075 650 2183 654
rect 2187 650 2239 654
rect 2243 650 2335 654
rect 2339 650 2423 654
rect 2427 650 2487 654
rect 2491 650 2623 654
rect 2627 650 2639 654
rect 2643 650 2807 654
rect 2811 650 2839 654
rect 2843 650 2983 654
rect 2987 650 3071 654
rect 3075 650 3167 654
rect 3171 650 3319 654
rect 3323 650 3367 654
rect 3371 650 3575 654
rect 3579 650 3783 654
rect 3787 650 3839 654
rect 3843 650 3943 654
rect 3947 650 3986 654
rect 2030 649 3986 650
rect 84 573 85 579
rect 91 578 2019 579
rect 91 574 111 578
rect 115 574 239 578
rect 243 574 295 578
rect 299 574 415 578
rect 419 574 447 578
rect 451 574 607 578
rect 611 574 615 578
rect 619 574 783 578
rect 787 574 799 578
rect 803 574 951 578
rect 955 574 991 578
rect 995 574 1111 578
rect 1115 574 1175 578
rect 1179 574 1263 578
rect 1267 574 1351 578
rect 1355 574 1399 578
rect 1403 574 1519 578
rect 1523 574 1535 578
rect 1539 574 1663 578
rect 1667 574 1687 578
rect 1691 574 1791 578
rect 1795 574 1863 578
rect 1867 574 1903 578
rect 1907 574 2007 578
rect 2011 574 2019 578
rect 91 573 2019 574
rect 2025 578 3974 579
rect 2025 574 2047 578
rect 2051 574 2071 578
rect 2075 574 2191 578
rect 2195 574 2239 578
rect 2243 574 2287 578
rect 2291 574 2383 578
rect 2387 574 2423 578
rect 2427 574 2479 578
rect 2483 574 2583 578
rect 2587 574 2623 578
rect 2627 574 2711 578
rect 2715 574 2839 578
rect 2843 574 2871 578
rect 2875 574 3071 578
rect 3075 574 3303 578
rect 3307 574 3319 578
rect 3323 574 3551 578
rect 3555 574 3575 578
rect 3579 574 3807 578
rect 3811 574 3839 578
rect 3843 574 3943 578
rect 3947 574 3974 578
rect 2025 573 3974 574
rect 96 497 97 503
rect 103 502 2031 503
rect 103 498 111 502
rect 115 498 135 502
rect 139 498 239 502
rect 243 498 287 502
rect 291 498 415 502
rect 419 498 463 502
rect 467 498 607 502
rect 611 498 639 502
rect 643 498 799 502
rect 803 498 807 502
rect 811 498 967 502
rect 971 498 991 502
rect 995 498 1119 502
rect 1123 498 1175 502
rect 1179 498 1271 502
rect 1275 498 1351 502
rect 1355 498 1415 502
rect 1419 498 1519 502
rect 1523 498 1567 502
rect 1571 498 1687 502
rect 1691 498 1863 502
rect 1867 498 2007 502
rect 2011 498 2031 502
rect 103 497 2031 498
rect 2037 502 3986 503
rect 2037 498 2047 502
rect 2051 498 2191 502
rect 2195 498 2287 502
rect 2291 498 2383 502
rect 2387 498 2431 502
rect 2435 498 2479 502
rect 2483 498 2527 502
rect 2531 498 2583 502
rect 2587 498 2623 502
rect 2627 498 2711 502
rect 2715 498 2727 502
rect 2731 498 2847 502
rect 2851 498 2871 502
rect 2875 498 2999 502
rect 3003 498 3071 502
rect 3075 498 3175 502
rect 3179 498 3303 502
rect 3307 498 3375 502
rect 3379 498 3551 502
rect 3555 498 3591 502
rect 3595 498 3807 502
rect 3811 498 3943 502
rect 3947 498 3986 502
rect 2037 497 3986 498
rect 2018 426 3974 427
rect 2018 423 2047 426
rect 84 417 85 423
rect 91 422 2019 423
rect 91 418 111 422
rect 115 418 135 422
rect 139 418 279 422
rect 283 418 287 422
rect 291 418 439 422
rect 443 418 463 422
rect 467 418 583 422
rect 587 418 639 422
rect 643 418 719 422
rect 723 418 807 422
rect 811 418 847 422
rect 851 418 967 422
rect 971 418 1087 422
rect 1091 418 1119 422
rect 1123 418 1207 422
rect 1211 418 1271 422
rect 1275 418 1327 422
rect 1331 418 1415 422
rect 1419 418 1567 422
rect 1571 418 2007 422
rect 2011 418 2019 422
rect 91 417 2019 418
rect 2025 422 2047 423
rect 2051 422 2431 426
rect 2435 422 2527 426
rect 2531 422 2623 426
rect 2627 422 2719 426
rect 2723 422 2727 426
rect 2731 422 2815 426
rect 2819 422 2847 426
rect 2851 422 2927 426
rect 2931 422 2999 426
rect 3003 422 3063 426
rect 3067 422 3175 426
rect 3179 422 3223 426
rect 3227 422 3375 426
rect 3379 422 3399 426
rect 3403 422 3591 426
rect 3595 422 3783 426
rect 3787 422 3807 426
rect 3811 422 3943 426
rect 3947 422 3974 426
rect 2025 421 3974 422
rect 2025 417 2026 421
rect 96 341 97 347
rect 103 346 2031 347
rect 103 342 111 346
rect 115 342 135 346
rect 139 342 143 346
rect 147 342 279 346
rect 283 342 319 346
rect 323 342 439 346
rect 443 342 479 346
rect 483 342 583 346
rect 587 342 631 346
rect 635 342 719 346
rect 723 342 775 346
rect 779 342 847 346
rect 851 342 903 346
rect 907 342 967 346
rect 971 342 1031 346
rect 1035 342 1087 346
rect 1091 342 1151 346
rect 1155 342 1207 346
rect 1211 342 1271 346
rect 1275 342 1327 346
rect 1331 342 1391 346
rect 1395 342 2007 346
rect 2011 342 2031 346
rect 103 341 2031 342
rect 2037 346 3986 347
rect 2037 342 2047 346
rect 2051 342 2191 346
rect 2195 342 2327 346
rect 2331 342 2431 346
rect 2435 342 2471 346
rect 2475 342 2527 346
rect 2531 342 2623 346
rect 2627 342 2719 346
rect 2723 342 2783 346
rect 2787 342 2815 346
rect 2819 342 2927 346
rect 2931 342 2951 346
rect 2955 342 3063 346
rect 3067 342 3119 346
rect 3123 342 3223 346
rect 3227 342 3295 346
rect 3299 342 3399 346
rect 3403 342 3471 346
rect 3475 342 3591 346
rect 3595 342 3655 346
rect 3659 342 3783 346
rect 3787 342 3839 346
rect 3843 342 3943 346
rect 3947 342 3986 346
rect 2037 341 3986 342
rect 2018 270 3974 271
rect 2018 267 2047 270
rect 84 261 85 267
rect 91 266 2019 267
rect 91 262 111 266
rect 115 262 143 266
rect 147 262 223 266
rect 227 262 319 266
rect 323 262 391 266
rect 395 262 479 266
rect 483 262 559 266
rect 563 262 631 266
rect 635 262 735 266
rect 739 262 775 266
rect 779 262 903 266
rect 907 262 1031 266
rect 1035 262 1063 266
rect 1067 262 1151 266
rect 1155 262 1215 266
rect 1219 262 1271 266
rect 1275 262 1359 266
rect 1363 262 1391 266
rect 1395 262 1511 266
rect 1515 262 1663 266
rect 1667 262 2007 266
rect 2011 262 2019 266
rect 91 261 2019 262
rect 2025 266 2047 267
rect 2051 266 2071 270
rect 2075 266 2191 270
rect 2195 266 2215 270
rect 2219 266 2327 270
rect 2331 266 2399 270
rect 2403 266 2471 270
rect 2475 266 2591 270
rect 2595 266 2623 270
rect 2627 266 2783 270
rect 2787 266 2791 270
rect 2795 266 2951 270
rect 2955 266 2983 270
rect 2987 266 3119 270
rect 3123 266 3167 270
rect 3171 266 3295 270
rect 3299 266 3343 270
rect 3347 266 3471 270
rect 3475 266 3511 270
rect 3515 266 3655 270
rect 3659 266 3687 270
rect 3691 266 3839 270
rect 3843 266 3943 270
rect 3947 266 3974 270
rect 2025 265 3974 266
rect 2025 261 2026 265
rect 2030 165 2031 171
rect 2037 170 3979 171
rect 2037 166 2047 170
rect 2051 166 2071 170
rect 2075 166 2191 170
rect 2195 166 2215 170
rect 2219 166 2343 170
rect 2347 166 2399 170
rect 2403 166 2495 170
rect 2499 166 2591 170
rect 2595 166 2647 170
rect 2651 166 2791 170
rect 2795 166 2799 170
rect 2803 166 2943 170
rect 2947 166 2983 170
rect 2987 166 3071 170
rect 3075 166 3167 170
rect 3171 166 3191 170
rect 3195 166 3311 170
rect 3315 166 3343 170
rect 3347 166 3423 170
rect 3427 166 3511 170
rect 3515 166 3527 170
rect 3531 166 3639 170
rect 3643 166 3687 170
rect 3691 166 3743 170
rect 3747 166 3839 170
rect 3843 166 3943 170
rect 3947 166 3979 170
rect 2037 165 3979 166
rect 3985 165 3986 171
rect 96 153 97 159
rect 103 158 2031 159
rect 103 154 111 158
rect 115 154 151 158
rect 155 154 223 158
rect 227 154 247 158
rect 251 154 343 158
rect 347 154 391 158
rect 395 154 439 158
rect 443 154 535 158
rect 539 154 559 158
rect 563 154 631 158
rect 635 154 727 158
rect 731 154 735 158
rect 739 154 823 158
rect 827 154 903 158
rect 907 154 919 158
rect 923 154 1015 158
rect 1019 154 1063 158
rect 1067 154 1111 158
rect 1115 154 1207 158
rect 1211 154 1215 158
rect 1219 154 1303 158
rect 1307 154 1359 158
rect 1363 154 1407 158
rect 1411 154 1511 158
rect 1515 154 1615 158
rect 1619 154 1663 158
rect 1667 154 1711 158
rect 1715 154 1807 158
rect 1811 154 1903 158
rect 1907 154 2007 158
rect 2011 154 2031 158
rect 103 153 2031 154
rect 2037 153 2038 159
rect 2018 89 2019 95
rect 2025 94 3967 95
rect 2025 90 2047 94
rect 2051 90 2071 94
rect 2075 90 2191 94
rect 2195 90 2343 94
rect 2347 90 2495 94
rect 2499 90 2647 94
rect 2651 90 2799 94
rect 2803 90 2943 94
rect 2947 90 3071 94
rect 3075 90 3191 94
rect 3195 90 3311 94
rect 3315 90 3423 94
rect 3427 90 3527 94
rect 3531 90 3639 94
rect 3643 90 3743 94
rect 3747 90 3839 94
rect 3843 90 3943 94
rect 3947 90 3967 94
rect 2025 89 3967 90
rect 3973 89 3974 95
rect 84 77 85 83
rect 91 82 2019 83
rect 91 78 111 82
rect 115 78 151 82
rect 155 78 247 82
rect 251 78 343 82
rect 347 78 439 82
rect 443 78 535 82
rect 539 78 631 82
rect 635 78 727 82
rect 731 78 823 82
rect 827 78 919 82
rect 923 78 1015 82
rect 1019 78 1111 82
rect 1115 78 1207 82
rect 1211 78 1303 82
rect 1307 78 1407 82
rect 1411 78 1511 82
rect 1515 78 1615 82
rect 1619 78 1711 82
rect 1715 78 1807 82
rect 1811 78 1903 82
rect 1907 78 2007 82
rect 2011 78 2019 82
rect 91 77 2019 78
rect 2025 77 2026 83
<< m5c >>
rect 2019 4017 2025 4023
rect 3967 4017 3973 4023
rect 85 3997 91 4003
rect 2019 3997 2025 4003
rect 2031 3941 2037 3947
rect 3979 3941 3985 3947
rect 97 3921 103 3927
rect 2031 3921 2037 3927
rect 2019 3865 2025 3871
rect 3967 3865 3973 3871
rect 85 3837 91 3843
rect 2019 3837 2025 3843
rect 2031 3773 2037 3779
rect 3979 3773 3985 3779
rect 97 3761 103 3767
rect 2031 3761 2037 3767
rect 2019 3685 2025 3691
rect 3967 3685 3973 3691
rect 85 3677 91 3683
rect 2019 3677 2025 3683
rect 2031 3605 2037 3611
rect 3979 3605 3985 3611
rect 97 3597 103 3603
rect 2031 3597 2037 3603
rect 2019 3525 2025 3531
rect 3967 3525 3973 3531
rect 85 3513 91 3519
rect 2019 3513 2025 3519
rect 2031 3449 2037 3455
rect 3979 3449 3985 3455
rect 97 3417 103 3423
rect 2031 3417 2037 3423
rect 2019 3361 2025 3367
rect 3967 3361 3973 3367
rect 85 3329 91 3335
rect 2019 3329 2025 3335
rect 2031 3281 2037 3287
rect 3979 3281 3985 3287
rect 97 3249 103 3255
rect 2031 3249 2037 3255
rect 2019 3193 2025 3199
rect 3967 3193 3973 3199
rect 85 3165 91 3171
rect 2019 3165 2025 3171
rect 2031 3113 2037 3119
rect 3979 3113 3985 3119
rect 97 3089 103 3095
rect 2031 3089 2037 3095
rect 2019 3029 2025 3035
rect 3967 3029 3973 3035
rect 85 2989 91 2995
rect 2019 2989 2025 2995
rect 2031 2949 2037 2955
rect 3979 2949 3985 2955
rect 97 2913 103 2919
rect 2031 2913 2037 2919
rect 2019 2865 2025 2871
rect 3967 2865 3973 2871
rect 85 2833 91 2839
rect 2019 2833 2025 2839
rect 2031 2789 2037 2795
rect 3979 2789 3985 2795
rect 97 2749 103 2755
rect 2031 2749 2037 2755
rect 2019 2693 2025 2699
rect 3967 2693 3973 2699
rect 85 2673 91 2679
rect 2019 2673 2025 2679
rect 2031 2609 2037 2615
rect 3979 2609 3985 2615
rect 97 2581 103 2587
rect 2031 2581 2037 2587
rect 2019 2529 2025 2535
rect 3967 2529 3973 2535
rect 85 2501 91 2507
rect 2019 2501 2025 2507
rect 2031 2441 2037 2447
rect 3979 2441 3985 2447
rect 97 2409 103 2415
rect 2031 2409 2037 2415
rect 2019 2361 2025 2367
rect 3967 2361 3973 2367
rect 85 2329 91 2335
rect 2019 2329 2025 2335
rect 2031 2285 2037 2291
rect 3979 2285 3985 2291
rect 97 2249 103 2255
rect 2031 2249 2037 2255
rect 2019 2209 2025 2215
rect 3967 2209 3973 2215
rect 85 2165 91 2171
rect 2019 2165 2025 2171
rect 2031 2109 2037 2115
rect 3979 2109 3985 2115
rect 97 2081 103 2087
rect 2031 2081 2037 2087
rect 2019 2033 2025 2039
rect 3967 2033 3973 2039
rect 85 1989 91 1995
rect 2019 1989 2025 1995
rect 2031 1945 2037 1951
rect 3979 1945 3985 1951
rect 97 1913 103 1919
rect 2031 1913 2037 1919
rect 2019 1869 2025 1875
rect 3967 1869 3973 1875
rect 85 1829 91 1835
rect 2019 1829 2025 1835
rect 2031 1789 2037 1795
rect 3979 1789 3985 1795
rect 97 1753 103 1759
rect 2031 1753 2037 1759
rect 2019 1705 2025 1711
rect 3967 1705 3973 1711
rect 85 1673 91 1679
rect 2019 1673 2025 1679
rect 2031 1625 2037 1631
rect 3979 1625 3985 1631
rect 97 1593 103 1599
rect 2031 1593 2037 1599
rect 2019 1549 2025 1555
rect 3967 1549 3973 1555
rect 85 1513 91 1519
rect 2019 1513 2025 1519
rect 2031 1461 2037 1467
rect 3979 1461 3985 1467
rect 97 1429 103 1435
rect 2031 1429 2037 1435
rect 2019 1385 2025 1391
rect 3967 1385 3973 1391
rect 85 1353 91 1359
rect 2019 1353 2025 1359
rect 2031 1305 2037 1311
rect 3979 1305 3985 1311
rect 97 1273 103 1279
rect 2031 1273 2037 1279
rect 2019 1225 2025 1231
rect 3967 1225 3973 1231
rect 85 1197 91 1203
rect 2019 1197 2025 1203
rect 2031 1145 2037 1151
rect 3979 1145 3985 1151
rect 97 1117 103 1123
rect 2031 1117 2037 1123
rect 2019 1057 2025 1063
rect 3967 1057 3973 1063
rect 85 1041 91 1047
rect 2019 1041 2025 1047
rect 2031 977 2037 983
rect 3979 977 3985 983
rect 97 961 103 967
rect 2031 961 2037 967
rect 2019 897 2025 903
rect 3967 897 3973 903
rect 85 885 91 891
rect 2019 885 2025 891
rect 2031 817 2037 823
rect 3979 817 3985 823
rect 97 809 103 815
rect 2031 809 2037 815
rect 2019 737 2025 743
rect 3967 737 3973 743
rect 85 729 91 735
rect 2019 729 2025 735
rect 97 653 103 659
rect 2031 653 2037 659
rect 85 573 91 579
rect 2019 573 2025 579
rect 97 497 103 503
rect 2031 497 2037 503
rect 85 417 91 423
rect 2019 417 2025 423
rect 97 341 103 347
rect 2031 341 2037 347
rect 85 261 91 267
rect 2019 261 2025 267
rect 2031 165 2037 171
rect 3979 165 3985 171
rect 97 153 103 159
rect 2031 153 2037 159
rect 2019 89 2025 95
rect 3967 89 3973 95
rect 85 77 91 83
rect 2019 77 2025 83
<< m5 >>
rect 84 4003 92 4032
rect 84 3997 85 4003
rect 91 3997 92 4003
rect 84 3843 92 3997
rect 84 3837 85 3843
rect 91 3837 92 3843
rect 84 3683 92 3837
rect 84 3677 85 3683
rect 91 3677 92 3683
rect 84 3519 92 3677
rect 84 3513 85 3519
rect 91 3513 92 3519
rect 84 3335 92 3513
rect 84 3329 85 3335
rect 91 3329 92 3335
rect 84 3171 92 3329
rect 84 3165 85 3171
rect 91 3165 92 3171
rect 84 2995 92 3165
rect 84 2989 85 2995
rect 91 2989 92 2995
rect 84 2839 92 2989
rect 84 2833 85 2839
rect 91 2833 92 2839
rect 84 2679 92 2833
rect 84 2673 85 2679
rect 91 2673 92 2679
rect 84 2507 92 2673
rect 84 2501 85 2507
rect 91 2501 92 2507
rect 84 2335 92 2501
rect 84 2329 85 2335
rect 91 2329 92 2335
rect 84 2171 92 2329
rect 84 2165 85 2171
rect 91 2165 92 2171
rect 84 1995 92 2165
rect 84 1989 85 1995
rect 91 1989 92 1995
rect 84 1835 92 1989
rect 84 1829 85 1835
rect 91 1829 92 1835
rect 84 1679 92 1829
rect 84 1673 85 1679
rect 91 1673 92 1679
rect 84 1519 92 1673
rect 84 1513 85 1519
rect 91 1513 92 1519
rect 84 1359 92 1513
rect 84 1353 85 1359
rect 91 1353 92 1359
rect 84 1203 92 1353
rect 84 1197 85 1203
rect 91 1197 92 1203
rect 84 1047 92 1197
rect 84 1041 85 1047
rect 91 1041 92 1047
rect 84 891 92 1041
rect 84 885 85 891
rect 91 885 92 891
rect 84 735 92 885
rect 84 729 85 735
rect 91 729 92 735
rect 84 579 92 729
rect 84 573 85 579
rect 91 573 92 579
rect 84 423 92 573
rect 84 417 85 423
rect 91 417 92 423
rect 84 267 92 417
rect 84 261 85 267
rect 91 261 92 267
rect 84 83 92 261
rect 84 77 85 83
rect 91 77 92 83
rect 84 72 92 77
rect 96 3927 104 4032
rect 96 3921 97 3927
rect 103 3921 104 3927
rect 96 3767 104 3921
rect 96 3761 97 3767
rect 103 3761 104 3767
rect 96 3603 104 3761
rect 96 3597 97 3603
rect 103 3597 104 3603
rect 96 3423 104 3597
rect 96 3417 97 3423
rect 103 3417 104 3423
rect 96 3255 104 3417
rect 96 3249 97 3255
rect 103 3249 104 3255
rect 96 3095 104 3249
rect 96 3089 97 3095
rect 103 3089 104 3095
rect 96 2919 104 3089
rect 96 2913 97 2919
rect 103 2913 104 2919
rect 96 2755 104 2913
rect 96 2749 97 2755
rect 103 2749 104 2755
rect 96 2587 104 2749
rect 96 2581 97 2587
rect 103 2581 104 2587
rect 96 2415 104 2581
rect 96 2409 97 2415
rect 103 2409 104 2415
rect 96 2255 104 2409
rect 96 2249 97 2255
rect 103 2249 104 2255
rect 96 2087 104 2249
rect 96 2081 97 2087
rect 103 2081 104 2087
rect 96 1919 104 2081
rect 96 1913 97 1919
rect 103 1913 104 1919
rect 96 1759 104 1913
rect 96 1753 97 1759
rect 103 1753 104 1759
rect 96 1599 104 1753
rect 96 1593 97 1599
rect 103 1593 104 1599
rect 96 1435 104 1593
rect 96 1429 97 1435
rect 103 1429 104 1435
rect 96 1279 104 1429
rect 96 1273 97 1279
rect 103 1273 104 1279
rect 96 1123 104 1273
rect 96 1117 97 1123
rect 103 1117 104 1123
rect 96 967 104 1117
rect 96 961 97 967
rect 103 961 104 967
rect 96 815 104 961
rect 96 809 97 815
rect 103 809 104 815
rect 96 659 104 809
rect 96 653 97 659
rect 103 653 104 659
rect 96 503 104 653
rect 96 497 97 503
rect 103 497 104 503
rect 96 347 104 497
rect 96 341 97 347
rect 103 341 104 347
rect 96 159 104 341
rect 96 153 97 159
rect 103 153 104 159
rect 96 72 104 153
rect 2018 4023 2026 4032
rect 2018 4017 2019 4023
rect 2025 4017 2026 4023
rect 2018 4003 2026 4017
rect 2018 3997 2019 4003
rect 2025 3997 2026 4003
rect 2018 3871 2026 3997
rect 2018 3865 2019 3871
rect 2025 3865 2026 3871
rect 2018 3843 2026 3865
rect 2018 3837 2019 3843
rect 2025 3837 2026 3843
rect 2018 3691 2026 3837
rect 2018 3685 2019 3691
rect 2025 3685 2026 3691
rect 2018 3683 2026 3685
rect 2018 3677 2019 3683
rect 2025 3677 2026 3683
rect 2018 3531 2026 3677
rect 2018 3525 2019 3531
rect 2025 3525 2026 3531
rect 2018 3519 2026 3525
rect 2018 3513 2019 3519
rect 2025 3513 2026 3519
rect 2018 3367 2026 3513
rect 2018 3361 2019 3367
rect 2025 3361 2026 3367
rect 2018 3335 2026 3361
rect 2018 3329 2019 3335
rect 2025 3329 2026 3335
rect 2018 3199 2026 3329
rect 2018 3193 2019 3199
rect 2025 3193 2026 3199
rect 2018 3171 2026 3193
rect 2018 3165 2019 3171
rect 2025 3165 2026 3171
rect 2018 3035 2026 3165
rect 2018 3029 2019 3035
rect 2025 3029 2026 3035
rect 2018 2995 2026 3029
rect 2018 2989 2019 2995
rect 2025 2989 2026 2995
rect 2018 2871 2026 2989
rect 2018 2865 2019 2871
rect 2025 2865 2026 2871
rect 2018 2839 2026 2865
rect 2018 2833 2019 2839
rect 2025 2833 2026 2839
rect 2018 2699 2026 2833
rect 2018 2693 2019 2699
rect 2025 2693 2026 2699
rect 2018 2679 2026 2693
rect 2018 2673 2019 2679
rect 2025 2673 2026 2679
rect 2018 2535 2026 2673
rect 2018 2529 2019 2535
rect 2025 2529 2026 2535
rect 2018 2507 2026 2529
rect 2018 2501 2019 2507
rect 2025 2501 2026 2507
rect 2018 2367 2026 2501
rect 2018 2361 2019 2367
rect 2025 2361 2026 2367
rect 2018 2335 2026 2361
rect 2018 2329 2019 2335
rect 2025 2329 2026 2335
rect 2018 2215 2026 2329
rect 2018 2209 2019 2215
rect 2025 2209 2026 2215
rect 2018 2171 2026 2209
rect 2018 2165 2019 2171
rect 2025 2165 2026 2171
rect 2018 2039 2026 2165
rect 2018 2033 2019 2039
rect 2025 2033 2026 2039
rect 2018 1995 2026 2033
rect 2018 1989 2019 1995
rect 2025 1989 2026 1995
rect 2018 1875 2026 1989
rect 2018 1869 2019 1875
rect 2025 1869 2026 1875
rect 2018 1835 2026 1869
rect 2018 1829 2019 1835
rect 2025 1829 2026 1835
rect 2018 1711 2026 1829
rect 2018 1705 2019 1711
rect 2025 1705 2026 1711
rect 2018 1679 2026 1705
rect 2018 1673 2019 1679
rect 2025 1673 2026 1679
rect 2018 1555 2026 1673
rect 2018 1549 2019 1555
rect 2025 1549 2026 1555
rect 2018 1519 2026 1549
rect 2018 1513 2019 1519
rect 2025 1513 2026 1519
rect 2018 1391 2026 1513
rect 2018 1385 2019 1391
rect 2025 1385 2026 1391
rect 2018 1359 2026 1385
rect 2018 1353 2019 1359
rect 2025 1353 2026 1359
rect 2018 1231 2026 1353
rect 2018 1225 2019 1231
rect 2025 1225 2026 1231
rect 2018 1203 2026 1225
rect 2018 1197 2019 1203
rect 2025 1197 2026 1203
rect 2018 1063 2026 1197
rect 2018 1057 2019 1063
rect 2025 1057 2026 1063
rect 2018 1047 2026 1057
rect 2018 1041 2019 1047
rect 2025 1041 2026 1047
rect 2018 903 2026 1041
rect 2018 897 2019 903
rect 2025 897 2026 903
rect 2018 891 2026 897
rect 2018 885 2019 891
rect 2025 885 2026 891
rect 2018 743 2026 885
rect 2018 737 2019 743
rect 2025 737 2026 743
rect 2018 735 2026 737
rect 2018 729 2019 735
rect 2025 729 2026 735
rect 2018 579 2026 729
rect 2018 573 2019 579
rect 2025 573 2026 579
rect 2018 423 2026 573
rect 2018 417 2019 423
rect 2025 417 2026 423
rect 2018 267 2026 417
rect 2018 261 2019 267
rect 2025 261 2026 267
rect 2018 95 2026 261
rect 2018 89 2019 95
rect 2025 89 2026 95
rect 2018 83 2026 89
rect 2018 77 2019 83
rect 2025 77 2026 83
rect 2018 72 2026 77
rect 2030 3947 2038 4032
rect 2030 3941 2031 3947
rect 2037 3941 2038 3947
rect 2030 3927 2038 3941
rect 2030 3921 2031 3927
rect 2037 3921 2038 3927
rect 2030 3779 2038 3921
rect 2030 3773 2031 3779
rect 2037 3773 2038 3779
rect 2030 3767 2038 3773
rect 2030 3761 2031 3767
rect 2037 3761 2038 3767
rect 2030 3611 2038 3761
rect 2030 3605 2031 3611
rect 2037 3605 2038 3611
rect 2030 3603 2038 3605
rect 2030 3597 2031 3603
rect 2037 3597 2038 3603
rect 2030 3455 2038 3597
rect 2030 3449 2031 3455
rect 2037 3449 2038 3455
rect 2030 3423 2038 3449
rect 2030 3417 2031 3423
rect 2037 3417 2038 3423
rect 2030 3287 2038 3417
rect 2030 3281 2031 3287
rect 2037 3281 2038 3287
rect 2030 3255 2038 3281
rect 2030 3249 2031 3255
rect 2037 3249 2038 3255
rect 2030 3119 2038 3249
rect 2030 3113 2031 3119
rect 2037 3113 2038 3119
rect 2030 3095 2038 3113
rect 2030 3089 2031 3095
rect 2037 3089 2038 3095
rect 2030 2955 2038 3089
rect 2030 2949 2031 2955
rect 2037 2949 2038 2955
rect 2030 2919 2038 2949
rect 2030 2913 2031 2919
rect 2037 2913 2038 2919
rect 2030 2795 2038 2913
rect 2030 2789 2031 2795
rect 2037 2789 2038 2795
rect 2030 2755 2038 2789
rect 2030 2749 2031 2755
rect 2037 2749 2038 2755
rect 2030 2615 2038 2749
rect 2030 2609 2031 2615
rect 2037 2609 2038 2615
rect 2030 2587 2038 2609
rect 2030 2581 2031 2587
rect 2037 2581 2038 2587
rect 2030 2447 2038 2581
rect 2030 2441 2031 2447
rect 2037 2441 2038 2447
rect 2030 2415 2038 2441
rect 2030 2409 2031 2415
rect 2037 2409 2038 2415
rect 2030 2291 2038 2409
rect 2030 2285 2031 2291
rect 2037 2285 2038 2291
rect 2030 2255 2038 2285
rect 2030 2249 2031 2255
rect 2037 2249 2038 2255
rect 2030 2115 2038 2249
rect 2030 2109 2031 2115
rect 2037 2109 2038 2115
rect 2030 2087 2038 2109
rect 2030 2081 2031 2087
rect 2037 2081 2038 2087
rect 2030 1951 2038 2081
rect 2030 1945 2031 1951
rect 2037 1945 2038 1951
rect 2030 1919 2038 1945
rect 2030 1913 2031 1919
rect 2037 1913 2038 1919
rect 2030 1795 2038 1913
rect 2030 1789 2031 1795
rect 2037 1789 2038 1795
rect 2030 1759 2038 1789
rect 2030 1753 2031 1759
rect 2037 1753 2038 1759
rect 2030 1631 2038 1753
rect 2030 1625 2031 1631
rect 2037 1625 2038 1631
rect 2030 1599 2038 1625
rect 2030 1593 2031 1599
rect 2037 1593 2038 1599
rect 2030 1467 2038 1593
rect 2030 1461 2031 1467
rect 2037 1461 2038 1467
rect 2030 1435 2038 1461
rect 2030 1429 2031 1435
rect 2037 1429 2038 1435
rect 2030 1311 2038 1429
rect 2030 1305 2031 1311
rect 2037 1305 2038 1311
rect 2030 1279 2038 1305
rect 2030 1273 2031 1279
rect 2037 1273 2038 1279
rect 2030 1151 2038 1273
rect 2030 1145 2031 1151
rect 2037 1145 2038 1151
rect 2030 1123 2038 1145
rect 2030 1117 2031 1123
rect 2037 1117 2038 1123
rect 2030 983 2038 1117
rect 2030 977 2031 983
rect 2037 977 2038 983
rect 2030 967 2038 977
rect 2030 961 2031 967
rect 2037 961 2038 967
rect 2030 823 2038 961
rect 2030 817 2031 823
rect 2037 817 2038 823
rect 2030 815 2038 817
rect 2030 809 2031 815
rect 2037 809 2038 815
rect 2030 659 2038 809
rect 2030 653 2031 659
rect 2037 653 2038 659
rect 2030 503 2038 653
rect 2030 497 2031 503
rect 2037 497 2038 503
rect 2030 347 2038 497
rect 2030 341 2031 347
rect 2037 341 2038 347
rect 2030 171 2038 341
rect 2030 165 2031 171
rect 2037 165 2038 171
rect 2030 159 2038 165
rect 2030 153 2031 159
rect 2037 153 2038 159
rect 2030 72 2038 153
rect 3966 4023 3974 4032
rect 3966 4017 3967 4023
rect 3973 4017 3974 4023
rect 3966 3871 3974 4017
rect 3966 3865 3967 3871
rect 3973 3865 3974 3871
rect 3966 3691 3974 3865
rect 3966 3685 3967 3691
rect 3973 3685 3974 3691
rect 3966 3531 3974 3685
rect 3966 3525 3967 3531
rect 3973 3525 3974 3531
rect 3966 3367 3974 3525
rect 3966 3361 3967 3367
rect 3973 3361 3974 3367
rect 3966 3199 3974 3361
rect 3966 3193 3967 3199
rect 3973 3193 3974 3199
rect 3966 3035 3974 3193
rect 3966 3029 3967 3035
rect 3973 3029 3974 3035
rect 3966 2871 3974 3029
rect 3966 2865 3967 2871
rect 3973 2865 3974 2871
rect 3966 2699 3974 2865
rect 3966 2693 3967 2699
rect 3973 2693 3974 2699
rect 3966 2535 3974 2693
rect 3966 2529 3967 2535
rect 3973 2529 3974 2535
rect 3966 2367 3974 2529
rect 3966 2361 3967 2367
rect 3973 2361 3974 2367
rect 3966 2215 3974 2361
rect 3966 2209 3967 2215
rect 3973 2209 3974 2215
rect 3966 2039 3974 2209
rect 3966 2033 3967 2039
rect 3973 2033 3974 2039
rect 3966 1875 3974 2033
rect 3966 1869 3967 1875
rect 3973 1869 3974 1875
rect 3966 1711 3974 1869
rect 3966 1705 3967 1711
rect 3973 1705 3974 1711
rect 3966 1555 3974 1705
rect 3966 1549 3967 1555
rect 3973 1549 3974 1555
rect 3966 1391 3974 1549
rect 3966 1385 3967 1391
rect 3973 1385 3974 1391
rect 3966 1231 3974 1385
rect 3966 1225 3967 1231
rect 3973 1225 3974 1231
rect 3966 1063 3974 1225
rect 3966 1057 3967 1063
rect 3973 1057 3974 1063
rect 3966 903 3974 1057
rect 3966 897 3967 903
rect 3973 897 3974 903
rect 3966 743 3974 897
rect 3966 737 3967 743
rect 3973 737 3974 743
rect 3966 95 3974 737
rect 3966 89 3967 95
rect 3973 89 3974 95
rect 3966 72 3974 89
rect 3978 3947 3986 4032
rect 3978 3941 3979 3947
rect 3985 3941 3986 3947
rect 3978 3779 3986 3941
rect 3978 3773 3979 3779
rect 3985 3773 3986 3779
rect 3978 3611 3986 3773
rect 3978 3605 3979 3611
rect 3985 3605 3986 3611
rect 3978 3455 3986 3605
rect 3978 3449 3979 3455
rect 3985 3449 3986 3455
rect 3978 3287 3986 3449
rect 3978 3281 3979 3287
rect 3985 3281 3986 3287
rect 3978 3119 3986 3281
rect 3978 3113 3979 3119
rect 3985 3113 3986 3119
rect 3978 2955 3986 3113
rect 3978 2949 3979 2955
rect 3985 2949 3986 2955
rect 3978 2795 3986 2949
rect 3978 2789 3979 2795
rect 3985 2789 3986 2795
rect 3978 2615 3986 2789
rect 3978 2609 3979 2615
rect 3985 2609 3986 2615
rect 3978 2447 3986 2609
rect 3978 2441 3979 2447
rect 3985 2441 3986 2447
rect 3978 2291 3986 2441
rect 3978 2285 3979 2291
rect 3985 2285 3986 2291
rect 3978 2115 3986 2285
rect 3978 2109 3979 2115
rect 3985 2109 3986 2115
rect 3978 1951 3986 2109
rect 3978 1945 3979 1951
rect 3985 1945 3986 1951
rect 3978 1795 3986 1945
rect 3978 1789 3979 1795
rect 3985 1789 3986 1795
rect 3978 1631 3986 1789
rect 3978 1625 3979 1631
rect 3985 1625 3986 1631
rect 3978 1467 3986 1625
rect 3978 1461 3979 1467
rect 3985 1461 3986 1467
rect 3978 1311 3986 1461
rect 3978 1305 3979 1311
rect 3985 1305 3986 1311
rect 3978 1151 3986 1305
rect 3978 1145 3979 1151
rect 3985 1145 3986 1151
rect 3978 983 3986 1145
rect 3978 977 3979 983
rect 3985 977 3986 983
rect 3978 823 3986 977
rect 3978 817 3979 823
rect 3985 817 3986 823
rect 3978 171 3986 817
rect 3978 165 3979 171
rect 3985 165 3986 171
rect 3978 72 3986 165
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__191
timestamp 1731220339
transform 1 0 3936 0 -1 3992
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220339
transform 1 0 2040 0 -1 3992
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220339
transform 1 0 3936 0 1 3896
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220339
transform 1 0 2040 0 1 3896
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220339
transform 1 0 3936 0 -1 3840
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220339
transform 1 0 2040 0 -1 3840
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220339
transform 1 0 3936 0 1 3728
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220339
transform 1 0 2040 0 1 3728
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220339
transform 1 0 3936 0 -1 3660
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220339
transform 1 0 2040 0 -1 3660
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220339
transform 1 0 3936 0 1 3560
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220339
transform 1 0 2040 0 1 3560
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220339
transform 1 0 3936 0 -1 3500
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220339
transform 1 0 2040 0 -1 3500
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220339
transform 1 0 3936 0 1 3404
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220339
transform 1 0 2040 0 1 3404
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220339
transform 1 0 3936 0 -1 3336
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220339
transform 1 0 2040 0 -1 3336
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220339
transform 1 0 3936 0 1 3236
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220339
transform 1 0 2040 0 1 3236
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220339
transform 1 0 3936 0 -1 3168
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220339
transform 1 0 2040 0 -1 3168
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220339
transform 1 0 3936 0 1 3068
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220339
transform 1 0 2040 0 1 3068
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220339
transform 1 0 3936 0 -1 3004
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220339
transform 1 0 2040 0 -1 3004
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220339
transform 1 0 3936 0 1 2904
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220339
transform 1 0 2040 0 1 2904
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220339
transform 1 0 3936 0 -1 2840
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220339
transform 1 0 2040 0 -1 2840
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220339
transform 1 0 3936 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220339
transform 1 0 2040 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220339
transform 1 0 3936 0 -1 2668
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220339
transform 1 0 2040 0 -1 2668
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220339
transform 1 0 3936 0 1 2564
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220339
transform 1 0 2040 0 1 2564
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220339
transform 1 0 3936 0 -1 2504
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220339
transform 1 0 2040 0 -1 2504
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220339
transform 1 0 3936 0 1 2396
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220339
transform 1 0 2040 0 1 2396
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220339
transform 1 0 3936 0 -1 2336
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220339
transform 1 0 2040 0 -1 2336
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220339
transform 1 0 3936 0 1 2240
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220339
transform 1 0 2040 0 1 2240
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220339
transform 1 0 3936 0 -1 2184
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220339
transform 1 0 2040 0 -1 2184
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220339
transform 1 0 3936 0 1 2064
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220339
transform 1 0 2040 0 1 2064
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220339
transform 1 0 3936 0 -1 2008
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220339
transform 1 0 2040 0 -1 2008
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220339
transform 1 0 3936 0 1 1900
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220339
transform 1 0 2040 0 1 1900
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220339
transform 1 0 3936 0 -1 1844
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220339
transform 1 0 2040 0 -1 1844
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220339
transform 1 0 3936 0 1 1744
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220339
transform 1 0 2040 0 1 1744
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220339
transform 1 0 3936 0 -1 1680
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220339
transform 1 0 2040 0 -1 1680
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220339
transform 1 0 3936 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220339
transform 1 0 2040 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220339
transform 1 0 3936 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220339
transform 1 0 2040 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220339
transform 1 0 3936 0 1 1416
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220339
transform 1 0 2040 0 1 1416
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220339
transform 1 0 3936 0 -1 1360
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220339
transform 1 0 2040 0 -1 1360
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220339
transform 1 0 3936 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220339
transform 1 0 2040 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220339
transform 1 0 3936 0 -1 1200
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220339
transform 1 0 2040 0 -1 1200
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220339
transform 1 0 3936 0 1 1100
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220339
transform 1 0 2040 0 1 1100
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220339
transform 1 0 3936 0 -1 1032
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220339
transform 1 0 2040 0 -1 1032
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220339
transform 1 0 3936 0 1 932
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220339
transform 1 0 2040 0 1 932
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220339
transform 1 0 3936 0 -1 872
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220339
transform 1 0 2040 0 -1 872
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220339
transform 1 0 3936 0 1 772
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220339
transform 1 0 2040 0 1 772
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220339
transform 1 0 3936 0 -1 712
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220339
transform 1 0 2040 0 -1 712
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220339
transform 1 0 3936 0 1 604
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220339
transform 1 0 2040 0 1 604
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220339
transform 1 0 3936 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220339
transform 1 0 2040 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220339
transform 1 0 3936 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220339
transform 1 0 2040 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220339
transform 1 0 3936 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220339
transform 1 0 2040 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220339
transform 1 0 3936 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220339
transform 1 0 2040 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220339
transform 1 0 3936 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220339
transform 1 0 2040 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220339
transform 1 0 3936 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220339
transform 1 0 2040 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220339
transform 1 0 2000 0 -1 3972
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220339
transform 1 0 104 0 -1 3972
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220339
transform 1 0 2000 0 1 3876
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220339
transform 1 0 104 0 1 3876
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220339
transform 1 0 2000 0 -1 3812
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220339
transform 1 0 104 0 -1 3812
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220339
transform 1 0 2000 0 1 3716
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220339
transform 1 0 104 0 1 3716
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220339
transform 1 0 2000 0 -1 3652
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220339
transform 1 0 104 0 -1 3652
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220339
transform 1 0 2000 0 1 3552
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220339
transform 1 0 104 0 1 3552
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220339
transform 1 0 2000 0 -1 3488
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220339
transform 1 0 104 0 -1 3488
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220339
transform 1 0 2000 0 1 3372
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220339
transform 1 0 104 0 1 3372
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220339
transform 1 0 2000 0 -1 3304
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220339
transform 1 0 104 0 -1 3304
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220339
transform 1 0 2000 0 1 3204
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220339
transform 1 0 104 0 1 3204
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220339
transform 1 0 2000 0 -1 3140
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220339
transform 1 0 104 0 -1 3140
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220339
transform 1 0 2000 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220339
transform 1 0 104 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220339
transform 1 0 2000 0 -1 2964
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220339
transform 1 0 104 0 -1 2964
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220339
transform 1 0 2000 0 1 2868
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220339
transform 1 0 104 0 1 2868
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220339
transform 1 0 2000 0 -1 2808
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220339
transform 1 0 104 0 -1 2808
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220339
transform 1 0 2000 0 1 2704
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220339
transform 1 0 104 0 1 2704
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220339
transform 1 0 2000 0 -1 2648
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220339
transform 1 0 104 0 -1 2648
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220339
transform 1 0 2000 0 1 2536
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220339
transform 1 0 104 0 1 2536
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220339
transform 1 0 2000 0 -1 2476
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220339
transform 1 0 104 0 -1 2476
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220339
transform 1 0 2000 0 1 2364
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220339
transform 1 0 104 0 1 2364
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220339
transform 1 0 2000 0 -1 2304
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220339
transform 1 0 104 0 -1 2304
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220339
transform 1 0 2000 0 1 2204
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220339
transform 1 0 104 0 1 2204
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220339
transform 1 0 2000 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220339
transform 1 0 104 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220339
transform 1 0 2000 0 1 2036
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220339
transform 1 0 104 0 1 2036
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220339
transform 1 0 2000 0 -1 1964
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220339
transform 1 0 104 0 -1 1964
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220339
transform 1 0 2000 0 1 1868
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220339
transform 1 0 104 0 1 1868
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220339
transform 1 0 2000 0 -1 1804
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220339
transform 1 0 104 0 -1 1804
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220339
transform 1 0 2000 0 1 1708
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220339
transform 1 0 104 0 1 1708
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220339
transform 1 0 2000 0 -1 1648
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220339
transform 1 0 104 0 -1 1648
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220339
transform 1 0 2000 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220339
transform 1 0 104 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220339
transform 1 0 2000 0 -1 1488
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220339
transform 1 0 104 0 -1 1488
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220339
transform 1 0 2000 0 1 1384
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220339
transform 1 0 104 0 1 1384
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220339
transform 1 0 2000 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220339
transform 1 0 104 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220339
transform 1 0 2000 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220339
transform 1 0 104 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220339
transform 1 0 2000 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220339
transform 1 0 104 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220339
transform 1 0 2000 0 1 1072
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220339
transform 1 0 104 0 1 1072
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220339
transform 1 0 2000 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220339
transform 1 0 104 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220339
transform 1 0 2000 0 1 916
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220339
transform 1 0 104 0 1 916
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220339
transform 1 0 2000 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220339
transform 1 0 104 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220339
transform 1 0 2000 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220339
transform 1 0 104 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220339
transform 1 0 2000 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220339
transform 1 0 104 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220339
transform 1 0 2000 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220339
transform 1 0 104 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220339
transform 1 0 2000 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220339
transform 1 0 104 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220339
transform 1 0 2000 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220339
transform 1 0 104 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220339
transform 1 0 2000 0 -1 392
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220339
transform 1 0 104 0 -1 392
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220339
transform 1 0 2000 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220339
transform 1 0 104 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220339
transform 1 0 2000 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220339
transform 1 0 104 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220339
transform 1 0 2000 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220339
transform 1 0 104 0 1 108
box 7 3 12 24
use _0_0cell_0_0gcelem3x0  tst_5999_6
timestamp 1731220339
transform 1 0 3736 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5998_6
timestamp 1731220339
transform 1 0 3832 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5997_6
timestamp 1731220339
transform 1 0 3832 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5996_6
timestamp 1731220339
transform 1 0 3832 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5995_6
timestamp 1731220339
transform 1 0 3800 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5994_6
timestamp 1731220339
transform 1 0 3776 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5993_6
timestamp 1731220339
transform 1 0 3648 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5992_6
timestamp 1731220339
transform 1 0 3680 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5991_6
timestamp 1731220339
transform 1 0 3504 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5990_6
timestamp 1731220339
transform 1 0 3632 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5989_6
timestamp 1731220339
transform 1 0 3520 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5988_6
timestamp 1731220339
transform 1 0 3416 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5987_6
timestamp 1731220339
transform 1 0 3304 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5986_6
timestamp 1731220339
transform 1 0 3184 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5985_6
timestamp 1731220339
transform 1 0 3064 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5984_6
timestamp 1731220339
transform 1 0 2936 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5983_6
timestamp 1731220339
transform 1 0 2792 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5982_6
timestamp 1731220339
transform 1 0 2976 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5981_6
timestamp 1731220339
transform 1 0 3160 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5980_6
timestamp 1731220339
transform 1 0 3336 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5979_6
timestamp 1731220339
transform 1 0 3464 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5978_6
timestamp 1731220339
transform 1 0 3288 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5977_6
timestamp 1731220339
transform 1 0 3112 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5976_6
timestamp 1731220339
transform 1 0 2944 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5975_6
timestamp 1731220339
transform 1 0 3584 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5974_6
timestamp 1731220339
transform 1 0 3392 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5973_6
timestamp 1731220339
transform 1 0 3216 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5972_6
timestamp 1731220339
transform 1 0 3056 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5971_6
timestamp 1731220339
transform 1 0 2920 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5970_6
timestamp 1731220339
transform 1 0 3168 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5969_6
timestamp 1731220339
transform 1 0 3368 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5968_6
timestamp 1731220339
transform 1 0 3584 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5967_6
timestamp 1731220339
transform 1 0 3544 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5966_6
timestamp 1731220339
transform 1 0 3296 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5965_6
timestamp 1731220339
transform 1 0 3064 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5964_6
timestamp 1731220339
transform 1 0 2864 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5963_6
timestamp 1731220339
transform 1 0 2704 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5962_6
timestamp 1731220339
transform 1 0 2616 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5961_6
timestamp 1731220339
transform 1 0 2832 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5960_6
timestamp 1731220339
transform 1 0 3064 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5959_6
timestamp 1731220339
transform 1 0 3568 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5958_6
timestamp 1731220339
transform 1 0 3312 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5957_6
timestamp 1731220339
transform 1 0 3160 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5956_6
timestamp 1731220339
transform 1 0 2976 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5955_6
timestamp 1731220339
transform 1 0 2800 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5954_6
timestamp 1731220339
transform 1 0 3360 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5953_6
timestamp 1731220339
transform 1 0 3568 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5952_6
timestamp 1731220339
transform 1 0 3384 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5951_6
timestamp 1731220339
transform 1 0 3232 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5950_6
timestamp 1731220339
transform 1 0 3072 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5949_6
timestamp 1731220339
transform 1 0 3200 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5948_6
timestamp 1731220339
transform 1 0 3328 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5947_6
timestamp 1731220339
transform 1 0 3456 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5946_6
timestamp 1731220339
transform 1 0 3704 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5945_6
timestamp 1731220339
transform 1 0 3720 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5944_6
timestamp 1731220339
transform 1 0 3584 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5943_6
timestamp 1731220339
transform 1 0 3536 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5942_6
timestamp 1731220339
transform 1 0 3696 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5941_6
timestamp 1731220339
transform 1 0 3776 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5940_6
timestamp 1731220339
transform 1 0 3800 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5939_6
timestamp 1731220339
transform 1 0 3832 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5938_6
timestamp 1731220339
transform 1 0 3832 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5937_6
timestamp 1731220339
transform 1 0 3832 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5936_6
timestamp 1731220339
transform 1 0 3832 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5935_6
timestamp 1731220339
transform 1 0 3832 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5934_6
timestamp 1731220339
transform 1 0 3800 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5933_6
timestamp 1731220339
transform 1 0 3776 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5932_6
timestamp 1731220339
transform 1 0 3672 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5931_6
timestamp 1731220339
transform 1 0 3488 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5930_6
timestamp 1731220339
transform 1 0 3552 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5929_6
timestamp 1731220339
transform 1 0 3408 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5928_6
timestamp 1731220339
transform 1 0 3256 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5927_6
timestamp 1731220339
transform 1 0 3104 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5926_6
timestamp 1731220339
transform 1 0 2912 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5925_6
timestamp 1731220339
transform 1 0 3112 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5924_6
timestamp 1731220339
transform 1 0 3304 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5923_6
timestamp 1731220339
transform 1 0 3552 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5922_6
timestamp 1731220339
transform 1 0 3312 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5921_6
timestamp 1731220339
transform 1 0 3080 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5920_6
timestamp 1731220339
transform 1 0 2864 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5919_6
timestamp 1731220339
transform 1 0 2672 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5918_6
timestamp 1731220339
transform 1 0 2704 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5917_6
timestamp 1731220339
transform 1 0 2880 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5916_6
timestamp 1731220339
transform 1 0 3080 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5915_6
timestamp 1731220339
transform 1 0 3304 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5914_6
timestamp 1731220339
transform 1 0 3536 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5913_6
timestamp 1731220339
transform 1 0 3656 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5912_6
timestamp 1731220339
transform 1 0 3464 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5911_6
timestamp 1731220339
transform 1 0 3280 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5910_6
timestamp 1731220339
transform 1 0 3104 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5909_6
timestamp 1731220339
transform 1 0 2936 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5908_6
timestamp 1731220339
transform 1 0 3104 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5907_6
timestamp 1731220339
transform 1 0 3248 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5906_6
timestamp 1731220339
transform 1 0 3400 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5905_6
timestamp 1731220339
transform 1 0 3704 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5904_6
timestamp 1731220339
transform 1 0 3552 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5903_6
timestamp 1731220339
transform 1 0 3440 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5902_6
timestamp 1731220339
transform 1 0 3304 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5901_6
timestamp 1731220339
transform 1 0 3576 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5900_6
timestamp 1731220339
transform 1 0 3712 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5899_6
timestamp 1731220339
transform 1 0 3584 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5898_6
timestamp 1731220339
transform 1 0 3456 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5897_6
timestamp 1731220339
transform 1 0 3328 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5896_6
timestamp 1731220339
transform 1 0 3200 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5895_6
timestamp 1731220339
transform 1 0 3448 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5894_6
timestamp 1731220339
transform 1 0 3328 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5893_6
timestamp 1731220339
transform 1 0 3208 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5892_6
timestamp 1731220339
transform 1 0 3088 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5891_6
timestamp 1731220339
transform 1 0 2968 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5890_6
timestamp 1731220339
transform 1 0 3480 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5889_6
timestamp 1731220339
transform 1 0 3296 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5888_6
timestamp 1731220339
transform 1 0 3120 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5887_6
timestamp 1731220339
transform 1 0 2960 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5886_6
timestamp 1731220339
transform 1 0 2816 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5885_6
timestamp 1731220339
transform 1 0 2824 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5884_6
timestamp 1731220339
transform 1 0 3016 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5883_6
timestamp 1731220339
transform 1 0 3216 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5882_6
timestamp 1731220339
transform 1 0 3424 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5881_6
timestamp 1731220339
transform 1 0 3448 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5880_6
timestamp 1731220339
transform 1 0 3312 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5879_6
timestamp 1731220339
transform 1 0 3176 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5878_6
timestamp 1731220339
transform 1 0 3032 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5877_6
timestamp 1731220339
transform 1 0 2880 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5876_6
timestamp 1731220339
transform 1 0 3120 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5875_6
timestamp 1731220339
transform 1 0 3352 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5874_6
timestamp 1731220339
transform 1 0 3584 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5873_6
timestamp 1731220339
transform 1 0 3576 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5872_6
timestamp 1731220339
transform 1 0 3704 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5871_6
timestamp 1731220339
transform 1 0 3640 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5870_6
timestamp 1731220339
transform 1 0 3664 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5869_6
timestamp 1731220339
transform 1 0 3720 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5868_6
timestamp 1731220339
transform 1 0 3832 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5867_6
timestamp 1731220339
transform 1 0 3832 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5866_6
timestamp 1731220339
transform 1 0 3832 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5865_6
timestamp 1731220339
transform 1 0 3832 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5864_6
timestamp 1731220339
transform 1 0 3832 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5863_6
timestamp 1731220339
transform 1 0 3832 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5862_6
timestamp 1731220339
transform 1 0 3832 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5861_6
timestamp 1731220339
transform 1 0 3824 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5860_6
timestamp 1731220339
transform 1 0 3520 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5859_6
timestamp 1731220339
transform 1 0 3832 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5858_6
timestamp 1731220339
transform 1 0 3832 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5857_6
timestamp 1731220339
transform 1 0 3736 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5856_6
timestamp 1731220339
transform 1 0 3640 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5855_6
timestamp 1731220339
transform 1 0 3544 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5854_6
timestamp 1731220339
transform 1 0 3448 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5853_6
timestamp 1731220339
transform 1 0 3352 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5852_6
timestamp 1731220339
transform 1 0 3256 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5851_6
timestamp 1731220339
transform 1 0 3160 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5850_6
timestamp 1731220339
transform 1 0 3064 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5849_6
timestamp 1731220339
transform 1 0 2968 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5848_6
timestamp 1731220339
transform 1 0 2872 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5847_6
timestamp 1731220339
transform 1 0 3464 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5846_6
timestamp 1731220339
transform 1 0 3312 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5845_6
timestamp 1731220339
transform 1 0 3168 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5844_6
timestamp 1731220339
transform 1 0 3016 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5843_6
timestamp 1731220339
transform 1 0 2856 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5842_6
timestamp 1731220339
transform 1 0 3264 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5841_6
timestamp 1731220339
transform 1 0 3120 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5840_6
timestamp 1731220339
transform 1 0 2976 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5839_6
timestamp 1731220339
transform 1 0 2832 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5838_6
timestamp 1731220339
transform 1 0 3192 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5837_6
timestamp 1731220339
transform 1 0 3024 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5836_6
timestamp 1731220339
transform 1 0 2864 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5835_6
timestamp 1731220339
transform 1 0 2696 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5834_6
timestamp 1731220339
transform 1 0 2528 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5833_6
timestamp 1731220339
transform 1 0 2672 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5832_6
timestamp 1731220339
transform 1 0 2784 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5831_6
timestamp 1731220339
transform 1 0 2904 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5830_6
timestamp 1731220339
transform 1 0 3024 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5829_6
timestamp 1731220339
transform 1 0 3144 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5828_6
timestamp 1731220339
transform 1 0 3216 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5827_6
timestamp 1731220339
transform 1 0 3088 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5826_6
timestamp 1731220339
transform 1 0 2960 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5825_6
timestamp 1731220339
transform 1 0 2832 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5824_6
timestamp 1731220339
transform 1 0 2712 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5823_6
timestamp 1731220339
transform 1 0 2808 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5822_6
timestamp 1731220339
transform 1 0 2944 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5821_6
timestamp 1731220339
transform 1 0 3080 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5820_6
timestamp 1731220339
transform 1 0 3216 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5819_6
timestamp 1731220339
transform 1 0 3360 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5818_6
timestamp 1731220339
transform 1 0 3528 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5817_6
timestamp 1731220339
transform 1 0 3376 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5816_6
timestamp 1731220339
transform 1 0 3232 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5815_6
timestamp 1731220339
transform 1 0 3088 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5814_6
timestamp 1731220339
transform 1 0 2936 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5813_6
timestamp 1731220339
transform 1 0 2832 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5812_6
timestamp 1731220339
transform 1 0 2720 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5811_6
timestamp 1731220339
transform 1 0 2936 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5810_6
timestamp 1731220339
transform 1 0 3040 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5809_6
timestamp 1731220339
transform 1 0 3136 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5808_6
timestamp 1731220339
transform 1 0 3232 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5807_6
timestamp 1731220339
transform 1 0 3280 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5806_6
timestamp 1731220339
transform 1 0 3472 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5805_6
timestamp 1731220339
transform 1 0 3440 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5804_6
timestamp 1731220339
transform 1 0 3336 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5803_6
timestamp 1731220339
transform 1 0 3544 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5802_6
timestamp 1731220339
transform 1 0 3640 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5801_6
timestamp 1731220339
transform 1 0 3832 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5800_6
timestamp 1731220339
transform 1 0 3736 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5799_6
timestamp 1731220339
transform 1 0 3664 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5798_6
timestamp 1731220339
transform 1 0 3832 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5797_6
timestamp 1731220339
transform 1 0 3832 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5796_6
timestamp 1731220339
transform 1 0 3832 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5795_6
timestamp 1731220339
transform 1 0 3832 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5794_6
timestamp 1731220339
transform 1 0 3808 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5793_6
timestamp 1731220339
transform 1 0 3832 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5792_6
timestamp 1731220339
transform 1 0 3736 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5791_6
timestamp 1731220339
transform 1 0 3616 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5790_6
timestamp 1731220339
transform 1 0 3496 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5789_6
timestamp 1731220339
transform 1 0 3376 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5788_6
timestamp 1731220339
transform 1 0 3472 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5787_6
timestamp 1731220339
transform 1 0 3624 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5786_6
timestamp 1731220339
transform 1 0 3776 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5785_6
timestamp 1731220339
transform 1 0 3744 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5784_6
timestamp 1731220339
transform 1 0 3800 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5783_6
timestamp 1731220339
transform 1 0 3832 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5782_6
timestamp 1731220339
transform 1 0 3832 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5781_6
timestamp 1731220339
transform 1 0 3832 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5780_6
timestamp 1731220339
transform 1 0 3832 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5779_6
timestamp 1731220339
transform 1 0 3720 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5778_6
timestamp 1731220339
transform 1 0 3592 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5777_6
timestamp 1731220339
transform 1 0 3680 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5776_6
timestamp 1731220339
transform 1 0 3664 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5775_6
timestamp 1731220339
transform 1 0 3632 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5774_6
timestamp 1731220339
transform 1 0 3440 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5773_6
timestamp 1731220339
transform 1 0 3248 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5772_6
timestamp 1731220339
transform 1 0 3104 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5771_6
timestamp 1731220339
transform 1 0 3288 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5770_6
timestamp 1731220339
transform 1 0 3472 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5769_6
timestamp 1731220339
transform 1 0 3504 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5768_6
timestamp 1731220339
transform 1 0 3328 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5767_6
timestamp 1731220339
transform 1 0 3152 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5766_6
timestamp 1731220339
transform 1 0 3200 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5765_6
timestamp 1731220339
transform 1 0 3336 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5764_6
timestamp 1731220339
transform 1 0 3464 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5763_6
timestamp 1731220339
transform 1 0 3552 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5762_6
timestamp 1731220339
transform 1 0 3360 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5761_6
timestamp 1731220339
transform 1 0 3168 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5760_6
timestamp 1731220339
transform 1 0 3336 0 -1 4020
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5759_6
timestamp 1731220339
transform 1 0 3080 0 -1 4020
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5758_6
timestamp 1731220339
transform 1 0 2832 0 -1 4020
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5757_6
timestamp 1731220339
transform 1 0 2584 0 -1 4020
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5756_6
timestamp 1731220339
transform 1 0 2976 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5755_6
timestamp 1731220339
transform 1 0 3056 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5754_6
timestamp 1731220339
transform 1 0 2912 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5753_6
timestamp 1731220339
transform 1 0 2800 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5752_6
timestamp 1731220339
transform 1 0 2976 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5751_6
timestamp 1731220339
transform 1 0 2920 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5750_6
timestamp 1731220339
transform 1 0 3056 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5749_6
timestamp 1731220339
transform 1 0 2864 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5748_6
timestamp 1731220339
transform 1 0 2904 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5747_6
timestamp 1731220339
transform 1 0 3104 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5746_6
timestamp 1731220339
transform 1 0 3328 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5745_6
timestamp 1731220339
transform 1 0 3560 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5744_6
timestamp 1731220339
transform 1 0 3560 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5743_6
timestamp 1731220339
transform 1 0 3376 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5742_6
timestamp 1731220339
transform 1 0 3200 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5741_6
timestamp 1731220339
transform 1 0 3040 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5740_6
timestamp 1731220339
transform 1 0 3320 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5739_6
timestamp 1731220339
transform 1 0 3168 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5738_6
timestamp 1731220339
transform 1 0 3112 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5737_6
timestamp 1731220339
transform 1 0 3248 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5736_6
timestamp 1731220339
transform 1 0 3624 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5735_6
timestamp 1731220339
transform 1 0 3440 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5734_6
timestamp 1731220339
transform 1 0 3256 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5733_6
timestamp 1731220339
transform 1 0 3072 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5732_6
timestamp 1731220339
transform 1 0 3632 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5731_6
timestamp 1731220339
transform 1 0 3424 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5730_6
timestamp 1731220339
transform 1 0 3224 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5729_6
timestamp 1731220339
transform 1 0 3032 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5728_6
timestamp 1731220339
transform 1 0 2848 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5727_6
timestamp 1731220339
transform 1 0 3592 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5726_6
timestamp 1731220339
transform 1 0 3328 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5725_6
timestamp 1731220339
transform 1 0 3080 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5724_6
timestamp 1731220339
transform 1 0 2848 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5723_6
timestamp 1731220339
transform 1 0 3560 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5722_6
timestamp 1731220339
transform 1 0 3272 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5721_6
timestamp 1731220339
transform 1 0 2992 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5720_6
timestamp 1731220339
transform 1 0 2728 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5719_6
timestamp 1731220339
transform 1 0 2480 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5718_6
timestamp 1731220339
transform 1 0 2256 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5717_6
timestamp 1731220339
transform 1 0 3088 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5716_6
timestamp 1731220339
transform 1 0 2880 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5715_6
timestamp 1731220339
transform 1 0 2664 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5714_6
timestamp 1731220339
transform 1 0 2600 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5713_6
timestamp 1731220339
transform 1 0 2472 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5712_6
timestamp 1731220339
transform 1 0 2336 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5711_6
timestamp 1731220339
transform 1 0 2432 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5710_6
timestamp 1731220339
transform 1 0 2608 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5709_6
timestamp 1731220339
transform 1 0 2776 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5708_6
timestamp 1731220339
transform 1 0 2664 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5707_6
timestamp 1731220339
transform 1 0 2512 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5706_6
timestamp 1731220339
transform 1 0 2360 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5705_6
timestamp 1731220339
transform 1 0 2336 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5704_6
timestamp 1731220339
transform 1 0 2208 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5703_6
timestamp 1731220339
transform 1 0 2088 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5702_6
timestamp 1731220339
transform 1 0 2064 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5701_6
timestamp 1731220339
transform 1 0 2312 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5700_6
timestamp 1731220339
transform 1 0 2184 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5699_6
timestamp 1731220339
transform 1 0 2160 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5698_6
timestamp 1731220339
transform 1 0 2696 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5697_6
timestamp 1731220339
transform 1 0 2552 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5696_6
timestamp 1731220339
transform 1 0 2416 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5695_6
timestamp 1731220339
transform 1 0 2064 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5694_6
timestamp 1731220339
transform 1 0 2160 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5693_6
timestamp 1731220339
transform 1 0 2064 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5692_6
timestamp 1731220339
transform 1 0 1896 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5691_6
timestamp 1731220339
transform 1 0 1792 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5690_6
timestamp 1731220339
transform 1 0 1784 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5689_6
timestamp 1731220339
transform 1 0 1648 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5688_6
timestamp 1731220339
transform 1 0 1896 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5687_6
timestamp 1731220339
transform 1 0 1896 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5686_6
timestamp 1731220339
transform 1 0 1736 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5685_6
timestamp 1731220339
transform 1 0 1576 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5684_6
timestamp 1731220339
transform 1 0 1488 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5683_6
timestamp 1731220339
transform 1 0 1640 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5682_6
timestamp 1731220339
transform 1 0 1792 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5681_6
timestamp 1731220339
transform 1 0 1696 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5680_6
timestamp 1731220339
transform 1 0 1504 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5679_6
timestamp 1731220339
transform 1 0 1320 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5678_6
timestamp 1731220339
transform 1 0 1248 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5677_6
timestamp 1731220339
transform 1 0 1416 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5676_6
timestamp 1731220339
transform 1 0 1592 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5675_6
timestamp 1731220339
transform 1 0 1568 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5674_6
timestamp 1731220339
transform 1 0 1392 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5673_6
timestamp 1731220339
transform 1 0 1216 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5672_6
timestamp 1731220339
transform 1 0 1160 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5671_6
timestamp 1731220339
transform 1 0 1344 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5670_6
timestamp 1731220339
transform 1 0 1528 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5669_6
timestamp 1731220339
transform 1 0 1488 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5668_6
timestamp 1731220339
transform 1 0 1288 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5667_6
timestamp 1731220339
transform 1 0 1096 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5666_6
timestamp 1731220339
transform 1 0 928 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5665_6
timestamp 1731220339
transform 1 0 992 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5664_6
timestamp 1731220339
transform 1 0 840 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5663_6
timestamp 1731220339
transform 1 0 872 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5662_6
timestamp 1731220339
transform 1 0 1040 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5661_6
timestamp 1731220339
transform 1 0 1080 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5660_6
timestamp 1731220339
transform 1 0 912 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5659_6
timestamp 1731220339
transform 1 0 944 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5658_6
timestamp 1731220339
transform 1 0 1136 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5657_6
timestamp 1731220339
transform 1 0 1200 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5656_6
timestamp 1731220339
transform 1 0 1344 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5655_6
timestamp 1731220339
transform 1 0 1272 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5654_6
timestamp 1731220339
transform 1 0 1424 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5653_6
timestamp 1731220339
transform 1 0 1520 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5652_6
timestamp 1731220339
transform 1 0 1384 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5651_6
timestamp 1731220339
transform 1 0 1240 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5650_6
timestamp 1731220339
transform 1 0 1416 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5649_6
timestamp 1731220339
transform 1 0 1288 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5648_6
timestamp 1731220339
transform 1 0 1544 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5647_6
timestamp 1731220339
transform 1 0 1664 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5646_6
timestamp 1731220339
transform 1 0 1560 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5645_6
timestamp 1731220339
transform 1 0 1760 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5644_6
timestamp 1731220339
transform 1 0 1672 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5643_6
timestamp 1731220339
transform 1 0 1504 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5642_6
timestamp 1731220339
transform 1 0 1344 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5641_6
timestamp 1731220339
transform 1 0 1512 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5640_6
timestamp 1731220339
transform 1 0 1376 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5639_6
timestamp 1731220339
transform 1 0 1248 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5638_6
timestamp 1731220339
transform 1 0 1120 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5637_6
timestamp 1731220339
transform 1 0 984 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5636_6
timestamp 1731220339
transform 1 0 840 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5635_6
timestamp 1731220339
transform 1 0 864 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5634_6
timestamp 1731220339
transform 1 0 1024 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5633_6
timestamp 1731220339
transform 1 0 1184 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5632_6
timestamp 1731220339
transform 1 0 1360 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5631_6
timestamp 1731220339
transform 1 0 1168 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5630_6
timestamp 1731220339
transform 1 0 984 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5629_6
timestamp 1731220339
transform 1 0 816 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5628_6
timestamp 1731220339
transform 1 0 1160 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5627_6
timestamp 1731220339
transform 1 0 1024 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5626_6
timestamp 1731220339
transform 1 0 888 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5625_6
timestamp 1731220339
transform 1 0 760 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5624_6
timestamp 1731220339
transform 1 0 808 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5623_6
timestamp 1731220339
transform 1 0 1096 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5622_6
timestamp 1731220339
transform 1 0 952 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5621_6
timestamp 1731220339
transform 1 0 840 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5620_6
timestamp 1731220339
transform 1 0 976 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5619_6
timestamp 1731220339
transform 1 0 1120 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5618_6
timestamp 1731220339
transform 1 0 1064 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5617_6
timestamp 1731220339
transform 1 0 928 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5616_6
timestamp 1731220339
transform 1 0 800 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5615_6
timestamp 1731220339
transform 1 0 680 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5614_6
timestamp 1731220339
transform 1 0 568 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5613_6
timestamp 1731220339
transform 1 0 712 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5612_6
timestamp 1731220339
transform 1 0 600 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5611_6
timestamp 1731220339
transform 1 0 496 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5610_6
timestamp 1731220339
transform 1 0 528 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5609_6
timestamp 1731220339
transform 1 0 664 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5608_6
timestamp 1731220339
transform 1 0 640 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5607_6
timestamp 1731220339
transform 1 0 528 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5606_6
timestamp 1731220339
transform 1 0 408 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5605_6
timestamp 1731220339
transform 1 0 528 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5604_6
timestamp 1731220339
transform 1 0 664 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5603_6
timestamp 1731220339
transform 1 0 704 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5602_6
timestamp 1731220339
transform 1 0 544 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5601_6
timestamp 1731220339
transform 1 0 384 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5600_6
timestamp 1731220339
transform 1 0 240 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5599_6
timestamp 1731220339
transform 1 0 128 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5598_6
timestamp 1731220339
transform 1 0 128 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5597_6
timestamp 1731220339
transform 1 0 240 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5596_6
timestamp 1731220339
transform 1 0 392 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5595_6
timestamp 1731220339
transform 1 0 544 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5594_6
timestamp 1731220339
transform 1 0 696 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5593_6
timestamp 1731220339
transform 1 0 936 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5592_6
timestamp 1731220339
transform 1 0 744 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5591_6
timestamp 1731220339
transform 1 0 560 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5590_6
timestamp 1731220339
transform 1 0 384 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5589_6
timestamp 1731220339
transform 1 0 224 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5588_6
timestamp 1731220339
transform 1 0 504 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5587_6
timestamp 1731220339
transform 1 0 616 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5586_6
timestamp 1731220339
transform 1 0 736 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5585_6
timestamp 1731220339
transform 1 0 856 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5584_6
timestamp 1731220339
transform 1 0 976 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5583_6
timestamp 1731220339
transform 1 0 1032 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5582_6
timestamp 1731220339
transform 1 0 920 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5581_6
timestamp 1731220339
transform 1 0 808 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5580_6
timestamp 1731220339
transform 1 0 704 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5579_6
timestamp 1731220339
transform 1 0 608 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5578_6
timestamp 1731220339
transform 1 0 960 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5577_6
timestamp 1731220339
transform 1 0 792 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5576_6
timestamp 1731220339
transform 1 0 632 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5575_6
timestamp 1731220339
transform 1 0 488 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5574_6
timestamp 1731220339
transform 1 0 360 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5573_6
timestamp 1731220339
transform 1 0 736 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5572_6
timestamp 1731220339
transform 1 0 560 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5571_6
timestamp 1731220339
transform 1 0 392 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5570_6
timestamp 1731220339
transform 1 0 240 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5569_6
timestamp 1731220339
transform 1 0 128 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5568_6
timestamp 1731220339
transform 1 0 128 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5567_6
timestamp 1731220339
transform 1 0 248 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5566_6
timestamp 1731220339
transform 1 0 416 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5565_6
timestamp 1731220339
transform 1 0 608 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5564_6
timestamp 1731220339
transform 1 0 824 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5563_6
timestamp 1731220339
transform 1 0 768 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5562_6
timestamp 1731220339
transform 1 0 576 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5561_6
timestamp 1731220339
transform 1 0 400 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5560_6
timestamp 1731220339
transform 1 0 232 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5559_6
timestamp 1731220339
transform 1 0 456 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5558_6
timestamp 1731220339
transform 1 0 576 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5557_6
timestamp 1731220339
transform 1 0 704 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5556_6
timestamp 1731220339
transform 1 0 848 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5555_6
timestamp 1731220339
transform 1 0 1000 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5554_6
timestamp 1731220339
transform 1 0 1136 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5553_6
timestamp 1731220339
transform 1 0 1008 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5552_6
timestamp 1731220339
transform 1 0 880 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5551_6
timestamp 1731220339
transform 1 0 760 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5550_6
timestamp 1731220339
transform 1 0 648 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5549_6
timestamp 1731220339
transform 1 0 928 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5548_6
timestamp 1731220339
transform 1 0 792 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5547_6
timestamp 1731220339
transform 1 0 664 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5546_6
timestamp 1731220339
transform 1 0 544 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5545_6
timestamp 1731220339
transform 1 0 432 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5544_6
timestamp 1731220339
transform 1 0 800 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5543_6
timestamp 1731220339
transform 1 0 624 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5542_6
timestamp 1731220339
transform 1 0 456 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5541_6
timestamp 1731220339
transform 1 0 296 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5540_6
timestamp 1731220339
transform 1 0 160 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5539_6
timestamp 1731220339
transform 1 0 688 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5538_6
timestamp 1731220339
transform 1 0 520 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5537_6
timestamp 1731220339
transform 1 0 368 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5536_6
timestamp 1731220339
transform 1 0 232 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5535_6
timestamp 1731220339
transform 1 0 128 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5534_6
timestamp 1731220339
transform 1 0 648 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5533_6
timestamp 1731220339
transform 1 0 464 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5532_6
timestamp 1731220339
transform 1 0 280 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5531_6
timestamp 1731220339
transform 1 0 128 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5530_6
timestamp 1731220339
transform 1 0 128 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5529_6
timestamp 1731220339
transform 1 0 288 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5528_6
timestamp 1731220339
transform 1 0 464 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5527_6
timestamp 1731220339
transform 1 0 312 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5526_6
timestamp 1731220339
transform 1 0 152 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5525_6
timestamp 1731220339
transform 1 0 216 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5524_6
timestamp 1731220339
transform 1 0 376 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5523_6
timestamp 1731220339
transform 1 0 304 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5522_6
timestamp 1731220339
transform 1 0 632 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5521_6
timestamp 1731220339
transform 1 0 464 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5520_6
timestamp 1731220339
transform 1 0 440 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5519_6
timestamp 1731220339
transform 1 0 288 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5518_6
timestamp 1731220339
transform 1 0 232 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5517_6
timestamp 1731220339
transform 1 0 408 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5516_6
timestamp 1731220339
transform 1 0 456 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5515_6
timestamp 1731220339
transform 1 0 280 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5514_6
timestamp 1731220339
transform 1 0 128 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5513_6
timestamp 1731220339
transform 1 0 128 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5512_6
timestamp 1731220339
transform 1 0 272 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5511_6
timestamp 1731220339
transform 1 0 136 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5510_6
timestamp 1731220339
transform 1 0 312 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5509_6
timestamp 1731220339
transform 1 0 552 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5508_6
timestamp 1731220339
transform 1 0 384 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5507_6
timestamp 1731220339
transform 1 0 216 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5506_6
timestamp 1731220339
transform 1 0 144 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5505_6
timestamp 1731220339
transform 1 0 240 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5504_6
timestamp 1731220339
transform 1 0 336 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5503_6
timestamp 1731220339
transform 1 0 432 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5502_6
timestamp 1731220339
transform 1 0 528 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5501_6
timestamp 1731220339
transform 1 0 624 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5500_6
timestamp 1731220339
transform 1 0 720 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5499_6
timestamp 1731220339
transform 1 0 816 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5498_6
timestamp 1731220339
transform 1 0 896 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5497_6
timestamp 1731220339
transform 1 0 728 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5496_6
timestamp 1731220339
transform 1 0 624 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5495_6
timestamp 1731220339
transform 1 0 472 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5494_6
timestamp 1731220339
transform 1 0 768 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5493_6
timestamp 1731220339
transform 1 0 712 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5492_6
timestamp 1731220339
transform 1 0 576 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5491_6
timestamp 1731220339
transform 1 0 432 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5490_6
timestamp 1731220339
transform 1 0 632 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5489_6
timestamp 1731220339
transform 1 0 800 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5488_6
timestamp 1731220339
transform 1 0 984 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5487_6
timestamp 1731220339
transform 1 0 792 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5486_6
timestamp 1731220339
transform 1 0 600 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5485_6
timestamp 1731220339
transform 1 0 608 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5484_6
timestamp 1731220339
transform 1 0 776 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5483_6
timestamp 1731220339
transform 1 0 944 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5482_6
timestamp 1731220339
transform 1 0 968 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5481_6
timestamp 1731220339
transform 1 0 800 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5480_6
timestamp 1731220339
transform 1 0 808 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5479_6
timestamp 1731220339
transform 1 0 672 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5478_6
timestamp 1731220339
transform 1 0 528 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5477_6
timestamp 1731220339
transform 1 0 464 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5476_6
timestamp 1731220339
transform 1 0 608 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5475_6
timestamp 1731220339
transform 1 0 744 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5474_6
timestamp 1731220339
transform 1 0 632 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5473_6
timestamp 1731220339
transform 1 0 792 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5472_6
timestamp 1731220339
transform 1 0 944 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5471_6
timestamp 1731220339
transform 1 0 1008 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5470_6
timestamp 1731220339
transform 1 0 832 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5469_6
timestamp 1731220339
transform 1 0 856 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5468_6
timestamp 1731220339
transform 1 0 1032 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5467_6
timestamp 1731220339
transform 1 0 1208 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5466_6
timestamp 1731220339
transform 1 0 1152 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5465_6
timestamp 1731220339
transform 1 0 976 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5464_6
timestamp 1731220339
transform 1 0 1072 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5463_6
timestamp 1731220339
transform 1 0 1224 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5462_6
timestamp 1731220339
transform 1 0 1384 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5461_6
timestamp 1731220339
transform 1 0 1408 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5460_6
timestamp 1731220339
transform 1 0 1272 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5459_6
timestamp 1731220339
transform 1 0 1160 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5458_6
timestamp 1731220339
transform 1 0 1328 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5457_6
timestamp 1731220339
transform 1 0 1504 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5456_6
timestamp 1731220339
transform 1 0 1344 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5455_6
timestamp 1731220339
transform 1 0 1152 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5454_6
timestamp 1731220339
transform 1 0 960 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5453_6
timestamp 1731220339
transform 1 0 1056 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5452_6
timestamp 1731220339
transform 1 0 1304 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5451_6
timestamp 1731220339
transform 1 0 1336 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5450_6
timestamp 1731220339
transform 1 0 1128 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5449_6
timestamp 1731220339
transform 1 0 928 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5448_6
timestamp 1731220339
transform 1 0 1136 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5447_6
timestamp 1731220339
transform 1 0 1320 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5446_6
timestamp 1731220339
transform 1 0 1392 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5445_6
timestamp 1731220339
transform 1 0 1272 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5444_6
timestamp 1731220339
transform 1 0 1152 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5443_6
timestamp 1731220339
transform 1 0 1096 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5442_6
timestamp 1731220339
transform 1 0 1216 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5441_6
timestamp 1731220339
transform 1 0 1328 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5440_6
timestamp 1731220339
transform 1 0 1328 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5439_6
timestamp 1731220339
transform 1 0 1128 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5438_6
timestamp 1731220339
transform 1 0 1536 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5437_6
timestamp 1731220339
transform 1 0 1448 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5436_6
timestamp 1731220339
transform 1 0 1568 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5435_6
timestamp 1731220339
transform 1 0 1688 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5434_6
timestamp 1731220339
transform 1 0 1632 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5433_6
timestamp 1731220339
transform 1 0 1512 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5432_6
timestamp 1731220339
transform 1 0 1504 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5431_6
timestamp 1731220339
transform 1 0 1696 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5430_6
timestamp 1731220339
transform 1 0 1760 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5429_6
timestamp 1731220339
transform 1 0 1544 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5428_6
timestamp 1731220339
transform 1 0 1560 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5427_6
timestamp 1731220339
transform 1 0 1824 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5426_6
timestamp 1731220339
transform 1 0 1728 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5425_6
timestamp 1731220339
transform 1 0 1536 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5424_6
timestamp 1731220339
transform 1 0 1896 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5423_6
timestamp 1731220339
transform 1 0 1864 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5422_6
timestamp 1731220339
transform 1 0 1680 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5421_6
timestamp 1731220339
transform 1 0 1840 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5420_6
timestamp 1731220339
transform 1 0 1696 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5419_6
timestamp 1731220339
transform 1 0 1552 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5418_6
timestamp 1731220339
transform 1 0 1544 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5417_6
timestamp 1731220339
transform 1 0 1712 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5416_6
timestamp 1731220339
transform 1 0 1688 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5415_6
timestamp 1731220339
transform 1 0 1504 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5414_6
timestamp 1731220339
transform 1 0 1328 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5413_6
timestamp 1731220339
transform 1 0 1560 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5412_6
timestamp 1731220339
transform 1 0 1384 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5411_6
timestamp 1731220339
transform 1 0 1376 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5410_6
timestamp 1731220339
transform 1 0 1192 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5409_6
timestamp 1731220339
transform 1 0 1560 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5408_6
timestamp 1731220339
transform 1 0 1488 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5407_6
timestamp 1731220339
transform 1 0 1352 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5406_6
timestamp 1731220339
transform 1 0 1216 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5405_6
timestamp 1731220339
transform 1 0 1080 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5404_6
timestamp 1731220339
transform 1 0 1344 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5403_6
timestamp 1731220339
transform 1 0 1224 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5402_6
timestamp 1731220339
transform 1 0 1104 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5401_6
timestamp 1731220339
transform 1 0 992 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5400_6
timestamp 1731220339
transform 1 0 872 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5399_6
timestamp 1731220339
transform 1 0 944 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5398_6
timestamp 1731220339
transform 1 0 1072 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5397_6
timestamp 1731220339
transform 1 0 1192 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5396_6
timestamp 1731220339
transform 1 0 1448 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5395_6
timestamp 1731220339
transform 1 0 1320 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5394_6
timestamp 1731220339
transform 1 0 1288 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5393_6
timestamp 1731220339
transform 1 0 1128 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5392_6
timestamp 1731220339
transform 1 0 1760 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5391_6
timestamp 1731220339
transform 1 0 1600 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5390_6
timestamp 1731220339
transform 1 0 1448 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5389_6
timestamp 1731220339
transform 1 0 1392 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5388_6
timestamp 1731220339
transform 1 0 1256 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5387_6
timestamp 1731220339
transform 1 0 1104 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5386_6
timestamp 1731220339
transform 1 0 1528 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5385_6
timestamp 1731220339
transform 1 0 1656 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5384_6
timestamp 1731220339
transform 1 0 1856 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5383_6
timestamp 1731220339
transform 1 0 1680 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5382_6
timestamp 1731220339
transform 1 0 1512 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5381_6
timestamp 1731220339
transform 1 0 1344 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5380_6
timestamp 1731220339
transform 1 0 1168 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5379_6
timestamp 1731220339
transform 1 0 1560 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5378_6
timestamp 1731220339
transform 1 0 1408 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5377_6
timestamp 1731220339
transform 1 0 1264 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5376_6
timestamp 1731220339
transform 1 0 1112 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5375_6
timestamp 1731220339
transform 1 0 960 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5374_6
timestamp 1731220339
transform 1 0 1320 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5373_6
timestamp 1731220339
transform 1 0 1200 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5372_6
timestamp 1731220339
transform 1 0 1080 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5371_6
timestamp 1731220339
transform 1 0 960 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5370_6
timestamp 1731220339
transform 1 0 840 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5369_6
timestamp 1731220339
transform 1 0 896 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5368_6
timestamp 1731220339
transform 1 0 1024 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5367_6
timestamp 1731220339
transform 1 0 1144 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5366_6
timestamp 1731220339
transform 1 0 1264 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5365_6
timestamp 1731220339
transform 1 0 1384 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5364_6
timestamp 1731220339
transform 1 0 1656 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5363_6
timestamp 1731220339
transform 1 0 1504 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5362_6
timestamp 1731220339
transform 1 0 1352 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5361_6
timestamp 1731220339
transform 1 0 1208 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5360_6
timestamp 1731220339
transform 1 0 1056 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5359_6
timestamp 1731220339
transform 1 0 1008 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5358_6
timestamp 1731220339
transform 1 0 912 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5357_6
timestamp 1731220339
transform 1 0 1104 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5356_6
timestamp 1731220339
transform 1 0 1200 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5355_6
timestamp 1731220339
transform 1 0 1296 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5354_6
timestamp 1731220339
transform 1 0 1400 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5353_6
timestamp 1731220339
transform 1 0 1504 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5352_6
timestamp 1731220339
transform 1 0 1608 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5351_6
timestamp 1731220339
transform 1 0 1704 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5350_6
timestamp 1731220339
transform 1 0 1800 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5349_6
timestamp 1731220339
transform 1 0 1896 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5348_6
timestamp 1731220339
transform 1 0 2064 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5347_6
timestamp 1731220339
transform 1 0 2184 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5346_6
timestamp 1731220339
transform 1 0 2640 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5345_6
timestamp 1731220339
transform 1 0 2488 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5344_6
timestamp 1731220339
transform 1 0 2336 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5343_6
timestamp 1731220339
transform 1 0 2208 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5342_6
timestamp 1731220339
transform 1 0 2064 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5341_6
timestamp 1731220339
transform 1 0 2784 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5340_6
timestamp 1731220339
transform 1 0 2584 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5339_6
timestamp 1731220339
transform 1 0 2392 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5338_6
timestamp 1731220339
transform 1 0 2320 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5337_6
timestamp 1731220339
transform 1 0 2184 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5336_6
timestamp 1731220339
transform 1 0 2464 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5335_6
timestamp 1731220339
transform 1 0 2776 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5334_6
timestamp 1731220339
transform 1 0 2616 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5333_6
timestamp 1731220339
transform 1 0 2520 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5332_6
timestamp 1731220339
transform 1 0 2424 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5331_6
timestamp 1731220339
transform 1 0 2616 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5330_6
timestamp 1731220339
transform 1 0 2712 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5329_6
timestamp 1731220339
transform 1 0 2808 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5328_6
timestamp 1731220339
transform 1 0 2992 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5327_6
timestamp 1731220339
transform 1 0 2840 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5326_6
timestamp 1731220339
transform 1 0 2720 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5325_6
timestamp 1731220339
transform 1 0 2616 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5324_6
timestamp 1731220339
transform 1 0 2520 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5323_6
timestamp 1731220339
transform 1 0 2424 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5322_6
timestamp 1731220339
transform 1 0 2576 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5321_6
timestamp 1731220339
transform 1 0 2472 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5320_6
timestamp 1731220339
transform 1 0 2376 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5319_6
timestamp 1731220339
transform 1 0 2280 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5318_6
timestamp 1731220339
transform 1 0 2184 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5317_6
timestamp 1731220339
transform 1 0 2416 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5316_6
timestamp 1731220339
transform 1 0 2232 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5315_6
timestamp 1731220339
transform 1 0 2064 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5314_6
timestamp 1731220339
transform 1 0 1896 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5313_6
timestamp 1731220339
transform 1 0 1784 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5312_6
timestamp 1731220339
transform 1 0 1896 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5311_6
timestamp 1731220339
transform 1 0 2064 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5310_6
timestamp 1731220339
transform 1 0 2176 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5309_6
timestamp 1731220339
transform 1 0 2328 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5308_6
timestamp 1731220339
transform 1 0 2480 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5307_6
timestamp 1731220339
transform 1 0 2632 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5306_6
timestamp 1731220339
transform 1 0 2608 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5305_6
timestamp 1731220339
transform 1 0 2464 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5304_6
timestamp 1731220339
transform 1 0 2328 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5303_6
timestamp 1731220339
transform 1 0 2760 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5302_6
timestamp 1731220339
transform 1 0 2912 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5301_6
timestamp 1731220339
transform 1 0 3072 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5300_6
timestamp 1731220339
transform 1 0 2936 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5299_6
timestamp 1731220339
transform 1 0 2800 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5298_6
timestamp 1731220339
transform 1 0 2672 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5297_6
timestamp 1731220339
transform 1 0 2552 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5296_6
timestamp 1731220339
transform 1 0 2944 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5295_6
timestamp 1731220339
transform 1 0 2776 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5294_6
timestamp 1731220339
transform 1 0 2608 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5293_6
timestamp 1731220339
transform 1 0 2448 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5292_6
timestamp 1731220339
transform 1 0 2296 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5291_6
timestamp 1731220339
transform 1 0 2696 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5290_6
timestamp 1731220339
transform 1 0 2480 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5289_6
timestamp 1731220339
transform 1 0 2256 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5288_6
timestamp 1731220339
transform 1 0 2064 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5287_6
timestamp 1731220339
transform 1 0 1896 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5286_6
timestamp 1731220339
transform 1 0 1736 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5285_6
timestamp 1731220339
transform 1 0 2064 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5284_6
timestamp 1731220339
transform 1 0 2504 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5283_6
timestamp 1731220339
transform 1 0 2344 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5282_6
timestamp 1731220339
transform 1 0 2192 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5281_6
timestamp 1731220339
transform 1 0 2176 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5280_6
timestamp 1731220339
transform 1 0 2064 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5279_6
timestamp 1731220339
transform 1 0 2552 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5278_6
timestamp 1731220339
transform 1 0 2424 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5277_6
timestamp 1731220339
transform 1 0 2296 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5276_6
timestamp 1731220339
transform 1 0 2240 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5275_6
timestamp 1731220339
transform 1 0 2368 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5274_6
timestamp 1731220339
transform 1 0 2784 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5273_6
timestamp 1731220339
transform 1 0 2640 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5272_6
timestamp 1731220339
transform 1 0 2504 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5271_6
timestamp 1731220339
transform 1 0 2392 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5270_6
timestamp 1731220339
transform 1 0 2528 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5269_6
timestamp 1731220339
transform 1 0 2960 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5268_6
timestamp 1731220339
transform 1 0 2816 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5267_6
timestamp 1731220339
transform 1 0 2672 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5266_6
timestamp 1731220339
transform 1 0 2624 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5265_6
timestamp 1731220339
transform 1 0 2512 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5264_6
timestamp 1731220339
transform 1 0 2752 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5263_6
timestamp 1731220339
transform 1 0 2888 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5262_6
timestamp 1731220339
transform 1 0 3024 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5261_6
timestamp 1731220339
transform 1 0 3168 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5260_6
timestamp 1731220339
transform 1 0 3064 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5259_6
timestamp 1731220339
transform 1 0 2928 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5258_6
timestamp 1731220339
transform 1 0 2792 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5257_6
timestamp 1731220339
transform 1 0 2664 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5256_6
timestamp 1731220339
transform 1 0 2536 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5255_6
timestamp 1731220339
transform 1 0 2848 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5254_6
timestamp 1731220339
transform 1 0 2728 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5253_6
timestamp 1731220339
transform 1 0 2608 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5252_6
timestamp 1731220339
transform 1 0 2496 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5251_6
timestamp 1731220339
transform 1 0 2384 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5250_6
timestamp 1731220339
transform 1 0 2680 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5249_6
timestamp 1731220339
transform 1 0 2552 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5248_6
timestamp 1731220339
transform 1 0 2432 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5247_6
timestamp 1731220339
transform 1 0 2320 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5246_6
timestamp 1731220339
transform 1 0 2216 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5245_6
timestamp 1731220339
transform 1 0 2648 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5244_6
timestamp 1731220339
transform 1 0 2480 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5243_6
timestamp 1731220339
transform 1 0 2320 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5242_6
timestamp 1731220339
transform 1 0 2176 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5241_6
timestamp 1731220339
transform 1 0 2064 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5240_6
timestamp 1731220339
transform 1 0 2064 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5239_6
timestamp 1731220339
transform 1 0 2192 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5238_6
timestamp 1731220339
transform 1 0 2712 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5237_6
timestamp 1731220339
transform 1 0 2536 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5236_6
timestamp 1731220339
transform 1 0 2360 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5235_6
timestamp 1731220339
transform 1 0 2232 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5234_6
timestamp 1731220339
transform 1 0 2064 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5233_6
timestamp 1731220339
transform 1 0 2888 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5232_6
timestamp 1731220339
transform 1 0 2664 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5231_6
timestamp 1731220339
transform 1 0 2440 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5230_6
timestamp 1731220339
transform 1 0 2392 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5229_6
timestamp 1731220339
transform 1 0 2184 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5228_6
timestamp 1731220339
transform 1 0 2640 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5227_6
timestamp 1731220339
transform 1 0 3208 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5226_6
timestamp 1731220339
transform 1 0 2912 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5225_6
timestamp 1731220339
transform 1 0 2776 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5224_6
timestamp 1731220339
transform 1 0 2584 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5223_6
timestamp 1731220339
transform 1 0 2488 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5222_6
timestamp 1731220339
transform 1 0 2392 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5221_6
timestamp 1731220339
transform 1 0 2680 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5220_6
timestamp 1731220339
transform 1 0 2680 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5219_6
timestamp 1731220339
transform 1 0 2496 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5218_6
timestamp 1731220339
transform 1 0 2288 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5217_6
timestamp 1731220339
transform 1 0 2280 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5216_6
timestamp 1731220339
transform 1 0 2352 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5215_6
timestamp 1731220339
transform 1 0 2432 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5214_6
timestamp 1731220339
transform 1 0 2552 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5213_6
timestamp 1731220339
transform 1 0 2592 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5212_6
timestamp 1731220339
transform 1 0 2464 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5211_6
timestamp 1731220339
transform 1 0 2208 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5210_6
timestamp 1731220339
transform 1 0 2256 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5209_6
timestamp 1731220339
transform 1 0 2088 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5208_6
timestamp 1731220339
transform 1 0 2192 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5207_6
timestamp 1731220339
transform 1 0 2064 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5206_6
timestamp 1731220339
transform 1 0 1896 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5205_6
timestamp 1731220339
transform 1 0 1744 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5204_6
timestamp 1731220339
transform 1 0 1896 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5203_6
timestamp 1731220339
transform 1 0 1720 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5202_6
timestamp 1731220339
transform 1 0 1704 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5201_6
timestamp 1731220339
transform 1 0 1896 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5200_6
timestamp 1731220339
transform 1 0 2064 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5199_6
timestamp 1731220339
transform 1 0 2064 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5198_6
timestamp 1731220339
transform 1 0 2176 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5197_6
timestamp 1731220339
transform 1 0 2648 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5196_6
timestamp 1731220339
transform 1 0 2472 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5195_6
timestamp 1731220339
transform 1 0 2320 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5194_6
timestamp 1731220339
transform 1 0 2216 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5193_6
timestamp 1731220339
transform 1 0 2072 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5192_6
timestamp 1731220339
transform 1 0 2680 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5191_6
timestamp 1731220339
transform 1 0 2520 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5190_6
timestamp 1731220339
transform 1 0 2368 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5189_6
timestamp 1731220339
transform 1 0 2240 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5188_6
timestamp 1731220339
transform 1 0 2392 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5187_6
timestamp 1731220339
transform 1 0 2896 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5186_6
timestamp 1731220339
transform 1 0 2720 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5185_6
timestamp 1731220339
transform 1 0 2552 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5184_6
timestamp 1731220339
transform 1 0 2544 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5183_6
timestamp 1731220339
transform 1 0 2408 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5182_6
timestamp 1731220339
transform 1 0 2968 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5181_6
timestamp 1731220339
transform 1 0 2824 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5180_6
timestamp 1731220339
transform 1 0 2680 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5179_6
timestamp 1731220339
transform 1 0 2560 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5178_6
timestamp 1731220339
transform 1 0 2712 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5177_6
timestamp 1731220339
transform 1 0 2864 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5176_6
timestamp 1731220339
transform 1 0 3016 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5175_6
timestamp 1731220339
transform 1 0 2896 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5174_6
timestamp 1731220339
transform 1 0 2768 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5173_6
timestamp 1731220339
transform 1 0 2656 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5172_6
timestamp 1731220339
transform 1 0 2544 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5171_6
timestamp 1731220339
transform 1 0 2440 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5170_6
timestamp 1731220339
transform 1 0 2728 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5169_6
timestamp 1731220339
transform 1 0 2576 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5168_6
timestamp 1731220339
transform 1 0 2440 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5167_6
timestamp 1731220339
transform 1 0 2320 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5166_6
timestamp 1731220339
transform 1 0 2664 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5165_6
timestamp 1731220339
transform 1 0 2464 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5164_6
timestamp 1731220339
transform 1 0 2272 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5163_6
timestamp 1731220339
transform 1 0 2096 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5162_6
timestamp 1731220339
transform 1 0 2728 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5161_6
timestamp 1731220339
transform 1 0 2544 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5160_6
timestamp 1731220339
transform 1 0 2360 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5159_6
timestamp 1731220339
transform 1 0 2192 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5158_6
timestamp 1731220339
transform 1 0 2064 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5157_6
timestamp 1731220339
transform 1 0 2064 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5156_6
timestamp 1731220339
transform 1 0 2176 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5155_6
timestamp 1731220339
transform 1 0 2320 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5154_6
timestamp 1731220339
transform 1 0 2632 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5153_6
timestamp 1731220339
transform 1 0 2472 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5152_6
timestamp 1731220339
transform 1 0 2368 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5151_6
timestamp 1731220339
transform 1 0 2256 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5150_6
timestamp 1731220339
transform 1 0 2488 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5149_6
timestamp 1731220339
transform 1 0 2624 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5148_6
timestamp 1731220339
transform 1 0 2768 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5147_6
timestamp 1731220339
transform 1 0 2792 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5146_6
timestamp 1731220339
transform 1 0 2608 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5145_6
timestamp 1731220339
transform 1 0 2432 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5144_6
timestamp 1731220339
transform 1 0 2264 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5143_6
timestamp 1731220339
transform 1 0 2120 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5142_6
timestamp 1731220339
transform 1 0 2320 0 -1 4020
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5141_6
timestamp 1731220339
transform 1 0 2064 0 -1 4020
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5140_6
timestamp 1731220339
transform 1 0 1896 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5139_6
timestamp 1731220339
transform 1 0 1784 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5138_6
timestamp 1731220339
transform 1 0 1648 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5137_6
timestamp 1731220339
transform 1 0 1512 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5136_6
timestamp 1731220339
transform 1 0 1376 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5135_6
timestamp 1731220339
transform 1 0 1224 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5134_6
timestamp 1731220339
transform 1 0 1056 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5133_6
timestamp 1731220339
transform 1 0 1280 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5132_6
timestamp 1731220339
transform 1 0 1472 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5131_6
timestamp 1731220339
transform 1 0 1672 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5130_6
timestamp 1731220339
transform 1 0 1624 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5129_6
timestamp 1731220339
transform 1 0 1496 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5128_6
timestamp 1731220339
transform 1 0 1600 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5127_6
timestamp 1731220339
transform 1 0 1472 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5126_6
timestamp 1731220339
transform 1 0 1688 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5125_6
timestamp 1731220339
transform 1 0 1680 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5124_6
timestamp 1731220339
transform 1 0 1768 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5123_6
timestamp 1731220339
transform 1 0 1592 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5122_6
timestamp 1731220339
transform 1 0 1632 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5121_6
timestamp 1731220339
transform 1 0 1808 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5120_6
timestamp 1731220339
transform 1 0 1816 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5119_6
timestamp 1731220339
transform 1 0 1624 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5118_6
timestamp 1731220339
transform 1 0 1792 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5117_6
timestamp 1731220339
transform 1 0 1616 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5116_6
timestamp 1731220339
transform 1 0 1568 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5115_6
timestamp 1731220339
transform 1 0 1728 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5114_6
timestamp 1731220339
transform 1 0 1760 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5113_6
timestamp 1731220339
transform 1 0 1600 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5112_6
timestamp 1731220339
transform 1 0 1448 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5111_6
timestamp 1731220339
transform 1 0 1296 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5110_6
timestamp 1731220339
transform 1 0 1136 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5109_6
timestamp 1731220339
transform 1 0 1096 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5108_6
timestamp 1731220339
transform 1 0 1256 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5107_6
timestamp 1731220339
transform 1 0 1416 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5106_6
timestamp 1731220339
transform 1 0 1440 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5105_6
timestamp 1731220339
transform 1 0 1264 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5104_6
timestamp 1731220339
transform 1 0 1088 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5103_6
timestamp 1731220339
transform 1 0 1048 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5102_6
timestamp 1731220339
transform 1 0 1432 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5101_6
timestamp 1731220339
transform 1 0 1240 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5100_6
timestamp 1731220339
transform 1 0 1120 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_599_6
timestamp 1731220339
transform 1 0 1288 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_598_6
timestamp 1731220339
transform 1 0 1456 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_597_6
timestamp 1731220339
transform 1 0 1416 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_596_6
timestamp 1731220339
transform 1 0 1240 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_595_6
timestamp 1731220339
transform 1 0 1072 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_594_6
timestamp 1731220339
transform 1 0 984 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_593_6
timestamp 1731220339
transform 1 0 1208 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_592_6
timestamp 1731220339
transform 1 0 1440 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_591_6
timestamp 1731220339
transform 1 0 1256 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_590_6
timestamp 1731220339
transform 1 0 1048 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_589_6
timestamp 1731220339
transform 1 0 832 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_588_6
timestamp 1731220339
transform 1 0 1376 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_587_6
timestamp 1731220339
transform 1 0 1160 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_586_6
timestamp 1731220339
transform 1 0 952 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_585_6
timestamp 1731220339
transform 1 0 744 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_584_6
timestamp 1731220339
transform 1 0 1376 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_583_6
timestamp 1731220339
transform 1 0 1256 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_582_6
timestamp 1731220339
transform 1 0 1144 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_581_6
timestamp 1731220339
transform 1 0 1032 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_580_6
timestamp 1731220339
transform 1 0 928 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_579_6
timestamp 1731220339
transform 1 0 824 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_578_6
timestamp 1731220339
transform 1 0 720 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_577_6
timestamp 1731220339
transform 1 0 624 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_576_6
timestamp 1731220339
transform 1 0 528 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_575_6
timestamp 1731220339
transform 1 0 432 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_574_6
timestamp 1731220339
transform 1 0 1088 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_573_6
timestamp 1731220339
transform 1 0 904 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_572_6
timestamp 1731220339
transform 1 0 728 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_571_6
timestamp 1731220339
transform 1 0 560 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_570_6
timestamp 1731220339
transform 1 0 880 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_569_6
timestamp 1731220339
transform 1 0 696 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_568_6
timestamp 1731220339
transform 1 0 504 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_567_6
timestamp 1731220339
transform 1 0 304 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_566_6
timestamp 1731220339
transform 1 0 408 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_565_6
timestamp 1731220339
transform 1 0 272 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_564_6
timestamp 1731220339
transform 1 0 224 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_563_6
timestamp 1731220339
transform 1 0 328 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_562_6
timestamp 1731220339
transform 1 0 544 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_561_6
timestamp 1731220339
transform 1 0 344 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_560_6
timestamp 1731220339
transform 1 0 152 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_559_6
timestamp 1731220339
transform 1 0 144 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_558_6
timestamp 1731220339
transform 1 0 376 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_557_6
timestamp 1731220339
transform 1 0 608 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_556_6
timestamp 1731220339
transform 1 0 768 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_555_6
timestamp 1731220339
transform 1 0 552 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_554_6
timestamp 1731220339
transform 1 0 352 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_553_6
timestamp 1731220339
transform 1 0 160 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_552_6
timestamp 1731220339
transform 1 0 288 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_551_6
timestamp 1731220339
transform 1 0 424 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_550_6
timestamp 1731220339
transform 1 0 576 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_549_6
timestamp 1731220339
transform 1 0 736 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_548_6
timestamp 1731220339
transform 1 0 904 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_547_6
timestamp 1731220339
transform 1 0 952 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_546_6
timestamp 1731220339
transform 1 0 792 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_545_6
timestamp 1731220339
transform 1 0 640 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_544_6
timestamp 1731220339
transform 1 0 488 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_543_6
timestamp 1731220339
transform 1 0 664 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_542_6
timestamp 1731220339
transform 1 0 856 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_541_6
timestamp 1731220339
transform 1 0 904 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_540_6
timestamp 1731220339
transform 1 0 712 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_539_6
timestamp 1731220339
transform 1 0 512 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_538_6
timestamp 1731220339
transform 1 0 736 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_537_6
timestamp 1731220339
transform 1 0 920 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_536_6
timestamp 1731220339
transform 1 0 968 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_535_6
timestamp 1731220339
transform 1 0 792 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_534_6
timestamp 1731220339
transform 1 0 776 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_533_6
timestamp 1731220339
transform 1 0 648 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_532_6
timestamp 1731220339
transform 1 0 536 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_531_6
timestamp 1731220339
transform 1 0 568 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_530_6
timestamp 1731220339
transform 1 0 696 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_529_6
timestamp 1731220339
transform 1 0 704 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_528_6
timestamp 1731220339
transform 1 0 544 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_527_6
timestamp 1731220339
transform 1 0 568 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_526_6
timestamp 1731220339
transform 1 0 736 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_525_6
timestamp 1731220339
transform 1 0 752 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_524_6
timestamp 1731220339
transform 1 0 552 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_523_6
timestamp 1731220339
transform 1 0 352 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_522_6
timestamp 1731220339
transform 1 0 160 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_521_6
timestamp 1731220339
transform 1 0 400 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_520_6
timestamp 1731220339
transform 1 0 248 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_519_6
timestamp 1731220339
transform 1 0 128 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_518_6
timestamp 1731220339
transform 1 0 128 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_517_6
timestamp 1731220339
transform 1 0 240 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_516_6
timestamp 1731220339
transform 1 0 392 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_515_6
timestamp 1731220339
transform 1 0 440 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_514_6
timestamp 1731220339
transform 1 0 320 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_513_6
timestamp 1731220339
transform 1 0 200 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_512_6
timestamp 1731220339
transform 1 0 336 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_511_6
timestamp 1731220339
transform 1 0 432 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_510_6
timestamp 1731220339
transform 1 0 432 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_59_6
timestamp 1731220339
transform 1 0 256 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_58_6
timestamp 1731220339
transform 1 0 608 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_57_6
timestamp 1731220339
transform 1 0 536 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_56_6
timestamp 1731220339
transform 1 0 336 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_55_6
timestamp 1731220339
transform 1 0 136 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_54_6
timestamp 1731220339
transform 1 0 128 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_53_6
timestamp 1731220339
transform 1 0 312 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_52_6
timestamp 1731220339
transform 1 0 472 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_51_6
timestamp 1731220339
transform 1 0 288 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_50_6
timestamp 1731220339
transform 1 0 128 0 -1 3332
box 8 5 92 72
<< end >>
