magic
tech sky130l
timestamp 1729042119
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
rect 22 10 27 12
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
rect 29 11 34 12
rect 29 8 30 11
rect 33 8 34 11
rect 29 6 34 8
<< ndc >>
rect 9 7 12 10
rect 16 8 19 11
rect 23 7 26 10
rect 30 8 33 11
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
rect 27 6 29 12
<< pdiffusion >>
rect 8 23 13 34
rect 8 20 9 23
rect 12 20 13 23
rect 8 19 13 20
rect 15 19 20 34
rect 22 27 26 34
rect 22 26 27 27
rect 22 23 23 26
rect 26 23 27 26
rect 22 19 27 23
rect 29 23 34 27
rect 29 20 30 23
rect 33 20 34 23
rect 29 19 34 20
<< pdc >>
rect 9 20 12 23
rect 23 23 26 26
rect 30 20 33 23
<< ptransistor >>
rect 13 19 15 34
rect 20 19 22 34
rect 27 19 29 27
<< polysilicon >>
rect 15 44 22 45
rect 7 41 12 42
rect 7 38 8 41
rect 11 38 12 41
rect 15 41 16 44
rect 19 41 22 44
rect 15 40 22 41
rect 7 37 12 38
rect 7 35 15 37
rect 13 34 15 35
rect 20 34 22 40
rect 27 27 29 29
rect 13 12 15 19
rect 20 12 22 19
rect 27 18 29 19
rect 27 17 42 18
rect 27 16 38 17
rect 27 12 29 16
rect 37 14 38 16
rect 41 14 42 17
rect 37 13 42 14
rect 13 4 15 6
rect 20 4 22 6
rect 27 4 29 6
<< pc >>
rect 8 38 11 41
rect 16 41 19 44
rect 38 14 41 17
<< m1 >>
rect 16 44 20 45
rect 8 41 12 42
rect 11 38 12 41
rect 8 36 12 38
rect 19 41 20 44
rect 16 36 20 41
rect 23 36 28 40
rect 23 26 26 36
rect 9 23 12 24
rect 23 22 26 23
rect 30 23 33 24
rect 9 17 12 20
rect 9 13 12 14
rect 16 17 19 18
rect 16 11 19 14
rect 30 11 33 20
rect 38 17 41 18
rect 38 13 41 14
rect 8 7 9 10
rect 12 7 13 10
rect 16 7 19 8
rect 23 10 26 11
rect 8 4 13 7
rect 23 6 26 7
rect 30 4 36 8
<< m2c >>
rect 9 14 12 17
rect 16 14 19 17
rect 38 14 41 17
rect 9 7 12 10
rect 23 7 26 10
<< m2 >>
rect 8 17 42 18
rect 8 14 9 17
rect 12 14 16 17
rect 19 14 38 17
rect 41 14 42 17
rect 8 13 42 14
rect 8 10 27 11
rect 8 7 9 10
rect 12 7 23 10
rect 26 7 27 10
rect 8 6 27 7
<< labels >>
rlabel pdiffusion 30 20 30 20 3 Y
rlabel ndiffusion 30 7 30 7 3 Y
rlabel polysilicon 28 13 28 13 3 _Y
rlabel polysilicon 28 18 28 18 3 _Y
rlabel ndiffusion 23 7 23 7 3 GND
rlabel pdiffusion 23 20 23 20 3 Vdd
rlabel polysilicon 21 13 21 13 3 A
rlabel polysilicon 21 18 21 18 3 A
rlabel ndiffusion 16 7 16 7 3 _Y
rlabel polysilicon 14 13 14 13 3 B
rlabel polysilicon 14 18 14 18 3 B
rlabel pdiffusion 9 20 9 20 3 _Y
rlabel m1 25 37 25 37 3 Vdd
port 2 e
rlabel m1 9 5 9 5 3 GND
rlabel m2 9 7 9 7 3 GND
rlabel m1 33 5 33 5 3 Y
rlabel m1 17 37 17 37 3 A
rlabel m1 9 37 9 37 3 B
<< end >>
